`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ww1cFCaKpEaygJUT+P6Z2OD0uzJ4IJG8iyHDm5UNlVWbTWS9KXjZ9jEg11wJmlv8lA2AVebHxIas
7nZJsy/GjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gy0/aj7fr+HoqiF2MKC2DdMRffpsNgkz3LCA0LoXsy3oP+ExvEwYs55sO8KAxVdJaUPMOFr+w6Gi
VDRBmTTzMTTD1KvHQEhDppUtYnGyL/2qAWb6xHvmSHDtiAjlHews7qZ26fM0sYgNx48H6LSqgFd4
hai7P1C8/gEiLdaec30=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hi2M/LxF9qgAZzAUuc501Ws9I83yzxDz1ea90Q5QjM7jLsFrH4fLD2d0WWY2wDTdG0Ih+QNnE4S7
Oq9DybBH0zvBRUhAQoExlvdlIfU3Jr1YKpM3lLPQTLIhhCp1eQgIZljQtMN1p0u0HDYYsZO5DBeb
LZHGhmPHPWGqNQ/iLmQ+PQu0B5Cb+1VKyvK7Ipxjf6wKC/NZlztCmWzwV4WC+jY2wHB2IofyzZfo
xRBIRCIpTb+tTiKgZ9oAjPNYVjgXC51YW/c8ZhnzF0gIdh/tD6GDSX/DdrrBN7Oz/gtduYw5jR0b
WsJx7lVGCa/mgRPb2+p2mjuutW8gGGnh6+Yo4A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X16goI57idQ5Yk2jq4rj0BhsplRtdzoYr8oOU2lBTTonp1Nx4fK7AS7KgGuzY4UqvPTHmPTfD5ww
0YcXmh8hr2Hk6aIz+aWFV8C8XcReGDrBhi5Np0Vi5hozuTfEPpWuDV7kTmarku7FYKZbPt+lsAsd
f8+cIo7ySKaxPnzoHbw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RA9GWDJZOdw/NASVbYOgehelK35X4QCDpOGKLkbLHbvCU34C5eqCOlazH25KMTrAHxM2lx7+fAsw
HHb2ZWqK4pB4ww23gPcOsgxVCyXs7Dx/H6E84snPbj5EBFAp1p9GZJoguz0skOVQzCSeso4vwekP
kvLqf3Ypkz4/BbGmeIV5O3MvxWppwuIHCb+NDzDYU2x9uQ7mLUtu7pYCzPfN1FeLiv9ttZaXRuYJ
ADExpcAMpFzH3bwg6Tm6wL+J1DzA4jLGZxI9jxK+L6xNTv2NtONryX7sLla9heWPJCSHR4TT8ow3
t3QklA4V7oRFEhlMh0Nv7QVOAHjukKSZ99LumA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6464)
`protect data_block
2JEuFaTgqghMsv5lmjCzRKFTRu9v2Bd7cfnnEymmK1IpMPqqHVgKVztK8UcvkN/cLu6meLkuW+GH
jEF+IasLsTsQoEbARf7iGoWy/qxr/Wx8iI4qK11niwKvKRzj3E/VIfcoFWMI7lDjskoNrB5ON374
xdQdL472o5haNrGgEzQCs124gMoZrq6ZZftrvXJyyhHqGqmNNfQbG065CYcPsuRjXxzPltG3oMhc
7n7pQE9F5O4ObyVFgYrFINih1IyuB6ga3CPJSEZRwp7Gz0bxN4RD0DBaR3vYvY1rH6jZ2As9bin/
g6/KlClzLL3bvhOho3i5jcTXFPp/oynSuLkHDQ51ZKoe4iiZn+P9Lh5ruWqMMwHt82cgnG4PNvMf
ATePx5qqt4t2SvCid8vOIsQd0vj9ObRA+r3MjtMd1buYDfwqMZz4PxaOcso+DKx3Gnjd9txsAm4T
Ux3rzFwS6J0ycTf9sPOLvni9MYJfYWdnxGP9YLcQBD7yQxZawpIY8aaD/wRcdNh9QMiibnfO0qf1
lRe/UTMU6BZ7EB2OLA64BAIRRtrFpIcWo7XeHjcXGzvo/6qH0a1cvr7RB/rbn0frDOQFpCRpbKV5
XB+TAAEIjE1X+FZTiMpP6XFZ9Ud9hVisNppUv9jiAmSdtEsK+Gf9JU/Pnx9WYBfbKv8DH9eIIKBZ
j6C+jkrjFdmQcd4iyvWlAi6UZGXPatFbo9wfgOGz3sSXBHHoGpBBKrFF/4MsYyRQR8ZNGAggXdXt
5cfnRPE47dTTaeqVaaE1kv+7tk+3OiAdgC6WAXYPJD47PYnnK8647/1mILbV+4Ulf118L1t8pPSf
GLqANMMlQPtk6o/g0dQxl/R/nu0aTKNA4D0+6N64FGPzUJ7HsFczUiEeT8Kq9Ve8YwAdYWpe//l+
Bri1qUDpTm2XY1MJ73mAcQ48d5XiZQo99qftwSRfURMgBUQqRqC8XTvB8LQr+nQ92oZSCkrdMfUV
dJklOfnWavoz2Zy4FHZzDmS1VjCJHPBpPnV3OSiNS+3OPT/J5ySkHkLkt4i8d/FBB3romGtkFMCw
+hyWqr8ijM6I2eJwdt9p6lOHmT8WeHm0vU0lzlq523yWVZXszm8PLRVAEOvkyy7CAxi/iRg7hDg7
vEifTFC+9m9L2cgCvyFsTwerEwlYxDFduSHMtx3R+oLFgTfn9Z763vWrireGJe2/gG5PtXUj6bOB
aBiIFYrOQuHKp+0eRCQLpXxSm+0DeYTG6xSvL3w74LV4oVXhytLUspm4qUUw0aCs+hiCDqk/1xy6
ClHf7lhD4BMZsLK6K99luo6ZV6OEooP2jaHcd2OODLxaAZ8d2lGo6VBo/kZobuGA8Nrw8BGJuVM+
rEPxAo71LXwd1vtaHtbpio3hJZ+GyiSoT7qqdr2Mu8crBTlZG19Rk8y63MWU3l/MImGiTAmm56Af
JA2qfkLA2MF+8gpQuKhnj6OmZ7pwBzaCrrdNlRN6BFNb4+UJuwrSivd+Od6UUptLQTJwbGEZkDWf
ecKoU+GP58PgOy+Ko4vY8QHt3egSOnsC3xXexhVJ98QcrU5adLFyBFYJ0jxRQfHoDAWhjErCD3j8
r3k5uUvqANNJ038YtkgFZexPJ4OU2zQvGQRGhG8t3I58lGrHtGDQVRf94jRDIBzKDZADr9K6DoMs
b/tMPaFJgwY3fbyWQcAGoz/owsxFLEtRF54I+IvK150DIt3R0ir0q+z/VPbTsRGejoCNC3ZrmXn6
z7bJoqqKQ2RGZZZVpw4uWuLwxHOSTUCkz4LyyMhjIRKtardNk+oMQ8ynOrXMJws9uD+MS+4h+6Ul
AmyQrBl1tDIjHdkA63Zw4q8UDqRtKLXDyYMAYn6xQ1GOD143NIi0Ub3vf35oyvilM8NGva5xB8Ed
0tr7qPhJ9VgXKHBTNhW+3QPmdZYP7NryUNQM/ch3s0G/VyfXD9Odw+EUChMN+wAC2cafCrx5pqhE
fIv3qT3wKTg+7RakLGbi+NghQyDyKOVbgyaTHpPlUnBeLHBqCM9htou643/A/6nahNehdCFlH3zC
glSSPlcsrZSNnJqOxtQMvidthVcXXQI/cNgx/bXRvbsa31pvPi975LR7JBMib8YDmlMjaDBb9r53
2CzcicwfknwjvTkdjBCwKVx5PGcOARVoHTqmAehlItmmlkRC2RKdgIY39/jOshgz9ih89/ND9AZM
0vDCBKrQ8LRCIPtIVFJQ4Jpe7dw4QlY/FK0x+KR2Gv2umLrZ3NhbenemV9+zC+XXsZ6BpqMSVP3F
q4CtjrEhAPooJU/xSQlYXYnsjdvNAluSO/USpTziepAZHplXTbIzjSyI4g6hwjKccWrrHhwiqZPg
omT2UyLj278bow5wrP71VWM3b+Ecw32nevJb0BU6zA7ZWIcD06g2OrbpxcAPxXYgo9c8Fm/XCZsN
29wA346i5nks5KjdU4aGD68c0pUCtNm9PCcf1bWu032jBJRXEzjmA1NHqgIZ0EGiZq1aixhv7pJK
x7xXjCFGjb/OqmwXQz2Pp7XAxwtyXCgsKwb/2hHowwgygc4LO1AmaA9RSKxl7nPaZRFiNBSRIN/l
i6EbBrTZVzeQtOv/SWsY4PcRmv8Ia1QN4YSwsaZT3wwWxhvpO8JfKIJIzH7iKYqLxbw5+c4d3UoK
d7uDoEPNwDplKyeR/QCGHwb5CeeqsRA1DpATiqIr1t5X90hmKZI44eWm7QOU/64ow3BSYpeSGfW9
jEq1veQCytKqoN3a547xCydtyWyAtSgISf+B1yL5ecTvfbl4+M47riNXbovtps3Ef5xRij7JR/mF
6aObvpOi8CdqlTmJ+4VwEvXddoibx9kMbn6Bpl8exOwExNyB9rQbKPLkG05MSHqTdwzoyyeeUyr6
C7kTllEvtKKvUtX8mJ9fXElK/4Z3ZX5XROuFg/hUNEsNMOqrNFI1LSTOqR+FspK9sxBBp0uTouWr
EFesso0zeUxozorCiu90+S/AjqcwX0kACxth7kN/rfks20ZspvfZ8gnH+X35k0+E4dMDQvRj7Qma
bf5BEeZHIFqD3yv2S2OX7B+WWEbRiIpLArzJ+N3IrH3FEmzySwofIw8Q2PArdTtcfQBeI9cZsNlK
PKxX8o8bvKN7PSOucFkn5/D7DCiwjnNJxS7mTbAdEhVwyzqQu449yigbItxnuLDHzHypXouV2q5B
ClXQ1IYhTnUK0teWBCq0PCyb5H2AD1shGtwHjzsiD2C6wsKqzw7JSD/plGGHVwRcOgmU3bxhOVoZ
Hd9fboYmMMq099emXRjcZ6OGx4nhMU3waJ/TxahqHosRthIzpSUvf+8dBUxGkck80DzLH43SrUC3
g/e0/UC26SutNE9CdUv+lwUMbSXDyop0cwd51Xqa7MQS57WGUbDpQPIk54VtxS1ig/IOJPQVSewd
9K4lp7Imck80TtjcJgV9bAVW3uTR9/U+4Ymxhmy0birEYdbXNLic59KvrqsHJ71zSgIbGC/4It8D
GhLfq1sHsZKp9LphwfXA9xUV/neFiYxqFKIZhfE0DyNFQKchXtYRm2GYVOcYs/BfS5W4dpORO5rg
wis9Xum/951bmUhv1xivd7/ppDC38N9A3aymgW9YddfYan4O5Vo8rxtl8irVxlr/pinZkP1FgSll
q6p/oyaHIOnF0TMzzWntDb1ZMPAPgBeuyrMnbaZSXRjhTXvdQOr9gipHELNTmIHQnqAPfqVjmBhW
3vEEFew4vrmi8ztQEkttIs8kplSPnNlMDyLeZ5EX5IYAcnfGVbdV8fVDO/t/ycVIhhU28+sua15w
C9YJ5rIIz+mEBJM4dOlLdmNARmsK6gdaJeQlutjXRo5+g5fDNpvW+HjbZvE3rB8MLX/DYg1lwJDe
V6k96WQwlX+Y+jzGrrb7azE1m9cAm0tWu1srtADPqrqUi1/wu2X12KH6+ib1z9hsWdBwbLLNTfXq
P00UTZlA5/epxUsfa+6e0++qD2wsZsONnQiKXgSocjnr1apKgQpaDBPzmvuaWLd8Sje0JBb7xKqw
VmK19GAwetFkLbORDHOfU3Ff2tOXVtuglWcOTlZPWrAAy2/nY9wIL2BMfqwEi1nJnKnefINPm91I
oDHC4vDrTD4EXiedydmRpDY4+gk8VwDc8eEriIWVUn9Hnl/KQ/BTAqcF7fxZ1YnKRTc2qloktVyD
EMPZwsTR7/KfRJVEBu0epOG9VDVBf2f2h3DbKf4ouIfHgqvKlK8y5vpEmjgZD0TWa/k1QD7GNe0V
3TYF8Y3BjvF6VlG2d1apF8bDmtt1umkfO6yPH/9Zce83U5ejd7FHIGJdlvq6QnDKIvC0I4YrmrTB
amGXJw1x9tsTjDflud1cp4yrT4Szhzy0bTZCtrEceg7L2BmzEA3V9lMRIs2j9QjmcTE51rK2Iq1J
W0lhjE6hoRbz9OL/+9sXHMMNf6G+Tj+SH3MdpL4OU/RzBVpqTn3ClyaUIqhKbTYdcnE8Hge56Cjp
zlGD/cuF+pHM7wRu7C0Sw2xTXw2/lpQPTf9WXoVI3ZuHz5xdyXo9bLl7niwfkRqpAavzrsFyFqzh
ClUYHFkj/cTdt2utZtQRbzEVJyTj+6SjuSUCnuqu4H96KOVyuCUBozTA8puImCKV7451rOgBwwaV
ODZP78HHv/BmKKNKpOuFVW8oCthgdH7O+s90jpKDiRr6cylG/ocrHxgv9dDZQUryLEvPrjSqLhzT
7gmcX9JZEGPdcKm0++v1iDX55r0hmxIInA1LgjzPr0s46MPheZIGRLqD8Ky6LjoxLv2GKsrB/92R
WUKctsAoCozzRwMC8FBWEZ7vdsByBqWQs7RgIW0sUW7rSTbFc2UdfPF0DXIhrf8UcsMX0ujOoje0
LnnTr0grng6S706lWLWt51UOVZjQu+1GRMBXq27Q+z9i0f5VK4Gu6IkOwpVRLhNIiDT0WdKU5d3V
4Gacv4pbAkj+YHoj0TACuz7WJEAKNXH9APh239D3EQRdX/vSiDHGDVm8fsDrL9ugLssunqJSICNP
VM7GiFT2ZJwfKVd99qeXAIQLeCRg1ig1G0ITg7oB7S7m68i5m335h2CtiUAceWiIsdys7immL4VO
0RkyJxaCIOk4JiA6dWGHKgLsJPg+LNWMvdl+ZG5dBG1Jxgv3piU97MeE6/HAQkrFUybXi6PjsQBI
4i1b+5vDP3TODubmqbvUxTQwZBPsN9fwOmXUco34QN5GezoNrmFjNJaCJkPxju2ynRNY1KFk/Fpm
jPnCpC+V4tyebluA7ggl1wY8agvtEwOhbZq6xeUHKgGVMW5IUueFds0gXqcBm2D1u+lBkt3FfWF6
FnpPvgPu0/3zMMB32f3gnw7wCq2eiJlU+VTzR0CL09EXG8AuREjWPCu7h9xSQbS3KuPaDXzhjJyh
0aBEJyeNRa/SCIR7xL2x3B3JGp4qMexGNP3a3ysWoaXz9iRuyF8Wgan4TI2KXaZvfe38FWzmVSpq
164vrGTn07Sdx6tI41N8zIclkGC6pYKRq0+sdR2WZdFD/b85IzdkXGyvwFCNcqfEbAIDb8BOA9Jc
CUnVz5rhq8Mh7xHVmOn9Aflfe2nuxG39VVYh7T8fNwxIcFdEgQl29zaE9UDsI56zqkczHFllXufg
BxeXV8c1rUKKyq0mDhWdMVRQqb5dt5jTIp2UiUC2YWeU7W3XNroEBFYfopp/pKmGCbHlForspZf2
hAbnR7BacUSG6LAGMoH997qgAeEPwMrJMzZeBWJp3RpH5A/WT5NEXHGCoi7CVs8fqYi1eZ2Jc5W3
bX4DAFbwjszMy9LgHykQVSIfe3kqIKfoqlPeAbS2eJ1OX2duPer5US2mnuqThQsHXs7FWBxcV6ZH
83+3VMCPkZf0o2uwqSc8qX430eYtPnCUqWfdzb0DL18Do5pETgwj7/TJbSsXipXI6tnYH4v7I6dA
Lxp1/t2ZvVXLGVifSuuY3zwyZ9+AB1HklyZBo4C0gHE5dK0d1GDsE0z7f4ccmC4+FzID+nzO2eub
mn5tHv6zZ2w6+ZnJiRd4rCozjCK5UCSBdoA+rgg67H5SLvDTeYp31HJyqOMVFwWO+AZ/B+gCznS7
AD/ZiNkiYSB9NNxzo7i21LydfovfjGZj5LyHJ8t6d5B5oU0t8/zoiPaC6Lbxe8xyM3d/o9XR4mKK
NYaciNpwiVvqAgu2YawshUhC+hQDF75jbRrpW9gRCNoQobIilNIeal+ymVDeEhrlCOPcccEIXT/2
sza2KfJr7meveTX04PFcKQE5Hgzk2nE5TOfsghY7Ml4v8oeBzmzf440c/p1KbzTYLH9oVxIBW+HO
bqYjXIti/XGtiFQwWWT+tQFYoR0twR3PNkmqYK4nb5sVeVfRwz5+5Xn9CGSel5j1GWus7td2Rpvo
AnbQGTcXkwt0pTEt+0ZWs0s233NrHXenFZjtMilxhFmwXSS56nCE0sQ9wEt94OwniEUkWZHg2n7G
Y8kBGodczsOVIL+5Hqt3jVQeVVdetTQF+8txDRJfGMdMjrigRo3e3/353T8joXz1prZYUuMhr0m1
c78uPHxvQj1ihqemE7Apzr0AEsfZH5ehqlAL0tgjsOpspH363C9XlS+QOE62yIULtdJzTcwEd6Il
DwPRoRV7aohrjxOGVqunBgZUylMmfgTGlM9ef9MPlp69Cl2t6mtmhomSI1u/uvhZU0RTZtxoBuMD
LoNGBfb6sPk/ys6AygZGM/tewdB/Z4Os3VIGZOL3/9No3pAAOia1MyL+CEmW/AqLgoKif2+UdMUT
Dz3g1PnPxJBRjCz+c6CzEjAm7bj9BuM6zc6jejEkvriU5oT7Em6qZenct703XCamUfmHj7AhZk4R
UpZB7AKykoyyxUYuGZBl4ZC9B2IFzkqiAGyJN6Y2grhnKWvow6K8fb4AD+W++UbQR0Z4klt0KUs/
1y+ed6UAEogByttqncKuJnPtSTBNrDn+dzl91CCsrn8F3MkUcC4pG+dKFDg1MwQX3Nbs6qZLpxgY
+/1JIl+JBWgBXuoMhjcdcjhyF369QG4yVBRUrtC/24w+hSWHhJr7TXAMGDBRxyoRPFA/mJ+xif/Y
uABOUBJZqoY7eLW3Q2pKJMSU/01SKcjTWOlQtJBv4W9+Vx8syIznNXaa6nlLBf4tl8hrxUK6sr0t
oGOhG8qz2t6qseUoS5h9XVakRXsrNhuZKLOyuVR9J91/z3BvbgNSbdT2aQMP+QY7XdA+CrT2z2wW
IJUC2n9gjjG56NUUCPsjsRamVdk0WzuuTsIIJjOgXiiBBOMqAiUrQAIK1ppf3yvsqwZmL6sweySW
iq3r4f4dVWfpYMNWDlPhmcBW3TVh65f6Qi+iS1323de9BcOiEfluvuISOsDUBzwqHeF1hU5OSmYW
GBzq9ndzhN99DrwLWU3TtGNLPdhYUYFB/PBY7Sddwbqr+6RWREM03M+mi2rW/bXMwTBEo3gw06s5
4JtdClj8E0Awdd0+8gIY3+W6n/9PIzqiifwRtiCvGA7vRPNl58CI84XTxzbWs4B08Qynf7wyyNlj
n2ctjqQKfo5grJHEFXwvB/at/qwG6oc/nBIVi69rXppz0Of5GnIlfVwl48l1wPsUfXD63At109jA
GH/yH0voPsWyX5VJfCSNkHTmUvUnI6zuKaIrKloEMbXHCEneydFZuSUKSqZO50Z1E5QyrdcFlBlC
mYgZ/2we+Lxz6G9/bmKw0PUQ3ePExBvMhrD5ozMj65sJ3+6SKIRyOIcpdYDkkUfTAHDehly14Tr+
G+r+VHDe+GyG0fZzEIzr+OH7sEW0M1cPu3hPZ9iitEjWw3F3M7B6DMpUAWnhg1ePGHC8YHgeNQxa
I2CvaD3TWX5DoeVYA2TyMprkzorBr58ylAQD/ptvP2NFDH4b5bQ8j5gjTrzh7b5RQyYFumbqLgih
FluDOkDT7s+BEw5QRc/0ebDspLnpIe27O05YpW9EPA+LX4of8nKGTgBO3by8XLsICxqaN3Aish3W
uEsl/UEwHJlUQe4UyO86NA3ix4Bryw4ycou+PcU8twf9AaymoUlmVMsYR9FiHz5xtpRT6MjUZOl4
HUUSeoCkxiAjYNuZ82CvJh3kSbWet3bx1piSAo9Z4j/sPXxbbRJTFwNZZZSTEfhSj4w4rbvi3BFa
ZagqfsJ0ZpqYUc30YldF0OOn/oqMJ4l0WYwaW8pmTAseJWeCF1um1seXtTYowmyPZcspU3DLfjLn
gDWiRWMq4WxcUn7DsDGAdLifgveOCsSG+8fgltwDcPhdnGXe+W5+rEgK48HVgoUTNv7M3mxslxXd
wqLqv8fw2Imt3TA6VCmNB9DSDA9r4SyJQ3GeVB5OGmF+w2cgpmJYki7u5FZLkS3+UIJiR/wGC8Pf
98lqe3QmL6IHiQzddyNYLit4CcUr6IYq59lHBXKHMMdJSOLC6Ylz/bBloJJn41fYDJNE9B2U/aH8
Dx2xatn0o6QXH5xDXbWZbVhUxsKZHuDFXkxOMHeX53O/qOMLy7sbPa32OWFkWO4bB95lgY80PXOO
Y+NKU5aqcMGk6INm5tzp2eam7wBVL9ofLXvVz6aZrSsYj5hd2EY4qCeJDQsTBRxmATVSVTDEOVyC
MxOpY8Uk8mZ6hBOaGPHQff9VBmaXXUM=
`protect end_protected
