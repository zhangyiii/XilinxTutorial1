`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 248960)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbB/zJnlY9bLi0AUFrGn2gHL2x2kzl
0IsX27FVgcMWfMmmyn4xpi+utfLsyFMd1KwCPbWyiNvtW5+NaAS6jRlp6ofWkgavuJbgHqPsHagn
UsC8kYHggKv5Z+4b0sG/2Lq5X21rpdy+8kYgZCpOxfWeFKnsV7oS7W6es/6u2eVsxHaKPsTHqXGX
zhNSizy75qOAWnDYoGOmIKtSuPupx3Hw6mbj+y9FHHbDtRRRCY94jbPBzo64MAig98ndQK4ZmZoT
5Dvy8UNJF15fBXlbCCc+ifpww63QnKK9K5kH2cr44YglyikpueE/uXMuDSVB1Sppm/mCha/w6Jlf
nuRwD3H4tjHdJrApmKUWmHxuFHkY2d6Uu7fdoV0Zy+YYYODtJu8ll9bmgPDyaf4PW6js/HdJNCBr
+QVg6TLiwgFXOJ2oGUisxjIcD/cxb4TcxxsYmIW2j9wefd97hR1LdUkvIejpfa0Fk5SDP50OlKp0
xGE1TR/m5SMgqG2XLjwTCjs99jiBwaiUckbmaNBIfEc4roeLvs34I/P64hFRozUavlwA0nkEoJtb
c+lHi1in+WUEW28uhueQnEw1V9Z0FWQ1nTUWAmQNEiqt/LaUeo7GQEibi03X5ds3LHFfchMTAIX6
EtnuFBUsHI4LkCIQIucsIPj8Uql1C8hoeZmyhbEUdr11GoFn5w2wQSGbFE2A1tpWj/ECzCGSAtTT
pGvQakQFOdp8cCfd61nprEbcYlFPwaqyw3tndLWCkc8fYvjDCLpxeHSU+NYue2ODVLPJXBGsFC2u
maKoPtcss4R4mF4QPxrlh2zQPCItKOUr2YlBHDgNuLEoHHRsYa/mpdag5O/zW09xdwnUBoNtVvXt
URa4tWLotuvOCYSkKYNnaMMShE5fsGRwXAlyKeQGvlKfvcE92ZlY2CN/Cqllr4xPvwgoVC0H7QWs
By9iZhdT6eGQLdWe1rviGN+xJv7dxVqDCTov4MZBz/8UCBxcrNi6LuXz5OcybDl4XDhtTdljMeEB
zn3sriRNk06XBr8rPCj4bNOB0Llz2Omym8DMfygJCR765sRnFhiPZIkprGx+Y4agfZeoUVZxniU+
pd4CqLHdD8d97180zDxPN6W+TDOlVJRlZ1cT21SasxPy/6iOHKAgTYHIOvC6OpIFqsgviqpVeykS
LfzYhXqc64yN5x+YLhIv61t5Xc3KBD8VZypIK9Gx2A49O+XQB+e7VuhQfmq0TE2opE65p9wVryho
vFll5cvFa+tYPkYCOP/DIo0kKyNB5RNK46S+S1mv56ZpUO0cMHvAfWvEB5Bi9SNEPFUCunBfxXcu
ciPcAV/piZcbI/t1FEJh+Ydv/NUEYR88MGzhmP+tQmtKmumdXckIhyOI/kpDmKD7bbipHGbnBV62
1RjcRowtIspabfmCUmGdJjYI4Rd2FCHo/EKpf9yFQ/NC7PUkPI/V4bxAJFLMgSHagYwO3UOT4LJJ
sMYTaSehUqqfj3pYohwhRyMBUrgKiHw2JtbFa0MXbO9euFN+uBqobB++BmuD/DZx0Y1SBpDBr3AG
b4hUwdxIQgaoqUn6yCLfjLLbZAKwT/+Jz7t/k1/5LVsZiL5JHljUS0VPnWIevU2DccPVL0tniaOA
yXOZD097P77OSxgkP/qzyjKpdbgF+Q9zE3+ahQwLPH/9O7xA57c8prD0OYySE1qRZ+avdnHfqEiu
JWunMe38JCRwzvkt4wBAwMQKeHWCnFzmN02QNFzLu3DIHL5OAnVd9rcgh/8Dowz2tS+B7rs/sJiv
ug7QAgYVqJKr0yA/s5hbpyOJgN0dDCzINSK1iRbJ4g99xD6C7apgo6zs6bOBIYcA1rCuhQDeP/C/
MNMtD0j9Zb8y6PsN9tyU3eHFbPBGSaQEjyXP2bA+D0eUCAbTTPpONjXCGS+kFziiz+iB6Gq7sy3n
RUUGgNx/njO4DXHb9e4FQpGTubiPucKXKhaiJ/2h/Ge5H6+fdJUgBGejI+i2+Ef+M4JheYVCViwd
KlFTI9FEoSFcdNbWt1EogAFJHo/EGlxiqpKSLBhPErJRVAFFEyIKVlYoAUPpC57FkhMrOTlKCU+T
zRTxdeWhwwmHyoBDVGyo3ofmXN3lA40JFovj/NeCvg+uz8OhhwC4YzBx0Fjys3eEUar6MQc/Ihqt
M/A5UQfnnOpoO9PfU5ZNYPZqnPlbbuzhBQtcAIoakYTEJCMyo3epKSB3znlg9uU9Kc0BOE4tp3JB
eTuERmGj0kP18CFMblg2j+mUUqNQ2gRuaN9F1XG0VkDPAa7YzMAMR9jTi9hadkYv4FsoFYvNqtj4
lnRM+deJavuw+3nf/o89UaC8ogrVKf7REwwYmlQ0QS4bJPRLEACwSfWkH5NQcUMbOezDBf48NtyC
v7lh0QTfo8FBJqTJBpu1WBp6EFleO3ALye0WtQ+S7oCmsrhgk4GYgzXiWrdnco+3TZV+h59ID3I4
e+lukmxQ0QDGRQJcShoCrekryJKmIlc5UQOPRiI/tODywHXhgMdeAQI3XAF4DzHbqZeX40ru11jQ
ys1cYcNkUp9VaqFuDaVZxWrqkH/Q2X71xW25pf7mZbI4atICSJ4HMbcFY3GlMecR4Vll0sF6XjGq
uJ9eJpsHelXL7M7w3xVD3oQs7CDoypduSPlJi+86+ArF8+cGat2z+loZfLGtSX3ertiCi/DS0Z3/
AIhYqEa8rY6DtjTFwukPtk3/yZiNcfTRqDIMxl453vpZQd2h+yOMHQZ0zIPFcDrB3sDCf/Y45N5p
+iZFCQRyWaGYAizXwOfKyWonRiKHDmn1gKdwJiTCsDlwC6E1YfSO22GDYO0B+BsV7D2sSZly7UrJ
D7xKbHTXuOpDq+JMVOD+W7JZYbKxB2/KKeJcuNGDl8BQv/e9MSH381hoqblwJZbuxRk2NUd3n4Ls
Y84GJyIdV5vTThzEgKM+Rr4zSD012kBMkHurwd/9oxuBS6xHvNEAr67PVBOxouAo0FLDkynIIS2k
Kp8IXpZN89N4n23Em1cC261nyq2NPWa6hDolQUpMZPxfu6OBPmgMxMIEtk8MviPQRArCCHDiG3WZ
6nXDAHYYlX8TYHXh5KeAOtVEdeiKp+bazTYv9De9Ffyp71v/Bf6F3gUPGfUodYNMK+AbHejas84p
4XSgHoZNxxEZ/FVTAoWeWN2jnvf0MQlDlX4EIUCDRTYShvVvd6iZY7kkY/1UvIxM05R94hXaBFv4
MIddPynwu/uUnZwwgizFw4I5VgTWSuPcbJhB53DMehZYMBZse24HS5GBMYDGc8TsqLRA33vtU2ra
EQeHkI2pPVtfmCQkkSglQHvaf4a+Pm3Ui1u/fIUdhGzS3pL0LHpUtWPzdhoEI1YDfvAGtvuqQ0HT
pL14E/07uKVc95sB1p4Ivh6vjDX33e7xP3z6pSFtPeDdAVHlF2c+wUTZwuRtxS4e8ChrzHZgCg1e
gepOcFTS1ajJSfwnvpgxa376TDsBwYDXsjL3kon5SZIJtW862NUeXLbwwZuFuHeffjLCGS0OVqpd
f6iBVGj1IdE71WsG3xjXPnDfC41JoZyGwLF7CtWfwPF8v/svqBm4cW3pfSysNJzSwQBg13ePAiqy
HhVpSqihs4dmrrHgcObXke7kkCnEyHEfZLbKytVPWiUHPYKJmM5LaEfof3VsMeCykT0q/K8WvBfy
PXtCWj2UIz/B9DoEFRWmQv2IzNb4qYf4ASL6g+NORcbUTfkVFCxN9YIX0NgoqaLm225LaB7TDDVM
rKOCPcoh5+FgvkH3/bzsw4ezseZddG5OPnxhOj9032o03jNxH8n+ElA1Ff8bKEnlngjQymman+z1
gTirpy2JisraJoLEe2mwPvraCBO6hr+VyI5dAAaNiGrXCcliCmxjxRi7/vq1NtJX4xz6IrvFk9QF
pIrmwC2V35u5UhFfjYErG4brolLK4itx16USvSjs5fBk8gVF7Uc50JNOjaiqiP6AlMBwp5Qp2FRk
z4n574rvS0DtXg6sFSomZBueqrLh7VaV7a3LF9CNANZle2uuEDTozfhAE+ZHRh1qEJuQcutJgEa5
/eU3Lkui+Azh+XGyWrTK9GQHakNdnklRhONzMoN4C3eTZNHo8PWb3BMoN7wbkJ852r+pHaIFk1VL
3yatkpVN3M8Qwot+Si0c4FPEx8lMiFSWTs06OJOux5jKC1PYXPwuniHFlVOSEuDSaqIjy2tGWpH0
6rrglGPmRVq43I4t14JMYTv1iV6r9JSlRJqoWI0woo5gMRpmLUo3xrl6g84DNv4a6Yf9TcqTqiTU
piK3309W5AS6Sw4oXxRiB4/EGMOwl0s0Wo3k8JD6cx6zU17zrvVHsHkP83JVvb7Kc3eEU3SmnRJd
wAucl3xH40IHFTPttpxcySG8skodBW86PWxnuqPuHRL+rJ956rwz2O/AAhz7vmyEAGSgzBCFSldZ
BeSr5r7J2eYRr0UueI1x0Eexyaql8A/9Zg9IWdh6BiAajtROQcULXhhiutkW8w+SkuPnDVPXxtvH
OdMvQ4Pt1I8rjUsA742aiB9/R8fvj7cB5EuZ0KexRWZBYBfzxiwr3sMp7ejJSQg+f4VUdjpGq312
UJOuN7rgroD7SibeoQG9XFElatV9r9DGvArjVT4lHxLhjT1vcDLj0Guw17zG/kkksTtHSLR126AZ
Cla3mCpfz4nRM0FGBpgTlS7duKcu4l0N72wsxKXO9usD8uyL/uj4f7NrJEAiGivNI40i8kQ7BYhL
KncfjZquZLS68OVEgTZMj1KAXhXqBdqFbNbCV9yKsHDd7W4ijBQ+EuO6092UZ4gJTzICboUBRc4D
MOEy5X0ynkNX9YIz4gDL11UvhgWG+Kb5cerivTdkr0k+G1yRXql0tF6zuRrbcNemcSczypjXQLxg
eDgU/9hZTmB16DpMSTH+N8yImFMbF21NrjYeGOYwo8jSHRkugwYiUdHWsBxtZDZM42AKTJm44wVh
d+TPS3UxBCekSw7+wZTGVOua0X/KC00nf4/RENzLbJBePe3FydY3rq5JQy+ZlpdvLkvdEHhDvm0T
fSXP4CdM34Hncj8yYth7e/HttzmSg8994HlsmaGet3XKchXXOpLTJYq9ILk/WoeVDj6OWLzKtdL2
6YRCI/I+BWKIQivVrLFMBfWG9F2bltR9VSu+1n3shT7wzzZakkgvmVG9raXAMfvyVLzGx9m7oc7n
lczCS6bKziQZwAjBo2jsiNByddI6MV/Y7fKUbV4gdHjsqdGLYjm3N5DkjLrRqh59o2DDKRzDSQLn
r7OMnPAH8aFYUqSINQn/N7fZuO6IxkC3/2U+grw1nKRZZtRefqf/KFpSB9MryIFoSZkz5PnZcjRh
D4eLKtsSQY8OhJUO9P8o2xc4pKrUz4Edp7TBLUNIQm4JDBjg3SqYqwLt4VBvKCCvTovg2k0orlsc
f86RFgBFxBXoQlFEkxXiFihQwQlofb4uQHle1IwLvfJI1iiBMZVHfvzzSp1Xbw9AHPQF9NWyvUWF
XvDrHvUIaXuJ91ucyuX/Ph+cazAfOSvVgzljegzE3TwoEGyFXLDDonfkZ4c6b0GA6h0b5C6Ejm/y
5d6dHLfpOxKmeWBRjMHFbbhlIwL+i4I24OQ4bX1ywy9TZ5g1f+QqNBnA7omJm9cKS6dGIAAwQfkh
hjd2jsP3h/kZmvRrpX3DnyAqzYKrgEgK1k0uIlgQIhWnUdk6R+D0RYdpHOYzcvUv2aO1xLeB0scG
Crr4wcosCynkDsMqyjMu2q8gptoQfVavJ4Du0MYSz9uYkgd+xunSJ4GNJWokEs46tj1j60AotIqZ
7sYj/bzXFDgNplOM263rCeNdpqSV/aog+epj2K3rbzlv0hzd+qkMARbc9S+iFKkHOnYTf8EdGDZK
n8LvGMAi97AlsfxdhL1ESIKoOfIOYfSzFDt+A7QNHrWigBu90CnzNVFqF6lQGibqJBsZowOyy+v1
Ml6MXvWATwFamHE+Pbsp6fK+YW0UZVPKXnH46QRtWdrAkJBYvhEt5yXr2pQT2nr2cvqcrNQm35f2
1GQNbxBEb4eTCJbzOTyqjPMv7BnnS03Aq4XGCZ+4S9MOpvoIso6KblA7wy6r299DgrxcxIZYRujT
mnUW4QDanXWWP7EOAFykOU6UFwEPmD6mu3rvc66hEeQSLvrI2j0WStLR8lSqHuTh9TUa00AZC1x0
KW+956vC3zw3pdR9nhcJxUHZOpun6PBtyMvXRFdAmd9/d5GPzWJxZHR6TrU10xaoX0wdwVFi8W1k
A4UTKCA/XlC7c+0CKOi1kWkMl3GA/kAlZ/CkEXT4XKf+BLxGEXQ1ZooAfJ22z//zdK5cDrFUlUdp
o+yVs/FUqbzm3WuEo5nGpkU1UrQcuME6TRh+VjnYfhbwitkyqcN8AMODwhx8APQKOHJGxdISJqTB
DRoSxFkf1LFul/ybE8WmLoz0YU0MGiNaZ9TADlAYIiMiVvPpvORvwRt/qVB7UOP+gkTE9y6QP79Q
uAIXG/Vn3Iz50/yHiCISPD2uKnv8eQEaTyckcyxgWvMPqmH1+C3+WDT6nCiu1ZDUB87Eumv0xZ0K
9KdD+yV47KMy7oFj3td6kLT5UnTjR6aRCODP+Nca9j/jEBUV8posSyJiGnw4l6SuPyc/BTJwbRB5
p8ljSza0ZkdaMISnUGzco7ILBimnGJ3l0h5pMysgIseh/L4Ii3N6ZGau4gdbeEYuA/57Gt/1ySdV
TU4O/1Lvt3scIyHABgNzmjMfXM866E2m7bbFJWXu4XJNjiO+260Vau0MzMOQ6PBEtSxFXkoAlzRQ
2HA5/CBP/mWl4Bjd9zofEtsSj2j945rcFqpOZ/AKcx7P3yDF2GZmjcP+S9I3rP21YxfBImt49sW2
Fpujdxocnj/Y7Q+W1n4Fb56LyvnT4+/TYIJi0NV7XtRnoyhl9oHtND3ESAUmseHPfIrmu4cz5pOe
+44DsoLbnGtKQCOGpiEEbo9pi2Q/E6qvU9pu44SyYQ/L4U/9HQqtcf3NXqafPnGUCJXObidT/LRp
FPICTNdzAcW2EnLQ99CWB5gKgF2EAcfwc80IPi6F0UxHSI9gRzqqLXCKARTwPjhNB6K5pBnaMh3A
stiEYjr5opV+WOCD8zV9jv6PD82M2rs3ZmaA4aaAiED/lEGkNRbp2ro2yV8ei7xdyFbBCJMpyXjA
bW3tTQRgq3Q7m9fbhPmJRTcCu5393oLV5M/FZ7ghtCkmJ+0jDGiliwzlVj5lKk6xH087cf0KIKsp
HhKKI3YyxSkV7CBFJTCUMeCRG9+EgnGvAbjEe2nbGEtN7irolNKFdE86n09yckbMxJNUL9ptzHEm
XijEc7/l7BtFqdg8cwQr8/OiBq61zUY6vQt9+FN4dfMzcUXA7xwJCkT4BfK22ec8BgHxkJinG08n
dObamNIYoKowfLLLOF77lN0ysAI4mXR0rc/9rWk70ANNkBVwooqINHaUloQZzjZ6H0CiIBogLjll
iR0Rj8dVLDAuqcx6eideq5eKVyiRViPivWh1eOrrnYlVt9b0+fi7kpW6RmsMHMOTbjIdLd2GgQGr
yGTmIaXYZn0j+odb4s81H+Tpk7+JRCRg/2dwBTu3RjP42F2l3IoGv1+vGynFB2WJLm8x47KokYC3
yXZbSnUdAseZzq6eyjb1pa6l+T51iN5zTVgk5IMaPGBmsfkRdHpV6ZaiMru7pBNfcSS7wnFy9T+/
XuWr+rkq/cKr5kSiNccWb3j/Gl34kqrcO1vFNdJWpsLagN6qfoQA1ZOx3bun9WozsWDGOav2aQ7I
DEgZNZLd9700nFxiuEr1cYcuLbnTVvqBW3u2Lmt9nHQ25+ZBOuZ7s5eyK/RkB5gCo9yoBaycN2QD
BdaaIWmR1iwhhAv0IcYn3NlzRH59dysFK8uImAYLWg2rqNtB8WXDcZpLLbs+FJCPlB9a/vy45Ysg
+31cN3LCUbTUlg+DdzCRtwbrYpzSOVEPo32Y7Fu4abM5GyKzGLomsMgir+3Y7ZXpP8ndWtIlSjmX
HXdbEfMZWytdCL+rN8rhhJUi7UrZSKy9h6cSbYbbvJK8TvmYygrrwDtofQYFjGcsH8j16w3mW2I8
OwDu9SwQJaYqxyUGdRoJ92b/sUyC7upsGtCtkjn14KEdJzrQ/QXw5Bi0xa6JWLqpLCqfqi6bpXSY
nqfv1XyR+4lfsQ6uGDynSUPRE/LBFd60BeiJcMS++WLQ6V27ziKS62HJbmt2BYGiRSuVSS4hyZLx
/hUfcAA+H2GLbIPt/pcgppXz/HLKfuX1RHyUwEdL45XUG387hSvEIc61F4UIVJpMTOwoR/CCyGp5
ZCw7RglHDGfJHjd9PsmavBEgsbEd7+JjyJ0ezbaAhnDIGNfiT3fd95klsoOuzXSEX8nZk+/RJlls
KOtJbhuVr5uVVStJ4YWGvKH+Dj8POsdiv3LRGNHO6CZnXu6O7LbzA0vpQ6ESjheILPGG0ZDfnxZ7
bS4AFMdwT3V4ZKEA8qA9MpJJzs480VLYOY2CHun52uRDCMHz5E6dQuuPZ1vOhK6aC5c8XuETbjNU
PZz+vxeBwsOj2cLQWXN9hwUWtdFSjijF9s7DPAuwSe87dI9RERK9SBSx/Jdk4my/pjk/3xuLZWGG
jfBw/0ff0Q4SRnL9++tNhKLiOjHFxhGhLtnsXp605cMW2soHqeC0enJqQQz3/3RBzan4LBtEy9B1
NSkRGUqd0xNoPKOXbI0dkD2XT2C8sYXwEApGsKDiSy3swPFntF0Zdm125341In2DWKTTSRQ6d8kR
jTQYJuL/GKhcJuEWB+ZBR8wreSV/YErMlKojq/3FwWm/hrVN8lcmh+olyUjNRwupKjLeuwipxdGy
xr1yjHVq5mNX0MEMT9SNacDO8iBrBturZa0XXa3aEzcc4iMizK3ACHhVKsB1CwxJeUGAGdF4y6Y6
ouuAlls4IYQizh0CjyLt0mDjWbcd4Fo4WTmRnZtwmNpRX5cP69lUq+CrBW37G9yFYVzjAdq2Wj7N
oSJwRvFLfpMTRHo1/t0ZTk25fFVzy6X/CZfZU0HuD1gjeEnTO9P0LvOWC9k4VRZAMhudGIwsJlpo
2jD34nvJzNjD4LZsCSNP/9yE/AMe0wQOUfZ6XYFBI8HEWERgWF0MXen6PIU8AzQ8gbzCXt9PIYY4
2DpgaQ5o8pQS8adujS73FZEmm1Sp336qzzTM/sS3uKXDQdtGfJ9nE3/xLSBAydcDyabW4n8tGplr
G6+jaFD6wfTK+4ghSJFH5NHsvy/zckzIqs6Mi/IVO5VsQCgGQ/1Gj+QLLTbZI/44lL+Y6O+7FyC7
5DDyS3Wb5zSUXN+rpwfKGVlWgkHs2RlvR/CGnor/HR9OarmSWspuW44pdJzaKZ5DOlUOiRNIuezB
h1si3uwxBSILn7qwVRo8swqvcWVU+GNOV/nEnThgpAGw5y1cYDEfzt1v58Mq298uyDvcUxAg1BYH
xdB9XLg174ngCyclbkCvS8Cb8mBDi7FJWF2dDD1fTHM0iv/7dV4k3TA8/Tt8bhPxQ5iGzxiFx9pv
SKTBum/fP5LIifgOOaVhleGZ6QsxtSkVoHFJRasEJ6hagE1txe4XgZkdiqoTKhaz7nnWECmkUsws
5QiTGdtExhsZw0xuHzxQWvPYmNThPaqlaUeiKBLshXKiWhmjorq8RLLC69kqVgSbar0wKCSMkkdy
eifAQSgO2dNciDZqT/utyE6BgXy2slY7Stfzp9taEvzV+VwQ75F1s2TLhAcrfpKKRbun0IFuqF4E
V4IQWyxyzS3KL+DfX9UiQFK9Osu1djVAadUCW7o3O91d+DoSz2sB1j+25JVhTCiu5scsGgS23CVk
BleU5yZKSzRdEXXDeWOfTNtlj2rZTnJjeesGcIQrXliaK/txccqruQAhYEc748t71/lHzz95qLyJ
S3VNpWK/qaOwxHryPRuzISSFXdbWoi+xTAdzEbtj0SQsH8JXwhNcTxGMDRXpJ1YL+/ew1Muvbyqp
nPTMRWRCcX3xG9IhBZJ5q2Qd9Pk/tk4GvtBmAQlJmWW5P0SV467QfodlJpgQFdnR5TOFyjIpR1M4
dFSjjFlbwc5rAZLFbpI8BLOGakdYgfSFvNPB4SEmR8mSCBaBsZ6CYd1zcY3CekIUD3VrrhhJC9nR
bQ5b7FEpvWO6/n5DU7WNORq6psmOMkAXtXJX82N1G68BO6qRaSR9uK6eoomwy7xuOw3FM8f14CmV
9ciTrW1svFS2ezHJqIF6AZIDva8VNYtpzS9NDXdry8R/nbza+128f5xbAOBQ+LqmZJ1e3qMN6LyO
ZEfawjzRTkOYlp4+0Hqk5LYRpS0+Y/1Az1l1kZlzTARSrgg84etSOJT0ONJaPeUf1PZNKt9NNTKJ
1wsKPanKpiNWfMpbB1UE8DhQRgRIzN8F7FG7If52RiEncEqfIUl+PVybcE1iNVRDpzEYLjhZC+YC
DgiqtOMPViEQ72ZlvGQBt0ccy55MW1nw54l+ENXDW4XHejyNnlyAhIiEI7yoPVNGjGMqKkBLNPHG
RXwsRfKbzQz/wuZKLvSt8hSBTkrr4rB3TbyuHN11Q0AFUzc6XglSvunlLXXNlJG3lj/tFmOD9nC4
1aYQgjGK6Ahn6pOr1N6aUqFL+qCYEXr/ya4ILK866EQp55//1WNtBKpxAFhxm57Cs4ZBCDAAMy2f
zV7DVMxpA/WmfOqoyBEtmw+rSfJuuq4Kf1/cfa87UYJSzwPKo9xiNBGttesZk5Gp/KjJsYB11xWV
YXD+ioUHuRbpPeeD3qySAclkQ9IvzT5OBJRIssJtSbv03pRg/amzSbOuKIlSK/CsEGOmZjK2vQby
QglpDtlg7Q7bMKb9XP/k7BffpQ1kLn3GEJzhCb+auXSE7R8NAYmmvkObZJd8DvjCknTOAEfgoZBp
Mj+JTz7pd7EJNc5HC3V4iSR39ZGgd4VguUB4uP3P/9fp/FoGOKSybL74C7YCXpTVlqj42De7xbnO
d1qusgdK5ZOTGYrQigViv3Yeb+9o9Mn/ppCJRRmhMT2bYDD0k3ruXwtQ/uEjfPzew6gpwOzLMR8N
EV8KdCJgYNINDZES/7WkSy4JmvUheuqS9exUr9XQ7EfKU+IBoRouRc0D2t2AKJyc9/tSNzRm4aHc
d9o17lcHoMo9AFJpOpkVTQrl3lA/PbgTgG9KQgiD3dlBMd00XOdwL8hf9vGSGQfH0twLPSZSKIcm
YaoG6ZofhVyfsnXrOoySWFLzbMtsB8AWUj1zrDv2OGdbXJKP2rnF/BFoVEyR2zbjoN1t8x9UbTyJ
76L95qGt87WxDccIVkmC6H8R6LjBjzxCOa8V/f29jG/jBW0ff1muktMX2uvQq07gnJDoQFVqMA5d
pn7HWPHT87alAnH7siwziHGsq6BmkLLmJTm8jKrt8LhWW2zO0TPTwiirreJ5EGHsCC+sQ7Hysvwb
aI0OfX29eSzJxHoOx0PAigqGbqd/E9H0GWhn242esxxQ6ES83kkPW6HnFX49BkGsACUaBL/0RWrg
FDMLqhzXLKzKAk1B90Xwxpdnrv3om8rSAnP+Z+F5s3cCZ5Z9l6BmP/JswDMBLk7CZeajMIUN8nCT
ZI0BlG8+WzPz4vhKGZRTcVyUyIKMz0HABlOSKlvz2dT49JLurQgZCsFOpw8DzxANEjTWvKEyfmnP
JJ7uXGHdiME1cUuZZk7KlgGdGXj+KHQQ0/d8YdNluy2L5s8OKjSn/C5yNnU5tejnjI5XgWeaYHD+
B2YJ3n5MvJ3eu15bBtWDwiahyPJyKAoYRh7rGbZ9yPX9c6UbMrDXXEMm9a9aMjenU4ejryBiXASm
cObTjJNykYyPLj0iKHsERpP3Qlr3F05BSAOezKg5GMVhDbCD+lHZMooKb1zxAoS5geomk70e+TJT
A4wX1gD74hrYzo4HwNPOtd3+XaLsNU5DV/coYvGShifL20fPFHsEsyW2wIHTAVpasc4RC9bwT8DP
pZD/mzfa2kLCRVQUaC7V5mYGyRYhxjb1gI80J/l2SWz6HBmsTY/UTV46UwozeZws/VUAzYrKcO9M
/JSZad6VeQ5gOuPEMhLWNiB1uow47suMF9C68BTtur0L22aQYzzD7Dk4+VA+UDtcgHvhnBM/7Qtp
AoSFz/E5FxtfYnvWTxBDa/5Pci6CK2FO1pyltCGGeSxVvmKwvsnZAkCcpkcOwrPmsxRKy2Bd+wVA
ONofCqCMzKZ4EierKj0c/HHAuagmwVkMhQbQhLrxULHz3zQd5XIOW2cKhgNO3WXoGUjPvau8E+fY
9/cpvYQKgHejQ/hPpUKbBliqRYfMM6DCi/7p8a3vSIwOeeySuus8JpLcFKt1EZTIivBcyfiNgmwx
IJ8gcSh4Czk8tyCQ1uQhxibwTOefF9b4q+qFO5UhnJSg/RlUqzghpwbtsmjA9kV7gUFDwHc6JT3p
XwjbeVLJrzfMqNZ0BLLA67IfpI/ZPJPMDyhLnV9+ElzcKwwTlE0l67hhTw+Ow39hLphSoQa6Ok2O
n7VY+E7NnYV50o6ehRyRZAzVdeLTzP897cqls6f+DUofWRqQXKwmgYyX6xEUVy92TAeGREgqH3d1
rjyVqzkxUjOc3tWCZojeGeSNeeFAYPUvI0uT0v6c5fMxSoCkvgcIQHzjRRo0VGj88vq7INqaPRSH
I0DGg9M4HgxhBnW28INGUjYO1piikAOf11rZEcvyyhr3djzucGB1smStuaGAUNOgXbI6ZEJhnh/z
FPjE4iD/4b+Z4mflUob/7mnLrtDof1+5o3KgWuW41b/ubcVrYF+ggIEneIExmD2THEMSUpz681x9
rpIpS0m5ix9UNkRoxC+8jXENXUxvDJ9btiplaZD7G4wExHdUmr+v42razhJi1WWE8rZrUSUqWRGw
SboRPf3go8Viqd/sjoOb8ms53ZxoTDPj7vWZ3mqd383LK3eEKz/M1cIqTa/907uRh41Ck2fQ76H7
e7EFeorJ+q5fjAnxjTivsCHkdKWFkjvW9/TbanJlt8FgkxOdJMQwuW038JZxay4kr0ZQ1Rmbf6M8
FAL0Wz+Ok39kXiy9Nl+iB2NSUX0dxjyBXYM/Cw6saIqP7fZfPsABeL+XfcsxvX/R4WsuYPq2YRaI
e4W4I8EPUThUZZVLkKXx6KKZRNcbQ14rYXMEc6/7iNG9OvrtmgwJnEXGfAR19hDcVkOpAztmA5Vn
P+PQdAbF+ioga8dfEFcH+UUV8Ps95yoax4xp1Bpzxje3B09ZBGSwCxco1tp1pZJbhwXII/I+QigS
CwZ0IEvmlqBJuNsZ2of1a9RNcONZBZ9VcCaahaCJnUkGl917S7mlqv87rx2ojeTDNeZdURqF6UKv
tKK56V9Ot5nowrL+W+Nl3Vwgr9HeRZp+TGhrDHTdONJL213cvqlH6ppBF80CX2PwDCRSY74V0G8D
86qqk5ROHEEqXzWASZN2bEb2REwKRgLrVusClw9LOMpZ4nRmq6CvHEngW3lq02Tk3a+OSy102cFE
7obVKxSf2J0Tz/jhiNcYIc4GO/TethZOqM7tsSCeeaJhPsG3ZKnrccmJndZ3ojJZmHrFPKA5Vbrc
XZEfYMrTWDNoa6WWQtY1fK80R+bkjAqiyde7geZ1ngYRfvxknDl1OLQG2itVFdannpNktZqEyRxy
/HdEbU/qT/Pc9f7kaeXvVEVNTv6PmRvXBstIhWWHOQHRRyaWGCC95KSRBktfcjd63IwenGIpa9lm
/JW/Z5FakVIEcjygX8mhT9oVdeEM6DsHqo35YZvH616aAZO7p4Th6TBEvfy1gVJzaSSVX2OonPCX
pRYE3N/imwtGHnB22+24FGVGTuiURbEV+uIyhM8YByOrhu8u4I4eoSJBwAsyM9yLaA8kE42xiGRD
+cynAT+kCjFg6THbyu3VXq9Ir8Cng7NO6i6oSvrosycrJBW+IYGldLoS9NSa1qqOLlt9HPhPYkhc
bNbCeEu2m9bsNby/VHgqWJj1jVB4ZQjRclrldoTaRZskxAKOA+w2RKdUf7ldtynlx8xn9vG8VaFE
bBg3w27BuqSAguTgTmwNFvk7+JMSYXIzShWzn3vJGrBCzCcHIfN5eSig1+buA306AICWPpG3pW2K
Lum7XvHURGlnrnk+/TRAxkKJG5npAfWFAyVPuns4DOJ8QDpxEsGEt3lNeGJpMgBjDFZcYYg1FArs
Xfg7ZpB2hxSYYCPHgMUtk6nDdZyCL1US23VMgH1AAi0zVE6fSRfNRJblz3jFpuNww+lCWCC2nJKg
ggINDPuv/W7fj6zz11cvbNxLHaELSvI6GWKGrpkwjuGlGLF3NtLV5UMj5tC17qB8fiAC1f8ehJ/2
FrE/dXpXDjgkXuPMRNFKuAsPx5D+bSAU74DNbPNibmK6AcsQ+X4+6Qds4cPMzn6tzJOUXP2ELEF2
Zv/uw+6gBDkR9AJxE9vsTF1tcS7mWhCMOb6EU+9RgnVJvn3tWJcpIVRUqwMro3mMBbG54yBJELpi
RVQSEOH70GhutZgyD4EEg2u9lPx8nLQBayM/Ae9hYJ4jfHeIkNqwRysl3lHfrjHLiSLOO/8tbmJt
moRt5ik7kXrFS94VBo9hcHCTMECWWVEiR6+DtBiASjPHuc53OMsk+nR2wakBMoAusTS3BAtlbZDe
D/p9FpdSsNrT321FgJdsbyh7G/FgCgHjKvpXDO2egCB0ZNmPjl6oDAN01jqwovsTQdw7hzGAV+4u
FrbQvUXqYlE0WfDMnqfIbq26sPQuFwab+tcP9Ye6QgFLnX2+S0vQA/urnJH3XjCFXOkjFyIeI8Gw
Mtcs1q8v0/wtnEFywmlqGJ8XFkrwPAcBBvsQ5ctoLun2h9ug/jZsTAPHCEQDX6LMpyJeLAliIQu8
+0A6y82Ez24TaKW/GKgySn3DL3j1zSIqrmtvypl/Z+gDii+fBqsH2Vb7HA2n6lxcyu1H6AkdQUWG
gVt9LLk+kETBi3uXZZtRaQKECX4qdzHWxJ4TSCQmkdhHAIju+EU8dhm9UPhddGlQmhGSZs3l3spe
z/T2+o1/Z3/laZibSus24YqFlU/nu4gr0kGRFdSs6iN8SjX6vpxchOf/y+d5xK1TzZM5yRRZXZM1
qmS4W1uX5IN24kna/n+Fi4XvNL+RnKIEvRP0Ev1sn4nF9EfynwMYBfmQUIpt8l+sx8YCJvtvQugR
z5FAh5XGZteZhInq3UxXAbKD24cDMobizTObH/YrvhnnEp1fUPz1voDkOxuXpzdjl8wW9Vgd6ctO
JE7u2GjjHDPOiDglWFKCdYWAsQGgIXl/t6x+2nSsrw5MkQy5i8WSFvjbRiLyHRXDQXnqsZI09yVw
+8hSVwSPi0ad+XC8kg1Xu4dFlDbs0rCktyDW5BvmYCULUnZZesqgMfTHkJG/S/OnbK/LCVn2oGop
tg9Mc6WocTk8IWirY1DsQ3rrClYM9gNXMRaGLIn+F99Ah/LLTTxsO7D0JB/FtBzq2iX/XnACgwZg
bIqCdZlgQ56slJLV7ihdvnaMMQjh0x6OpKwQNRd5hQUfeMZdZHfBiswecRQZBxNGgss2NHj2nLFv
FI6z/SVIMJ+tr834ziKM81kFSRBzKtD/0E7kzN7vOSS/JeQ9qRiM2+uveuV2vc4vj7AhJnYNAeWW
lBJoT876npNc00//SHvLalGX8/rMaSWOFnNrtlOI9fiw2GRyLgCQSQBJL7STP7BWmu8B4VTHDOtk
9Hwf8yfCAezvdFWDBuTWe4XCX9DCIyCshCrk6jaVhT8+JFTO/2jzYCQ+jv9bs9bb4PkrY+X7XLLW
wWBHnDd8hPS7JLTyy8U8h5op0unZ2GzgBIGlsjtbPcPCrkxSH5xX7+7LFQgwb1qhVf0EIt48Jpn1
kKLAn1X7VHiyYMANpD47MSqZgpslL9nvl+BlnoBm30AeC2xKarups74snD6aidYT7+Kb31S6j/wa
Dj4Nt9hm5w0bboO/uleyO9UuljWNZnajGc2Xqg5cNI8XrrEBX8salfwtQ+bT/HCQWLdn6OMr8qFO
LTKXKEdnOT0h9B+RAEBH/SSPwfwHY08hP4M2FfSqhar/ihC0cw09mVaCHCqFrfKfR+53hTNIpT84
5BWh6F0NfQyTxFWWCrs2oqR5HfWGQvcgF3KrGTsHgrXdaf1sIBDfXCkv3J+liKW3ddmYPirl4pd6
qx5UxEtk0uXH4UbMFlO3CzAiaH6KsU8JequLPh/w7YJStlfzMZ60wQtPE3Mv/vWmRi5jSzxdxA0d
AQVKfQUQrG8tFuAjWI2W6MCgpYGxQ3KhsRjz83/E98K0w8fH960FY5Jt9QaLH+NUCxknHOLiS1JS
+P/rNJoELAVsaUxN2wIeW/kRd/xjbbIlVwjKgmJ1T+GuJaALcJXuUyJ5D/pGruFw0LaM8elEuGQC
THj9kWLK67ExY4fEqnbWb8hWS6QG1cMa4uyNC+3tEHpxcibsJNHbTTlCeUrcbeoNN+hxksptQEUd
HicvMX7PikXsJDhCj2AAQ3RTCS3YYTepbY1JGrW71KcDAML9S8ODUhSnonjnaIcKLQ4QtNKzGFlv
WRvo55t6ZQQhA7vhzIV5va/y9l1ikjeXvAXbzkOcZRosi+7w2G3sY0qQxY1vUWbn+dGmvPpRltjy
Lz/At8V+Mf3z+ujzQQTR8FJui0lsazmf3FCqlMdodj/yrPLJCmyMRdSJ0J0rDT/cKenbqIW5Ezz3
LMvghzzW4uBqmDNaiFaLOBIM62af4v4QW0rps/MHBrLfBk/n6sCVnCMezkDhts20NCiisHnkvR5V
hpW3IStaFZCOvRVoU0zc6nyW9Go8DqN2lvWYNXbNuCxtIFopvoU45cVqV01wS8eeLg8vCqhwryW6
wet1m7JbmdX7TyA3TQ6sGAB/9mRdyiYc/gqXnLfLLY9Ri/uH7moU1Ae1272/xObO8vCkqdNi7Vzb
MA9+AVGeM1+Y4IauALeIEW2J9qbMKfY73vMmgmKqQNjIS4Q3WcXGxDZz5euunhXEqmuRHWjEvSwY
+X86RR5XORpskL/C76b7jrAll+EbfM3IkBsPsm0mnmeL79CXq70AbeBcvI3qCLo2bSX83B+F8Avj
OHoI6v2gbx2wPYorQ9cY/9nbFiZzHcEfY3jouIaV+h/P5dfKjrIsYM2kMsztq6GOOAyklKAW92G/
+iBJIQoepJsfrsDL0Mrk9F67bLRahFqcutnzbEFVbR3pt0KSuWfzAa6VoJKfv+d7tAMkU2d6whB+
fByy/4w4DaGItabnn8NRYZLxORDcQ9IHGHfGDgpAmgmtSQ1aSqU4SFMFlbX9d7NVJI2QP7paHgeu
IgoeRHfiRk7FB3c247d9YtS3ZKALmucHpKwgyTtTY2KNyoxsHI1iWP1Nywjuhle+ocwIjSTKaVx6
5H/hcDDVCPtviYPoeGlVN4zsqj8q5NeCRQ1f5W0iu8nxfdNqj+VbAZ40qFAaFM+0pj5J78CrPBxI
NH5PHeOm22QFvctK6JYMl90wgzoUWukaKbApzLhQXqMoMKIjMprWiIZg+HQHTMuzVh8z0Nji6938
CoPsU39mMM/tetor08OPG7/UtqxDfMdFr7bJn3uPDz1JT0aaLYBtSxkcTHpu+Udjq54tWezMFsyY
Ldel/0UXj42dh0x9lZKHygJKOda7xN0tzf6saYKuQrK7a/x/Ips1PEkUlimtF9NGnYV89VoNatfq
qPRvrgk/MqTWw/kstlFi0KsfbBpQUj7Pqk85Iumhz2++n4g3zrTgNBIqwitIyHzI5v6KdoR92KV8
ZcmI5z93yFui5KBKeo0N1ZAo64mb6VGyKKzbyv5BoBiAX9hnO/UPKlmjCwhMoAlg2d6O/u9LD9QW
ZDt2pVtoBSTODd+CGAbqewCXCX8Qydn35UReCnU3klV4gNpFLaVrFTiN+ABLAprBXbGo0/C+dqol
IwHr/vk5VnAnNaLJDrX+aRsjuLksIuFJhILsc6ndZdJQxcY1xuw9g9VBMx5ia2JiJZ+tlWBqUmT5
R4NVxPbcdxNlip57YLrLC/8MPHY+tWjHBeSYGqv1ilSrZ4hH7cpVRbAtl7cAQwiVDuVsDPgVnQOa
FPebzGzHcccUuMv7wCUhVRELyKDBwY8YShVRyxK/6xPWtaJ2GRuiwvp4+SAqmQAVPR7LIbntsDiZ
LXlZKksT3pdolvVastAdhXz7V2n88aFiGsIvUp0o8+DhXWrbiaHz56msbwwNhv/DCkh7xppIXbJB
SB5HxNUuiqPBsPPkwVo+Zyxpb8+3qdssjZM1QI+kGzgD9ubSRzm5j/mdmu7lXC47QIaoD7btMSni
hQxEfKVhIqsfVIcsU0FF6S++I/n+k2O60i831KPlDTiasVokCdIx91ax2Y+8sTu4l8QZYChWVjtT
ITZWgwBFQoXg6XfX2/4nzOprl+9x8mZaw+VfSzdW0t/k2rzgNkmRo1o8wMuKbT+TdkFc/8jta6tv
dCL4GAduQJUi9mIUEZECQYaPZ2HfEwKroT5LetTLwYFrWuD4B9oH+BoD0xmwekTU4PJ5YXq7/Rz6
Is5yCgt+nyqyDzT6hnwSyc8f59YqJOU94OrnsTVC6sff6KY0hH07/xZWwcJmvuOJF56n7+frlsry
hieqP7pZpB8F9XnxsnTw5TtJ3qO5S5VnpVMlih8YHYOBBgeisClZQ2hnWyp1jiku7/TOUPsrjYqz
mUwfQM0Pgl5gsss71xXUdpRJ/9L5zYNNfOa6isDKpEmQXSE/WsARQo1t0uYx8BNWTYmaBq5eb8bh
wzcb+9+3JwyeE73KhfIJgWezkfG3iENaAZDKxE27HT6FUyusl6l5i2l4t/BVP7k1YcuB+035DW4x
1MRSoy1JHomPyJzPelcTT/c7LTlEZf5HjRA2lRmh17OJ4XRFxaHl7f1S7iHxL7Knejbp8Y/XxlSf
SEDlv61iYuhVXRC1PKFDr1orqnT6qFIJ/FTCu6r7OBax2EOymsYsX5QD4D832Mqb0i4y2ESxQCvX
pm6r8EGP/kPhBjhHylSsLvyD8sjDt/KXDZNWYCYRc1sp6k5Do5qM6p6gWEoBoQARyzpZteSUqYri
IYQk56+Xf616PHPsD/Z5k+x8IZLXvcp7HTdpwxgTnhgPyr5m0TuQ26zHptdqDeDSqAkFWgu7oMvf
Pmd93LYoULtiq/e/8OHAQ/xqxzKskHOFMPQm5XsHYJ0ZEQlcbK0jUZH7wZRN0IDqCKQq4Kz3ZxHD
DTTsLFTlRO7X4psO9IlHj6RKqYehJ0Z/KCXO+OfwT1Jry7xQQ1Nr9t4iB8gzLvjGhFSmzX5Xp6Xp
1T4Eksbfs714+Pm0kgMmZfH7+0eVb/KkRYsWcqeK9E1HPFqTGx4oRHi0AEz1QBM98zmUcgSOqkFC
3G77rU/M9bwP9s8dEViyWPbew6S8RymmbYhshy8hHZM2BS5WrsZL1xdPGv9+5DOMRX4wU+uRXqOD
G2sFKpHzcogi/moWmT73Ra3osYS33/tXjdloxZbuVkSf1hf5SNYA8qRyqgglrFWkJZ3Yb5jxKd0V
XRYvpqYZ1buAIzXoVo/UznQJSJHaHN5tUVnBxthw33x0vIv4EcPf0Vr1SNMoEOADwX5aBEcGOOeq
dbIWiSG1SAOeqJt9rUKyNGotcv76ADieJ/wcGSEqiiqdoW4yQhAF+tGr0ZmE0iHk/65wfJYHpkDS
YcUpJFAIa2E7dTBPD2LB8kuy3Jqk8Zs8/s40jQxMuSHDQSqFhN80cuU2ER7H1MzRtQZffXiWSs2s
zDQa2UKzWzm8sw9Yli56TZhW9RjLtSBan5g9TLT8116YQoBU9MXDIhVKltF8S1zjxI7l02COWu/h
OLdw9SpFn7ykLLxH20b2VwPtgDWe0YmWufXvCllqVSw4QETOOuC+Faviazxuh71pld4KbSmIvSjs
yqjmb04zG0dByOV5aLHC5M4Bhs25Y1hv99sMQq5tbnCSDV3Ea2G8rcu0p54REaC1aF2GEYnGcJau
eKJFeW/2ztbEBaE/R5I3PwP9hM4NnPvPJ1jX+xs7T9HhYIWu3ZCfSldxGGRDQ894F93PyRhr2x5k
0D6P/KW3rzVMaFERIFkjrSOn9sFkD/lKvu43d0qe5ML/b7KqMJOSMH10jZeBNxLbJ+MeOmIwzKgB
jN+IngK3DTNmly4Wyip2c9dfd8F6XV2Sc/oSz4WV9CAuwlGHAVHwRAbmxnDoJ4GbvWLNwzYWWfuk
mvacRvHYp0JE0SYvL061UMMah4uYDg0xWDka88fPQuv1Mg7JOhlfne/gPx3w0f112FLadO93TNWD
v1M2oJIcapFYB28XUMQ6OI9a3/4DDNRW7kbv+HzuSW+sT9huo9naJ5ZpFDonIrNn6caaY5hQfmSV
ihNGhkmG1smKx4Hn9GWkrX0WCw6BkHcPkwLrcGZVTuxUJZs7CBgXoWV7P4ZD7KXsn8jw+kU8OlyI
CyXmpEVDbVc9NVT893y7NJwSh0MBFJ/XJ8+yNBR19/wdXY8kiO/koAhbTeNjh+a26PIX+hAKItL7
9Z+mUhPq0g6lHLhzGGreH4u3ygsJp5nV/Q/Z2nxRNo0Cjsr5PUcFebz74beiklP+zEAkFwA6l3ex
eWnXgAc4lGrrA5hc1B+gA3zxbNrqSdFL8ds/+fTC/Y37V76rv31GO68v7pPZ84zhN7TSiwRshuOC
9X5IaynaYteoe1bSQ2yZgwDcjHKpB6yj0zIWfpAE1yNTw81rt5nhexPK4cY5zTxiHgeNwpzIvAcj
DsmgWvM28xJvajgV7C+xYlBnjxbST3krX8HuApPC9GpBspBEBueo9GMwGwuOhdfx1k/ux02BfBxr
2FF6PppKFL6nWMnE7qf2hd8YkY6a5EEIZT9CnyZsh7RGT//V3sH1+fY2/MV0KkBioKKZxYjECRdP
Cb1A6hLuML6M/MO0PR+O6jlx0mwEiC8xYm1XcBwtQmCKX9yT7TOCBVKk1Gxas63FzalCuVkjJ9Zu
hnmNrVOY4rC948TbXasmO+GUCLXGaF1bVhoumInMLCmi7FYFtcyupzKA2x/VwuEvoivpvqG01OCb
SccegQCXbbTDc7oxQDGdTtxcQ4Lo6WiCM+DVgjyVyKxduKWhrAdbu8odMnnHjNsGH/Qnc8PpJKBc
BO2pykBjSGoRJLNSHqOLg41/ehX1COZV9mQEFpYh0C9wlr95i1tTGWxBRiuSAe9zX6wUPdrgsTzx
8N3w+Fzy3UYQyeD8BVcPf6VO7mmQfm1MtnzLxp4er/T0LTbFvhOvxpdtbPV85ZQkYw7IobahzcSb
NN+6otylEZ1fcxir9V2alsp2C2WbS4fFu1hqzqKyh0IjOEqXo6U4IRyLEG8vZdaZBWu3gdvL1Aja
nzZBmkSSP84W4ULbYGBoziMhzaLGhCQEFjNpo5bMZAXxqrvTryO6E8/0wY5HjQygVyKpR1Ms6hPt
aS1fB5ba0B9Q5pxzdV4r/W8EAW1pcgNVN4cnrrzWtZbhtWVug+7x16S4tl+CpVKQICeOXMl2AiQI
b0E6eop95ve0nBqWeJZSbLGZOtYvJNwZ75limspl7ohCGIPi0NMnUWFmsH/k8MPf5kHz5dy7wxtA
avpsli0G0VsNSjGetZC6qe61/mPT4ImPaw+fOoTXkjALwv2y5pJ6HBZuDxV1pIyn1ztCVjronb97
yN5P79Y0untbSWfEltxUvfo3lwtSXiIEkyho+R4jSa1XX7+XO/ru5HVdh9Gri4pLk7SxzBd+vZRD
DOCPT0DG/CvSq7yLzhQ5OC05X0B4dXJZvIermLQo4kG7eOF+Eo2cKd8ugRbBQfyItWaYKv/SjfD+
2ItHGuiQ7kKElQuU4+nWtLXmSEgaHf1Aj72zLX/K1LiZq2pKYBbJMwob+Pccn23GsG6RiG4iI1v5
j9y5TehYVPJRGsxqVKdpN+xhkmL13dQWU+QVtu3syoT4S9L/dusZTUn1V3s83SdKTpqF1Mv6tE56
OkXclC/rG0lLji8mETBVvEqcQ4lhcMluirMC8Njj4kiKPQu/i3dhZNDfwBF7q1u4pIonda3AJxDr
fU/t5EFmue+JwL2eLyD+gYkw+L+N49+b7b3RlMpJXpme+e8aZ9wBxjGPjSXUCFMU9i6exmNmaLNs
3Y25xG6yWxSdg2Fh60Z6q1q0+XShUpAzQFHJI1/RfLchzPpSwWJ96GoSL5nZC63jA1j4R5QUUpiN
t5QyxeZkTCIGB7bzbXVh4oyNpf68hYFfJNpaunieibAoilpfY+Du/ICK9NcKsIKfaoER8BdvNJCu
bC9+UO4Vw1PHLimkg1vQm+mw8SH1K0HUfyK3R8cx1FmaDpPfE33XwZwHzOFRxwQDL4PSTh3kuAGZ
D7WDgJHJVLr2GDvQcFqa/ToCYtnN0jSqWE/acgjnIGzCIEh9F/LBPwxU4+FU16QUJKI1XGBbkERp
HQ02iCrw99FU/RX0SDL2Dc2vuw54Hs6ccb2MNwhJ2d3iEiMUmE9/KWJ9Wc4SUECuLxwDZbmeecIK
BXsPAl68ZdkagQeoo6VlSpXaZAQaxmzDyDu1tbwHciCmrW69Vw6hHtLkTPtLWjFj2gw1x3E7fZAJ
JSSBqVEQVT6Rvu9t1kCupgx8d+jxXGb6+EVPpftpd6J8O4FnLGmTIspU4g3BcKuP1HGt5BxciHo4
VT1PGNaT/cT87m0S21G0P7CS50OIdbaNptrNrfxwz9nSVuLiq/FT/lgjKFvjuJ94lhQxwNyHd31P
zRk7AGCQNNqTemJH3skQ3EjjT8SFveAb5F85dyVy+htMeYVPBBhWBxcvjKM6f1BWBWbACqNe2zLc
PTNTa3cQqlEeL+mLoYiKz56L1kgZKngcyg9V5c0pBTccnMG+TUUOdiBqv2ffjF3xnUgJ+97LlOCY
anytsfMWFxNc9sQMj/it5ygY28k/cgWO7uhcZ6XPdPcIepHwYj8iHFRQOKC7gm8HCSWWG++G6QyE
GXwRKMB1tqa6UE4Thajx7PlLVn3hOFbcgBbtPgvKtYZ6/ldrUGqrhNc8asd9VWEexPQku/yJbRqT
RpNgh913vxSHKX9uJ9l2lqCKWxE6wLnLAn/20bTrDPM1XQnb8SQKR7SkEIHQOyaRf1cvjyHRQvii
fiYxwz7o84jqTndaVCv1ZvIS0qIFrO5KqIQ6T8P3scFjm20YkylEI0CCbilT4pP7pOhUCgDfgdVn
3TRtQZAQJs3HlC7k2qTBid+k4/c2rias790F2L5tJ8nOW42y4lfPKf9Sh/iWh6yi82OWaXf0LAd+
5pbU6Y74LxJFQt8teNQN8CXXfkqvWoCjAjnQPYVILRHPbbBy2hHKpn/TRCLi1hJ02BEya6pNo1Mt
1YJ/I0ICYKRNrVm4vYZkux7So0txpL2wUT4xg5XEGp3lcZE5SaPMt3FG2s0tn51iuJlmrSRh9bro
3g7aG69ZqeO1yHTnyzCHCIq5mgPe8MZzIX9fMK1jjEmL11i9mL1HF/rrm4pVB6Xy0IlEXXdKMmhl
gsrk5+YhMJiwMWmY4FJF3v4rAGLno0wtM/3KuABfF0MQQBgzNbsEuXVaQZtZ5woOUd6gsxMwzOiX
MWXL2TBeoxUehzdfvhN30BGlQiXWPLL6jkrzmc8j1ktxRiJ5I5+IG4lTLumqDJYpDNwtZhsaVJ0E
TTIUNLlC5OXF4aXc7GS3C7pOexILgq1tmlAs+e3GdY/wfBf5G3O38vSC9Urwcn3+OAbckhLO0XP9
DnQGtmuSGzWr2nBJjourqpp4qGtrCd3X77E6YE+ufdpazZVzjfjoBg0WGN0lNrSTtklCWw/L8rM+
FS9nYh77dLP9bTx7gSJ2ECBEH+ZG8lSN3EqC8hwLcmfS4dfNYXTZCM00/cWidXEJeOhyQ2obb6qx
mUBpbdbNaZj2RZ+ZHq0O0WzpGJsCy+s0PSjORG0dOyUjwIFACfkvwQUtTjbmbLYSX2ETdwYkNCL/
sPx3n8eiHXkjLhBGZvKa958FqDSs1MTUFMg14OduCTK3BXBvKBOUfl2tYIRERK8T/d1Wgdgj/4Er
WuPuYUVK5cERWbyTmyalYz6POX3IfKhAeaK92k+FViFxM5gjSff8ymI3FgwFuSepw6hIdBdLPyCa
tetFFlzofhBMvtuKBaHy+JbJZcPEwSTGFFNsS4VTyI/u/eJ5/Vpq9E7Fz3LgmsZC3dgbC/tKv3Z0
bV7WLLbQkziWzp8FaVIIJjqRb3A0RKHcf9GgmEArmZSVdBc9YR7WyDujqvIRknH+yDvI8omMNQ9C
FsszK/id9MQh16cNE6mJjJXJYEbe1TzyGzIBCjX7EobHy783luIiORDEoYlsXZxzoG0J+DyYOkMn
Pvfq8eW0/Ym8iVUXgSGx9BvsVMZ+JYM29FdjKLJznOvtPTPd6laOIS2okXgsVJ+tqcc88CSs5et2
ZQGTQb/FIFT1lEL9Uj+KBU8wqirVmdN/sp2FDkyM9paeNiOxILpUPR7rjXwuL8KkdvgJwNI/vClt
sRkV9dSZE/0Xs3203b1lnpsttS2ISMY5gWRs0BcNKyhuI8FNdoqJwsLP4zl3Th7Nof8RnzXzUoLU
5z8XKBuML3RMLnNL+AaGcdAi/0mSj0d+JNyxaMU2oOlzjyAprIWcgHVsg324rSCv1xMlUzuUB6kZ
e4beFigwp2bNV1aLSSKxku54oKgxjBWHR3u6bU74IiaLlWlSF5UxCEU5gD4AKsXaGl6DY4duBW8r
f0pk/Sdf3ML9MaFIslKP25llkoV5verR5BCQ3kdCJve2ko1rk8XZZayxrdXwQ3ApinnqgIp3935t
rhtgw7rWWy57uvhq5WK0wbwb1e0TFzeSeaIZuz0QQPCN5ix3kEYypI8gUArCAA+4x7Il1ptKXamH
2w4xdvdaovltLJOEobBMwchVST8JoHf7SOAl0CgN8NKoIAIjsNUZoP5yE+VJidBOU7fNtz4/hgBi
QDc8FYgbDhRjMl+lRAJ+q8WvvUlUjnSR9VluPY5Zz64bfIc9HsAJ1WtDvzkhpuqwgYTK8M7nzVi8
zUFJRZfdqzKRuT1rznPrsNm+IGjqiCvsjQymW5807G7lHRKOI5BdrwcHtv4JmqjbcC1Bnd0Riytt
htvwzAegXtgJ6bGhBMgEAYNt0AU1/AK2htcIWiuiouyVwxe3XZlj3m+9Zbl73eybqwqfOBLX/fTI
5TgMS268TMCLqojdkiLyQmD2tRb5/uxj8wfAWvKJOkC0vNHliGojK7GTLkSuVzagNYG7J9x5Zpqs
TtjxK8d67KgkBv4RE0wj+udo2tHhM0Nage+/FGKjllSAfSaaDYxMqJ1JDOnivjcal5QNcazyCAeX
4iYlOePnPUBePdqY85o7adEF3erDA05XGVd4AazTue17LzEq/N1cKB4T3C1tbNzhe90hvKYO4Kl3
OtXMchfoAP7VGk5GXi1W5UmE3bIYehEPAW6BIbV6jlqlGYm73yzieuhNgqmcX35Zq1CokY8MjDuC
G5TOibzrqW40gYcLqGczdAGbgoKFdqkMM9Kx5Azg90LVDI7gTWxH/yj3L0CrqjIxTWJbL7XCHf0M
aczSkff/5ekCSRXBn8/3YsJq8jvk2W6efeJ0v6YXdev2jFoueKNfIkwIwtl+J7856lBpV9x2JutP
Mip1LhzGJyoodsJDmK2mm1BYBkhYu3dHf18zbqebJ1s8HpCsueEsc0RhxOCD7+GBQj6lD+zZ1XAo
ClqIPYz7SDNCjP5z+rav4koig8sdWWwhu7r0JQm7M7Sxe9gdETs3r0wc+AD8zU7rKPsU9R2gRHGQ
l6Ivd6I6QEO3+5yxiwYn5O1nWw8ZORGLiUXf3fk2Gkwqe3iw9WrQEzTZWQKUv3W7j3hni/14Klqu
k1ZX8CdOzOGW9zwVe4fW2cw/hlRyqtoXroe6CSNAzVQOqzGQ8REojAFhdOmfmqBlv8RUohHt9TTb
gzaa8TSXIpqZxcKINsEmhC3EQVX51EtXkp2ALX2OU9O1y3MovkG6d0slmQto8Rpa3GVKbXIppZoJ
xPLHFHaVOQpZhMStAkyW80N+TVVOlCAjpMp/yskifIuT9mBoM3QPAFanraRSHf8eGwD3ck9O/TN+
kMcuCh20npfqJDp0EaVpboLQrJeqfLvJ8UIzgxe/+Fp49I/MrZ6La5TcadvPyMrw9f55MMYLnyH3
50zfG6IpQof6MG/mfcLQsY7a00p6d8p5TQuSAukDglJmvEU7Uu1GKlF9SluvDaRT4bBemtsyeKwr
RAQRt1eoFOdl40VyGFyOCG2mZnTX5pNwM6sP6G1pUI5IPzX5zN2qxipcKTMX5kmVXpQO28PsCwlj
NcLzRL158WkI4SFAz3lcBm7hDP25ym7uIYGrxG9Wm4p1t4NNLu7VLQfrs9XfV/UpHMGE18Y/CEOH
JdJLR8ysQgKoXuiLrLSRqkRJfeNOwTSHLcOlTKwUYeUpW/1PNNCrR9+DVkTi6sOnWQrDAXmZe/nN
6bHEe8GEUFfVc2yggS802HlnAiUI8F/7Zo6zel5jYBohRY/HjUiEC3bqsatp4WClnjYZR7CZulFJ
tvbi/fv/4dQcCwNR5tY17k1MKuP8ZBytF2VYv+yxARemRtG4DjRnznle4mpAwyOXGKmLYMsz4ar8
Rcuji34hyO3TqrlTNpADGxrjEuw3auEu9CUlx1hth78jG+Ukr9yWmhfMZ08czwJ6r/+TIm176mso
kIyXcvYu9MivgZsH6ILV2H1crJHJ+qYonCRz2A4l3NO2dJEOtgAZFgXF5Kf9QoWrpIkqsCnfC4U3
m2c306VMfAFpxQN9C/+sepHdrwUIr1U8OTS7K5w1uFhdYOn8uZHScRlbgTgohN9aZPjmyDEx5StC
mpPIOV6lUlqrdoUKuaQt+1nLlerRkqI2sk2RUN1pmBEQz2lNtfsPd/06hGLIN0R0TRPj7/1hKm7q
DnVCI65oTYprwysF4/uouYNeZ9MPgJmMTyJF0VMDbI6ltQ8eSOacYN76vvcCJS4jCFt3X4Gmqtz4
dofp1H9bPm6wfu3HZCbN6m7WWRjjgh6/AXU1W4LTGK0rOch1vVzmsYEkxwz0LY4mGj9xWnwCQ35N
rcq4QxZ7pk/mZS+dyTDd3JlbwkxitP2xHTQ8k7k6NY4drAhE4BLQX4Az4haMgoYDPI14+Q7KUbqa
tTHbBOMq2EeeNlJeL36jj8cpY7cmE7B0D47+XRRYg1lU/9hWn2RGOouPgeE2pY9VIV9s2JC5RjJp
EKh2WbeictaJqzdbnu9p5MGhs2Eb4260zEEPm0T3Ncr0X2HzdCIXMaG/rC+b8DMxoGL+vT2X4vCy
kManzaFs0xKUNwdwxUiFUS/Hd4UbzjfVh1pL1aaTLmDGoAQzMhyt5ZY++jfJTN92d0/56AopOCuJ
BsZQIhFbbVJqRcUBcX/dUTu3HS8ZWbwhZITL3kTe5V0yl4ON6CBTExMFEHFMFh9yKkR63qQolG3E
x28jJ9wI214ENyUoeFbTfL3B8igp1f6XZcnC+8oZOMmGnK8ndxP64obhcjXl6GP1825cuTqTnfj9
Te5E3vA1l0dNmy4ABafTRSk+70TxpdqwLpdbMdSbm8mA0GaeifB/8wCJd9aJhdRQ3ZuNn6/3Tt4T
9SuPgRvcQBu8TMhq6aQew7rtoI+mMqghtgAPsEKx2OYHqHdJSwC26j8gbG0K1sK8TBJH/hr+/Kow
xXobmA4JYr0z/OAoF+rdjY7usnDdqZkyS2RC7JsEUSraa3U9RHqMMZGUTbHeNbw+ni1iJ1O/pPWF
zhaHe8hfFM+lATSMi8AOvdTv6ion9rIbmXN6pZolMLKobWRM/5h3UYP7E2vmRTO/E1AcN0tJyIs3
SHwDluSimUOkmis+qcJc+jtN5kf8E6/L7cWQtvf3ILmfdBVWBDx+DFFGZ6uGdkRCk1Eo87Qqkik2
NesxNgfAp5McXpiDEDRQngPcW0W3arYgC5TG4IPJSdszX94H0Nizcatm4Dltb2QsL5/PXv2tEjc6
bNERpvVzkRLexEy5n1MtUJrd8k68l/4JFRVBsBqA2KYqiWMdqxqQmTZOWOPPBobRp3KwBvDzl49v
IHHGSThYMBcPYtJwZVXMtH+qFIV+eWF4VJ3kj9VE7rt2JubPhP1DV49CVin4LeW7vV/WMuM+x/xM
iHWp9UbP7uW9KtNojRkpzjEjWF3bzuld0xqOis71RyK7dInoiiPB4wrwX4u94OP1gSy5NHYOKow2
Nd7UrQsp/jEtvl0h2FAJiJzSbR5Jy/euXC7jy5WAoZCR/TvaHaRODv+rcLNLmJBPHjKuyHBYiapB
X26F+7pH4q5BLmyqYX1FW9zHRx5ezt7PjFeJF06Xlk5EMsTCn4hD4IVM7gByTItm5Q28MFTMSZRK
U6ke5IYefrbTYtQvhB825TjMq1fx8JnFujgXthLO1vi1EWTIIxF3w0flniUR8ubuJofFKZ2ilBYO
SSgLER6Qzmmt9HptMLeQtOFACAhI4Bcf8CZ3uorYd3xsL8Phl6kglEsKe3BLu0a6nJp54zFkvCmC
kvp1TwNd31nogBJR8knxmkO0h/Jusk/B3bbpED5li0s/M42xWgB2q6bg9z46xf45Hk3f6Fla00M6
e52cHlOfbt/JkjHy7DiSAzzoW3GQUkR0cS2B7qns725CtTlMGJyxvF/utypVVXC3hMDU5OEZ81/l
EDG5Cef6B+dhVcGWLxQf0hnOko0T6sLGhOYYk8rm5B0Qi4u0u/4a0sxqbxStGJ5+RFsilMjF7fwF
kO0BeUb/Ne+41lzJpstvnIDZCJCVA3L53WXJaChvLKBUyAN+hsRBiXE6K6E5M7zOGL2zlYcmc4nL
Qpx+OfDd61tkOp7++CzUatDEoKYv+6xhKOM208Q1nJHP/iU3zBraciF4vAhftkpL3+fwhpCZUgoT
AfHkJhvUjUYTWKb0y7yGNoJW3KM82eV1GX86GMauqTMY1tkgsiJVUoG3ytigsR98f+tsvFqlguh5
bIvLbYnBA2qp+tdMn09LlHbSplo/5NgmNLsw02+ZwdPNBA3c21kdNwEGgrrAv6RPI/ANTGjeuzIW
xAezbqhxicJVEEFtpGM3H7P1m7sx8b77ksLDs2dK4uIU8I++wNGKhV82LFneJ6x1rQjayuzit0mj
veJnHN2ESb3CHMNw31kzO8M7p8NUIaueENL/inOscw6Gxqn8XK7GQg8+sLObbMmVhpnnD8koZzVE
gl7bdYTEN8lVD9tLJXCsRtlYrpln1qJ73J7GKUBOzZUwmb3Z0aofkXRJmTGw1lez5INf0iTKYvbP
c+b0xQpq/pB4bA74CbEuHam3uSGrhqJZ/E7YHteEr48ZfLsLUsxxDxuLmUbxfuBMs7Ym6a0sJsB7
b8AyZtb07nyl2s4UKbc1PBsnzLiQ5xyx85fNiUrJvDGZfI55XRtgCn6apDVF+guIKGZbRxmsyU6Y
k9DGMAeu6dwp9zk22nIDjuAg3zb/HBM0JtHPeJR2VsY3W3uFGvrmOC1Pm/Ak8ZDPCN3+RjYeVraG
CB/t2/H0/rodhrpBokR3ltKJsLmKx2+AjneiWuyK94Yyipg1WwNJ8wdLfx6IEKD2wWbTpDV62jFn
jgDO3fwYkJ4Hzv5MQ9G1z/Gyv8eVl1WtrRgm0YDOOkrtT+EloHOW1MEqJSJdU3h3N09y5W101iUg
ZUw4jxx9DYbo5DFFoB/JbW7xv2ypWWdDKcGnbdyNkZvPfGiA6io2tP4zNmr9Qx8FnieA/gYwMUyA
mF+OpkYuXAJS2ity4sjvAKsKhDGC1JCYvgsvVi3zGRF6H+oiYR91/nEhOjYbsGH3L6Rf2pu2KlOs
nE426+qAIp0Y7ZKgJkKl0YIzheiDykXWuZM8dVvtWqqs7TsN00mZhofBLjtG42iD1FiMc4Nsi/Ve
pYgzNh9rMUI9Mb/1OAOx1OWbdrSmytwajNI/LvHtvA2b0JTVpHL4X99dHYq9Qcg9QSG67w+9fP/h
eakCfUh/0ZJqIoOfcFGVF+DdWlOgeMDKP2sAi8OCHno17IOBcs3/LgpfTe7OlvErlShoGILuv66X
nwZi8zdvnuhYbXZgFB7JCi/qqwbEofrEz+kixCOrWN0uwnWED4xucdI2YIu9wavK5oVy2dWWuKrk
Hb6YeIY57Yp4U1ocymkw6Iiv/BWfB3Mz+zFAab3+29HMtLfv6Ojx73LuiHFhtAJj98spQUb8X9hj
/0xH53v+XiV07Qgbh9lTH4cM9yBM88YlprL33aOP5PiEHJPKEho6E/1IrpYQ6QBqaKf5ulImOAn6
+AursqhEwMe8Xa2OVano8XaOdEJm+rzrZn71yW3FM+OiQaoAYjbDDNlS9m7n5DuShUc876uzneLE
1ASjcnKJuxY9zzhWMx15hjEGscBvJeLU4pwhqlubBUAq1zX0h6sQn75lD1f6s+1zJNXQ63+2GF2N
g4lfK0/PRfC+FqokH+pRLVpTH5Emi7Alwj9fyy019Gg0KStb9HWBzb4eCXGnu8geyQxLIu0ztZro
j40UjgusmhvK0BQj0Ob2+TgWyGkEjlMhRqxje0Yn2JYwFIHHdQgu3bQ++qPvsi1JMK1Y3oNeDn/r
zNVgrtzYfnuQNCy6f7ScmmTqhK1bB+PrfH6GWGvsXyeKWijwK9bMqZ33gqvx8rohdhnTmKWLZwT1
NtFejUFLfNQgK2TvcBriLX2bBF7AsobQVDWqTorb0P1mO1gFvptqhb0zyV0au3T8b/OUBQMfp2+J
hu3joIvNSX+szh8CsVU0nQhpeziec94/N7LeALcvdbFuQOUh8I09KhGzc4z4WG3NzGxies3+ngwR
voknMx/ccDHmIQUA63WPKRgh1pMleiie/AoFJRsy1UTOOQTNxNS6cS+nYhhyEkCdyt+QLnBqsIgo
ktTw/3sNpBcCRxXbio5Niu0VdKbKuIFNKCNx9e/cGSp+vA2TNnipNP+1GBMDr2EUba/EkEzCWvLR
GxUYvplEOaZySyQoRxuu982Z4MJ8pvEty+LfzmRi1dOEGsvMc4+bibDOkNIbUfnzVmXISX9lMHhA
vLuvb8wEe7iKyRC29TUcnzGRyuCep3opiDv0R0SsXw6QBBOgrtXbqCvekN3+kM1FjlnN646ZTl/k
5dACPoRSWkCXBdaP8J4844qth7C1E9vJMJsNHSvj6mIx0AWg4/YPb0V1UvIqcK6Qa23yIMfm3YB/
syDrs4iaRjinYv1S8QwqjPDHP7VQRUVv5xEi37zQkXusr3KTrPYC7kMY0T+jR0z0XR3HW+BL/lir
9V5BWJTrxvfBGwIpYldE1ZLt4TrwGnxLm/RIkVijQGQl+P7dSwaYG+Nz4vXS/0K+QXTGhpE+XV/j
dsxBLXFY0NVziF8G1zNduoaIe1ralOhvw6eSPdOIFsQYHVfyZI5ESA3uVUBSmlaKdfAKpSBuK6pG
MlBsFwHNUNVmumx8g5a7KfUfTk6Sb0K2VGgBOcAoaeXJkFippC/BFDc5UsIUKER3WBX2l9b1wou1
NWglvwwn3+ewK275Cke/JrdEV5imVKKlLdWQbNTAdOFw5YOJjNolzrwZoDf5RpWNSRsuAR88v7cy
BMkh1aPuk84oDX7oOWQTgpx3r9GL4Ah2UiR9F4e4RdvHnd21F+6a3M0nn0uxPa9SOtqfVLtO7hB4
D+A8FEC5fZFKmiqtHkn0V7ets44IQmjmMtNV9lssKdicxC0swSdbwpj4A41UFtWnP3onxzi4D5DN
M5OAO7tWS44m5EW8e2blszOqx1XOax3cCNCJVaXWOHq13u5h9Ke2IMM1kBlSC6V5K1JOWc1pCW3B
8J5ECLLj9a94Zfff7Zn0U1dpjQrSIylmVGday/ftmfGf71pJu3nLJ6i66pBp57enCWQZR4uHLWAm
dQPIMLESV9dJmMk1F769kPCbJzmu6GX+rcZIdMo0p/Fgo9M2J2Yc0j34lv8onJN8LNSD/DB7vqk8
df8Q1Voxd5yQgHPRW7lhxeUum9cX3OSNqo4TyOb0QhJA2KnZmKdGxzj7fnx4LPa3s+IbUtNpJaOd
OJ1sJFiSF6tYIaplwo0FXXc8jKyPViNtepfiWlcbWMO95DGPOGpAxlN94+sIMSu4B+pPhQ3ffMI6
jNmhqtNeniPSwYktlcijOMRGef9BHfFsl3OK+/TZq58acn6qyqO8DgqlfoXnCeDH25E+tE5qhBRO
/FifxrOlAKvTJwzkgOhiPXEIxdAebucS7inkuZWh8dMECyufcNKNx8wvfFyhI5TYUoOLsO7ylGGQ
pZuLj4kmzkpPwYiFAYCvnNTkC1QHa+qjsYlKSqNkgGtCoHf7AuWhaITKTGs/lfz31Yuk0S3D+0ga
rbSN/+BGKirubs/KUva1KZbewKTYgy4B1Cb1TF3sGEMHdcRxzARiCiu0z46HB8TItkV9k+KTcrrK
UD4ttH28X1owzESDIG7L0WB55LSRNv7lwTC4PQVdnxRCBhQ1WMpaI3+UOwvcCkdScr65UrX3q7hg
n4pqYdFeaCUJ9TC5XkTUfkGgUUdTGNq9TnV6AzezBKs1Mxai5S4O3nTu5LNOE0Eu8lwXWkOrcbmj
V4DtMK1Mlm/zKWGiPaa9MTPDS/ptho1sZrf+d8z4XPLX+fWf10AxDAn9CmQJ8doV38dl62edotUY
/Mec2oQvtPaJXUgFg5xUS2NuXVx79mB8QPPC3dP7KV1zqfkm3qStZD1cT6c0iKvHt/HKZgMiqIQK
EoDxLrAdcfx1KFu32y14LuMhay0GSO8Yy1L6ocQU1+MZPhCiQesF/cH7OgK7HKAaRixvASRqapJX
NGQMWfdvR3VFOf+ffMr7ThTARsMTwc0+mdxklMRCIO05Q8sVfkEqiectCq33wquikh8K61RMHTcP
BWi5U7grRJwYsBm1TqTVPizQZIYO5/NdYdCAXJTrPP+Rf5q89t3ZTCS4OWHPgNJjlnC82n/wCW3o
J6NnLVkx5bfmryVj1D0zXonzznzV+hmzzUSzdNqVhhbb552LlCDZ+0+TQbRLS0RhDgiAkkBU+ge0
yic+8zQzvZEqpCRBESGlRByeKTUWwSJyn7Rx8MCiAdfwe704MPrg3kecYZHy/d/yqPjM1v3INFx0
2kQI49MciEjl+UIYkG7XFOeIslZfG81J/24ANis5VXFlaLb5qyFK+eGd/2EOOC3SVTZyiGaMY++B
2fnlJJH+TepBWUyjYNfyPTrLOX0nFm24GH7myndkMjbh1FkTUkvMh6Yy48vd2fTG4u7/RPsMCAaf
cMA4AWQTdxhh83jKgPb+iJYYEQ4sE2DFzL6ribm5HblLDYKx5eiSxCpCn6V6NcIkxj9m63+Pf3RJ
uAsWf+ShNOa5OBiA8JxvGcxBIxSGY2K3XRDPhIliOaPYx9jBlEPff+UnWc81E5waFgBsY1zDlh7b
zHP2xpZgpUn+Yx7g80l6U1pdjZkENBjKGOsE+XmV+iQu7v5FmologdvosxMWibCHJxPylxzoDMKr
CqxBmGjlKfXwjlNq9ZJPPyP6xP/Kc9FUWtpym3PCAgm/0uGyhp0i/nukoxXobo+hQ3KM/L7rOFNz
GcWYu0ys3xJURUhDXpSxtffFDN130YZCguM8inDfW+BwBi3fJGo5oowdv8G57ahytWwc09R91ONd
DVBQ70iuZvDDYeAJrATvhegoL934wY/IO8P587YE1wbJtRWGXaUF+7RGgdP0i0rGbVhIkSqus4J3
ePVS/l1IInF6kE+H9HQiz0VeZB2eQmWbybiJVHTp+hnuzcHYYXaSZHcAqQ2rvhxffyL07FZz6B4j
VtavW//qfZaq/T6ahOH1CM8DKZplKrTYp2Ixqj45/G3LAS103uzk6DxVj0/46vg8e76hHlQxy0hv
XkiQssIPiTywyJkwykKbGF8WHmDU+v7Ho6LPJdri1kaZEMtIaHMdGLUsLhLcMNyUPLK+TO4b8GKB
0I6E4b7bzoZD28dRIWu/E8jtmeJywMBQrZdXplxowi6jQsHMWAAaLTNmoPYDfP67QrYE11+ETXwB
jJZkN6se+kwJGs5ltswyIZBVSloK5R1vTjpIAtoE0gBsrCuNiyIihCAOBVLGa76OoRBHlnVkcifS
SV5TYKcGF37i7JAKkAczZro/P6pPoLH4IYEv7PJ0DOm9cO/dgwpnJdZKOxvgRvLe/ctCUJ2eIayo
GoJynHvBsRly/aATC+WI92HyiQ4jWqszirR6O2A/5k7ditnL/g+e5w16cQ6XLgyzwsJigsBdemRZ
hLLZ3shnrXKcO7PgHoVFuNae1OxbTPf8Zt1HByG/IdlqDB0ZKzhgzltcAdbo8RMBMW1ln/uOe6Oa
j9597WhjqanGZAp++vamN1nEVyoen6jM5fdH74kjkLNKDbXJAqL5u7X/naBrNMKCfuutLme8OlcI
NkUhju6VABaxv+8G0URKdSHAM+B6fBdRiC3iMCpu+2V3vOhE2n0SA2gNRFDdvmcx+jLW96d14Xkb
mCtSqXBMLmBUI7HNY68Kajx3M6GLBQ3Hn88rYPSqEfRE3Rva9aaAgXfNx+mVMW499Uy0mkTMBdc3
3Qc7nHf+3S9hKOS80Sf6KgOPxHFc/smtzG0oCxQvIg2pbiCeyciNxgt1s65FB6uqQhdE6YHr8r14
QB6rG3U90zhkZQ9xkYZp/i5py/k3AHL7ypjXsT+kpfCgLtlkSd8KzDiovi5orFQwHJzSigiP7Xrm
3iNzmsULWX8RUwpAIZpAz2R7IXa/ccaVA2VL6kyxUeR9j2C39Lf6qAPlsv6w1llcPTJp8gNZ8o6J
GfDI3ZYLTQUqpQhIc7OVLjorIJSyvmJGF8yntz7hZWRBxo7WQ1Dm1B1AdqQNNFiXKm+U7LZ8NZBP
7qtdyfH8QL7fuDON2Q/MyjvWiqEHK9ra20kC+7um0uH6rPT2CvaNH6TfQe3tfyJpv/Et8oM0Ssej
yP9/zvEmnu0g1K81HueldH4flfpArNQFyt2YQlVr7j/ACsImm6+rAi2rvPsCluJg0Z67k61b27v9
1yUENspFO1ADeyYY0byoDhMFXdO9Evp7CK+yDAU20jjjTLxGArTT0gHFu1smOXWivmA3w73r3XP7
y5X1gvStInw1n4CJ2uFniYxzxMMsxy/FCVeD39IvbwZjK4A3FQ/pTa0/azu9kVMnCnFCTtEzpw3M
eF8jAAF7DPhR4DeUc9MPXbGMHVT4dhFIiV8bwuTh+pnjhNY+3iYfgyBHo5f2c1mFSAb4Mw9nv/B6
cB0nyRQtv1KTpC3LDR7vSn5O9v7ltd8fytPaCdL3cx0y17dh6pq/r5cYbwY71XfiVunwM1c0/aHb
C1tYAiVeZnr/WsvZFBt19jmpFiq7BZhCyooE71KRKR7+kHJl8ZL+1LZjyvsgfcDkHYe+M9COKE6V
nkBV+aIk3/95yzmTm+nVP34UttsQSekKNfaTsYbkDnlwMYFI3p+Gaczhqp1FcrCfAgRrbzz/iq86
k5mh+k2zh9RldKmRYGpFvPFGb0d5wBsLpJvzFx/gtK2qO0LCCxveU/t3gES+khYrlMBtltcMfjlg
pAizPrD5nnNFytl3GcQBVc0qYN3LOO2Cl/Y0fKX3dMUxps0uT5B4KTfv922hT3Mso3fKBaDa32Dl
oxUPc++D3EBgRXREcyTlK/ZKi3a/0U9GcXlBj5oKVdEWGyzezE53NMmQZHsmaEDqjrNiqArW6joX
BHjP+GBr0eZ4wdT5PDEcG7fM4yLQ1ADiJTXwgYYXYlwXG2Scn/hiyjKiD2N10w2V3QBci5X/8ww3
CVcaZATe2G+00gtwb4iqEJ3Hd7LVRL2QhXeUlYsWQlRLU6RyNMxo89t7B4LBlIOREC4uTtutdgYL
EkYTiLTGkwNhiEXilYmIb35KZViZNKjbdQqcZBcu+fgM3hx/GTc/auB4nfLETaH43mKAmoyxR/Ng
zZM7SH0flvHnJxYekpxDRFFtqcOa73YdYRH08O1UjeNb4yKRw9vbclGMdSDKuQQdg3MtFDxqXcOP
NT5DGZyEUwtye6C8ZSzXDvOCUuFYy5ZLLQC/0zK+Z40d7qFG6XDQvgrlu/gMWTxfI8y1RAmK/szf
m9SvOMqPAEXQhOOSwlwNvzT/dBr4ZLu5A96ES2EbwBuNM1JU/p4B1xS079lvOnq3PQc2tN++ztn9
TqI7qmR7z5bfXeYpPd2qSQViyfxDAhrQ4kFCAxXy+Hdbm2rMNHxeiCOxJeQdW+k9Q9uZO6pB2FMb
cKLzNvS3wka2fttmqRcOjdp9v2kPo5lTjwqymXHBj+kTrve3qdhmVF9kaNBz/LjBGZ+Z5IaHUTuM
9HEHmQr9VjaIgljL/NaonDLLCrW+8JFEIVPQRGH32jXL89raqBQNTaub0TupH4/OJU3+4r6e/kza
VyteJ+IOnuVQkr/Yd/DHOkIXnyNkSyqYxyfutGBO7rYtAGm/sO7nupPWw39riQwhh4UxOGlVYThv
/ycnOI7p4WuoKPnia5kdy16WHlf/LeCIagHHDpVchIv/xvEONiBdxtk+xYffhP++roEi8pmCdDTg
X6qoRTkvMdNcNxb5JbQWDVnXUUjhB7JYjVSSoTl9aNea8G2SregkixxsFWWJ3zFNQ8r9m5rmyEPl
HyxjIDz5QeTwLO2mn57wbGL1yy+0QrHtB6eFI6GH9ICkSDTCrpG7i7J1dI5btitC5P4p9pEHjRuL
f4g2IcMFmJf7PJg0cgGVx78xNsA8Q9YMKi2lQRIX7wvslyIyg6WsWl8M7g7kg9EEPJahRv1ywMTV
bON7ZiL4u8CnxpLUInr0zvAybxJFbnLfxDTu2WEida+965UB29yZ/pH42nDs2NF9CFVWT0vGcXtT
9X4542954qlCDdagtCRrLjH8kZW9jiv6DlzZznbEMZtiCxiQ+ZtXXi1N/xhRODUcpgScyha4Icjo
+5JF8M8VNKs/gTrBZAzNxqoFfXJgWgwLIcFWGN3BJsN7CrC3LJkk8qIZ8zB+4rA0YZJhGJkTIGUp
NSAGbe9BNg4++sZyAYPuTNiE50UmC3JGxzeAj7m9s4hL8GJFNzrp0ex+F6iY1cfrQDJ2r3KgH6aL
Ut6OeW//GB9ClIkTf6ma9pC/0BVYigWiqvls9BGcDW7WLy6KD9tf183211EJkPU6zlagCEtCvz+9
9pRZ2WZaK5E5wkHU/eCoayvOda4bvIanMb3cOFX3sjqz8961Bts50CxBJRxp3um47zCFlUV9UokJ
oGx5OfKZTPthPE9y2Nhf4LVxeWYccBtnGzDhz2DD2JFrznBEYYeo2OeB0/xvRNOFxeNOfL7FLvt7
aan0rNmPZVYVqg1ORwacCBuQg7g5KDMsgYajb+m+pa5+qi/0Qr+fBRCAq1D/91QrdXnKCDHwAXLM
J9CTkcwbccnTdlp9RNZXS/U0aWlWMhmG37Fo0bY7ZCQ80GGi7xmPooKPbBv0Gj3fpmyO5QfZ8z5S
1CiqXT+la4EeKoDwX+sJRC66vahiyxQGzGsfrfTrvWXiz9PUBIkwIHWtQdjtcKmiPEUq/U7PFk3G
BmVJGNc/GKUfI2uh+tO/UDtaHUd6Sph5a5+KqYBAiyD/jCy/CihecYuWQ3ZhFWW0AJBNxwc6zjXg
YRuRo3V/4f9xlGzVb6NZJW0xZpHokTrcbDPefXN2bhvOP/Obo1NHa80yCn0lV2VDwxqZvHP4ftBN
D+ruceLDzqpvTwTcdJ4WWYOCoIf81caFT1M8X8r4SxOkILO/4tTosnQRcGpd24duWNNV0jR1S8Ml
a6btNW8DsHWsL+9PzVq0I+ikP1A5RN5DJ43SVw95Xoak/bod10uIu/JHun5G733oLEdw4vAxLlXo
Ly+NyQcFwX/r8Ai9cC/jGpgKuTk+zYoXttWcGb5/R6tmhMbEpYSrXnBTZONeo6WybfOSh40t1Lpp
8iIJxRP7kw3wHdssVsgH0awW8fYPsWGcUzifkbrquUvhu+hKLHODPT6y2y6Nww2COjFXAuB2uIcj
ewFGLGg+CTNsr3a0Z8P+voN6/9WKWszq03GoSbscBPlMkMEt0EPX8m26BXzxOIs2L97xPZOddom0
IGVPUqZEX1kjYizMDthbwhLRJF39w0+KTNurAnd43JLBz55ib0rS8+UDPJndGmCsad5eahAhK9JZ
J/EgTo2luOApAIOCICQojk/vN7/uQ8EMNKYycqqyIRTMfSzpO1C8pQp8V7ISNTX2ZEGXnBLoZNGc
qVbZesn+uol0nrCrLLxusfoF97/9Z7yBku5gBHl3cN5adMX+hJFxMycU/XhEZZZq30MY4h9thVR3
crvi3ZdDagVYavDe2KiT5Kt+dVJWZEl9+wHARVIaIbvpUfbj/JpQ7wVhLeE8Qt8jK+FtclzCeU2H
rmxcke/xi4KSIwmy7lj9WDt4fwgB5nWkdXkJ0i/38UF2qndO1AIj+ghp4tr7X3YC/L3BdkHiyJi4
J8iJ0d5RLXiec2mrgsjF8D3zC74+cShBSW8mF85LU3AFjnc2enlWCCZaOVImxZp2p66Dae7UNk5L
7V96y0Zte3djOKhjcgFg9bYcRENHENn3neuym+Ud2q+W7x9mD7EdvBRagejtoN4xAhsIsXBKe1WV
lUSQVR6f0A7pzfqqsbKuK8Epl0i6PbSfF1uV9upFx+dIVv1eVBmozJ22roTfyvsvyVRo+QKKQZED
4ISgntmnK1gSjf6MJ+hFqOuVV0szuwqzcDb+9x8mKkYlcOKgOAilhU+PTP2B1VQMKOV03kv4H4bT
JERRamcRrqEUzqlweAc+M0vzjFvf5ShDXiMDbCQFFCjFIxRhqM9h08rT7iBxgvtO6nhSCowj8ieJ
3S2t4x7uZ+JsB9e+1pKWVncpeo9H4JZhKz90OQtmB3Si4waWc0M33Uo2E5Q7Cnd3eUnAUguDPi7H
cBH+5sCJE4rMggt7FfYm90ofdyB9uPkkoRkIU4DLEIvwuIzi5LdxNF+UtWlx6wVy4oE0bNnHyJXy
YxZLZGZ/GTb7fjMSwfBsTXuGKWlom2zVsFzSMCo8FNtFc9rCWu74EeIyB8obMRbNZox3sjc0Xo4f
MO9A/Se28I3EJ+jRj0BQMmhqr2fidWRAsYG/qRN+3057gQhXBCIlo1Nq908NRpIRdHXpNSX9Bbls
7uZPV1MVvjgPn9mII7PEoQPGojTLB/fzOUexdp5M1OafoKgK8drr/U6imE1cA7rYKtWX9Kavixpx
sgVq3GYNYalplKYtGwCubbipyGiAd3tczksVxcLYmcw1MGI5GKIGU5351GKpBS9klN77A0F/8Jl6
IOw7ejQiRKqaJLCvI8gZKzWbbO1YajWniU6ULz/sDtUjxonr/NplBGzzyFCDIIJpDIKfw/Z6eI5D
+jkw4b8Ga4eEFIcKS2ZWggMCFMaU38RN2kevMHxhe7gil5XaZ0H0A1PXas8WZMP4U///NIh+Ckag
yNWck0KIxNAuhE05S+3qT2PCIJeAbFQUP2q5czcrt2XkwgEYYPmiSLhwgs6HVVJOlSsR2oWcZtSI
j4DBxVjnSA7a1skCyBR5x9b/zDSGIzMKSIlwMuBBbDJ4jEVGbRNmf2DHeuXkhl5+08OCXMbt5ADS
YeQRh/2B4RrEDXS0jG1q0a42DkGLBEHt3wqvoAaCQUHFjNLOkQhrzBCntMibVcnI+BPGpBSs4x7z
RNEOV4XJ/oSygYKidYNqZdw6imm41nz1cebVLr7tZUqhKAUIC0Kz9dJ5AI3T54E+ilFaTdIIu/Fn
jsfiO2kXUkM/68RYE1wiZy5fyOrGOZL5ddhgtuqMvICfFrqO93qqtODyvD+JBYCnXw+4xXlDOg4A
oBBh7lrNxpQ7WIwh2PeU6WIru+4NuNBANPfHUaC5u8hiUmrnC94rSYi2xPe4vRzR9bgJa1h83sfq
FJzDyoTVjxsYHre7froz2YuQaRVh9xD8zudlLYHZpOgW9bZ9cu72CfDCCMYozgbve8mkoDN1zFSN
4LtAH12NESd0LcEr3Gf62ffWynsVE9Gsc2rK2vs8z5IUUVqi/9Jc0RP7Uxhm3Sr46lXFXl7D3DdY
Sn1PMnlxsXyfESmQ0KgfQWasjfr0WexcDA/RQ+AWBoDiL29ItJrEwsTL55GYAUiZVTeMJAbB9NFv
Yb1aXK3f2cpxjrgMrex9o0uqNLJnNIfKUDAF4fpK/N4sdXhvm8Og3RodsFtGFpO8SapBqzcJ7bFi
gXZpmH4ADRq4Gj7ZQZjHJeGBzJfTiqu5+WHO66pfw+pTznOu5Izkz/ehsbwUtp1E8f3RoKO0KvzW
TKauTH62n/wXkEFoUKYd+HzFdUvO7Vhn3WLJPo5j2b6PCHW2aoThvj8UnKpJgxgZCZPyY96La0qr
iB8fXXGo9jWb1HKW/jXpm4KpGg/ynKwUjOvpoqc1MBgBQ10+rC9cK2vrXknlL4DBTdZShOmd/rUu
ZGFduurulw9LPc+pBFOo2ZEir0vvRbb2ni8retagmuvIKXp4i+9eDSXhlxyZqugDcF14gcWM9Vmn
FiK2Oq/y9b4iPpqeR7XKusil7z7L1ldPAue3z+O5EGK00rX6kz3G/eYP0/LuYrKQmuzmSHZorXsH
u9vxH1wAgBdFW/IdA8nWDWKpCojgZUfV9jN9EwQUJyf5UyakzLSG48B1j2DWZ0h0s84jPt/CvZUg
+k51KX1YGGOmmxf1ZXvrsBYFla/oVqK+bpD74p7xEvQHfWQkSUy2sUuV5atUilZdarEyDC1i9FCJ
Vlm8Rs30qJkmyuTItKsrCAP8mFs1V7vMj5S9TbIVs/wNwIBGmuTpDgJ6pOoHxSZv+6fzMizApdW1
XGIEPWcecrmN2UReo9X8jkmCqD2B9eWXLTpAVFkjryuaiUpaLQJKR0ehbtHvul1WjQ4qDQirS4AJ
zWoiPWhv4ZQ80zthlZOudAn5G4Hw7yYS2ols1fIVdu40J/JI3zlRIUQB4jHYcrQVj5bRaZjRSI8r
4aYJHgp74YPFREJBdby4SLOOWD91jiT42kIwtQpdQnVwU7AzVPJXogcoUXUcgVyizv2aEH9FqViT
ZT0WlTxh14a5nQPrY4qM1rcXTzYxYiVbSMnswSr/+z2gY1kDgIHPYiKaiboCFo5hCziwLhXv0H57
bUxVMbnkAJUZXFfZ46LU/SqWr8HoGEfPvRsV+6Y+bbQZKFqriwUunfDHG130zEW8aAK8NfH+Gx7j
CsgQYlJxZYU6/XuOD4G0/+TT3C8oPazkLyvt/4vkx6qWToTb66aGYLvgWjjDP9Dp2wgqqQM6HUyb
qRpivU8y3Mr40JiCj4M4WSbYdOZDScd2eu6XngAORL2z1wNrzMtMlsVL1HElydMuNijx9SaH0ai8
RkaPcU10n1ET1Bsj9853+Jf7krzzqxayP3MCTaR5KjIWMcG8bMZzXoeszSXbazK6u4qof7Gw2bPN
scY2b5qly0MmEfYpNIQiQtq2GwpHkHkO7OX0RbEMrR+AWDq1Nnz4XzMVRfwXmlC0fnytaFfeQm6f
zhYWDfy2ZwhjH8JOX7rjlTHgYl4OOQIoO+Sme5E6QuHZwJYhoDk3DNllsO2wwUnERJYbu6j0wcQE
d8wQO/wkBIuf4fsPmEkawkYVi/y9BwT8KSxl/8Qs0auDP89qjfwbDAfUvI2V6tJPwIKFYV8dvtNs
qnP4N+z9QSBOuWnx76Djj4MmVIi4dhME1mr4ZNnVMJroHxeZUDb8I5dA0KKFzbdxttjRqnDjTyKW
QJT0pTk0CxFK4jdlk9b1Cb5mscQbVSemjltLNo+D8cvOE+icL98LvWoVrSEr6pOiXgnfGkG+Sydi
izn8vyCZXC2/fyD6iL2cANBTKgkO6SXP9+PsLgGf4GMbzkZdRRzoQOaqts4iTDPfNLGu9wwuEmQh
gV+S3nnbWlEZR1hqb7+E6T8VwGSxl5Pzn6AkCfuwND2uWa9tn+9kBgcMZ7ML5rWXzZuGGgmw+kWQ
vt8VxJ17godswZWXtrW3loSvIDGqCRDbN6SIAWAA7xjs803WgrI3yjO7OVKlVVboHhGFSbwuOhbQ
somD3i42PCo9nPyU6Qx55R/HzmTQ87KW7QQ8CEzruI54IJCzLqkSDhSW6vc8kbr4922Cj9000XCV
CAhC2fST+1STarnGDKUXfT4AnCQ0QnD2KUkWqj1cX2LC8g27AtQW6Y0h4BLBfNaej90A2fF7ZkhL
nKF0qZrrtjoFDrFLLcOqMntmihgB46QsNUzSmRXeXPvMvmuSCMRYplkCbtDhfYF0TegM2/TZ9GyU
ToE399VZGphounHgaT4BKQrh3Bx4VdeoxuD9OvAT10ROl9LtB/ORB719SOWfO5WAJAyoUBxvlrhe
6ckG8WqeJUv2n6ZnSausFuoMZOki0SEW+4/E+8JJOUtm21hSyAoXqt0RgCpzCaCVRH1CQruS/Jxi
FkAFQJxgra2U/EzjfazSZpSfqKhEiC7pT8xEJmFDPZBn0KV+HvSLZaeUPzbsnRZNg5LbyAXoz+kN
B9XR0pZf8ZyI3W/XigwKQsgG6ssdThz2VYfBa2YsuMsVVeijjQuPRdcHcknLa5N16kHCcu66db43
NCW0zJ4KIrt/nqSy5o4Qy2c1Wasazta+kjSWvfYGBA5bF+AYhM2mpM6ASgrisu0D0C1tsdM0JUB6
H6D48IzK39HCNLCylLtQ0ak2N5947wGdRTncRR60Bh7eaAcxk56GIgVKqqWx4y0chvraB5Iwupf2
f2jCwFrHVInQQ/UwDw+YYq6rm40Du1DLtOQcOlWEuDUTMQt0sItRvszBxw80qGq0rsDokSD9BMcd
PlzAvqe1Uu6A8+CV7nF49yyGIr8Z8U5AbtDs9cAXVROv8Uba1y4HLMh+CND2aiEB8GdhK50TAJ7g
2L7tDVUQRCZ+iBJBLc+xLRN1i0JO4Rdo3mioKvtvuO5+sME2UZ6gUw7+0pnY/iUCvUSWX9G4t2Cs
QTQavMWg5geFJ7J2RmjkiEEkksdR/d3K/Di0e7e7kzL718XDOYMDNCpND1GWAQJ3R6v5sayztbD2
GOApdcFpRa+cbAoXrfCcp8B/3U1soCZanhVmR9qvruCO4D0H+Oj2YwRXnd+yW+Cuvb+q5oYFCZZd
woU5jChtWkwry+vhZjMpNgvYS+JvkA0I1X/G7Zw5PfU0zMY9FEuf1P/A9+l+3FIsw6KmFjOwHq+W
lYISfkvd3eC5FzVniw47u0g5s1ulHd8m6rfsv0fUMMGwX4yFdwAyfKvypUvtVqwWiwapr1S9C8Hv
QTcoglU+p02jv/2HgO92q5NpRxh7a0tYW6wNQoiIaGrPa7Ihld03MIUxKTYVNjqUqv+y6dRJYDNp
+NMaZXsRJCibWC2Lcvk5OFwi0eujaU++RnJBO/n6UZx8b4vH+4CSyX3s39zKI4jZYNCvIDy51NhF
l/pwNiflYa9lKvnP8ZouKs7cki/FLJGiSlXJO5vEcLZFAOtFy+kBdcg8XlK1zx5CujTR/7+7ZNdZ
5Y2R7dbiwLXy1IJfEziNFQzaHAc+kSm7f+twd8QY6YZZvA6vQNj4ONTv7ZRTsJNq5NxMn70bWCiL
m7xxaiYh4jrMHzcL2/TG2bPOEpNGVk1/a0B1M77XRmtKc7h0FMvdAr9nG+gOP61Xx/A0oEKXEoeH
kZsaA/ArtVI0Hog0cu9vo4ZZffV/DWJaq1UTd6xbWSHlvm46AoUMcnW7yza0PadQnMEAX7WK2+pn
CsingobmVAANeJCm6tPZzGGKd1i5IkM+4MZH5IbHDcMVqd5pNQaFn2ceMhNcJHmNgooixLnMATax
co5YAZRDzdsOYU+vCqOOLysICt7Aa97teTyGKBDG1tN1EV5jwVhDMK2Lo984ScwlqyjQPpURJ3Nk
A9DyIaFQ7+bjbmIKRZE/dDCD0YCoIJzEZaKIq8Frx0rGz4BWPk8mRRxtXft+0cDc+cReJ4orNp9W
8GrtqlAiqUduW84JW4olwQmhp/mqJK1hU5qhyPvyz3HceEzMgWZMMtZPu6hC/iMwfW2yF5+ao51+
bHUgKS/dVqE+6T9OtsgaNuEv9XBvSX/9RZipFoJiep3oiz7civy0Eb/MZeJMZLrU67r+yyXlgnBk
ZXzrCbrNaJUd5LpiVnapaHPirIBIFN8flRC/ZX0FZ6c96lM0u5lWo4xEsbttYqq1LdK/37uDCC5b
m3obr2rqYncbxgIqwiMg422RxwDOfOlwKzig73n/Th7PmnfW9wJa2L+HrHCdzOzTjP1LHHs1qw+Z
XSRpiZ3tMBEww8SCESnXMMDmONoPw+CZW7Muw5Bpt5a08tLZWMvVA1UU58rIOTEAXBmnk1SiIOGH
Z7hSGr4MZvf6HMj97OApJDWR9W3iSnObl9lGvY3zNe9q/Us6SyX/WQSQrbekF3rb1vcgOpu+JMtG
2oKz2kC9jOkTEYfOJcPtMPUImtPMyMglam4RpGY9wFJc80qHh0HV1Qu6Fvu+ul8KkFGx3YfvDejL
bSTCo7NE1IBMXRJ5cn9+y8vAYPcJTDDpG7vKy38zO0kw/xg8y0+qUiGQHA2waEdUN2hmiWFcs4in
/G+6yNhnWULeBVIj/RKEBDWiZPN2M7YOSGzzWcOEVinaL6cRQhmfG/sVUQWRnuJCj8iqy2v30S+A
j1P2B5oRw2mTR85+5bQEhNmlSUC9YAcwmUODU+PHZ216kZncxz+63Q0UK2fjvtS8Oa9XDLjQYgfJ
vovIK+s+wIuW3Y+VLY6B2y7qJKYsYYfYcEubZ4TgqImbDoj37YxmvzNsh2dTREjGZ7lXvblnF4Ey
Ie/B2J+Az+rNkx6rnlQMbrB0AUl9X9K6bDN6mW/9W82ejG6tE9NPfL2T3+73wtKhzjkzo6fl+QX+
MsuwcROJx2OoId4HSkrC4ZmBXR+3xhd1d+Ec0e73dfY+5Ep8AvR1u6SJou+js6EnfTaoUUaFtS6G
zIxovYOjITYyAAy/BfF8/eQGeBTn1I63Md1HsC4xHVMs+nHXha3zPRpj5rMn8ugxt3LggwLh+5tF
e2UcxefqhkV/ll3KDIi5frAbmOfNIeCHP7dXmaHvCTTFwM0HMdFxRQUN/Y8sZw7axBs7D3GZn52g
ET8HBbGWBVZQJmo8NUf24lib0kVEf1Elf1yMXUXn2B6Qlae8tdchh+VaPkrBjCFMLQSrvZa46zSU
zWVuz0mMrxhIOvwqfTjG0WevDuEFH2OdS+GKexp3ukhujbmwDjUDxXaP4HrMGf5Pi8fMT58dh+0o
QDoCbyZRVCioluPzf5QX6rrS9lashjzMepMDF2o/+Mn+D3P3Qgj7OBpi2y5ZfOwhUtk6R33m9sh0
QVu4iZLSKqLQOUMe6tvB25WQ1/Z3mFSFBKnqMm7fUFJ80AVKxOvGSkyE74fVjc/ypPDOTX+d5jA2
e59PQV/fW6Nza7R0CtptQ9BgrLQsWeJkUUmWgRq+urMk2Qyps5CNRVPo5nm9XqiZyrjU63m5d05p
uy2q2Eo/bH5+V7vLrn0Q5ljiYEl1Ts9C9z6uiGkIRcTEBRb5s5vzOmFX74hL/xQv+S9/TSXVzyMo
wkdnQqa4wfCVzOLjQ2YVNYT54I7zlnBs+aNpa21jRD3gOFpKP3k/13ti+TiZvutkAprO2YK72dXy
aVuISWyzDw6hBHSFc+Td5sAXKX7AVtEGsxX9DoFoAMUvOWRaNM3Hl4Vr4f09NaSA6RtlA4n8BPnV
/9l6AFGRtmJRYruIGvl5YjS0ar+b9f7MC9m3XUCW2LZQCWaDs/oGTH1qgNEgSp3ClC8eatcuwxRs
sjyhAmbdZd086k2BX0u66pFsFQ6x8N5iaJ1G64y2ECdGILIRY31mW5X00zLJnYhpzLks2vwUP7KF
lq24iai/OnsqRDrzVW/7IlThe4Zf0khvUNY5U0XlbQscLahwjWsBAwQdw49yOIXhAuvi6IwSCxwh
qgIGnAMdwL2aJmtbn8QIDmfDfdasVEIgK2j4H15+V8YXQ+xNB1ySrvxMj9StdjfX7ARytaeuDpHu
p0pV/IPIDBTnOP2QO/rbNWl7By1krcOaHcUv36qJMdD1/YO8aKXk2hOSXF1mC9Q8fRdqq1Ec1d+C
DjVNPR817kFXmKs+0VsEDPCXKoKJc1TAetD4A4Xoz/VO3otS4w2a7hDw7PauIKCGDTsBUaXEjpLl
MRpH4Fzg5Jj+vOTk6gYBA30WIXh3Ir6O22hLmAuIRVbPD8OX/XfQ7U97EDg8s8GL3uK7g76lbPHE
iCSGjzGzzYk3s9OCRhz8KZ18jFM4K3tcE9SWbw3d16J4ohh0B5Zkz2cfD9t5kOUFRkL47hpTap7M
aOO8NonDQRSKl63tJ/IGDlsG5zDO5TQyoyOWXYqRJbbOJD2wcGr/0CXud3uiULAfErEGUEANTk5h
FhpaTaf2vJZgrhkXrpynUeS43/O8MfOk5WPNKtjEcEvfjMCmr9SIabq0lCt9SU/L6U9vp6TwMI5I
yiDOOH2K9WZ0zlB3HZeOJCxDHAC4qzQgAAy6UIzSoVobUvhPcVkoWH0Qb9CupCOTXiB27JSxaJdA
WlcLEm4X4KsYU4CQGo7A+E5B1nGT8oEquCRNfayHGsCxHcombjkwrYN3wF7SNXHFFLnhOMzBfj+R
ykQZD0tXarR2hlIlcxAtcOPhfPU6LN6uDQazZv74Cyv6EXoSO/QuEftSxI0SjZjf/LM4qrES424H
G90Xz+TnGWOT+BJC5qjAB4D6OSWn6HwQCsVPtHxL2mYav0XO6IVVjUykIEuhg+ZvQF0uFqexXJvm
v7i8tUw1Ym/Ft4EOqJebDtrbEFIRRt0PoxNVtLSIcrHzCthEvQsp9yuo5z+lLZYqI/7voO/4T08l
WyWUb8x6+ydSjtk2jtAWSisb18QA9WfzGCm51bZMDpB7z8FL5v6h6Suxu+AtTni/u1BgIjBx1fMj
lmHRpxP/RBRZl0YW6v/qcjTaWkGvRZMURn9FfwtWtQzY3x8h4s/Mdey0IcmT8g6R1QUmDrKF1+dZ
kbrmF+oNslbeq6LcPzSWmYrMhgsxvXHtGX9SFcUy+u2KSpu8fGdNZdzTEQwK00zgWoVBQNnUX9R4
KAsdcF1Qi+KaK7Cg9IXpp1WDtG53C7Jujn+Z5V3Wo5wldj6YjVaew7TCJN2Bm+L2/0DEla+ttwEW
sCWHA59b0MJfvQmp6gJudhbNdURawm232I+XEItWg8mfuv97I/tFhTpxWfKrQb3LIINUJJKICjj2
XAwSleIW5K4PK1z/a7i25DLI9qswMahivkKS8OJJpShj5JN/QUVQSVZRqWqOLQvChld5Hkoyxe+b
CI73f1uVmBP/ZV+GeeLJhFqtsCTUPkxDLASywynj/r3FwrY95B5+6G8kpn3F5mIm9mDpHrv2LUTm
1rL9vug6fokhaCpcBmh0pmRuXsqMuuEvDE3kGQu3hO2DMD6kCLvj3m/L2HxLUsELBV/D3daJC2vg
hp6CVYNfU2l3LVCGpfcJTB/CDo/GXIix5x6+bkzlnkPUoplV5/QAtImS/KZFsY16y5++gdQotUXT
ybremZyrtHbdYCmFqIAafHdu3vtRpvXHqJ+hcU7ScyxRNShtqNqYVKEovzmQV9dN+taOjTTPPsOR
w6X1wYG2zec3o20hrtcJ6YzNoENSRfXMURg3D3UNyjjBr6CIcyShmASy4Y8kJKPlb4ggX2zdDIHf
A9wVR60CcGDud05AOyIbZ2hZ50pHANi3StzfdK2j1yer/QHMersbUGMtAObZHp2fMH4OrFGCixOX
bYXGac0+MBZD2VR1jSZC+FLnO/ZAJCXA6T1ty8VoFMnDNOZlnfLhYcFm2KT3pAJn3NqA76cj+dtw
L+Hc8mFhFf0ghDrEwx+JMTreOZPUSkm4TUAEYNjPYFsuishZvcQfqSueZQpBm0B/2WtGs63glvL+
30eyB9qIFzG3F1pXAhCi7YXFwRsUjbjioZ4oxYHmT8ljNESKcoGDompQsySeDoW+E71rFuaF/gfo
lm+9axdpVl73LcFTXdN8+yachduhI2XJSSMP3RzRCQg7y3QnaKCsxcrX+2JZiTnyMk/lMgUUxel4
8WbNkjRY7xscG0ZIkZU1/P1QdUU125dJdYX9S9vbyvf3+ewS+LXomX4uiO3pELPpZsD5iIpqIlNM
/BXS0ZmHR8W9r6E4849zn6yiQiIhM+qPAskM5jWdKUVFSQOGSIIAsncQpwf8KYY64dTGGdolnQh1
u3hFp6tN1/+GDLpWzb7S5kekl0f9hK6tiEasCDOA0EM0sk0QxXeNn70kJewhSpAC9fMLBT5FVqsf
GLNTwusn3gAF7/N5lue6I7+7DSNsO3cjfrD62OTeXQO7ZE57M5tjb1J8tXHA+ySZy6HMOwM0jbUU
pjxLtGynbe4oD4mib2LrR++GX8bY49BfO/SgUdde+W5wXOSShAmxUSEKXLS5q5DHvN00k5YQg+wG
UK6iDIRmdqFH93gj4Ss1cymjSbTqHjJUG2m9Yi13pnuuWflCeX9WtUWNf/5pH0p9Yag3OvLAboRL
Vs/i9JSkNFx+STVUKpYZt4Ettn+oXP7en+tGbR9RNwryeSFiDMAqib8akRuzC6y4mxLu3J5jwxzC
lQYwaFPYOjeubHdEHsw8Vi1/3OU+saekFU1D+ipCkd6qrPD8z8UqnY9hNGguGAi+TVHBH3ZdTPSP
//Z7hq/sxUZhJ8E3in/LL+Tj9M7qsuZcF0+riXcUlK7xRi3Ptir+x1U/ukSdRmGBz2wOaU3X5L5n
UpjT+opPE6HpOjMbsvdlcXwAQ0VaKyLcqPgkZdosi+c9YbqVdVqY5hBDPmblC4eaLQimAS+IgRU7
4nW/dERoLdWqjkJ60h0vmAwQl2qeVFzGr8N1jsvbkOl3XLEEIeEPbRhWLHKNcnrJgnKJ/rE9adl5
s0GOIEs4zIP4ml1y/KILB12xHGt11zFoT21dSDYwdBd96PIdMwSBxl1wb6KLkd1trhborteVNalA
2uR034pVTARmGGAE4tfilYL1pKgU5dF54ihaJv53OtGRjHIdYgJ6xp2fPUc28FDGxMRTXVx4dCj8
ZhlyVwH/OF31JQm0hZDJlvTGVO9g79kKg4V6V6tdzB1R2TmhuQyGyy/KDW4FFMxCHj2VH9AJfgW+
sPfkjPr6giz4HGWVBDjlTPjRTfI5uUjElKbfb5PWQ8S+nYf5sr/L+7ySk3WAIBdziADK9OSKe+Bs
MJuQ93SLlvINopdr+BA16IMybY1lqiujzjfhkIW/O/m8qk/lIF+AjQwOAIsOdB+YidwW0Z6HWHYa
ZgDjYpvhwht22J/RvjAz5U3JbbijHelHoNcFGB5+7ylKlhZf9onot6Uu9kyV2ubOb/ECWeUtfI+U
dRBwfRefev3HwJQ4+tqO1ectsFiQrMtaYVSNkwttAKqqPMgJaq3KNcsZOINMGbW89pXsJmdBf8Px
5nVkeHczMpJ5jxYmazjM4Prs74PDG/EOlTC4HQOr2WTtK52P0bespw2/n+XCHRxRj662KPO4mjEU
a3AY2MqBUt6NYg7tRuuqRwSOhWaM27tE0dg4AVh9U01SX4idDTk2iBpRpgOoKoSxRKvZuqQm22hD
9sGd/WBwVE7J+rtFKuzsfLpwOm5VE9Suj25vPnOE6mSXT+SByh/GGbd9Mi7Cj8CMGj/Qn3WdGFIs
+SbLngfMDpg047a2D19pnf8S1M00wWaoTbHuUBggwofJUy15pYqPWpxC4yLWDPl9Cx8khgBgiYRf
M6jC4w7yGEJk3cDjXhdic5lHmm6dcI7MUqVrJ7Q0EoFKNpHXtMp+sx5HT+G6k+8FQmYLjTe/tS6p
24pGLlxTNURNpuPWIbZJWwvGZn7XwsrSjKW2xkkm1mntyaqIIVoABaPnZHaMytExmlRl0cAQslcp
cnCDUK7E/4Hp5CMNdZjxxvE444KIquc2lM9fK86yhleLwl+VxFEA23aGPFnLnpE4vDtAjIHsJf2X
UsxHnMLnwrKqOaPjlpagkei6CoZ7+BZGEt1covSrtsKWoDedledQ0KHe66kulq9wqMHh5m9L6+zH
uumKTQ5QFaC/T/dyZnIe1suIaznr+wwSkslsELKTm/Jx1H/77XrC/BLBlGNTJgYoeN3mXcmRbZmx
qDNj8c8DQle7D4kOmAN6nJYmm8JhSxLWNW3BkGxKC7nAIsQ7nui+UjHkS8/Y3NjtKrDDRuf6AIYq
7N2LAfz/IbqeDoPS+ocCzWognI8Y/6iyGwfK9lzZJfc7i5Gwurbj3kpsGFufFdnq64t802tL017g
QkE7rols4I52WVgGrn8oyhDW+VTHgdNzdf7rREncUw88eEg90Ydsb4m2frsqQ1EFXATZIe+wMCqx
Rk1dIn2Ie2PMlHyt3W4udwgBu1TBSIDOPTDSVn861DfaDQDSYWGPR03BJ5u2SkWXRLmrXGPBl9yd
1uxGkeQ2MWeWyP2yIijg9mY2lz/tyuOjP67/KAu90vIw0HDGbQzoyP5nZyTdAMUBheqfooN11Bp+
eGFo0k5AEgla1B/1BSvb6kMG77AMIH8KET07msmQwmRaNhNCRqYtXKNuGB80AIo5jBnlyGBGZOt4
AtFLtCRg1/whDAhSZ5EX6vJYlzQnkOx9AB0IFr2AdLHlEVpBlvs2uVFBlk1XUGOk62pNis+1qOdL
EzSNUCm1fhbtMMHIswvDVDcX+OaHVTOH4HRtNCgYFUyCzXEqC6QLE0wTOXsvIBNxeTMcsdy3lOIK
6Baaa0aIF9a9wW/NR8ShzVOdnEW+EyE/LEBpwuJ+i3n9KyBzlFH2vzxOT545UsCL578jDzCiirSh
qVkaHNOXTu02pWw/YGT6MlIpWIMY5q8j1BaF9HlmoyRrFzYj0yey5GGYJtQECdjZXzK7VjyI4D17
Qis1lapF6LRsMqj7+SEheLEa8Yo6YKojXxMTTeyKvEfRRHw8orHPkQPsTveFbdwHEpbSfGG2HWmG
dGfmwgJHkqH3yrAL38P6zov5+JjINRRi/GGMwYR9CesYN+kCYU61rYTcP7wNq/VUDGuUj0a4PQLy
IHZyKaC9mfSxOUvjKttwR5Zar55r2uaevKJFV1BCI9LYjighEEAFYLp3WSg0hNqZDMzVgQg697Fr
eVAU1jrQcRuiE2Cscz5+iWP34omfTXfibF23cALbklP7XfdfnFbFIsYcPEEKImjBDJn8MScJWyT2
Rq4DI7zShvqn9BFLq4JNMWDienYfKihKOdR/Zme097Vk7JPtoRoiZxwYldFLr0OOyL7ZodD5HQSy
YWyCzfu9LM+Dzqi+UHrCyryx+UKaBpNjQwFix5zTkXisz7NCl3TRIY/R1/tl4EY/JDWuKMT09GNU
p6jKZYDL6n6FxfER0+cNSytWIka/hzfeqDM+Eput9xVH8XjHDwGuyYxQgLrw7dvp5iSq4hgNNfJD
RClmgTUxOAsSyWFWnq8vtgPmhH4kPf9PXEuASwTbOrcsNsIac+7Sa0+373+fSni25igAsY/KIUZZ
fzcqbVID/OIIfF0HXEUXiLgCaTn00xxXCDcH714/jwKjohqNgwfz8GOtFNJcc5ltmhlATVrZ+AE0
Fd8yl9gsN1C6d/teXPdzZms8/pWbDgKMNm19kb1UvuiCOqLmRLCV8EbP4Con4Mkeu85VOirb9CSR
X+hI0bQqNUprRQXUZiY3xzEBzMac/9C+qiL81rnfaA+rPGmaEA3aDIGv+sOA1u1Wcm49635Zn0cs
EyCYJT1hdQL9OoXt1kQT0cHvyCIvaSchbj4UDlD2aYYC1ln3u7WFIclezsQ9GiqiWOJXlIzNADaJ
a2axsNAU9R0rzhFkcX0TMZ4IfrblEWBzTzhlePwXqD7wJnk1bUyw+LGcdQhbYcSFZH/LAOFMZZo7
wyp4Pe8L/ZXEttT+A3Jq6DXjQ5sRhFNftyHD6gUfq9AYoscDEBUXcGjeUmMgQPQWWFUBwqpna12M
AMfahF/+Yf+dBKyCx2lpUHkHBZZzEqfI5DILVetKgPoFv7tbxtwU7VQR3MLuQYEwSzr+159TrQKN
ikS2a/tqliXXu4zNa3Dck00tvppTrcu0JKRjOyQaRJAP97XmY6zdCeySTdv+z2HDhfUY7QVSmnbY
grJ5VEDVZESNRLvRHQQdLVtmdelBKIjnU8reXes9F3mgNyRnPvhvc1cYhKYoNpCHPqkeRpXNuXmV
7YNoXIdh9OyO22QoDEKjJ5ng0zP+U5cIEoICJyodNg4OmZlJK/80xP4ETUW9DUTGs5rQmJXTb/0f
5+HTtsOPe0m/v7H99i2eRImVxYnVQIxw88svvjwhtCFZ2dBNMb9AGvixCwFMloqEazc19IcnIJcf
lpN9qFiGF+nwxzmkR2GJqQa9mM1vajsxkyxvIFusmgnD41LRd2xg+ByXBnKoJillhkyngbm8SzDb
dHHJWOso35Dq7Z/28KwgMDwHxK1N470FikC12tMO+vFO59G0P11omD8nprVDHD8OTEX3VHEd+nbT
2jaDKAnX9D2Jc7CwZmDwC4fCVc2mLZfp2JbX2wkfSI0RK5dNXfarU9anE5On69vYhqYVCnb34hD1
VUjbOI/zv0mgWeDhNJs9RB/BXM5hkof2yCfpB8Y3JKQ/zBQRrJOsLx9r6hOz7okLrdCWcaAbU6+0
QZNl7pKM7lBLQN2wWri6EU7U71crFVFcv07pi+QafPcPGCwX0gj5sUsCL9TxEfup06L3M8zATC9B
gXkMlpZHXxSmycqh7otXxiNzjFIIgBeitTYm3qUhBHJBxdNjRvtulL+KhgjyKrkjuD5MGLFamQDV
uNj38JWGjA79azLmZJgaZWkIZNJCya5SsUpo3wyFoPaRILCP+Tn/nc+Utz/JVmmG56YY7W5h2l/V
DAwGM3vZtmUNxD3cOL2+bGS9mzMbrzbp0QxlWOeUOA8FuwtqL2mObv12nr6H4OEUobiVU+XJUBLu
x67hT0e30hBc4Tn5iC+k4vZp3pWiRZIPEbHawHWenavtGlLFKBTzz+wwp5nf/WFex8tTEYnh4PcK
EFFWjFvwGHtDUrYl5IWDDYLW2V7C2fyuyVTD2sEfMDyPaqEESy4PGQANksBd7fqQB9/WJL5AWWra
jiDV3H7hoK65ouiIFPwP4BNZCumfOMmpYabcUpl/lHDHM/kM35XvxBE/U1jQs40qvIiTp1+6h6V9
YjvhFr8UqgZMYgZRLpkqfp3bOpeijZWY+HHXs2g83sHwZd42Eu2raKEPdWlkkPaLpTU9CXMujkUc
0kmGOpaymEOQOp9Gnm66fFlxVW5IiiByLw12DiXK2IiefzSgEsw7lXVInvYz8yz4ovR2UhB8ADg3
c8BtJLeqVDmyKoiiB13ozT9QTKkH6nmKfx4IeNyqAucnn5BSiqIBfl6hALrLmieelr6Uk+KEsUG8
bgcEOmUHA44h2Fy7MwTCcE+zZm7ASCXQF5pym6uNVOprDEsd+JBLrwCsdK0Z+ZdMar92jcjMFYME
YZVoywlvM5B8kSgwIKN5ay2YTWbTT2a4XHvh/YCpUc8+UyYrSetbMcU+GPIJS+Jf21D8DDGAO2gI
imur+rhO4wZz90QrMigBncPpjRGI+nTSwS8gMiR3Jy5YP007E77nk/vDQY4aQj2JZ1RvtwQF/EWt
GUk9AwdYCAEWjMlia1iGs36qAOiEgvXJ6+77c0fk4H2tZHCeN8IaS3xo/Unh/g7M75PkTI7WP2H8
/HyuhBHcvVyCmVq3ye3Lq2urjP39iyXsRUvif1Z2PU32dTmSIHSXdny7kRmmrtXYPFRcsEcofbuH
rthmbE7HQPodE9JuisPeVOcxDBUHLWWcrkFsvifsAS7pv30Qjj7J8stVG8KOY9nprI3JGPWnM534
0Brd+epa6YEwZObWsz2XyapnwZNIWBOwPeuAORq8og4rEjUrfjLzQYhTA9bBaYfoissm9v7Cba3X
5gwzeMf8MPdwQcK+ufSAXtkLBX0H2ZRdK862DApgiWSH6rSPUOJ6/MxqGn4EDT/uJkCmyEmwvynu
gu5PWgHcEZgjsOCNM3ycZHY0oGBmUn2nI7iSoD3QptGLe0rrYFCphFGxAJsvvwX5bCXIuFxsvNin
2e5CEo0lAb6IrhToRycMiRA6++ssZT2napYLI0bn8iCdga7uWPvMX1IgdWT4yoLZ12NJ9+OnzblP
zddgf8nunuq86QBPwCT6KQaRduagvbxbsik8/CuX9zJCuggCzMqcLmDXB+X2OYd0bF/BHZB98ap2
/4v5Ml/LY25pW9ud/EeCcs6Whol6o616ZW93JZG4lfyaH3Rgmjz2bXr7PuOmzBJIh+jGrq99cRWr
r8JKBCR8PQZFU2SCIqxKyXw50KfZgin3nuisApJcggQ4pn0QhzXm6kuFeS/d8h2MKcJuD+nwCt9G
A6EeHgbtBp5xhvJ1I4kckKuktkd9QRa+DMtIPVn0UVUX45I4UtZp7Q0eKP8DXjAEtXkJn2UDs0Yr
brZt1bTvzD4asq0GFoC2TzYNe2zB77x8rT24RVI5ePqcyPESICuqTxYTrQKlL2ytv2AMa9dKcQp3
eIPKt6D11kzg18HjtcJO3Ue+2ufIHTKX5GhECrRxPU+OWRsBs8OCaCKgwWDD9GO8h/atLcCx9fzG
GfIuz/rfprrwL6dO1qSZ2PT+o6Samtp44rw0J9hffjTCh9dQUPtkVICFkxTxCH/+fv3NO431Cpxg
VUvH5+1QNg1y1tXS5hAVNOh8oMAcZcmDfidiKudonM19Zv9iT+zsoTtA5MM6A4XLtMIWYrybGcXB
LjfnqHoWoQoAE2CIZCCkoEin2L52wtUfZBqf1M5hc/Cb6cqRMP4eloaLXqhTge8TaRx89oP8CfT0
i3laQ5ReJuGOfU8+YKIHzVuDEuVSm5jh7QAqy/YGx/M89hT+SgRgQfwk7u88bM/+8HLY+c4bcdf4
/UxybJ2Kfj+rjYzeGrGym/J6Wt+PgVtx2i8FhYo9U3UAN2A0PoBHNg21Ku5yZVCDcFMLgKn7WazU
thH/9k7Zvm5OhC1HGQzd+Ahi/UHqMh21xm36y7mrlrRbrCowDJSi4csRRaHssWLV3tJq+nEEGvMy
zoU2k6goiHuwhU0Kwkc3vnNy5K4rWZUQmW4itP89og1bB+HC4RV/e4K837Uvvot8S2738XMlOc2s
3HClBSaM3JUzlf3mK+eNLii4vNxwPLxaU8LzQkHDU5A1jIlrjVkCTBGNaWq0pCfX6OVuo+EpAV30
e9BFDjbMqkiwJ/cq1D1IoPZ3v65YvEOb+N7gxk7/imsvEifMtjK1NmYZoGwdk6MziL3koZWuVoSG
LhelRoBKVbLdc3Xjby9iZzZJeUZTHUK+7vMHUMoanrSBuaHlD5iIMEacnuQxQcZKDO3aIxJ4PPPm
dJTowk5kjM+M08CbLJfV+RoUT/kyKuABkGKnTCKGbtxGGmf5uLSH5a7c9Nj/J/ght8B63b2yrIeX
QH0ehDXlWx86NfruxLkTFWaGci/azmPBNU1n2Ohh9HTYfRJOYgiej+aHoZGY5O+FPh+9ygxBmeG6
CDTvJ94JyBU/FkEMe4ij8cME04bSzZEfs/CYSzGVa29OgS3OblY3KoEz75fLv7mIJeZPivLZ5Muj
eHAs7Nrn3VoqQUn/epRx68u/oA/RlZJF+Uzy0CIJQzYp+LxNFM1hsQwLZ02yxVml9o6IP/szEwNY
rf5XNBaPuE60UOWmuaB9dlwdJo+wAVBF5ICuxmpN3rFDU2yxTO3WI+Mm9u2MVmRFmVWVDYjanbOl
T9QoiXQtA5oIRRCheeRy9ztFABLiGMEgLrByD8eBlYtnHKeQ+UjiO1Quvbb7vRf+quw2yMAyETfX
jQ+2wYr0xRy+xTacOf6Jlh8kfxRlTllfy/H2bVra/Gm/QIXooWwkojSohJtq+C3D9SMX5y3ImyWI
39gqJGMFsWJn/mkOzEm0MMVIk/eRHWputVzyzB7R+P/DefWMhgoh1gC8UxZSxdebGWogDiLSq66q
EU8wY3AVYjbP7XreqTZIMWmQ0FHNjugWXyXbTRMuejwlg1oEI9X7+N0MjdnN6x5xltuVtiaD6aKU
1MH6HhszI6dnL3fT6VudL/cJWhlPKCA4Bv72udghAodyQ3NClDStakt6Xf2zav3dnrxcxXxfUqpe
6CPaeSTvbqhOPVF064R3YAw7M64DMbshHQ3GX2r3JAEKHA6EQ1bjVCHOnnLT8lAiVS7+1mdZKF8p
NTjUprenetJoqYPTNXGnyIhPwDKac6LLfDEMKV+aEq2Ppg1ke1Uj39a5GZnW6tFvlpkoMRpdDw60
upaY4HTry+MiRSXgOtXAvMaQ497/D6z8ANbkF6OR4cePbRAw5MUmDM5cWaoMrt0QioAgBp43AY/G
mFhMJ2tKD1zvnlH2LT7Oy5dj1bXrpRIY+AMOWdn53n6+ObdxpG3Et4tGRZS9bFg/fBOcDTG7gG8W
uWxfT3RXhAbzC7LUPw4S58ECqEGbGa6nzZKnNzIk0e/h5u79T5jqqaOzLkrGj9WtabHcbFo5/ViB
3cjruzQh6TyYiFKXQW7r0X33PIa49sKGWALOOZSo0Ldk2qvly/NzR/QV9dvb5Oynnmo15E88MCVA
cKxhM5GgHYlJ2qfxSMwgFaKLzYYz4j5RxNggyB6193EBWIEMKwhhpJ594WFMIGs75y2eGodvIMhy
dY+f1nU4Tglr1fPBHF7CaFFsu0ai4k01JQF+HawLS7AkeqPQzCBUY7iVZ7pXsYkw/H4Ck6iiMCl/
jIqnVFN4sGkpr4UbpicvK4R83DYsUCoZf/8YKu0LAQXLHGgql5k5/EhLDS8KF9VKTjeq/oTKVxTs
uCfv4EyeF+DOv3eK7LfeOHq60rkvhWmTKj0aq33LWXVf/9Dc5khEMr9+xqUT2wtduxgltX3fz3LF
yTmGUGx9HrAzPuyqbUZTcFS0MNFaZlWQpMv8PGbcfV0suk1h4TZSuYwbsoijgCNrZYej61K5USZu
sgznZ3/xWSGEcTwEu+hucprLBV8lrXxr+DdYqxxQxq8fTNwv6hv4kubkBrTMuGTJ7+BfARjVpP6x
y92w9G2LhJgp6RBaby046dBWni2kV4vKcJEuseD9gZ/6h10vuJz5P/R55zbBjkJaAAMI5bPasni0
aPavSemGSOPKK7GRt0IA24NOcdnbjoYTuww5C2Z04zkzYeAXDNziXDKIg2HPB5+Fk+Jzc+szEoFC
J7Snns+rD/YXk/LhAxwmiAcFUsyHTBbbXCcgw6KO0e1lwEJMibnfDOwXWadIOj0sDWcrM0SY3jCV
RxruPrTPl5sV5EbrqmKMY5i8VLUW0ef1ST0Vj1TIBwFIiP0Yoo2thUtbco/peZz6ZCiMwQQEW7ZU
6vz1fjItQjzvGuNRmP0fUkMB8QIoOttRRwtFc7Fyi8HQP0Zw8khnMnM0Eaa7MtVnL1XC4DalzT2f
Qliu82AgwwhaxGCQaDdzwKk6iy2u1G354m40aK5JcvQD4Q+lsyf5H9dguF4CmSUUPicqEq9m4WWe
RxTLMPHlZ+E2LmGQazTVGvxnaHowRK4oW1OTpSaxiWaI6VMBW1TyEcFKCXqr+yp7z6SOJ/R46CRC
ZU1F3jGNOhK/tI5KneQiowd6q3zLu/PgTPsEoPzzm3gTbF6hOK1vFCPjtt6NmyJBVNN1a8OxO7DK
tbJkn7snOI+QSHMRHevu9kMMhiNWWeYtK9NNMCkNURxNufNvXCvq9FSR2SThZ2ZRmidzgc3PvY+1
tEFbThpyw0TzXSUEfCypaiqsDfI+LiHG2Xh6tDYqzaWLIkkkiMReuHA410Fbb6Rnxh5PKjTIDxfp
gd3N7pv0EjGaUdUfO9lqsSew+DMiM7y5/cK7osWg7fM/4j15/fXdYMb60YXHpcuaSJSm6ddC72mf
1F9ItFQJryDIc3CZNwGv5LdVvy9M9JDG3SgbFMdymCmKt8KMHXj3jqqVk4tLGcWxaM6FonacfXhQ
InXMVLUiSbMBXfzo7yY2XdwDcA0pwpHO19e3BAJH9VUbgDuShlHf9s2XAaWFbkczdVrEZUfZn5+V
TaAdadRp/wRlD7T94vlXoQBA7qKYJzGu9fvbmAxTEFa0C0+Oi8KrQ/hoLaQm1MSbFUOqiyww9KNF
OKQAL02FHtQQu8z0vUVcD0eJqeJlJ/VvL7z2L3B6HcA5rOOHuA1M9fZar84hBNCrdm6qqRt1Ge+c
StFQTqvvSFkJ7UI/97xN+2u8AxAK6n7oRHxLSsVc5Nrx6EFopk79MK9C4Rrj5fWtx4Cbiy0zLW/Y
W7FgkPvJJ+vsrrsEkGw6pAkAX4wc3K/WEqNntC0dk71aHDT3q57N4g3dx9/ktc0QKAiLgeBRXVWk
nIs6ZgUPvVcewrtHomjqbS5vHT72UlCakpUhGgFGdqmtuapa+7LV2pmn2SL8WWIzt/MT3RouWuz+
/hTpLrlS/opeFC1SKAZTMTBA4lFdkNJSCL18eFXQPrmGHvVAlnKjlVhVdEM9HIEhHfxIerbAc2Zc
OV5VRqwG9G6IsrlJ8iiSVyMgCzmqK6YoRWeEwe93ssNv7qWe+Go8giqkO1PDpdMy/BdyYR4uUlvG
JqP7x0IZar0FNbKFrPVGDw99RWJTkQC/3r1IjDY255XXWMA/h13+EIpK6on7R9YYompi0lW51W1o
7SwJsudnlGJFJGl9hgQAqEhOv3XKPhROFwsEhztPwo50mOeWhh36KgpChd7PSolIcNwz25nmotVD
9TvTmU+cPA/hRfOqQZy0JPFhiqYu8Z8ABbiNAjsoiaI00REy8ax1GNFmuQ2q5pbe47Xf1kxL+XYY
CjfXvfgI3Sd4l66Su/Njpvy9RZStIGXquDv2wjbkQEN2ihV553iqUBo65hRiQYupRvkZMcc5nHr5
XXSmWeo50etH0iERrHELkCXZ1AeEruqvivCUGHHHd4TvmgC0S3Cr9SPPb2k52GX/lwXCkr7C2r7U
OlrD426Tdp8Sk34LtiESwbNfk4MinAxJnRLI/IwgX/5h6dBOZoEcxwTF64/lLtDwklCwjJahMGME
ZZtjUVmaJiy1Q/xawT7Kc8+tE3qKa8TSNE6dYNeKONfGQiLiAbKXvuUq50OB8y8/ayzUHQ4/8NvP
KyHVXFL6sCzm58yFUMAOMWYnhGQBaRKvDWARuiP5tZ3Btrcg/TTnXsFT8dbBoO+ajY738gvnAN+f
4SKlRcDBaSieUry/G9j/98sFFdBiYf0321kgUX5/7UILUioCb/bgoCnIW6FOizc5It9GSNSHm9yT
vRDVIbgwsnqXBqp9tobelAx4X+dzgHVLL/P9Tic4zQTe5Jf3ciCOXkhZEoe9ZdGClL3wZJSE4vH5
dojJHb+BUu/qE44uzIoI18To7eiqy2JTJgFQ7YWjKlhQhmwxH1Q/oFvATyyiFGI7+9nVEiNmgfgV
arFomFdEJWfhP3Iys8R9i7A/CxBbA+Y8P1vmvy6H6FdVAnU25VUQ8aaiHx/MmS6PXLGq2/LHJTbd
XM8UOIHnYw71JMxXw+WN+KN3bsbJ1bMWbDM/0NJv17/Pk5cGRhq3UzEuaHuY4qXU8dKAwdGUqdEY
gjVHzaloF3Dh5fyThajPst8esTXlicq9gMV4nmJU5S7+W7oe3FzA/Y/upfL1yGrcbq8fq7N0tG5L
X47DtmubTpKCCyMhsJwIhgsjrktYmZGpC9/EZ7QAm7I1yKkJ9fqoJ4bbHpY1qcg99uPRzwkwn/0Z
qg/qsprtnDp2+QY7ZWo+KJXN3rcsDKnWWGUDynOrkutEOuIYJwZRhuL3fNqVVPh8DoZg3C0aR5wZ
G5/JfMwG4L37zdfFbT2f539hWKcDGtCq2CVtm7zVOI1ROx02R7VN8HM6Vo4GcRZzJqfQ9JYUKohz
NNSYVBOevNPv+ynCo1tjVMBsGehVITi0ZHUX842lDHlgCjnDx15B4DNbTzCMTBg21Pm/jOCh2sXx
rIkpohykaxRvRjFmzInYid186nKQVqcyFpxiL9QSleGF3yjhf/VznSmlvhrJhOFdH3QOe0oD8nU6
RiBRxGj//QHrF+Jjfg9lOsQEU6Ncd9kFDxDUreuahnXBcBFhGNZmESTUSMp0SLsGfZ+177fTbJ7J
qBhfeLLAQocNAkFFH738ixXSkAU3yogNMTfAvM0GBnRlRA7XsIdmyRE9dk5pgEtLQUwQ4ipxjDDJ
vVfu9sIYUGG6bFo0LwxzpUH1tc9r13EgXl3ZQRGvaav9rmhx8UiZWvqadVYpwLvGi5YC00UzuAH3
dGkIzcaX8Qdl77TrFe+byRSOZAdWBX4NNWnuPmZorP5L+8PLKrfDDZH+HphixPSFbTRCthorAzat
iGkLMaWg3zUr+Ao3fB2q6Ks5GZ7HLC6EjnQAgGDMO9VqQjnxrF7cgP3qn//Lg67huGig0PBywL0t
ii/QMg8/dKRtEVtPZ5H8SiboeXUtNWVWWXXWd4ZPQuXop4pkgZCB0LFi9ROjrozgUPyyruHOSFB9
ay/hZbXG8lBSMCBs22fRq+SYL1ZzlGbElTQsfQ8q6MGuDrceqzz312mzbFnyYVcalq14qwj1alj3
ReOHpsB17I3dMNvurDhSzC14moyb/UjvAGdEOSXokoPuRuu4oEavgMnpho13jdOQ14HikVjyEz5L
TUqgwRXPl2tQSmRuGdRHUsh2spBvhckZ2pBGdTEsWjnijF2flKjUaKZeE+dWvnfRM9Oc9sN7llCh
QiWNS/OWhOhAU57lyovXSm89pdKy3vFaSkWCSOzOW0Tar0nwhb1ImQGBmlJF+cjqxlkKaVsmfFgm
lue90NpRn5vNP3Bosm1BcP+Wso/w1sGETtozvjUkPY+s0Ji7Gsvv4u333UGyDiMTpATRNqFkkozn
jIQ3+U46NeMEzLnLdLEwKvmhJ82whBsRQH6S98oEEAxCulBtjHcDHu7YUAa2p/j6nqf6SEROI3+W
t70xUVtFrfmW25ChUWXN0jyTke1+MI1HCgfxacCth2bzHMcVFQcaNepJkzTv8xEdbhuGQzbtE8iW
y7ldennvzr5wTWPtnrwGugj5AY/HqNbU1XLzNgg7sOwPwEkrmJ6wT8TbtPyIPM4hLEv3bV5FPclA
ty15og+ITxqK4zRIdxvD+efeYIWrttfy67Dh4bACER7kWn20Gm5wsdqenuRJO9tsIqQrqBN2bndC
+JcqsQEjYfH+GwNPKU2GZ3jB6tvAZznOZG+Enjmh8Lce/1ivrBXZiWILYSIovZ7ylzjGJID8iNTe
n+b8RTgoPHSTQvxK9lFzrLlZD4wX8xsgOK+I4FzBV8Otr8jeE2EbfnDC2Vyy9IAxQlepDEmypHer
mzMsVWvITlDZ4Io6g+3c1b7EnB6BB89QgX9YfAlDkq9dKlefvBqvL1m8ny7W4fGWDNjfvDT2uCLi
rznCgdWDCuhd8COjpyyBBwuWcu0nCn+5PmjX+wbweqNjG/7bTeNm0rvTn0UUSxSY2/DrdulZ+752
UP91RQJSkdWU5GE//2iOYR+idPwH/Zf9XlgFpNt5WMDrI+L8owDXEQe6qeVXaEd12QNNoxp7FGDQ
q78TBFQX1b8m3Tkqkh4LAjBDva7TD70bf4S7g4wueDyh/X6NuQ2UpYjOodRp1FKfmgS5hz9DPvUc
dvJYVF6uq/4r6wtlNYa3Z1vKfkRTSGezaf1Rl39zLIvdXet+Oihr4J7OZ3wh6LI1CCyvGiXFY6yZ
MSBepOBrLsW/8pX7M6Z0obN7yGfdcWi0Hk3lOxTXxTAvrd7PyrZSQy7oRPzweVSXJzYn7Urjpav5
yFlUACckg2N3hXLIA6hiRwkmWKUJduKfHl2t/qt5dpjqsH09lyOt8YnY/iHECt+TCk7zGLmZr9hd
aI1f659Q0oxso5o3vOYpM2NcZ4K5L/xdC2R1Ut2V2NrFh9KAy+C+YmM97O2I2AB+Rsl6/twHrEVb
WbG2ak2hFs8rDH3WdKrv4xNWdhEEutYDiB0QK3yimRCTaMXIfzFB39H1jRbOZKstuNcweCxcZYqe
+ztIQfqd8rVOWPJUPTRZMTlUk3pA4vkCSr4hxIOXfcJPPPjiYhr92iuoUQ9EzbBshx2yxTp7C0yv
E5XIOWywrQi0zmmMSpM0I0eyvyublQJs/TNGMsqYdIkn9A7bu8RjxrrladdqrnxNtiE9sWZ1Q7My
1OEakJ/TG/86C/e9ZXAifTcNous9Qm+hEdqxTkxFLQpDYNSJ6XRTro/wxnLhHiIZwZmBLVtVd8Oe
bR0QRuwZegmm9u9M7mKmDf2/GF+2xUtT85ZQ/e5gA3AKWR77TXKn0VcZk11T8L/tZ7yOmUJoxcCc
FtrE3ZMCHXClWG10VOE2o1V5j0JiRMEolTpL0lU2j+qK4DkYx9x1aNC6YblcFE74nrujL6QAC1uu
TT2EX+vIqUQnoidFRIy6GFz4hvu4lBG4ASEJ5gdIfBoHEGgMhPbtcZgQU+vHnSUlaWB8KscpLCx0
SzVB3r6WXuOzUW8NAMTIG2832vT5UYeRTmOMze5PnA0kiNsifs/3tSaefGWYTORNSHCHuO8vDD6J
aRAzmAmrMofTC6t7V7x43ZJkE4PUiFYkbnMbTpIVNMEMHr/oHRrROAp63AVyON+PV8g2v4jl3544
741n6AiVQ8ZYofszVHJ1uU56Ta1KN/zjvut2312COBc83c5zzf3qudHv8ot7PXrDFREjHk8OsAmm
ZjPl58vTypidpTpRFUE0LEMWkCefeEXk8DDicU+qN+JfaDAvdZ7Z25ORZmF89bCD+Jj8DKC+hv0A
fm2E+ltFvkrj7Sm9BwW1WUUrci6Jt0BjX3QiK7yiTVCHcaW3J0T26KxjMFQRl7r9AQlElDrYdppz
AfFWqU2Mh9PjZKN4mmvVtU8Jv0bvVz0PI7Cmgcp15TWX+kzJNma+9pwdjzjNKaM0dp9yzK0qMU66
T7bca2KeKvNslvDfjp+bbwTKO9F3rrQPKt+DucmGuYdDtEBXI47qxIH17+BKNBhiX12GyhN4Jp4y
mUhHnlZIWpVrNVicGD092Bp7xLPjmLdDfvL5rEaWRxKcDXzo53DYcK5wXgEV9frxviGqSywy04wd
JE+pYklwSkU6ErVUxoEFCUmWBMWvCwDlRtCCp/hIKXXR6j5/MsSVD+CGpreEylYGsGJCaYKDLiLN
6lIYcJzWFB5Yv5isW7l1176KZqbCXmVgQ66joteAMNvRdAfriUVos/jNJFYTAav6QP8ZTxdaXB0m
RdbmpFFVi2F4oktFOKGxAQGBSZMv7gYEeiuwwC5HB0wOWqPKZPlx2TIt/85+T35le1/FixdQ7q8P
ESwnTC1EIifHqwLzEcsxPaKvjDJKDMpYgRA91sEXz0xkMUESsuZ2gHIEdAsbavXEuQBVnJqo0dDs
6npHgGK81pbdj7ID9rkbnnxAvXyYdsZ+LKkdKT+DQA7XB6abUGhhgdO78x0b0aUwi7l4jb3Q9x9e
ehzrI9q8lA/zsQNnReZeaciZMs6B6/MViLS78SN+73IdKhIM5dJbY8tAGyJR/kXyOjXfIw6gOZ8A
cHSe7hhDWi8+LGsfC/jj1ahlV1K6+zO2XnJ/k+IYtNNOF1KEKulSdALU+IPzbtHJzdlz0irc0586
B4sG1Ik8NwVUYd625QSYV4pGx8P3ZfEndTQ5D2cs0uP+b+0QZHQksu7ZGQAA+4BeH3cYrBx6lcVp
Y0NSSVb+9oUY4NCd7At22n9DON1IUz2vkzaKPHXAfLctOm3OsjxDjDE12gKBRuXUKKUCAIvK4NOe
RZ+odBHcB3FZ04qBjdu9fdzrq1su8WMwxRzNoT0O8oeGSP8v0fYqFfmINT5cG/aRSeBlkY4AdYiG
PZAYImavX47KVOZJunrl6CCSzXa74sbTBpbhSkE4L9AB91tPccGaXG2asoOjbL7mJq2G62f6SUrx
4sY6JWMtvrfZy0uGqGpEFctYvl4RYsACusUf3f+iKVYLWDjW+uA8PEACvxJrMaKGTWPHlAI46H2M
srj0MD5OxrWsnja03JSwMu5SeN3tAGBXuHrA1zker0PJ7dmbMpb8Ht/iIYIMlQ7/+y6bxR+2Tmpb
deFuAgnbfcVuSj8AhWCHnoXAQlbopLFUYL+1ItbYlqc6YTftMVJ2eVu69gC3LFaY6bdCLCRPOP+l
QmtggFr9krdC6EEsa34JunzArX4XvJYuk5y6c4rtrfvgibMEe+KErjlZcTmv9HS1kwEl5ZaTuArj
zd7BVndgjgDiFf1mfK1m6z2gOEi3yuBUvx5892RXPI/tKY4BUu4UT1EMWDOpDDntzWh8jBLFg6Mv
gOdVjxrupdB9Pd4LKN+0fI8e4Fbf0QQxxgUrrkjidCfRf8bVT+IDuHZrPWIgXqugRgW5u8+WmrjY
QsdyQi6uX6dQSFViGQAbMvpzJi6q7ZoeYaSXEkGMapMJaJ8vywH8rIbB7KIn8I+28h773EZNJtJY
PPzcLVxlAVhP4A9w7qw1TRVqJEvWGcJgIJwlkXr5yqx2IgJugt4Q73U4CQhEmVdPSIgx0W/ybeYR
V8PeO4VOnN96rH7IqEsYLi+6mVPu7TNIzWa5u4Bn3E5F3n35xXdbz3wQdcGBHPYLuejjIrVlADfA
0kr2T8ZzxWjWch2qaNVggRRZ7cWaIMS+1yvB9MgUisAgFRruH1bQ++LyVdE+ay2zsHeFoDUWLlty
GISCvPWKexq1ClWPgpFCJVUxDxGzc+dY6EmmVNvIKhmHASIRzMPpvjGD1UNFeu0RkZhq/s+nr27r
vOAf6O4rXKyd791N46w1mPzJRHf63sSQIGHSf/SZXzRiSiO+tjb++S/viXH4L+SZ9V6ZbMK13rWt
qaUPbpKk8g2cJsyN4v9OxW6Z0rJ1lH4h+Qii43FVxXS4AsyOjwf7Ye4FSLoJHXdBfqSzroYaKxK0
4KbZRTeHPm+hp7o11C+u2TYvnva5Dxf1cqDp604fvZtyMlkszmbHISe2bVHEzbWTTvkKdQilCViv
R3uXlC5CW2tK2klAiqVbHHHJPyiKn/qfyce5q2hcI1mqNwzTEXMHXD4Q/5BDAqq6bHZ+dEzajW7y
R7RDs7pKOEChYFEWbRUslqEqiLhWmJTdxewQBhKor+D28SrUVXwRJZ7QxmYyjMrbuE8qodFGZp03
w/jqRLuuwsiDJHq0q9Qp7yY4y50+FU3B3cvrXsilXonGV+lQjewNJE7+PYRB4wb7TfZbstlyzUcG
X3h7MMO+bedDem17sOEnNyc8IRs8+fjjCMg7csDEMgW2Yd8hR5m3oxmo7r9fUIFwPSU3s6GqXJFZ
ZX+yRfnB/3lwXyIBuZpqPLJ5q8HLejDYLjFoloFhFFMGcb/xTI4B9vnHYjWpK2O41nHGze024PQU
+EomqGhTNyVC8KRu+CK1asvdgX2f2/592qZ6LrwL1rMOUowOn7mnhKpo+TvTLs6O142WaeqkHnIv
7ZZGWSFUVkUMPxqL5+rlTqGLNoL6+4czwCRgO9jDKGx7iy5Q9Vb+908O/2vcHhr6fyAq5xSlikTI
OVtXXQO2fBUTXZIv/qSuwRuxkd6vPaILHl+Ws02sX0bwkFSArp6Lf8D0I2M3GIKPZTS7VXCdWBpP
4AaWrzl5gfGNAbPwxUZrxHzNOTXO6tWe6V3xjGmCBiZ3A0R8/XTk4NwM4zZjPU1NNbozaY1j6arC
l/AEU0TxpiWR9QnBXKVOnojo3e226qFsWsnks3BPUw/GmhyUeKMqjfRi/M3zOOHcMFsfa5Ii8bWj
CCFIVO2ujrK0AyTnmEtROLrOaCG5yYC5AmK2O6snTZ1J+NmBsaOq07nYNyXz/0EWSeh3o6eEou1w
5lbMC56WkDv5QmNpJvjBz6Dv5k9kUHX13Hl62FSPbp7qZWN8C2Pwvrt8NOLZ63W7OjvKuE7Wbg/E
1KGWTuZlTll6Cxd9HtBiF/bVdywFEzA5wN8pM4uX7oL5kBPRjUmdMZpJCfyuKrs2bLN20iHfIObg
0Ek+7iLuhI0v+AMDB0eeNoFtq1SPHuXPWQXvIJefHwJ77yteDCBfOp3wHgnEja/QU0hsgz1YWqw0
vnXiIcGOQGDGnSwTXazAEmI+8cNIW40QyR6wd44YWPJhDaD+4mvxm5KXRWF+VuiT+Aw9tvUVaDhT
n8T1yw3toIRhL0wUPICMh4E495iGrRykMz3iVbP4b2Er20JBN6y/5Q6mFxSZ9M8tBeJg0rhDgV/U
/ZOu1IsjF9udOo2I8UspQX7OPUzLplEvJLQ7VGxFl9fnL1LIvtWVd2UkYnGBq2Lgq64DEc5z/0xl
HSo0sXxr1FQhMLYvVzpLcizTXXWV115L7WXzfQjpVpubSpEGfAVoy8k8boS2Iwfqi8G21RjYTE2Z
fvtA+GItKf2+t3fzbGQI/m/tP0+ZV8CArGjEjliEKR1n0KzyYB07M0ErREADLVS6i5OyUGFoQHWM
kMtM4KmX62DnD2rWlWart5PzJ9SwNoxfL6AqUW72/GNZaI+tIKjOpXMSTH685YTpK/5brdEUGGV/
fG76eO2grRIE6ZXkCrk1zoX7ggD8z6FiH6drjPex0Xj0rs2v83X6i2OscSztv4jeIyVQxruTM45Y
lbMlNPzJZdCShbF0M2+eKaZAeljaKSWh5BPtVR/7Y6TQc9vJdoznVneLj2rmmxI89Mgz/I1FNI5S
aiZLo0I0EwQppIWD7hHS3I1QH40PNZuonS8KXCTYa/5QUNWY4pu/3WukzkS5d+JAIhgDeijk4Z6b
n4DNnSbqrn2eRgHx+sldk7/Pnouf8PH+gK7llpmVLnVdGwXhfE9lY6GFuX5S+nID3ATnfmMbSTjW
y19ID/7Q0pJDEFWNmGCKaKpb74Kip5OTBb2eX0H4li79vRF05fUYGuNOUilm9Yuvb5dS+pCeZ47i
kD8IEA85wTPmZX91/IbfL3s0Z79GwxWn7vfCz66UiYpHvJAlDsa5YW2e6jIEudTvfbTvRKFLa6rk
LwUu2oKFosQW8wv+/HVFKuDL/WpiXuwbV48wC2Iythz38YRLOgrhvCvUkL+7srHWu3trRvaEALz7
Zmaje9W1kmk4UjTng74vOo+M2nVQXePJgjNBTLmtKLfO0+eNgMFvOfoOtioNEIMi/HGF9UUkEDxZ
9nULfF15SgcjyfXogcuy7M5MF1wnYwvFORkz5h0dnYYomcd9QSnRxNdrZYaqApZE1TfzsVeHWdt3
l7lfyUr5ZUDMLSeTBC2wwlOWrJFxTljczA3iE3JD1ySets9yGoXwp0hR1fpEWfbBt7LXlBeQ7DXq
RkLNa68UJNjjx79y9iF0U+dopmldUw5WkSVKFb0mSjlpOlThs8u9TuEFVtwpHPjGDfFi5Hys6I0U
rIKcQakpmnfCSet8axIOLiCr5+VTRx2iqL0sbR765HAqfvAU2+t94Kp+pqaKon1yostixDRfvbTQ
KXd2/F/9M2fbo+BrOROck4bi0stFCax8jdti9AqnfGSwiwXRR5UEP03jWWn4TgGT04HKeyAN3ZiA
/Yo4ytUcTbFGDothRsziG6ev/rUKgzo0F2UBr+wVZ6Ampf/6y1FjKAerYJZVKP1Cr5C1uTqRdRqs
aBmzR+yAw3DpSKL8P9/BTz52YEM8UJVUoFkv0Es+/pU/8lCJKbdjCMYG7jzUxo0GXS/Z8L2R2dsi
qq4nGjBKSSjsqfQwnj/o3YCV2t3GDG5XonJs1m4jwlz6kgRRsmOxe1Z7ochb4ak+E8g03AZPvlbL
a+1oc/C74ss3fPAubZuA2gXKn3ebdsh/uhwSv79zc2+ZveJnYU01MOOn43DlY60LEZMQ56rldImp
lHQihMST68MTpEIlOMmrGOvIlLlrkNa2plWceX5PxCmPnYozAEB38oxImERrCPGXGsl05Lyu49KL
Iy5P/xlB7ZfQIaBLNv9N694af67YvERx9N4ifbM68cl8bhoxGlonJLxUf06BcxSXAzE4hOyQNxWC
a81WWnJFF2J7qTGG2Dn71UOkMG67tQ7VMRSnjapt+NwJkBgOTsM69SP+kuelYlw41ClOGFB6jbse
LRK0WZR+AsHujRHxwAi5qZYlmcFNrEJsKfCOeoi9l3N55QgviHi3P3Ha9F6GSQl5zmymJgUhe2Lz
FfpjwKriuJJyi3OZWjVOH7M5Dzh0YrIMMxpnymzkeaaLn2a4dJYCOgb3NFBsfIY3otXuU6fFmDUH
f6hIVBUMyUsHsuSzLYdsB10NHQTLAj3l536ooX06ooPRZfHPy+T3SttDwKLpJ0JT8MVzSb7SyCUT
YKli2TzY5JdlKKH7AWKxaku9XN8WCREqKcZcH+4MXSQfTSYtxLt7H5xkcCYv+StJAtxlciZ8p9Mx
n3NrhEjQJFK37UC/CnXff6ax4Qew+dG+A1IMWZO0+A2GuivV1XEc96L8n/zcK7zNyZcWgM7M5tEn
dyiABKV8oVHev9FxlBFpUW2FzUbJUSQ3dVjZ1HEHupKUKLWbOC1Mu7cE42REjIvcMqpapTUFXcHt
1lj5D8SoMRLYuG7Zi93NjnfRlgYJ4nIu9GSHAqJeACf5IhteY1XA21EQALt0sa6YP1D68oTet5b2
KDfO/onpXnfQ0fUDpUGZL1IdlKDxE065obWPQ6AU/ZMf1q6kiYP1IS5URWBjlxUtqR3v5fJPEd9k
Q2J3p/N3Psccj5U+PUiKbMBahD/nhXcRFhoN+/GfYhWw5azLy6uoUC/mSchMObtnEMpkJPyivFC1
85rYhCIbOgUUSu0pnklFS8hDAmU6J/AV3GKgCgrAEkxrXj21nwHVf1MtepjVrYG3urHFCTQo5zhB
mcmxR+3JCh3I2HT25LzE3lCPz3DWDjBmY+0KGsAidztDRBFkbwZa8lMutWSQspktnz+aT9nNbfbv
ocVokQAGt2UuN27WljQ6AYHxztKEseFBcFB2PZUzk9f8aXmL3xMaslbkVaxzDN+SlmtM6dD7nCqX
3j6CV9IlVkbg0zQOn5W6a35bIFz32uogBAUdMoS8Z53h4l0tkTDHxXEFv26LnRPifCmKRoZrVZnT
nCBpiVld/YvffLZ3QOm293yd4zgEeeGEupB0rNLap2FbxPL3XBiPbqAlDXK7G5v5AZ4KMEUye4+N
jDXjs6LnMYMsQn+vc9Y3ocvPrlIDCwN6SlMe9004gdiIY8UsEE2WgN0H1OC4E7FHZyVEgiV1wrO+
q/cGUonctbyLilkMdll5XT8dfd6XiQAiJ2LNcaakYNhtkc2YxgUTiKOd9Ornn2Z24UN/o+pK335p
MYPUr8c2IW8vCbdXjbsquOj5AW5wwG04zlqzD9EIq4wGjwwcv51jhVgVTL3/FYjU1b//0O4sYqOr
4rO/iq19uWQMbc5uQDEg3tfYbFuqTLRgNP5Efl3lsmuoeDbZLUmJ6uV9cIn6YZ/7WaM6wP/gXcgT
j+QWf7Ho43Agd5EOGNJEvtbkHh131pgiCqB7daVcL5ej3ztsRKWAX2xggTPde3sWgEmy/rbZ/BLt
R6t77QgIJyWO24TzLTD6RT7yE2m6mBrCwFikV8LBEJ04w/gyhYV3iO2FNMsUCwRDx/5psjhuUYdx
GP/bfMZD3E6n+QDGPM82I/pdkyTrfVcxa3xBMXA2K+t+AvxMxreimJxsbokcP7qoo1umJa2g3YNS
0qpLFkS4CiCqrbRs7Zxe5sQ8t5DxiL5xz8YX8tjmzGQiVMXAiYoPhPzhvXUDUI5PKsEY1L2Kczk7
38ay9zkUm0cCF8n8UbUZ65sr50i9Us1qDL1g8VVOY8TIqby0Y0kO93B3dE8hUfc27Nby6BPz2MEA
itt5u5c6zqLw64VR7aOqpQdP5xMxzrIpljQA57fiLbKNqgA7GeOCvnWKa2m3SFdMi985F21mIqNS
ZlGosvOkBQbkDDYBVoF+zxCHTi+vWhjRc8Wgu5NTTXhEEA4wzas5yEo46NIZr0e2I8fEqYu1ymDB
qbTLLFEZL93OFtLE6GsNA/Ml+C9bsyrXuvbKsQoPHNIwET9MzGSZ+jlLqkkysmUZ6hE0zAfP6tVn
h1+1AW/0eJo2qjy51QDJTFOHTbYWemdvNTSZf2E7FLOg0qToyWjqQ12PSg/V/7782Cq6afugPQcI
Apxx49Hta/YFxe49x+RhoBnRU8XmuBolOvyydo8EP56pSlqJfgH7ZZ4KmPy+Zwgof76YLpZxeMwn
+lXwn6RX1U0zTwsuPbNEvfNzeZJ31IdATZke2+Vc2++PEuJANmq9VVq/WGo5K6RPNj5P6eaV8Mvm
N5d6TX4vSaEoOv250kQfd1JDYIWE/GNU08TOTDerQ9CJM4YuRxuQttqS0ku9D9Aha1BnUIfgRlRR
/2kdDu62AdV+CcshzP96eWlbdbotF+ozPuoM2Sb5L5gD8eUMHKRZKS4j+SXhEe1tXxt6eOawHamD
TApNCT8wIWO3yRWfBtSq1Km715QnfViHavuoAf3+6MZGrkVsUgtVw9x2b1WoFvYGvYxEenfanKo8
4fd2a2GaLok7qshoxJB6BP3IAlSW4Me/7RnHNBGtGlDGo28JanUV5NZ0DWk7BT3YbIuRujfRF2MF
7g9ndXCLajT0G3+X68YeqoZ2SwPkvonIoRvm2WGy9YMAnMAOWmjVshMSn/traHZPikZA85FtIWs+
QS/CluZ0XQjn2a61kukrp9tQHNepjak7aOG1oQsKgY0iWcZOWGZ3s4EMrVMJYe7B9MCwYIDT5cyq
k198HlP+HY+l0XqMIEC17qDKKU6Jr6/33Bzvz6e8g74CN/adc2uFCTPGV8aGRrnMbNOU81ez05wT
IswZMMl6fqpim1azJJgPXwMU3oczmoTDo5MYUHHmiqvA+DGc/B1gOtl1TPs81DGitBCeHYv4FfIL
cItLSTKHqHC15K+/BgEx1xYITdOjmt/hjG5rPc3EcNgFesaoV5BaNg5bT/YueTgdEHaVAIzbTpNV
2vuF9MB0d3zRPMHykBijreJH/062bstlvwAeajh3cQ4mQszodzfV0Hwm94yxW0sxWWomHUVX1L3V
KzcJwegEXIVihksMqyyfe4Fno8mKuP3jvIxbbK4FiXfK8QeE87+ZbvDYFevv/qM0b65zzzkdQkwF
cRjOshCtC9VTFbcSnNZDx88DxITQBLFuzljhymBcV11LczefkmEFwiYf95fho+t9slkNxptb7aah
qxjBMvKzlQEsQvp6AIaVBnL5nn/5m0qP34WWSQ2g6thHpbmcBcQe4Nx8kBy6GnUv1B2GOCujb5nc
YQhntd2pOOmRcTgHbxkleORXhRKsUDZjqT3VxWf1D45h1xNEJD0+EQ0Kg2BNCk5i33uz5ap4UnDX
EK6mGANQZBQqi6Qdv0N6lWQZXmX6rgYdvvHJ06wFIPVQS99HucT6Z8fGMoFEXvkBhpl5LejVR+6l
Vb5wnAJd5EbXYp7aHIlNFD1N38VaArIO/WlRSDly7R6AsYnH8Mj6hSM0klGuawq1r+GID8rNfrEB
2LyU1VrLFoUMCdDtSIRm06dMBJORQjefTfVZ/EcFLRrEpOmxGm98DReoa+NN6HJD7grRaButMUDL
ykKPoRHlIaUwLHceLksj3hQs7F1K1pcQmwYVk7TO9ba4Uf4t+uUPV+lah+ZzJuRJNL9Awimj3hMb
tuph2xufx1lr68Ed8ZmfSuKbKQmSa1v4s9QL0/cNRI+uhOaDT065JJilms7hPD1i2lhJBMg5m0AR
S4cQYLOf6SF/ML1tcBakJgFIHGfPToSvAAKSC5lZ0FMKU/+fA73ZjsVJGcgmLQOhWChOApXni51a
JdDmdrokfkkZ5xEF4ALEcaPdq9rdp25Immi+t/cdsXmjeRjCYn37UqceC2LBxdefKd7+HAS9W/CG
X/xBXJKa2PYSShakIzowMTLhfEgXxXLAl47f1uVJFt6hXWkVp/OgLI7uq+Hlb4Rf1iG9nqvHrzou
KLKHAmbhWcHL9NSVCdlhZsjGARST9UC6x15Ojgyf1yNAGP0KpnUASVCC9wbE3vT4Y0C/SNssSPlb
7XR23UI9jACrkLZZaW/OJHAjXcfhraz+efNqCVWJIgl/t/e4Yftxs7IM0OleJnF782N8kACU9mdQ
fwICtANxZNM7/BO/o01WtJf/3nVo3Dh3P9rNKmb2LpVsKiYwFq97vLxIL3lZ2Qw5ts8h0vZJzh2g
Ujgj5CtJ4cqxpqJcKYvSOFO6l5zXT2Sg4gzQTUYbNm/K2X1aMJmDgTrHTwosIhLQBWOIg+jNoBXJ
6ua0R0zD4ciUgwJQJVcTj/I5lQZMgfIpsMj/phUzXgSHDP2IU6hjMZ5q6HPHEYOX8T11igNgAEwJ
KQUu/2Y6kJAx9ney/qvgu9JUyYGZzb0D/rInvMI3Szsx+sdeDnqlEX6vnuggA7zWw7DHd7E00zru
cHxKj/p9wjxI8FYmNUNBduaXcgh+y+kyXYI5Z1NyXlJcr21k3q161ms03YAkGJaQQKOLkctSO935
molU/tBfo7GvTR8cmDLusvt5zjeAVgBOBOO4E4PqkEP9I4KSZ3CjJoeRzWxbc9QXZNdideGNvFkp
j3p70h8xKmjovyMthd2JnY0jqcwMtrgrFucJAql3uH6PB/XkZp3uUoO7VmNcs1RFOw9L5QGIHTJZ
ogXCl+nS4qX095OX7e4zRaLSdw/npiVCy3hjSjqvlYvWQsK9bEdlIrQB9bH3RwgDH4Lfk+fl1Xpk
3Ils2dkp5Pk6bPNi/rW+NdJbk7krgV+QPF+r2Yb17k/6NjCtj/7ZCsRmOQHQoKCmsEbfD34sH5R2
X4S8kGQYG+ZfNbaL+BzhzrUKqA9aq6rk5UyuspeKqg1zFo8HX4gqjSdcNH47Neqt4oNLrnqfE/2t
xzUJJXFGWjJvVMUFoVhh19NBL8PE4mvy/42UbCndfJBvLPE0cLVwoLJlnBlnqB3O+gt767+6ts4m
No9ju+IHqCCz38nIwDHBUbXbuv8fBW9VErkqJ8QaOf23JCZjbUgaupBYxoB6ohvEvuqZ8XpBoN2t
NQx6YmkDKSDyNWp/yCZz/lijOpshyM5xbFWaTZFpgJuU5Zp82rJFw/0AgXv4aIr5JjVUKS+cLStC
/zYDDXR7pz8AncKXtV2YeM07Vhbog8BoVtTKgLESFAEchIbwVbxXcXxVeaebPwyWK60R+jiQyf4C
33t5b/C5fQ1FRalkwvFE3sOjcwWehh0P70ri7iW7tl9lYBgsxCIQ/isPMfNWz77DwWe5Jd6CpUN+
QwZqs4fA1A+ep+h+RPOhuqnKUMAMShYwA0pAMSw9LNNQ9nxlu9SJ5b1uK1oUIQSnP/GU9W7bKXIw
LtCqPXMOw1mVoPbvYyvfdRihMR+exLCVYRHfAL+MbTMtYQM9Qb+eUxV8llHvykYfnnnzFE1Hsc5x
npTEpKkSY+mCKw/wrlGbThwcQ+Vva0In6U7/LuASCWAlr5xyxS82rgaypRW+yF1mwiCSHsFwrngs
BVY3Lcc2NoEKQpC6kV0RGr2w+PKlrMMTowyzqj+IRGSY90OovjqZaKA1EXtXGWBUrj0Pg60gnTYz
gUi2c3eChv3ShGCANNpBK2vLwBnGYjePsQz4Fob+4JHZz/AGhnWTDgbwlEdAQFG1PiAxILGOT0r3
JTOdMvF5+rYLqYNGDCQwghQlWrcOwWHTgC6ctvBgytqnXevTNI5qWtvPjoy+TOoXUjZo8Y2hTnDR
++wwo78vdLF9s3eeKsWk5ewaIdYQw/Y0QjV/RLtWmc9gm/IIe8UtCi9Qc88LmXu5CNC0urPczFZs
mw53npkXh7XvHUzOaGfAbv42E11YGCGQRlJs8FgS1HoW9gYIf6DARlY2e54Do1xhzO6Vi4B1uOw9
J1bEXjIpihjz1zL50XTWIPggMZJVB6Hus+zHROREsVzquZ4jz981dEtRzxK9XtZToc1hh7hndihS
8PvHYn1k53RS8FzFI4Irfnef5SI+I+4gy7KbWcA4ITmR+XDKCdOKguHyf6QE2Cxd/jxcndDgg38l
tGRtIUdVidJJUDHhxBgnP9Hngo0pu0DXvz+yzUv/7jz1HRWrfGL6qL0Z4WMuT90H3AB1wX+r4pJ1
/xouMRj1eJvIsJWE405yPyX84hfpDCX1xp90bovy7eh7y3Jd5MCYs2I2ubd4rkSNKR8KFTOIqjc2
cORjwARsKF4TVNNWXlR1refEZfxIlziVamKjoKYxyHYPlgd+a6+Culh2FHoXlasKuuySx9uHJJYE
J/HTxgV/nz06IJI62KgH+O4qc/uWQl9vmv7L9zCqVIODamEe1uJ+n4NjrS1cttm4GuJJzIYhh3Og
DPc0bP1dGbK2+v73RBseTG3d10peJavEATcwTLw0UDE9m7S88xc2a2MUbxUqVA6oe3MeWQSnjBRN
WOIrEqEw22mCm3eTFUwrcVOgcPqOOzeOWaQ8PaBqFDxPZbMkwyIhEP13AlxrH1J4f4l+lqbRsdU4
4SmQNc26Bu0q2XCV6u8KaEFuKWJAdXaa8LYyXtZNPlTP2Jim+SNgKYuD0Z65tlZpWNzodnSORGwr
wWyVsBTnRtLpDEavepvBAiX8DzPOiq3d2yA/NMkbdTTe1VHpJOLpIoKUVNNNTlH3xJGqptWKoz0B
jYtpW6kGoA1PKvNLfw1NUp8fvZnafQbjKk6FWLCKLyezAz4T+gvw+Grjh2h/tj/EKE/eawbbxnyf
e7gxNrzorKRQdIMnk9igqF8AVeFgFrXem3ay37t9EZfKGBRe5xVHVALV5bRpnyeYWE3UwOItOvhP
gsQq8ofaIPWh0QtTOVgUxXRlirkp0OWtEQKzZL9Mrc6Sl62J8x9W/+nOETLcF627KuFfZt8T8Blj
dUszCqUtnp6y8IuNIa5o4DloCKRhslIRNnGFMfFNJMJ5vXj1fJx39XbMEMReePsNU7WZPg6gsRl9
CAAyAb4iJaG0xXq50g98BjiOPqTmZXiMY+pGUC+4Hu3/7h4UnaSxWY5+U3L/PScKyAAqGi1EzF2t
p4EDVIx1S6LDv0iVq6cuXSaUUJ8b0TRZtxjqbvB1t4+70Cz9BLymgGQ4y9qqz6BDVgw3FnKKk5I1
o+izcSjBokHNR2dji6jplsq2l/HjPREGBbgZ52iKdKv9fweyrEPuM0kLglJ/NDAU8+HMrZUdou6Q
f/J/WgeHYSDxMFEWqc3YDd06bFtfzorUKVvV3Cchr6n8fGqXJAaK+0RBFl5chbWHTyWmvGmZPPUq
rW3vVtCIJ6WLlCStxfcAZLSjlF1cT7s0bgVM2Kbar/KVV0YBQ7dkbohiei1aOz3Sn24iNLx4kiIK
RhpiPHpKKXjFxl7ccqlU5sIqQe4hamg6CWUPTQJNbZ6QZ5BuOwaY/y7uX1RvVBt4YStOHwtYwY3v
cuMNclZr6R1fGLuauL/HsLokosKhzhjTjuBg/S9n5EXikKoszrRwOnjjPKkaK+bu1mnVyySQi6sv
ytpV2nWsedb/n7PSDXqUuJZwEK1Bw1Y+7B9XGUscDkpFVVj3JlXuWGQIdiSOpTbwi+to/IiXeOLW
ORpUJxeox4QGskfl/oEApAnJuxqUXRVq+XuLLNj+OVO9hMs1nftT3Su15xvwxrDvZAx5uqY//jDS
HvDWDPZxQ9qykKqY3yFTFU1ple/+K4EV5LjgkQDH757DVr1P2LfAbM5WYYnkYmtggypEZlivk9gG
gFwWVFEO0Pfxd6GXyADx94KW+vZcTfddyxHMDQ2B6A3S17oYHmcVcYbmSPfCAZSqyVG6lZVQ7JyB
5bUt7KLfSzi1KaQC/ulQSNOVPfQ8pOvf6+i0sNMcGEKzlDP3NZqksOAngCt8rRz7Y8lqopzk/izh
gG4X+Y5RfBz0zIcbSKzFBhbNPc7uAOEllhICQNbGk0WMn0ZTMm5AFB8ImI3Lhfsbno51WSsNNi+w
hoY4h11yngWG0uX1lvPX2IEaTIL+JLphbysB2KqiqVh2vQfjFIiQR0FmFFkmRs3ti7wvXaHFezmX
QNd3bw1xseEddXngsxJkIy2/bCWHyZ7q/SQZqzCmoM3TtTUvhlXrNztJoVYq43pazFOKasSMvQi9
oahCt4ehJ5tcp306Ezjf4C8p537LCjC9ltymnpj7pLI+SXJPbQ5ouN4IGvu8UPS1DRDplF3FK2HU
VqohMntlMWWoLZz1htxj9r4ihsMfmNyvM89CHxyqgm3pm2E3Uzu8iwniMcLmrPzbKDGj0evlKotW
F04L+SlfCiF6RKmcHOV8tp/0R4dObBwkBGVt010EopLdHL5zaRy/b3pCc0c6EeJDf/OB1uxoaBXg
GwfPu1XBXzSKPV1AVYsnluz4ae6vAEJTmxZng6R5KP4xO6PSRT0uRLeykrc/7srF/IEc4RUCgkhe
C23YgOdK+pr9kovAxVFSCqiebyEhU2ZHgIfvCkvK4w8W+Ok2kvTuBp4adChwm23JgArw9KAOQWgQ
Xh4ta4qm8PW8EN+tbPRgjsYoTwMyX2ZXyLmx3sUN2MQKHcSa8LxupfU+lEvFvgt/c8zBFRgZ45JU
Ha4DD2nURJxXqbPubEfm9Mjwt9Z0koTYNgSzlSMPlaPs8fH+RL0Mlk9A96BhPX/8KVCPqTWfW8rk
YEzaD84q20RuAWUyyOFT963cmXpeVIlvuaInPb7k3BCX8dn7TvkZjaRLiseyxOPuM3ILeGKB2w2Q
BbjOthYPEaxWAlp/n+TWiLWdoVDhDVUuIlCfSaT/Bo4nUCuOlZS1jEtIVyTghjTyHBoZrNQhbdoE
FEaBzoUmm0yFt29gupyokmTzlqf0ksvVkdf5TC4a0i3NWx1E+RQM/mEf5YkTmU2l4YBvllb5lSla
6YsmZVzFz0EpmlkoIGYSkEX/gQyzmYfcj1xzPKsvmdxcYfUdl+rdUIY2EMvRmIsY3deQhG6Yvuw0
O25HEGcRleVQ5AJD8x37SaADB5KJhhiUCW9787PkgfCGVJAwhPMufeLYnySDdaBF5+LUgx9b0Cul
9TlJ/E6QIIAQETmdH1KdA8dXqq3DWD8bZLcwlFQyW82Hx9xAGPCvqQr+fKmWd9GeH91m9xVsIbdq
TWLQHY0Fl9JH770QxkZdJctCFjoQ0iLoExEldZit+LaP3pmTRXSVu9z9HGyzqzJ5uQPGMJZ1xtBb
aV37CEUwMmVVXRSJjpJ42N3HAFexf6Loe1kAtpCmLwOqElEldHHMwLVZW60aJ7ijAuiMobr+7L3l
rzbRoBLU82oLE4XNzpTuc2eaGlY4WTk/EcQQHoBtySegJWOQw+MmZy+RrgS4fWzCbFdgstW1V4Dp
IwNlvKms/g7xVGy+vPzyhHjZqGOrPO28r+Dt/WrS7UGI/L+eVzG3C5y/Uavt9BnJ7Sy0jKJhXYrO
aKfG+my4zyjS6x1DGKShZLto9bVr6qyNlkC5GiR/F9BFPusXJLPL6+OWWo1InGha8OIcnrJeUP7x
QEAxaELXMRnyPnG8Cu0nRSBJ2iqXtCjTOVkvLrlRtzlqVQ6BXEEtVDbTRjBePIfPfXOOOG9N8lg/
bWC82Y2DV9DtGq+3n+OFC4z52LY/orynWlbwmjCXjcg/YWyqGi0bNmTRlP0pAvXwQzFslqyO73on
ynoRLTFgoHkEnGD/3hXA7Yk+Y3GDffQnkCPQjsOr0GLOLiHS69zWzKPQ2PFKE1wnHL2u08LHvWPw
Zc/S6QyQA1mdbxFxUVe9BiMOe5m1DhHnltnEQlGQezpa2uUl4adoGU5BGKD9NtOme2kO7oLPrAoB
Zj7M2BBtXQTS6iufUH3F78H7KcXQMRQ5uF+a0YapuVtADxuH55geLsAM/Ay/44MptmsBE0cPf60J
ktGlK872eLSY7akeWCJUQVwPDBxn21ZMvWNemafvVfuvjHrLMQDhVgdPW+cA/J9SL/SHtBxZk6/H
76Grc6HJSqpAv1RDnBelTDMwjJyOMGz07F7RLHdyGIPk6JfWqCK4rv1C6yhrMX+3TjiNtj8dvaGt
VWlIUxa7bT+/Cp12ByVti17pUbJXmFU4mA86eFVhfOOTrAQJvalFq4Sv00W6uTFDiOpqX5+LKRnK
ju0yUkF835MZtZ0LMz9uMm1yCDcr/kzJfPuOe71lGVYD2ZxXAPuZj3GxGDZXnVMb5yGvVOG33cfJ
NtUdYwazFrK9zPI68Yy+Upzg9olayUfQxRrXNIMttJOzbE4HHs/4zTcTJD1tV0pnqB36vMtkrRpM
oI0kmNsp1nyRtiVpN6MjY/igSuW4WIlTEiKC1WZ90ejWlbCOGpCLMi0b9G7fcHYjNlLuauPVQtGr
5cArMppK4lV3pEvg1Af8l+zn6p6hjVf18yKq9lwI7JTJlEjJloewJDwfAbtNJlyScwznEbmm3PaV
D0cECvIXtJbUGpCG7S0NtX+HOZxCwJfuiGWWf5coy+Fbuj9bVwrMVk/GbU4cfrTOegKCXvkwOqID
//+zbySmOYfOXDm8vZOCD5nIURqFewu769TGD1f5E1CwvQC3EjtbXxfrGUNM3A1aIWutPDXhJzdq
ztXHAN2X1mZU5KstTbB1OL4dwDqqRg+IQR1zlIEmFBnA1K4JhpvYecyabmjojJlVbngA9GiImnge
rvtYeaE1/nBCHV2HgJLz+ND7SaVlH5En875O+qVBGOD7qLi6fuMxXmHeYG14wSuT6Qy6ofEUISQb
Qk+z7TuSp85TiR0/qN414fG25N3mOS+xrAkLODYb2E2+YPpz6H38u0G6yYhorzfw/di+bYhjNXuF
YJS93sEbxKrE7PxjnDZ6q/XViFHu/KLl4Q+YNX47CA9yU1hzfDm2dYKnF9OnMronczg3OL5GP2KM
sJCeVql9yG3B5iHHuTGP2O0DEeeymkQYGCrUlXS+OLN6BzdF8hEV7envlED5ylX9aXIL+PRnwkrP
azcPCZIF5cM6gqs12q3bt17YjZurY9si9n/BNUclELEms1BTj2kRCYuLmYkEA7nJ3U3h0etsCV5G
NejxSyss7cP6IF3yCP/dKV6UJnxd1dyPIzLorTKxkUTVwJrpF62xvJH5MaBCQMxcScsPEDbOQB0X
JFC+eEGJCUvpACRatVXya7UUz2zcAkgF99Ool/Xn1NdqesdeKgkUde4YirPVLiI0Med1a5ieVo9O
SpNDmRvt/hOWSvVCm5b+GJuijSlLfQD3Vj1+b+WOCVv4JzmgEX7iBboLdXbWzNpTN5v40pl+OsJW
SI1MYcaNTOwmTymCVd9SbgtUSR0SYodn+1B2cGRq/tZMT2v5HxgnY8WcUDvYvktNGm4VzrevghJ5
FwB0bNscdGizQX5yULqyx6Ig0yreqbB3wzS0kFYxh1whShLNSZZfzHVI/pwC+o7sYCh6dZJhdZIT
1bFzfFHqN6ZLsYrPdSEJwq+tjWNYAlGUGtYvDaRFdh6tIxT2ezfrskuX5SRFZWULh8PjK7BVCEjr
ojAB2meElF0tl1rDAG77w10k/zwk89iOpL6PcvCKmtcKYdpusZ+zt7JKQY5ERcjJNEFfMxsl4GV7
9kZs3pmck0VO9RKAR9RL8fYBqNIAAl/sJtk44f1dAZldVdPmlLqpWjU8Xj5Z3lMbamOFpL0RgKRi
jgpCqovPnt+pNTSGgdrrwkCED/ufRTwwoLKPprc3KG5J7JexZBXq8Do60hgGvIfq/1ct9GAoxlwX
LfMqyxl2DwuVUVP33vYQFk5jgYJnzr3//1gjJTKUdlElKG9wlozn4v39wwQtzhMDcDCQKfZoVHW6
UYcByZx6BxbAsCGOEhZGcHX1WCbKx/aNZ/YCAkv5mLo2efLKOEf6ZrUoae9PU5G5H92T9Ung3iiT
7y1glYTr/yHDK5fahxp364/G/ERcpb0D8ErOSAcsByJyonhqoUh+JTiXmbZ3taXmUNiUwOM6lKW5
8IGY4NHHNB+kpLKk3RG9dzqBEpY+dTO8A7LKZYIAB/2TjHxaxU58zyayWw5BYfWRWFMAZHmZh1Km
uNR/Uaxahfm/4epVcKMFnnrbhzX6Nb1Mdc1SCngghsozyvR7bT/8rWbUQ4u+uIg9ojMd8sbujVog
yCO7HQWbtrquNDrHANlMhRymB2vv8+t+6BPWWLbOiPNOPxAukyq5cO+ovj6FZjhxiVb8dF6j+Oud
qvuOTDLqo7cWjD6hFbi6TT5nfHKD6+Xn5lCSYMu9PVrd0VccaVpNf+wKmFvaBKo7hNWf70xW5Yl5
5KEgs4UE+hZiSEQyU56pD5g9xKsAjTUmao3rRQBvYJXZhxvCtBIiAO/6YdUoA3pVO+g83gyUCDaO
6zb1/TsB5K0Yr5w7wl1JFTLAJW3WkK/AkGRSQulb1VhBuTbWfIflxfuNeqc15JbPIik3hzUCSt0u
0NWLbMfS9HFAj0TsA0OpwvyAmLgy3qKa8Y7gsYtdm7xFVtk+MzJHj4CfwHakN4WTOtVSfjRqqOza
qjQuyvA0i9m3KQ5LRS3g5eW0LMTrKJaXStQk1ngeCSv/qvc1/8ZOWk4G7qLTlpkLn/QrpxL+pZ8x
8qznYnibJf0gR6/Vn7bNr1Yuddp/N90rGbCLAHKvqoIb8d9OujiEzpOo9C0gcm+HKx13atFW1M4b
zey/V+KYRTGUJKgV+rkW9fPYxJfCiO0jmhg/ef6S4NxjhR4clVQ2epZmYDYlOd1p35v3eggYRlnu
7wTX4WPqlzzW6GVVe3FLPpcUxUfjm/HlIPjUOdAM8ym5jamY3QXLu1gAaFGTUSevp+54bGFt9Q9f
Gveyy8HqIhUkNxXyY/NYK4cEMqqeSRPqOk5clKmmgFS26KzaBQS0BJE5qR2pFLT+yG0cG3Rtt7sC
ws4hDGubvsmW5KjOUKQg6aWQB0ed481njzXrIayihFwG2CdsMflBUKSKt4e/AgZw2cNhu30QdfkG
BfqsWTdjclvyftfFCdm8dy3lOHjC0Uzmy1UYvZV1l1PSMmXx7Nho8GCsZtnak28253lDK4PZkg0Y
upK6QxDiqwAUUrHazDiqhnAar0/zgqmx/YeqPKTKIsVBjiZvmRJLac572khU3Ga7Tr5EZuY0CBa5
2lItZVF5gMXs7GynNS1VVHgf74VKLWOkEJjr4rT0ebI/rK2aAFU5G/H+C89ozUeM5fv6D+XBBr+e
kRqWCwpyIn2v7D9qqwhwWrSdx/R9SsQ58iLk3dAiMw32kpjHURqa4acV9X5rPqWI3BhPZ8HCVOwh
lB344t4rx1UJKlvwztY1NCCI6TmcumihN6/i56Y0OjPSkQtpYJEy1xp7x6GxmF/plWboFeSA58zy
FNaN5PE1hx46PqQSV5PopgVvNfB4EBhgui3mrFF8bCBSWhsaiM7pjAKHZUE3/tPLpEPDfaeqAs65
GHxATibbcFUJiqoIonL2Xpazu4EQGMsa43tEK/55fIEzlpi84dJ4OqVUPE36Xl/vdqpDxca+zDMA
JVruq4pp25og46fyG0qCw1iMFcYcnsGfZSISXX/EcUCGH8QEbOqgtTA+tiwJeLlfWjHV7RPM7dB6
XuVazMHTas4eAJlegYlF0LR3PNumFWqsikjkDtFtePFyx9r4IfjXSD0VlGZX0yUn+bGDbyAv2hoW
NqVhBRXwYAaTzdXtllan6n2Ed8DWSfJglcmsA7XZo61NjLF11nZe7bxVZ7XX+vc9pST+K1WEGWHD
Nr9X7IbK276H/VIMLiPBZnY6ZczmBgCsvHSXJZOqA6s/nk6+9N2jF1ID176oG8S2UIogKSqBCWTg
jJ+2m/BPXYhAj/NAlIvFOmBg9o5GNaplEnD5UarvVKm9yc4nS0IvOQEvf2Xdl8XoMYsXkiw9+89z
oUHkgkr06Vjj9MfAbbk8KlvDvZeK5glbszwsJ/nZrP9NgOVJU56YvuFByreVdsgY8zEk/mi75ncO
xDdRrfn7USC475BmaymBtYeZmjduUAHCSnIZYosYP23vkASxSkQ5pNPpVl7cjVkWtmOJ3tlCGNgT
oLRIONIKzX0/Al4XlyeQrbMoRW1ahGRGPTtuPxkFY1eOc4DobwhBebRJ+cmly8SVLyxh0W/enPn1
xZvPqXk1ZY/R/lCT/99+mQJHql9PLjajscHjDS+IUbeiMd/t4CO2MSQ61FiPbAbtPlJXx4UfGAWS
7+Aiul2e05aOmL8CkDedl5Zwad6eg/L+8CpTYf72C/H/DUOiAifmRGNlH9jE9Aiq/PFyChY7EyfK
1ZIqUvcRBqasyAvF1JFjW+/aMJU+lHs74nxUeqms2jGIFzdnSauuhMLYyTgCgEseyb4wGbXwlA85
NgnVRJYrHBsNhzljHJHJ4Uc9iWIEFwL7/DZkCRSB9TZ/et/14mHxtQk9fU/j4C/3jEdQxux//gTQ
mJQEwxCk+eI8iw03iGxTBb43dDLBfF3OFfXoulPpkxQ353ri71ItzrhjE7UQE6hLvIaFq8UiZXq6
UvvVUcQTlCJMBPgF03cyXME4sWffAAyD4lQVmd1/vC1RyjkbnsL8sLhrp/VkJkQpoWdORpVYdvEk
bYVjPv8vveluxLuYB+ShVg1qiZcJ9qntepy8W7ElaGVYtEcQTYspoUl0lie4pKdDK5XjsrGfz9Mf
wUEWe/D+wT3PJo72CPybbesZ9ESkgYkQjmz7CeWPConT06UCRJ5UkKbkcm7yogPoTcK5kbToW6t4
/MEFVwWrxj+krN1qvnYWFOmcTYPLd+r1iMHSZtoErfY4HobPQVOZRcrVEE1nuX7g7IuSdzEUIZ77
1SnSJs27cAwWPqGeZqL8JAb+7E1yLdMyzF6Hn+xTekEVo1hWiLW4VPy4YKfXCFb6nTKFbrvWpUDF
NPlYO9r8foeChny1L1XgtsMlyh4B5JjlaZ4xDP3HgJ2RL7G+4RuNO1ONTw5WEGqrz2L4sWSyDUjV
mDDD67cZ1JMTPdO6M5VG1p2LFvgGZd9RsJkTBPdMproX8VRCYLlvWQlhpK28OOl5CcENpyYSHQLq
wM50AjAetISFuWdl8+b81VmWQ2iX08taaQwipX71A+3SMskPy2KnZvg+IDRe2I8DBeG2u4ma5ATf
0yHGu++vv3k3ZHz076umEuLMP1DZiyQmsYtz/NZVBL6XHmwB0MnXsgFa/HwwcogiKramwWYmuSnn
AeClHQFcEUDfRgSlm/m2dBBX3cRo3TrFu72WVt02UWpmmJ9xqBex5+y9d8U0gV+bgxyRBlQa9OMi
OZUaI7gZiSwrMYrcB5k9YAZs81xWpMxQUg9m0++td5EwZIf4a5WIveCi/3+qIwdo6eBzR2/K2Dda
kyBdqh6mjrfZVPO9bABQ0endcsaM/JEVe2OkpK2CwgfBvyWEitEbo+FLr5Vgu9ONvMbtPeMadlXk
8NRxqIXAhu6+eNSq02mpvcHwwhe8is90J52NHaiI491MU2+scPeWPRsXmCKp6GNrVyY/Jwa9O5JX
Vs4a/XCygV+WM0Et7x/bvu3I2N4Wc2G/9U2mrlob8CkBtGgIrGHfdPieZBVUhP8k34bZS5xG8yNS
3QSSTxYzYR1cU8yi1G0ygGFja8oWsV8ogg6tX0P8EUoTtVRxxnwLITh0DYxzd+5YEbxICVMTv7KK
FMZTXdfwqbNmi2QOenstWwRIxe/HA342rlzWQ966uVAAsjQG716g+64UpYagJxZTSFixzjiEu2A9
/bT1r9uiVm3AWo1jiXyH9aj89y1IIBnA/vIRPhVPqCmIDtzG0778R4nxITTFFz2Bw+DW03qHI9Td
cVrOd8Ikm9jk0qm9cUjyAKyDw1O5zf7Ur/1OiKXY6C8xXfTOLsdUVoikMKeaNq+1DpstMa0KNuwR
2kn08fAS5b9wPcG+G7u8Fp5GkGystGW3MnGubuhBxram1M+RzmPHt1gHSWDufCnaXH9kuBXx0e4f
HvlAZVAM6OLdKr9Y3EQM6HYWJ+x7hYElg1xIGXBiEROe3yLSn1nhGRYM2cS7YYWRkWJ45xQt5UiO
iCQi0dbXqUgcKx35Le+lyGLJIX3ZKHCtwFniEAJa08D8g/CU4kIrSTVW7dQanr+yaa1UhHOqJypS
31DtUrUG8tkmnpsyBqdqfqiz9LKR2MJ/JZEAzO5GdPxneiXkQr+PJOd04Ag7P4V20/zd7ktaqT6s
i8bvoEetfpinLAVAMjXyvnjdIZ+pqmDL5fRDCGeHz7RBLJnpMyTugYmKtIqfs77Bf1krXbpYZ+4F
4sKQGT65gTUnpdMDAFrWKUQjhSv78dhlIvIEtJCF7VfAdE7VUQEempi5XgoEiv4gwpuO0c5bhXJ3
hjz1QMPC0ZPYNMqKyykURCqazxeK3poSEpS+d6zg2eUpyUHaMkx+ApT2EnPG85DAQqdcvf0DhvG1
MUQ1oNT6dcu1I6EoCKY37O+Ma9mECLMZFiZnza70ls6YS964f88eb7TAR1RNAXu5IlvuEuJqDg3p
ylDcmx0zzpw5oAu6VlzgiHh+H0pBM3WUqTMeaUa81BZ1TEGC/Idlp91KW7vjUrLOvWAQWt75zw6E
R3OhfaKrkVomTMBhtlPJZ9u01NMEHB/HdaevpFPEu238kNSW1Ht0mf5JJJOaHqXqnV8WrXLDQA1d
NY41OvU8TEf1k0kGrk8oF7YgYYTotKAPdoGYPm+bk1cxGv6rtSsa02CfzpMHCv5tqUCYVF84YLQK
XUgGp9oY4KWFQEIToR+Po3My7aHjeV+E7Kq2vCS57FFkvgVmQT4Oy+OSu/K/xPxMjRNFFtamE5Zj
AnTVapgbXs43ZOfR4HHgnw8JHLbqCFj+H/jcVi6CEO7tdRaTjB1i4DmmjB3vK47Vg7bzb0D01Bf8
oSb7E5rZLHSUzt9rz72zqXhrlxT7aYrCVeFjZQodfMMgugFSRZHItbZBsUmLFcjcTLgcNPqN/cfd
M7mzXrJjCDX6+LhuNGIhxPPyTZnv9iBzmNQhVqQX3bkxZuNDvOJFHhkUSxPvIb9rnj6j/yeMOhoJ
ukjDO/+M1vZ158MNHzV+3trlaz2xdFrfy/GrBvOAKycz01coUOwAtBAsRuOr14HKIHZaFPVaGTNx
35Cyq5GYmlsbwBzT/K31p2kDxhMoDSiMkY3Jdx799oaKIe2+ne8nZYbjko7NNk2Zgq4kOB0bhAqG
9CpOLIi7fTQdwsbNiHqAL8MdFMQvFfGlAJXTmg+EhDykYVuD3hO7ATZz8ygnnb6p7ZdUO4Yzsyye
4chKyUy1L6aXn80/lNFPWLNNAnx1M5I/EEqd9i9q9lpHRkMNe5/2X+mIrHA/AAMOJsoh3dCsT86I
vWesteF1OFREOPMJsvOZ4Zm7r5hvV5ssQgM3Zrus6Pe6uj+sWd3Fpryqh+4hn9zMWGwlxav64lbY
Km7W92mESBWLQTHFni6kTEv73BaX9aW2BoV6TFrNIEfYpizAH+OwYeYYhv6HXZVWEbwlzhVbMENH
PLfmXGAOpumSVmfx+sEtPMic1ht2zq7u+e8ZWAjKsTIMUut1SPGE5+IhvmIYnCtbgQrcdTgGEPGo
9dQ3/6hWRwULPBdjTfpyKbfHS75ty0mZNgye3pezDOj4/sPc6U8+Pa6bGKr+J+HW+MlxoP7Js1D1
pEkfW7HeKBj5V3u39DJAUUa9hrznWSFP+pss1zAsg/gAVmzN6tmC5EJ6UEaQBqZGGudSqETE/PQM
/45tAs39l/DGJlGMUuVvei8cU80xLQMkYND5tJjltpV2cL+Ae83oiKpYtGGSLtLNA6mwTzsj6r6O
HYZauQYTRrm2v4xsBEC0uWPKDxjQbJLqwM9Pjt9UA3UlciqwZ36qfKIjwjz/FLsR2x5+zACJbtEn
h7tk8WA5Bw6Na2yawBFVV/B8j+3C16hq1sdpGM8gfOhaY5ULg4xMN7ehjHpkN+sc6uECn9tmP1hT
+utVHU+LUGrO9K346p+uTY90pgBmSdTqgnRgf8hUb/Qi2Rb9+uVNGqhI5w9aVXsuqDY+ExZ4jOeY
VLNS+cDDRZGxVSQZvoE+b43ZcQL26nvgqVb0JpmXk0aXzkv6wNTReoiDpeKN/mp7N/9u9LmAt/oB
S40pAOeIwBIYEwokDSgxMaDZFLwus9INr7V7sGf5LGk1ZLO5qEdfHVoMh2T46+am/3Jz403XDc91
iNzAblNsArwNQBlwvhhJ/R0FYZG7dXZDli9hGVpxw2RQ3AM+aEE8iOBWiq+In/VVmVMi5BfqA9tO
u+g3U4JIKQv1Em38xD3U5o0aIkoqxcouy/97J3oimT0C60O2xmtzJfzKJ/3GVImY+0UVj7q6ixuu
blniF8CWrMJJTu6/Hl2v4NH5aPYhLMkIr1aGgU5zzoFiNXDe8s0OXHluIZjgfryXahhQ5Yd5sO51
ajVgWCjNFU2UgoAXf71etVQu9dcD5MsGfDWyuEi0oBgqCXO74m0zgiTKbYfgNra6zE/JD8h1MAOQ
TeI7ktPE8nX5s5UDUu0qDaB1UkpMH5R/t6w0E7tX1KnOeEu+kw0ZqdhPvcBzahiZUZgAUiU7d+Vz
unxYoIntQdcBkyzIcfVFPYst9UgAn199Vpqdr3qcYvDEW/Am55lnWr9DNh+Ymxg3bxpKAh/ozLeh
2SdneOWPoNfIA44TxMuDeSuBKRafEwhzolPwx7/gD/NuOk2F3p4OelIIO0ZWnyKHaW6jVfT15hvH
sNiG46xZckOwui2+UiJzOfEUXl5mfS+GS/lPxcgmSFRkFDLW4BVNom6tVPG0yEccor8bfd1p40yQ
Rin4CZPYXdjAV46NqPPS4sg0Mdb3bZLeMqdTuLeMz5MMk2KaIXIZ2fKyWd1SMdeqlC6LbFaomNKS
JYZ2uTCUeY/qdScdwF8JU2fRdEYQGwxAtElgFn9cha9Tp6QstMpW1jVszw125KEbFdHbSuHSn6W6
w7YQcoRMMzhq64QNnPk15aMUyPKAx/zANRfYrFJ5g14hNNJ1EmyIUxIcj2hAazJjVix67UaO9us/
6eaOSbwW80ux1Nhloaqs4MJFcR/b7yGHJ1S1VNr6G80F6LudoChT44VhmK9+KCYztWlDgmXBsdcK
2+55xKaUJyRejHzKDOymrm+RQ+hOlPrMwjlcMCdxvOwoaaY5F3X0mW1HC+/XA6mVn5L6MlEhby+m
jw4mSlfFZSeUlXcNIxUhDKjRiJjbuJxS4JYeqK5OnJvUpHnaZNqVpwUtaZEKn0vMmvDbN3Z4l9xx
eBxDDupY8IrGvlzUdmRu5sM4uHj+s0zq356LEOLqet648syYz1Vn/+7JYiTs+FXKdYOd4lohvj+o
D09rXMAE7JFys8AbrL57f3yWyjWr9D9jKKiLcTGcmB6LnFujn3bdGpoCcC2T/g7LSAQMrQQ3MRN2
ZjkbWiOl+EAgpotqoMlWqJY3fgNTMwhJeuQz8GwMlTXRBH6kcAnnhb+xYTFfERI4OMXrFmX3xbo2
zUPoSKwKPLF9Em9yhh741wRvrkwnxzcjZpTeX76gRckoFt49AzTDh/lw/hAy5Kv3RwkHzDKHm2/B
xPawuTJ1ZspKJHS+dIHGLkcAySKtxjr4nQ+Xp4cTlZgQ/79AFb9dQ5rhLjUXPrGU9TX+VV+0riOT
gZSIFQY+HaxAe4zlSBYyHjEEnvgkTPapTdM+GOmXw31UVpkdfDxCuVfw56QTxhaNM/ttiY5S52ni
PaQpPL6cfhCirpxdInPRfnendDo6nvvjqN2ifEgTx5v69zq3bvum4L/VSccHdlGvw+q0QO+UtdtQ
WUzf0DVcgXbNs7lBFCG3nVV5AN5s+7EW+G2ckkUO5aeZKWOGqkpY43Kp7kZ2WRsFN2IIlwoEZFeO
asSqT1hPfEbmDZRMGA1qdClmHPS0zTCbbw4NFrroadiorMYt6ny7jynWq1s3JEcvA62C/c9B9Qt7
VuE+B9CdV0qauW3EF0QtSIn4efB7YOJfSHrnZPB4LfBf2nXnMx7Q7xWDWDf71XkQI7Se1/W8ErFI
DXBmvjGJpj5hiDOnQJRoFePRXZtpHyfYXnQVU0fzR/h9lQx9776Cfas6Iha4/z1sBQiPQArYf7w0
Z8OnFT+rt0v1iStcYtwRbtO7Fm2mPjJfnRgywFFG1X4qe9SC6uKc9a17Hg1kKJWsXKjgl/GxQOAa
m/gTM9OIWLk454Zef0vB0b6N8h/4yEtIVlfbU2/YPjfUIuc54GS6pCFXGT+7mYFm+JFe8r6ejDex
bn3H3xEaZH8NIagtLVvecje7cFui0G4RYT28sEawGt32n5/r8zs/27vUYH0OyNGIi4vcJ6SVZkr7
qHTuvkZt6gRJNPPun/QzDdaXfvoebSSa9Dn/9DcyejKwTpcKuDQH/OuhH+KF6ThzOfiOE1zrw19u
CPzNkebEI20Pu6WsPl1CMzQTpf/MpqnQHedk4ZoxxVuqn3w942QqcsjhBfcjepBgZ8HGwrCjV5Pd
2WkhvWOVjtLezckXSSOyiDKdsl6O5BtYbh/yy0cBAfBlTq/NTcsVp3Wyw2IzyYUsTfuqsxJqRHf5
319h7YZvim46DJrpNKWTOzL23bylxhe1ybR+XOShzEbgf6Uak5ZTfcWBdORIKaxSD4BfwzZ40kxe
cpfIJsu0LO7iijhsY+iKez2mrIS1byvAH8LGNINA9f5tlLWdXUzL5PkPG0xmtIUe/J2/AG86bgzU
48kppZFdXZh8FWbSEsiYelmJ3KExzD0CCJa8ZxnmGXR+jzVlP076mU8go691vCDbA/qrhFDRB4hx
V2NRRE1Km3tVBP/sYU+yLTa85VbFNRx75jN2uwogwN1OoYO1BqRkfFTUP/XZOc616H9rRWnqJNUE
Gc0fcmt4M6GcqjHR7GVyyzvPToLFZEFYbAMxp/Ijk6+iOxpRVRw6nfByjd237HhtrSHxfOpS4AfF
tUekeQA23vZNMp2ANovNASXWrm518/JPKTIJPf75FVjvBMv+WKzLnN10QwSJIVnhxrCRP47vA7fK
iFAg8bYWSHDH3PSC/aJjdcx34OBC5M4inWFKojAgi5Y3VI8sJCTu2AUApHg3x9TnbPcVl2f9o87c
0ZOJ1vQLOQ+oesWV8qHJgmCEOXJ7bpEv9mQ6ExheoMfvq5NoteoH8c5p/qcj1UeeltH+TWIGWX9A
srP+hWR49AWAJ2R/k8VLiJwOxkNqD9y8jE2+WYdkntkXrskgRxzqCqUIsv3roOBDpWUKremmpMwC
ou/HrJYL5iyQQb5kt7OEOxjCEkNCGy6wbwi/uUzdAhBqURDdcu8Fvd9AFIbvWJ2wATPTeTd4E+kk
d2lvDXcCzco5yN4JgHEAHCZBUXOEMB5Ez4/Oh09mMOBmBrDP5mAiIa+S9CmPQTkI+yRCibn4ttwn
RMlqM8b4aMYiHGGDwWeJ9nswzfiUCGxGbBOBf76Uu/psYRZe7TW6A8WkiuMIS/a6x8gODK3vOI3M
2dNz51sYxlf48FnqAhsgC+0PP5Z3hQ+d1a8Gv6MSSD7skTgcMZzncOXVFSvT0/I+RbjMjt9JB1yT
znr11M1q/a8BMq9tmIRpCjyd91YF37l+NC3c6OTNNHFzcPxZil6nPi6ltc/IBo7iWXekkASQBvfU
9eS5nADK7mZ8Q6GK8/iCBwgrqU87yobPMyjfIfUgKaPgE+j1583Ca/t6oOowa7+hEGBVSchFnX+x
aF4KPXWRBSu11uUUJs6WjvM1awQEBWY7LpEwkqN+uFFNMUHy7TPBE6cC4QwlvJzJZY58iQrZQ5uo
YCYYfA3SDqvN0wiW4NA1gnelKIpWYL6H9Sr4S2ViaG76l8ZCW+v4BqI8fELTWjqh83w0P3O3blJM
KXg8+SsvfaZ7iFc5TGpB6gSJFcUBcxszhiJrOwdHR38ZnGhMp4xz1q93H6yLJiobgGkWMxiCHVUK
2Y39+qUORxGMdCNFusqlDN6T8VpudBHxMKB/bmXusXgYEtRTETtx1/5eY2nunMzvUoX+NikTOLbV
hQduIVXCf9T52RtKV/RHTlmgB53IBRbe7qY3sgXZWPM6hgaiUdWd/pjh9AA6+W5Xal09rKhsB+GE
2BqX0jVKxnPrLWQwDPGoFkTcNeJ8HgiNOoIFSqAgcN8GzN8NeiUfPAAgHWrcxuuYmOu8DjVFr44d
s6JKqtE57lcTZdvAtpjG2/puFUd1r25x7CaYu04erB3gcsJwXbRCsbzf1cY0fQ31XEcRdzBmO0gR
+gbjkHf+qiXF37j5Wnucy9Tc00MfBqOCucsQlwK6VVsIYsrRjrJmCJWD4d2IKxYbf4oHpxlqebMZ
OHEgMauohCDJqSi/ojTcf6PZdMHZbIs0om67N3V6+CfvA5zMQzCROBf/h27JGjnSLQcwbFKA0dMy
/l6sDmB1usALRuHegC4Kr2S9N/HmOe1DleI6oIF+kTg0kqQ86M/XZ7b0lHq8Zvj5h1g32TuPAhP9
jwu2tAcztBommFbinvoZUYwnKmomCPsbBLWjFOMDR22xvlhbweUysqSpWwMdzuWEw8+vNfxmVmew
HxoD25NPoTBfYlRgT2Zp7EZl0ijH5FCvt/2DEtz2qfFaWkmBNft7Z/8Bl6NdoWXL6wq1JoxNE9+w
wQD+Ke8o450fR/A2NjaeIzM3xNwtW990dkFHHFjM19LsDL5MM2KqQrYGpiuPqFidPxxWL9RSQkaY
YK8rQDbMyCBe/Jd66Ii/bDlvsAL96SwcSilR4TzkzEFmVaiU0yiHqjutof5lz4vF2HxDcOHJ+YCQ
uSii6F4sTb6ECBfX07XAaxSKwzmnFBeGP45UjC/zJ0Ox9IgWhXA/VSEmZ8suk27EQFayXSG7tZaZ
qzrgq84k9aW3H1mEKwEQ+yeLNPPVAc+7LOSF2nl46JDRBViJB8OMYoP6I+6oF5OGSKD89z3bwnlD
QtOFsljf0yJ6+VnlXE8ki8E6Tn3fSHrxv4/8ku0k6TlxR/ZFL90Bq+Qv8tt2iFUGHL3tL3HD7Qm1
7miRZRNPDv4EmDwYwUyJypOpjFyEqsWjHhkxqa3cycNbsiqQGBmWU/53soz07Tf4Fj/2PJjNdCMQ
jaPH0/CmMVhoKbC90h9JbXYAOrq2f+I6MbPg/YIgus7CsRSXZJovgz4/j/itoIPkl77ZUeXhsW8K
RTuh2Gupimxa/kWTB80G2Hp5f6kydaI1pSSavzgUH1H3ASPIn1VnL++yMNbkCjVUC4sQJdJiVWua
+6C4XfZpeWWYGZ73H0QfGNK6ehmYhhu87/19jMSkTA/J3N2vcY1gsx7Z/Hx1FS/qb6Tla+ZrQTlo
ZZPVjWWUYRWxy0N0pMgrXKfXW15tjaenvu6QwI5dRRsEbyLX9gujwtcmLMtZilAJnMpwNVVKdBb3
cbEWvt8RBDLltlR+iqPTwr3xrH07cFnBN6LJG2X86tir7k/ivUvUZCxDgi/tzMJLbtXxWcZIiCB3
42FcQNK9PuH+SmU02sFGxDvf2gAb16W0p2DIteDhoV5PA8jQnkMjTbQ2gFsuNa46mgl4HHMf1mTX
a2Oi3prMrHr+BIi8fuG0eCw9HAyzbyiFKe6eNqZ5F5G1LdBcDHNJyGREsFtLIqJmn0F89dyw7/LO
7vEF4Hrp0MP9ZU/b/xd+Ne9pbrVmcTFaNPAc3oy7R6nkonMVkK/5UikACK/qXzQur0SbPO2FNzIn
VPA1mAcCa5zllx4cZa4HPoJQ22XDZZo5sOJtP5BGbdbxxcgtv6LK7HVcyihgLvaiYEvgrn7k5xGo
likF/0JlpAB2IQzUwECsZdVJgEjUq64FAOErZLMkR30tpyt5LHsCRCkkRTpTvIGJTANWwLAlQAsW
mthS7/EXFddwNsgGFOogKbnulCxfRocXG09E1bY4BQxZMugJNBMZ42k+7AB/z+64m0zV4zU+gzzA
2m2F6InwXy9GHNLzuZrjs6PeoAN1//ia1OIwmIlmilweSLyQUyX4trOht9j/syeXKJh8z12C8m5b
7fRhU+v9WJUfuW3DOiOjbR7ezByGIvcyKPUuFnTBNAyaTiTFNUfPazUp48XYIKVqOG043u090V3M
TzSvv0vEDQP6Le6dhPzRnyAnE7e2UZIbofGo6djd5a8J1m8jYlA7Q8nlvGmh3/1UNPu3nM2GZvzJ
I5xKYh5S4CML+E8u8w4rZ/ZlESBJZ4ujVDFeEP80MC/OInt5xSOJkj8TyFpzEuYKqDhQA3u7aZCb
LMmcqG37c5gA37pXmzjf43KS6Ko9y75iAo1fgIwU/kGDXbH+tY8cN6fCG9hOk074Uuk20laACb4o
IJLdwxUtBCnYMRYxiaB9s1rg2w9+UrSusJ02TRhftTCSKSwkIVU2Z0m3Rek47BHgVJBdVDoSsf6F
5uojWQWL7P3H7AP4qP9nOHGO5I5mWRfgrZMa8GF4LU9Pv7t7PptIpzI8OsYXbK/lTX4VbR5f9lm1
MgmmtXX3KuP+f6eJULWXT62W2pcCcpvs0qv474OmIQZyb/6Da9RwaPMY1363PZFoXBC5IL5190sT
TENSll3n1ahRYtXFGQX++5DOusA/zjXG7rb8DwSsBLB4mCEYVCMhmKFpSJ88CuBuiujVUFPEkMWz
zvx6Fc4/CcspZBN3R4ck3MzbeeHEwDjrx1OpHlFpgWSl5IwptfkW6mz0+HDTTefkKf+ND9U9+0e5
1xyDTTRiF9VtNrb5HrET44TN7SwfSEZgWoRMeI7LOT6j4hopvBgFSBZTilGNsl0e+aUvvDb3KM5v
l1O7wWe90MCtP4d63c8qyZqGVghPtCNzhG1w0fZ8g/q/MsCFmOVxQH250XRWmv7RuWRxgAl8Ymxg
SbwOL3JCGjNlggnIsCwQChEfhGaemPOAxT3YbwWNk8vP4bCuiWuWOrst84NAetCTH7UJaXLKQD2j
cP4bk7OABHk4K3wEOj1W96G7w5iTdhqVyM/KpHzjLbHRVr8mDmvD9zTrjNcmh/HXEXlZ7Fx3f9Zf
cG7qbEjzIV6kcMFzmC+3+KXrzOjiG8k+8BgfzhEz4hHiScDiIxy1Ee1jXrWTlBh7bjikRUYNcw36
uSXXlJC79SQk3te0OQUPqpMqtjufbBywIaB1scZ9t43ycmHt/l4hurzYek1TsNjdMnfPx6gAANt3
lcqPuMSqAo/bS10R8kWxW0IRMlnKosWBPkkiYMyO+WQTjxMo8KUch0WVoZqiE7J6eltvk53Kzj+S
UETtLpDFIfgmUapb+W/34ZzDwB6ytuiSukIlEDIxF4T8xVC31RCtY66tSALO721zRc05f2YWOLmL
Teu+Srl5UZkvKe0TllUqEdIFmVVK0gO784CMcrq9lp+m17iMKzEL0+YssYLasr9i1a6L8TyEsTK1
vaQfegOQTZ2w9CK2ZdLEGhzerTVYkE30Sa6FWNi6XBE1+aKGMM/qA/E4VXNoSbIVPIkOsZQblEGr
Zatizi++c5uESx0XW/ylAIxjd5Wo17xCaqQwDsvB2YEmOfMFaBfp4tygT7CTD2toNwVncyyHxqWN
8mtjmkK3rFQnLUJtmL9YPsKJNgvqi+nWgXFP4xuu0WxzkPFvFdXCQegR2KKFZYJMv4DV7zdHLGna
zsYvXzbO3PHm7aTiuQ2jRYzZI8VD6LISqpQ7q6fPQPi48QJgkJhmaQ5N8To4VDiejy/PuwkKqFgG
FxDrizYf4wCOYtmrMuUt1KxO8lMLt5PkpPeoiJBFQk5stMKT3A0zcprbZAdekFOEPKz1hlZV+8TV
dLEKCXbrZOm2qQLSmzPyoDA8zKOTb+vN9MMRDRlSjSGD11DSm+wR5j5y7a77/0PopfjZXrummK+h
BCxoNwfDbP83d2sOeXSBWl3N/h2SZZMLvH6kAaRBjaNq2EwTsTttFC9fvOayYxCBQOtsNP0vw1lp
3y5+Z7V9eWfCDxlnEReKKgx+FNWbuFH62x5Yu0sB+HmGL3SuZynFDEBO+GkyKOs1JHXvDYtZkCRa
btqypA7Nv8IA5oKemDbSysoZVoFXLTJJ3sicwnisaoTZBvOGsqu2+Hyyp71S736ZLflV2/sqtqzM
FDHajroonryoahQG0hnKMb24OXjUD6ah/+Y6uaY/mCs+077J+1hTn5mxph7GamGIa6ZJTxH7uywg
P1c0ifV/t6zhiBqe+3FT7pr1FMGO+dXbKYAIvvcXetWFUanjxLCcahHUYqqqq9Ji0iDapKjZv+HO
bqFU2vO7UnBfOFsnPIe2Zxbpz4Pe8g+VMcuZQ8r5DWAPRL8x/9jP3Z0SxVt98VFmihDDqYgO5pN9
Vh8kfSk9z6s2Z8eqQBsD+BfwCrSohzAXCTqgXg9OayXg20Mz1HPfCZRrbTKM1Eg9kI+LY0U3K2WJ
fHGSvouoRPOAY+jpqLYBr6z446KAujNUyT02WiXdQZgj4LXjb1661GPf6gYW8QgslYytmHIqlZTU
+TqPcA8QQbSXz1Z6y/GUYb7xz411kw1aD8ebfDus8+vH1ra7FsZ3o4l8i2+516uW+gyg5p/GN3z3
w68pFSQYDwhP3TNRn6oIO2NWP1z6VxABMt/ZkEb33u79rzXdM6N3QppRRthLJNo8uvXySOT0smRw
Ot1PkGmhzlCmUsnOKBcwbVcAWlLOB7MkEkvUdj8Ud3OGimYIn2JwYC1tvlyp4T0EYUlD9Sl9Ds94
aDmDCNOYt1dRex0FTklFxI1ZBFnSNRb1gM7J5/9ZOE3VJUznAbJZfBdDDkc+wRiZJDmspCef5EM+
2psmppAvcJxPH+8ilPr3FdlkZ/qqZ58uyEtYj2fOTS9m/YEb8vMU0htBsudIPNqE8G9OJFjg09SK
kkGXx1+9udLhoLoJOQWiTUOpvs9m7SqG8qb/UGgBHJk8buA+OV97s9K9UZDnpZfOfyEZwA+WzNxv
xHOPi+6Piz+FmqN6V4KfBMHcFDm307VdKV9BfzAQJCfv4z87Evkjy9ICilare3ocH8cOljNWl/mq
XkvS2FOS6IHIpibzHTxn3CEFKgnCHDenH70riCzirEF/vTYpbUMKYDguWAhHx2WhhiOJQnIzp3F+
DrgCr4HDGo3LxNCsp3P8JsbYq6fwdeDSIKkoaYFec9mjguS8kbmDLrZDzEYe5ytz9OXgJSBQufvg
/ZoUbB025YEcNx7xY2pOftpJpoHSIdnRmpThXRqQCO7+aV9JDMlwNYHcf3n2J84n4F1LcACVXD/s
lg694V2c1EcF3VQXffpCuJ1A0ywhbBSed/UBmhkRxNOteST+CkByhB+cfPp9GTRy1DKOreCHA6mK
FfpaVk3rnumSqNPEg/D8fED5jVmQ/H47ggUqkiniClxGFsgO7/bAvwyYFQGXVn5HgABe8Uc4r/KA
jzSDNPkhJWlN1FEbyJlimtsUG5zz6L04IZHK6N5QZ0XOWrwXlLxzowVAVG9neEEma72UCNIOAWIQ
4r091ThGZjAclWI5FRYH3MVP25Nk4Sgiz689rOog+F2pR0oVlNzyN1uD3Q/OlfEWccCfNN7t/PIK
4Z9EJRzR2RFtVs5qqP1821R1NvzvQOk8atd+qeyJyU+s7wvpvqxkTniIU8SALEq5e/ZH4cCcjTyt
g3EhKBfw9TObk1S8H8X3+rOkYUNik0eliq2c9glsHpu/WKYGXp85E3Sv8o9Zx/CLj8mfzby0/rmU
+Wy1SA1Bja1dBGesVVM+hqZ6P2PifHkT88raEwkuZaEVhoL5eZk02BwMbgIWW/+DB3sQySBP8Ra6
D5aef0EfRqbkRJzuXfhqw7lL6JI+KAsaR0xz4iqK2gf/0qoQXVQn+VBGvUJM9aRarPbbuU1Do/cn
KajEdcCoNyL8yAe6LDqwyzc+H7HfHtnKTJtqVQB9MEhPAG7cMQTsBCK7NxWZszeQLT1TKmphxTYv
ygJTIqcZEwYO/fvEWSCVohaO8HC8RlnKyWyKEq38vwIJxgpospd02eO4oQt4w+zlCqXEye5MVtpu
Yzeg8drmvl2qXxSApBESpt5aohK+Ud50PPR20rfohL9ANc4vCVRfj2i4bx6WgIGerJ6fZ/0Vgt3N
Cr1c6a5wQ+2gmicDwJRmWpYnXeL2n/t7rphwGnJk02kNIncne/DKI8z6QRskAKEE3IFdn/fgcFLW
thJzvIVjKKf6qm7BS5hNznqrDW1U2SKPnjsqRLpsit3Nlzeb/rjrzwPGTL7V+fhjM/5vczULFzwE
+NLfcFxSb4UJ8zxLvjyW1sEOl1NeuD+qVPCzGGhMVCd8Q5yo45+2NRJzqVts0QNXLbHwSeU0MCVl
l2jKUt6FSVEiTTE5oD67P7jNZW07G7NAnVdcjdaBeOLUsYNpn35To+uQrM+W4q6RO1DkjtYxqPQa
NQu3u4qiADBXtDMzmtgdlORQlalQlziSayAdY/rv2227mm/fdtN2miIeBXap5Rq83gogvWqpMJTk
LjRTN83+IwqpgjyKZRoFhRp/ADuUv8ulmGvwBpeMggzJjaseAkKgW3AawgYZQvwbd3d9JWHMRxCG
pJpqflO003RKQJ4U8DZng8oVO7MKGb4NSz2bHVB6q/+7ZFoi5q/fjCboz93rcI1NJ3F9sXrfzjDN
MRq1hUQ6+RfwvcqO3g9EKpDoZgICdRCW9LJBJE25tuIWydZvtLXX5zjdgzRbTgzlOzglN557gvyj
VTcZNpx5oU4uSY2S9RLYY9XaG9KUAwrRbfjlLcwrKGw/w9gJEkRZDkaE85aY8Duu0iTbJWgeLURL
jbc0b9ewU2lPI2diDkv0PwGDUCttZ2OUiGpxH4P4JH2MtyluDAKU3qtm+CirNQjhSdp0lJIbQo24
jKJDO0jo/035S+I+OwVflKmQxo5SmEbn4o6Pu4y/qbz4GK21d+M42ZFnfPX8QuwpGb5G4zZ6nNhA
wZdRShUuivY2SsKM2tPFLoKvbcVv5TKbrP4VEsqRmyNK7wg6Qgw+9mPX1OmNN1vSCev/tsSvYGqq
XycQO+wB+9tpUQ5fdt+ZaJ6eLfHzQqO+OcfrC4VYqOdP5Rm6gANv1uaOHAOtH8+ww559h3tMtWSg
Y0Qwoo1B7nHzyrFJJVFwUHXRD5HQOL47AaMlt1wJwfXb09I6PKyIpLSW4azxFniTrvzfR0OdxjwT
2d7mIA2mxHcp1HR31T5RFgj2iGMnpIbycuD98vHw1cHnrZWUY/LvxpojWGWFgVnfcNcRJFhzqh/F
PgZD9SaQwAvlNmwuyB84roT45eS1sgUu+Pttn8OrYbMdZDmuX3UW66pNgk5w4cwk/RJGbeNmO5N7
b6mvKNPI9aDjn0zlP1X6ZTLKf37SJx4P+k+zqL2fmOiS1dKB4VG5ZzgAmKgMKKhH95dOwXqBkgrs
G+68NVBGLaSK+W7hdjKTLOQ2ZgJZNrexvg5atGBSw0DMG9oYh9V2OQnRLTM3yghznHmvAz2d+6vV
Wr1IBda6Y4Fh85FGvd8A2AYEYjpoKRD7i+uVGWVpqSI3sCYin1Qdvmv5l7q9/IBtHbGXYNfA0fRX
+Wi5A1jRweMA7YmzzTb+wGzsDiNBDRx1iFn0p3w9CjwiV0v0ubhSIDnrlhcZfFDZFclfI1S9zmKU
1MU5q/d8xaqFW/DU3N+quxUTFS9P+t5emq5lMr8qLnctJAgCvzCYH551MIldcYOYFnR/4s4PFXBm
yiKkxpc4AE0eLMzxKLTbB4XonMOq1wLTBT4QVpc6LdpfvmSvd+qmqiorjKZ1XS81dh3Coh6B6FIf
LJipofVeDAlOQh303rTCETRGv2Jd1c//MB00wzHQXO5K3k0ibV2Bq1IcQbEbbo0seP7hdtU1CcNO
22pzHAjlY7q2PCy3ro2b6gTjPVCcHjH0Ip0n8H/7Sbd2N5y9UxF0YKsOXEAJ+ThePDbv1+f0BEXD
z49lVN7KqpyPj2m3/XUpypKGlmYFSrk9yxrmVMyqZRxV+ZRuoyNLMCuedqF3gj3kcFgeSq3pDVvB
MaH9FGGyvmJQ9Zxn9SRuuchByi0SIQi01Mo8N7nU35vrdrjcLIvZdmBvJs98TBhMds2v1zONBWww
TO82K6LUUdY1mCrd/XN/Qeg93RhzCxFQjUwjgDpCtEO3anP6tYhYuMpcE0BwPFq2ezlLF9rNBkwm
BOqTze/yicJpmGo+aho0sVeZC2l0UWfjAfmHi1Kj75mTrK01xfrwe4g3ewS9lZDm9DokO86htIOT
9f3NHxjkXs6jCOx8OTajOGah5zL7gqAoFkC2kjjfFljxwpWnfea/d3URVHeB5Cjy+tOTfHx42GlT
Qwk6r4nocBLf4SUcS+Jd0dkHJXMcKrvBa8WkVH5ZF2Qg0QrFciQd8DbprQaFxpe1mxA/0wNeA8g0
gxLOP3rPSLUwsFA2z6LPisqylSWYm+smEMcvGksp5wBYFNeo/Jq+nrZZdcAwOhnMsTjoWT6gzNDJ
kku5AJ8JwPjmwQyfc5PCHMcIdbGrXKNIETtSnZO03X8H1JxqfpT/e7AgtuiHAIp+gN4UNs9Y8Znk
ylqYnmcCpxR+znIID5BSWGKSfYrz27eX7DaVTWoKESvu9bArm42G+FJ7h2Cssm6w7Uc3dy2M/snW
OeK6x7pyhqh0UtJkgL0PIEm9Gc7a1k2i6VM5CJxsWRvsZ2CHNDe8ApASnrNjkv4szj+l5PThyjL1
xpfqqAShD3YB/IzFL4bBuf7qsTrV8LOGp6UbepWp67nA8iZ3oUMHuGVuUjttIocb0xAyS7CRFRAa
jsbL/PRQXvrmtpFQJPS22haE1SV85+Ty5RJDQI/u1s7x6kG9KxIXz97JD9Zau9PNI4/95UqR50rX
O0oq7TCxbO6deweIgn9dayJ8fuXdEwMQ8A+Ig1EL8WbeMjKiR/B5CcjXfmtCkTKbVVZJCThvbm4m
01CfZvSCN3IODyt4PREX/GSaWYSnef/QVPHQ2mw97+UovC/YzQObtq8VzGS7vOp0w+4XJ4uyRbar
jeMnjGtWTTTT9xhhYGyJ+FNMLSgt9uPmrOMuE90ojlNx29tuRBgi7BOwvrtb7xxDZVTWfrnQD6f3
cmjX7oyz7NtGXmoDe9AImjI7jMMh4z7f/6+df+fyp/vEqn1oK2VWIhw4PtzFg+5xRqM+9EYNq1w5
AZ6kEMitGU30uYi6f9C0WFZOw1fanupOAb4XXUmWXohOUHFbodImNJTjIv6eNmGYFeMbuDpWlflO
EOGby73Yi2kMbwKVEe7wZWXo5ZINvx8F8HAUMfB1kidouwFpzRQCNMwPAT+8o1y6AXXYAvBBjhnH
/hSCwuOkePtdoDi6bSCtOp0ywGVO6DaxXPEiEvQrJIyOEXfLDcNVjdEav7/u3kDDPlfUVo7ItHnt
dwqEFh6zHRVGt9K6tsSBkQKQLeTctEM6KumFxF24ga5sTQTEqSp5w9eZUXaR1Wypt0/M3bS7SJn1
mN6HRa882Q0aLhQOTXU/ryRaoacHEbl6Z46s0RxtIlWpuacjnm+DvPI4eWmp+TIpHoPImF18lWKs
b9+D93HCQieJt1GWWXgBO19c6vpN62AFYhu9ea5kOWxurqrZK4Jh2goP06rJZGOoO6Jly2xS8v3F
1O2pWPJGVDKyLcSynpTxOaMAohCtcVTv8qUiuw3yZBtG2zEGTfFqTq1yd4s8C2VGYBcEkYE+1g2q
GecRcUp7EvLSKaMhcBub+zTtfcSCo33mhcxskCaXeOvRIUTPb1AqAYin5EoeMjVLEDHAB5DmP3it
A8iTSCB5rFF3TUzlJ/CTPyhSHqoyfeJXtWu6KwbdQU6whZECcMiM43a9pPZ06HsPz/ZGz9YrKVYx
OUQivsG0cgbyDWf7JD1/Pxrezyza37vI3UoNL0weZcZye9qlR1PSt5eS/fcRliNsK0pb3W4BPXEW
3Vx3ll4+FbgeODU1Et4mWBBpZUXUXZW5FkyvdZr8CE3YsraYx8+2K89wKTjR7e2PI1qRaq64HRjR
G+eJyyCvoJlX+VIDTw85I1TzjWX3VQADJSCLq9RtY2ysLWLAVItvJwcWAIdHHHp7En5UK1HeJK0E
3Ha244pzph52CbcfLlgp2NVD7ac7SyyskKb4KHSuU4MBJLvabMqaoJL3wYhjjthjGR07uP9qrGI+
/8LzQrFDbYCvusIz8tcbpIn1z7Jhc8SpzVSFgBsSCPwCRadiJZarH2c2DzlIHRNtQbHzXmtMJSEO
v+h78vdf0wuuI89GrhflEgCJscgmtKnWw5urJ7W8lGyzyoIoNtNS7wbCaUIL/pU2w3Xmh5KQeS2+
P99W3baO/4f96F/2xD5NykwElA9OlgPuNhTDW7pNqIlggTAnSQq3NRbVYutHMib6vJk6iGoLKVqz
HD9UVoMYz4eITYu/C4HPtRzGKJ0eZlGQR6tQgI1urks6UtMElGDUzH03PlntN0deQ49jbZOb6fo9
mozm42UuWqSNh8PV814jkFEBkkUgTOU0dsxHF6B+CiV7U1zufbS4rJaC/rYoLW3SLH1SbyRp1wQf
fQ3epw1Wr2PN654kSQFVzpYJObHAki0WGbC3Jw7jn/GOFc/TyMmEsZKEPO8dWoPQIUHZdaZYzzH1
0yMRTql/Ofuni5KttGtEiPAtK1k8niIU3QyHfUU5Px5fByuG9QwGiywyjRVQnWUBv5lwrRp2Mnq5
DMKS3JSjrTx4J7+iJnXyqmZ6fo+e7aLBLwbdKx9bM0xkgGyUzvMQkUV3lmbxUKQbjErLkl8VhIX3
NBuxneRXYh43Thc59ePaW9z52gNxENN/7owBDr04BkPg3E4kwWgzdM7na8bRmgQHX9EHDpPzL5C/
6YWiheo4cAbhFpdT/LnXDqdGg39QHaDAAkrZ1JV2NE0iQBclsKBFb3UEgwthnfC/kia4MYFkEtuu
k1BhfXOuHbpu7iWB5ZuBK2HJslphA4XvrrW6cXnktFrOcdMPm+yH2fa7J1P8NOhXhTbHKhzlf1fU
IUppCEGNKlBvbw1L5r4CbXmeCIYTaUpXV7hVOjWQ23kMp57nddsjpoMuEhDpXWa/a2jVvLjOcZy3
AktTo6zdUq3QCVwBQl/XbLXDB7KA2HTUseoWT4Ud55o9PvyI6nnajJHhxlLnvfdfMsTdVA7xg1Hl
i0D85UghgvvF6He9tgPg3dglTOSABW5B27hDPyU88cAm01tyZ1uVMMYJ9jGEYf/2tStJIChIp+Gr
0W6TL63/8XjIy0Jf69arRQoguB6bnu7idln4ZQt4d/aFdiMbKS0ButNr1iKKM2cQUY3FykeumBMS
+hPk253X4EFqCxGvGVZERCUvTkfIotIiHuK1Hi3+gtrsqTf4MG1ev/bWeiMO8yoSrJ8nxcDvDldS
LNvtGUe/ULResPVyA+oi4c8OnZDTPAnZJS4aEhMlltWI3GNfMT4M8uMNTqhK0C1F8yD7IDwfax8Z
0nrRypuxz/9Dyhee9kKVakOgsyU9ww2YFWa3+fB7PcNqG2N42ZFncfP/Cu4nDTBJZOU/vtu2slNU
Bzcg1FxqKOMXJOdS0wcM1uyOMRwPzNWeJdq7EsA/SlToiTJ1w53r47q7uhn2AiFh8GlGWQvuQTML
N84BQap08b/Ii9vZmIHdz1GJMAeTl5WzzP08ch1P2F5+i/nlUZu5gNgnGXxfxMLD/vlCWq4Mnt9+
mXjPGa09WQG0aKzhiVLnPZ/Becnc+dEIa+ddE8PCITHP1zPEW4ek4Cq47v0B7BPDTPBscTI4WNLG
/lhM2wkXkEpETvkBhEXAWvxcW23fEoo8Wi3XUwrESYhVN47ACqAGVenMjjdwoHFdimLbTAuEYP5b
KQIP1uN3LQ1RhPyb0o095T0TKUj92CUxl4biZ+n0gyZ7vl3tGMgNvuMWtVemyulvoFc7B9s/nfm4
DCtJ15iso2XsS90e85Ia/xjGcAUHLfSXP8liCaLvIS5Fgds9JGgv/OyR4sHGKL2QG3gL5ezw5hFu
oXjiSJjKPKBSzlWfUDLrKZ6gRB/f+3qFmH/oLfmBeCoBJXTrspXHWlT1ETrJoSeSZny8uQetVrco
OtkMrd1p8BVhPPklh3UUUDjSQPXDPk7eDPCNNurwNQoRM9wbwdpTY/fSPZ5HV98CN5AThQNgPtx+
nQ2K9mkRsumgA49EhPqYhTOg+8lFfnprfjDjhRniKWuhz8eoIRBTPMHRxn9R8WzgNPl7RJU6TdXS
fgUJgpJWLQ6AKCmeWXSnhtluTfteodSdj4nYTfugCAIgOm8T4YD77gxG/ScC7qrnODbuImFsAU2H
/hVItXKies/PCJxnVjYHRzlYa5QVDlVuywmY1FUcLFMlKEXGlo4KKWA61CUc26C9qHEeQwY3/Qax
XMlertTmI08Vp6wqiXtSmmPUntXQcjyIdh1Q9sDSyvcEXeexI/rfcZirI9V3358cxpHaCsSaPIsL
8e74NLLmiwYU3g6/r6iCnDFlntFmoyseAPdKaJAcUyDKzKAP49BMNx0MYOQakzQgDqzvjhN4cu6k
0IzlS1Tzmfr6ZUKd9uUnqdoHZ5Ab+yAQKTFbXMk2D2EMLDeglo5MPh/x/ca9vKlho4S26i41Lzkb
NBtOTOJhwP5p2ptmkxz3r4VAA+qavyAahLXIGgexMc527IhigxQy+YEjKpKAUttoyhQsIUt+ivFR
nlwMl41sfaS7KzMUpPZeCIdaqKjwVWRjZcKSb+sF55cpw/EZAqNE0+PVL8dHT7RtrgFo/XK+7zXu
FbpuElSMuMj3k9Fcj0pNw8pU1ZV/tHGZp9NYr+VCts1LSf+wVi3GoVBdeUZwZHhVChoxagifmUuk
t1vvtAw4wSioo6QKUe93KjaxGQQB6Z0jQYrz6MWRtWkmlaHNFaCP+To49oGsoyRvNSUFRpI7aRru
mWU1za3ix1bXZ28nt+rEEHzM6QfVlhrl0Ja3ZW30FXdOQHgOcrfuVZ/WTeeSVF6y/nzphhHX3uDm
4VjiwwtHgiq16xO5ZO3FuHeaTu0H/e8K8WjTb5lLxTTMZ+J3Q1zsXPgWDUO3AbFld4z4c22Ar4b/
JwLiADIIboFLxM2egNBibwp/1yU0/KL8YBI/OB9P5Tp92gNdS+pqCKtQCHdJhEUKnY9JQ6lNjZM2
6YfdqOaWLVLRfe5edQV/vwwc5IlRlSDt5DfYTH4NIPYeDkIgtyhQnVlwmEv/tg0z4R3Sl0kqZQ5U
vj5JQDQPMHttQh4Dmd04cj361Hb1aQdU3mKDlsdDlGGCYxLehimfYQT/lzpZddrfG5yMUoM1wZnt
HSZIMZMQuogqqSmMmtDuq5Oplkq9MQYg2b96XxSPt9pz/cglOIaPKv5Li6yMa0JdK7HVUTwrJSWS
m0fIoEDB3GEJ3lkDYeva0UB3vLxlAuAVkj14zZW5ImDPpPxTybKcp5LTrk0QfqlJ0EFKuVYS/x98
UneW/6eefXjhbs4MO8Ppa/YAXF1YvqFmeeBjq0yp0erAhKVtclaplbwxxbz1Eb1E/2+KKml/s3xn
sC6wYnyOphdcOSxmzLMN6i2F7F360IQZxF1N6VWghLQlN6/6cNvF5I79z/0JTIraEmBPPGAvX64q
UIaea/SwAGllshWa2SGLbg+Dwy138LIoEnrfvsZE+AOhQIbl2MfzPxvy5on3L38Pxs/bLmassOAn
pgSVIZCfVhXv+eKwDUWiIPtVYqenuTy34AA4oXHaGzfv3tctLcvzbINSU/gJ6SOmM1HviptlgLK9
6i6Z3btr/MqyK5ScIii1mz5kC2Vn/ZS+6WU/SVANqIvSBLtI5XEhOnVNuxVdJRxNAYoSlITYaGy6
1hjLCtJUgIgImQrvy565u8qgzoIimldySclQMo1v2NCbRd8toyasDoJev8k9mk19/BFNICwhvlpM
Q5MJJazXxhX3yXyVmhyWF/fct+l9hV+M8qAFrJzlE49+0+cUyE40L9M+5BqHUFZjddgzxAL1zlou
nx0g3ant41Zn7mnxuVIEcnQRbVvqLQwDu97nh/URUyEU8H6BEd9uGpjw6MmzaenP8QBz4t9oi6mQ
mm49CchKNHCNdgCMD/RpD+3eUUd9LW4J2tKhCX0pr8i74yyqtJ2tNQOXgMihzYx9I7/h3p7LmQrA
cNBv7KvZHXVu8QU+LBXDE5iKzNkxMN22GVtiqs4TnDzwvIhu4E32TYyLuf9hjCTmSeyikZiY0e0V
Nq6tR+gsS+0DlUlxn5Lo+Ag+xksG0eiczmEZtlpC4dcpMlYdmOElskR7VftX4L07HS3LnK3QvSQU
FZ1p32BBbtbZ4Thb8l1taQ27tM0hzaqYgvJv8P4WIZPEQ/AHRKZaP/XHOAjMoJKdOprR7sHM3BME
sJmGbMyd3D7bWz93DlVKPT3ALI4s70c4bCi3PGIBQzgZPivow7+Hg8Uy6FMQC52FMe/iJh9l3Ogx
3MYF1iuBhhfotq2Vgzm3C9en3YE/UzHYMzi+Z49DOP78QwJGhLKCe4ABtk7KaAnGPoMfuEK/5N+q
L2zEEkXQ1khLim5EOD6wFoXHZMzaTsRDXW1WSNzrvvRnetunrtV/deUOFKqY1JIzo2ObtLX9+LFI
ch3cXnWUvR+7sMuYfOK/lfGT4BZO/i6XRzMefa8AgXbfAqB/KHdyrPt5romApMKk5b3Yo7SOmZTo
8Mjaom+tojiw+Minn1iW01wUhDCeD//tRiGhikXA9p92iIkGg9gWa0teY+9nygENNGfRVZU04kF2
GUonNDvUd3GHBWwpKjSaHBL3Atzw8EUcRcgGGWQToonJoAevuKE8sRwgJTp9akdijgx36LUM+n9g
wKBYyO+Rz6tkUCjoSqQrSCMsQk/GXFd/HRWHxWhJw0oFcdRF3DVzzX4XIletqFeYYyK5et+8JXyA
yUxmsOp9MWd6RjUcfzz/e5PKWEIjzh9qChlAkDzC18GvHx1SRKKWqCJD9FGQ5f+gr+mxLFzYpi1S
hMdh4EWEhUM1WL4OOWGyuH7UdYD0x39Xcgy3DeXNQqb2tQHKGyEKsEn0MLt7x1O9KxZaFDIkL7aP
3aMtzyDzQv15VAJi3zllH+VTav4Pgqq8JlOF7Ona7Bw0UhPf1KYXDCbf0Nj4bANWtp1UoxC2lPkF
b0dlEueW82G1F+yZTnwigbonSA0HpUpJ0m7Uq96u56pF99dvpHGSc9ezgEhK3kRHQ1Az3/ZXJE84
rNSa2wuj7Hjwqan7ogVrd7SSwCoKPXVGx9wZwujs2RRAnQJv/zcwCW9bLeo625K9raM0eA0n4vu/
F/E41lpved8SQBOeS3qeGyxm3lGnxRJj+J6reSJ5/YkG4IilJ1UjMqJRRB0zwABeNGaeHG1MKB1/
w2wxD+btC1V22l/UyypgDXBnRyaDnmu0Twocg/0OvMADukM6/nFCCpcbfBWIOn44+6km9ZU2+6bD
H45aAIgNVzDek0l2SU3lhqJfNEkl+0VaOR+AVpqCud3lMzygXchavJ06X4GjMsCw/RA8k0F78lKv
c/lFaJUGyJo2EmRTU0+CBGl0MwPUqvRgR95CDl14i8CpbUjIGxV9XrhRvJ+Sd7pDmhNKtdMeUOSe
mayHXIfrBTI4JmrVPjBY6fVvIugnGIpA8WXSO4FZSdPu/X+1poUOL2pKOoEDUNs/Urc36Y4aahNy
vUX3lhTNHDdRdyQCJZK4bwAHCz+wIEAG7kO4BIKw+ybVivaFG4EDv3Hcl8z97f0OIDbBuPP8KH6E
xgkGoDzLvQ05ZKqKt6lBWAw3yNcN8qO0oGWkEUKjDVAzeOYD+64MRsHJWe01/fmMCwi0Efy3EX8S
lLB8A2zK1m05WQrl6T5WP2WuRLx+oSOHppfcmriZPv6WXft3cJ4vVeDFVbRxDWnRY8C2j84UpmJN
7GbGWf9DXhwPoB01SjMCD6oyV0NnC1JjWaQATJ23VQlHLZyeM+REU+gfcjySXe23DznrSPcb7XIA
4E7ozaokACol2Dj1z9L/Dfc6hrd0N1PodUmk1Gkz9pCf1VaSJwoT1Z2BmBMHkS2ERQZWxFNMNsQ6
dpR2rF9vKLb2AddY+2B/vB5bYHv7wfUVnE8A1fZ2/qC+OXsLG0AYRPuwhmzH9SEqqR/DcCeM28aY
xccGgO4joQcvn8JtaPTSQt911uiF+iGPDuf7pFZRUvT1qDe4dM/KmVK+KrfREzUp5HhygKUJb75e
TZFQkGBQJBnIhDbR9z6lZatcuFCNRTc/MNW5AKTYggsf1kN0Wh3nneZ+eTEoADBNSlRsqi5qwvQT
Xm74RBvI0BaEtjR6PoqAnTGTI/MrPdtYpBF2a6Czq0fgweiUGM3sIiHq/pHC9NmYMmiv7DHJgBOL
VVXHyd+KS8CQCedJpJ0pzri4XcersCJXTBWN4c1+CcW7YKNgWo2H8flt71275qIXiXx+9oZZeZv+
IF2411kZuezLkerjQm5L28eOOjJceguVXt8Wjojv9H8N+AzcySbmj5NpD65rwZBJ8owFfg6lkgl4
lYaNUJmg+QRZ61KjJuprwkwERYtaooZnkvb86K/ocPX44kxLKSAFXQnSj/pwUTZ4UaGQ1GsFLV+o
fFd9qCMbMkF4d3nEzenIJhEHY8db6cqTnuNA7y/qXUJjHiwFUePb2wslsr7BW4ng//QuFURHZhab
pzJP3fNKSQxt8L8ONCUlRt/UBbgAvz60Kj9Gq3UJsarRhfU4ZYav4ngcAljJwKdHaL+NDvhOrInz
pckLgHFHI9Sf8ulGK/1nFVtvIbIAMMR/9UtwFy/Tjhd6SJXeKbAzclVIEQCXECSLv/h1pL6QQ6aB
tlxoVquolmWx44Q8SiWCApFvAnXhy4l3gTFwaYVm67mAvCWlTe6RQZIZnha/e1DG7xzs9nOO2uBG
3nKJkPgCS7xlxo6VjDeWnnuv9Hao6CV42z/H6H8+Je2h2zohOODLUa9aGmYN73RG0W2Dn+m0a+jq
Jmr3w8tOiBZXTqklQ62hr8i/e9zoYTKBNH/foNS4brBSS3EvYXPrn1y85BJk8q4rksL9rUXt67G+
O2wm5bkrp0vPr1VzRfa7DxiGTwadPiaiW21b9IPCkeuzaPl1LjVEausnBJqG4cs98MIOmAKuVAvH
CAyFb7v/3PLIVj36tK8xHC0KGQj3umvfKxFHrZZTcCcwfszgQXbmxhMDnm+4Bgv4x9ktcVPWiWdK
lt/wRuLdqyEjFaNda1x5NhZyi6CzGdhCVC09rXzlsIuvqyPhQBFaiPQiMbNdReE3aw+D1FQxsHFF
Zs2AaLh+77Z/cCookh+3VNEvrItTz+lufjWL3ZrISPj4iJMzrs5y7ga6hJEh8U4VfoM2a2Gw6JUt
KzbjcVcHHEmtrC6JfCNU/HCGTLtJ/z/FNVi+tgNgRfs5eHxt70tlSkbJQzU79Btequ7rKNyT5575
CdeXLKC65/NJKOnF3UFClmptK7bNOeCJTAME7WOszSzo0o4LDrucXS43ijVwtMslsfQn8/Rw1Ote
FFE5mzY2iHU4jDUFE5+DH1hy3cDNVAKLyDnGx4EEFGbdUYboB9jIfHabSDkvwJI11KAvHUMLgsuq
58EHs5UH3RUCDDiaTa3EksqWBaOHXyGcSBxxlHkF2sbHnljnVVedMwlMsD9Zl59VYIcS9J9ewkqr
EZ43BYQkjQEMlsFH0rTkoeClo/oayA/tidaMMM2s8uleQLxJAn6D3KwGUxJs5ZmYSifn7jJrL0Yk
8mobelRmdEMT/05f2HYOzcLAhPyTN3sryElpSIwVyBejuhYbQ32r8VaRDjHibIcCxBiaJE70EeJ+
U7s2uviqXyX8qkSRkgF45MjPVeVr4m19Cb2PMVr48zVibJ9j/QbU5zARKimf//iGXJ3By4+DlR4i
Q/P4lOg+oM+aGkoS121mp9bXpnZNiImh4m3SSwmGg99d2B6kSncqnrOs6itUyYyihyG1DBXqGEjW
Evr8aWbLtd7zZSL83YCBayz2/MvaSz2KoE4xynJbNphNliN5PIs3GXQSCaTdebSDuapeTmeh4pJW
WEYLkGHvMPC+HgH4Gz+LSctDIaCl+A7KLMkT6m/l+W0zmWB/8wy8GaLIobJ0+lWBpcBcpnlU8GCV
B9zJQeTCu1C8eWzPvFHklbUo1FLpnn6D0nuLUe98SN/zALPrku38gv7NrWCM0auDdTh2g0qU+JGX
ItR4try0ShHhcD2VGiY/lihXGCv2DrW6TE5QdbCle5obriy3qnTA6GOkh6+zPpwsPOGcYlAblQsY
/jMGj0kmGe4WoKsv7GuXp3SgumRnjUm9NmQy+5Ggk9x5FprgxJggUwwUZu9FH+C+gYyIPCRCEx62
ZHfy5fFukQj7gjRGOfktJ0drJ3OIoNC5mMT/B6E+PYdxZV8ePTq8uxW7jEtnq/QjQfy559VLPTia
5tcYpfRMRtp9xMHvn/CcPfbJH01o2IasFdGNnk2qS2nLeYyBiu3p1X10giNKGAl+fHUVXOEf3J01
tGBtUUEllc7r/1AUtGt57tGuFmYdHHKjetkL+ae1nXZkUc9U9rT2vS6Wx2mxJDPZZ8x+RjeUHe61
JFV95FiQNclxV/sy3JL84dKCBTs84oBJ412qms1+j/USxJCPNUFT9k2kyS8mCqNnJ54+B2b8Pf2g
7bvYYUjbrrX9NrxUwDecrlEKIHSe8uaSmKHOcpdPUzNa99A7MWpg0K+7DjszOajlHWCZujZehr5q
K8c+BgMcAFUpCApan8XnpD83ZoFUAiENqvuMyMmpZhTo0kXPYO4KlXN3b2kQHOBSJIEK8RWe9+md
U53Xwzxi0Ydoupv7BZrUM1Xe0x6vDPpErED4jaGET4putA+FK0rS0nf2/Z0WQdT0DuyxhmSMfSix
UJ87Cgl6uY0K/Lcph6NdtwYl57vOnlWIjxeWz/0luJn5bVkR5t0Gjzzn4wERQWEZzkZPQS2UKp2k
KgxrXDB0D4EjxuKeE+Tyuck/8fW/ktuaLhgljiAfL4tiGfmODjBZliRj+SXI98AgbRuPjQtQHUjE
lnWr87kG/SME2qjaoJPb8KrHm/re939JvidyyM0ue6WsMdxPQh9XFSZtyC99dQdFO+D8lbITygbn
sPElr/IJfh77j9GLq1bYcbmcHN3OkdIN6D7Q/sEY86ei6qlEhaGeLntW8apagMDoblblxb4ht82z
iMe3u8XwYnlnBBC0Y0uGt/g/ukt4Tosxb0CnVw3wW4ybxBYFBcu3IoAQDGR3p+ofBCuTlm7sZewQ
ejBH1tFG7AEls56MtFzaKuSSSs1c6DXv49CHiWkTrzltUxumoflkTsgQMilsNwBkY4LI9Cn4ykWK
L+OIICY5BSZSmqKuadfhdclklz9ezbzo9z4EaqnAbx/bPQ9jLqffRMxb7pD/4bmdjdn3FVksE+xk
e5VjMso+WxCjLwYf2z0AGD0ieACspxfVTckfJA2rdHod0c9rtT4GUkVzMzDKVEW0Ogic3BFUbTiZ
ANoD06qh0B9Yl86YWubX18O3H53EvgKIGTLLo+OFC4vHnOJYxZU7QVI5DJ1uXYo400xSy7SBYAmI
uCjshapJzes0InxEX1c5Q6ugKL47G6eyBbgvTdpYFUfslPsJLFAC9zuQtuJFvnbvCDWslnc8EqZf
AfYD7uQlwKQGDClKYCaFOShmLC0A2b3eU34tjOYh5uk6zvwIQlKMKFRWXxbiqcEbIrBY3bdCSQ7t
6LEuba55Dmc1qSBeJy9vPWKRbuBZqg9yHP4ulnvfaBRGmZHyhuwC2IblQS7YAaMqcXVe+1I1zdVH
KTDE6vyl8pKmo+g5WnLrtfEhWAhQ06qQNE+yLq9g6xfk9UjU7S3TN76I02y2nbE5LVq2TUodXE6B
6JfPw3Oubmnqis175JTgEM/9C64GmeL+5nmf9Ce75E760WKFuFwCKsgAfdhi4BhSoFGjjqCpg9VC
sGW5Qsk9/Z+RqQ80An7yAioNbw78PhPdfizOMdoKmW3GqMeFpngSRX84aLMBzWv76sOfxL4enFLg
wYe2vlyDDQ3c/I2dlnHGU39HWkmwJ4lTgJKKzbxyuh24aCypFT4+jW3A0Lu8Y5YJxtHt4SKttKKh
LhbphAs7TvJMOIQtsRxyFT/+p8sfgJat2KaMc4+CskkL8zlsBnK+E0JPjxTkodwzpj1H5fbVRztZ
WHFdFnl7mrH2n9nswGYJBw7C5flyV+M0xrH5UfvifrRX4i3gWOVcQI76ylg/PfBPPsHixsZAArpC
xOpRKVGgSj43E55kv6mIOBK3QaC/S/3C04MhaVHH7Hon8Dk+ccuXvh/6HTN0L2HLUQPV+aWTE4rg
PyDw7r5n283i3Fv+vXpcBq6hHaV3TplzKZkA4tKoo4eNRDYGn4k33ja9U9GT08wn3q85+K4qKGY/
6IgFMdLlYrrHzX/+8LnGokf4yHcK5vXgVQOJ1PI/8VKNpWLnQmT7YqMAI0NP8dgFCrQ+3gdepPh9
8vnvcYO6BFWeZtBK4eDbro2nBTDTX2oSd/XxEljh+i4aYAvfejf2NIuaQf1IIKds96zUShLoBDDi
3UkLttT7GZzguw6W9Eu+hA3ylQWKqgSRejqEq5x1Kh4PWkwCTk91GPlmrkik1dHTxuSzQNU+SJFy
nuGz0FFeNgsUbqA478AV+dyT7Cox70/WPBOIqkuJGAICkDSjfmlQZuWOElBtTwf3fjCXQv4/x4sf
Se5+Nc90dAe+cECJS1PsgbAzRjXFYpR7S6HSGCGtiOPjK5FjcSDLDzPkb8JYSheB13Tpnj7fR1l0
d5Xxt6q8NQaba7+amoqcMg+Qzvhg2EeQuJ4L6ZmppzJDZFeq9GVcAZEjVBvGCozSfuSOVdH46VfG
h2lARMKlTxVBcqGHfcr8yKYCVf9BMcVVCPveXR3I8DLZYitso1Zea1c9sW/JhcYsksL51hJo1Way
JsY2f3rMq3wqW/sAO61Ud75llS5cM1sCyDMLD0PsIxu6iCYnyhGey3t7+jCs1gm+r211aT9LhD+V
NAfgGl/H5HNJag6UzIPWW/Qskla1HHu6++XYo5Og3YvkaT/ysORSpVJhSnXGxD8/UBnyST5Gr1V6
Ka3BaW5Z6falYG+5TKQDpodaX/kvNvmuXnaMFt7nU3oYr3xybUStX/wm9XNT1KXWa7rNKKNudgbE
j6PzpAOqIzQ7MczQL1K4kndcdyolSoXUOKLi7wy/fSrmYGjGyvCz1K3/zyEmd61a9yLPrHppPK/y
UEeeWapSMjchwjNgzzjrQ677BCzfXW+VOkZNTKPie2fiCjvksoMUhhVr8YR0ZYFKeb0UNMFKeZh5
g8PUf2qaAMjpek05DtS2QzcRSjKslOJZOTK1B0J+ezpE/3Aty7O/B48vyBqQiLfcfK1WI44FPOwT
FPjKVPY/DRhjtZvpvJRPbDuibe/V1EQNWwGesYX5o2Ql18An7fW4VbMRql+7wvN7dlAOsFHk/bH9
+797e9lH+ICYFn4Nv87T8YI0PR158gxWPdb8j0FhDVYbSKkfhStTlSc6sR/Pf302CjNAcEnNOuNQ
vw2G0d5pv4VpTvD8VwhreiHM1kaGKknGBjvu9z1Vmg0KnSLSUCvgOznmUKXmCxHVZNepZTfdYhu9
rPMyxFPMo4Mthw/hs4KeUrh8b9IlwiTtOMAzTLYShgQQwu/AOch5Tv+E/mVil38ps0vuFZ0Drq+t
dNRyDjuENPRkzTGy6GlVIgBRXKq2lhyyyUQs3SmHM6BLRY6NVMUT5fgwi4jxLJmzfgvd8W1VHubo
GdPaP/wSZi4cb0cHYAEEfxIqxKUPI7tq9XIqxwEnFRaIel1BnrK49ykj2jFINVB2hZN4XdRAyLYg
POUDnvJlVV/ViFpFzHnZ/rFvkLeOQ8btGbCcrpmAvEkfE59/v6/uiweYKVwOrSVnk/JAFFFAHyR7
2FGpVqLD4cxyuOK8IK4C537os7ebUHzihuonN5WU2nCmFLhWiQ7HFW2pFruxIgMLikqsf3F10reR
T4uQBBxY79PQqY9PvRxtnAiVGv5AXHrTcOUxzXMGnPOynQ4598cfMNr+Gp5qWetzNfVq8bzUm5aZ
EJguijU/sXYEclzBcnMK6x4wXYnGbQp1UdSQ7GqgIqpU4mGKJ5/RKy2n2xqLr5LOROqhZ3jfuiBh
8KEh/YA/WIhDEeBdt900uwB77ZkchPE2CEYlF62RpDufxFHt1Qnzp7/TGSC8fpum3QuyOyppZcJv
Nye+QK+xPfaTdSClsWB70c/URueTWwQKZUlzemJx4LMV/73cOIEYIXbYEbpdUXHwOSowshz6dfSE
hfElNA81MObjNu/KSXSPX2TCSUNH1IlUuP1wqAOI3tvefzV4+b8VK/ZT6zMDwfTNJxsN9iU1SBCY
cF6bMvl+SjXPCTdFc9yIncdh21E0+YeoCPqoUiN+oM6BLzZv97deQmo5v6M02TG9St560QXc0que
a4uxlVGmuEufUIcENgdBDqpdi5lEKfCdKz3FuLTrfcGwWEJmTN/henq/7YID4jD8jawuonaia606
JEBfifwNkPeZwwGZoUMaVDVHje/9/aphQnC+LKdm16oVzdya67ZPYwvCM+kLOlTHhfWUCNpj9bwX
E/zCPVGgwBV0Dffo27LBUVEdHSbZqIKoeACd0gl0dloS1OK2PWg9co1x7Gl85/0CMIVKBEjGqInC
9uOruBxECAkyxaxQhjYMqpTB2WfPzSOca2GvjUyAVI7DSa3PSDBmgPNOolLNEWncEFVW96e+yD56
YwSunp+45jpIciUROyqJYYxK7z2Gl2VmTKVjN8CF1eKQi9N+C2flJ8KwS4NlFbokQAxwl/itC6zY
dJNmGmT3+Ya9RUfAfoqHfk4OFP5u0gZ5wGtTATWrPh6Mubnnha9oksENaJlh+j/5wrN+/8fgNFlp
EZEILdRK3fPvwrsW6dMgAqKgyNH3BsWxK9sCvV3kPIM3OYvwEqDW63K4fkdvYE6VcRniM1gNvGKh
6YAY2/osOIfkpZJ2MMeic2wV6bsbBZEP8Qgbe+NMEUifnoKEU4mpugFhf4UGX60IcZQ0R1zbwPSl
qub7dnDlmjTK0QCdGpNOKSzZrpQ+2lTsWr/lRc5shlimlAh3dfpxhyFFnhJ6SiYrvAsxzrC4tcfB
RtMG7ug7XeqIY53nD4pHVkq77ab104JDbCLDbMGtdT334/U9ksXkSH8BuPM/rkBuf2vRzV/6mM+Q
EUo6Pm2dN7pH+5I08F5+c3duPM2W2Qok3t+d1Og0Qe+Xja2fu61NzrYmDy2WmlQvdOfea93RWI4h
6pMWcBvMOvTBsKPPdXS9EK5adANVM2gew5irZvphhvwqZpXDlStR8EglWh8tak5EtRwSzxsdMdl5
m4kcQI2HaAziWOxYXJKAjZnDzX4CWW9UtEVOOpc6kcHMmMl6OYXPrr+c0R8DKXirOUn+plE6xTKy
MEgKiNhgCvL2IWnOFqNlt/Y7hNql9YqjYQeT+RHFzK6usGIu9Iuib9ReeQyD4FVc2TMroysIFhPR
BzRZN0Nt/w+ulTdJIAc09CGDu7+RqmkhuQ3WMwSuB8yelXs7GElTznTHpnJGSdfHVhDUu+Yv/wKX
RwRDqQhvGMVmjIqMZLFKKdglyxcvEG+rexuXb4EqHeISOfXpsKk5QFW7vHK268QLiW7Lf3YWbA/g
JhtKHITItOrTUqElumbEsGsNGzKEdxG2iNbac0Ecey8/mHs7bZl3fsl0+UJl3lXmvF3Z3qvagtYp
1e+XQAe3+VD+gc6fKbfjAK+eobhvaMIkxXJp3oGjZRgVOlQeTfMIRLbowfdMgXgijakdm4BrycZ1
scJDnkDwks4E5rmFkvgRkG1b+qUEexAlgzqEzIi5hX4NwRay1sYo2OWKOfO4jflJk92M416TIBGx
cL5c2lYcGKSFTI/AdSJPVB+AtVYRitbNXkJpK+ePKzDWgpNvPnnBzX8UU4tqi7P2RELvoskluTup
FpRW+SizEkkyMWXinI6ATXoGcCg8SfeOHU3kp9KzOEGu8pc0BEAJQ4Uyl/eMHTnG5nYy4N4T+l9J
fIoMUMIrKiwlIriva6n3m4diluQv0tQnNpKGz+n2jNzGu58j3+B/akgX6PLAMhrESGW3UzOr771G
ncsWDNjyTHTf5YKJWiMitd0MDwHVrF0q/wmbYNPtFX4hI3o2rgjG4XPvmsKSWllx/LX1Qkemx3oC
YJ9Hf/FCng29RI53roWQdKJ/gjifBBL14FJGuonG1MwQsOzK9mBSTTBH4hYDOV+/vBy9IVK4UHvd
Fj8t0q3fyaqsX6rD2KwALbjVg/SGdiz630XBEusibAqbkDL2NVS7onWv1crgYqI+b96hjzdrDveD
FG8Hm8GoaV0fTr7AUqI/4u0tA/2A5p8apqCy4u+3VbHB3rkLc8VlVhiFb/ofhYBeYMvMokq5MBwa
UcLjG1hfyJpNCVlbRLpqxOmGJXk/1Ww3ULDSZatc+kbM4GxAGUWdIX+mdVH1sDW+OafmntGP7J6s
63Vsqp72lwc03EZ2OVilhWfZ2L4YSawh1PLjVYAVIRDlpc/04+9QwOVM2bkKG/TjdDtVBh/guvMx
MDSZgIOcoUot3IfS2R4U5V56ioX9IB1jY0fwppohcIJBAbyDHnmmiTVykOIlWe+amuXzDr+pHi8I
8iDr+WXeFH70kp9nyNHxJqPnGDM+Ur/rFUL8Z6QX/3EtBfBWSv0KXPJKKYmQqNMNco0Ev86ZhK5U
L6fE9NR6NUbZ13ZUc7QzZFnmiDU1LpBML7x/zafx43kOAWpB/as53DbrCJFLSEeDyQ7raDBY6Gni
zNR9tLun30FpPtOYYCrn3w8cNVwyzJWl+VTUeE8qQ1UFUozh4YrlYj0aWzXaXOWqc2T6rI2Isf05
ahOG9RA7We9NqnZN1tjkPHEgDSAML4lTHpUxnEGxqpns+C0xuaI7kKsehrvvEa/pjrxkBpOctPSf
UzZ1ADu5woh+lrcXKCgHfGPZDzBAIvGVyCdIqvebxnoRzn3Bbmm/qxt5m12rIuxilKXUnGR1bEwk
xXblI4CW4XyOV9hDo7AZoZpKccqhJpDHuG26NUb+DXE9wQ8tZOGj9kBFpE4ITMjI0aJYyN5TcoHc
iCnYpSxkdwz55O/hzlSHIrsb0JvZXvbunNfQeDvStjzqJODnaP637nVdIhvIbjx3W+0TT3oLL0mI
95Z1Enx4WKYNzYh8Cs1+odPEd4HS9hmoem8Chns/9Ubo7Ry+BHSljdXYPHLwfJyBPcNgTKER/uYr
d3i9x2AgFHiFiwrHVJ4V8sc/j5Y8IHeq4kunYqt1wQ1yxWL7vx+NONAewYYJAOrzz8xTghtCkGSg
x2znif5MVlb1x+HGZi/VZ2ImQDsXUfRSRYTtXdpl0Nb4dWFUef4ET5oDtBwv5DfBK5/T9X1yzulY
TdUQ3iGR93yhfegUMQjo1/8Xg5E43bFHtPKdamF36nQJ9Ssf+zlhkAqkV8yttkmcbiqO1iaLSRq9
ZBSdXIOpFWkogdkgR0kJpK/wk5wGb1P6ElitZnMaVlBupTppKlP2s4Lu9LHmhbqXrqEaZDZABALz
ekBZMaoInNnc1R5IzY7asooZKam7rBg+rvFx/g4tgYGiQix+VAh8f44Vyls2e62ctsY5QACyafho
/SHCMgmF3Or9nF/JnQhrJKXYXRwf6nSWtfswXLT0na7KuxTBX49pL/EdXyu0yo3CDlVoIemBJruI
6eftCfR0/3Huitz8/opeebtlf0PZ9NaezFreow2e7gR3F7wq+oZiR2R0i2jJgy+DzxDRgm9yRHlN
sz6oUOps2q/yvWjafwDyw4KHu9eKeOd+lI7YaoavBT0rK6Pf/pI3IOZo2iM0bjPd08u9x6dZ7vz5
/Igh9JgbrUqQ3LEyU95kjCGbl4/ZfRovCzUFuVqcO8mSb7ye0CLR8PvZSkFmDKENBQOXGnIB9G1q
3RLihpYwqeun0oISz98zY4XjNY66zwgRVnkdvqg6nvSDETkS4RCjamGonIbjNS47CnERlsldBnq4
Y3mOfO+ww3tWymh0QsU1vhcGCqLFHs1uz93lXK22pcTxYXwH57ORAmJ4xZJipaAXAzqPda42r+CU
DmFsMLm19ddWE3HsBwXU9s0VdEib9Z2kQ+4se1GLhx8Ru5n89IYp8jy+HtKVIypjQ0gFDmcxi0Ux
IHhD+JF3n4L2zWr1jBZ1v7oRcGyvkknCIkRh0CBVOMoSGqG+UzFKA9PRG09KXHi6C7BsU1NVqFyS
jHt4mlC84Iul4GvQ1y60746AFzAmC4W4fIP0ZxMRfLhfCLegIK8M2oim2B0MOlJ13yEnWtyORZyf
aWDaP43Ew4xGAZPY5ERCnvna8OTcdgtwoySt64uDuWnXv4K2uJ7iYk0MdPTH/fto/yedbIHsQugf
km1OVForGj8DWGn4RGA9WfQFscWkbdwwoc5ChY157fGNdkHQDeKNXajwnXa5yjWVelZ21jLM/al1
S1raRpHehWFV9MGPwSeZfKUe/pqCeDgsIe4BJBT7tespWyMlGJCGaKa/UFBRRdXMjLoKYhobzrvc
0aV0dMngW9zF52XM8cBFOGqZPr7jXoQ1q+81XlwFJ2VkL5ebuZJByYxbCyLbL+w54u0cjWPPjqlU
HpeMCtkiG+TTP9hGEbLSMx61RNa1S6ZMabCdSFXyZTxXZXOIzdgkpIJ/+S6g4zn/6g4ULZ3oDik4
YgU6TpBfzK5wM3HjSqnqW6UwGssqsUCddDKXK3A7uWXzOWlnUeG/040cWvXGGAu5vkPaBQSV0XaP
Vp2835lMTd7ytcn9ittK3FfKE3URsVKZGLsygbEhFplgq8IckqMnBTzD+OaGrNq8bVsgM2Y2rC6h
r7CCvhYytylM+wwwXgN9HL75YS+xsT+4gRCNruB1vXRfxZuJCuLmQY9EODPZubHnMhwwoc0hU1w/
vIm85RDMlEF3sTvnL3OndmfCNewpMRIqjqJs0WTM0D2+kiIeh1g6ynld2yZawV/fNSr5TnUe62In
4X1Y5TI6c9uL6awchEfcX9YwO6ogxSw9BVCnD7nEfJiWn91CRTmvd6mfwcnVN98HdcNXxJE7fSBi
rz84Kbi1bvV9iArFuzFMFzUcrrxBMeKPyn3Z+LRMiGE2qLlno+BBFahL05eWrtxTB6Vxl7t+41MM
33U7Ql+DPJ4Nzlxo9+o0xrGb32mUwSTat77r2agApE+Vz5G3DIyEWURmVmpnE2G6clTwZbRcsW7J
AN9UGxSUleH5I8SCJ5pdC0xFJ/DsUAUnCzvkVjYgYVfWuYJ60RU7kH8MVoKE36RGPP75nlHuWqHK
DX8PZVRCMhVVzvrqCFBQq4/ZJUsnYpUW04rHh1rWcc0bH8KZpio0p4NI5PxoA3I2nCsV68MoqxMc
GcM21zgZ4VHzTk7iP3gxWutqOjsIYxyKXNV4ZVZRl0TRFXVjuRVDPv986D2Gjrzk/iggKGL0K2LY
vHgYilabzYN8aexfSXU3a2aorMJhQBS/siQAfrWb4KvxvOvuvBQ/YOsrsX3GN5zfHHRlUfhxlBEW
hDytASxtkT3fIQvUXomSoe7iKALPWfJDrAR71mh2VJARZ4QGJIC8nOfFE4gK9JjfSWs6hfqIKbKs
1xAOcGoVbrAN3JWCjKQLdikiGL2oRFBZRwnn97jJGzVj2tP3CLv/fFPl+UdaokbF6Izt9rQXfvIY
o0mBDFM3OKVDTfmUqSNenxu/fNLrDJ9JNLWmdUTm70qiT5dXBQfjrwKUI1OHmDiOCHmI1pMFMM4W
po1sDsN15WwrGRTviW1mjwA3auPrlw4FthgMlmrhPApvsLd4N76tWicwY99craPPYNWqJ1OHk8Xr
xKoxpJPHNcTlGi9i3TVJ+j4J0ZUGv9et2Nh+XsJ/2GUhCfAoLTyWxFxnwaMYgs6XRegkwd8an4Sf
3KDO8LUbKc6s4940QaZTClHwKw8mrhW1dwL5MvJYgghKUP+xBDPtWfeFY+7ZKQhciv97kyK2lmdy
4qJBlJUQ7GLTGtBgy+yi5+cEh8pRwmyk/itIsZIuxaRoo7fSHjTlZuYHh3L89oEvIGX3SKkzuRnZ
6r8j0+yi9G7xuQrKZGsXdZnsBjIOPkeJUzg0tkW1wux+6LiPl8FipltktEVaveUiocATpUEJtHag
yaAZb6mdHESmuR1SnxF/iNGZeNU0bMLrFvUbxEN3qkWk/2oYqDIJe6zrHDrUxMx8oKTTqlYatZ+b
x2BNBMgZB4+59YJYuuxMhi9/w70/PqyCrdNVNuh1QW7Hv6LpKd9luFLzY1edaaGI5IcpJ8HFeCHo
7NuZvvn98uuvACJmiOSoO9Lu7nTD1rzA8CHrjUWUhQQn7MLn6ZtBmua/0QSzXGD5o1UOKcxrRIUU
fPddIMautstWgKdwsOF1utyIIH6e3DfWFADzcod12F7eE4A6VJI5mcvLX6fOWM28tTFGV+UNVsCE
2hSRftDFdgjIFPKDECCqwnmDmF6h56uh4+6i+8Vv406JISYiPgdRT2/IvjfQEg7wuzPDgfpyOnKg
KcNdM8TbKN1OSR5MSnCDbBoRC14V/DMNV5046pztTAMY26ngdY/eRQtpS0p61uU5gp66sH0pGmVm
+6354DqYTAvVN9cmiljshQON+cLgm/K4bRh+kVZlvMCINKBTAD2nvnEzkrs+MQw/osVu7tR01ids
TCtkgkq9SLz62COzl8WFWHTKArKJlPRIs9iYyfUgUrqSRkxR8YlPJwbsLvgQEPg/vjc07/ytzj+c
byiGyUo8NrtgLVYyBqu4NRrP6o0QaiiWTd5hoc6RDZt2hUz3v+GCKJ77KEGpwUOiFQE48s6D8VMb
9LMmNG1w9zCtxTJhdBCSI8IOWOkggT33QQhxD+6l/V6bBn2oeL391wvAEBF5wd34NPx+DYt/wISz
o/hsHgzPjcobI7mi54jaXJ7Kl4WdnocTLeLKsLuEVJQAR1y6jD5cxDCPmY+pCkmTagm00hkxSpRo
0yHOtphPd5spwd/mo8RSKcFYlYXqJVoP0DKXD1eNE42LKnJDDLPcb8i35OJcfLEEFtbazl5bLq//
BH3/dIYCWFVZ1SCgPKkqyd84urTZLKyiKO4kupzhNW43jgclutRCyiuAiER4MwwSXIX2rxgrexYL
MEsEtKWcEzCg2dIyWLptpk3HcU4ZiEy4+PZeFiNpY1ruUZ+oY2RYBQKlTLLDW5vs2pT97uBvHedq
88au5k58uyQuK8cRtLyEISbwx8bSyPtqByaA8pFkiKu61j2l9xYAPb6/fRo7wPymRehYE/YDrLeD
u1J3gG7cLQHARVdHQDG44BE63m675p2PLcM62U/0lKSePPg/WWg5yLz3XMefqA6Y+1fV9Nif9ag5
6oCZieZvUmDYT8nb/G7q3cU8p2OhDUzjfz6l7Q1eNOQ8zy3i6f3DIc8Ity6qLuSjfBz5rMoHzhg2
6AoM1l6nkdDwQ6ZK7fxcIo4ZNSNyI930JwQq14Cl6OsYFGK5eb8Y1PJnjl5P2nQ6gwP+YPE+xogX
SusnQsw2uvOp4bV/B9u8i1B8GvW7mCPvLfLE+7ii0VdR7OXHPS/SHoU5K6BNjW1cbCsJ/RNL4pdC
ZvN4eNu0aH9kdnbRpwjCoDt2No0HTbsjSiEsLJnlTiDTXPKbqM/SIf5X15JYSfdiw58KVEB5ZIks
9ZV3EPLmBM2LJ0M5FtJqM2zpm+524o/EfxT3bcf5MJE4e8QVm6iTKYACNwnep6iasyONuloOPZKH
kGZHFwgB5gvNnNSQvYxhjcsy6uQb9LpN6srI7NY+3fRj+nKDwO1LlgDCQD4crM6ASwlrgr0hrA5f
GDY84mEkKQuWIbFOznr/Ynqb6Y9zdsO3YjPtZxyuNGFMhmMvoxa7zDAs5rG7PPJOw9allyxjplxN
avOgS5lsizGq7sYQcZhntRMlOI2MtL4pa9an4sE4mdtpFOUNVd/zui1S1zbUYKkBKowGcTR/lLxT
X8BOVhW/5UrwBRlTdPPUQ4C+fxaFEviiUQ3Fry3LXE0a93k+kjo0OuwwzyzOeCa6UjfAf7LXqNVt
XWJNcPKP7Pv7kcG4iNt1XStdoTeGtctoM3DQX1/bwHA0RegL6r0hEdjcIznKxrVWESS/Xrw4Wwlf
u8yZqsLywVq/Rcpm0WEUzFO7v9w2IZhhRUMewvD8E49AR1LO0TxVE6yiNCui4CpCek7oGz0YK2MD
2U0ZZJXyM5oZxgAj7yHIyThzuVuyX1160mQXA4JkALcaYa0eDKDC0LM9qSUBeZZCDEAGJmCX3NFy
Pc6LHzFEHxrMpo1ROCGHzsCBt31dOTFUuOCwapVQU3peabnQYrpQb+u7bUh06Hgl6pekubNQB4rH
DLyGxVkm9GTuNhH38yXVS7t15Pr8PMVZ0chtDP81JJ5fuJD/OG720G3X7Y0rQTTDzFk2jU9X/wIn
xVQBcIfGHqnW0/A+8z+tI/hsFl/J2fF9MefYKaG3BK2JpjfVLn7M8sSxKN/54Wuu5+iOjr9U5j5M
Ocp3LTmGoCDn4EwZDSsJZXy/bl4jjFkH2G4ZnD39bhEonYFKfIAv05r9k90l2pCIOyY7WsEI7r7N
xVk131JximKhnKU2NPMzcXyzRKNcoVizbvMAx7Z2RN1jxYQXfEGzm/WkvVxB0CVDepZp3owIltft
w5b3n2I16tWK88HOON6a67N9nfGcqtEx6RrAnm2YCanCsaMM7+Neghu9Y15XZVISSe5ejTJEKQAv
hEaEhM90Q8MKZ26NoK603mHcvmzNIFqQfo7xMj22noKlPFxTRhTEBq8s+9Hx2wBHV5pz+Kw7L6GN
A7atsvWY14rUg25vhp3lRqCPBAh8fMsQpJtM5FeTGBULfu369fWCUS8rrCV73Ae8oCcWafD2eVUQ
j9fOW8wNHCbOsfwWK6bghoSNMMvf+kn8iW7JcPsGmIaexPRb6KPtzJuKvULM9MRLF/iKcsYAgoov
iRChSVAKkMVXBLzeB5zPJ1IaDcAsuqsbEAS3AIi+qoipf2kC4w7KATrxBovQFGgbyLv4yKCR8qh5
R7h8Gv2pBDbxoWcO4JesQMVd/4HwFjc/dPAdbtTJvYS/4YQnO2U2nZtQoWf3iX5n5ysOw6+NU4Wi
uwYEbJ9Em7o2zCDE4LmTwN2O2lDr0ZJdQ3xmsL8qKm78uSzkcXWwtPoMPSW6uWLlVFtvgS8OusrW
wGZwEHPPHXWg9m8x2gTyGkNtUlUjS1F+3dDfBrHUQsV+JCe9D/RY8Qk9LSS6k3P8QDDWpqQomsxr
2G7N/jMH2fUkrrNBoIXTxc+SYwsrF+rm0UaWTA642bA/fXYLL6faneP1RijOWl1b0WPBZB87eXE6
9I9abzflJ9y4svod+ce1SsLCN26hF+/xBvGzjbJGlqGBXbLY9GB8bunstUpsUJnsY97kaluSGpAr
bjYUqlJWapB/qolimT7DZOS0fphcEn/PBWwRwbh0ZqIXINM+IO76iEcjkFKqxftoNtK3SoAG2mqo
zxOyRR1EHaHp21Y+CZzbu26YwQA4d2wqA2tlWxBjUwAvwB58s9EeeqwU4BhzTWjjiIegbGKAtG4G
UeFMkdXPkmMSiJyGup1Qht21ntYpoTawvFOy1tr1KP/7ojHqUzsMmC08LtADgq5sUot5d2dbgCtx
8/HrbOwLHtDbEpO2fk6vEzI2ZV8mlJEyBOFznH1zyXAcvYo6x1CXEkDO2Oognkj+5akMMzE5NOvn
quTd0O3kwGz89ymgVoiAchvIGBrs4E785peFtCx/Y31Oi1u2ztjxJQvZ+lNZl3+2CKz5UZMwDy7d
k0fWCGNuxAsIvhN/TAYRDX/EHcL0XJBkvdQX6avjuiQlFzihcFerNDGMsReF4iwP6g1Phq71SXUh
z7SK9Cr7xX5HC/Yu7gfjs629gMX1Q3t5ktwuPhKkXUe1YNgGQ3H7et7DDvJcsdP+HgJZy1LSxGkR
ZaKZufset9dvTEr3OPFYxGSArFr4s10jpK3e1F4yVGz2Qm9bvKV4uSmOWo+ksSZtfb/ONeRB/yom
G7excFS8iuT/LpeI/+xA9UMVUm5ODwhJrVMoph9k3rs9gcLCpAY5U7p/W5J5MSjvXPSjmvTy2rwN
lPp9Ss3OYkDiRFZUz2qCOBip6LjzzJOqJTXN++DhIj5J+OBVeX8Ujwg6e0kpMB19RzHr2b6fr8Ow
uvWUQ6TEO3e+mGubMuxaIHm2vlPND16FNi3pT3rhpw35yWALcNvytlDE0WuOScWtEK1uAzQ50VQq
zFOjF1wN8oYz2ON4UF2JcHJSmiczdqQZCnN0U679CbFBfFsaf8TJeELIAgSOwGins9hrIP1wAh7B
4M6FKy5sFuWx9M/KE8d/f1Dfa/VFe3y/7jgMMT1Pc92+AQ5gI5AGCmfsBe7q7pLmIDrU95Cce0Vb
/73Dj8i3WbG7MWDnm1e6aCCHnuaHLG+HuvyAXAd1rSvUdNhzMT2QCe5v1ntub3k7woAD7Pkv7X8x
XVX5ALUf3M/SR8JsQcDZR7sfuSDh1Lw36m0zdl81xmX9Fqf3VBw1det0B8kD9ZEpbDVJ4VMbgHog
rL2TShUv7d1gG0idwGbeYw808+LZ/jjoyAQLt9rYaCFcRVMkJH72d0IeToj7FQjf3B+ateQ6nepm
Q+fq2kEBG7z+WSnw6ZjoGvZpl7V5DdpNALjFBkLTyHeuRX5CLFn2arwJJu9vFIPwumeFBtrvI8UX
2ZNJyrR1L+B8bG8FHJkAxCgkfgAtN+hKnl5lgMxqh4ah2Q/R6mYdiwQmE5AP3AGh7OF3Y7mXOdE6
8ZT69jYjBeS5Of61+GorY747yspxy9W0zmDBd8RylCrhuuN+V/43uHG2ARpuygi39cEUTTIi8LdI
mAFiTUuBnd/44xwdNch9wB+Q3T1fJNg50+DTr/Hr4Yh/BCA+qhq2Vy+8pjLCd/epPn1h52z2puZu
MY5MB0B37+92fXQsw49hA+KLiHJWm1UWouIiHrcGWKRArP4CwI2Gh2sa7GPmZdR9Wx2k1XYyCy3K
q7DXLp+VcHbKJx05uJbZzRDgaBORqlFCyHifPCV5TIbDTetDwnt3Fkr4iLBzMPAIjxUTkQ8SPjWP
dJyz+WiJaqOTFQRhGqxfHtWAer78I+NqdIr7uBf7eyCS+hqQ9guEuXrTCTmau8jIWMl7KkfzAvf3
FwAvgM7BQSeX7aKbvjEmL3F9fh+GJY+/nd2ct0qo/inGQSVkyQ01HPAupnJkq8VY9pZ5nq0/ntpR
yK/9Wk0sqnQNLR2sd6TUXMtgQXB0SI9AgjDHWcWXEMnTkg17SsOU92o9VfH+GtgVQNxD6ZRQlWig
d5FT/jTweJnPpTut+dMRRis6Zud9gxo/LJrA9zBmfrzfXNqxFFFTWbG5idRts2aLl+3yBi7/4wex
2MMx+6wCqUbAOqvZOh4cd7xaHewmr/8g6guVLW1BZJyLeiz+c9ugv8sEYSfX8QSEMvBr4qY+y1qy
fU/W6XeXQ55ClalmSqiBnvQN9BbAGLn3R7OS9GkaO0z0Uf+XDlSOypncUorF77B1RlIUp6ucm7od
AvahdF9tCRk4i9YnU5yRi06p2YueXc63eDyLoWqmzaCit9EacFxpYBIQAzMOZr8qqCdj5zqQ2X1d
q34/ctJrV/z4xiQfNnkrnkNVpRXDkIDB0CAj4sviqNKGolKZwWX8S2SIzKM70Powtl8q9U4rxyBf
4tA6y9MRFWW8oedy0EoJfszdBC3lRg1LoKwWDZKEXSr1EYsEP2ZZqTbMaf0++YVpkXdRog+xgzxr
XwPXZ2M7FdrGO5CFLsJrYPY1jXh9asAJ7K8eEI/pnBIaHGVMvgMxOWgSLhQKrL3NeSjBspO3miuT
VcbnE4J7YzMEW0nEiMD6nkWo9786Hyba5oioNOpL70oWPJXvCntoPn9Flb6cmAwOuo+TPP0dHLJQ
2rRPtVXRL5NpnqmTPSJPUSSWAnoIE2UAkWkfbEOkInIEez9DF5VvwjcWUlSl/Ymia3ryVWxmwLT6
UCmKEODiYriegAy+i7oFX0LN1asACxsmUgjc/ERyjnAd/aqdXT41btOUir/oLt/qI7G63fsSX2it
DDjTSB4JxOOvGzzSzSbVz/ReJrtN5muBF4OguhcRlVUMbg8Xj1VVsiq6SPAkyPacYFSB1HPA6f2E
FocQqw8Uc1Ioe1ZCz6eCC/eqQN3U0m1AYPkg+UGzikO8SBIkTcubocJNUG2VmdEu3efxspPV6N+/
MyPZIkHLo5szhIoF9IKZa2UPGEgTzvLQOzfIIVFq96C1DHYw276vpOMjzjXkuBUR82TocgPT6tGr
OnNDZNamtkfb0hVMo81/95oBJlUoA01ulMbqj4wAQxro47fJ7mOrfE1zorfxfvRbGuzDGWDR/deM
Q+saszWD+Seq+IhduYARwhIafa9YLINI8ofIpk2UZGDpIAloEo76XlED/Swsy2RUPBK9f/ikqmRI
yZAxd/OKrS3CQO1LsA/y9tGdxfnyiJ7J9THExcHf3iMFIGSmtxXMA2GlF5Hk0bLAsSKWLX021nmT
ulPCtn5VC0hxXsb8Ut0sKSX98tgvETf0hSNvpGgBjE3/TYkufjl+XAzqgDM044tJx7fzg/DjanQR
vRf+n+/hWbkde1tBySRThGeZjIZdJK63UPdmkIUc+IfcqSlOld61QB4iXV6K28sbpinHRlHoSNl8
DsYxmB1bmhf9ErFhEg97n4ISCnNl2QqF6U8dGpG/tRaa+xqCzx5SP6UXrFczoq1tlZ92v/QNn7/u
3yPl12Gk3cOHGMLjdxHWPtINcXFTq+mGuNhsBcLJNbVbKXf5ad1fnxXqCFXK/enrxjfkUI57NZpc
op+TGLdbutuP+Uk9+GCO8y+7DYkkN/noml7hEjzvtgPQKMAVWSilp1AXko7cCSJupR43pgByN83E
/tP4ckOOOOPorVqz94x1zx0aNgrZdNV9YEYLA70qhDU73D5q1h+E+VaxB0Sc1iDUg4vMUcH61EYz
qHHsCNVTf8yoYTqlUpZw4zsW2wsrb/ssyaMTiSwy7KcalH2IRW8+n0N6XLNe9NJyTBU++T01YQh8
oaX7JFq8huG+8fvTGBsQiTOmhdGGMh7hSB5XZ9dFXRa49XMf+CKc4qR50e3mZWbsYV80iWZp6IGX
JA6cUNA0B3YphKGHASkxlRHP/cJ7+bzoLD58szUA2p1YedQr2+4Wx1YRnbm2Nw57ienE236q8Hpp
H970akRRUJ1MRdrf0jPem+BuFS8oM5Zd4f48UyOfi0T7KL67Xo4xzkR/p56ag/QAR8B2Atum+5XO
wEbvouBhx2WjWGqmYOjydhtD9WK6Rb9KtdqpsQ7QBudWrxJmOwGRJTmCwgoPy40kXeH0zY1eI8Kj
e5KX19n4Pv7u1g3iJy2RFz3xUT2v0CQNO1wbVJZiRe2cxYkhoaj/yG0SRAKlqWOjweBCH4CmcvaL
zt1l77rNKTcjrwPX86kLrihalRxuoc7zDkdT13srterm3GjJIX2gS86DpT3GbPkokPmxL6noAbjt
hjYdliYWtrKFCvxL2LIpUXCd5cD3MMe0+/+V8JasHZYZ3GwqRgk2cXTwsgDITcx1mICNUiXnJD8v
fRatjqifU18x/aNzfhMFOJHLQhWaGIO3NJOdV12YL79GUORqv0l75Q3bAflKItbHWvrFUKf5waJt
sVw/VmrfVsvpu+NLzszNMKXTfgrA86O7R4m11CpBrKKu/ehx1+FhDgMC5hWYRT0bRihIZKuh02gU
0FDwQRty4GU4bQ0cyzFqEqDq6CV5mliBc5jw72NdWNvI8rkz+hkFZBRWxw7vX9poz6kvQngsy4uu
WoxZe1zkY/fWQbhgK4Dx2GLZcvjx/Vc3uWaXbjqyS2vMB3F5IxF85H3UFP86w4UcLt8PIL56NUyr
QO6RX8pBcEnRmLIOzp9PEG4l5k8K+QPQuae5mLrIGqOvMxkk521oRdMxxquvs+JicgHB39w8+A0h
/k5C2zsqBj5WN3GiI8nQapRUwPW0TBbjFxYpi3xsMIEbA7jRAO/7nN55k/ulrOqYuhw0gWoWmECN
ZEWFAl7WGADH7D48ZBmgVFCsbprx+rUcStusxc2b2dnFxzkyy6ogA+Wn6Fyhe28YpURKxA8cfLkz
yObn4Hf5uAp5XKbSNyvjrMuWMJE2cA9F3lgkUMQdJULSPrtAz8HyPvbl0GhxzHuDqVS1pun4nssm
BAIdYk8wNWGxgtEMrw2g4EZSd7+ve0xiqEBAlS1ukO6lOvIymozrnIUkljoAquxYwWaBdiEXbOQT
CGN+N0I6tkZL3t0cQ7nVVvO8V239QzLQZQZQmieNsGRNoJdkRjhklXVEGkxSNhJjHtUsxHJv84x3
kUHGeLXMgJyuelfbutxBW620jn9zQMDmtXmF283oMozdwobv2/Vy/eCe50Pd07EZpQlCcGOq3NLf
dz6196UOCYbdwR+VGi3TBJbZJ/ZXVt3or2Vx4MFzcWjbR/JvrRYIqHFXJX9UNsgSV5gS+Ztfto3z
H+JGvZCq9qYvSsRESBecC+QJiKGSQXT/sRThoPf12RIW4xwelAGnGuEm5q+a0I4DevDtmCKrAkw4
NDL5ypfXdxjTXxpoP77lfwKbFy3B8nFE2l2bIp49K8B4sAfZ1F1Q9eUhsPFjKC++MmHnrw/GZePd
JGgrNLJ02bk54aQ8Yw2tfafe3B7C4gK8WLQMQzEGGPJKk5o2aOAp8rI85Hvt5RSeAxaMYb5pAdp8
1hBEbrS9+Vj4sU+3qNnHRx5r6i/53Rvpo6Cajodt9oA0oILz0UYyTwmGG4XaLqKeIyogu642Md29
8szf5UrorHgE+KIVot+jwcXmPuhOY5Dx0aLGZQQ90S7Y1dwgzaT3RcMXxUIBbhFRWWwOXUP/Ye0+
GhTiUBNCUZTDDf3/EPdcvsoc/TmfbbEVyDHWS2tJe7Dll4FWQc95biGdlwEsSOn4taxuy57A03sm
6tMv2Xy7mLILZ1ctFXsqWz4olUzmQhkrqdevzbRN6WI4IvuudoMXDiVstELXeBM8cd1tIcNrm79E
Y1DEa4Qvur+BioHnGZosgTpyLxDvm8eArLrkl7ODvCHSv8B3sAC6MNQq73ebPn1UkL2zmhxH6D3t
WYkjD6NFmDbzeOHal9PlxUJXJMlTrbREa0rMh1Ld7OzkZ03d5sD/F4VhlmjUwwGbotuSgJ5ODbmw
ZgWK98D7VQu5OoaTIaYIdz9I6eOlvRDwE7Lmt7AZ5p8kq9kcqjc5makEWu/eD6+pIgYcPPbYqHkE
Flz42Vy+0QV1MSCTAM4WKE84hSJxdC1zGsRPI9e4vDXPokfkbEZdHUXgve3N1iZsD6CDT0TLg/hv
al+NyoBu58W0fcumNLRU8jLHbBpZbJBZ9JVsDZKXE/GUuIvWWtkN+qzMg3kkVCkwfNN3DuJfWNu6
ncXrKoa8F5esUaYrI1zUElnepxuXV0r9OiU04zGlr4LPKd9iKhufejzIPSFHPD2lPF9LldQT/sSr
g1+JuwW+6p0d2/yfb5IzQCMEsQVZlkEXN1VY3cD3YpK6HRmJySZ78S7eLWR3cj6IyGTV0sNPKB0f
NBAnHRm4W6emP4SN56XRBSzrZTR5fu5dAaIu2qExuZTAWRMkCeuIUwIHnYHuqPfcl16xpknCKbQZ
/pgPAkH8uIOhgbmPkp9X6tVWkw5FDnUqo6KhfESh599ihLe/97N4FRJxraqJwzDODWMqO3LZ2q/A
Uu2/WMX+TpMbsPqt2BtcSaTB/IBGmckuJbkSXUz9QjvHn487jVD/j0/SXMaCbS18mzoTfNHtCUDr
3rnOekQKb/+Y2crzFPvEvrYg0qgO8kZHOPvxjx8QfWOiG+3hNaXDOFpZxNAxcMMFXxx9nolroerL
/PvsQEEolbK8poxwwwUCn6QUu0qA0T79SBdEdA7qULyWrBno2HuwVbSfd0r+kSIromZ+KZGhqoD4
rRpW2DWB1CrwCouaxd9jtIYlKqGH0/JjI7R5/8GSLkHsqRv4fJzRSGXWDJbH42BlwWEAH+Raphos
znNo+NuS5NWJFDXpyO7yvCeWmEMwUwoRGYeItrTchP7IXBeVYncFNJrg0/uJK3RM1KRaWdLvMQxK
mbWAEUHHT6cBcCchDyuQ3MMUUCyrmeota2OY142iRqrLXXCVEQeZZZdH5K8PbxgbpQl0agR5dwqM
doTxdC5rODMZQoeQWDPurLKh/jD/CduE0hwpVOYUOV6DUxjo/T5V+r4AE1S3DQUiSATauvadYRCy
odMEiJ3Ae7t3+0KuUFvsjUiaXxCo0EGfUskXzgkuVLTBj/zOulsArFYFGHLTcaMAynSVVeBjGqXK
lrPIPV6HY2eAKA1uRm13m86JduD+nLb/rj6Y2QO7E/KuOuKq741T6o4PZs2TOg3gF7CVoQg9EjdE
/ldEX8SvUbjtn9Iyt5HWGrmkhqQOG92aP2pcAKDEzM5bo+DTptPFwhLzOvLGevSZKwpoH0zbSoJH
16RQ+41BaXx4nCiyZGJbBQG11AWCMM4xe49VKVx4mGTzAdp/W4BL5dMNBFDE5up99JVm8oaRS6E3
jtkUGi4TA2qXm42jtDmVGyDI7ulQ8TyoP8NM+I+5RNxvaYIFmoiA0K6hsun+sNk8DFFRs58hV4En
5b83xMKIxr3tz1qaRYOWhntK0fc1P5geykVATRrQ5+bdLaGFG2Tta8UOwIXm1reqlI1tN6Cthim9
RtfTtheqERfsE8lVqmgTARePMuOJ2aP1ursLPQp+cHy3GN5IX0xMLYXHYD6/VA7eD9OrqQ5YX5ix
HDJ8LDYJXBiI7pHws4htxZuzcfl0hYea9lwosCGykgiYxz083gb507jZq6cp/8wgP20ZcWNNxBNc
SQpIzYmCRk/sILBqMZEhHmCb6XtKHI6CTU2H40glmOn/givXRiuQKC3UtBi/JfD0+V/FoybEHl1g
2VrgHf5WnRZwSVP7Cg7hlKN7Mcl8LgMfE9mITY2az0plc9DKw6LmEPtdFGROPa6Oz+r4zbzh20sW
fUAHWJmQS7JjgBh5jMmv2EuA4b4cHEKZMu868mhzlVS8qIyLVg0VnidV26OEmC9XhKCx5KuANN9m
4VKrp1skXCsdpBIUNZ6wNpIk4oUAO4eLnVCwLLwzDC2871JrUAtVmbM/yOGELfjFIsLem938dj++
K5J7x8AA3XKXw89Xcc7iCWVlP7N3G5tRSR+n5fk0gWep/axye1X99fY8rUEmyOnjRhFIDp+jXXcW
7m9QkChPPtkMwT/Loy0orSrff9coe3BkZTXOA/aS3C/ShodxTQBX1A2d/ms9QHGCyayCbZ5oAK1f
KUQn0EL2UkJqPk/1ADj9is0UQOzgPmF3+izSvQ60Y9fppqE3HS1KbRb+aBMbLJ2DbDBT+kqMWPwq
gez2WBFf2OikcVEqhioeBsdZ3N9uaHjFggfKLpTV0yvVeIoOjytYyROg5AVTREWz5TGZ/XuDfB/g
wK6RMN/JP9QiVZn1/137TAkhmmU/MzShfmLbVbvgpHC2nOlN1fv9WVGfOClAY9nqnPZs+pEbzUVY
CJmArj3zSjNfM/f33xKSQ3uNW0KiU/J5c9N6hQUMeDG8tCfB0Ir6cy2eLbccA1oIVa/VCMmIftcU
QjwLxsxjoVVPAYzcZALkLk4UwyZemXZBvGYLvw3+66C1wDedC1hHuQrTVZO49/MjVnXvkAx+1Qub
5gEh6uQXRhvZ97vAQXURhlWTn8jm9EMYHzs+EIcdfYHwpj1wTUbv2Jw9fVGPVOKOMp0w7NbIn0zp
C5FatcQMYDfnzLb643AtZWO+0kwRBlwb6rY4YOtLXnq+OchO324uCiTjT3Gxyaxjermqiu95vyuO
GOZEgWCPtO4zDchDh2hxaJGQDCFxBo2hGfM2OHDatsaz3WimUVVP9IpCNLwLnWv5F+SQ6R+UHQDN
AaKlcRLD/s5jsWw4VT76hkg98fjnSRZuTP3LvoR8m3Dc1XzX6IJI5tzpUSZreo9q2v/mbk5tSY/W
KzdLhOiceWGWxRDNMde46vxLvdwYoIoiH4YS2sUZSgcX0It+/IHthJn/8dPlMtx8gmX8svrUcHnG
mDumRTbiAjOU9cf56zmt4WxWfbrmniywoaez7BFuogqVahTajkIrEZ8ZW1PhG10W5nLbqyIvvKXL
kpEVmMiGU5VQVJtNRT+/sdpJy/teNGbWM3S5qAamanc2MUYHQmUV4ancTR7mDTCZeWlhjG4uClvb
86Eohyil6KXSFQgowut5hBEqE3s5QfhNJP1NIzt8qDHpadl69JfUb6pw1fmCRBr5k5Jpcht62/bE
SUgKfMFW1CHbQbhY+hGHz9Q8hWHV8NvtUBUXkEMBqGu/G6NjOcHGLV5xEqU7EO82F4wu/n3QUMov
FhKrAbHWTbASoRpcHwTzInWnjx9CorlrhhryicyjZ2D78JM0bAZqKDGc1BxFZ9INoj4RVaBlk+se
VCF+thSB01QpTnbR2O0PMcEAUv3DfV4agiz4Pw/py8ig4bTwGrIBnq1gOV/DXKOM6SObjN2TRPCY
l5RDb/xlwIYHLGuDrLjr+CWafoBAEKislDrM+6m9vevPqE3ZNgPH1555RFFPYnITlG4+ogCFGScE
3vmaMqeMgTVbYkQCS2DS+qZCjsnRYocgzRzfgIBebzuA0Kdqh7SePNoynLAp6o6xbDazBmdeYC7F
Axb9jCikFYA0Nw4FD++MunVxZuZd+TpSkOLW7iYN5B64UiqNfUNTw4rOkGlYbjcj8W7IsI1Cwijn
uThZlcoKkRnrSSmE2ldfo0Q9IQiVmaTN8riNKTOupNVynexn6zSq01CB1pAfZo0B9KXzdeg38D0J
G6KRbbDNXTyF6j9NcXC0sWQ0YQrWT4aRSCrwZq/aOTBlHr+X/24Ar9LogOV3t4CXuB+LTrApgx5t
+hz27bux6osG7j0KqNbpfvA9OlkFTqj5XOelhsFltOS6j9UQ2/vQqF3AWLkkaJWOK1Vs7ok6GppO
eWmpyEXbLzcZAT0Iq3puvm8M0Ch+Rmgzivn3ufQx7a9gQWqThQufPnl2JSxY5zYh7SNFvW+lh6Vi
fnd288wxL98G51+cUx7LxjGI2SqiGUD4KBPwOCduXFShrSxZGpEbF0TWR5MvGha/4Fs4XW00OYV/
8mSXDfaKfOVs9ZwLVAyfXrb3QQxq9QrKXmSg8aWvC0eSC0YCKVcR+g/QHQQZbKrLE6zRPBDUyf04
4nFT/YfCe3bfVmHexzVmS/OzU/5Ijge1dk5iAbUUgG+5vsg7viREvurCmkN+7BUOCXzYM3taHy4o
d8siYjJMx5kg+fyL+YnXwi3mcv+eNd80LzJ3P+EjlFQ15nS8y+Se5Alzisw6adVlOyfMvDI0ni+/
IDySVj7fKXJHa7kX5rOqNlRoZ8tIkGM38pNJvXV0nAoi6SeOWJ2vQVwS2cc2122pevCwD7/Gvi/T
4GILc6imlkF2GVTctTz59TOsjGCB6gr1ZpaTU4bLZOkt+kiN6RwzCOR/dKH8lbL9DtFLju9iWIOs
WEK+Kn89GCV4DfBVzcZwVqJVOfR9TCA5sEUIDKOS4ty8NcikUkxfo7w06R2ypr1BKdlR3o6jfELm
EVs9DnTOzDK0rIy/fxA0d1zrLnpxpp0ttGAWovXFF8yax0PYnV5iuYgGV0fKOd+mMP/8OR2D0nIy
DPglLXIjdlo6fJxkMCA+ewrESn8GgDO/YwrYKXM3a3OjNl98OlnUxx4ju+kqgBL5KmQfXtUr/rCE
hHomcbHDXynk+lr/nF+B8YAR2HDLrGBPodRS/QMbRCe6tiqyIJqbxj+rVDu0VvcnYyhoBDIXA9R9
g1QYnN8wgKGw5Q6X7P+vFE/nUK/lnkOU44+Xrixcl+M7Y6TPoC96ft+9A3jSYnU/snddPVPfg7xn
yxF3REKw8ei4lC+I7mJVgzCT4wU4IlJR8aADw/KSN6MjKNDnZ+SDhd22b2zJ4B0C56mOapwv6B2a
fXZ5YuH9dvl/btl7qWPbIRrNQVgA+9Zsmcl3SmCe1EYklHzzDEwFqevMYqg9Bt2uPC+CIfoH1Iwj
z2yXDXh0efemu6yMiqRKWmsJNTfzahoyNo5IYBausKXY7nY//GqIU9USoXqeSm8/92v6wT/RuqXt
yRBh6c6CQVfK5i0z8GbSPwLXbasr5w3QbguXDgOjIT0m7WxKCczVje3N23DeFke0+ApGLamNb0fB
L8/1xeK/TtKS3IWmNaPwNDbN1IYBdGUIqsuotB2dWXjNSBEur5dO69f9pCFymEts+qTiEN2kj5C9
MSX1023ev2VU+75/tGajwNE1MeNsmtwjLbCRU3YIoz3n3Zy5O5P1H1midYdGRRmcAvlJcaBiMaY5
bXRmHWIRdPvvCKgfXVHY4onMi8TdFhrA5lO96mgLLAmAvVddK2+kdlz77qfzSommuV0zTx63mwXL
OBeVyM3jtJJqL/VMXG7o4YgToT2tvRvt6MLlXW3P9v6L8FsjBKo3ngPLOXtCzWc0nWiE09GjUCGh
DgealDr7wq60TzfX39mUdQtzPuFP8dgWdG+tm44bDzQNYzqqkSFxqGSpHFydUHMToLrFu6qKwVCC
3scnPUyRM8qPi4Dc+4/qRBM5Zc2hejW2EkwDgQKBI95q+Gx2E+dKJPMeHCmk+IowIPAc2fBZ5FUl
/nN8yo3jiDzX5oKbAcuNGE6SRtX4SS2LvA3nYFArn596HrcUH+YBsgaOyohncVv/T+TkuWlb4h+N
yIQZKUOwgihRc73ZOOBD0vDx5XlB9Km6Y0I2dVNfpX3B3gtlM1ffqzvaQW7cZnM0RPUHYwKFAIFQ
u0qWlhG5GWZwA/pCkY/Ewysjft+mPGI3RMTrxhZXqyjDGxivVcUvqCuKSdVyE+9gGWHsn6FVBJpb
AytPIarS7lbF+Wh89igZph1Da9SZLU+YAz2W/wc2T1LIpVZIfgWM7+ggOHhtZ7kDkQ6A72vARPO6
u6d81vw9Lq8YeSVk0kdO+iGZOmqYJVJofo/8yk/mFdJZ3vYFGo5cz0HhlKjZAxEgdwHFa4Pl6R9T
2Na2DEEgIyTOHc0LeWzSYpKkx7kstgAnYL15yM7SX0QDW6bcibOrUi3otr0OqLZbZaBxcCY8gdnV
BUixvfcpO/J0TWoM+iLH0W3CVJlVxLzTmK49q0+cOetb21uNZRoqBePfRmWKU4qH07cmhqJ2e3cF
7gU74RZXCXfIWz8O5nYcZCL6FMxBiFLc289cnREa0iQwqG6/Or840eEJxGFwYM+kG3grOtSKPbRI
OiXU3q/NgVMEzDX8UWsx/d64kMkr1Z2Pli4jFdRqGrOmYkNMOpcpboM5INq4iKpvrV9HyBk/btRj
rzWiJvVuOARkDSlAXMNlC6mBTiZT5y6qsmf4b912xQUFFuhzL5b34qFfxb+TTrDOH0K1AcObvJpK
1h4hC0EKt0q0X1qURVW3MhyRV2mFjTOVDyRM9CnBkYL0IgHvSvLhqjsYI1ZCSN4EQsAYfTy/2gXg
40f2dgR8JNd1EjScHlpPIV0GY8bRbuEyGtuhWV4p/xaxEvuw86bT5jARja7MSGJgMOIGw8Q+Me0Z
H7HPatHds0T+6o8a9UI1W7Lk5TxKjpqQbfrMP8GpWHXL+W3/OTpt+yk5n3uDB7P+q+NtUzEcBXiU
HG3ET7k4GsWpPth80Ur8kKbjbvQakb6A1xlldoQV48aK7u+SVhVZhhUZErskY6oFp1qWpwweiLOK
2m5pBuX8oXZlpW9vGNaIqqx/9zna/L3isQGeDFHQ1bby5LT0NP2xyUK4DN0NXo7TfkBkicbcSfHy
AEiBIX2Y6S9uBtg011bAdAX2UEAPxarE4ROsPHcUgGhVkxiqDfasTtV2H7tz3ODyHUipDDAoCzKR
N0ubL2hqhcBW3AX11enQUoS+dBa2hvjCxLCxE1PERFO/8a7SZqTBKfl/ar4qDXB9fpyQcTZztgSJ
4d6KImRUlHO8Qq8uh4/vOqPVtxMHyFpjBbFPOkwKiGFBetJqly7bmPlBzJUK8IPGWOFy6BfUk0DA
mu9ti6+kk1f5KYtLAGykEYH3GBIlE4HUULauYHmVtFPZnXsqB6bgVRy4xrE3LtVcMTYOvyQxvYIV
lDUDr1hxvtSWStOyQ9g2SpCw0l1RumUtiu052UGfe9zkuem3Rw4TW8+j3CIevbzbu5JJCZo7y8kd
7zxwgirZDUU5qQd7L1MWy+pJuAMxxcsjK3ELqXurAvGa6l6z8EDgRmOdPvbQpjsCXeSLRxZGYKlc
bXnPtYkgCS5Rp6G3kOAJel+w3T4Nbji/Bi6AioJp8Ayuk2NTIiAUDRD2SX3lmeiJyO+Ecz7trrtA
gD+/JNuICIpPzLHAhnyQGnpvigHaDqyB4SYXGNPoowlEt+jXkX3wnzqS6bss/LeNagQefT99iLHJ
Abqbg+k3HD1cpHHbfczaDlvchQMkke1wgTWQrs48Hh21TLyHvnnZZBi7ur35K/b7xZTlSiKfoNl1
NmlZw3OkEazUHCrvhaQWoJFi32yVWkN06jViowVT7UaHg06GdBmkoiD3nRyiAj4T/Fi4ksbtlDCe
0wxDQ8YV5Uc/hvDsTXOxVJSVtGaRqWgVahVdPgLKQvyfToY/IoypjISGOefxw11NkyBD3GkE0F0f
6gqW6YQhnOQvULwq2Uxa3vhRk6zEPgztdw4Fr2BdzlT5I4jQczjKh15tTqL7kH+ZxZAMIcwSUDvA
Z5o6qfM4o9klaE1HfYAwu8sjyEhXCrEk6qceTS17sVu+8PQmJXFnLWYWeSG/g4SWo8ip/XY39xFD
qFxZDKdHK2sGbMd4ovlEbLaoDO3XSdkw/jC2kL63GWXRs/2rxiWktQUSpeZFA916PsQLEkmECMdD
WXtZImbbx/db+6mZ7nTnF1cE5NJN9lswo+0EbAhj7kTV8wa2ZIFpgVt7qauOIfzanUlfk27ZJF8v
DVOAECvUNFcwlsqDaVAWT8d/NUvSXpOcIK3v8NTeC02uMohWVDcoURlITxm7Pa5X++jDlEk6rCce
StYROc7Ar69YF2jC7HnrBjc9cenSHJzrZcMnoGGe+Zd5gu5WzWF0kokV3cXkGpjr6ecd2lm6htHz
CdKw/KS3zH8BVoGX7fuHA61CL14k7mB4+h5/++uMp8wULPQ/KruUl5dedHiy63i8o4vvqX284SxP
pE1BpD0Luu6q7mxVGPEkdhdqbWq4aV5L9pM4+i48eHVq0B4MIvPP+IC59B/WLlk8spl8XAvcDhLU
HXwiTPXeP4gsGHx78UGYbXYXTziGBM1LLyZD54aBGlHxVvEaLP/rz708XYXiEjzy+VzSoOvoCsN+
v+xx5BaKKb4Wou3+oei8O8ogfHrEl1G1/rkd6XlwKTicM7l7491nUw6Vn2Rsy0+bW2BPX2eam+zk
rvg4AaZ1gIMoDtzAkXJOrwIhdVnUUnGAVe66wHu+C7MfWTT2Ibf5m3NWA+k4PnxQimVlPMMixgLp
RZWIRJA6aGVBwaMdht5m9y5GcZVL8yoImB8G9xeGIyvPwQwOKx06//7FAWE0papx5kvLe9Wn0uvB
MZ+F4ibbCw/Ch+K+kZUgWkPBncpnut5oPAnjfml+cVnkZk/6dXD+u8JNLup0jzfoQdrT/4Eqwgjn
bm+J02rnpnfsOMr7cj7/4bSiD7WX/SLdVRfYPgkbWNA0pDgpDSDhP089BDOVG6/L0/3qaJDYmEwO
EmBGV2xUXeExZV9LbfiAYOG8bgqb8dzUrCvXEgPAuLtDEtas8INTeBtWcszmPetT3uWbsMn4GqJp
xZOIe3c6Zzl0MteF0mbS+n60angDqcOu02Tlh6pgCYFZsmOq86iseUNaZiaukw4WGx4Y94zcklwg
L6Cgi+5Gbu5P2TtkWgPYBmnFUR62BrgWZgYT42aw3ttE8aRATxlS0ND7sBdblGLODzLWcpcNglFU
PUsoGWVXNgiVZcOieM+FkuDTs53vnGOD/x78vnO5+eUTrE6lI6X7QPFlDqr9OfqD4md8RUtm1xmS
d6eGuvQFX5nBXIXpxWu5lHJ5l2GFITDrG52BYrSj00svnvz7R7kqk32HbWe2gskAt7lNq8R3N23M
eiSXTpgxqEq/hNVWXxBoHnFbnHxYQG41Jjhm2Dv9JP760U6qf6Fh5MpWzC7X5KEP+OtCKjHnt6VK
Kgh/Cmb6bihTWp3gBd0sXsOcb2yxBKU9JsyJU5f9owydEAMNjkJkPNk5By1r8hod7YMUXieyHcuX
ZSZWhw0FQsFz1sGs/BlGBuRTDTJ7gVmcAZnj3yF03kShJ/gfbGDLs9V817By2F2O4au6IOiigr6p
+ylIaqp9sln1neWBCRlg+QaG5MAKKhT3izX05IOw+znngPxHu0umk01rktfTgjMKKjqMxpxXKTNS
3sH0MHqvXoSq8FrWRrGEl1DijMgplTT9hzsMYhAMhBa73QmTaqIDf812h1bzbAqamENFqDlOIwFP
bnmu6swHpm8erQocndE6wlOEZ+aMM0tEOFl4b4PxjCV+Xeg4aeRaICe8bMcfc47XnM7bVKJXHSow
PRQz7KHgHgW5UVcy489JfI/MBbCCPuqwfi2RaWeBEbsNWj6fFHm10XE3E818moUeyULVtOrbFo2g
1oeGoPCvo1NRnqxtDDbrNdE+ixc5LuV/2bjepTN4rL1YuyQhVCmSVwzXRoZBt3kBnhglPZPysIIJ
jUn1YO5Is4foG6O7+vZ4HvA0tlXrgatKz1g0vUSbsbcaJTvs5jvPflOTLlZunjjHVIeqAuMNaPwt
dpphQcHXrRvU6b5LYcPcPnoy2KkCf2eHCUmVX+cV4Ky4QNd0n1q9HIynWczAx+s++ZoyFKpo1WSS
T8Xo5hLBDOfPlSvEiRmQvRivR89X9n+y83xw+Fd093J7srRom44Iv7+nhsla/ewywW8Q10bl+H/G
ucq30RaMSA0sWfVcGzSoB9j1xncNz+HW2LJQTqAswu+VRa21+ca+S9b7FezmsItyyWD02vJzx5kU
6CHRutFyrQuiqp8ztMW2rN9iSL50NVUUP7QId+nNcbNJvwNGmGSThFA3v4eAeD2Us5bf6TwTuf31
CDj7+M5j+hBn1nyCFiNLmQXTkm6IDSfSDEb/EDO70/fGjrh+uhbirAWoFZP+JSVYFZcHqW04jEz/
96zQR4zKcpR2F+q5rDGQf/5vJSVr1z8UixA+Y1TOFbwxMVb1GsGU1kW5+3ttPnoUp8QyaxNz2gif
w5fIrPa753CaWOlFXnM4unnmrboe+w49qaGL7yTx25n0tamxpNFQ45gLk8NFbJpOtQA/m8DxUDPe
1Y3FWxzOiAIIU7Pft1SB2eSd+7jKPKJLoWP72WuE2BqhixbYYWv2jUcyxlNZwPQ+7xzE116VpDry
AEYJv24Epr21A4iF5T8pHN+EDtrtv6TBdkYWW0Fq4gs8/3ZmXu1e09f1+stKZkn0UHDy+bJji4rE
8eF8xDY7xFOlc7nxbL3ouSwWwFPHIngkQb+aLZzMbpebpkF+wvUdBIcKfi2jX6Xd2v0dlBsY4abR
aApJyFmqyDmBidhl1lJOgHltUfDkXFudKZRntImoCiU3Tc3aIWGe/W77SwlknAprKuGPghFY/GBQ
pH0SIR/xlTKLooubiEdSmAuUFv6g1DP9Y9fIcVcSMILr8A7wnjlRM7K2dqTmrrlt0jZoZejHfZIt
awkrBXnWJvaKpFB6YsxLsTWUumY+YuZkBROwiIKfnwBB4PUjL4YUq6Z9dLcpHVN3EHTi9sQj+/3b
XNGfger9GHSH7n/3HK7MFXF5vtRIbc1JtQA/c6vfwJGTahVCYLMnojl50QLnDHDHiqBf1piZ2jgP
Bno9Nolk+tnH1DVK7CIp6L7H50T5RvSl4ptKmUrSDa5BK8/NqM6d/3oHzriCUudRi60T8AYBK/9/
zbXx/cFxhNl6dHN4gJbza2j9tsT9apLyQZO56KZWtC9XCFmihPg2VoCXgtjhbIn4fbe3YtsHeQno
lBNyJJC0Qejst2nr7KzvabMX7nuPMntA7pRJg6R85tM5eIpLgNGLDXLtt6O5UwNiziT1lgqjn3sx
3Rb8Siq3ndHECBpne4UKX5JgymZUu7Hdwc43munQkDxhLnxEaXYkHhv01RvX2yA4DRscuNkzKsbU
uacp7MpDc7ErKLGUBTjd1Ykmut+o0E/kNgI1rZ4GoIh6V3LdzqvXkiivYm54jdLL8cYs6USFSO/g
OzLDmPm5wwwuxJcTz6Ws/GsmAfoP7xBzFsILQ2MVrwKMHeQSVHvuVrSwC6B5F+WO+RX8F/J10SKw
Ap7+sfeKLc8twxxumA95GZD2e/Se/smtoNlsoLXQEl35pcRcUhsdHpdGR3ZW3jBt5RLso+PZsFky
LHUrJBfwUNSu2+nlDtlMLRYTrtFnoelnoqF8vwkIpPTHChSnfaE6QcvCevMTEAGGGm0+RzC0KLbY
yfXHaIreWMjLEQLkPrUHe6WVIMb0Dx361Q62zEsn5R+hyVDXjxwnWD6Eq/lhAr8O34wcGF/PtdkH
rwQLMItShMF3vvUcF5kOzPxA+Fl8KBGPd0rxtgf+8tokkxr2yWLziZgwG5a+fquWGl/Gk/MYcmWu
EX3mQndz+QJ+uOpXV39aHeiJL2KULuhFJwyQXu+zcNkMn1bvEKe8BUi0zz0NVE9glWOSin5KHy6X
K5gkSfAZsVd2ItuN04ryTTpLDluFOsCg+iCK0ZMvyzDi3Vmy2gNh6y66SVW6Gy9WWLvorsDbquGr
FF1arJ8dLNUNvg75vF8Vd0s3hcEnWIIT8yUYe7jc4ru59AGu076SsZLR2NJv+DRggbIWbNmRSXhw
oXJps2s7KwYYHTxGe5NAAXSGhszO3izveFZM3FseDhCxuh94VLdlDE2GBzdrE4MfaQcK2nWH7ow6
ZGSYpWER0z37LDG2hapauaPB0FTXV0wz5KWhREyfY11amc4DDQHEgzcF2xaytaobHhq5NIJdm4cL
QIXZgee4Hgg8cOnQodNJsmoNFgtwBRdmgLiw0U7an+nq0ntkQq1nf6ahxa1FGgAqDsVX+/qxw4Zk
GlQE/y44eQY8TElQGmMQ1VLoq5TxBHK6ciiV/Pj5bEf284rXvR1q/mjx8Wo+4fHqPaGLlTTSXUW+
z4efXiSV0WrH8NwyNNqogI/q2MT0xauE2NJSHsSIBdbf4dzuoF9Wrasurn2CID98QH7u7okA7cGx
k2/eWkS754BZfLVv0dehwj1eGYQElMEaYlx4iI+1lPDlGoJsqqPpO9O9Q2vR46aINqf6pUe0ji7V
2QXiSDdjvB0Iyt4DsHzSDldviAgzjlPGHigr+IzHgzYM7bp1HgEG6N8NzBSpBys6hSrdSsrosL+/
x2vBMfvAU30k2rJbjBKyPa5GwdWDb2ZbVnGpmkK5PBgsId1kIKXy6Olic78Fv2E8h7IerYMto8lz
aXiW9yhIyP5IAOAe2bFX6wGCD47ewqzYuKGF/amAWymWiSwzUhiKzgz8qLO8mdl3o7l5yUbPf+Fh
LYycswux5RmjnlJmA8Mcnly2orcCotvplIlAEcnwdF4Evv9PmWt2Nry+ZVWzRFvijXcHxGsshg0l
Vs45pykSCFHrCquN04zv17z3ZvY7IvKlFRPubR4dbFdyMDSyQl8I3IqgojTIp9ZlDm95p1KlasoJ
xyFW6kiJLTG2Iq3Twes408TCC56pOxR6XW3mwz6pkoD1j8IOGe69F/t7oUzvBJZ4OnGB5utrLt9z
Do4CoeyCIPHCeGwRPIwYCVTmh7eaDk3MgOZU2iob2s0XwCDdDMLnsxClr2nZ74de78tQbHiDdkJB
YgQSKpWQRRX/mGEYnjOcy3+aui6PEfmpZj8epGhJLlHnBmeM1GjE84ASLNfw1Xmz5wqXxlHDqUF8
7ti9ai9Y/J6KokyHUWVfog2+RgYr4ypV6eO+w1A25Nf6gP/W+z4jXyBw/ZXxO+oUt6kxktECVJq4
Q3CKLMar5Vy4ExFn++2EO0EuT7nS/d0x68xJtzIVIfbZnyOvGXkfLT4FNNpRl55ZVB6UPCxhDhy9
pmcoFTmiVGTsVR2RkGzzS8KD4naEL48sAeQdrt/SfHnntQKWB9ujtb8cEuvtJgHwCYlAF/dJ2UM5
sxYJ8hU1fD95tSltHYROf3YCJ2aqrqiyVTY+SRLVi4cx+Oot9L4iU1adblVNi6KrDa1W8+uwZnac
IfmenQPiSGJSHK7S6qTvFS9tqj8o71ZVAftaMOVVycr5HLYoipFy0r/4WLMq+BLVbxNo78ukSeE+
yWGjm7qeeyNYYxbCbpdG7btxpcxCKPW519XKmSevZmyUhqSap2KeX5NTA0+tzIBpU//ht9v+hckU
jzOCVQ5rHen+jCqb20rkq7s5UaoXZGLj1ZCxMSvgGingb/rqkW8TT3SrdICpdnQGUfydggEqqNwJ
QgrDOB0Zd2yrkb6OoG9YqUVaLkegNoogW8UXBdD7N5Zo/sMFceH/ykhDLKaEfm0RH4p9KVxqow9v
73HBEg9PcG75weMjxWmry1RVqWc5QUkyHdRYL7sVfPbZZdYozm5zPc1IbX/5MGDpG+klbavNH/x1
6w9AFaY064ourNMmzTx+fcpUzyP23TkId8hQjYBOVAHhAtRcmuvtwqajM1xMIJcHFVcVhFfCx8Nm
B7CDJnnQqP3TIsdZDJBTXMR3g/s0Ds/QsCHGj2aosodjRZD8q+qXApQlIvWZNqXjCynbM7C6YFEX
vlzG2kNgXwC2X0kl6tpI0Zfsj0lkQE7ucuy5JOMpJ3XwYX/czPseGzrKYY1wMm4OwYRYm3nQIwj8
SQjZeEbhtUJ/qgPFGgnmQ0Q+4msx5Jzh+jZukU9PssAIOD4ymaK5oGfSEEjhUdKHwVt6yUDfdNH6
ZYCYiYZKU8jXyMit0CaMmgS6HATELcTzG/6ZR3Rv/JQ6ujt0UlXwg4Ua6R4SK0UMObXzaiV69evk
MDeVP9faFwlWCj4EpEYtR+s9GxH94Zwcta4O3PWT470W3Jjddtq2sjaoxMZokfsupLz/WvRlpnCP
v7RXUBsLm32u9fuAeVeAwosxxeigjDg8HIMCw3Atkd13yxop2/zGZ34v/k5PWFhEcgtl369kUjwm
eSDwoAL/JIxoxJEEuvyTfFXplQwOPzmpblWzl2oL7gEo3lNPSpu9NyTLBH9SYRo3rhOShwOC4i3T
kFeEImCWBwCPaRu8Bn+FH9wCi5bBsrhsnTSkn/V4zE82SkGPUY5g8gOvg9vsHB70iU6mCFRhpolC
ZupE+CMO+EteV/0VL0b44KSSp9oHq+WUHxOGpHK7KcZ+sNwgy+hH7+Ol5ZHmyhqYzrflL+K/QTha
1E7v69tVX1fCfXqGWV7VmGlXrakkMoI9p1K8fEUkHdnZZ7MQDZlI4iw4mtyrNmudqOagADQXhRHV
0T7ZRzujWtDD4xu3Ed261cCrj6vDlqvtkW7YKNpUh3LqySSZKiM69SvBnNDo0tSO/k5j71PuvnxW
1J8n6b02s+MMOzRaShO8beZPcCdjkWTgnwpwJFQ2ki22nl3wyfR/DbpnPa0pFigli0LksfhCrYnA
umX6L+A0kebLtNDMFQXYR4OV7bbBBIipMedUcZe/KHTNz2VDL9ahoPDaF5tC0m+INeT2nTBQ5uKU
XzWBXUZP6/nIiIGTCVBrVhbYBBlaS5bAfg3T1AgOz+HhGjOd3COi/SgkLR7btKFG13W9EQdduj/A
nWlv0H/eFWd1oco6tiImzeSw5PJrp+MSLRZoamfD3+4zg+SesaThQiyCUC6kmeKQ6kAgnZCZ7lEo
v4vIFcJgqdSsW2+FFMAbvMvTiLOITDrXUL2tfR8zskAqcAeJ1j+0S2X8tRDs6FK5M9KX0xRjOK7k
+e8VpPNXP2DCSsdPeVqFQp80DCXSHwCCx8D2itrJlLrvEabPGoWYswWw53dB4wvnY9FtDt8uQjd9
9eaX9eDz3ITFxKzqkSq/RdYNw7/3l+GcTmeVyXgmI6UosImpiYqd4SIAGzmrLO6vxW3Tc340RIsX
BTH7k8BZ0PYBs5SeM+6jAmNehp5d77rwIKKnFmefeUdsBgmWROtXLVGoxMQi0EZPZjb/UHkebTl5
b1SF5XYZv9a/xyKSUB39+qsMes0f2NGCLeGWyKpkOTJnnh8WEL/2XbIvSV4sdnKAZekaUrmnztyi
wUoHnwXX+HRiBf4tXVuWuWTuZsWejddPPmzbNC/wPwtY01zJlJFeDYpjGfMpoBt4cRAC0MPCkLHY
Bbfw11XBk+a6wRqw/KVNUMte7P5MOSzEpr9h1a4ccPyd29tmS6yl/bZbSGtt1GdUHsvskqC7uqHi
RgnciZZ9+7LpxJIcL4xsNZszOEqeHuGWyD7CjANapnM1kY7ItakPe/fbM10XRJu21cQEPma9bPoD
/r1CazAKhpZEO8Pahk2Nb6CuQCeLqPtQjg1FCCNU3oEz8ON0DhpR7CwaLUy7KCCaHoO3PH99LzOk
lkA/PFhG1bKFFFmFx8ILxKQecUmmDARdi3DRMzFXDLUiom9UydKAq6s3wnjSqn0WfaByKKiJMtEZ
oQoSPc7HIKGnGrDPHJQNlhWePniRhgOhrKDze0pt0wk0Uy696pUoOXyUbVktJ0vUdx5t7PFV7Y89
kxKbhRBdRLNfzv8ytrvxgxA/0PC8roq2emnp/tRPtLpNmpTyPmq42n2E5Uu0mRgmNNaH+nFM3CcJ
OJGguqgkrjwOfCO4bUxSaiLCG+QvtPqB+2C9Wbty+eKKho9QP3YY7zqOTFrez/gQIOvTjraDPhgs
irF2OE3fhBWvNu5Un5THhiaH587sKVlMREGLpkt7FxqrbdcKN/YA6jFK9AJT6ZZPzt0hRY+1V9vt
lrpdOvtBcqMap0H0cjF8HU/nn9o1+M27RBb9n/0UzJjJpq+D91YneNO0jSQfdxuHd5HW23VDDMhw
SQ74tvPsc5yzOh1osIM89dMqYzFOTkdSgmbDi4wfwaYzaJMrbcZ57Ncb/7PKa9EQzZp4+hHxD6a0
GGKirJO/5HJC6zQcuQsiTNWyPVKR+8xYQg0bqgCXUG5U9kzHKqCasoLHN7Sb47hA90tNrSRAfdSH
TX6XkHTtR3UUxnRuISligKFaTymHt8Eyttx0SSifrqKI34PVIn3pNYkhvvlOJsxIWwdO17fLp78F
yZ7wwGGvKLibuIt+X+XnwkiJZ037sNurLoqGyG9iDcSwT8FIp+WmxO6vTASwICSwYSEQFS883Th1
HLn+HiytdIMP3dVNt7gD0rrfaNSUlFiUzL/Nr3G/5zt5ZmXtsuefUqcESxgvEQ2CJZkBHrCm7GC/
e5cg8mSkqOfagFMlycGBhpC/zVSoNs21wMnC812/qUtNGBVlaGFRiFYGC071R9hmyUnswO/rRaxt
yIaQ0lHvGeCWGZwKG2nFsyN4vbB06ByyFP21a4ODwZy8o2z5cqLvVvbUAagWYtbdRZmxgWcpDIIE
4pA95J15jBWOuMmvYFo0oBsQJWRoXTlatTio7EcJdS6DNy7PyPjH068MNP+V8JnzHSdZIeTjsnwi
P0M5BmRfKmHSDgJM9q+X1crHUYvrwrGB5hnfqVyIDJ47bdUbOxgFrWfhTHYcyh6g/ucGQ5TNznNr
saSmjP2u7yVNQvvGMpGoeYNHks1xqbcv1kbAlQhG0tHvIUF6+yh7N28KpOckhx5UQuYOPJORaGI8
dYwMYLiHSMXjwvgWu5sBpMeAqKFy+wjnXPw7v9Fe2R9W/zPtKxXO4NMOFxdEPntomxcEF05h6nth
pTr0ifwhkj+coOHfIVyTf8mfhP7vMU9cE7JbK4lFJw64PUR1ybISUF9vFVrN6ZF2VMWnzafP4G5x
4YI56WEHL+CG/JQrjVjERh9GGQ3/h6DYmJ1Z8oVin5VIe9w3PQA8Cf9v+Wh6RrAJV0R6ORl4mue1
sjRYlBTijiza7eKY29zyhHZrSVA45dJOWPaElJVa+B7+fWlsPUGxIknNvwbJL3EH+bNgTjaqNcGG
DO0PBS5rbpvZmNbJ/yWDic9NNHSW1rbuL9vyfbn+0sqaCfpOlEXKY5O5t7yzijG/9vvCxjX42KSn
SQ5u61PkL/SGjwrmJMKkySB/bHZ9RqXoBVwrigVHYYG120S1dADtoZnNrDfpR2ApReg+LIUppIj+
q9qOgcRcbz9BJa2X3d1W3Ywm1w+0lYD2XpBfvoZzfn9HVE6QUXweihg7lct4RWXcFCb4CxcYcZXJ
mX1VWaZL/8xOI5iabteTyFkCjebF67PbFD8/F2f6Lf4/T8aVNXcMbOAtVjmGEOI9hLHXOtGvfp8N
+Gw6wZOWh88h4kkN1eTWPRxWyPG+VRW5H6TQzNyJrA/8/efR1yquP9yjbBF5poPpX70OtWI4ckwi
j5ghSJlAz7suykEVvHrIMyCt2IGGi8eEJJatHqFH309fiKkS88iMlkH+MsLhgWAh8ScmHKeY5Cv4
1yiccD8CKlGilDWya1jaA5EHOQUS+soPDhdgT1wBNJvCYe3egIBxXbY+wsEcSL1tbTvyfJK+Ppxd
CcghE7scCEuSPEGd2wu1FMFYZdojkZJJTEF8OozWIA7hZvQgzQM0iuBcheDurlUSHDsAB/3+TK2o
n/AaVAloM41d/6NMcg58qTvv0SAEQP8MUcy02Zsoct8s1QLxoj9lftJn9edhX2uzsCnNETDWJQOZ
LadI1M/KLrb14c+yWPjcRXif3sJ2t93/Vty06RwEnnxjPjE8xd435M+EY3acPMNG09l0BHyKHRdS
AEO5Sd5NVmYLG3NJD4qq8usxnZOd8Eu91xvr61t5LTvGICJEQIM/wwDfOnebyzJqm33SPti+Dgmp
KAUxMocxkMUzDnbilYPF2Kg4f1ip5qslsXsYzihbjvGEj7N/QK2T7TAhgs1n7588zotUQXrgPUV9
Cjo0odmTHjprQsJY4bXgorUOACttvDFaUGhrEI2e9jl6vJM5htyr8i6Qe905Fh1eBvekmREwhjqP
AekCnv1IQ0qioWgxs92g8xuV1Iym5H6qaC6OD8a8oUmU1JorEkyfiUM/9IviRY8BbNEXNdhNJNXj
UkuqlnOxx3o/pSO5pR1gj5Y10HEawQkkBRWMx2Z9MxH8gK2hex1bhK0iW8h7zY//WrhtHB/FMbLT
WP7FM51pZQ6iC3KtugfHD6CLsfX1MF8pOpuKZCwIZ/he4sR8JF9QkcB8KbNfBnMyyDYT3YU2sGIY
qanGiqEAfJqYnaW4pKGjLF1/B2XABup67JWat43qzeJDFkGrDJQOg3cnbUEhqrAd2z1oYaDrZCJX
UTWgeF3P+iUfzgr1JXFXePpdpdq/NVUvOcwt7lpeAZnpXkVHt1OlgNn+IOxsZmX2QXS4AWwFxxvz
EBNjOEjhkXVgzwH91KYCUZPqmC+CCz39qRW5ES0RZ2joTCYm+oM3naeRyyZr8AZPfOY/DSZtSTXf
MP/cWJs+gjJ1ol6qVdQivFm/icWM7GoSGtXX2duvyziy7OeV5NtpWANzlm8Of5RJCIAeNdOCtFO7
nU/4+vrRiZexNDDpFtIcOMXLb5rKlNPYI5LgdC92mTK3qgwvbJnM8Q4TddSfzrE/+mN5WLmHCELz
G0L7ys3aAcZ/IlIbkjq/DFIQziwpmH8kW56HrhxnGnNWd8g/1AAsFk1WCTwcGNu4R1viwSp/K81n
AXxyS+eliQYC/cjZV3yJJUwOoBCwJPQxhCcO5FMaRSLrPqp6pDWP9FHVVQ/YWcDb3HByfAT1Hekk
b8lBNqBmnmQIpI1mEdLSlx/oGKV/hn1bc+Bz8+SVegUOblVsEcWcq58R1WYGii+EiOwqEKgXSptY
tn0nJk241hvSPvpCEHPdE87lvZ3dO/l+pJt1W+wvGec22ozYE3zokpQrYYg0JW6FUB05DXs3NCZh
NFSB4Z92/aH5xcF6Z8iD0QGE/HmF4xhyDDd53HPcrUSxqOsXvs3zXr7P9+nvYBMRy5fJlTpd3GyZ
Y61fJgdOp4kkzqTACirZeoj8SeDKgBlKS9iayqqWw4wKiIRxY5IQMaf9nPN8udFLLjxmqiHjj4fH
3VGp8dzwRDSzJKkfGvNs0WypgLEPrHyTq0lLDMAZJRg1PMhkEF1sLhwpKrpmlaSKOPF4NrhKqKib
FfRnfzx8GVvN6Gd9/jU97WNpHZ9nWMSV84v8zJe0pTQip5gZd1y/KEnmv3Wg2IrN6KrPr1+XyNR3
cQVau90OW7ijz//MZ3IZtLrIYgr+o46yifMkfuQ6OGeUeFsaz57RVtEn7yulSZFJYEXa4djqUOZ5
YllqjlDKGiLLwNBOqWRysPCRs+7vFvx/rjzSVtdDVq0glP4f0JPnQQIUbTlkmO0P3DzO9Iyoz1sY
fTBZYZu6rEnySwYhX6z+0GFija/k49dGZcpd1QvR6VfEoDPC1CuoYVFc3JAAyESzgeCVxHeHb8G1
y1hCa1x+4M7TZ/pjyW9nkma7VGBzVJqTQIFob/i+5mm1jE+K5MSsKIZFq1/KQLlOSJtekRF2sJg5
pGwrNTanwhLQyI4kuC/Y8p8NP6iRuRn4UbI2wv730S8Zz21t/yKK8czvZ2tC2HZiOymrZZCjaFmM
p3PtWvlJVobF1NGHSYUyO8DUiL2JQWpjPC2mt5z+2xdLKGMdbvNVvn6mPIHCNRFqxMgOvMyI7hOl
2zk75K5vI6F9sjsvHS1cnaZ6VL56WRLlrq7q+KIc6DaMKgHvgNpJxZadIpNMcgc0C5rAY2rnULTL
NgAwa0hj6aORZzHp5jgfKrc5ZswPZpTv4bpANZRlClqgWxQX/45SAUmDE64r6hIn21S6Z/JnV5Jr
DHeyd6n3iOIjZ1xrlp0mRdifHaaxKgJBu1YhmOAPWtKK1c1D2EvJlpIlYBQ2Pe+1gX2kcfyv4Chs
404xYo5gp6iygQxoylgF6o0pO4hzTaVtbiciZlPx4u90qCHqL4VHTXRhoGy6Akf/a7/RlIVKYmwx
I4X/NTLqrEiL4Yo0FWPVTUC7S2llip1DpNwX4lvJs6Rcyvh5bj0Uvyz1K8oEf/Nd8Sm0abSvQ6Cv
6rOVRnT0aAN8mN87Gwho2HKQ37ZbZstzNO8TtbxxE+WeIT1PcAjEJ69uXOgtm6AAjo/FWUy22w7Q
PFthOFsQPrLH2RMypoGluMMABJ6l5q0DA+zmFETHV/htxQDvLiPTGfWvPa9e2d/NSI3lPLUs0iD4
UJ+D/h7leyC38cYh4lZJZSayaaadXQPrpgWgC33pSIoM/6xRIfyYbWyMBThcuVWDUfhamnmLL680
qlg+pxTY5SYI81gowvfbPn+mtpi1fwsfrODgvQl95AAr9YWAriku42mDxo5R8aPTZqzYaiXWmisG
esmdD5b5k8rURuhOWMvxk5roB/u20VwZY9SD0n/DvELX0c7hz230c5/VLU6RtBy1R89H4QgHzTD+
jSi370Sbs2HgzT2iHhH5ga0XZ//YYdNc90EwbYWgV5l7ZTy7tEoRTz0yS743aYGxmHnQdOoRUuza
uZGgkx5iyzTosqg/z8m79ysPsQA3+d1YJI1LopgOVFsUxCzgDlQjSztIFCWkyNavJRmB4UGS1uk4
i2MhuHOY6auJA85k6ZDRC9bVsaDhg8JfE6UBsrcuyEUESd6BPC2NYGTmnYs0ig0NZyc8TltWD3Po
i5VUgf79CGISm8EphTux1eEbu0qiHKhoQWZ+KzWmS3UZ56sptMOYEa9G6G/nbXqNaqBYCd0Xjzhj
YBB1gzcoh5VesobRSfACe2uK0EonY+FAOFYCf0TdYsVAg+p2y2tFJVwGsBzNpl6GUrW/qY7Z+UyD
aWkP5ZErny5Oyzc8n73L3gcpiv62NkS8g+CE8vSKyZYOCpslTZecUUXezZENlwKtZDjNsJHmKJET
4ox3hJ+uN8Ks0emXV8CZdIO65b/UozQ0BmM+crrFpW6gERjVmkyV97fVAvAlZuRKWJeeC1x74U2G
8pLwKFuQ7mhnhI/0TbVYCX/h7NtEkt1eUJA7sXksCtm1PMchQSHaerwlC+BRmWM0bW/bdBgm03W5
wXB0TNMbGYDoFJQUHCnKJyHY4VIJF8+GLYefZqODHdfefPzfKUqpS93yGZsB0wm5Vz3bBKkE3Nc3
niCKxMeYfYBSmgvJudfT2tN2x/nRGGAv6fI9wUSHsxuYWX+MAnS4bhHo00GsQ17t7C/dg5rnXBjZ
ex1u3O8JVER392HUzBPniEYlzHTi04z3jqkO6zKQBEJeXHDmuY0H3jAt7SdxsK+wQPzqEfyZpEdY
QHNBgbEeARx53eDkfQvq5UJwUMVKfO2gD/MlVMUYgUeMUD/J2H1OdvY7JTkRcv40odg9ESvYPfwT
wjHMDKKLe3T1XwJ+05JxYqVHq6XNL2lPoEE6ivupSJtufDDB2Ao25MqinKzVZVFmXe+jjvQhrRPV
P8kYrKpf4BDvXU4CibPhM4XsjkUtvg/dsOQuG6zX2r1w+EhTMiAyd59DP4fBriLuGFtEFlN2efCV
zIwC4diMaAoy6bl2qPSoD3LzncQ5Hrym5nn7GzmTq9etbzWPAhxb9Fvbq0JRzkSNt+kHWAVmZF+n
ZaDkjYotTWWfWgK3xkTItoVRgyFtZTKHC1GufCbRP1sTaXHw1dKoVXuyX1pu5lKNBqM54OXleE0u
FXd76oqCgFT+5EAOwNCd6ptiO20zwjbtz6RQrdCRhsKmSehCtal0B9iht8l6TzpQwEtE4qV9Zo2s
15r8MouGQ1Ds0ZYvDZJF1hMmGxOMc8sCnQaffCecNzMLb76o3n2qOHlT9NPVoQrqYjuLe6pqdgG6
SynUaE6U2B9iVR/gRWeZDpyB9f94xMfo0hc8DEhqAICmErxYqHZgnw9KoxoSoY01pvk2/Fu94lNz
I25ZcbQVdE+gOujpRbGn6W9SE1rrwOA/CokCO+zZw/oq7DOoaaph7dc1YAMT1gB9ewgwlLdNzeTq
ZCxoc54I7v3mPRlKk0kfDVJUkSw37hWAKgFvCVbkKrs6CMurRupBVh+QyhhXmSSFyroVqZ9BsDti
SPXELVcSsGs46SiU6nqGc3j2wf84p9xOt36f5HJkys3c1e4ya8Tk08yW53L2JiTQIbogBbp2ynqp
sfcg4fmv7cV0lkuSx/934BjFw0xMqCyLam2lijH5baG2872v7nQ9VcatY+NT2KZ1XuNw7eBkMeeL
8jIXb7b2MC/6kctl967WUl0/qn1ckyVD3/QpfRET+nimvhrhE/BxbOmiEtVIzicqMVll0miuLFVr
oJbUFp0mr0MsIu3W+PIcA0oSH8RKodUHimyDHyaYYbtvV/2444S3XnEAmKchwkVUmUftWKeV2rlU
B6hbWps30LIrO5EmL9vbfm8bPMUNYqf3FSr42e+EpzMKDPzOOEMAKrWq5yrZGpoASFyzKU0OVtmU
y4koOj5j1p9r8k0KR1YoiXxeTU7bL/gX1Trbh9tRSRMTffIkobpzHzw6HaBVxsYHnUkuatVY63jH
5wf73KgHuBYXt+nOQwKIUiW8sRhmQsKOCe48WI2u6EKtCU83ilTkq3UlYGOwe7xG7IYpURDcFiXX
AnupSEepik8ZFaocQRc2kXwGFLyKsUF++TWRt3TY7hZgfQvb57Ne/9by6kRZB2RkVXBuVn0e4Dx/
A4bABLhGg7vGHPo9RPEtZCvVt/co+6rC8ZBtW4QJ88M2LQiAHqzRx3+MbRoOVQM3CL1M5yWfL9+r
nbi8jEYg84vYl/0rM4USHSatJNkVDh1VM9qy7QtqUHTHP9zVG8oK7uV5GCu5bpUfWD242BxYtzNm
sVP2YCmDXqDHQAnmpA83lgGGJoWxgc6QfZNOrae1dTjvwkRVAIMUOqyziyqDuhS+z/OM5cNar6Y1
RfrOvPWFMmQEDAVXa9ENhzohpPMW3FqvPTy2EhQA5cWUGNz7J+wqXLxLnpVga2+wnc25ILvMB1E5
FOCCH+tVuAl93raACZnJtVC8BGzN1yxTp9TP6Bmf8eh1KVmPNbIGInOVkWcCpu7aTehSxuPyao/k
C7m05UifxbzyE0N5zYD6No6Oc9QA2386SJsVXqJdcypLeXd2bKrleUqj2mQC5rxDwfgzurRAXJMu
xb+yXxeG7wE3PJT4paXMSNdecfhkmwroJLAfwFAe6qfrqh4GtRTjMfbdExDtLvSGswHZU41+qcFQ
5VDX5oDTDTJZCNbALFv0GD+aTOTX3E80YefTzv7rqZP+1ZjJ0H0f03+Sqa4Xf1CNDQPyCaKvoQWn
qsSxee9r5u6mLTo/QHAXITL6t5sU4t0y2+0clyWvhoHNym7a/Cf6/p1HyYRa4rrDCBQ8TNnqjdFz
cgzLv/qsECbG1bMtXh9WPzATay5IC03ToPrw6iJa41lHLYYTHYca2/YAU/0/xEOLt+CsYKkysnpt
DcllBk7w+3ig0dXcuDeIhtU87lIDcJ68ZI0OqsRMdKu2fZk4d+awJ3IYOSsvCbUsFAUOpvKDiMka
kezibaVFpzvrZFfGnivzzBSSFrQDdXTMM28wPUD4XcB388IPGkgIeFuTmaHBhHREXFLEYnZ0wNGV
iiuDA31j2jcqCI8n7hHwcUf40GA9RsimOy+AcDhx1a8akfmttktbgEJ6UBRRoVzsOHrdU7AF3LOE
dU5lbxa7mBevs7rDxTBi0mvr0M2GuqLtda1wEKpZd7RxCV3x4z4SLBkD40BDZTcexgdB76Afixg+
dyCbq84ufbigNmmA7houNdRXhtKqEX2BMz3fLv9FMtMxmwygp6H4JUsiVvRQcmwzjHC4TUdtOdyg
svIGvQA7DuFDgSu4CwDLQbAeBvek6DrV0bv48rEmThY8u7Kjaem/KEjoSkJCR0Djy/68bysHw4mn
KmL3kCJd3yrL/Wz9UrGxpymC4hFANeZe/r82F2an+qXLBMfF05ckYBwVd6AT+UAhDu/RU9qujTUt
oH4R7GWGLvjYM/dvK8jDcdiM1t35uxNY2Gi59jcNVip26hQt1gTaowaeWFNuTNyvQSCFQKVX03bI
TUweSagI4CbEznJ3qmVQ7UNElWq/j3l+zkg+HzwV0xpFWKTqZ0+In+mMe2O0BKUPZRpqpJYFHOw1
gBJAOGBtqQfymIzIgtUnY2sCwMy6MTmsvj0tMsLeULV82uOFrGIPfSkxvfwtRimU2Bxpth1qQZP5
gSfSLpFK3/7kKJNn2ATB2mWFitAje8iMSdYL11GdvCJGPvmw49jK4yTlkRyiuIHhnx6BUPxhl06G
3X2yVqD0kqAmwnlbPwMsNVzgNh1wg6BvQdP+lV/VxlCEtAe8ciMFsN+Q5UkCJiUMd3X+n/KwmvJ8
AaLANRRoDrtht7Y/+jO4WyO6+up8g1YK2/Q2rnY69dZzGylC0O6Jt0NtAWecxCsBveRZaggPzVvV
H+gbzrQBLrPafDCK9YVdXqKqe9N7A7PbiLaUmoMxoyfSRPV877bmiQ00wL6u6Q0fRPJq3l9IJ6HI
M3UV1Iq1sJJyJtjL/Bqej5oFJd7szetNL/8ahOt67QGs/OMQtlDuOExWX3slWVqBVBarCmLQ6M6o
y9DWEC5Mh3f78e0YwOuhjAQFBCHV3wdJ8kZOzL/WpSHRi1UrzDWDyoUIxy7CieA8IRg9E1tEa4Y2
8yPVKxDKRLAp7P/jnacsdtXYMcESh5cLXqsxfoy0xRJrMIG2bcpIt47MrSBRsNnxQ3AIKC2DwnNB
RkwlHaC7X+1XvFtp4Sqp63YyLS0p5TLVoX5Dr5LBLxi+JCyJfXZZhCByLhZ12BkeD7bCHqSsweLh
YGrpGp6Lwoe1yj1sHRLIhLTf2vxe9Elr2PhG9qEFzaA3YEA7l6d+2zpvz+KyUt0tSJaapx7f2p+4
Fg7umu7tDF6NODP3oeOq9xUjWd8ufyNfOtgUcles/1hI19P1QJoEObPB0c+OCGtbc5lt4XleMrOr
Rf975w+mlMHvcZHH8g+Fc5m2PPysqIXy4hEwWmFt3DOLSKIflqpS92iZCj2Lu8CkdFhaJHSnF2Jn
SSRzSqLpAO0JQIQP0FTL4ouvCr3bzme3zmZN9lTleY51TrcXWYpXd+UehUDxhiDaZGWVidsDXNDz
OCs3JKtLSkiJZJzf/fSrKY7yy+Yz0UZlzAyczI7sCt9JqGTkO1JnNXBdI8lz7JbRibf54uEUOVaa
CqnBBxkR8ddJzivNKgfBh0sZcgXwdUImgUdTIZOkhC9k7S3TNSQVolAq65uLOc2IYzB5eAmltacn
GQgxALQVE/daXHXxQ+w0TERPX/k1sIDsLp/vevbMHH51KVWatwGSpcZKfoU9fv4dXm5MxPFVyGF7
tZ21RRqSU+uc45wIHBPn8ih0Pd+sYBxIRCXNOGKsvQaXph00lFiL94WVBUMjQ8xyMUmqEJFXXPAR
yVxKFFPiZi6tFxLyks6jwsoWIzi31SdBphbyHxvAQvmUybVIy7/jcXXgFCDu1LQDGvBKDfMsFIt5
Va3QlvcdIxW3HEUiGDqFfd4fYphm0+t0jJVwCORTsSBTpFpXQZ/ioYsuqTihun7279WdacNrOJtF
mEPGx7T4mqzhr5ADDYaKqeMQ1ywk8dkWJuGreI5SaX8donrecncPBbTbGTPEpmzB4CrBAMHJq1hp
gj5tJCEejFm3E+wrgzXtmJqICqzWM4imfWVvHQNcPxE39T+79E0HtWZDASrADLxgPr+1L7sN5u2B
ig2f5kyH5LiQT1b71dbRDGggRMU0xo8tuEeIGzTUstN0jA4/p5T5lkKE/e6Ui/1XJQR+Ju27Et2q
FO3Met1FXKhtpKfcofOzqGV+h17XRi75wVxARCnjXad+nYK4xgxmV0fZb7UE4SUdYKJMrME79V3O
UimJ089v3+WYbKrgZBGFyus4Qo/2K9/ZCwxESupUSX+LF4QHnjNhie3+hGdmObZk+2i2ckxdyu3Y
X0TQpF8ZSkSF3ddX4BzZjY6QsdvpYFF3cAd5GAEQcN6Nl2sS9qjcmaBBepZaxmn0Y2Hvg7T9ye44
NpWf6/M3wQvu0S6bu/+B3WIuTmbmGh8nYyg27uQLxLheeBVepGuLgFATQ2uujb5Tm88zp8/udjc+
Hxg4P2GsfiExJD+GOThV+NkJfycQNqrx1sLib79/4zH7Cu36Cry9PXLYfedp3P/ddA2bxaZjblc1
6leEhaSeeE2EzDylxP8FXhLlKlp8iabdD6EU+31cY9kqpj146n0PGM79J2bd9F+LoYK3LjZxJZW6
FpXmasnP2WY07Fts1THQ+7NqMO+KqO+F+qFJRw2ETlJxRvMkLe2JPAOq4FhOnK/svdHB8kyZnfXc
5o41rd5q1dZN1r7T1yBvJFtlwtgSckX9vpi3XenTfLQ5ObSX7/BlaiidO9n6guFnXindXBzpze+l
HFSAMpbUxm7HZmImYDaiqeW3v0laXcw13KL6EdH3UnHL9DLlo3Ut+jaUAeC9ZF3J9lGdwcJcd+4P
77S/s6Nasm3HqfjnYI8AUj6vl/gblZV8krfu8wfxkikDZmcD2Ae7GSHzIQicpyTj7WAw4bg+loij
e/wVqln8k2ScNPhcFkfPDC4CX2OvrjKh391J7WMD/oXbbFvRZG+iC6neVHU1st9Cprdr+ElYlPXE
QKXvUNk07EesnXklI5R4eNEafECd3uTugc6QgNoX+x8fnI2kUnXi2/JYlwCbYkXUearOPuCOlkuA
WT2OgGA0S1V+jEICOKlOCPdvEcffvST1BbEvX1CYtiNxO0rGoIuPO4s57K326cNB+jql8DfIIBRx
4RkH55vLzzBuUS9nOIA5NnCLMzCXCGhVjh6o7gO5BXbAmpK+gXMVLFA+38yz6kcIO3mgnR3AB78N
W8ihhePuQSRXaf6Yx9YYpkj8F7r5AQrvHhAymIbeJRygEq8Lhj4nVZYBn6JpR9Af6dyYXokRn8P2
t3NkBeS7FsVnGBklEl6UIK180Kw/YpheHnRcbalQ6FG/2NJ5MnH8KfTuX8b7SeLIHGxwjXeH2DmD
B6jO/FIS1l1INE0SrAvPpT9pUvE3TwHK+ohXObZfEOTp7DgELa2cobkmGenyPuUQ+4mO1PZu1wTB
3wITHSRCdPmupw3f2xUxV4OXVpMy6Cfn1Nc/Q6VzjgYLLw8Chn2d9ADflbQh9FreZwz8qfK9OLKw
E042/w3TsYZqQi2O3Gr27Ll1Gzvtz91He462pyfuX+kT5z+Pg/xreR6MZybWizAmJaqSi+6CEAPl
err42EqdwtLsMZhVH29AIPIZoF5cox7yAe/Y/Uoo53oThdg9hZ2Xf67D/rgaM46r7h37/ts5m8/H
27Wm8Z/mbQLphVZor7EJ678+ffQn9pCMUxxB8EXBRuBFZAPWLU7xLy+A62eT8mnvjqORSlNI2Owj
ZthaaK0fKUPT6FrhScDHSCSCLmmfBAmgOPlLU7c0z1zWr+hJjc89C+stOraHedUuj9wvdMh9k3yz
5fQk9XwTwAxzyXpEKNVg7YIWgxHq+mT1C6Tpmaa5nrfBzy4y+MxjqEZKv42gaYSeJO3qA4MTRbM5
jownrPddtRtoUuaALiTESZzYoGwd4UlPlgvPOmvUTenbKllxLtkPcM4urud3C9XvW87em6C76oAl
n0NtylT9k/lX2Wy69PWUTv0wgYI8JKMSoEi1LVOGDJIQZbdlfetSK07Ql9IZMG1BiBlrWCLyq+BH
8qF4M+hOPlM0fVcI4u4qkNaXrdMsqzhngzROJtdfI4i6Iu5oq/e+niSHrqozpuYo7q8rlRIqUnCW
lZHKCRJNvn0YzNSGlTA1cHF65AE4mviIEdGVYkxDbHH1w/nu80bTKcX1kZboyLZtCc55A1jyYZB9
DygyCO+Mtk8a1bwEU2fTShH+qRc8pleTIZf38pxP79euVI0aBTyZ7kVq8+8JLwahKVENkAH2YsX6
v+nx5NJ686Rjbc/DAuly67e+W6TPA/zNjCa5x/1rY5YV0GIrO9TIyzttMVcZVwQ5Z7YY81zWwCwj
+zk8t5SDQneHMf4mwuyQFmJsW+qjwd6AO60fUTcjngQlqpoGQjio3BTxkF0wiTu49on4s8/dVD7R
03ollRcs9DjVgUwFs2SrO6bAx3IV+WckLXWA3SDxaStqu7VXwO/vZjVh/hyTn67WUOYPW2AjTpS4
WCTwB3NDAz3YjG74XpYKIJcIOJU/0H0/yGRcjFnsScgjzuZma2gVrBG9jj7tQc7L5rX3g4eoJz44
Rf+fJwjoLI9LjgcKJpSmiW4HKeYQJ9nsUgiun86OKZngIKzI83tl9UbYCiNLucAB8ntpEGWwrVzK
1WCx4bOmf6tbfs89eT2QYmnXFix9FUIa7nCA/KNonV9v5b759bfzcJjuW97qqEarbrOA81MC8GWg
lbvlVEGuAsicukquQEI/g5ZIsNXYPi/n5I8Fa5AgIBuA1WmLZYt/2hN1OmeK4+s5OVj6LkmFH/rm
geK1dY5h14/f9EVhryf/GjtkyCqoXQrhsWfILZow/5eIHc3tyPkPJlmigsNjL9TH7/3kyYBrncJ1
SryfYLrFEotziR5xaNR9nfm2+OLomMxrVpbgL48ZFvu7yu7VJ2qMTGfqdtqFjkblGDGlQngWslKI
dfy8kOVlg6sTF/k6jSp8NiczIyFWN7KxWWll88ugplAwxTL13fQ0fjsM74iDkarbeuduunXOw72v
6z/Xi3iPC+AkU13DCA/sPZJre+nEwkvqXvj1RLWyhkiJtr0+55Mr/4GwnyIgsVeu908o1hDyxUpg
rpePrGGGJcX1Rs0erBVD2+pUYHG2ioDeEX9SaTFIGQKeg02C6kmReuPX3hZYm5bX88nZwqqCLWQJ
0TSaicV87H+tFbHk0mAqyP7ORc4Ukl9UuEkf6AmebEZHl43FHbnPwIJXd4eDXE4Whx2WTVbgHCQq
MvL5BcQFlu+56RZ/QiqhpVwqXsR7sDKsYtwPuPsuFPQKRZ7fxvscQTEP6bKNJpaOTfboqjTCOl9l
TmStAWCCd+ySXWy5HhBgFdy7CeJWGoy/Rq6ps6kZphAARV5f8VjDGidgIZBXyqR4o1jfawWrpBiD
in7a9mdcPE2cJG1pz/I9isGx9SX1oJfbvYG1vzIWsetsppbB7KUl2blEVlfLz+k1zlOc7+hN7Io1
vXdZt89I+7B/hjCkRExDUpaHMJ28IXpxJP6nVJbnFK3PZja0/Ro25AN3e1SlO++KGLGbpd9iBZpe
IBXyShwsfhKBYQyqS7ZFBEyP22bPzt9RT4yZpWKCcJYAJiNg3vu413LP+5ZZSengB9ijAvbNRQhQ
vvbAcpTHpfjk8nPvoyPxiZ2SINTXIyZjxD9bxr/JdC+PS3xhEzsIuerBUbDmDxJVRDg3SQQBrgky
HANMr2TH2mcYCJFqKVcetSq4MJcF4JckXD7InrtYOp5J8ED5VyrUBHve9A3IOMTvb14H2TB6LdJE
MWHCH1tLPsV2LCOJJGYsMXiSuxoDuzHBPar59gqBv7sePyPDHfe/Ir+S/YNe3anv766+zkwKMCKk
uOssKGyKBR3JO33Og6pdzCN1MNvmRezH1GP2eUdGtxx7ucgEkV3HDfwXgXVXE4VxgwCDrUsynOMV
H6uCKdujWnGGrUlczhZZpMupCj/67Hun6wNymOF13j+jIYh9lxl/yvYNQe4oKX8LiR7BE6cyPDdJ
Y0b0Ln2Wt6BLs6PE/r6D38VOySLgoD/M64FUNkJceL7q88p9Fqy2Z0CiAPnp4w5O94Zv4GLH6/fj
En1TLkYXoVInn0RyKX3rWYNoBOZps2cLnkYtZpMLtzo9QIQJaRhGlK31gZE3pc7p8+d3DS69XDTf
/JcyWqLEhhbKL1CJ2fBmeGsoFv7nfsVJxM0yMMwpzOnnf0Y9KnpcrBNNPFLSDIV+jnktV/Vnb+Tt
ywTFqChglbxLAnLOtkxnRTfvnlnI3Kr1Y/tE4wPYSn0G09OZIvbLxX3Rf14wHXgB84rZL9v1DHtB
jwiZJLJ87H4EUfuh81Ym5utvoomHj9Si6wUbLYEZ8HVW0ejuVrFu8zCcpO5ZdBZND1QTMbRVPmoJ
d78pZd7EKDt2FfO+LhDmRyNtlfmTNjw0K+AL+D2Og69kKz0jwugTBNak9CmZJQ2QcXgCgigB2CpB
qd8k4qVFhma/1qlquxy3wJVrHSGs2eydTNelqL9bOyjtwi8TUulSJmPfuyFvZf8TjMtAhPj6m34R
i3+MSuPVo2aW6dGsr3QPeNEsCYOhLn9X5KaH0celebkw4L4tBKgotcXZ+kJTSnp5+pocHIjXWohg
6lNJXDWjUKSZo77n4lrroLEVa/h0UWbejEyskyZicL1hDe+uic+DF0bvPTgZb+dF3JtTfbIoX6ef
h653ysZKdnJAWGEd7O3SQ0otBDxYADKF/4mRO62RRxzLzWNlOOPquJzY9NJUPaeoLmgm9OLx8gfL
hRwzdB0ymg0HvNKouHyXIdEqTTm6lAxgimgrJHQno4O7RGfqqbyRFgxzys+c4lFJr9QEIaC2rRsd
k+a0zfINCgSpLW3SM91+hZuqsay9/i2ozSHR9QHwqR4rQ9J24g1lBt6Bf9wfhiOSXpzZj3uHbScM
E72NX3eobRJ8gXtKq2CD75wgmpUxKG2tJ2m1kUUtI08ZfRgnnVbRhzyBHH7OuMt6C65ykCHscUWR
Hq53ACN0dWKOHlhi3Jz7fty16vYHWOKivqGNqMw17zJZgRAqwbve9LPLEpbpLmk39wXs8cB6JF0/
I+33eVDt8I8cYxW6Bz6gKBQSAbFwslgBDIQW1hAQCJLKmexEVvFq588kLMxczsKG5iAU1n6LbLM4
8c57Ewhqs7NKEkSvUYdrS1tC6UyjR2P+04InR3GtUyFfQaFnE6jYbdPodH2jfewmOBZn2MqzyiQ3
StTNrQiwiRfMNjYezACGmnU/5yXHSpQz9JC3nIp9ZsrUgtdaMmjeguYCdDzVSHoP9MqaXlzPNgys
NPyZSd97hpaVVMUuKIOwjalgYylmvrya7g4A4lChevevcuIBhCBtkCF+I0NC2TLF9OHOQ95p0VbF
UBhu8DIYUIwFeQlwElnjG1YKlQzxcPhgFJ7VjKlrT4ue1Qa1oFs3HSQajTdqTSB208FgzWG1QeFo
oQFRA2emk+ygXNwcEkUcM4MMCHVILaUeVo9fqRJO/ZvmcSt4a1Ft20uNQMAVv/ap/I9wtmxP3X2X
YGoCUSGt/JDtpbXeg0pF4q+aOD46rGVFDITfyTd1wng6DV22dkERvPxLo9PLkuFWUX1Rt+dAx0sT
lbkOi9TN+4qybE8mGR8v9Fd8wKW5FW/YOYpggTzPJ+O3hsCgzM5teS5SLs6AVuh6lS0Niu5v/hVa
H0O2Im2mHU5vJLvxxxyLAfavJ0a3QGczR2PrgxZWD607eJQJd2QUyeMQwzoPbstFtkXARAwaOg7U
hQDWW3CInf8mxCLaevoIuttJxFc0ZZSGCY3UqrGW4pIyPwVvVc7XAf07Gcd4I8j45iZMPSfnXNoZ
k1iWTQ6TIkcUNEOG9fv7qoOeM+wZ8JhjKtIV1JpwZIWt5fKi/4mvuG6qcK7BENlThd2EDRSeRqni
/um6/hsU0GA4qan/HvOQOch5Taf4sJd7XH/Iz8mFPbAZi42ZLfHpcJAXlYpp35/e1uoBzKSCsFFE
uC8qVC6iGZnNblIz5im4G2UvNGX5eT+867SvPrI1d84hOGjQWer/eGeEOPoIR8CvN7M/Eq3J+0Jz
Xy1kzzvwcabvcaYwhqR2bIx8wKHG/lKHe/ErGtFOPMPBehX/pLBgKFzqjdcZLNd3jFXmw+zSA0yK
af2RWzgpfVdSPSuIJBshk3rDHdD8RZTOyNIR1si2whBo4CN7cG21pOihSDMEFEugraSqGoVg8GMb
qc6rXPyKbZ7JhbCBeoeMnAGbRxYfKM9reWSiiFv7EoC+AhJRi2N60fZmitaQ/esCJZm2yJpUMHbR
T+3Zr0gPu5LA2DpKgO5229hfSaZ3IURjZHpqPf1Jd7daZVxTDYmjuVcrwgz/UfFYQ8grEeg0kDxm
yssHIWcsgMeuyI5QVkMrc9SbpUmDkciEEtKh1av2SXMbYzGZLgcaitRdkuxoTjAJ/eERFvp/vonj
iNHPY6yYA4ByuQS9uJ56lV0+WUmsjKND0BwcxLUJTu2m10nfiEF6jdhk7wUHb1IAt4xtYJ1hB6Xi
K4PC4BBiXJwqqNym677OESDthtnaOn7FfkvpoBK5OoR87TRIed/Smx87G2Jc2Q1e2FAiPuCj/gXM
4lZdeaGOobVCa9q/COTG82PGzZoa3EUZqkb2tgZrkk4RMpoHtdK6KEctsl+y0x9r8Y6K8/0qXBuC
4riUZQ8ycEreiAKVKkyu6BLk0CCr0sTY8BS9+AcmeHabtXMCRYlr72ze5EVIJE7e9Pafel31wVkI
c6TzdCbVdxA6fBy4wkBrf7dU1M3OGbN2bwlQLZFf+cIzzTnVKPIa/odqKtsTfIv5lzHilIEks1Zo
oeJXIaTjJoJsRDH1yn1r7JrfNdKWkR34mH+eTcxUHDICKVEpToS+UUpj67OMC4XC07UEtQbGMi6k
mxzP7IAmtD/gDHKEXz4Za31msCORWgz1v4NeIB2WAw9+LB63L1FfS4jkHCkhfIDZ3tnqdf5bfSVF
PKLcteWo2SsakECLW+ToEsX0cCojfaqsrF6xWJ9r+XaYJxWAEe9p08MFSAzvsLZ1cF6dCtXWKI+t
WAVob7AKQEp7Uz345pbrI3NVo3HO3fJcPgmzYXYiOLQFdeyP/fZo1vOTGV+/xC89KD236Er6XhXQ
sFhbl9v0EKm1Gig+mg8qn8FAXHTod7Ca5Z0LH2mmGN4PqsbBfjhHbRR2s2ZuA2eRXqw2J0q3p9of
8pHvVg4de4StJCzPNpxbG/VaOGZ/FKC/+/vFfLDL6XdDQe7smHlIY1e+mKKFsx58B/PD/tvNzk9J
SAk8SKE8tTCX7cSPVSD+CaNj+AGPJym+ahQ3pTmpt7xbbVRm0GXjrvL0Kcc0yG250JpW3UXD55dV
KtKIZsqpa+Gv9LzyWGvHf89SSz+gq6BgHcIxK2L/415wiqUtAi+75v4w76am6wdrBpdkrWBbG7Mj
E8jkSVZo8InkTK+1TUbaawHtkXbkslRvDAebx3C0GQLlrNn1pWw/nEUxK0Di/PBDZVgeMhlriBSu
ywsaa9kRoGHFiQPFbORCkX8JU2yvehcscbGLSUQN9g/40Tu3MWQaeESkPTj7sqkFLlSQHw3E6tpD
vh5y/pwf+aJjEV9eeF7LmouJsnTU3z6ytV1u9ZnDJWos3mvqkhEJnHvObQ/iqZz6e4FPftRH4lZH
Y/rVN4jsfFd931IqZ2FxU7ZJnANO4LYxz4sq/pe2q6sQydiBOplRClLVYy0OVnWvE3K14eeLyH8s
lmRG6UEMx3YiSmbhxEE+i4DTfXjsV6RaQU/JDDxun14YrDTrCMUdII1H/oePCKms7YWBwBzrO94e
3/QIXpBMh3mXYfWwNqOL+xY3jA5uqMZgMCCz/CAN2PLC2IUyKu5iPrPHReKg3Leej8STxCoNWsXh
oZdUEXOzloJT55GUA6ycVAJglri7+rfmf5nsKaSwvGgP3PobOQ5B3BfXrDxjgX8tBjTvOmjqdcE4
N+4lK1RqVgLnkCWprXLDhzaHnuJ6/azJATANTUn39MJ+NCfqSfrdVyW/8HZJqCTn4l3fo9meGksy
7XcC/2WwF0vOJsgT4gQ898swn/P4xJ7IXMX3IvYb8ScW9/1gzBDSFFhSghWDiJLkUnUtknzqfRHA
mQUJ/i/Qrbz9kvhHIfdgHT1Ml78N2Vkp5Fyq+biUyRb4arfWnTRv031WwvJj4APBOkgN4Tx/ob9b
ZUPyxF4iue9s1EuK9JrEMBiP5eXwfkqe5ER9D0dHVQxhbyXn4TcA5i7int5rNFyVR6LmwiKeaHap
tfZlmsAUUryRxQ+sLtzaU4mgYpjCJHVRKtNzkLKwaVwNu5tNvt5qoMvr+sbt9Sed063Rp08B4zCi
rIzQLANm/BTdecpd3KO8sH6WS4Pm+cvXJLtHT8fsRLnRBX2ZQua6mFgBzZ4/5kpVVatC6NqR8AX1
yezPdLjI4vvZM4l3KTN9SN/ANuvT/Dxcg5JXoRTEzXy9joVmfUITfG7UVAAASRtlLaN4peinZPEw
zpLpG25QBnnulb4bnAwBVHKn/RUbUIkqBPVk3Iso7oxUSREqi+RDHWrOKv7/lQc+x2EiqrqMiNdS
xpPAboo14WeXPO2GYlLyqpTytr/UduiJrcLv3jiCsszehO+lUXoigcqTKjJshvwuvQNNxT57eRtN
zFcv6fD1eXniFB4q1DactHgaxpY6ctZWbybgsZJ8iUyxOKkG1aPDzyVF0RNE1Vuv18C06V8OTZwg
pWuxpgpDXQIU+pKWaG6ZddZULMalRDU1sMLLEj6h28LRkPOfdSC/0e/KtrT7wRoy2jDgEcLZ1h0S
+1FQuFNQ+K9uL90IHD8cUe5MIK6iR7iN3Ckd5z6zKg6a+a0WTMuYfhxMooptS+3x43Er1yp0OP9N
vaSGwJVFLBXyWa49w0mqj4NXLP/fVmOQd5sqWVSdv1Dzxda+OCI9JEBCucLEOqm3kLXUryMFl3bD
yVQRcosjlWYGZvfJXFMYBI0XTl83q5NNpXd695eC4fN8DhNB7pIU4jaBHGefHletepQ+4SDpaXAT
yLPXthlTIiw5AjFjPKJQc2zrlplIXt3aRhvgbcho4FRLqWx9ORByE80V1J40yyu58/2j/6BRFN1u
+FFaWuMEOhFGj9grhGfHTMfEpz2SprB07rZiP4mrso5ZCc3Dpnh88eet3S7Z3NpNPg3UroC+FfaW
VgQzW5rtiR3D3Z29VW5MaH3xH+WqGWcmNUZjntneKquNV8tMKcc+v2p2asOl9+r9/sjFekQ+Ye2Y
YbBmwuud3yqyKDMjFEdBC4lS+uWTa6N/zO3fo7jw4kOFaszKIimxaisyUEQ8edCmN+n12HbZDCcr
ypW8qbbU3OuAE+UJMTQJjcOzcPrAGtrJUSG+yxvjECHwm6T4tfgpqBCq41wapp+x9TsyKAmgOSvT
PZbZhLFzIy+Wbkif8AIdtI1/tHraABEF25BcOqiMJhi7CIArM4pWREBSdsc+8JQxnUgC9N/oQZCB
iFfj4o8WBbt3meNtqpLpU+wgU8e1hQKQpsfi1G/RyGVbVeCJoi8UDc1Pd+UvYZZrd9X3FwD3V667
uZ7dhmlLn/oDzinEo/Yu4QCYo/MyUB21LkrbtSfxJiqIywIestdfR+SB04KhCLisdtS/lnhqlxm2
2CTltcLi1/WTeSog3iC6F3+uOSsQi7J0ZFCxBlU/M9keOIdQVnqBrLZE2UqFA90zkFD5oPsGwQAh
R0wNhnTuRC+O+rbJZsyduxZLMj7ocYPQCqBqX50IHgdYQrdH0zOodrbyTB7FfQoZxTJeazJ8q6lG
58W3GtxuO5kF7PdkXk9p2Xf8YhanRWMiNiEr7iLOiL41fJE04c5bjYg1JA86dLyVrNx8E26AJYEK
NXe2CScPrYo4LDCfJysetBwvcdqckstZb4DgLvBbYUKoSk+7BQE+G6eQ8qu7LjGF5sYXpZ8z99he
Xfhuodsv/1TYnhO+6AYFck4jxK8K3wTbf5tYXMZ1KjNLzR96vJb8jz0yVR0CHjlz7R5pVXLzP/Wo
kZ1oYWZmpr3/g28pqU/+vAZe88jS7H85QBRs+UbanSUJRG2J6Yb6q80VoPVQmCkH1wkm7Dbb0EWq
Xmbs6lW2XpYTWUlEzFzJOzqeG2XK2FZlxx5OQdXXcmjbITyxKmhloZR+/mLz2rp4MsiLj+Cv9DOH
0Cw/v4ikFhqx6EPDCnvW2qxfR3nvI3MEb/M8rRpGITQTXOBQ9emLQHZKTWmPHxU6pXE7q9iFro3R
xIHEUWcUhX/sA2GiKeOYqIca0aJ0haikv6rd8l5TIVbREVTDOybWE3SKe9eSaXKahbsN42lH+vIh
GSxPmxMIlZSFUZw1NV9B7KquYV+QnbS/0500gYHnT18ofAsly6eHfCRir0+45uWoybd6mCGtCjQU
cjxWJH/xN+S3bl678tmIhAloD6wD2CASeC1sS6Cg/uUn/U0QBb/52pr/veIQpMF8C5cCSi8bp1HZ
xGir32UCthsD2tKONPt3RBsf0qAD24lkLijsbDs5h+cQE8FTOYJ7nh0zyN6OCseOxtwDjRihS/98
ob3QLVXzBvAfIVezaVqwso3jGH4WiLsuxJtnfUr2rgnjV16Wv5EZu70wBaJP4T8NOfaXxJ0Q9NPH
Hyxmmqy0nNlO1Q/QEGKxLqxr3wIg17CWvFHt0m/SsLEHdFyArWNAsTKE/v4Tv0Fha6J14iAilsfo
eVxCqvumofzkaX9cYgCXulwtl4ExfYu/uc/hs9GpU1Ybk9RLlUP8Mohcn5BG1RllV6u6eBOVpd7/
XygwthzchMbBtydkvzwSRV27Oui48UspIl0dWXgXpijxib5RXOhL8FbntRa4oXDQWEXqCoR4+5GK
YOgezY17HLEXmWdEanj+xXm88Bv44Buf2rp+5Ab33aCW935UrFpE2txpQtJc7Sx7jMS9Ks4/gE3p
ke3L7iER3HBT3qiH7azDpyVr5LqdBjfhKCcqsTK6p5ZJc19CxbKkDi8AC8GidB247FlR18g0chyD
X1CVe/VsBXee/5S87xrf82B+XTc86c6sJbtOBCjiRVp/skGg3Mh2U6MBWt6WWusnegte20W3kJJb
DHUOuMQusxSmmXMZ4A1Ast+WQec1Gkp02ucAyQHj8ulq1tsFHmqRTogitIjqjeJgnadS+VtIWGpQ
nJdgqddWkLsQ6aNYx3mHgO9O7eOFfi6otkn3LdhyzxNiY+oYUeITuPfBYbEGejjJm4R7V2J8Qf8d
ygAknhYiNymEvfUtKC4OzSeIBB7UrmiUcYvs8xHYig8aZlNJyc3id3dDAg5qEaLC7ioU5oCjIbzq
z07Y4DjIk8Ytf6orJkU2RTAsgZnB6EEwbNNKyvKe7Fg/yjrjTkrLPZuhI6ciuALVyg3mu067iMO+
meIhI7klbfYqBl3TFW6JA3mmPFZ6XcpT3PkXClKxofAFCWgkaD8uv3RtRkzB4YFm9CawdA9cYnPZ
xj6+TSVSFuzV+MwFgmOtLYRvIBbxFyYHwWsIOa+/5s7+ZeNLsWhqMFx61g6+ZSy+dRcV53KtJ4MH
TxlJjCBAagDB8Csv5F9RCCEeBDh18KC97dwneq5HOqHeBzQRdueascZdiT4y0z4imelCmHHOAAgB
A5PReYabNQckvmd6Iwt+zH4ZZ7oQNVNOhJipet6rnaEmFHH4kL58ShtWFHbepN0thnSx/Co9Awb9
ImNkgbjzCO5/b5IoN7YYRiax7GBKmneDbs96dDkJkkF9h+nDXMroCWtx2PKpxY7iP91AIfEQwMd1
zb2/1OttGbXsrdGjpNeonFKVDG+2jQ1Qqm4sY7iJfqIhVJtrKaVGEVUwegd0bg3ObdUImOfRY4yF
U7JhOZnTxsqpFvxfYhMdM6mOieAudu6GVlkspBSajsR8ikvLYJlVLkExOVJhKWOcNww5qJxvSzuG
aInXXgfWFQyhZH174zon9I7qMizJJvqBLRaItknji2QkJ6DZ8rCIQB+qQ1RsUd1eaoaOOkhQW8oK
l/WF9jk2MT3s1ghW5SRKwsu4mgcJwRBr5YzBh1b7Lk1Mvm2FXo8K/1wT9HXjKN0NphxzUpd5XiGl
ealgaPHA1UnNEGrfERbK7PH/kgZBTFIErNTBqhZN0AY/f0F2ytuv3aEaBcXHmLGriXpProvhFLhS
/Dm/zbV6TycEydb29rP6iSaCsj2AtbSOsmzQcIy/sn4WJ8TZ/TPTXL/gWUGctHIpaA7x/EYgxhDw
K9lIt88GuqBmjeJTiW10SJ0zO3rYLFM95G2fjO/HjpTqNcZT8VyGEPvFQ/t7fT+xlSUzVEo6j0Su
C/Vjw5Yzy7+rKX5bwZJRff/2ejVhLFn4PqhwKUPtaJDrq3cTiGm0i6SE6544EyMx1eG+U0FVuafc
pDh/KZQRh8j7stiKsiNOFTcDY1AkMXl00RJDSLFjuE2lAGRubXvrX3kbOdUbS/lWHcmTX7XqwDEf
Wz1Jw+zgMDpi7uCHxl5JEbJM3Tkagrn/qksxoE0xVGLa6wQAJt08qZ9ASi1fbwpXsXB0tJUjTVXJ
7LqMVA1+vS0315WRjYPLANuwH1YPHL+ut6hJxwlg9GIIxestYTBrgNy6BEFMYkq7F+lv/pLHXCCu
g0+6JMFOuIDUG1CdYvA6Q1IUNhwZLgCPwOnlWasemfDRwGD9Zq1JpbNuRDNRLNVViRrRmh6o/q6W
j2y1uPj3s+GKmNkmQVd1cXGcpZigBsRSSNh4Z6WZ6iEIeP+kyCJOzFQfKcmO0YLJzZcoqUxQoBsm
/zrrrgR0HmLOetqvIUXS+CAcCGP4kRb1Gu5s+QlUjURcFme19phRciQKFkQ9zSvZWU/CJ60kSapT
Z1IfJzaknd0CCwXelLrUHwv35SrluVO8YbXsjbK+CI1Swx3A9QGKA6JQWrDUuSOJgiMwjffSLkf7
Wy/zQRE+SAaj5b50QKv+rVdGYvLRYxOMhy2T/ZvqrSRgH62mwTe21UtWvW6MkmIc6K9m6/DZAGCt
2WSBSLi9K7Le3DlCToZFlHwCY/UT4egSgnyZBW608PO2jWmA6rJvnrsWOJduWgM+RjqxlxYll3NW
RsYAh6i0MTXI7y1TXcLLjL+4DAK2+Ap7DjRXAxHM4fWvihjrQMSZu7ZloyuNMUPD9WvZ7R2Rew4p
tQXMUv1IWH8oh/EVz7FPWS/LxLb1G+NHCcIuEULy1oK96lILs3jdTG0eagtRFghRy6QgCvLTe/EA
H0F4w4NBgOBzOHyrh6Um1rO65828HK3ZBl5Z3jNJOq/ojjugLpVS5RBOLTkaAuNev7CdXN6aUaZu
oRJzXRGYrT1uxffKjEdaIx96MAr+lYnK4WEL2S7GoUV2g46AtObsxhTK9XYdEx3B+NrA50VYcisM
Yiu2nHJa7WtNB2qCVpwPxAObcc+D5Czoo6vFqYH5heQsxCWXzMr1AatnsZKArRuBopU+H6yw3uPU
w6vsZVn7h+lgzIQf5VT67pQbU1ZYGSCtE2f+KHrH0U0aD5V6Jdm1/sl1oZKy7HvDNVr2641ExOuw
Iyr879qi0e7J721n9Sel/aXbcAIafEPyshPtOEh+miRy55O7+Km854I1kyCwB7uYSQBDcADsFfwX
EfNr7L3aT6eoVkl8v98kfYRlcWcf7c8h15e7i6jQxw9OPv0E/6A6XA9DU/QgOr00Srtmh5Urre9c
t4kWklBcK9p8C7wp4x0uY/r81UcuoRcbB2/jJURneKQNtw4tLWdOdb2lU8IW470/GQUgLwRFXwzS
u+meGYiX2p+fiI1q3Z8QtXRrBGPds836jtq64PKp8kxSxXT26Kf3h50MXmolJ47LVTUKEc4/rfHf
A/ndpUS6DIzr6pq/E0XHDzqzEbTIFQNDThWDmi4aXezdfNLwNJwDDZrC2WqYV0J2xvpml7LL4/Ff
C9vYV5ntltAl1clphQ+yuJEmcnL/lhPV5BQPaL4fYrYKZYIqPfa2Wnlnb3YYBY03vta8Q1HS01RY
awXCQq21fsye10VcFBhiQArcyCmdVpTWu5pq1UZPjdazpfB1kGsZUl9xYxpHq+M7GKP3jaQs/TI5
XkBjzb6SNlP37chxTRESDnuHwqB5v6L1w0h5DV12A3yOQ3yYNnueUUElyp90ZXRy/PoNSCYpFNS9
BTsiXLeikg+FqryRM0oTVAFAmY2zvQGCZQ46CIRIOa5gOYTLwl7XfnCRapC+BKFYVdcxEld7CpmR
lIkgyKezTI0FZNL8FJumX4VqXufYuc6ZTeFwxVQ3tpQusqP3tjlCUoPwTLECEu2zwA7HC+Y6YF/b
Qa4kMSq2gEJLDkDJNEkP2CWwfF1hG9ujf+GLnEkaXijG2arRpubZz4sBE7bGwC9vQrGn1StgfbUg
/Y02yBdcJgWtXksS7hMVtZ2h4NYvTJVaMSjgNj1nYkrwtR5Z/Sz0tAR7rThMqo7BaENOL0MfjCXp
Hbu3cKhWAinEAbwdGTp2/1nRQQ6Y3ZyvASbl7M6T7kKhapAUg6hqVl6omBKLRbB2y7+yD5fzqtr0
TkdIBFGZsbJThboJEhAoXxUi0jG4OENyd2JjEcR5uNK90POyg9i8X1/BVOt1IQrr1sXkAocgVmph
QKHClgCN2C8mooinkb2HgB4gim4LGEEdfzQb6PUFOhSOOtELlh4n4YqCPjLs/K4PhK0Vvf/IJUzL
hYxXwvVou0MGUrKtZbNoNWyF0bfq3G4iLZjx5ykl28Q1jI+j9CT5I2uUIZBqUI87BQFJw9MLchQc
ITNEHagKAXncYrZOGTfm2YfEbdRAid8y9OSXSPnD+7A5Hw+N+H3+6CI23hmSbsYBanBopbjzwzWx
eKyw2vsJNgVI4CmBFx6ZwFDKvKCsP1tcey/ubeCn4J4qacDKAjAD0qtoFL/mvpdlDPHvE9kl2uuu
WY8TZZK9nxxtpfx/Bpb3v0ODnkZZA4/7XjL4H2g3DPROJxaWtyvN3+Y5Armwqj8Da4Ae4bAFtDx1
S7yKZnD6FN9O2V3Nw08TsVhd0khVkTtgplVscTKIJ83iE8p+vA3PhoeEmOOBq6Muq68pNUeQTdKQ
NvwQE/pmHNylmdZ9+Yjez6xkJu2unyN7u8jSPzPcUioR9qFBRiMbBGCfA6GP0QSkUs79FyEvzbjJ
RSopAWHSZi8qzYmtZBZTFam+hWDns9W/Ogax8yNVYe480D1vAqIB35Dt6FS56sv+nJhpVQ/0FzHr
oHZQUm1dxhV5KeUbbDRiMbF53qRCgifivgKU93624Tuv5ZRduoDgvsa6orAapeLvE7tq2bbJvosz
uEs3nS8pGjMfusMI4ApUX4MDXYW5jCV4JqAw73M7PkzGPgPiCiOFGUHAkgm7wGyQqjisGktxewjE
1IVTF0/tJfwNXKig7qvT6YHsqTWO4P3tzafHnq15FUcuyGko7roKFr7WYqPgyLZKI+bxaAhI4LK8
+lASWGQPOWRBA3cZRrZ5rv5M9MChsA54xFYTGKJbZnhDsDqu+/uiDj5cNWR4DTw+IriHj0mr0iYs
DQmCxA2a2dtwXTj2UZdk4fpuiZvTDPjV1Q1abbGD0ZSBa8fpnmmI8KP1ZaNrdsyTjSsGuZvF52Yu
rCIeu3DuJl2conRxMsx/THHlURyeE0Mp7DNbK4lYnYcfeTpM6K9XfwJzmtxv/ZvcLl7b5JplVVJ1
fddNoDopdi7Q8p86SsHvQBMFc4cJ2PZGTEQF5nBgJ9D8R2v1C7Gnk39ZuRbX+/ZbkTV97s/B62cx
LO4cVZLk2BLUs1IILdtBkWY31rhaJ+PwdYB5vVeEpXSWIFFxG7yfu6EIRn9Vr5KAiMPJd+8UocjY
SDRPVgirubf9Qcqa5r9Ab1Uf2QOO4xUA39GiMDBNAEVJEdBlKqmcy4aFxCEB9fY5v0EdZ2Ak7x0O
SQbWB79IRkD1/Wt7bpEOgSemFvw49aBVisVZoA7Z+lslRzz3za7dRx9zRGvw0NS9ocduWbhUa1s9
nQtXa44p5q7onP6VWHxHm19bYx676GjiExgEzGF5BL9FDdrUx8k5gpglvFKghTFfbrl1AzIt2ak1
jPxIf2KrigdcbXLGEFHstfFK81/NjJzAYgtpWKZvPZ6667DGq5YBJyZu2QnLNoHNewELnKWNcWxS
k/c/9AVe+wU95fPswAGKEmsNp0NUFd+OnrPacYUydPkRBlJeV5+T93SlmtIyqG8fgY4Kmalud47b
ys/gwvjIHxKo+CWH8tQ2D8sArHzEp6EqLAhQbYIxq/C6MlKnrJo1VABl6LsSeMxUEGa9mm/N3WfV
M0IqVRzrcbfMi0XK0U2nQv1WX2OUi4vub5W2EFeh0kRU0UNV8XqpgNPs6fHrVcP4pV+RhtrxlS/I
d9ALCq+hd5SYRRAl6/Ls04PKASHZSXd/9xPSVOxOSlDFf+k7b2Kuc3rl25SbKancrD98nNeO9UqH
SLSZs1h3V9DntqgIGfXwfDdxapdPIWVPh2ixZ2BuCIMa1vEHgGR+c5LP5SWUjpY/DUostp+DosAb
kcw3+EkEhOgkbIbSwrzE6tmdm3NSknKk4czLGz3yZwskLbt+MbgbePjqwI9nLB1sk24sk2DAzJZw
aKUXh3LBv5Z01CiiSNCTNXQbpmYNiqaqbPs5MiGCS0QMyfoHv9EjdyutxPiaSr+zBsnRqBE4fxWR
+YXN8Ulrs1rLk1D//Fa+uIr/qnh15PTFE9DmL48ClSG0U69WxMcwRT5sU5dkGH3R9wdzufwSdVt7
eop0iOk835n9kZPQF/dNrdW08ztpV6/N1up8whKdXuf/3CT+iYrMY4utTkgE78s0lOC/SCsjN38n
G8ZlEk0I/R40uLT8VbJ2NZuR7HijIolWq/WogkSE37Ia2bhsk7UMhfY6xXpaPHRhvAvnEk1chI6b
g6Y6VHDBcrVjdo4CA8u1VIhzlIe/k3YX7KfVEFJ2IEpfb48dsLurv/58Up5jjMHpEgBcMan29lN3
1AIwVkuM49w97qrVimubP4TNRWYWqVDytBRWUqoGFXA2+WIhqYF0StscJmMrBpRdDrbSti2k9HQP
qSxDAttMbO1HKTZ/GJp9TDgdrp66m8pHYbOI+3Lp4aeE4dN6bOyB3wRkuVRCQKZKh7WkVGiqP0AV
1PdF21oyv1jT27Hmq7svzPwnXgtmfqyccG7otWvqR3RtD2feuG9+/xjCfmdb7yGyS/odMzv+gjxy
Dbtfw0ROgjeaM78P6tkN5Dmo0r0ayOE0aiCleT1cmXmvY4P6b7pdXNroTa7HcdtFC+HfawaO6d2F
IB6w93h7h41CuoSC2P8Tn1oBzjKlzw1SL1kNyhnG/UZ3WkmlZfUU0krEHSY4o5sTcVm5VHALM4i4
m8IirfWwIWoeK5i/8WBQSHAU7n3USt13QBExKoBKKMFmUqy3B7u74hVK24bUHD7H8cTCtJkS3DpE
JqufLvE5gMXJqQut5DvIc/CkfvfRczoIyPdx/0VCcg+qdRW+uIpqj5yUEdYxITRowIihoR4b0+yG
IE0MZ76CJ84/+sbnRG0wcq5REIgmUrn7yVe9u74Eh+36gsuoDKT82W89TIISw8bTiPr6DPYhpSq6
lq47RLw3bykFerUgG6aBoU7Vn7tyy9oTEAMHWnhgvE2+eITJO3paAe7x+ITjPYjWUTADwcMiDtmO
GCBfvmcGsKXsGOt9RY1br9pBZVYR1a+AwAdAPs1CcepXHgiwCxVkfi67VcECqfDB9k7kz6sjcYQi
Xe0nOlR14IgGsXU10q4wPrXI+3whe51Tsy6cp60i7p2PIOwwXx57Z665n4Ph0fJz9/TN6KuubdTs
uySbvg5FLGmuAiEz05PXdqgkCNACjQDUtdOYja5yCvqobfHRuuU7r7Qxpkp5Kdet7dmY9QVDE2mn
36qtLbHpoDbflTnOqJ9kM+AiaK8zHSIN9rwVuLkuv74aFELDyjAO3yYg34g2Kl6ql7Ejf6YxxCD4
3It508c17iy9UhX0UiOgtAr4e5JqD6uoenwQA75Jc9mvcoq7zfNO243jtg3PMR2va6PpzxlhMdgH
EUOsTnkeXpKSZydjnszywk8RrsowYFGaADsumiJPyc8CXLOvecjVE2pcvgPWbyUSl2ztqxhYIXf7
d3VWstdl96aAljQIeGT22RjIZD3rjF0SuAAq7Nf1ACpg+jVvHcQ6YYL29InaHbScFxCrP3R845R6
h0z+XenTUBJZuiKomWxSVkbztA8dT7eqJ99Ut9RkLz8ibKsRL07RZ+tNo7v7d81A61FIHrKc330g
g7WCecaHbH2LOzWHO3ygNuILB0uk6VGoPIlKOV6jaHL8/zbIjRe6k4oH4RibwKH8OD0OuoSKGVMi
Ll3dBkOU1FtEA9v5OyJsRgHbVVb3GTbRpgadZUqS6hxdBuibArampXph8vLXsS2YPULz+YNxfDWw
0GjcHW/eHsLiemxMKEoJk9iKauTGZ7VABQpr8JOo+w9bVDJzDQepxm8JGyT3zcV0/sC3cqw5wnqW
Thm3Qf63UX1QQbCV7NIDKp8+f83lLogxetT5IIW2syY0DwGygq/hoRR8WPScHW5gN9V/NKYf+t22
Pkf8eo+2xYgEWZJoUwYKbyR2oTTwRQZ0KDpJlDuyVK6Mhe2vcVcPwy/MKrQxwoKtGQqpwyuYU1kP
cTvWjBF7xS0SaW5Vbvh0iojhx5VXx00na+n55lPCMY5befdL+7R8Y2le2w6tGUeCja75JeSThIV4
BmNDHQcJgZaDYHOa5myyj4qvkukH/rDvTPQtwNKhXrL0rsNTEZSfpwqv/kY/1bIC7H2NuUZrJaxj
1PMkCVMQRoJKSbBHJDO2IjSUTTpCP5pgsR/gA44mOFZJMnfaUfhlsKy9vwUC75feaTyFn2Rgq9fj
gJhjKjAufTwU2ikKVpnV4tSQIqgom5NEWVt7goekzh4EdIGmbiCuzk/MTgXB0KC4msU8KobHfwYf
4nA/QZb/KiDb57YIr91umgnLQSqHAKxO3xbaRIU5GHWvvBGmrAbLhsck80Uor2tGMgXu4HBwprgY
L4i9y1Cj/y8hnbKxaaQ3OkNTs4IXEtl68i0WiuEv6ttzfb7jWlcW1w1P4VTZp7f3MimWFY05HMe/
p5XJh0fmL1sX5Ez9xLUifZJIb638QoEfX7mWf9PIqCuEbq82qZHIbJe/DQ3bWiqZV3IgolL/nI71
bqHC4AIXE4883icLw0snCTP9dVXRukTOFkVT+r9Cf+TAvMmemQHFPH830nf4fSvRJjN44g+rQEFr
Hxf+XTFRlKixZ+SFxus3f5bLb5KUNv6RBewVrt+rXJw3BjFKh13PK4AU537P3DjN9tFTAfMwQ7jX
vGKiyC+yR0TUO+Fq/rOmnUZTrOSaCmPdxNkwmZqRiZvwmRKAR4mDv7xLBVuPfqcz59oPWeXx4tsW
9HQFYF1bkyIpZngOJpgtNEkkEFjChhDjvevXePF5rxBxWzFZ8orPai8XDvaQv59iKquS3kb/ViPn
dRs1S72CtqVWIX90BAKy/OdD7dEAiOUlSCxmCAfDozvzxp4ojjVVNWyCrGn/3aEgHa9aCQp9Ntt+
3rumqBtwLA5oBuyMjBkY9+g1z6rwcopLG2rqj5hpCcMxLULUC5zoexB3GkDju39xhx31JeQB5/Ox
jcsk2vDjq4Uo9E/nBKW5FguTrP+vYBoXRbwMDEcg2rfmSBq3aQVX1mAvsR9DYiFEXRaQuvG4opCp
5EuNVrpCiMYLAFFjR539ZtcK7F5N7G46euXmRvGQTid1YXT23dsWFShIAPRZOLBPzL6lVqZZ5MGh
67DB6Rpe8LA6PZgEbzL4MUb9kDYiJ5P9FFww5ZgMxWAS5GrqeIQ2+IjwQE5Lp4UclJ8H2RLOb/oj
4AySUgiFzXeEO+T2Q8pQRnQxF/DAs+lW9m5flMzePS4elbGLOQcPzaGO912DT6+OQStEDdP4Oeyk
YoaufhLzheewgI7gUEhksYLnHiHA6orSjNMlS94I5OtK62keGTqkem0sey4/s66oJYAjoWfYAfEp
gjqq0LINuQ+zPFAPvCK2lra8ESIMJCp2umBEosx8/6jMhB7H06jA7+eXpR8Y9iB6DOpk8WYr2Gow
CtB2j79g87GlE1l5FtsJiZ9MPZdayL9tV6pTuFIY0Mw2RGsE/yozkUB/k0HF6MML8AVpl1J8WoIK
w5QHCruG6qGurpQ6ZNT+DazMyKfmhKl5tKKdIp80xJwFIpXu059gXQxGtdNEvJoKPK9ghg+092OA
BOVuq9kiCcw+SF+kLkBVSqp6ANk0Kc1oX5IGYUh/VaX8tSnoHRdJ1IaVgeR4o9Yyq8weOMyGaPqr
GsggGondu+SpnE8lIue4F4UtfpGhgzaRK1ezND5XstswZmpN8KkSJuHmeNvCzGH5j8F04Mb6abER
8g1SkNmhwkxfcE/IzgoK1ewKPECGGwkf9cgQ6zTC6hAIr6ojeihMtf2UBgv32Q+lsFbiG0vBfyQ/
K+S7CbOC+NdOpG1HQzyzvY/MFHbIt18XN/nw4NWvCimEn4LmnVgogslAN0QT8Lvie/tu2f9XGkOo
aIz10UqsokEteWo7tw3vkaqD48kE4E1oM4gfPoeeo7Woa2VWRTn1+1/5JXlSi6B7BzU9PaurXxOR
H800aWhY7kCsz7ZU4asX3oBz6sXBVfDd9hEUOmXEv8uih0ltLS1wbLRKNrH99Di322yK5ZjWhP85
+Wc0avnRP45qoX1TPU3icoRkWWWnevSjrr1hfEBQOaojpitupTg3uhRsRSG9BABH+S+6X3Fo+ABG
TwECtPyuJjjQrbfPH3XMyCNxY0uJPNf2Od3SNiJRFyRXmFKIpLDPDAQZ03GKedjGOmt2NWi0PUWr
urBoUV4j2ySZOzLqpxu9smuig1nXbsfZBrCn1yYMoDbkxRkvMi2GG6kJN8vLn9cwjYD7IFAgSUOM
l/wPeTvTEIeS95IutovGEQhFCBnYoXg8MpZi72XVBdPqyyJ6K3KaVrNL7gAto2Byfw3Uc8YvNZMp
JIU5zLzZUYhPbGGBNxDSR6fQKmgHpYo14yMDFqWFzLyh/4WIBJ33h2KFxh1g/zOdWVl7sCNwOY72
u3MIZehhQU8/krNtGWv1cxXgQmYDWdveHvLh7D/h3zyOlWtpQTvbxcVtz2sVV8V2bIhxGmN5zf6C
TRpQ6HcgmRxNAEL8Fgz9idNVijmlcgu18IppyS9zpnvxUQvUSuKjWi1xSfRy/BXVRun05QW7IRSV
uPL97Y1Wy1SasXWtVj99F9v1ve0DD09Mx+opHKVLLhxmfit1yZiTnZEDJLnoQtwfL3RPEWgEJn5W
0vM4+4Y1WX286nyE59Z6L0GKqr4KrUZHz/ReD+HNQWC0xML3I3mBh31fu+vjn/JXsNryZ6rX9fOS
Rno6U0vfOKCjBlvUTcdnonkABxjytP6I4HDGFvq6pagkFV91v8BTD3QU9GVdBvWBGLfruakYpm4g
H8o+JArJAUKXYX/XuT+1GiLomJ//dc3bv4pOr/qrNLmQZijvATbgAv/QDBrTuesBu2Ii+LMu2mke
K+98HouwGPfbTtRthRnfWR+oC+EkyQ2Vm5CJb0riPZOy7Ewmllc3f+A6DLpYtidA4yz9zTdBdUXs
eZp6ZfLYnlJ9SVWxKbndd7ZFVXOyDwgUH7HIqakpNvLN6E8qbwF6WQZ3wka0oqBKW9+3Ex3Hk0ph
Jz2NtCLxL3Cv5mnXgHgSaeDFJ0ZTMm2pQ+QFwlSjNnRA/v3DXwWzES3dGzxhPOv8FBNM7knH4rIg
3odDvbCK0NmNzPmmvlrT2TFyy/5Gds31en+ysl5+vmLaf1GKrUU4q1rTvH1+hQxeUptu4SnvPj9w
ACkZf/8ha4i69Vb2XyDa6pEtKm3eou9xijcOiKlEXytKbVQRvcDEoW7QDiuMZErGuGZ/WIwKkd3Q
mbH3Ey/7BZ6LCvS/VGzmmeUdjpe157hVDwEgb9cTMyHsOsmBztpBUPueJ7P4fdHbi/yWHfGDHJSJ
0gC99wOjXNQWtfHC4Iuq3LvtWPpvjxVIBpAeMMduRRi6pU6ZRFyvECj1gG/ctw33C9bXKY9tcTBV
5KUuDgA799sPgleZMQGIc1IsP/o435oto2KxZ2V8w1DuZayUWtPOLwM92d3Zn5Xev46AYppQaIjI
M6dsnkh9paNhEvuYv7M9d2OCVFQzKS+l1pM+wgXRGIqd0D3M3MaIdOYW7vx0UinRhNsh3WdtPsMA
Z7O/EbgEnBWvxxFXGIrCTaBgBesAbNi4OWX/ZDfV8pUI8uqOxnzSlet2JRaUY2RGaEfSVV9oB1Lv
wYKUWIlCBih4ujxpGa/jNmmmB7VzJA23Ahzl8hWMiqIGcXuf1n4kJBml+OE/kU2jahqnZX3rcvu8
oUuQ0NRqyMdG44d2JVD3op0xd98A9uSOpwzsMgHCS+bDWZ2kLyAkG3wNGyb+qZyIR9ciMIfxOL/v
9aeCxbqrkbqjPxCT9GD2Db3TuN4Tu7I9WyI99oqtSLh2PMXDJpL6je/E0AoKqVH/VtTH3p0CXSBY
oeyoZU5BC5roiey1GVlOZVmn6GPLY7nDlraypVkG1y2kc7t4tUiSjRW7sC+DPxhds/dH6Kny5J5T
V4BFIh+1MQarij0Np7MlJDWaCn58PsPzHjUDKH61prAfJfs06Nx+K6sL150IhQaFm4l4ahjnwvfw
koGuO5C9y1kDgmcJNedc95rBG/sp4X4P//ltJsi45aKMp1GMbM05UbAuVaoFunubzOB3b8xe9H/7
twPUFSs3JmB5cTktgjpbLoKrKD3pMQlMcgVtuIdWMFgF9cpDlE7kiQHWNyPAJU3yi7B3Rdbj7gyE
mQrXKTbT+d6pRKwqpxEdGpQNxSXj0HDLxUQ9goXzuM6Ih9LzoTR1g0Gua+opWxL6sj9IKbpopv/I
zrm3W3bFnJ0BO2yW7b/NLvNgUznWfez1MezhGlWqeBDFM8vBAXsjBNy0n0M7APhQewJBJ24Pa7jI
BxYP/Mlj/crlVNHbB9I85IarzyL0XAf64XdeYuPpB+es7djVqt7U0/3WFJmE3N/NOBLifzx7NOFc
pGNjmfF5hqD7m4vK+w2I0ujBZG9X3/XPwkR4/aasJnpQBmC4HAOoVq/CTvOrvkseJbCtUW67SFw1
6Og1Tw96LxzX5ECUwTlc6HPXZT1bnCV/brPUolkTnsaTqv7f6GJNorYV6v2TFif9GDah7w/BraIk
UD2aEw+25pE5Uisrrzk/6LqrG5XT29RvcI20j248gnd6OxAfvlx1jlEAwdDUIaxvAOCsrtTmrofP
xCxopAF8oWtXUpISBfmRoNih3HD3gw/T2dzoZbfZ3mFVSmlQ/oYeqEEFM1rmqNYN0p3HIejXUdfC
/23nOdb9OdLp8WU2A4e2tth2HOXbohJCIZQuAtTM+pDtxjKqh2no9Ilo3fd4pjT25M6HIZPMcJaZ
kRbA8OVKBwzbHcz0OACsP7SwXFgYVROS1fhW5yCTubxi1X9UnhbILXgdt9s7BpGK3yYGyUsjJo/Z
LPOsdumCyEnSrnTqSlxd9H6/wqmpK+3tvP9+7bFdCNfNW7Hg0UsnjAjHlFw6BixR76HGET8R5jYG
x9lJlwi/lynMlylZrcJCxX365zKVWv/LDwcRBiGcvRfGXW6lxCRkbxOmbFUmVawMytXQ5Zm4jE2l
OC489J/tDAF0fkVW3wfNMPugawWOzMgk/cOiB1rYfrti9kSHvOQjdfNSndH8G4Uce57qemoKvwiY
J4iGmGdetCFPCYDcC6nasOCfSRNtw44o4tVvNj87LTmnZ/qh4H7WFRIqARArXoZXho/6qxo+fOwB
4E/kUWDi2A40FoZbxBqv7WTyA2C/4u7GVGLlxK6AgFVNaDck+kVxBNESjW13WRZzi25+tDe4cAmg
Vkpf1IWNmWVeeSXRnEEOU4dRGWV1v0epVbQDLjN4h1qKdcY1n5SwMl1yFwnd3K3PNZCYjHE4ebyA
/6ggQrkr3H5CIo7IRS3O16o2p8kqfn6uEhDbyG3YNtVUZu5GorQ/ye/UFgZNh1A3MqGMFpYZ/UuL
8L3XitK1jaAMZciOtkkUZQdsQ1FxobWJnS3xUZY5IxzkkzkRCOgy6fFbsHxepQaxw302YfJtxADB
hhAyOJ/7+v43MHesym8QeARHaOqe0v85g5Zr/s3m/fUGdEr/RgffFtW9wB9HAMagurZ5+ygYe3Ej
KGlExA7lV4+oJEFHIRbBfbQzhW5Hd0OKd9S1uyOMJCywz/C3Qh0IMuGYWTzAyWFfSu/7WBiaE8xo
gzFF5lWHi9XogMO9Tyzgp03KWoFdqrE5/4oed/ZzlzRbrKZIuLyUAwtSTRzTmq8dTAWSyXcrlaNG
hOeuBzZdgKOQ+DVLXpLJiGGgihSqf7b7jjVn03jSa+tXHnz+8YRKUCqRy9ZrHq6kuAd5Z5Kp73J0
yNU732ajjIOT/x+E0lL9C4r9Ov65ZnWuZtw8/mSHWgLAE9aqc4zmjHYHsR9oIDzoROnyK5DCVLY7
NnHBt9vS+ok2OJ5LJeqyJuu3HLdEo+npp3tPTcmfa1pWx4B1MlZQ9ZhZ05WNOc/zBUeVs4mEZl98
ElOiKkQM3bLIhM4HPHa6ss3eJfX5JfKEMDFqPXb29bmH2COjF7snxgaZ1vajZQTZPgiug7LLEtTr
VQZldbWDgJIOOl6dv8Up2eJE1j3VPaDg3opLQHKF/hTOmfxKWCd+FOBvD/ba73cP54vubFNGpWAT
4gm0tkaEFi+efmyj5+owyHxAx5OmaVdqB7oym0QyQFCfumOjORE1GhvphWbHcHcZ1GZV4ckfnDCv
YWQo0FkO32bp9Nx44pPyru1Vrt7y+HsptHO/Aq9zaUnsz4wsxkGFLzuaPgqUzhXMUUHufATYa0X6
1ieiUG+svDmBYHCt6YGCV1JKz3HOydMWsgVkmEcQPRdRJM6gUDL5Wm4P0qQEsCqrepqQ+a0pUAUI
BaPMhb97vWmpJH6OkjGCRUYgbjrMrH+WH4S8v80MPW76F9ibQrInLfB9EFuwOm55kYIhcxHI77Ca
zkZuUeAxmMhP1wp13EJ81l6sMZxuxC8HPtMPccSSxId4asi/OeF08NGc2mnq2tISm++Na34fgSjP
CcBJ+UKZorK72ptVb7mcVWy9p85Wqv5MS2afOquu/gOgzeSIUTCgvE7ZWWbwcX2X5clMNI+zkd7Z
w2G4Yq6CB+Qhlw3abFz6BJEJASonTqLauQ3mShlBIkyZpaDec/qKCNVt39E2pQGNgJyi316kUIwu
vVFaS0zP40YZw8t4DCEL5GMBJykJEhmSHVMzpH5VUTXX9l9K52UeZlp4V4V7X99m8IvY/0wX+nAD
ejOMVvE+d7+HkpMZRJxs6yFvheNq2kxyadVj1CTdDlBJlXxV7h01xX6XRb6GpmXuYVqM4BZ2XplD
xAP0bZGkP8LzrOMWcKtoIlyfawdQUqYojwwoV4rIWGW8n6LH2klDMy438et2ThvdYeO61HMc3W2a
dbgMD0xT1DCcddzgECsBBy9KrhKoniuw10+4OSNJISz0IMAX8ep9eQ+CphmI0fvtIRv1WmyDzBof
n5WXfmxN7vNu2PVcOsFOxuP3jYC0t53ffh2H6OzUVlC7o2YCHxfuIhJ1k19t7QPh3q6INz2CNSho
RIcdD54TNP9pRHvMsvPVTf0WMkl/9u4wWmf49RB8QWmxazFEikM1L/KBNNcz7WHrdxhcSTF8/vjf
AdwIwd3Fk5tXKwGCCYVJJNmpj3ikT88kFQTdDsuzmtw4uXx1Yby/yWXZCQ2GgCSO95U9YPVibMTM
wnsVWVdRXQODgoUqzdxe8ePqU4+dwiWVxv0C9qBW5ZbRln+P7DJVByvGMCc7qS6/WQ++BzykzdsH
jm31QV9nlrKWrIkLNEU2+zW+sWPQ+/+mNYoDnqjZElDsPA02liEbwFhj66yZ60JWoMUDRyWyAtzu
CbWppk1ejn8pkns4UNTKzAvCJcpwYMnCmw0QD05h25I7zoO1Z1v9Spw1VNX/2+otCxtIVoyCCJRp
so67Ss9XnAtUT+1qAGcWVF8TF4AvN6ugJQbJumvvxaoiG6LXZXJk1FZQKwPi5BOlBjiCCvWzC044
nrJsccWsS+awtxH58WJ8Bo7LGMY/D2y9zlw1wkKw5fgJsqreIY7/fjqFbsMVXj7Bm7A17C2Wm4ew
1FQ2zOG3TDwLh0+4dA7oSRmAEY3wHEGSBMWTovKatXO6bo7tNVKD7z8cLMOsqSIT/uKwvcZhLsua
sJcDkCjKURirZwHBv8spUsSE2Lq7e/b/L4RnCJHJMULF7jX+fLvkUKnr8XILszxLaP1lHLYqEb7V
7f82dlswU82VQbNIi4WmRXS2m/8Ck3dPAkRDICgzMHHHoiwDhzLFW1ERef/0F9z0ACbEcx1A5v5N
ejey94zsLOI/xOY0BSkISsDaGs3vjH8PLEF/uncNoAEqTz2+nkZi7pt42kikBY3R7ny9YMpFrdBz
T8m+lh65DuL81oPm6smJgLcgWRRKfuTtu51Grxs32nlM27go972463lg4mrqSKnZWN+4mEo6Ff93
MLOHJH6c9ERhq+PBFdQsDyqAbt2t0d22VC98be7q5releiXwH6xpM9/sfvDHaZ7X56JfVJcKvr8y
zJc6eQWIjkUrI71J0RMeKUVyTpu3B4VvEWEMzygU7dElT8JuetWMcKq4GNetZu/YWH9hPq9M+ReI
3b1gbkHH0AhnQ+wFXMFoPCjGmLJ/iYf7/wdhIpCgDgjgveXB4FM8dqA0dpNU1tTmhHIYuke8pysI
suroZXiQCtiZnP44UjWpZqJDksDtaE/40d6v0IINPzaUqlmz+0gnDPe1Ejwr5/aUEH+y7iloFXZh
8/nXFsODB5NttzqWDfMR4fZLZZWVeX7MGkp40UhAK66EsJZTfnKhB4QyJZ+G/hJ/JiCJjPtsvzrR
2+4Bc3+Csg6c5aPfP9gAHm2ZZr9JyyGJt+0UIUUzOOIpffrSsEoihBCeMFB+ytwOnopzXUURnK2y
jw1XQg/6eAMFkVUAlwn58x5a4dNrjivVvs6QEbMajYVRLKhuKTpgvOS6zBhwO9+BMvAaST8N0LaJ
a44AArxFUytLZE1UJtU3YaTID5boSbj4beCePwDSWs+r2aWeWEWHIRq2qNh8U7sKLptQAtEi/pEt
k+OuDCFw991vGB+QUugc48ueRmJRRAXMP2daTj3GGfVaUN7QindOOV1qYvTwjOh9Q8jbp/3AySOe
dETFfjkKoGE07c4wUL9PPuKVIOdEGw2zkhExD1XNoXB8qu4muI4ZwUcH6Jueb/37IQd0CwTDT3vD
O2ODKt7dao56BKULjjQaBOFjP5/LG47WT3ECEcXMwD6bgN1ekIfNRoTV765T5HUZW8LuLMd5aQAo
1h1/aJxfVSSHpuDSMA2n89nGmSb5HtDwIy9Vs24gHG39aLE1nsYVUQZP9dqq0SrrsyFp7kqY/eSc
mi8Qfe6tktf1QzOM4we15XjPke1/xy1TathsX/8zS4Hv6ZaK2DHBn/AvIBKjJHY2JEs+FYqK63Ba
b9DIwYhNjBsBXwAH45xCU4Y++ErD0jzIS4qYkJ375lsD2Z/lv3HoQwmwZwJBT++iWomMNzUrs5XB
pIRDR3q/gcJqMvVmJ7FdhCF+wynjadEXVyLd5kZiJbNMUySAxoG5Hr1c63tea2m2/7Zf9d5zA6Ml
p1cWg9uu3NX3JDQqPCExfApmHNArGkxI3/TcK2RmSj6O0NMIMDp/frVANfW4FGLNd15X7JlARSRx
IiolVCvwlqkVKF9Ji0H/N7bUqQHBhlyeVsanWpvAjs7Rc1ulWZNwccKhXiybNPysTIqPbNkzK4HY
am3l/gLVru4tB0GkvpnNShVD5LfW86VFU8wnrXhpNGdwv850vWZlguK6eG8vw+skBH921sCUuGSd
1wZlBO0YLavnYS/t01reOzU41z1te2zV7Qu/RZKutUfCnZ7W0hgBVTk3hiOn9zyApT3jVUfrNsgC
BbKXzkyu0paIv4WceA5E1YNeYurLcrb5vHtR1HlseDtu5LSlsfzqOVpXH4RyBt+8ixcz54lsTzTZ
imaRvIltwAJWoXG8bFiPn17zO13updqbbthjl/7NWFMt725U3ZaByvwkakY8tldyUadNtZsH+OxQ
SPFcXWoTcp9sUmndysb3R6CeM6IUargDOQpGD9c1JkGRn+4Emtkm3gvzOQhXc30ZDX3e+tjIfwBC
cP3+DauSsywhreXuafTo++fRZQo32pxFYQj4KsTUeLkuVxkiVpGSGviohQJNTAcpLXkY4La/e/Vx
bkaQUmyjh/iWppdCJWKbeWHwPgC4H5wdQ/j9fX0Knnib9wHjut8EiJ+3qvH/A/XZPpu6BihGcAKz
4vCL8neHXxYOONaaf/3/GMoZC6cTibKyWy1a9/yLsNtafGuSzZjEWvZavMDGQCUCcqT8gK50aTx5
Iem7T9ryMD629vNrU7i2Vy4SGtAYFSWnxqD/WEOkI1TqyDmb2wqS3OyReQ5gKmBDVbzsaERX+H2e
Kn37XKKy40EEGcWBTet4nv/WLYcY6OIGHPomAF6nUmVkyH9Cjab7/wUjKbQ2aOokIJouWFp+UfVn
R6xg2/dWsMzyH2Olw/a6TzoEFi1LrQLfUY5dRIBYTl6Pedp4WJ97ftUEqKc2w9+R16zpVIMUVDrh
WO9lONCtr2im0uJxWkVZob4OhRYBkQ9m9A5QbAqIkO0PDRB913V0KcFgpd7eOKMw85PhvWyFlEjt
joHXCKPadAER4QAjrTutHa/FPQglNZ+Mp2oInWgz/7Zd+ftl1N5xVLHWMy3dk5SLAIjv9yVgqHmg
9xTqnyAkv0065csBLT7GYx5uTfvZpyXHEiuYDpxcGbj27raTh8yenZpnr1gcznXpbLxTRnyo3eBT
utabnCNfKhGiWF0+TDcM865Ucw0siFy6UjDR1pcbHkg3gTxvmKt0tvfVULx7qJYW1UxjiCZwgVFU
dpEu+VWfbbroHbwv65VNHgdSF/MMCI+sAYabULtqOY8Kz/H0iJljuaWh2zkLEU+0ufzh/37kzyE7
3OTR8iy7oC+eREL46licI/88nQXQXNMH/eOExADGH8e922bkUD/tyuUpSXCWZMWLv8zzAscfwruy
ODX5Sbirq5mryNQwZ0TSFzu7OUgX/PfRDEQxrVJrt0bFDhlgHExULzXeltWPQShvol1YTL6KIuPA
fjWRTRlTxJJGqmn9p9tbpRKkNx/2PxmChU1ai5CgdksEkWepEGaBrWiYYkl1s6WWybbPlRNTCshR
EfCV83F3vdat5ZX0yBeTnyYBg0htyv3agBjjQ2nmvz9AyokFivlaoBA7znjvg0Uiwk9QkF4kBSlh
ncA+U2UONERvFDmUHDKBKaCnfe68IdyWxQNa8yIO3NKZpxoWLs5tGN5b8bisESoIPzAG+Mt98haW
986clxnfsoLLsTMj0d8lVR39WFHA0wxm7QJeZbgDYw5j80bz9Nmvaa93q/9qThwgJiDEzfsJ7rHm
v/Gr0NHzacBa3UKgOTokkDuUbYWOZ3YraYWPfEpfIT9KbenoapaTk1MEbyM52FHF141xnyn8c8Jj
bTsh5kjC+2Pri2z+xF5YVeKFazPCb5D/4ywYPJWhZ8YTSvG+ggCdSvO9+xXdD4+uXMDXcyyBDh7K
pvEDwcWx3U5HzWb+MQkZ57lnkje6T3b5r6dybGdu/nfD0VK2kTlrZeJ+0EpfjzJ0dh/Ah3zngjSe
slF2o3mCOMnj9F5lykSbdsMux5aVBsUZT9/Ry885zhJBeW24EqtbrjaILCp4wN0rVxDesQ04D0TE
3jzmcmxSFw7tusK7N6FVI/I9UyjAM5ttbYLaoP+GHHOHI6aQUnSOHw0CXrEG4qKtQ5bXo7rHxEBb
crG4PvIhy4y3ve7YnxaoQ2svOYJRkO+lOZIv0VSJ5mea+l06aM6OQPiLKNGb2POSVhOfpk2f/k66
EPDYTRh80pHIf5EDK0ViCqu9nLWzQQj6okFWYPq+YDsDmUl68Oca8Uq9WZrUOoaeiA6EHVm4KYVK
vjuP33NhovOetwBl813eZE65OsyCR6lzK+F2Xqb1uzneqXQ9dMyOdmi8vwyFBcpM5ErOw8FoXFAC
RuYPtEysOhgGbHaaw+vqup77EFrX/NZ2+Kr6PZ9NCBWkqk2wZhwVNT9nDmhgjVSnvoMRlkjUdPUm
LsUD0f0zmGN/dLoYKVC6uR2BONgWB7I/+4LcakTLyNLNcJdZbSvIXn2ufizK3+/pOk0MK18vPqcM
466kzWjQHhxrJs7p2zWdTxxRoPN6poXsNASk+ZhyDbAHy1rVlyfLleBqGrPejO2o7hSs+FeUGEtP
j9YWOBSU/MyJcC+YJH2d/+7IHr+ghut9yDBvE7eKpozy3xnDw1xqmH153L9t7cFvogjrBeceHdMv
CnCN7gOtCcZWmYQyV1DPROFaxUvcAjYvTfnOy7M/9xTFQshuQEBA08nHyDUkxjYE5WAAbM9On1kb
U9XKHmLJDTgtPNrzTlGMDoLCJOI/PrBgeNGVhbTBwvlEQJ1VZ/BQWKPHXa1w1M4u+vu2LSBJ+7fU
wXjG7CQfJzH5EOOyWSW/kMw/LFvBVuh+xEc3JOLmXFIWk7zL0OdEnokzqLase4Vd6m2whz95AZXA
nC2qynWrtiut5bCHPNGmf46odReRPmsRUUxldsOv2E5TizoP7x9XTE4+e92+0kQJsJh4ESKojLg/
Wg84EXJpMAwDewKoMxySKtPb4AXEBpTNbf8wI4NkiGtzBYO6uw/VZfS2RqvI5CTkwc2/YlBqh/UJ
5YCcoXYB02qAzPaXkaL0AviIlU7bFLGLC+GfaLp8crr+zkuFSRRr1uMKLmjcz8kv3/BZ/egblHxb
Ze8lXQoN+OWtKlDTuqRoit4nJFiMy7pcwFSK5PxXmVzFLj0R77aOkk8Dot4/0v9bOgyb85DhFRpI
z0tpth6CcHbiGnNc05kT2SUdaHPERU0diC91EP0so3xoYgwf5WNFZIbHUoIlmW9+1UsfeZgTP/Xo
m6Zga6JzHQF3Bl88XGMy9BxDapPI7VVW2lU4+k9Gqe0/YTtW0+ZzJ5mpaMBbJHgWaIFDFKHZ3foU
POsDomPYCHXsfPmABdp4hCv7HeF3+bMMOiZRUBbv9J7RqzylXYKHhAbekUMq4qzIjKsIBkD15dPH
MPn4bh5ekR/3hBZPJzoynHW+ilDGtZQ7JjCgzCBKhY/9Vh2Wz9UZFYubkQopcM/vi7gefIUIdqp9
SQ4z9YUpO4M9l0Hava54BKbmwhl/wnQnMX8ZOr8KQvMvygxE5sEg5VjfPCFzlZ3E4qp4NuLXWYQX
wYzYlXaEqNU9/3BDM2Tc1XHxNAKmqCXeNMsoWqm05T5scJ4Veo/JbRd4EZxcrIfJ2sl4dBc70DpS
BlUv67gMAWZGTENz/fLU/1j/B5qG9CqU9U8vCH4FOlllzAhvAN/5sYekfbZ6cI7S27tIHKEg4IPT
vxwBdYsfSsDrCjF5y/gCk94i7QuDCa6y/G4RtmOq86ltpCuD1nS046IX74xsXMaolpvLCoR9xAjk
lgvVcgSZMNV2TpVb/tYO/8soLAqV5YcM9g8YzikiOUPpj8GL5wgnEqyp14qX4DaV3/L0tuRWqIzH
sfDIQ0GdAC5ct0SEm6G9kTUMyS9vA7Vl2jVy48nsaYJWE852hT0xRn7KDZj7rR4PCA4cgGtQ3Jkj
M9yX5/o3r67mEJCc/Nwi33QfJEq3tLCMGJHkSyZLLGcXeGApM2ZQ6QAo2n4g+/bkfDIz7P4Svcg2
DZQpKySUEnUmCRlajNjQsgLE/6soO2/K9SZSwndBU3mMVSitdETpVKlgoYxtW7iZnWbfF+byI8Hj
G22HApOntUauU690mJJ/bFbsRgqsoh985IuZaNPt/JXuICinrdXUF2pDPNFShsCrf/7crlWurUnO
e4RpimsAXH/PIziavh2Hh5ZbVS25e62DQoGqzZCS5M9/kAaFUcUaGj/3j0WFLr2kssFyhQEtz9Ib
PeJEjfLgqHpuzPYs95CIIl92WrgE9kOqri+5/Z1w0gnG7PeSl05blLpd4o/gC6/ofTkytjhvfvra
GAqPMphVXOafMCTG+0ChLb+garQfP+DAdAvtLRb/LDLisN2zNuAYesKzNA0e2gq3wcvO1NVJAzkr
hA/MvIIDKQJ8AUhOEo8wCcCnGABxJkdKAmTrXm1/67UnliDztdBOM5g8DkKIaPkBzmKV56iQkUPl
BZpWozftfHBqa4G578Nx9NB1+diL2FAYeSGMp64FySgxG4O5BvYclg1LLQQynO21uqQWiaFJtECL
04VksJAwgvtILuiV3nMhATIWJZ/IFjtWtcIEENO1Z8OKF5RA4anUlaK09VXoJUUX7Xw0jkQfxB2n
f8PITvb03zXbLijGVRi/o/lHqIQdA/cQeIBMR7yXP2VWm0JnCfeh3sp0FEXMLtwMpTLIT9jEjp7O
03sAr0+lKQOV6WHpi2bn7vRcqi4kewx9tKkr9g3CN4mdMqOkMDgF+muzpQ2WlNKADd3+IEmNMQZ2
uVw1D8NfIAh/yiI91oT+s2rmmATwdfYX44QuEgJLIUEo42d6ip/85EPAHiXqeu3GzIeYcgZu9xSy
Qgn4gnmqawrjSC9g9/nADxsJwPoeiRvVsqU3CXzrRrSzOMGwBRQApTKwE3cUJ1dryU5gbaBG4a3E
3CMgp6AZqm0KuDAUBCux2CDRvCzJ7tKQwSuTIa0KuayXFU151XBJegH++LJseenYp48GBO/G9itN
/18qeAEx6ygWUPyDKHiog+hnl9KqGJcatsPcHwf2nWAQl153VitFyB4knjl+lQnpAuwQ6U9DpHvo
+8w8RieIYJ5tIoYtQ/gd8ioeglPzpsx/zcR6ka7KdcHcZWUb/NWW/mCacqITP4Yj0SmDR+vUAo3X
pubqm7DDmX+iTPVGcNm8TlGYrI077/5hJWJWLLienqbtDZIHlU31PlVGMxcXuccIGkvEqpmD05hD
rXZnzeajqgcgI04djZBQy5VQZZOI95I0f9ZpHC0Au7y+EHJU6xFmi+ynIET0e7aNYVTgJwBUFG9y
4Ot+BrxX7NFyoc+qtlVjYbjNj3IwiTx4X7xA/aTJb0T7E5OqxS0kkurULD3r092t7vC1lOk7FkQh
fG3oH0JlKvM3q1Un2ZoJfs50aQ5ciKedOSk+rASDpOrxJhDbftZOGhgLWDgKNh2ZaiBIjo4B5nHM
adDwPTkWjgPvKCrYrHDM/rBsb6zC0AyL5eMcxNJuqTsiGQO51goUt7OBePAct4JLv/8IJuo8+EG5
pyrYwKU9DaOHicmg25Mmyl9vBQqc0w6lkjUBlUg82DTpNvp+P2Tjvso+AtRVS9HyZTCiw3jk3sNM
hiJrXYk6+QZe5XSmgngXgCgDMJm+X3l31tf5lzbdS+fqkf9E68gko1LkEWsKiSoW5DknFAfaK+lU
z4TA9WA7bpLM5EwiusuOk7si0hvSiKMOeZevcbk1XfYz0PU8ihyM0qY8uTDx7a1X6QnJniA5YJhb
B1trCSgKrByIx3XjIKxm7ghGm8uPaWxawp/JXOSgj0n11p7TvfdyMsNYwfPaasNI6a5hvHSjg5C1
LI3C7GFFuuZnty26q4JbMV5DSQiZ0IYwEZ8g3RICib+uS4o7KINHyBGeYF96E5gdZ+JMjwfWcIps
mrRw9cfODOY5KZ8od52YID/u5Epm8kZw1rxt6+fTL7sncZkYtwOumZnb+4AQ+XBYPyNAVVr0Zww5
onN/qrDnaFzjgI3nzTk6dg+Y501BHRNC19ESzUP3CxTnfrjoYAgQwpYnZ1WFeqT5aoqLmv3ThDsn
fEcVJX0BtfG1qRNBcrt2zrSW/8uLFPVqaMQ5EtaasSDMfRLUzxpkcIOBw7+YMYhZrHNQbSk3Odr3
yUHOhALF4Nn+v11b1nIDGpHdZM+1HY2F8dNKsq41XsD1qAmSv5eic3GImv/kWxCy5Xyahyd23R8W
CgqM307QfN0EOuZelCW0jtA9wiVk6p5cZ3Lz84KL9AIhk3mMsdVSIVE22KCQ1tRajF2a7MhSxfAT
MtJkBb7rvkwpHCitm6wmhiRq3ih8DmfI378I9aBrJJPlMFAWZ6t3rYHvT4D4/4hlfUwUGPQmk99a
cwbUJdEY5X4KVLwY2XLWxQHD9a4TaI770N2K+t/etVauxx8QoOHQXxV+vRn/KCtmblRtfOiTJEDM
Sov3PyHac1oNVeqE0wKAy5tpC7AZ3Kgj0OY329vm4ej+l5Xs95huCQKENXsfMx28AlkZHsaXMV3h
4/RbbdX5E0sJE6ZvpZoS7wQHPxTuIIJltmA1WQzwT0dM6R99J02iRV/cpTuSu1jpay/BT3cnG/bL
4qwZMB/6DD7T5WvSTr/zYu72IRaDHiCYmoOzD3f3CGs891OGsHgTwvX8qTW1sntT3spPmPiN9VYm
FH1xKQDvvzZKtwJ9WXu1KQMMKmpDqhNApK0JUQxXIeWSaMKNEL+XX8DkcWrAxZzRJaRqmjUWHhQL
7XwK2Bmk6qLDeC/avOdTj9Y7N5JsOtPrQfTgkUG6f6NiwdLRZJ1beHveUDD9uRuUhtkHEJK1fj55
pX/Z6ZOD+doiUVTJft0x21pMNidNTPOEcctCI2u3AiOX8byUM+cPhyGC02+ud8O0+06TWkgMcFkf
lSJq8s2uAU3zUk72wBDWSgV0vqRfJQher6Zp8GPDmjLyvw7mLL+JcFlDjsCdIzoE1r6I0CtBywOO
SlqZqJBTkRpTCvOaXMLhMBb1gFAzj00zdi1Yrx1BNpCZHIwTWTwLxsMPAb0Phhqdqe8mvux1ATwC
pCSFHvaO6I8uyoX5IY1FaM47CgxyvwZG1Hw+QS96HZc0DHuk2nCY9ZIIWSPQIJMCfWQxpHOCS8pY
lysLKIG64ulQ/VIIXOdg3umeJXHprEirFbMAHxMsmdGiVQL5Eti+Cz78d1XbZ8BSFrBrHvcM7sVT
LxVQK9RiNdNnAD3uoacbZhu0WklwnHbm0uzXbYB9R+76UmBsk77UBkRxqt4H6u472Av2Oe+JKVWw
F9lXjkmYWaOYiJltUb31dUvPvS2mHp91o7o9yzF73ob910V3+mmLYRSRBZS4eZyrVnQfBO+B+06S
++MpuwfnJQ3Pgs8SAdQ2Fpos3yAUn814irxPK7PYoq8SKVfLbom+mgWFODVvF7iuKLImFyF0hO4/
EMlUD0I+xwbV7zWvThmrgqCZR+Yn9k97jG6K8+qsFcsmRHQj8diRSaJuIx2QbgVgvcGwRJnAfigY
FXGt0TIGJAq2XjZ6Tv0gSYTk89jrJYdkHRFIxF7P58BGwmDhVadXRHWatx2djbqPrVj2acIBcg40
+gFxrelp5yr2Efe4eaNxl4DaVs0/0y8r7HLRKXAQR1GXuq0lZPxe4NKwNTfL6TR98j+V5Z7KRB2n
p/5cOvdddsbAPpi611vMnNsNqJakF1DX5xZC8gT7liGWyfyh4vEJ96xMvjofEEg4EeH6q3SPef1i
WHJ5xX0TJfps/8+ROn6/unW/V/yJgyHfO9qPAN6ZYA4gwg86GG6IICoDeaYB1LlOd6jbdBrEAXSJ
V4Pyb7x47bgSD7D/UjJ4Sy+8FannsFKH0zbocIxnUg3DrDWFoqn+Fy7UHjKxc14KfJZCOoE01zaQ
Jzy+qHhNlhGDm7gK7aNrIIc+U4sfBLtihfu/kxRhLNCzYaw4F2ZybMGI1ZYTUztapVoQIgLUgzMD
AyM3mLn2HW6oCyHKxfEpfJ/66CJ9CVnb2nQfUI/e3YDL3FqJQFsHEgXguwoNrPRfIawk2ASbLWpw
fGI+E4a5RRRWdjAcSwQqRymP1rtAEHckgq+vLu5OJJuVHDS/FryCsao69a/Mh2/JjtBlyqtvva3A
gY8uJTAMf+URd6xfiYJJAFuplZq2DSM9Mxwejx2s6gc7QMSsOnWnMBmZ8xd+ZJGnm35cJDC2+OtQ
sJzA81pMNXuxb//vwwySgx2rabiRTMYDH6OQQR+kRR1Ea+mqA+TwP0GjqZaJ//eNR43c9gH4u9Y8
47VxhTXU0GsDrpz59wgXoTPJxXuzkEaol6KwNIPdfvl9ntHSWrqOWD+7X39JVBzNaTRMlDWQFoQy
SOvdZEMcouiQO6blYwI5ren7mVs013574Makzu95pCXvB7EHvG3jReI/w86SqGWFG1fP5MLnkASq
lfiD1GEhOETls6cpiRhZGIUtYdbe7xSUAOxYsoQ4KSo/SzEzXgT8fDynC1zczHLUajAKtUr9+HGX
bNNVINbgl+Y16Wvn1fnwNOSkhFFWC9zsZar4hJcHPXQLmTMr6JCwJkcVFjnNLZa5s/ymyPeTNLss
+uCiYapEE46jahMN73/oqcewfxtLAS2l3AUSDzh0/ZtzxxF6NX+Sx6orlDNJDaE9AdoU6sxdjGi5
d8WlXlkeApWOkCf249Psnx34m3ylDpkQMqtucSdcVGDXMBc6bmhVcll5Tb2/2vYTfcMPymB6a6tG
+eWzvzObS8iuJCpg52p20YFSgtDEANbp8iVo5c88/OoVfn1RLOih96o0vfpgI72hhCOfakXVoUFh
4UM1ZRyqxZDS9q4CERCHFRkTy60b3kb549UMifw+dCg2kb/E7mOeA1v48leCkA0aMD9bwN/vjTvS
po5wILUxi646ehbTAhbafgo+qQDSygnkUzmo17bekuVmCkhHTO9EaalyDmbqRhqhvv0fofPRDrCQ
WnOTfVCDraHXd8apfaBBjnDAPRczpew24kIe4eOotii1AyPs0VB2AhkBuFXUEnPmngk63tmOK/bF
Bowsbnf81dlbswUgHyolEywyhPWF9digy6l31wrQFuj+8gJCeV/CU8Tc2SrfJMrlqz+tHgozgKr4
mfq04AO0xyjh/FxVCdPYuxACAYbxFvJBqh/O9/F2Sbxa9BXTTbfLKb6F+TheErQyAHPgO0RG9g46
xEchyPg+AtL0F/4O+I9vRxJ7rykiUuKYlCaEILegyOdHlJ/PSxnzlidCc8KkLrnoqdSqG96btjPt
AVBk+v3eLHtZo9sf9+MqXkR1bZaNe2XvOUyxCxThcNXKqfo469kWQkYyf2vilBBbnoLRyVNuj2EI
WKMvXBWsboGkZrIlzJzJ9457XkvgYuAIuyodeNHx8CEpEhQMagxb8FfzG9WbusDEEj4aA2AONcEn
V5L4TSrFZO+uzzsOZbihwqygOKv2nwk3/3CR/r2J6jSUL+RmI8S3jA6wxzdHc/pS1dNRt2unRdxf
09WebjxWi2svnBJ9V73R8HLIKgd/uZmubcXH2OBxY5Sb/MTspX+Jcybaxcyh3Ys7ezlLW/icyWFL
h9ldCJ/qlLMFJVta2lfgGrYT7+AcT4/TUShInAabskfDMVvuDfrLbPSUm61L4zgNwIMoe31H6CY6
sTYxQQobGM1vzuWREcIFybTijY1SR5Z/ooEsvV9mTNORRyNyYiW1WNoyMipcGx4e+bw+CY0D+N2D
upj+36vqfKi6eE0pcaHSs2MD8jlKFdCWAM8etjXfnrB3GJiANHe+mYHsautqwEYDMBpVthL7O9S0
PrP3KVj7iiU/zcV7AnofhPHZB8/p3V4QmIgQejiUGWCvCbPZ2mpHUbc50RUxnuTaDhPJHpcGgNT5
D4EgiRZkuzyuqkRTtpA6beq/Rxo+w1JOw6kI+MeOtLlQKMIY0rm+Sb59feNpc0n6CKqoVTjWUBdK
8TrfYyvl8Llvk7HlnlwZCuXDiH5IixWirv6Mn6rPAy+6uJzWFjhScK+glZTcsNlNyOLog+DoB1zh
+zHccSLy/fth143rwpUwUVG+Q7ZHA1xERLCYWtMDTxG2hBokO16Ii7FSrfllMxrrqqyYn++wtRMd
HfP4SD/8ES9Fao5bbGgpOwgaXPBPUGVZwmkXtAMWrZy5sXoMh+SZx1XYJwEM1sqYTUcsM3xLrXCS
jdwJnpj3ImVj29fzbDHTMeS3QcPanitB5a22R/VQ2AdFkH4BpV/k2BL9gDWyEfm1dcaaB2pRuqwh
h/8BFR5xS8j/QkftfXLydO4K+cV/N99t6OvFhHB8TVQhz6rwISdrYFgQ2YcUwt46E/LQxISdhOTS
p9qQztqxL6GiysK4fJPKfv5N61lmGonRl7zDN0F3mWTKhtiVuo0lKFw9ySAVKsHvxx2QLuwAID25
4f40aBPsNREE2/gk0yLLatJcBYJg4ouxPQPa2ANGcVcuHOd6yWdu8G/sErtBjcG8yaQVE/74BXJf
aqvPHscmej6Zj6nl5oat1MdcZlTYw42NWRUAIHMlB1/Vu2uRUnlp3WJRrS5Zng+G+xML21QmVilS
6kYWeadV4K2hLZHGJn4VSlgGBhRqHSiqBBsXl55YILZMqp0RMbDrGocyUR7tWUTOWNU6ottbezQu
H9PykVurL42+MGdtIh9zudCyAmd93zIxZ3Zx70ibwBUaEJ0J26RjCpd/oWfp1hZ3EvzJAwUEQ/nV
0xsbI/fkIB5kg3Ni5CTyLeGgnWlJpbx32Zw9xYemHL9iCjZ5eSdTDskWvLyxAyVLoCH5kVyshjEM
REc67AY28VaGh9xSv+T48BBGmyie89pNXCudWEFSrscnYjw1XYUBvPrro0dFygWb55i5P2R2CKpv
WXk6GdlkdJQoxs5JFV29Yayx8LDR9eHQKLd1Pdg3rJ35oMScZarmG5z2qH6jTEvKXZZCj4z7Wdz7
l9GoD7MTqSE+ee9xr2/pJeAEPDBDhQT9wG/3+fhmix/t652BqGrdi18OruXKsaHnkDZwx+3Vq2na
BSSAjTUIrC12m5GyQHQTD6dB8MHQfSdF+CExxu5AsiKld/RJ7I1JG9hB/QDm8KB7J3TROywKp9b/
a77uaBxXbB/EDGrKx/nom7JZt+2nN9slP0WZospc/Bq/W1LLCD+EiZ4Gqb/Qt12h08axfnfg0CyG
Hr1Wz8D3fZl2+MLEY61nicFGsLxVFHopWabVMWCgOqtBB6opwcBzc0xUzOO2hEB/R0dqjFaGf9RO
KAURcepfIvKJc6hPmCBjeAxla00tS3cMs357hsolGO47bhbtQWN3ur5/wQOAGGyfUArDttNAUunG
r9S51alWoT5yP6Vxclqa5yieb1rghVpxjl/NldEsapQ8tyQp4h55fRUK7i1pMvR+s+3g26temOYY
+VD0FRouMkap5SAPSf+ZNPRhjOgD+14/LgT7kGu32xyUaTLcDXitqYs+V92egiaGgyZROpc45+0m
FbtTrickzSwiyK3rCpUwih6v1FuYfCVDSfofdV6ed4eXCi8cUySRKUTF5Lyd/FCxIB2T9aM+Z5NH
UkNUIfW91uyMnDZ3yfHoCAtYxLGibAdpYy831vVJAnu0eMD+qNC8REFIipeaAW59TITsqKqZNlvx
qmTDQkp3jw2Hh+VeIKOJwhcmYmiR1jgdS4ogkwx1Z2hoqht6QVvevj4SKHrlDvEz1zqH1rbK22Yb
b2Xyf0/9E93h/CAZa+4SjytvtmCA6OPtMLHxScZGI4QhHu83wgi/OrjdMoXTECdsNwPw3f+anqvL
r+NyH9aGXk/7FENrB5Zr+ftnfyWONQkhy4a8aVvNF3XGQHPL+azG5Hd/2P4Qhu54OaaRli9ZjTP+
WXRa3HRkr5g2caG+v3uZDGwAiHHPmmkerCVWeBUanKkMqt4ujNj++A40P791WBC8X2wdpIDkxpwr
wEgtgzkFcYhUGK25x7NtCTKuSMU3ogNcliULZly5qeJFXrZ4gJTG46V/8rSlDPf+pSVzBlLw7e8u
Tmb9eQd83eaTnhVxq0hWjMcor3nsRhr8rVEQ9odG5kO5S2VDyTeqvtkpHEPGWF8yd5YvXdic7mEx
D9rQvIK0nD2t0y7YnOyABdi/Dq6JSuLiJzdNbdfnIbiOQgZJd/8Q+YMZed36n2owuA1I1ps8XE/G
SOAv2MXEJRX/bqiTWObsGRSiHUpjS7sgqmlAYZl0thZ/t5lUMkkmvmCpvYs6YJeKfpyVj0MYpNBc
z04glRP4p+sDEu1tkBRLFmQtnKHhDy5g7PbyKq5jTmZHVITjOkxjx8InplZqAJzKkL6mWDKeqh4h
TJjQFI1S66dqKlNE2whiBIYxtca0VB/U4wrv/d1q717yWxd0e54v5jXRt2zxtAHAOR/pwl7l2i9W
lm4yARwj4uFSVpvV/bSTdgkvoy07WcvQT3DMMdXiwEoZZ+5oDsGAeOSKkLvMXPUbvsB9vqg/3q/I
8iLRimj5KuaFe42jW3k4vkwYneiIt/3J81CirXoinOGGSmxha7QZo2JgXf2jx0Jl9ZDoRWkb7D+g
yMktxHjzqQFAFO/f9wsUjllzf8Kv0/KFvbTnsQCO1eyEAaBEyzSDBfnveTfOCeuroN31cOGEv824
9jbYXgbmq2a8WZOklkZ//Z7hwORHxP5HV1crNldisG4XiqSx6WiAcOaHTFuhIWoTufOUHhzPple6
/Cpl9o5h80rEWTQ+MdSK6tSEHonuNjsEy/2TInGgKJAs3WcWTACXK7GFLIYboVgwnVtmRkRO0Wgw
c/DN3ZKqkzdJVkqJOSPymasr4rwy4UgX8GhTMxwlmTpKZyI0OW8sEln0WkCWoS3ROJYU8TLSZhhP
b4B6izc7rXTKkxpwRQh+EICJZWfORSK9c1CFOzZKpSWUdD1JnPqglyvLfEryTUeWy0/5TGLhCQxI
pXOLQJMxbUpvXynUcvTlzliBoxn2LCh1K3Y7d7u/5YJCgp9aL8Agq2rD7d2ljOJxq6Zxd4737QhF
gURCOwa4to1i3VKL2Hfim6R/z7VG3xXWQ7R3FGrq5Pizb5Ben8UBqYMom0Wikhl5QaMtMup1q7Rz
rbOIYMR/gluQspLZCEf5BUfdtnIkz6drtEZT9OpTz8iaRq4fWruX2E3VXhUD+7CrT19R3S1MyfHM
JE631Qr+Go0luuQw/JwGLDemZgy3uv2KomYWMjcuJsjM/44ImhIRTvJQzXZl48hm455V4durUUPo
p/zI2b1xNDxYNJm/i8FZuNH+8LMMn3uz7LOQmFmYOzXqhrlsVEn06ISQoDmXLLdKeZjryAHxrwi6
R17/JrL91oMEmmJrCTb4umSiQVNC7+2NQ3pTdjc6Hp/YPX2m2WOV9PFrqT/6PddMMN/05CZG2DxS
k1vvvpDoEGLobS9k9nQerhA8STm9ld8UvPFP7DsBSV0h0NdZv/WtdIPIDqeh9bD5LKwITy7jY6YZ
jrYEsG7TSSYSTbyujwNnyevYcZZWBHfskTMUTrAtznMtomtbLyZeVLXe1R/4i7SOjSjDq1mfKM0q
039u0UfKLUQS/x0s/ljmfwd1+gPAls3mcMaEFJUm21a/GJgW5rxtNvFuhosMzuKWZQ8dXxchW8en
1Xlp3rmN6uZuYaj5Yjd6d88fTNPFdSAZoeATDXzcvU9lFMtN3ngR0AoTH27xOx06j3cNctfFt4ML
2Gxxg+jp9X+Gf/rx5QaDW3CQFhR8BmNUkWB3s4T1XF2PTkH1/MHqdDevpWl71RkQLB6xMa/XurN7
RrF3P9JlLyDV0ff7omR9n3b/jrQawzt+ryf7cCQkCtZ1ilxd7eyvDZqVYV+UKeXMTgAF2m0gu8XK
SYx7qUy0vfIwsUw6e7JA8qDVUza+5Nnb8izfv4aev1dcnA0zJ9Xe4EqyznSQUKycPcMXL9pPE1M1
BtYtxcuIrgHNIjjxVeEvhnnLT5weM5t+UFXcSeg40Xv4qQxsmreV+xFkuLOti6AF6Xp/FZoOZmi+
ZuLS6icYY2d4mBzkPHNojHRHhGnNFkg10F+v8iN6B1FQwphuG9iFV+2e/tfjMtmgPf/WemSqnfhu
XK+XbDcifSDXA+slYEodJ+eF/DZA+xUYgloB2TI4bXf5jn/1OeBLAGtsHPXrjxUn+qxhS2XU3wxz
2DB3utojYwKROSgtQswpvJ1NNmX0swXKM1SpCBhLAAys3Z3v2nrndi4ZYUkT6WIjbIcSK34ZKiGl
16aTBswrmq0ZToQCU/VDKgKNN5dtMrqHP5zvmWY2hhpJYd/JNBJ/Bhxq5UkDt2bSLK05P6gqc+Ms
3r6G7/KLwvHUFj3kv6ABPvQDtGXqvWM/REyyUIh7GQO4mdV/MhmOA5yBtrEKnQtr3nGexPDS70jN
QcDJ3ty2u5Lw8YoxLJzAUzb32qxO9mcjQf5ELWgR47tIQcku5xzahqiNElJeBcP6Jo0WGXWQiaQ9
H8NKBCL+P1z/OA+NiAYeLo9XfeEsdTfYvisb/wcTaNlxvyB/asfUk0GNSZenN+Txlr7tsKzB6I0K
UwLCEXocX2cnuq76LjBct/4YmaKzMM8gTzvnsxCANzjqyq+kNJ0qCf/LuVDPTD67hss+1+KYwfYp
6bDElsG0YeITPL07wAxPAfDWQeulYd5eB0p/MCAjdLplza7XrL8gASAAmbXnzC78765Bod99LJKI
es0JBnJawly7GRa2Qx9dxoihKkRP3P39ExrtACQ8pZHs7JODzrtRy9mnTrEAKxyqQ9k/cmnjfLRB
jgdTG+alFTRIc2/lZimnLFeho92DtcUlXHCe+8uUbNKWvKTzXm7UfQdV17mOnxLzxhwvYFfIW6Cr
7doP7R+i0GlaHqToRnbY2rMhWh/X6ghLDgqZmGvByasWKBa6UBKtLeVVEQi9DlHMES6BJ63PSnif
nX0OFVG4sovGdQsnI2XhFchLGpEJ04EEtS6YPoGH57iqG83NexrYg9VG1TsjTLvzOK8lhogOJEPm
a/R48Q1/76R8fuT9waqgTMT3OUTDTqGHej6Eph7H69NjS7VRrk8CeYzaY7Lkqm725TwB3d0HxjBZ
R3PEE6FlRQ7uI3UrPFVI/HJbSy8SgZ5eyflDFVhhomJLeMDzuANePbCe9Qtb+po33O2EmZWMHw4T
02i7RGuZCPE9q+sS633zJkLvk1yLJwJW60FtlhyUgGntfxgxDjCTfWIXwXM+7Ro2v2KXy0x4Rtlq
pUd7TqbtNeHXgGN/ts0hR4AVCtODEGQl0p0bVvuaP0ZQB0XJRQxz4RvqTLo6cbMWw92jaZKeEnwO
dW8nhG6WL3DZBW1Ks0gfZLzIuu13sIxJb9Wy6QExNT1H/LMfW2IE34aiUo6IhsCw69O1Wbi3/Q0z
QNSWWfh28zbGCxUzXHS3FNg97t/NsdYTciSKM48CHRcSOrD0mVwq+ylvaj7WWH0l7XnLs9RgDT6P
V/7yPEKYjE3GV7+L9nQNupodQDlQ6P0sh0uw1FxNFQg+akOTNZJorDeEHkJ/c0Yc5ddkpalEf0Ax
mjqWTKjEAOVReNt5qprk4VrOGldYElEtf2UbRjb/1E3xpDxO1AnZQMMkzx/y8U27ftbyCDbvJqCX
2BHQth7XxZJBx2th7PC+vbVpzGKCZfThoJ8CYlwr1OmPnu+j9qbAJG1M1FLnZfyU1icMWMew/fhw
UQJXJ6TVRBr+9ZgANxLdSqhwQkVO9vFPYy6w/m9I0V5jhldAyxv+6XsUmt+14k6RZ465E58KYEV2
PpWjhypG5hmmpELCSqfAyHF+CJGPVqCP5gTGdEZH5nSs7u4eTGJTjnSG5tBzQrcsYfU5mBrfiA90
UMc4gkB3gSV1uaiW07/zVoAFVKC7dM8yXa5glQdBy/F0WIjMVZUsusTQGtSzlewTSMPKUMDLdBA7
rsZPp0LiVP6rGxLkbrR9Z/NJ0feesFbKtK+iXLXCEWHdPc5qIOCidBdgvNPtxrLHTOtKLPOpKRuy
QIFS07EMlg5kF8p3fLLAyNXgqsPbReqf1CyPtgGBcP1E8nnuQ7Yo83ioTh05aqXb1izaq/fwEsoU
4tXjjjbhnZh9YS0+WL4UzY0uDfY/z/aW8OqlGhjkn5bfT0ysC49oG3n5T/EtOWZyGlMFle/MT/Fr
f3KY2urWoZgXA7Whww92u6KyFPMu0RWhXYKjXvlCZZ2lgRbZCQRMRMY36Ost0oczssgaBvSKJeRE
CJH7LMUieSV/NzZXe5IX75qzcwFXfeWvgQJIl27buWl0L2b/uKszPtvnE0nbpulU+dqXq9qZZLv2
V8gBp9IIY7+ePbVRDAd4NtVF2L4wXfojlsw2aDiDvkCcmOQQBK5qupKR6aASWej9Sj+IKjRX9oDT
ZFA0qSNmidPf2DYHaDLKa+1la8C3TTqZ4CZI/yzBrB+EOWB4zjnxIMnFELl7idei2xS6BZu2jh2x
zrz6+GOPg5E+vUNb+LNcJx3V9s+b7aT4Ggw5HArO8dR/9vdMlf5ApRpbsV/NWP6dbJY0Kab35G8j
PygMZ06fVrkLUeHKs16uK3EmAlvyBkGTZmotv2/FUMR6E+VaYqeENMl5o9crJ2W4v66269TMorO7
EBg69BFJMq0F/RHhrpoAc02KhTcNzc+mC4O6WXcSW2TFy1NcEIqCLstJQlplXtHFBr6LsnPMHPBT
sG0I2FP5ZlUo3CyT8lAEsjHceWaYSrhQR6s4pj/gw1c8J595fQxkP4pkdNWsjgGAjfUse5obKAuy
H9hFl3D9uy4GYdVRFIdcyrv3Rs5FlMUm8+3UrXjmuilarNxNaSZ8LPF+qUit0SF3Z5KCbh3vjRND
gYXNmEw32N0t4yOrdG8H/HHrW6RXtvhNXrAnAXyWbveXa7UoYVkvvRzy1XC49+PH9pjDBheHHXAj
Pp/GWnsXTsFmF3sE2QeeQ0zSs/EqL7BurdxZofQtf4/IgaTHuSg/nm0GRpb1xyXu+G86Q6LtLQxX
iLdpLPUuHpmH7dehMj6mEVHL0SIlbJPphkvK67DOF3E1y7Gucgi6p2ZjAUr/6A0qibSbT0zYFXWO
n8ibIeFYxarBshtagryQAr7IoE3pbjD02tpngT5N84IDNLvkVfPoDSg4G2zUxlUupFiNvf5R9DHN
pCQLqFY2SiEJB3y1QqjY4jCaY9NfNgCmywrJoS3rQSS5xp9jBtfaN/sASsnAcfTwchRThC4v7ld9
MvEa4x6oi+f5GjVxmI5bQbXx8MYGb/Y9sYConkIyUB7xd9cI9sBCYIx6nDTWe5kD+SAtbS3NZwEW
TRfgtaV/SaL1CgT9zI9ovRTNQGY/Bipu2C6qJLqX2JwgC1e8eS7170kQVbWVhUCJWx180S9PXgLS
LMHsYFB0kH7PIZBgf/MP+9qOMaWY7qxyyu94YAalO7MXI9QRusFZpUzftQQkFKdPmwsfwFHkN3qn
K+Y1s8w+ahGgVQwP7I1PQm0rnSwbVtNycx69qkMsRhdQ2eXr4UMfeeY6gWFUjqO0gwarfB6nfK8/
c3wOAMpPheDesWPAgh+we8YXWx393J4C4DoPaaRQuv3lVb+uF+vY8pq+S7TPkvqfIqlqlMkals6t
bD7yFvXpGwT8QwOx9Kq///oNwKF64yx8hoog9gzXpUVDCdUw+P8Zi6bjNz6r+T1lwicqFa913ZdJ
aZFqp3Os1KhcWWb//H1jBP65y6Yviqar9edT1s778q0xhHQOy7SzuS4iM4Oz/BmZ+b+9yoPicpsa
PBkxA1XVs/Yn71Il0QU15uRPSC93z4rHZT7wkMDJfmovQPpytG+URO5ebC98ziK7SZUZ7vURwKA9
QxANmETcGHN6hHI6c8TEA1AkeckNikTbs6FGLeNk1ufd/GqDG5iaioocVnGRvzudzkA8rchaXn9x
VIZie78/1BGM94R6SRVUAEV/QJEkTLAJ/ZZLQt+Xpt948aS+tyLVPagyC0+p6yCoYzZ6CUysY7jR
5mbo5zX5+ESE2uKDD/ZnTQlSe6SqMTbZVDdIRrPVmIuresisFLJcI1oDeS51ltnlEKF/evdmTk3r
flsZ7Rpm3LLvim/4Lnh8Xt9INLhyMjSqi8mjCxJapTd4u7UaCk6BONsxwP3FQH2cS/rhAvMMRluS
2ke5jZxkpJZzdS5qh9ktPMK9J0awTOVAjmvp0SB6hANt/X7AzEmyQ1fVUbDvdxdydZAaVA/UyWHw
WUNmrzg1IwNCaF+xt/3b6/rXFLoztCX5t4CK/LWMmkrxNVmWFm0hWF4r1HVLG5eftmFbOgCWfQBG
3nOv/kDwLilWtsbdwz0+4nbjgrIeNQplL218JKsvExJo8NNtllwuyjUQ7M7vahp/eoKGoevTHCX7
pz2tN3ojMv4Q006IgfWSf94m0jl9+CU7uNBILYrVMVGlG5Iv6YNgB3GYw5gpphnfzEteEV5RscCr
7ONl0pYkkhzM2nrmYGM1thf/kPQVQ+nKI9VA5DOH8kKB/b95sRdMveVPVDVxqLo84ca9CkJJMO1Q
TzGVQLcQYl0nUhKBiaQuCuIrcdEkf2uxYbZF/j0AbPESTpzad8lLWlFIPxddvaBnYf+HX3iFrF4q
e1SAHdSAxwxIeCDG37voXrsmP8Qy7Xb/W/lWsHv3XDsFAtOB0lTNHrRkmHdZc7Pt5PgxAeI3m3EC
xY34SSHYEXvlVioGojlibRKNMhGnPEYi1szEsUmjuLBTrz9GmTtfPJcZLawyjmWaBcLJZjNVDz66
UimkGqKWtdXQB4oUNLsNUDSJ6Quptift5vti/MednUm3LZQFJJIermfgjJv3CbnAqJ9Wx54TYx91
zCMKfiHjk1K/KuPbQbOWbGN11YTBVVRsaqJKIlV4FLJTVuiylmYUdgADWIdNd9w35x29XExlaaai
NIyqlgAsqU3A5xwkRUbu2P1XNSd553sWItYr7vAVz897Gr7oOmLTjgJQFQd3JneXXxgK8E2XDh2w
qBnHV0Woqig6rXU7amgJFm38KlJ+Ymw8hwQJbxlyI7BBgH0B9VDdsg09NzYZ5Z5K2RfglUXAyDoM
1r+wPiEcjA2wVp5s8FTpKBhPITxxHoQ3O3KiS0Q2e4WpLVIiqPJnXJxAQcorgLCXaF9/fzp3AZd3
mIjkYkP0nB+ST44yJqSj6Yagds+HnxRB/SFd7wlej61Ql52m8/Gqxr2fMEngAJf3PMEw8ES8r+Rj
mSvE0WA/QgczBnbq2vOGiy6bZ12t/SwlSmVrW6nxTJxBHKOuZGwPDev7YkEbS3eDeSkuS0XBFEKc
0z42eTE5h3yR/HJ5K3Rpe5yah4C1zo8sXTvbCoW4QRvHKDNEANBVJbwaQxvaCwOP3QFx/Pps7FpY
tzJNHoBdA5KALo+zuQNWKURMvlNCiMERzI4UG26d3ipOIHgsJMR7JPc0OULXi4zA3LMevkZbDY1S
DgJU03UgctWpYm+i4QDkA5pX+Kgey3w8P7+C0HyEOP/fO8hgcpLTVKLC49iGmMPHNIsl9dlSxUQ0
0K+5aGpGgZmvnXXfIyVhGjCbz8mcgcJjCL1HFRiKEGIhKQr2z2WfkO39aaDuNjq/yoKojswhNAjm
pd3QWzQdiEt9u2hHQ57e73OcgQkv/6Q0XyU3zhF00gEyoEqbpMaQwuMJjuOJEIdyx8sJnte905k/
PAtDaac4rLiQcLFYRKXQdLAI3QDtHerRFOaV1yDXAJpEFPWNeChKIgCwIKbjVPX/wcEdZ7yPTIKl
ZQqMtLtQ3mW8/GeBxhzawuSHr1KQtip/kF+aXDO1xSBKsRzig+j3w4jGJErqtgnJwtuos8+IGz/y
sSmXiUoAIo4b+/KLcjm9vZCuX1hN8O0oZhUS2DrrPefzhnf7IzueSXK/OHnSY1KBjQrJsGXq88tu
0C1oOADfBxATUMZA2pYdQx5cl8GwpFjvUTOggZxwtdsvbbUqU6LYQ7vtiIEmOCZzdfuCxWo5YmmF
Rrlzkm5b6BvQ3Pi8WP6BRPuyDSGQ9/tWnYeBkhHQl1FumYDQevNnKRJSpKFXc97UqM3IwRani3gu
4SIIfQdhH57Ls0pobe89Kld65K7fE/Vu/zbI8ZIRIT14HaUyoQLfX6xo/HLzlp+ckI+SABFVNOxJ
Bty7DxRfOPS5NDbrdOKJzDjcRWRetWF8WqRzyZVusK/Wjh80HHXS3O9nBNKOIOtRV5e90RUVx9dB
rt1S7/5LsBsgiWtXV5jRcV+oTg3ipgldWeYZ/inFc51GhOIp1PTVtW5duHBCQU1dNSotV15MIyp1
m72T+6SzJAUBvLowGmh72zLo56a6bwqu0iBu2umcSjFSWMDndywjjBEJnR5Q0X98fWzkbeD4q7Rc
cwH7TNb9tfRDe7byMXstMLuMmdBv1KUHsSVZZk7iIPsbBa5eVb5VcO18RdaJXHI0PwjeUVzW16mW
+geW7eYykMuUy5g+HE+T1jGpHSNCyew1rLlh6MGOQhL/y+jLiP9d4FUQGPstXsaJXtPKew4ryBo3
9wcJLBH2NvBfaGlOKwd5eXl8kG6c37X/NfLTZ7l2rCPqk5xrNBZm/3LWDBJVeX7MD9dCgNZzqdWp
FU5VTMtGEbn7Zqo43u4ztCOI6MQorygtUDrac/bYBTgMhUNizB/D2ObH9nCtPpjQHBZvgswjWc5F
AKxt4V6if6Bcv2h/3HoQ48pOXZbSp3NwnKjOgL7DHXcF3rsYaZi/AIIOl7F6bLcrTkzaUaS0iHZc
+1HYEj1GeETG1236uaM0FkItk1YRpDYAIZjyJgyJZNaLY+TNG97DC4gm0O5SJjDOf0mU7Ty4QrLa
08ZHVjMPzZOs090cmbmRYNuepzV+TAMdKj3DdNF0alQJRLnhVqSp14uocLz9qTi1xCPrrFqqixZA
69aF0Z8Wc/OGOiItnWAb3QxQKg+Rz2m+GzcV+hYbC7YThYBkG84zhNHObgKzNsG2nwhtsvFwLiRJ
uII8TKz+j+aRBWkLzUamGfpt9MnWp+c0p4DGo3nc8OKPRkWGuqIYCZrW6PKLWYg7vFwC27gRUe7Y
40Efhs88W/R+rsdrtIoD+MhYrpDLMFGh4op8PjQ6JJCSXKVM1Lx3v4ZMueKI0JgI6iF4Yj8ki/eJ
vsVn1ecsxzOgBC/FE3mt/vSKz8zkkshtA5coCqbmx8Y90NcSjuLBGhulW7/WOs4FmyFlCOWulziu
+U2H2J7UJhxOtLrvrcwJCivywGx8vGdlp4DS5EEhTdytrwv7JN71UrcBPwVZgXVEGKi7vE3XtZxk
vhBvXS4nphoeoU10df2OwGacooxCdis3QokZqc4YGN/Ia2/IBGqojylPKqIsJt1ILfIYk8ieeTgZ
ZtnOduh6r7GYAW47lR9vz+R73J771LlVZAxg2R0aYmGs6/jFYCmNb6KbSMqKCPi0BJLekVt7oPLx
6AXwK8nf9Zkin9v4GirNNkuSQt8sdhsiimxlwTBTuEg+C2iw/i2lqNLZVKqwO6GQdpRGlZVN9YJC
70cQvtuzTr2aXQqDxvm1FJxvyf7ifyhwncUe19UAzmQYQkZA1TEUkrSTg61sHu9yZ+7Wk4E9bRzv
FeR4HVOR5qf396EwN8K8t38S4GDnJZswaBz4dwq/WLKh2F1SIhslF6r3EN+k81gEACx88NC//kmi
8oExkCkeEGi1DhNd4sXfjU39nj1PGPePGr5SuXy/8I3zeMYS+xSAwR+h6ne994epCeFXJnxuqk4G
/Ha/qKxeo+lzt6sX5moAKyi3Wte8+VxxZvD2/Nfh3cZPdH6dpNe+ZOcR7vi36xr/jPY+YZAaW/A/
vc1onUDas4jAo8q/zIkll3Ch75ZbVmBq8jH8BCTqRBtrKxB2sRWhN7VGTswwUiJDz6p3Jlg1WlSe
CyWQXWJr69IVu1Z0kV+ySoTvNoMI9q2D2mwPGST9t6ZB6Lk410OI6hh5cRSQfYCBlc6qJn56mMgN
1yZJsI3tEEv22LFLtPtfwQ2qEiaeorswN3UDdJ80jK5nZf6g9OeMW2s2l+XuXmIOTyYFuN3eSxL2
q+o1K89owmIqCA0aQXijXuK7ciSm/hGYakR+hsA3rK7j7os0S1eR6JZnqmF+oY2Dfq+teCDtxpEG
LyWLqcbougIl2sMQy8XlSH/lsaGVq/yZ6Pj6psL0JnfhKHk3k//axs7MKbiOUzGZViGwzvdwiyi0
sRd6QJWR0syfyBkGaBixRMFcJalLC3/TWd1T5xZPHcqQtF01SKWbx9mjLB8mttRlf2OEKQdQKrLv
D88+gbRM7sNj7LBcRCiN/fYlqwZC3doRLcMGwvQDDqKfY+/h7VxhRMrx2kamPlOU7ZOhviNp+AXQ
Rq4d6x4iAiLVYbs1nm06cdr3dwRrd7vpSCKoyxx/7A1bM5IAFcXgUcltmozKKuibwtE3y4djnooq
Uvp7N6JWmpIX6YcymULlWxwwXh6/A6DPJaQqSkcadC5O5Do3SSk6S9LBLc2WCsiJD2Xj0WFaX9y8
b6fRmVnZWdOCEnfItnFuKVh1/xuU/3xk7YpkkR90v8BY6mRPQy+XrnJMFc8SqjoKOC+vd+t3b+Su
KUvNYT8Au1kAhRy6rAl62MSxMIbWELW79qZE+MObbXDvGnkUK5UcqQsgYWg0+fwFJGP0xhrac74I
u9f6MmGUY3RpcFmCaFyvL5M+d/qPQxhlD3FdU9U/8GEAmjViu7+tQivJBUe+qXX4fLDZbaRg9rSV
MYrwAjWIdnNogrWyqck+4rRXY9BMO8df7Q/nCTcqUJVPV4VzK6RfLHvuzTTxtDHslv4608hX2W7m
8+O93f7q+iXaEpcMqG5hT2e+KSRqnQ2y+snG7q799822WfZ5PCuWTSQ66nOxc/PbEbSDt3kH6kXT
WPWRifK/Gc6OOAxAfpYmC4aWMrjYPok3oGWJH1HJ5v6rD/L+3i9q6wZyrtyAmN4h85ASmBfggZ/M
v656Tx1EZxDSIW1VRaPa5Jhu5GTIb9+PdDkLcS049hxEm5P022iBiAXLc4HmR9AVuhqnJpN0kT4i
YX/V09u7GyEToCoDlATW/Yt1C2+dah0C4/+vlvahhPBI/Ree806MugzdNEtQrOcoVxtAHzl8AN68
MQceAMkgchRhUb86+naAkFqqIBiy46xRRS3i0NT5+7peh6RbbRWl3eTDvIMCg6+7O5bwVr7B7LsP
g21JGJ/EteD/nxCh9igNDNcWiqedgwyM28SUsow8YmQCwbB4f41dFKL+Vb0VpVfjUiI1OVyz35MN
JL70o3fmkP9VUIxvA+jO9t4jEnpydbWMhFSh5elT1s7cGC9hTpnfr77tT2hlUUYkRqDh0ILTyPT9
9P8ngiQSXtpuoKztKoicQYfMJ9wJRYUD4+395ULRmIZmGFVNcw619iAoKpo50Gm+QqOknwRabqJR
UgKOuprYqGKLdcTCl396DpPXQAYX8A03H3v5Eap2HWG6imL0BFiQ+UrN4nJmFJQKX6AcXH5foqQR
O63WDVfXDsbquK8mkr0gSsyxz35k5pc+C87sBgp5/Cr+78wE40SyV+zWBOw9ZxqakA0ZRx01ktFC
uMuapidyz5Tq+FjMTJf7e6VS5hZmrUlhA5dtFZOVIbBz9NHbP5zSB3otI5FTyseVTQwVLd9ZQB80
FYiAgYcO5jlt7/QmNYwbFIhtBbPlqa8vcx6BIBuSyz79WYYv1mEmQi1lBRy4GCrlUv5FA7vJn3TO
5GtSWZfpMjGtGBo9upnGcKrTmuhodwWd3GyHZH+Ss0IwybvyYchlHOKZ4nKVXDfHFioIk0DwrAxE
kt1yO6BRlXJ0RVImO1PL80o219ziZ470M8U4rxrLDn8pqTOCO5AZCt8x0ihZeooRklTKKKGZ+NdC
8tIB9aggpVtoRh/1R4+ch/Eqyuyoyzzl05zfkruZJEpzABb7W5l//3iKsY8lIdPQKMX2E6Ytg+BX
Bxsj/SRQWwpkkf3xE/hOtt/2tVtBMDsiGbZFmGPMxEA1V98Ybr/sqPZrALvWUa88OTmwmFduZtlz
AAtqzgClWzElo8eCFAOJbtyWpLlQLQmTv2M/3lU7L8SfciNqm5cTgp+U471MqG+9EV9mhGi1KGIC
ab45+7F+7TR+o4T33Svy/AKkmNMyB9Z7yps93+9pes8TufIupb4NycpoUJYAb3DUce/5Bf6LFUJu
G2wu38T5LjUdLJoFa14UFtnDHsUXEhRO4pCG2FG1k6IppF53AALnxXOZ8SymsiuQ/GN02O5B+T5h
GXEWsmQy6hwEENoqJI5XUp1V29lGhVitPoNlsdSsm0y1EQiKUbXEqoZJM4IlGeJlrCdTW/FG73j/
36vM2DqT90XB16NfadWjkQapNdC3fQ1oK0+g2rzNb4h9gFN0rNl+/3UVP9Vu4gIKJmg/Cv2BhUwX
83//0JhWAzLXmfCcWHM2Ul1jI9xkwucYX+IcU5WmkhutlIpQNLtdI/h4l2XRqJT+ZpOl2K26WLOD
y60LDn0Am7tQygTxW6XNBSATWe7zRmaO1LAO752IUed6JuRRvlLXNSeMACbRhwIq2crMWyDIdSJx
ehMlliu6Jdlc5OVmFxr3MMJVLlaawoJb4UPwgDTHSn3MGuq8JC+76PQNmwDEjETi/IIt+dhk1crq
V67eT6EwSYhjsz2lGeUN4Elq/RCLrJx7f0X05Y2h2XGVeOe/gEF5gFZF5cQpGFhaOlLhDHnDl1OT
jdS9y1AoV0yxkhq1gd9VhAmYHV9SiJ3OwE/0mU9pGWpGDP0y36otYeSdWmWt9RbvFtoe6Zp/ZP2C
U03H6lS5cZIWpxEGBp/tP1d0ucjj05FBq3dl9Zj5KPxb5o8h3awto1nX0NjKKjFX5vLRIaPc/Mda
JOs304Ln1WrXcHQYv/QfODT5cri45Wjo/m67UUlIvdrBzET9oDFrbT8lM+bjDoX7k9Lo2PSYvUom
MgPibY2oMn8yx3WGt4DJfGVf0SCyptXaduZbun9Flm8Kt5+oOivdPWjOTd7i1lEhVlAubfoixo6T
Xy9kb8Pa2SfthEj5NpzWEQy5yIw0lZoH36D/KYrX3zUIYi6HOQfTBY3Tzw5L/Y91uSSUKGp7M0vr
Ly0XHLh4PWoxHOXdlLjcny6QZtNE2BOCtT3QtQWmzW/ntpMorNDqs0dq+Yzdwbe9zYDKcWqsZ40B
4lF4xwxjPRnXC38zKzUAk2AJL+81s2vQsxm/2QayMKTQ0dArjYgNl2YC98t1ZpVU9y+JQwAKTyRN
IhANhtgGy75o65UqEL8SDdmnhpEIndIH+wlJF4b4weoX2ljbT//f8N8dbqekzuf/t+NufPq/Ok22
ZQTNw84ZJxbj5OgV1TiQIeeDFm+jvgA86ckdkl59V+tKcCZqq1CAO0fwU7PXwNikfPHambJktw2J
J1T8qFDGGeK6DKt1uxhc7ks5QzUoJFSWNpR+yrI6Va/t1W7+c49RImO5vqirZA4PyheV8oMMiIqJ
t13O+xBBtzPKFlW4kp9o2yPFVLsXhfFq2aPC8pfLWBUqpTesAPraXL4iS1nJWXzjv++g8SY8h7QU
kxVpWb6HyQ7dUJuYCzYXcy+/UfgoacuexfKqDT97j7OCgoB+jgf35Eh/wOKpz+1OE00Vks+w5D1m
lZEG4w/NX94bVT1gdpxTBploDExR0Nbe3qUC93RKefKVcnQMHnY6ivnEAOcAlLLo7mzanUqfWbcK
MgMtSfdKUodQtyPE4Dqm7/UTsvnugwce3MVmr8Fuzx2cPCDdZF2FgjT7w4Hr1zE2MQ5CCDwJJ9K4
X5wbQfByOV+p5HV4oCBLnoTR9LtH1nsMGtYbwIKD2/hxOSDJcT3SPr501IAlYtrzFzdjVUcce9OM
u496iLEt+5rdGVyzhycc69epkfsuTScXF3RKdFkBxluEfqcqWhqYk/mGul+lxeApqzR2xPFjdYvF
LO1edMo3j9pUQD7ouBFW+EgKL/2NFTpEm+5BMGt3K04BFTYqj8w1S04L0PQlbo3tQrJEwRFvC5NR
l31gmN89UAEN/vBrJcqx3lEMo2hAD8XRtc/nUvj2AbXJOjJTEZ1tvITpGdRqV/kBsrSr0bmIF7If
qtmPC3OYUvf3Nassa6D86cBGGspytwNQbY81zO52cJNg3Cj2t4LG3ZdGnCoHc3PornabrS90SZ4E
Etf/KtLhpMtHCLnPdDhxKm3e0lNLEg774YB4gLp5n6BIuFfK1Zf0zGY63l+6hybMx1gHG97IOy9T
qKATjENXr09OT/sat4mxSSikwNilh3wQPIfEpbni+1BxAsyNtzyRQghGQzAipLa5VVGDBzeRmnF0
sMWUkFNXEC5NtuCw+jXM7n2hBwS0yVb0PHv5Lb+2a2P0P5S5oQYcsKI7WDdIBrF3ibCIiKpmmwzz
hn3wIgHSXsxa9uMFIoyH3vYCbh/LXUV0tpkNX9UD8NApXQhUny4I7zklx2583vkS6/x4PDH5eUzQ
VC5rPhximug2vpTcDxpTQnplokF2+1eBZxvXol6ZIjR1FgEKeq+h7SVYxXkuemB46MfAdgjKZyiO
NKb81qNV1JhEaMh/ylHKKXg4LnFYEC66a7EPXIPjwmXy7jNnCCO6BJKFRGP8BbgADFIVuLeKQbR+
yaMkgyeqPMYmJvc5QFXvklAidqD/84t2XxCjUYCSAczupkvo/K0a01s75BTvZhab/fCm8uu5SvFo
kjq+r3I6pSBdykqVBX9xp6nYrf6Fqv0Yb+WFywuwDayvEGmK5lzI+dAicPQ0gZL66Kwr8SpvBW7s
+uTBNFwh/bfuuajuawIqNxH6zVtb314hoBWBy5O21+g4LkKpjgsM/iBbrwegAZDUBrr9U4odQ9SL
xL+IJMzkBB7NujqxtyyteVsxOruJ9tGFZbK/an5NN2J3LIhWcPS8PEDjMInyRjpPg8fEY1+FfwN+
oQuvWbt86TxCo7n/Smh/sqaAugtFMfAgkEhBr8HvNfgH0rOY/lPQdKIYgf1Cg5PyCzSDKR1UmB/i
oTg47eCiaoA3ScmUTDJqsWFEDkY0zvV3GvBpJ6kEVymre/fBpX3TlMJRkZBAhmxhxTBiHLZhOfv0
rLeLtM/RUWcc1DO+k+MOQM3ji6EqnEW+5rTJqqnbAINIWaZm0Dp0jXdzxiy5yCbygwX3bt4FLnlZ
YWyqPTkwhtfGfNBtf45k7CQ2v8Hq44zCQ4f7xPMj79Cz6KRQx4E2jOmwZPmcksf7fPIESrubYV+n
r+bVGnxQAH3hd2sYljDmkg2a0okYk+aB1OjHzu78PizPj9nLZ35J1YRWcog1QbqXfedzA1oDR7fU
pRPGHEUNMtOP5ObkZq4pvbcgttME1s8Rc5CKKyzX1h0+2D7lc2m+rVuKX9rcioeKXDJbQnltBYDt
oVEcwMf4Vp7TqiMPwUkkJeod3s3GzGXa1HzmRI8r2Wa6WAc+WvJ6p8L5IO5jnfEk7i+/miUoC64u
I1tA+T/Kcy6Z7wpC8sRTpyxddWUtiS0nFdsdCSOCRYjN3lgIEODN24JqjQrLYHAquqIfo6kNRMx8
D7RL/4maaWbvWY1ZFJmbrrUxGDL1TnViJjx8fQad7kLp92c5LC1K8W+Cwv1ggEONkiz/BOgVrj4U
bJNE+DPPRFSk3I3VJ0f3/+KNuQ7yZavMy4uyCHGEOY8qdX1keEVjWCz3xnNs2FZJSZ9vYbkzYZPw
aEhAeuTCVA/9494GcpT7OyZvzZ0+Y88rzxCZdZmq6Tb3CCo2RFze9JHWx6h+RM8NjY16J9j15R7d
PQ6hyKGmW8tRdYxsGPquJYGeSTkLie2xtjxqlV9ynrjKUVz0KZ6QRR/4d9n8y3Ffig6frmiHgSAT
jQ+iewDf2U0fXRIqV3ZaPQrL89Q3OsCHTli5m+JTUfmYDLNKm8mkOKFHOGakwiNX1LwHrsTFXzHd
zUIIsbPc4CSYbd1STrt71nPWaQKmTOUCUM21aBTBE6Y+rIB8aRIOGvG0Yrq8481/Y3NrSaqJuR8F
f2z93wzNbryTeJ7x5XLOqOJmOdZjYnSNrqOcvy+ZQE2l74xvAb9JC7mAphepgF7UFwvvQYd+/5K4
KJ/eY05Nl6L412IAqCImdiyolfSSTVpyG1ylW7tPu1vARRr7fWCdrWy8br9lYV1otKe/Rx05qGls
J+aLZFiBauHYVIgpI/OXDj5Uj7UmrdBATY6f6HvDNJLablscw34YSVZ0NzgnUFTCKVUwgaktVtvB
962bTI9YitB3ghlyd+Q4mY2n6Eo3hkXYtfmIFFW8hjKxSngNW4Cgk+AyuP3qi6MwreefIdNuTB70
ihXu5OFZJPlgfL8OrRf92iXP7CE7fVDgqDixNRALdvEWETQKeP6CYJv5uuH3XgWvf7Q1TY47xy43
+TNmTmJaMMB+RUqonQr+I4NCq8PLArS7voNp+oDoADcTSk7DCsa68BErBnb9aH3A4zQklH0cwkAa
FSIbsiogtoge5Xgu3akLwAHM5zCSbOD3yIC5B8zImd1rZulPC0WJqFvJHQRa3s9hkozCUlvUP0K9
twO3MyTAh5G7LmXPLWiHVeOtd07d6x1qFX7DXfRMo3evhz8jS1C7QTwTItp2dWTIePRCCd9+erSF
An5xOOMhLfgMc6HpRaU4R1O+lzunoLmg2EDw6SKAadJVVxqdRr6WA44unIEjAi+Ha1H9wWukdgNl
bN4q68xPcgm/RoYPW/VAPJhejTm7/eMpi9ja4EMW8B6tGdMvRP8U0kyQKKUxxJjyKz2dPGHhWlCp
4CjzWQzv/Z+ZeCWr4OcpacgMS1GqM9ts24dXlz7E6++fj1Z5ugkBDVeVPvdMq9ON5CvCP1rzvOI1
JqSVexBowKhQ6DRD7B9Lybr3SOtiMxcuiWm/Mi9zz1HAem4cDSePU+oeqIJATLTYcCihPdsEzd6e
tS3/A9VB2sfEaQlr2TMXZL5GiBeZ5O654gbVsV7FXvj8QNdjdALj6TTwZBVECbOuBi1v5vUZ2wEQ
SHlnP4JVWVwI4/tJV1SRK0J93KwMf+Y9DJHUGS/zho8o968gBgzIOR0HzEc3LI+uM9/KgRRJjbAd
B4qwpVy5dXc+Je2T0W27IaH6drXn5EACclRR4WK0foyDscaaSCv20hKB6yqTeB8smKPe9vekMlCe
TjwzjkAwV5oPX9gy+OT7j0oNJlZf1huAwLpyx1cW6HSOJggpWLcqHx4XoamVqMYsvDsS8fi1B9CF
tW8z0Y7lwzYKkxMmG3shTBKb8SEjtq/okYLvkHBVCoIeEp7HmTI2z3WohBjj5JnhFGezkpnnm4j4
zsp8JC5KqNklo2ofZg0cYNk0nEKlNWNWGMYNMSAetQNiPhV+Unk6F5BoPj7pMIN6bK4vj4UXEmId
p+hHOu/50PgnEmnVYwmJKhrHPNMeCq23Y9mMcOYEDENsbBRd3SCNg5AW4elz2PPgOnpmmMYIxLAQ
Fto2MtsXZZwn7jcxD0enyxxM0VuAe3J/g13bCO5kAVJ2tLFSryUK8G9ogk8ZuQUz/JfPt7lFSuzM
jF2h2O1M2nvCGK0YJzQv0g0zaZMnc/PiqVEYfbW8D7TmE7lDzz0BZKvG/AN7eIHJVzsW1w1mjgKi
XX7V/ckNTmyCAcywz30uP12AmianDpwdY5JRRhiT/uQHAVTlCqEhMRi7Fs9D2OtoLU/4Rbaf9J2d
aWv/ikumg24NueURnMMsfryuM8gPhZWkUIq5o3ymJxCzDcU1PSbbfAXBMEJ1QDcVY8yBVwHWkGC/
O6NOsIc8i6Ld2ednBac94m0CCp/hcqziULF2tVB73rjaKF1Tg4+/zX/e1JsNtkDg/1d8u7IKujOi
AvjOmJXgZUmiTpVNMLFYnwMOKsz7+vPNdRaJd4CyNOVSwpMIJxwpELT7Jfij1NSaPUT1G+OWvbjd
PSRP2jgTdqxdIzZiJJoX0WxEnjP6VeVRr8xBHKusiFs0OVoBUVg6WV7MwExkoIMDx4hLd9eOYpAA
J6Kg+m5/clgTq080mjIEl0mp37chtuXlSSmrrDBO0qepzJWPVp+xtrHz0yG+GuuyunCPc9UPYIv9
chKoubOJxK1nPz14VIkEA286wsmEwVkmh/bGkL1lnvHE2ylGTlI6tHwrGNpPxYjvwnUgiHry/fil
swCwd5fM4V4/mA93/OO8oyrqm3F3KDW/bY8xtcYOZI2VsZEk0mBEl4iEVfslMNQ+89vtQZ0s5s8r
pwsK5mCra8k0DA7oUzbZMpG2P/Z6PGj111BeDCrsChLSuXE9gy3jxijBnYj5X0foS3zZ5MlgBRNT
bs70vF3kpCi46dbz39dh1drNqoYlVUC5aM2wi+x6WyMnH8gn8Ye0Q4KAVfTkO3cK3KjuycLe8siJ
/XZcjcR6cVV/YegLnZMGvUrOVr8I7hd16sv9KWweRbrOPuNuayzZ+sVpFEXMnrFcv2aMkpFjObRJ
x0IGoHBR+AP7h5AF7XKtdUkfMtz/f+lPzwG9mZj/+Hvil36QPMKpGXHse+f2b8HEE+uSEW8TmTno
DgzTkhzWu19KdT5JgMj6ABcoFHJQqHq7X4kD0xvoG7kQXpT3LlglJQAGfPggxwvv4eTZGb4/2zmw
GtNudYf/mN0PzS31AIbQoLOCI6jiSCazfj8iHt9waT1Or9HsESkYmrPCK/o2f/BGf8PwjaCesJf8
mF+0VcuWX4hhenxRzkPvRK7bQgjOYq33uVt7h6a1BH1gyM7jAkRHKwCpjJ4Xf4wFerAVlWNzNw7L
ey8+gs/j4fDMNcmarbhPoCr+TByADvsJend8lnyFlc/k872YwTWk8xrt7hv8vfhV84HxjKuW6FQZ
nAI0W3CwKZBHTF2VRZYGT2s7GwBD9I0E4CY+YdzmNrbuuxraxrOJu4MXqnKXBr7QkjDr9CQdUYTm
cx19pU+hp1Osk1zVeJTPytMMwaD9Xj824hMI0piWYDZPw4v9SxJVDAkjsvqFMaAGD921e5yJiQ8I
DYUX9AflgE5pjpWH/pw90TE9RsWlTfuyZrvY30djvhIO65Qy887MhqAxpdiqRSs9jY/1+DX1ltgd
hvQ5wSHTnszFjHNtC2GbUXzB255FtBLWYivlKTJCYA+VE8lPZUlRsExIXg4zVsZixthohev1uYwn
UbCvyZQsALPUddUZz2MriOyLn/UMTu01G3BjoZVqlA0G84ojENpx3ItMmDDYYMF7TS1JE8GacQft
R/pKffKXWBkzDnwVAu7uxGXeqYxPLHJmjipET/q0OD0dnEjs9KvY37t+2TA4BN8mOHNgJxpuPK3M
D9BtTM+oUdZl0cp7V9a1nO56tpF4unap4tTYOIDVdiXpdy/xvHa8YQ7eAPTfNZbC5D/JYzjdB2ul
s3KpbNs3xxFj7PeYPyxAiXSpbLJYWaPbBOp+zYX3Qs/w+DIkNXizZpfONz51051Doo3onxLYrf30
q7O28VuBjHTxa3yElU8qHBsGdfVdIUvmpPrQpygVWVF3e5E+NK7EFI7EePy9q7LGWzjbq1gT/+U2
6FloexHbfzw5FqfBBEmE0oRz/q4iZ+9uuZCcJRmVuEVusCgZQaLKyUDAsYUX/c5HhkjxapjccCb+
Id4UnIbGyn6iV6a+58SE3cZS+N3wwylj6OI6HQ5pWbfdVjXEw1q3StGyNHRfhqNmfGuqSu3PgYd1
TSwMKhiCkW9SiXebFK2f4P7P9aLa/EENd0Jx3skaPyXmwuoeggTptuxFDGTCquC8jDCiW+3J/2XR
DD+UG7M7Abcl0pRady11jDrRpxSfIsYNRZpHlI3hr8KbX8bl0zHMq5vEPjNEo9U9K5pVj/thjWvw
EfYwxe49OrahqH1y/pmzzHn9qpNLwAVTJ79b3li8ToJRcp2p+DPYLT1cd99wVvxvJ22mZi5lD3zh
q6qzJwVuTEtOlTdYsbmSexKDRA2KvNV8+P92+VWHNKgikxrHKIRks8Es4uLqffku/vjhB+o4MZ/Q
SZgkeuWZ6SNYLTfNdFfs+GUVFHPSJU6R3kgyiz/fI41QNMoEnKLFijIWWDR6RnnZfOTUZh4C4qm0
jShYhHa9uYhN4SYRgplPlbPwQ31SVJ7e/jv70+6iJai9DsaAMdniiH1qJO5VGgxO+3BSAKa0J+lE
bKvr+JOWZKtIp2sRUORYOb8g/97JCk9zS/jUCiMaEiQCS5CLFBUPKa+M5EBovijrQm5O+SLrbYhg
mWQR+gOgg/BSksZktAw1O2uLtsYOzzIKDDUDEy3Q5WeF/uI/HzBpt2rcrjWKzzc+OtQOmzP16CMK
Ra0iHKzWnrWJ7pCf/Zv64aYL4+Kyk4HqieNY3w5rYPqKwD5mgtMrsyyHzAooMVIRB/Xbm/W8kw0t
pFQtvwxxkBZt7K+jIenmnYaXrz/QD9A2oTHCqQHkGb6T3E0oB5Narv93Exb7zMu+nFT0lmhd2mvK
6PIOap0+z6+HmHJEANIGFh6L44XR7qRrtC0ia8HIR9RJ6Yl++1TcgtCLnJDt8b56eEpnXBh2d+cU
KpxeAaVOkGHhVJ1g2eWL4oydRU3WcrDnWr/SgXg/r4y02IAyPN4IK/Wqx+Hoh1HwxX9daoS8l6ix
B9XdCUVrgyz6UGG8Eh49RLo4th62bE50MGWpnzUcWN+pUyKxsZK5Fc8hkE5y6uI1VbNCWSO/afdv
6OWZjeYeBIkROHEW2Qiu297bg+Q7RmuXdBrgGuhkzKNFFLQHqj5dPPm0cDFcdoFJ8wRC8vJ+W0Bm
5BUsrhaDRnpO8vsnxkIib149iWHDdK46AVYxIwSljwttmL4KkbiX3YazDLbc7Bf9Iny4/u2H2RTw
K4HyX+irltzTA2khxkfw4oW8vzo/DvlG7g60w6X4rF19ofqv+98fY5c5yZgZI71bCPYnq//oEkyk
WkVSeIl3avZCZovFwr36DGxjku77wdlLFIgps54ZD3LOYXtFXMisc6aw9j6FNnyVsXcl04lH+8go
wVsq9iolihhV4VwtdUq4pBB1O4MKuS3vP5+51gWr915AEd5bQJ4pjef7JWiag3HcuFYkGp4eA7Qg
ThLvFPwwu0TY8VqlD4TZUMnxrwPHPZLjMmf/38ftYuj5OwssiKuf8SkvV5LrcUXxJhaHWKsD/xSd
BCyY3m/HpEh9Dkrg5mcrUSUkzQDb8l40RJKteAFoXkpHOpEuTII/iwhtxgNv0rx9JEVVVm9AbU2k
QEY5cEXg2GMlgQEFDYQBI+iBxn3EGfCUDw4bDhV6u3Q3GG5SleX/eS2YfCaZ1yZ62EOrn7i3Vw99
mXGXRZrXE3ava0eelS/OM71gIOTEZQC/dgEI4gkm2yHuO7tj8JJg4mKTFb08DbssaQayA+KT2Lpn
lp5DImq5WwiBBW0ctsYAOVzpMCrH4Zj5XdXVHxK2VWUtgXQ8v0lkUATx27fX0cAGV3hOL6kKwk6E
QQoLAqwOxoqa7xjphh5+IqjbudCPqBs2EmMBT6K3a0gR5WKcDMm4Gi/B6e6yJVbYE5cyP1rBQTFu
uDB59kIbtiHRWZmYYePZB6r328cYD06TdfT8w6xpsJBSiYH0DGFakgGSHJtpomoltquhnO2TivcF
Fw4baX5STH6etSgqJCsHWt8uFoLlqtJQyuU1tWTHYEgfsv6kDCplFU97J8ivJFY9noQA/YUwVzTG
jRjuWKlcpES4K3QLkDwdd/etmsAGkZJ2h/QRN2J34xZaKuAHQocTmhYSFrFZq7ylSmN1t4S3OJdY
1AzY41bGzZx+1rXwcuX2fitU0Rh3+FQ5Tau3q1zK5rqSvjmXZPjkWYJVxexn0mQXv0e9eKMEddKG
sU2J5y1mnCc7ylid7KjE9zBn2fhLuZzwcyZZs9NnL/6ZnLfVLvYNcpXwQFOookrSzRqEV2POVlUI
p3KTkWBmpiWE3M0MQ8rqOW06BTGgN/BV8foW34526TWSEyggim/ZL2rAzLDV2feo1fBmvaLmCW57
pItuA3qDgYHWRffXPwBjpcmv0fiNkvFY9p+WxRt782fchdB3T+R0GItMbjBLG/kA+N3B26Db0Ckp
UL1EYIg7YtQ6Uo39BtcQou+7hUPv3WxhJjjNuPUHVFMu5DdLOlAB4a/Hu9+/kAp2w5c2ybv2peXu
tmshuEG9j0n5yO0C6X/eCXSOOfIzvM3tFJxhAHjk4CXXcIqRLutLd4yqVr8vdmHSvvebOIJhrcCM
Ih9q1cbcLCRGx8dv3yeoLjV5l607LMkesOMUQ8InDpLECIPiF8Jyv9S/kV2DHZND4m7eqmi9XoAC
lJ+aAlzIMOC63+AGzC09WwoNsVC9fDT95ea6vtnAWwcNOfQhOSDHlGMlOYZTACKM4z3dzJNyT6h9
CKktrJ/PsdU7joCjpSJFGmYS6kfplvklMb+QF9a+2drlDW5BPqz4RVcpi1LJ7LTFstQoZbzfVF8e
PE7zipEu6CqYCRIPYOOumxjxz4wZAsLHbDxM5Pg0Ke6wAo6CQtw00yDMC02tSgKNlZNsoIa2CPtc
OKYh49rrhV+ETII0VAlepH1LyItp2pWRz5tF4OkgSGCiwAA4FwXWxAhImbZg+EoHJbfN9Pyw6L+k
a+1dDTa8iWgPRXgTOPDsQK7R/YYHDw4iBr8jPp16Dp1WYdWdestLDg88Lr4DaagFzYc2oOuWARwM
sPvFp4fJAK3k4i/MZ68NV9JRgjueH1XoIheDDXMmZwRJI6oqxGNGeBzlISkP/uOXAwqcoX2ssHfF
aaQlSMU3zNbQQ1RICCDIUumClhLOXzKn2iZmcSuqs5fVrpA+Mx5WbPi+FIF8bFTRXyts5H4nW9S6
pQLwMz9L4gRjw0wy23UzsdPdWi82nYW8Af6uGSuw8P/LTLw7+SNqkeh7fCJlQiXnC1MFFVkMn6yO
Sw317NBlZwmPm4HvsV1kR8D/5TiZqwEeikwlgXtybuWn6GOgV3aaVzROLK+IEVns4+TSenVPg+qg
zaH2WNpc7PK00GDGuMzbbgQnEopEsjr7YyAthXibOWcf50PsuETx1daEfnlu0gUlAJXFHXRwwDTH
C8D086FTpJaLV/X4hoYNJG/KGFkAZQ4p6HMdvKEWY0enlOAMZdcaVOf1jcN/QNyTRAXRGyp15+za
ht4gAku3HXbWDcEPCnTkDAbmdyeDNK1lNjIWzR2+yn8O3Q/zo6RTaDW/QZphrJYZF936Y8+/+ghd
qj14m7x5yYZ0FUnO+vjv4jClaxwo/WD8d6uKZjVvvbN3jMH+VAsJZYDGlOwkkhN0Conssk2r7ws0
oxGUWM4UTdVuhZpv10YKHBo+A5Z0wqNiK9bBahhAln7UyEJG2X3BcrRNfm7rk5eohThZ14ybqyo2
CIbF18/QS+vwcKIcpxdRzx1g8W7Eks6Z2N+I7lqoRXCQfRKY7m348pmFEP0odMjrHJ3yJB3AMsyD
qBcYqdAJEjuO70mEw6CKSUryfs6OlrHHqiGZeoMwrmp5H+VZK/hDptc/a0Nb00Ervtm0RvECxVXV
qavFSlwkIW514yEbno1Morb5kPlvPHYlAw5m/2JGJWIG4zJmb7MpWiv8eKoFIM2/4+nOLBtzf9uE
llsaipx8IRWd+8HxpDvZPzsJpjjYX3r/TqB0Xdf7hIqwnZvhaC5BWqSpfnBj2PleDNOXw0dc5Zzz
cvK57zOb9Hyry+3vCu/qWw7TJcXyOOaez/zW8Egkyia386LET0LUQDXkuzw6OOxG5hO2JcA5tqGr
U2jOku0zhOZq1XaQcXImS6ZVHeAFbj7m9tsoe/2ZrxsJK9UaWM9pTySxrL9QN1h2CJVIi6k8ATUa
6A3slY4geJsuemLabnQ1ImJCKB3BETRiT/sMBBOR3mogoLVIA3sDJAQKjgDarJLq5ERhV2DyPjVZ
Nf0ePDoTr183VoQxgK8TdAzDfeUGFn84x0iGF9Y7RaSk/DSB8xas0+ld4Cd9SJjbZdCcKKBhA8GL
dx8/WN5UUSyxTX1iq/HHJc6LmdDrgcwZiTytAqIVS9/eudGTtHuDnTkoRw0iRzLaeEyXEPqIM2GX
iwjgPVMNDJ2umrVotG54J4JdMdQ+Htdn64+p6u9HYWowc7rCGGtq6Z7t7RLj8FfeReQlJSuqppdm
YfPeGqcxNWW108QFak0lloQp6x4kAF51x7KUpNliPIP4jxqzI65Wvyd0ZeqmoFsNaDkoq4crfM5h
/TdFJH4tkG9tecZmqev16/WwGX/P8y/8e4qJzekIMSYpQeZZVcLGGrFdC1bWD8ZIR3mTqh2duPR4
c86rLwhI/5LFxEZD/jPnMzWBdkR1y7SWFVMx3s14oishSVfB5SUaD3qY0+rlYj5u9VoHOdNT3go5
AC4LmOzga/iG9a1YaCX+AynQENZzjoJwtEmv9pksEVBx5fWVmN8KHJqXTvEzLZSrZVaff8iiLgt5
Er9Sx14/fI9dp6t9Gr3ppJYzYmbAXxKnYieK8esh46cwMOZZ3C+mQ6gbGs6RB0gn+Twy5d4M5e1u
iZ907mrJ9PaAAVVXnRB5hglyjGSZWhurHvVfImcvbkc6WaP5i3GzptDxZtc5511VCbxB0NG02vL2
lzwftvyrTIbgN1+JJkenux8pKva00tm9Akatq+liSCpos8rUyhmbDaV4P4ZhxpUXetzdoX9cxAX2
XCwHCiHm40npxCBA0WSM7ic3cSPE68ANvQD7ZLSS+er850XVHcQCjid4Gat+5H4sawcccOL0318D
UII19w555wDZTggfcglKvkkgiatuIHPjB2WEBXG1lb0qeGs6uBUB8qDBD0pr95oqrjWz/qyoEwtk
IZh0klTePSGVrHAaaNCvjRu078pJSwXnxYhGz37WYDMWXC7xjJ0bxS2iUT9XzOwrAo/2EMP8T45G
QeClvCMXoPiykRQws/5v71wsjgG7JRL5y/L5OdCLF7XCUo9fIB3AKoiyJygtalFpI0kHB4wAi2YK
gKlPtjOsKmePYvuZOzwz5u4VDsR9blR5gI0A4TA9YRdWDJT1PefSFM7yZ61NLUJIbomnMM9e3oC7
l9aY1o2Qd5sApKqmZ48NU/0KPiV/jk0yhRqRdbcaR1bNaIcdSkbrix+MqVH8RdqFuS6aovDMcRMr
0JYghmyS0OJkCOMF8ibeO8CAtSk9ayL6KZVaTEfZn/2iR66w4hGE1aqLhZw/wPkkDuji7gtMhujI
+NBFAzvzrjQ6mP8sXLHWFq6pGqyyeUqDt9aGZlE2ACwRTCbv9GgsEcYxe9uMfrdMi3V7mVrzXtKR
g46iZbj/tZ568Nv4ZwF9lDF781tkhyxaskRM5Vkzl+ezGcL2PeeC5iHqD9JNg1R3Bo31tmj7mBv/
o4bJAiVc5iXLHQdZYZRePRUfdPUZI7NwmmY/X1KEwYerR1Ef0L3FdeXJ6wZY/EuStrsMj63MKlLW
GgerWS0A8BySwRk77SF6Mf3ZmK2/74Zm/4vBVv5hSDv8yZbDd52G7LTGsfbLHc8sc/UzQUnqOaL8
K7JXSbfOw3SVYoQw8/ZFtoaSAuPSJWxz+KSpDkuTr4BX3Tk+BcW6TKDW3q/xeHAXH+lKK+w6Y8WF
pnCb+JQP/R2+awP5XVmIFB2AgL5PMTk5tJtN7lsGYEJ+/uIMdofTNlQsuvVW/maEeqySEJfAOIbH
Hqv6xM/Aa/KWC3436yBblT/XF13NOwte3GvtbI8I2Ybga/RqZEe0SSe+7XhIMTnJjBgnb+OGxCQ5
0RtLtLQ31dOgpNuAlpnkf7EpXnMDj0Aasf1OxAmEij6lvEVv7sjG9yD6sU+bnuCFwcY+JMjzgySM
wnv5mLcsMcnwb99QONS6lWsmiK2cfU/62qw4vymqns/gLhdP5OYfd65HbpQYsZM1Hd2D7RSWV8HU
PEwrYQtqNMFGGoLN+gJcJ8A1R1q377L76MBmrkSiKIAR8IhOV6+t7WTdSJL1Tyuwu340kPsBzvFF
yDa184zB9w/XAhhzO7jOcWNPxZfva0Ut8kihpWTcYOuGimvf94uuNydRmVbNf32RmBXq/YxzQap/
dShzIIB45IRN/EmlhCMXL/SW/5MnM+IQhCH3fURGfSVkUKWCcs5L/Nkk+y3m1T7LN+jsRx2k+l7y
q1yK36BJRnJS8WnBamjXM5EoNcAyIQOZpKFEDWovpRrd3OuYbHVW7PBmXh00gPuTzH8lQeC7/n6N
acShm6C/OFPTflozGf2xA/TORbwgxgljKRad9D28xlwEmtLBuE0M/2p+1aIbKngckOuqXuWCTqvV
9/OV4yxdM24xDUTGHi4d1tX3UmkJJ4s5zz0GqCEurHb4WMXhSNQ9th4qgaXBzQWdL3gFzboEZY3g
vCpxWrp8Jyrt9YGEouhutaZCdEN/+62You53yzlbeuyIo0Uh8XK2O3ku8XD8RIebjktfQYWGsqUU
GycoU55mMw3Rw0Efsun6D6pRH9c3M9+0f6YDLBijS+79BLdMTT0TrlXaiBkh3rfqORCm8JiNBK0m
GZwjRi6I+hJeuD6SOUSotYJSrx1sgPznBeQfV4Wde42ISAdbu3JQ09O6MX8fOnbZDL6TdFOo+PC/
JXmPRVfq2pGT0f5maFuv64pQvpJp3apDKNjWbtAsGYKO3Zz5Esy5If5MRZWh4RIudlqfi7JrnH2r
0HYx0j/CpIIM57SsaJ0kKzxzgYog3lbsZopkmu9UV3ALBZWxeR8cYILV+WIgsTvX9BFlghIiuo7a
w3ZUqgDLkxgzOXqRqxX2MUqHYrywG4QR30pXJVCCXeSILaDZHojkjvzo1QGmc5It5n4oLN2fH3Ve
W/6O4Sg//+4IVNOsZPpGJFGyOIQzBhPFgzBy+kuzzCaM7GQjF4bVf4rtKsY6P9lJjANyh1AHz3zM
FFddivp86rGDkhCUHECPwJfIXQQUd0/BHAzggI2ZmAFk1UNWW8fAq46xsR87yqIElvY9FUai7TVC
kzJM439Pqf5z6qXmgifiXJvYzlirNqhMSjVhth92TrfWo42SbeHn4lSCGM0zCRIQCOcAY00eqfFK
h9UZu7XcTYd9/amAtGJ6CWTNrBa7OXYhspw3C/gJNvAul94fCeA/+1eptJbeaQt3L9JtAP1dhph0
8hlQfwdiU5Gnm6h2rf53WlnStcQsc3IxbJblblxf1hwn2IVB63HKTGVWL1JyQCwA0W8bUoWMqbmu
phQbsuMnp/AeCnD59XXL06a7pfHcY8k/Ckz6lv5TzEsNDfah5fdiRVi27ILLQHFzw3dbKEAKz1C/
Rs53oNX5+bGQAnvxWzOMy7lXTZSrPnBVdMU/EQqvBmN9fZjU/OzFSCwyHEsXgJJgEv/Nwg79PLd4
JP6LbWzDsAWbTaJx9qcbQh0SrMNPf+jzVcuJRTYFyP5hUehUPxCEa1jd4ZHVH2YtH5miFbctAwzT
Ots8DHPlrkTFCXAp29yU8XjzEbxzDWyaEHn4ZPuoWs4VGaM9EXiMNJSpukNNVinGWUFlOu5n0oti
k4kYI9uXIiGW+qi2T+xZmKvK1rUejX08lk2YVpwfZGJEl8+TERk66y0A3HweTnEZtr31cHAdrTPQ
UkvZFYibNh6xt/LXsGN91q70vGbFeVWxgGdvyDFF0OBn6Mf5G0pZsIudcikDUkGLoEL+nRNYuzJk
zdKDnnRSdZN6zEU77/lGfVCyxEy5jEebypTMvzRrF2cDswAOOiAGj2JP7M3qo4fPXh2ULluRPMte
ySyvyFoVfI59hkpywO8fbnIVs4++T/99p66DuFjxRQiIZcNoQ3Mjm/36QdODTJXvigwy/JkuJTHo
BYt2ABXJ9rUcsMQTsMjpdxyQeD5ost5ijGtWinjAe+AlepOmaCFDahzm/Vv3VvQV8e4Z8tr779yE
RJZu3YfRuppPZnl2kge+wAKdVX1Sy1fEh2xnfTExSzzHEAcLKw43LRXv/w+13codHuneZY1a0rHI
/ns++Sxum8kVw8FQbos6D9p9aJzhrnxRPdtWRb+X+OXAlTW48zEDwORa5142JtGKAOCyuZeWj6fQ
SJNbdMNga/sVC5oEA9qg3n1RujP6UneFwfQEbKKWixdh0SCKwMIL2q7f63AJFlPYiNDaodfElkx/
agBjzBGFBcn6F8ddzowcEekczWYQku/YxI8TxvEEd5Nyg5gI6c0RqyN4TY7KANswtzIvf8rDFoPu
zZ11nMivlVB9+fRsbuVhYTWq3FM0LHhzEYwrpx57jtQX/fIhpILOA9TWvk00X2z95mMrSZtP+TtW
IAXCST5yx2OXihmR+kpf4WR6uGIdIEe90bFOhBwEYQix/gUnC/VzTuaP1ZGKGiW/epErTpM2WsAM
qF5fZGwXnVqZFQ/clrLKcye8PGhT8YsY0orE9Fxtyon6OJ9A2TV2fwK5zF3PUVpJpo9na7JM3hSd
tsxp+N1eUpr4zZQdYLMo0Ibd6sN+qzmP7S8Hh0t/Mh6U4IhLcV0mup9VA46oarvU/EmZOpSB01bo
l/iDibQd+pjVr25kAYn+tO98F+Tj0JfwuxehJjkILPc9RWBzr3TgFJsOFNShzN7Z+IWnP4YhKUdm
MUbx0MtTpzHZ0BTKcPZPVvXYw8sDft0sHGPqrmNbplBHaQQ/FwlEYRRTT8FaZCiQPv/sXU6XmLgB
/H2PPgT8yfUCha10o2g55HQVDU75Zpu0n+aoorl5RFJq3H21BoX8LAcVLjSsiMymmM+SQa+hPPcE
hWKybBMAsfigGLJVlgiZRpk0t0Tej5iP5fCIa6Q2bXl2o67lYeYU/gGJDVMpYRH7/HZkEyu04n3b
KP0JJZ2iAr92H74dmuPvwHk8wI4lqDybmu2iN/634boYjrXdDJahVu3F49mMVXgBP8Pj9LleUGMF
SclDvmuSuw1nTHUPCgXtK9NTuHgbuhtfCqDl9QPT1VYDxOrw6hHSLLKoioQFByGitpFsc8kFhyq9
IPxmZUGka+7qy5etkeP4WxB7ce+vKlGL6eZg/zf7igjH+srBG2RurqgWWaPnM+1NeJ+F+bfta+aK
ARkOyeXbZRhz4yLe0MJ2Gje9y+c7D7jAFfoSoCmPvXRRsWcQb2AvlO0oXcUS7gZWujqt82oeS7IK
4D7SiSMRx+8FZOfU/atZAQ6/B1OD1dTA69sBmdAPj6ZlIylwX85qvuDgu5nHN8ENPGLb2UbE6cvB
0BuFAMtrNTyLZ9hhaf924uD5Vk8HMoDJLFWqz5+N79XiEk9G+loC5rGGz4/eXmQPpwpDkkerBmCJ
Xb9qTgWjoF6NwL9twqZs9RgiJyQKL19GW/E4xUdNJfsRrx1+/ckKEvbwLEBmMM0TNrvQKG4Ak9xa
R3Zr9Dt4YAaMV2wYeyiCcu28/sCT9e6kJ1DOwQS3mqsf5RA4tSPoMdyitloJ22CpS8Gu7vd3RuyB
lXK42Hv8x4LpvJYO5fR9y7mYLUudH7vtTmExLa5W5aEWB/3TURU6tQroi3MrWRK+v1T8i5ojyS4t
JghdQY5R1860UkDT5cHgB+ZStavGPTsYN81gyYGiiKs4XdtUXj78O8X+xmo7LkoLeJsVvuJkPXaA
E0pJmOXH2AI+N7jent6RcIIyHHVTQy+pN16c8h14kk7uj+XeyIJSsILWkaDij8rUDE0qxTE5ZuOV
NlII9jGmxsH0tem8wHV4FoxLzEsxGdyxKaXWQQbEnNyGvNtMpvOECAWQVP6NGMzlIHGfzm0amTij
f2Iy4hJ9Nh91t/j+YkPKEYP3VFFsV2rstcedXTTRgHt2/p8wMc4JtqT/FWE8pX5j+MurHEX7teEM
wsvGLkVmOiiPeEmPQ+OkDMTvcML0JD40F6ISp7nJcP62i7rilFMph17XLQxPs/a5MrWXlo2pJ9Nc
g/HN/LUPpwQLtEJjLAjiMZzIZNfuK+RyyyexzmCcd8SRVYtCsD86bb3sslOuCk5cfp1VMwGPieIp
5N1NUodXJysRrK5/x2Pchbm+xfyG0NlMYNggcbetmVHqqVEYuJkpA6doUe3+H4rhz3DpOWop2zwJ
eAk1IJ4WV8kE4KlEEhwiAdIZZfo8TZmDfSRL/+b7W+Q7iCbwgUSmWUtvmcE9Uq5D36ZlUi+qUT8Q
c77kPHI8ny3V/xVh76g18e5jPOBYA6PdCXO4EEmpL9ymaPoKnMD2XSdhNXR9QNv9stPgBtkAk8TN
7fzAW30OXE8sVspCvPJcDEcCaxZoAWExmbpkoC9UoLmooMKPYhbeR1ZdKopc27zSkh1Aizyjv7hs
978S8rVVIhYeO6Eyu8+He6kHLLh+gbfwv5vuIYRwuaxZkvw/247w/bL6WCTPik7P0zxAsmOXOiNb
hAFOJaT56uamz1u1TRdAqBMD1iRSIt7YQd0p71SxUgq7H3ZJP4zCOnd30jkzkoyDzs+yrNT7wfwZ
fcXZJDFqojpQEjVqR1ppSqGxNmLC9mUE2vDNzhYC3z4Zrp0bBBE2xjr+/99Q+wd3xtYniP2Sm/HD
pV4GfWJt8Tw+QbR9b+qf9WjccwPstozahiQDfP4gcHMGE5WAf5DtQU6QAkeNQfeeaJchcS6CZJjS
mKVwRi2qqpa+EvVCUqg1eWh3ieMD1JJ3bE1ItRRdJsa3/vQ91i+ShJN8WTM0MR2A+4hyXPsjtABL
0NSjvJtqa9R1pIJOSvC9opCZXLYbWntkUaKT7llbi5Ewxvaz/B4Tntkt+V70ZKbMnni/ZF3H9GHQ
Q5SKYGSjhddnBN1TlrOJkbkAN24UFIVoSiReI3QBWMOJOiLGAzwkrmOac4J0AEplgsHEDyAAW7BS
5jX7/p8bsHSCyusgGJKlypEG047J7WQ8YT9F1ROMXEopJmjHOaucy25uf1WshBt8JlYEktzYmbjf
VFP66ezHQbKRZkmsYFBykczVlRFjrVq46YmvDBKwmZLIU3GBYzx88da/rJg4W7jpKHwzZ1ARdZm0
Ieh5OhB0QA9J7Z97m7I4O3NQLpdQGunHel7J8I4WjiJ4NDpfPDIxSzrFvK4dvRRn3A+CJSgbBKP3
PUWZLMFi+9YEQf0RDyXF9wMrDad/2bGEE0MgVFChywoC0L5kNqr5JK2MXHvNhHXIZ3rg6ePHL0zq
Di8prs+fXuxN0RbQ3S5Y8CxfvYy623+PpA4ltr1fkpY9Y507KR97H5KUitZWsEKpY8Dp/CoIsJAn
3vbkd/eBbh4i7OGjBsJRkcK3GkykCRN1e8pu/mHvbaByerpkdgwWoqV8SCmDVlvSPyGPIG0tyxrd
xURtUaOyHdiAEQw981GhNW6MZny9AeZlq8v3ICjVbWi8HXXHAO+GJap9v3AHbV2MzIB7R2PynJHm
YKaKJ+WWJm80PJPDAqKXWKDsMl7Bawiqs3s4kcjKeVj6w6GH4UQuOCdj7XjwAgOGQTSbTqKWhCRw
N8aaZW5qEOYTtVfX42Nr9gARu4kHjYZbGqAuylCUadPeCs8YhpUIhEGyXWfS6Ilc/foGgxV8KNSz
Ticf2anRyyQeREhptYfCM6/6SU3iUZKG8Eo0M7ftFiOc/CBXTfLDZwjsIPuil/PfGDba/1b8M+2G
zfbA2uJpnwffdmuzdpZ1/E1ykS+MLVEj59HYlME62VkvqQmY3Pp4EMxma9vXZyRe5+zywObn55T8
D13rwH4AWeWDdnyqglVtjUfsOBoXCcf2msDV/efc+T3PjnvxPfFUM5IDLPsC/+LnttKjHUtaO8K9
FHiQfPrUK/Pd2BwgX91vOcXowDABkF2XKDOumXgV8T6EJTEQTZFgISgjaDOaZMF19lf2S3mIDgJc
YL9igTQVIs6B9Ytzb6iiJh+wCI/BJMluaEfOzyjRbwdD4VayAIZ3oOHhf+pemlah2M98wysBddaJ
denJflOjFn3Hhuo9m3t+dOkxjSObZNndLFg9IML7aYYBijrOXN4XzMUimB6UJM3ChojNhHuSfxQq
JF5WJBC8A5VWNDbctcjuRJJ2Pd8MPxT0eoYjNSPgalSEj9INCX3USS+4qSx6mh21Rj76WUYgIvq7
aYct15Z8fph8ZQ8DKO/+t0orSrC6tkO0aUOHJk04nHC/K6d2xsvTxLDpIqmLthysgh7B3AbTXFF1
APcWPJAOWKsGAS7a45YlTxCnnHhaTwWpfKsewbqPmTezBLyoPurSk32BA6fv9PQC78mbgPOnttwc
1iEOQZ/yGCCWj/xBIpvXg4leVmYrAHkLbZaLXEOwgh1F9UOBXc1h14G9t5oanM9dIP8mhotAWHSV
5YHami5nfanXCJ3D4UxVAvCn9b8z0wWE7ezWKZ/FEpSnlToDAcoDfwIJynmXxiliz8SwuHiAzFpk
mCb5mseMMjAlXoaFVrNdVtLvU5aFPnFP1FX0ncUTgzgnjcEV8mZRZ4PYl7HPAJoWdCsu4F+8kQ5p
1kVr+qGDvOqoZWOHZryfXpm3odWteqDBC/ow+B7AknHb0Yn8JZ80/CV/necSHLuYB4dbv5yrJtKM
Qo8xrUTGs8WHCeTtlXf+u9E/3zBAvXz/gF8rTfjSyZeOOEzyOjo3/LLA16BBm9yWqxB8F44kPzlC
nVS011WjuqeikoDSbqlm89mK80DJccQYlkPoi3DfL5z8iypUdhMa4/xRUiI2+RpyiNny/XmdFtjb
LgQXqumhep3Sk5cVePOJ6zPELwqfFBzH7NSy27e0q5cIiNAfB3l05Lzp9Xay+lPVJPE0xGeiR5/q
YokZPo8aLKJiE9ZuacOtb4ka2Fb9FKTV3jg4UjTaWJi+fIobMd9P0X9xZ6Ivs6rMECdM5UMyXsSX
BFzVTg6AoyzIo0fSBe41+yCqe1fXdIcBtEGEBtNcHTuPX4EP4pkOTyj/F43qduDkg/KIsvBP5z5m
QhclvZ9xQBHkHnrBPJAwQSv4u9xCa0d5CyLzZ93hp4OEC9GXU8qNgb3AQBnj7IUdmKxdZLk6p/Hm
JlciPr/YB7MJ/A7tGzXlejcAx35Gln5F2Mc/LbXfBENPyY7OSk1O9Iw0MCnDXdmYyO+igbEFKqXO
M7hKDjcvC0x9pLDaiUqfozFmaQEGV5xV44hb8zk31SXdS93FGx4BMutwMEjq077odd3Pkbg2OLvj
3t2Iov+ngWsbwx1cQGu6kM1SBt4rqMpYfMMGh9TlHGOH2gAd8aY0uxTDoH7ESVuycMD6qrxme405
ySpup5m6Lflax+JQbb8An+mOgK0ld0PQaZP7RjPeEYTmIj16q7E63ajVEv57ENRDicur3VviKI32
tsFXrl6WlCRjqpNjv95h017YchDsqRyrnku9FJG77G+KMjZi5scV9SRtDMUPEvsfymKzLYrMpmaW
fwQYC0hR4Rd48PVUwPDMPJX/Q+iF/Oyqg8QX1S7IUWeEQmh1WnMOfn6I6hWInWzUIVsDmBrTlgA3
vgIAV9a7CyiFodxnp5We4e+LpX6cWC9zHjOt78dyh56Q9Hr/CpRyQ25/B09DZENXmhy23FWgexgy
mU4x4Q4Jf3y6K8u/AYg1f9d1s8THQn4JKBJOSQ2LeP4TtCHZPstJDAzbLC3epywKldBPK7i7b/Cn
yP38kuE43cYpOD7zsb8k1DN9fqwD4rbIztcBqqAxhCl66zJy4yOuJhdfev3JgOVJjJOGmvPUJTi/
ZgPGLjT/oHN35yjQyOdhhsiNJO4qS4F7b69zysAqJsG9rh2mDaYQ8NYctMymxOahb3m7aKkEmbSK
c/QfMkVLMZ1KKcd8+MuuinTI/0Fb6XbgqaDphPxymLQ3hG0u0pl1y/alFxWkdG8oFo39Udpg6GEB
X/e3q+oSnyP4J6/l/ZEjGvbZ/+gzszCh6nJcw0ORRqQVsHGsxMKUoHrA9Fn93tJkEIiUSDKuanfI
y9I26mENrZ70YVVoVl8RQWcBIMpVmdnaD3soiqo6Ze0ijxvoRjpjo9WXYM68/hwhms6WoR6c/dKc
hYgIuGlFAyxuNJonHDpCUAe6sWEg/HHqTYLgsefC+SjOrr8MwuZ4LUSA0ywBXdLdOtOuX60zRtYs
arT4YPW3tXLWA6/Af3hEPz+T2Me+yUMEpzHNdNLRZHwXsMkwwE+G2ExX0A4VfjXXdstZaGL7HWTk
pmCmhRzbQHVgdx/dw0re0ZP7xiVo37Hd4V8DrSGV+6uVBu3irrzVlFMNkJ3Aq4hix6NymtVkkYnj
723JrOAI0a6aA/F5Izp0pwjKx1Cjz4aSh9pZJRXXifRtsrweQsw4xUcxJgfMGiWyJbfBvR07Opwf
A1qWYvrWL+Wz/wJbbbXqi3eEEyiNhXP040xq4khheIhElnrGAb8Ln1wt9XmSJj2zSNJRfbLA1END
UgWY15M8nHaQ6x3/d4RnjUyvhN2yRVovbuTiHBBkjvHvfzt+4RlaahSDS4exhZVkGAdyYoV2gEe2
NCqF6mFU9hGDBR6SKxOLD1u2bFIJBDi44iYx0Mm2sfYpYwEOAAt7rm1XEXVtKpumAVWeUkmZRQC6
MiYEoSMReCT9cKbNgPOyZLhStg8sTYUhZUTpUaPgsbIo0VxrZ8e/XJsNoPeiG57SEn/On+X0gk0J
coIrzHzBmUMe4XveX07KaLyx6NZy49MdQ14/7T99mqeQRaag0TVBBGfLeUu2QHS5/29X1MK8gQNh
QSpQ8aCMZaS+xF0o0Cts2kqtW7G2QPl6lbqjk3UI3XCn+s8z0tQ6my3TbWSwyR5+2oC7uzu2wHSd
EuFZRPqruUcayLa/tglSv1iIv5w4t94fXVRMUUhwPm5SF5k9WRG9eH2ZteOMa/cPXLAJ+EyPhiYy
9ekg+f65bxGjJUDOqMHXu5hAQxdxUiAJzM0ya2700UN9QmrO3Vm4/YUtw3rOEU0ptLhONtYU55b/
M5w9QVC4xSUM31i/q3WsOSBnGn0IkBet2d2bxygcjc//6c8371Y+qe9xbrg/V4QeB+0rKiN3khnE
oAUAPM0WpoVm8xo4gB92GbD4HnXbOfCISRQfKHpR3a6nzo37aNm4V3ULFUyU8EB1WCHC8vph8wpq
rcOJz039UnpSaPQ34xnP2UrX8A9P1cRACgM+mZicDvVNoQ+YMZahToscaaylavl1tBAsvgup3AvB
a/i7MPwD3QjkAye+eyt0jFFU588F7lrM4/b5OC2ZxxM0MfjmaTKrHAVoRejTuauzdT7zIA8AjMX9
jxFHtBnxKj/bjkysAZ5STga6EeFRzUG7tyHZmC9l+Q12VutZd1P28LNSU6aTXZDXgYkORdZMNOHI
yqw9qt77sH1y6rvFHXyPvyUAzHxGOuUPrrzUPqBqVWKarga18bi8WAR6dwHnmDG8SEtlpNJie1jm
0jLzZA7bhniqznm6hqMRx4CGdwoe5NFrxQOJlKngm1llBvuzLxN1adhrMGUKcswwI6qq2WsLj3HR
GKYqVHevaVnCoQ4FA2ALR2sczIgFGVUaZsSUFKoJDZWOZjs8AVjiTzbBPZC3I9PXwbPgWtidi7tX
fW8gK5C4lR+G6rJjxKrvGhGoFR+PabfjIGrBKYrW1SmYlPkxyugZcKMqijYzFh1hFl1vLEK3cd20
Ar8XMQKYDSxqr1vVNBdfShTe5v3DQrl6Db+HroM+kmKJCGhSwQ/R/FR9Fm5+3KDzD1sMlklTKU3Z
qAKwPDkFJZmiG+AH3E9PY4KGNTZ3OJAPN0fL38pHDLklb+siT/9RH8yzUAdkqcRq/u8f7YX29U9E
gfu+v9jX52/xJFnSNw4d8qJh5qvx8J+HPQK7rSwpHCavMktuBjm/zXzBZNRzq2uglZbesKKZrygj
j1j0VR8WjGQ6NlMHFTmloX/VpeLcGv/6q/tJwqNiaMUTFN8Aq3JfjVH3hrI8HHcT4HZsuBhT/pVq
TLjJD/+RDHfSkrRIgh0V6vqBpuQtEJ2YGMw8cUhHN94CM3rnhdU7G70wwRqfuLi6HeNpdT0fmLTo
F7u1DsobN70oajs1G8XKyddfYEQ0Nw+FUL0Fv3106nyBVh1nyGOFWWZPNGuNQBlBrRpTceFgUySb
5WSe8YDLyYxX+C51NRVbCKYmEV5TJODj9DJo2qDUzFfWnDzLWXt1wiZG8ScZostVZKtZzpRlSFrm
Z4ufjecDttGFPKsyekkVtJpTVzoIqAIOxmHs0bMOcKhDE0vxV6jnsPyK4os4dUaQOLaEmh7MhKCQ
vGE95jksVgnXd1/LMTE+KuvcTxWJ70mnn6sPoHte2Ujf14IxxNdGvQpwfJvqySPdtIOwYyfUuPx1
ZZelqI1YazYOA38gegTN2bHlihFk6fJmTv7HsHNAG+11XKcYSQuaeBsdejkOSx7HfLD9MDvO8DOV
RhhbEtrM7Am5HhFlFFnKz2yfNUn+XTnVn1/4R+HvyqspDVpDsgyKXbU/5NUnmSBfkT444SJxMjxb
SLzu+5oVwWkBpuhT/rE8lP08aJvSLscnCVrSHJNIoB9gmG3cCvmURy2x84Li/i/p7hVJYfhoezgF
87zcTqRrxCT+rM1du3L8OTE+t5CshwtgFWVN/eSToQtKZifD2jO9RswUeoFJlKO7zIt5lxPDE8tO
a3f7EQcG9K9UDXQSs4UpzQPgHbo7JNsIdr5Y5ieAg+Znsa6Tew+mHOwPzjC/YL6WgRAi56aqnWrK
jViX99EMfuUpq7836/ngKjmUDLDuB9BoToatDu+oaELA9XoUutcdN2pZs2+sIdRELNrWU4eq0Pws
e9roE4ZjlDtHZoWQMBOznLCjhvJ05odHWGl0o/ibo/J+KfN8eonRJ8JAMwRjBbA6vSIVjLhAwbb/
DfcCdwsKV0i71NlsDViqOnuVzyIS7QYKptpUQbIXW38lUaVHUdL9ZUXEMvkfx4NCJFeef51AuWxa
auxFb4GC6cKrk9UCxlQJZcIwO9JR5ok6dHxveegPwC1FYeMOxwsn0/2Fh8YaHvSOXomxrc7gXwB5
7BuK/L6c5Gl+P8aBI1RGaWR+fdP3n/Jb+3lhEuJZRHYb2baiim3G9ArqY6wabYmu4FvRyyTs4qwm
TeYu4331GyPx3MnDqF8zI4oDEb31ZpOp616ZlIYYhQqBMVepI4o8v9c+LsRUQorAUWaXAzxrv2MN
SmsPTw8wVtCqrpmDwZFohr+E+4ejc/qTR8sQFXFAtE69I+AsmUDSa7adorxUh3kk9WNmk0RpRVGU
OcvQ3ao4CAmb4/AsysHnRDyidMm8PuvSReuW8sh/hLZI4PwsYtk1pLGCthsztwe2wRGLZvKZo5RI
fED7zYpTpc28q6UHskpOkg1kf/iyTLBFSXu6Kl9zeLSEg1YJwuyObBMdv0gOqZj+8OvqKO6yybE3
XDvEK9mbTKKvMBhe+Ten421vzaXLVw3DTElnnyBKL89E3WGUPxS/rMsKOMIv31FRwd/pczgvfMLb
rGWdzAIN870/qISUAfLP/UzsZQbiSIZ474WOctH/m4jtiCxLkBiKkQAmFKI9v8QzEq6uMVWy3y5V
/m7++Kev+FSSl8D5dVTagVroaD70xapxx4ssr2To4RQlthhat0Y+ePJXLFkhqfCRRBP9NQEkZrD8
zNT5qXujpAmc2EYb2qbmiYbeJvsphYIZAC1hkpJ8VrkngkmpROO7ymzfVDVoYIok+bGY/kkicKDh
cqxzU8Wr6vYFVU8d4tZOdTjLBuJGfOJEE3v4vCI5v2/9pIvzQicBPMCS4zYzCoto/h3OAX4euQTi
3PUEqxPUKY3iicJQxx3yO6D0y/4braF1B3tRa8XbayoAUIN5bP7/21TmUVuT2yh1pHhvA54TgQuV
mEZqgjorfpVvD75Xc+tPyefevyftJ/On9gdC/0V1VxYHK2syvXlLAEizlg2+1eskCTClUig8zmTE
YlxQXeoybFB7sT8VGdzKuD1Mu0kTHESBttacfHAt6SLUWWQjgdCE4C3eeGNzpWyk25rSuZzVPBWU
C8Ed3oV5+VmUOd+1AB+rKlJ3ZH8UENWovTG/riPM2/hG5ISOxrqRiVcMODrjYjoJg9ejhMoYDU1+
24lc70eiEmOsY+GfM6KZ1n6yj719ofsJrYoj1WB49HkW/F5g30Qe0ti3cQKL+4Z19VRB5yakjICf
ceiizFOef+97r3PJFDAgQVpAitnooRDDG487InxXYCqSjC9DbOhFxzz/wTW5bWBxa9JxTnRBt+eR
NFknv2UTzgut2mhtWhxURv66gLMapwMdHXutM3tHByfu9gSqszvlzVKXLbnX1yu0RAQaDk3c9oFv
vd79DbYYsuQs+4hQSfrAo2dxP0mXnTNjpTMhONlWYsn4DjpI6q5BbIc0XcJTGrn34raVZE3n7Woq
WHtzIqUzfIUMiA44TdYIcIRxQNIOrocrR0ufnCd0dZ4KZIabpeCn+8Mt5n02rvuVgxkaLd11NKzV
1pZUh4WyKV0GirOOUBkRzYRD21LrCpV7IKJpkmGsESe6aCkQrRANtnSuaKhkPIdaR9IS8sEJLpC1
iN63Z7qv6Pvy13bMNpVnwINZoVlsTABOwrg75Wu5BKBtB1XN9RuQG8Y709sWL9LMGk+o7u1YXGmk
oFeZPelioIDQWbvc3Nx20znFeL8jVHQN5sc2ZE6duTGl1JmjAumPAQZDdoEZ8uZ3rCfen2ICmJ/f
eiopBr+biAVMRn0jciKCu5KTRc0G8rfAdtdhLOtSibWbGvp0gr8XHYhmgspFqZ2ieRBahzKUXnUp
2o2/PO/AH+pJqxC1IU+eGR7znMqggfDuA4l4NYYqkn1D85UXywA4O51RcoXUup/t+6uIZw6Sp0FP
8XwX6GSws7tppfvQX9tV4tTolD2s67whPP3PYH5a4ssDQOUPi81cJXbZyG6JZidu8Fxl0S4EnXR3
l1QcLk9XVpa08vqo31omog/m6/RfAU65gCq7OhcMTenW6CS7OXkFPAF4AjA45YQM30zTF/ZlTr7Q
XXt1E7/t8T82iMkJeVBbR1hAtJBtl3/2SMV1WNm5hS0Z21on02+Ldjz4xQnFiHsqmQ1OqcAXCXsd
NtRO0ITS2iHwaKmHG8cW0g19vtDp/vPSsdUzc2Yn54FoNIZjqpE6GRbN+T+pmyHrdEZIKICQPivX
padf9uMh7fHWmvwQcIGUhY556K7OzFGI0Fek3fYU49gGivuFCEfG30c9vtnc6VGdUUfoUPeSyiBk
9RyVxSTuvebKWhXVDS8KWoPpdl45rEwZF0Dg0rJVtlMsblqvX0yRUamxbNyXoka4LzNwYN86xJrK
UmusG4yMGCJRS8EX8Tr/k2CQRmO691ClQhg6vplHiS6VbwrIKVv2kEIdpwQ5/aLSN6eK6bCTIynl
3nGk6hkYKajQu4wsNAXcSUaov0rNuaZSKyZvgA3xOPWKU+Q6+X62/mP3XRFUDAh73ePzfbUVnSQh
85AXoOILHESQ5zvJzkFqNcexys6mgdmD09/4W/BPL7xpXX5H9uPsQGQwYl5mmnEnaZOWzRIyq3x9
sXoCv/GJJD1km97GXIpmTEwq0zNcAyQI06jBYcZUoqtVnlfXYe1ppL1QBTkAHUhM3AHtYMikbiuU
2FJczn8Kja3F5GW7BTvBex/dtkccacI09ivuZO7pdk2EibGB4q9v4hmfWACnJ3lmnk0iCcoxRSBC
WFmzh7NImaKxDFTqWCyLpyObusUZMCaESaiaZ/8MNFZvX1ZJsDWfyWu48XLmz4ho9TXbtPlBsDDo
9N+BbX/fdcC1NB/Q90D2S1ilN+o0TXni3e3FHgAr/IlPmuNf+osnVqeExg6K2R1BYkYpbX3pNFr8
O2TFyKbuCnuOplKCzOurfjFpH7RXHDQRe38DTspC9ndkstU+apR2RogBo69L8T90xEJs16RAH0kh
WZPge/zNKj1LtvFZKRE0iXWT9qQky9BpxVfYPbgO/nG1M2xTDUHwyWky0kCxeksILi4K3C0ab2te
CbV1ZEFh0fJ4RSHSGO2WzRRukjLC6K+o5DyLR6dehKMDHaY4XbQnvoYwQfPdCyLeDQuAhR92o0fo
jByq0yxhmwpJEtiyKX2OfHmcSWOh386xXBgQHgOAMRsYsmoFNNV33fIaRbivWWyPoEAwUB8yW1lO
yO56e/yuA5vh+49Drc/F4tzn24OVmO0MlPKkMqNnZPbxESjIc3gBNProlR/RjKSntlK1CE92F9sM
Fea9JTgodH82CMpO5waCBrY51lWjb0PErqeMIPkfOKqLOdtCG+BXibUSCpuJkA15CfBQkyJxTOR0
e+kqEgqRkGtbTcTpLtz+tdW3GVhlxW4vhV/WJ1LPg/MYF43a7QUhoF70C7SL8nt329cyRMJ2lS8r
fXc45xRzAoIj1iqnt8y40Sp9Ac6lraNLU1HaMcl16DQl5evav1+snCJc5clq/qm1V9gBYmoOjv/2
ZTgTAOMKiexSN75cz4aUrKxGGuSo4zHUiry/ZurEsqNnQP9qbnhHC1DoUOV4MujyRdJNzKYF09Fw
sz4fRUIcmZJjndPDRH3evDYT0BYWUnUT8C8vhcjk/qoM4j/+KbpoyrOeLD8OFwZQjc/sm2y8caOu
KVmq1P8mYgipig4UDGGxg95UjYzR8v4xEev5i6B8mJcpAlA7NwAbLbcLjP3stjOMuBB+OAsXBaGR
lLfI/2u3kgMMOpknEjCIb+Rq+vKMs5y2w92Z9MS3TsCSKvB3XwJnHWIP07LszPjyVQeCL8uRe4EP
HyKfxCRh9njCKkiiVLWv6AbpDMntLKQRvWVQdSdJuwSedI0YK6cagKkVS38mNEqiapGWF7mBIUKn
ZLd8Jnq5GD+cU2wO81wQtV/LtQUAwsKGXUeqJz1yH9NssZUcWHh9cHPWQYvLewwVXnqTq4wwvKiS
u9897HJ3SVLg6fTqPj6A0mbhwUEUzp4Img0cDa9CMFKtiSAD1/DSdZMqLdK2CcVvWaHvfQ17d/jx
3ZFcPropyy0q8+BVLmKrvDnNhcmLPFfKaPxm4KYPaOKN0Ot1VtQwjGpvgwlfbrtg+akFDTGhuOLS
orjgxb6fxmBnwoJrjWfM/PRzHBgJ+OirGP1EV3oEFU9RW1QYGJevHmT8kzI/z149Z7rEvnKTkM0t
xMHDr94rrrmXbKSJAu0L3Ozm8wKZauDsVboJJ2yy6nhd9u2rKK59TSRRh9i9G/Fgzs9665eqEO+Q
Yl554pJo9HFGUTyhM4xnskwrhZTc1dHsGKzjcYVEitguKSvvWxj3hSKRmFD4jvp0BqQwBQYQCHVn
Fz1cFPI0Gbuo5vAlrMaHQLurCNBzfcguBX+rEGzPg1BQmZEklq3aXpvXjj9BzsTueRK1UP5yBEq2
+bYw4pSZ+Mad3EKPXbE/rdRcTZElnnlBDhu998185GR2HxWnv9NopIvVQMigMqsST4LNDsrqkDhI
GcPfiDA20iBNVk9+/anuiwGrKvb9RJX096IGUFAqLRrwGEGXTuQoK593np+wzYI+ZlkyVXtfp2tR
E0v7nph4ZjrADNhyB9qJhXn5mHwP35BK/c/60vadp8VFs6qRI1FJxEoOpAA5z9KpLG6T3EIRVcXW
HXAZYqflM+0tcD4R1gYOP5qm++Zl/xi16ys1wLaKGmjl52wEU6u4H/KwC6KYdf6y7Xv35ou59o7p
pfa0m3qeYYuflWQMmWN0YIJHkvbLvuzDWSc9uvlZ86a+YjMzwXN3pXa/2zQEPZMFd7cTSoldoge6
LbhEJ9podli+vI/KM/QRGNZy2/SY9UfudvsDNsoK6vQj2yQk4euBNwYQ+EorCp8NXE5DHJ7Nt5+r
j1J/clIXyYzoX7f7Sln2vfrag4XQxojIFeZt/t76UwipAysX7ZmcpODLDAd+AK341ZtiQsv5EKYO
50008J8sxUro9bhzzJg+D4+UUyFLZfezhwoEb0OgUGPm4Pjxc5ug/Dq1/ABLiXZ58gYVZyScLSka
W4E+qzbWjycZhEULFRxksLexjx84fnXvpEfAodFPHM1s3KM6HZhKgv5InmUADHdE53PHygd8WjIs
3V53dEggtKRkm1lpwRkA6hd/UtfHUO6UW373noGP3IbBPVq2/aKTCOOKETn02fT0ezH0fxuTNaVo
lgY9MQnt54RMNjjUnLm1V3Ui/coIBVUWPq0wfBJbSn29YZBBCH6Tjwq/Iw/vCyryvjSImSHXPWED
l+XlnVQeYANlc0FEQGOIAJyBUZzsph57s9rrZJGSMrWDRXWkLORjUNnFXgf91US1SZkffBep716N
/MQpggMv8qMegGEJQbkJHeSXYMsUi4SICZHpKFnyLSVPUrLOktxGKPh1ESKDVSt9Uf/72lLw9KI3
CiajcCkVxvCor5pGuiEbioWhUDbDvvQS+4rYqjanduo4jgE2wrgou5NTg7V/MHFJyBsspsgShWde
GPukYM6C0XQdwZvRW0mfn+04nOWH0mIUXd/DnwfKoSXXrlYXOe1C7U7sDkPJfMz8jwqaPW2Qbt08
6+5zNA02h4wsIOWHYtxC9kS2dvuiwfKcpKv0wH9Vn/uvoLiInI+12NzyXeIt0lzRRGjmmqFdQ0ce
kUoAZj4mPR67TcdIbjB6BWIgEaX5nSWRiI48vGr1BONmhFBpbYVu8KKDqYJZ07GuH85gfzan5ps5
v1IfoXYeADpp4WvVVRxKYQOoj386CcE31xXFefsJP190m7s95CX3IqVybXNuLWSH70ZCnLgU5+1e
B9UtmxS0T3gvidRn8gAqVKgg8wDG9oheY1NDBDjvea7ZiAitCu2uP7k7fWRrjN0iLU7NnTI/IYUT
XogxF7owc1y46ZJwsduisci2VhAqMyZEdSEz2gnC3OHkb4kFS/7EWkaz0Jz8eSLeWLu4RU1+IKbV
+UNRtvhua2aDdukzQAC8uOfLMt4ZlbeULA4vd22dphNIPcKKJjEEEJkZYj1c4sLxXlZreL6d601z
7n/e/f03TpWyJ1HgenEyKtFu+S8lzWc70F4wTagtPUxiInEPGChg2+jaZSZoQkt2mRcBoB86EIYy
dQs6kQTsi/pgi+qquF9g+bg97XZ7eFoI3jZsGHBfYSoB6CKcF9LzP/dtg0spu3PtYtPC1gWXAMyg
Wig+m1RfRSBCDqH+aa3j9ce+ZXWCvues43Lggvvl4T7Rug3C/as3mnwDrEALkk7MPaJ5+KYBih3N
LWNHseLGdIZFa5yL/qvdfJzQxW+8jzmlJkMEERIefaemfg/WTfZc0Ws7awl8PbqQhgOJpCJ+yNBc
H+mN597PuKKcMGNTy/aFskXbkztiyAwxHK7z37mXWa6IZs0UPmrissrSGasPYpimD2nAWRa8W965
RbV0Pf3TtALzHr8vbu6a8tj+lxvzwKz+Cf5SO4nVe8n5i8pZJZ9vQ6YueN3j/jJjiah0tq5KzHO1
d1bDjA80G7m1aE/kHXYapZQ2mlwAJ0EYIEoHkwVgicT4jonUGb3Yyv5XuyocorIcRK23w1mbzW2a
/GzWdfN97aducUbFwRfE+TF93/tIH6ldNE3cVoFHRa3NOXm1eXSB4IN+520BNSizjL1ZEHYncCG7
JaBwW4neRWWpIkzs8y1UF0nKqOt2F4NyAMQN2gOevYsPovtuUvryeqn77eezzhFm8w7EOeLlJasS
kbZCPC6fo/4Ctsjuq+2lbwlqaLBCxjbEAZ6lhQHuG543LAHrU22Ib4K0do/gp5enk2zfLJQ9Cngf
ly1kyl/JFQrk5kShDUR5ED8MwIbOMya13idJzzOLco2liv1lebMSBS77hsqmRil6eNtm3lj57MXX
k9e/0BPQnmqqcbPWV5yMsVSpe2csv6du1P9BvyfkzglqK/yWtkNEsRlDVcBxC93plJoWnAdMEBHB
hdiMpDJl+T1LGq8f8gCRnFjQUgjLy6IzVEa8V+ytMUKWinl1FL9jtaRi62dEMfmincXj8/bQoocv
dq9w0Sn4YU8UX70eZekl1KZq2T8wvddParZavWaMDWDdMQ1NmDnloWx64wbNvJgG7UvGCDFpdDD7
tHbnQq9Z9yGCJlbtifCUQJ5wR6/VFe3ZVi078AQJfmHaQBQjawtIqYj2EtCE9MOeYS+c4Nz3HJv+
hfSAL+r5GXinjvzZb5IPWEPpv1LwWC0QsrlcmumxoMzXA7Kt8Zuf3T6ThEztai64RX3Zrt+3cauV
wtc2q4ujSmdVHf/a2I+WLUw9U9s+5pWyD9O4gX8/MK2F8SiL/c2DgE2RTvFycN6EfaePCfjjcxHw
0dXS+poWt7AeJ35VIr/ykkomTHnL25Q7TaOlk/U6ugw3EtJ/2IpvWW+d5IZdEp4sA7CoOujQOkCb
lFNCCS2lWHnEe42B1GSy/CUh8NFP3EwHjRvJx/U9C2wV1+Dzl/CF0hMKjyU4hadTYtrB5bSeFUUA
tXh1+k/P8fag8Pooh7cCiv84Lb6jqEH9XGjxDZOzeDCPmApyDwrcGqGuRToGkYRGt3Gq+hwmQKUW
5S+x7cV7tE34An9WVyOfJJGjpl2bnFQd/u1v9ss7yspgaLP+wFuL2SZ+hDN7OwbhYleuzP84Fgf0
8+beG+SamkyJNWmSzcAsuazYafQbmeQkK422T/S16ea6Bw7LnJ8DMVRGXHijsoZughLJuLAiZ4LT
8XR769p7mgHeLwTXH1avg5L5UxgR6WlVCXmrbqfUE1nKBSntAuT4PjPA4fVoSpou/SAnpHcAvz/w
7gdyLkI1uHbuSLtFWGB6ietMeq6Lv6/gfNTS+/MKv/Sgl+nbW5mxE3Ze4BJuqO6TCjZyg7LojfW4
G6aMsOL8RSTWQxM4gwkOpw607L7Zcvj2Ub8VGm7rBuAdECAbkm80sA302+x0KPRJ4jUlaBfRf3K4
mCGgC7RcjE1C65E84GHcL6REQXUaVoSmQqTllChXIVdYMJ4cY+Y6+pEykfeCJN9SOAoT/CBdEk36
CzGMZlDEq61sf9kLBV4MQiQas+GJ0qUGa22SMNLMa7Erbqag4Q9GoADELhvciP3ilifectNaDEjL
k13TVY8xN/PgdvhMK+LF+8pf/E9Hd+OGE/KrFmKmTWUKP0NN9ovz6TGFj83ceWMZtB2SfOHbe12Y
20wEPeyBx5baxM4aAgIrpCW0LISf3Rn9BdCbHt0heO3cAccf+c/l+w8K1y5SoujUEVnNKDF29SLp
Vjgxr1nozEeip44zUMmGTVisL/STyhADZ3snU6Yw6cCrwXSCUABvvCgxldKBb2AQKyrS8ahl/zew
KMEl/GiVoUoCvpCIRCJW1oPTdbmSgxVYAjenZaGGZ9TlYnc8aA39hU8KGiml/f4xAGdKowWtRYOo
J1N2q4CmcG1jMsd3HYnuffcwc8JVJJgumYwCT57Jaw1mc+j6ksG5P82dtvhXl4GFAs2ct6CGqLHj
zr3DMnBArV495Ii1HiK3oahiILolq8KxlJuWXysJ8QRbnpfjNweDalNTBigRg0xm0quhMkDsy3GL
yczcJqjF4PliSVdWErQ6fz4RRxxuJjYPV7F1cmkEDyMollaWqKCMRG0y0yumVSOHLC3qNysWqjXW
QYcuGNofwnp4g/f7lb0xLjul40A5CNsvfmrLLrYZDLwdc95yZ+mNW79AA3KAWQytAaUbNbKEv4x3
LxBwoTM6atrEnJe54ZaDD3U3dGd+V70bx0Et9qCGHuqc5VUKg8eD6XkceHdawzq9xRhimmTuc1LK
xte68oPjr2DaDJRc3ygiTmtbTFfAOg+Jb+yu060t+iRn6M1AU5fELVleXKMyU97oQqUvf0WwRP1F
nWDjA6zrh8BcfIqKQwTlBKn0NxPV7q9Aa1E8mk9WypjrOzCm8TTJh4tONEaDV1v3RnNUVzjy1ax5
iRn1Vi4k4Xrod7BW0jDdHvi+NWoM1oob+LQgr9afy6cTCxILZ9dWgmafYRJvyrAkq5J74SmfKOT4
sHXuGHtJKBEDCZcL5cWRVwnT+vXpjEi1/t6CzFQGbGAn6mWagp0Ro98C+z8TvVOlTf4L9FMd7dnZ
81cEposnaezUDfGh34MhcQM9R1VT5weSrAD4k4iAIvn5Te47Yo2rSi3QuSt2DwzHHF5ProJgxXJh
avlNhAexZl0WkgfDliC5tzUHcfRqX2jHL/aikq5lhD3L7kT5bnycZrH66gJ1ShjC8bUnQ6nILC/T
NDkO+Ti4ZiFmA9iGwHYduKMVimYGBUGS0pgeUE9cH+lPpWjLpOhRamOXZuIdDR8JOiTrplHyGbPt
H2chSP8fv+QbAH9b6vnaY9Rc81MqKlkrfHEa77SecmxE0RNpBz9T4g5yw4tBrgTNriAOOB1VBIp9
uGkX64j6ZKrb149AYmyn8F/R3D/gp4U0JXCmBwsLpN70UxjnzaYNI90ET4Xis4SjBfuF2kMwjcc4
re+f1vCyshtm1GYNl2nk6SMSXJ69zw43NZXCkm0cbf+aQNddFFt4lpLWUQvOg7sw3vdaH/2wFNeV
mLf+KiA2RmZ1BdbAqbKoMjHBjvlwBJxdFmizsDE9D+Y/egCvEZ+oCBiCuiCDBqyBo7rflGXZhosT
VAoGX0pFfEz8uXF4xCld3Q5Ugz88JyDfMMXimLZeMhKNZdYDcZOrJ3xHeAPpEPBshLmwc5LZTMiX
KgyfC5tDbowxRVCPxYutm46xeYzOHHmNH8tCQ95r23DmTbk9pP6yBcDFJK4TlXxFMFFl/CgzeQib
C74vwxod4MU+oA8+vMRbDgN5bQ1bdJrgx9nIMVFfOA4Bwj25fUqPbww+hnAWru50gMBjAjJpxiHW
S/sX1D+RKhFIrwQFSZChxw/wTNvwzcGt6dHZAfbNhR+2oaqg4ZTO9fON7zdXaTvYBJ1IUNWBfXJg
cV7qnrDLmmfHzqzsX2lpyhm+vOaxeQG2jR22SqEo3fQMyFXVVldfuIPu/2Lv8XRMKhlbLGUKSBC7
V0Qy2GWtqkXnfJNiEz93/8nE560nTXDLt/lYXP5xzzDb7QoaXyW9pRmqwLDfOxyWJO/zg+rgayiD
umGS13dZHlMViHT6sqpoFL4DmBvU/yemTwP5bTAPxB64LKV/5IKGj0bcMWinep3MprpwYgnB4lLl
RzIWngbxOMZYUUDzniHFn1ERCBhYgKqvip5ZrTTHBWpbzXo986iHYwXJ7RfP7i46Q1pdsy/+RX9i
oxT4mNbu/GPz026RRYtO38EkxF1GEdKpQ46d5M7Zm2Vxhwo9GbcCegaCaRqARtjwJQ+8ih3WvuN9
VJNmyt2HcNUCLY8qfykZB55EvW5EKJEh1dSzb/LdSePlbWQDA8fmGlLF8GGbjOrbPUnNuYT84E5M
yJivlpQW2OFbN5TRSMrrPBaWUwg+vdx3xKEeXpeECNBV5WMIG4Frt9VxXBbb8rifVsfwpDD7R4EK
mVs3M4bMaIqawioLdeUIvCb0EjAeG7F3CAozBVDJ+dmly+TznmA+Ba+uUyuHXV87HcBzr57IY03J
RbFRrRjOafroLaIoxfZIHDaKvBxVXUp1IMYaUBn34i1MfyU9A587LeQyDKP2RMe5EkkuFY/mcITU
CuoEY4IeuEWwRn6X+vLh+RT460JlKv/V1Qgumdj3TWuW/eJq04vr1A28fGgQYzi+XgKy1jsPjJEL
saNgA621gZhYnsMINCKoogX/TUdznXjK3lekN4Z40TiPNlAj2fd7AipfAAVgmpJ1fUMlKxQAhSC+
hDDKEuc5lLUAoqZUXZT+uQpzmnDdr9cM5Hwj6GlAmEfchovpHAJIzxVfIyqyuQ1n5y1baKtvMo4h
m86Wb7qgeKDUBDce9fx150YqTZgLK/w75VLGHoICqDCii2n0x2hj2X1XBhKsj13JYgxOMMsbWeS0
KxdVzr0GAebtYTKdGc/PahNAwZUaPulkJu6tUWMEbvspzzfKDXXrYUSiDjQhRgbyAOkpcaNaKMNq
QgT1nbqKRgrJi00kixIhUyo43U3F1U4rSg/Z3WevdMGxLCnla6WEWJ0BWskK+9cNjhESh3W844q3
KWMh+zpITsu8fIhvHrzVCi6AjxEdJduBTSCyB7Ws7CYxzesPxoc7VZKImtwbJhc86s79kNVtqyxo
cf1qO0KKxFSb0tTL1qCFJ1Td4V+3FNAa/vFE2laeuD8m4XBvd/SZrJPjISRvP7QRUTjqNHaT7A6h
am5NeJLqlJ2gPdvRpGNwyFg00fed36Wd0gUkdrrkz0VvWRQmdlZ1KwOCH/csB9k/AA+H2lLS276g
5MbR1J+YiE0cKgY+jX2JMcvvtpVj7ft+KNkWtvMkoosjWCPO6FoGSXSMf7xultd3oOSqoO1W6ASE
b7ELLLr066YTdLuXuhGKASwR9kvcFGHjJcOy8lqU/ctb5XPDgeQfB30jMDBPfz5JejILjOpAm3+s
/sGxidQjXch/fOfR+PawUTYzQ+2RNnxtq42Z+y48QglvUbcqRkOuSS9GZbxIcMRjf+3M6DjYrHwK
nMpogIea/LaWe7p9jtcwfg0B5ju97/q7NSz2qd0tiAgHozMia66x/eNCZNU+JE8VeXK4zVP52XkG
j0XQdJrF8iUxaBbktHADHcVjFIOS8kYKt30/AxjMI4X9C5VqG4NNa1yA729JwSLfki7MYNdKQ8vU
dr0tHD0A54aQGo49z4TgtEDOsKtZ7pREbV9OGIAUezhZvZteFrpy8H1nZgT/ltrTJ1+x3aGnvYaF
gQr6+Y+GrcvHXWi3BwzzPu1Z3/BU06r42tf7RuIQAhzc857VC6p2y+CT9dLk3C66MoZOf6p1KWua
ubk+sHbAjo0xZPtsqWNJl2QJLDqFqwwJCPYNrw1BD759ES64FwYuh6qS1TGH/Ixq2MOibKPs4eIY
YUaGlWQXUqkt/tOEV+qlotKs7Oi7ekfQISVAWqB4ovTiX6F7N938ouCkxlB7sfzxvAV3ZuoPdY9Y
hUkqHGZGmQc8BATGXIHrAxzAkhTr7idDZuyq0zVo9viHf8eqgosARpQRyveago2TYULQEE/aUqkF
csp4cLgp77O8xDWrhdhy0beJ7i9RhSYn79CT7qU65PdQfMioo6q+Ikg+kzKqkUHY1n0QsGzBRDoa
4TNas/HQfYF3/dOBqJp/jLWhBw970krinH3DX8uKv6YfuT1oQdxw7NdSV1evVUp+K82naRjlRM+o
4JYqMfHza1wRvThN9RWXxfToWdX/h85L4czrsP6xV62T/se+CyFn5BJtm2CGzeT7gKuztuizK2L+
HLohFW41qXqtzcuRjg/UvOA8cDaWi+lktXJ8bpJX7woPSaRkYvj1YhAj2y+tnQ+8IDF6vnmyN+Ub
x0mkb34HZ8gSDSLPm47Rn2dMpux7sHWSJJsiEqmLP5B4cHnHaMz7AN5L2IRmQambOBB7mqC6ZgC+
28O2VaF4QOixdhf5UEcGXkSL5I7k/u9IKwmHrwLOmkWeptDFSLumCMLd3lczAVzhnZr+X2i4yPB9
x3R4gT9LXClPcJYegRyr2IvDVx+kz8QjPczTr1CdwekPIBHdMobnwTvxEo8dNNNY2FJrMGLTlGy7
MAy4WJrjSv7Uwl2bYipE0fi9xrXq6zAE1xDItU+abC5la22y6E9YQFXxgDvetGpfsxpB8iuKMpjF
cpwCWI7bGUSlSqmtzIRjfEcXXzCcEmXukytCdUd55j+TPF1tKEFbAHf8hP8Hf66cuczaPI7yWpSd
OQMPk6sk8XMu9XQ3YtaVDI2gNnReOOjgjK7mczWNuittvJSDOgCx9oTOhc/l1AVvVcdcHn33tWv7
shNbdp15cK2L+UqqnZB2NbWYY4KRS+Z2KAfGpD0of9QiKWSOhc9+WdyTt7KYoqJWyh4+xvPaajdZ
GGnf/3qvOhS78MxGI1ptsEdYSqavrsi45n3zYD+LY94kh9RJSef/T0RleNz6e2mbPRBGAbvzJQLg
3iE7ikmUOdmdfEgzx9j1Z6/vAue9JpmQfV2FmXPXS1t5zQbU9gck5q36BS8+euKY16CEiCHv7lHR
UaW0dctfWuEKUjowL+ngxLdzv6jmzMF4gu4Ums3/qL2k2Vb+tNTsyZRTg/SxCkigefQr1ZzgzJgb
jU0eWjv1kFv0T2mK+0/Sbodd5xSwqfaA/cPHAuNZM6d6G9I8D+nEfAl5Z2awOYu+KRnIZXgP1/Zh
0U7nFr9oTd8Jo6PlsKPj029YhA7I/IBJAVZrIUZW/RFzKOu4VyQ2mRfhTPyzGyQIFd4c4sUwPR55
CelNUN3isK7tIhFCNw1cs7BSMLNiAHn1NYFVU4V3vBGJIMnG2DnuZgJ7tZ6zp/yZVXhREKpDLxMz
oeheAF0Fl9ufih36ffVrtccEU+JT73+6LRm9cXZ6dZSV7lI/IKyqweYRMiWW0Qwu4K4yfl8YcjBS
CrddRajWMgyCX6+UxTT4RIxg5n0gtOxzurH03fziWW0vazD5dynAuWwXV59rXlzLaMY31YTlVJ0K
2bUkvhkG5g8qssHqFJ6yyii5QWVCMRVNjfs1JJcLBYlvlW46K0MVTMe9S/nVUR6UbVgRnpTz+Ucx
VgtfIkVJ3KIJYlTyUy/mo4c7RvVGU4GnlY2cj4NWVVCBTUAZoxhLDcFbPkbH05UTycgbCcktB/cW
3Tzj5ilWQiUnwOrYlE31uDC+H9nrGh2ywDJyx3b3x0mS3rUXyKzYhKmVYG+5wAz0GH/oLYhZS6E0
NdckkLddDfC985NYh5t8StG+k6jeBJ7LfiMksTaSsaBBF4Kf9Ffz50Lug7t9RRN1IceCL96Hruaa
Ijh5N2SDnLzpWbGE0MdMuWwp8QUggJY/JBT2LAO/CSXKgTsPoCEAvoG+9/UiGoKGXCr/OPSrA0HQ
iWrZhp8sIDHYuVjA+7GAwAfyDuXy2uLRZYRe1ClRk6so1Mc2/Jr0/LXmLEGl01ArQ5Bca/AVi64j
wM8Z/+wMoMGlwcy4/sFzrS4nVfrlbAAUQP0uDU3nA8m1du9ng7PtNNb+Uuy+7KVcZGI4woAimTG8
f9b5LBvsIjtZR/s8MKvC/DXa3ltJWLQ9Er5OhrCPL0Vil8Sg0Jq2XsJCEfRLqwoiZO8GtK0A5fPA
T+REDcykv/oxMN6/QYVpYBfda2SUy/CFrui5RotTMmJUDPag6qsXE28YUhauu9ghtv1lWUdMsmtL
GnNO0Tmo51eo/YQaS1SGyFd/v+0Ujq0XXXlbVy4LLEga4XNRm0fhwHfj/gidziC9ingk0FMGctKK
KfDjRveMh51fycqzr/p9DXItZD2aB6KUdhgII1xrjCX38klPldAmSIj5DmCz21r8sJ3fWXcoUHpi
KiM+JhUXI1v14YnCjAFE2JBa3jRzTGeUajItLMLV7LFMMKuG/msjB+leDsZU84ExcgxrKG83U208
BIMPswwBtikZww/W89R8N81q48t39llVK1l1ALWcYhn6xJaMlJpZk2mWhlbtmNYkQUtP4gsSbT1H
uIKtkg27al9SAb68/zIm1U0ZUq1JLfJ95EG7DNJ6k8rZmCz8PNCzFRO//wqd7Kq2F194qRS5v5uI
bTdoQUx37Mq66nZN3rKgGLKpUxCBJSr7oyNVWFeKngX+9lF6jn0dfXApEAdIFU395I15gxC4QDDg
U9nH2HHp1O/F4KQhHqWIguxQZJj9EtXvAgEE3f5aAvFP86xqmBffgw5sQgVw7sjAC8MMtQTqNmJv
EAHAtw04ZRgWJn0L05sgaAPjqGFTUQk0SU4PPNFiirPJrELFCCVbwtCO8gTm9OuEljvW2xPEKQZZ
X9QyS0gkkNHPl4ZRTNF/7dCZ4irqip4Kdw4hprDdqIoE2y1UE1to0okKvtR+NIWDuQiKTOkCrTLO
EE1mFcB/0v+/YV3BweNKrCkLhLFOroopGgL6VV/DRQsIqeF6LPU6psrL/rqYoMpmBBvbLac+gnAq
7XmayUBiRDigplkT+mtWqvdxRI9lER+yWBsrLvQLgtJIRSy/zrNVzfRqz30DKqcy63Iaklp2fZAM
TCOFpGLNGpyZobWGRJhrLyzOovTRm52MP5pAeHW4HwFc/T9TAEszSKLIlCsBWnYXRLdY4+w14en0
dx1wdVQ5CndYRpdWvJIhy9gnt3g//+dC9h1fKzZQ2ulZ/1+qe5XsVMGcP1XOOhm7o1l0sCa3EkiP
usc5hqu9KetB0mCQ3Mr2JH5IcIAGBlU0MJHUzuc1PxKsHD643nvsSqRpteMe5YzOP4f4yNIsA2NY
7gkF2Wqp45B3Duh4kmbLwl+VDmoheoVZYQmBfkN0fJ9fKQhQCCkAZDeUjeQV4JgFP3G4hDuhwHF7
9O0UhIUeYQ2OvDBJyBucxXT6eoyD1qs4UpqpQDznTHp5N4QRZGXTV/MwqUoI0JBOfuthig/OOsKU
Vtn2wnyAX1I7eQXUmdTB4Rn3W/hfrCDEaOXf1nTpMPbGmOO08Zz6ie1zdo6w1gri2uUOKMQE2/NL
q6KnEpvbNyIzp6haOgIpUBTZ0pW8R4E5IK8HzGozR/ht28gxxBRQRRmJJvmavjjpphpBdScMVGhN
+2Cqe4EQLvFEM6Al0YLzhKrh+FLNd7kZKtTorzP3lMaFcgEi9OicGV6SXCIC/qJ8/NC6PqgrZx2t
MkJehAr5YCbve+EhHv49NpV13QSRu2ZnwYPLNGN4GLfgxjeIZ3qrh1dumvwbQzmPKmhdBh2McSMG
1/EZt8XG+EK1vpYgidaHyi7e+ZI0HKiZ8eAqJciU4Ienk2QblBI1Zy4ncUA/tL27ZFBE0OTw4GVy
rotamVYO6mJrjsGrNTLPXxC/u77IHLN3NaD86Lo6XCdgmsDQa/qAqPV823u4Szz2wklec7a/ilQw
Gk0giuWpSx3u6ctC9Kvlnl6fiepamkMnLbd4yFXQO6daUXwCs1bVETp+arch4L//SMnERrOQwp6y
3UzQYxUxMbnYDaa+QnvYf9VmOLCvj7cykx8osY5MZk/p8rYFRsGfpTxUCUcAGpRq+gRXdDy0kJlF
0lLC5tqPxg+76c9RzSh/kgLpvo1bFKRlWipxDZ+CY8whQ+pxn4C5W11gT2B17RcCVIaojvtPymlv
8t3ciBElW6KMN5r/zFtXHEDZAKjkhMZU5UXUJLjwO2O8zSiXFQiG63WnLEjwzuxoUH2lr/NvSF6K
or/kDiSUVKXvwaaelA6yvpHdt4HbfHjc0LFZZBdEsZX/SSOx7b7lIBdCoMLj21zxxNd3rdYxZ7TK
cJbAdimg+7skzs24Nl7ijOFmrs9eNntzGZ/1dDigSvncSL6EliLaX9A7b9Io9TUU356wELf4M29M
HpWJkqzVz0L83l5yG+lJ7aN+TSXwfkl/yoC2bcii4bRo5wLA2w4mCyenxjGiirK0+WWEasy500ol
lwlqHCFguGzPczIJpOKB6SqQzS+/R9Y7VQu3BkBvhcpzCFm4EV0aHUvLwpe1r/z4I+U9SDtktaAn
81JkTclr8JBJB4kuwjP4lGfKuDzouphufr3Y/4S5ln/0FaiWThOgjlhffl6TopSADKKb/phzzTN0
qpRvQBfyB4ZF7xV/Ftx7FdkTCWNFjBOf5WxR1SPCkshR74EX15NMi9GQ4RLCqLz6u0OdJIqZdIT8
Cwc3W/f50qYXEh2Zf+FUkqVT5OAMLf8z+1TW/D6ZZnMgnAnzAMBbj51o65VcDercH3swr7G6cZT5
tzWA8LPzk7dlMsiM3KmSDMC5+SWYxulyyDpLnhNGM/0XVq/L8cvDKb0g6ywm1P9Uk6JK3396UHG/
PCJMgoMqVtJ94FF6auYS6SltXBYHqV8ccoJUp4xUgw806fVoIVHh7l8XNWX1M3alumTK3QuMnEu4
/MnW4b8MV6xCcE5vC1zfGdKThrzi+yEMW7HnJ/bgZRVg5y7hgZ3UFfe0t3nKU3btEp9gSWyOHd3f
IB8vl2Wkm3oytl2HmtfWRDBW+ixz80jOGH2VLGqpnZu+HKrc+QGK0aq6JfazK9lJnSwLnpk5VUe2
ooHA1SLAdDPkrmHpA4gPQSLiINBVxF9KnEDB00Nr7f4bseFxuR83xZYIFGMGULnT6CBKlgaBhqnN
ABm/+mErgXOVxDUdQrm6kNf0lSsqgmu+F3CoVTMXOJgXRIcsMFBbEV2yR9T9bP8W/Q21yvJxnNWz
Ze07CtLTgD4+xMYaMTIs4q0RYrixmuBh98DoK4CcNHzXCTtu3E7MotpNzyqmW7uS3pjVQz0eNJ8j
zCDTbB5F28yV8+y+s+o8nrLiwVY6T0aVaddyvxHPDdn7RymXQCw0j46DQ/WcomNYh3RTCHJWzT0F
YgDbMCN/Yn5aBc2mvRCAjqi79oQAK4KbbTtg4k+liEMk5IPturRWI5q3tt2d/AVD75WA6BbJ+mX1
9ZysHoYJufZINFFjJljROU505Y2iUZbNeaQWepqQkP5iNhnZ6tUD5h8RICJzL2QjEHLL11eP+cpn
cZyX2XE66ZSIRhFcAPq34bQosVTeNWcI6KS9rjU62IaLv19/sX6BbaAkCLkOMsyiaUGLhzsQak6E
kZtqhOVyY3qiXO1zORmbZjRGP9d6IskHncSeImT661bxCrOsc5UDnpFxO1KfS/jx8IJVupGnxnPp
09LpunBIf2yMy7oXUYpl3EMjx2AbiLYAF/Ws6q3qHNcXjyTZj2cZbCmsRiTy2CfSasaX7mSgmuU+
InnhzG9TiLctoYiyd/xYgpZiu5JZEyS60bIm0wOYNuLoboy0vKr57A3sW7xsxVf+i0Alu+IUC75n
HjZG/xxUMssTOeDqn2sF7v9yMMDCmWFHRuzard/2VnaXpgbmr7d7ubZnu9IqgkzYxjAfH825tG/1
g84/3CrKJz+4/GCUDm9t8vW4+mpeEK28w9/CChotCxi28hGD7tn1TB+/KOHwalpNNCfIZTRr/m4O
63xWHXIjf8XDSVifxNh2ovBhL7kZ8+c664XODqmC2AKKcM8dyysY42QDPW5wjIaxXuN/2nOI4lZ6
+nEIzFrZjj6o9+ZiriixCQlCqmUMat9kKV6M/vEIGjqqc2CsArbo7KbZQI953qZT5OGvlHVIPLya
E+4lacyC/R1ns2Q0mSrCapXh2Np0wc9IpZfAo/Drkki/BK0EK2AENcJpKtfBZfUMFoMgHiIEsDMF
EHVBHB8MwVLatWb1b+0XUg4XyCDBws64qTvl7tdWY8/7goT+vWENbyf9dNwZcrm3ramtlZ6vFFgn
wcOv+ELRLX2QIMHtM47FeygUijy0BYzuqE9PQkmRfU3rI6TD8eQk9JVlpB4YWc0MZOsj799zecd3
OwayLsPOcbPbc9h4xewXIrltRfYR9QHjd2MnwT2lB7idZwLHsXbn/s7S8hp5HQTmuoyu7p2VAWDK
wzgSiZGzm4I2aiFssL5QlMPGO/1+ccPFuVYsL57cUN2QBAgjeNmj//btlWPV3F+80TZWRhDbtpie
Une+95bC1SleyPSUNTaksxD0hcrhTr+KPo40RtsxX4jknkZuVZVNMpbMwIYBeznO9zP84s4UOx3X
/72tQqItCfFWdFlBlov1YxBsdVsqq2DBV0LQzk7oPorp7XgiP1XbJbxuyPHmVlGPObnfp3U1LNtb
0A46POS47eeQu37RZcNQCVbtRp+2NBqWFS4L2zkIHwLpGFQCwrIoRpxaK0wy+k2qQ0x/69jWzfec
gPmyP4vmAxV++dwnhn96p5zxVNikoVApLHmCUyIz7Q7MQdCI9JvZyH5RhqrgbwnquDJslGoXtRPi
jYzY0FbfvQhQfNyID5Bn19El5UkiicU1yRrl7y+taywtV5qSnI8R4veLjmotd+Hlmw1qS3MzZRPi
YK33qanYP1IYLXLSEuA1tTY+Mkt3GMj1nxAAgX/pVHhU9wSDMcmRsIlcWhrTRN9NT7vmqjXFoo+s
cRbHB1k+QsKJyjjVRzxsGWITecGp/vdwxki6vlhhYRcLdGnV1qwPTpk6Scl2MdnSy1DBoKn51A+M
EpXoYxAi1cUPT2uNKVtqe7KIT8yZ/Jf6f6ZrPaqSIzX7VA5AZM2uMjJ7b4OrTYt59VkIZBQiU0yh
CFPHsvZIJL00cJPHWbfECpwFJ+DPyJi/OLncgYOT6PRyzN9I5ursrVkQgI5QUnw0EeMPGi3biRL6
YViuT/e1ukGJ/lODLad8qHXgtmIIE7I1caw4/6xcA8xclONIIorGqU0aUxLhE9Z/CbYKVHEwkGM9
3kkNjM6mXyUbWFH5zex65h0rU60J8jwcieihWZX9mIcXd0ijozwSQT6mbZ/iFSd3wc6BK4vkwGrb
smgW7Ay24a674xQuTB476y64e4tgZ7cvDNIrxjep6OKrS0JsqU9qlm0P6UMWtK4dhlXbStvzwbQ2
TFpNeU478el1q1Yc/flbd8ol7dOv1fRV4zMHB4niRbSQv+Bi7m3ucdjQmhUXhh3l8+98R7+UQEXd
64IXdXG/akfyT6oSLKmDLQjRfdRVqKuHEWFT+gKiThUkDTYxBT0YfAjEroTaXCv62v12tbH2Bnva
Im5zCbq8e1hgZQVevjpuXznkxd622kqaUuv3Dw7bBiKh4yzdE6XIEioljufBReQU2KQInCv2XxxM
vl0Xh3VVYpQ0u6c0h7d2wQfeOhXX1mHwtfOnJlENGwBEQfwy8Ogpgc8GZSlxt9TNU/v1iyzjWDjl
6Y2aa7AAUiS2lKufLmSUCi4oo8cWaIC39xIOmOgMcUN5ySvyg4QnP1ZbztAJN8khWeJUreW4W0pY
GsiTIK+tJ8I47tx4RFC61wej9EFFrj+ZUZj+DWlYVb4yVJWN8LYXai4RlFC/4YbzxZIHZ4dwuaoZ
b6MX6A8bOKLZ0nz+17K0maxNyuUJWzmmQsA8JCELK/O/hJKUpGrM6CKgaRBR2Akb8LyLhL1lsjXv
QfHoplKLzsJoIQd1L7Q0ybYI4prbQ9SLtIQN9eXMkh4Qf5783zyj/wTNOGHMFlidgnBaa0ziftDR
laJH/KK4tjahaGNS7Ty4+6LA8MMLZ1HBoLbnU0EuFUvxzQUHDrZ6MtZb5BcOHID2K9bfFXgTv0nA
jzuqZCK9unCv8R7UMAA94mlV90F0fOr9cu8iOiQD24VYLEmuFjlM/xw7A2BD/fN/dXL0ga9MlDYy
phzxJwo/zXUSmYQ+h0bUk1pQWFKbucXPYAQvJ54y/iv6AEIt/5pT5E+bUifOnd//HmXkcdikDdPQ
Imt1mj2w0kIfFQ9T2JSHmqszwjHqVQG4eKpZFwJ6Rxe4SH2Yt/5w6v1U5ivs0BI1IjLYt+r8c5To
G47jEjOZLi6ZAdPEl8W62826zbF/Y0aa9MtVTmctNvgMqybzIIUTiZDGBORS/9/BQ6nz5rK29bsv
4tS/klywQH0Nium7YG7IRTMsQcJsRqgluACk6QGFAyhp7vC9FEgHn5/olM43HD5XLj1bKSeP0Q18
aKPbQl/RMQIMMxZ2WzVRh/IOjVsuPoXa1LMHKbMCTX5OGkdiwBN0UXAVVNzpvY3AKElw3nXZE9dW
NFbvz8+2YcRwOWfmfHyZyyOBcMDeMkrS0FzRsAx7PqRkrv1/pLpTfWQq1wIRce0I8O9t1d6+tZkk
ifpNXF/ztuodhxrPYZcVShxnjDnsUAvHO2WTS0KT+WUgDz85izj/4zY9Ft9sO4PwU1EzdAlBFoZ0
014gotL05SacJ4A13YlDqwzh8cz9adQ8PKa2q3pKwjq8RAEbvZ6bhjVawmOd44eDrnnZxqmJuaTK
FT8KANgbWdfY5DXA18BbeU3zgtiRUOeTT4+2jvgaQ2fhoFILDpcfUCDV9uTmSn/vgpTkMcq6uv2d
rvH24h/24W1d/sprJs9Sa6OH3dS3Czg5XNJMvJCliMrrI+zyslLmNzyGBxxMiqeeD0rfhBl4siXe
61TwOTuOME5tCI8aZRQy8OYYZuTX4rzud2dyDRhd+KN04U1GOsJM1XK4K6qsv+sLzeT4lizDuYHO
yDedNsiUOcQhajgwezfov4IQq9uj+b8rItfR1mjAK16FzHqXKWJrAnpV5V7yUpyLskmTFGvr/BvQ
n9TXpLmd6hAkLx4EqD1jODmL5ZeW3vOQhd+YbkqjSWY/MqXEQ9FuvmXSGG4ReHdQkMWCWxZFWhYN
t5xWOi+F1SM8SyisykEPvkUsZe+2hNZhHMhzgXbWFpBp8iu4AAnyE7Yy29tcGY98T9SAs1wW1SkM
0DFkPbyhxhMFVMqQMKF/FNLqt6xJaPzqfVsfnfiUIXNfhv20dhIDJhoSLnRXFWSiCTVYS6JMZJKi
HG5yCaXMwP3jOwP91odHdKVmHtnHQEq5HUocueESdpEo/ySrSwmekfhVgkmMkI/MR7KIwwFoquyH
ZHaX8NNVNRxUUyLGRnoi1l01xI17j/NY4eGv9WoTMqbZxjYCO+jdQw+02iK5YISe2UMZAf/7qkLh
FVYSPwCOZbrJoWARr+BHXfzVCIPAiZIv3m8bB63cMhxCGL/Vv05DxB8j8W0L1WrhLCIg++5i4nN8
KwkkRA1RY9QOo3It+FcpchyqQqJSBg1UDeN36KaTbG8kcXyOTx3doPjICEgno57SYZoIH8d5zGR3
fe3P2HGpN7RWnvBCSlnhfJOA5Kxe4gRUME3z0I1rNmbvYzbmzj/qEjxHptr9lS8J5tirLDMhY0Wz
j4horo0ic2SCMPb+7o4wUdp7H28db6RcKWhIJRVGg3hQlKc2EIgDq7l20VA6V5hyDlSsFFxUVV/I
ztSyI1OaoNCSP+N6kW1yfx5RAYUBLedQcDfOM8kv39djCCHN387uGFgkMhLiZiFPPLH935186qBZ
2xI7voemnJDSQlxaoAdRKZ3k0ivothwEJ4h+ZR+AA0xgWavC6XKkqvA99UP5s7KNPRIjtVWowRdd
cxo3vAXRM+Xs8fVphkqMRNqIlJD1ZYDNUyiExFpTNZ+ZzkIaLhDo4wW5myc/i7sYsE7nv6K4zEiT
AUM38QUQQ6u3xnXEAyQvB6BBgji1WitF3U4u/VbpMcQbbPMPhwRfY0PCifP7Yz5/+TpUoRYOSXwg
RvbPGqpxG+Mwsb+AU8m2wBxumj2qHiFlnDbgaS2QpKKmjeK99wP3sbuEL7BkkCAxskEj2so/sazs
aX3hdhDwbrosnfhX+FtClXLUg580286K8tBmEKRIbj6caRxC/3GqUt9JsNCFpCIp+PSakgBxbFbP
wKvU0OY7d+7Tp9TwG7v8MUsu4KXkM7cb593AgpjrYPTL6pUOexfgy0XxFka+kGurpRpKUzVrgEPW
+RdBAMZryYXt7OedL8OPQpW48Tp0cYcSVk4DpvyhNdJBLvPns0GI95u6cPHjiKFReIgTdWBDLdB8
XEb9CoVVkwJrQS58hHveVTh6ZEScihKREVPlfHhYMD97G8SbWyWhU7rdn3OL6NU5uzagwYdlvweJ
o0mXvNkPINPDk/vPQGoPnzJhfPgd7br18ENGy5URyfA2AfTCNn3PECsuyRUZaZCKtc5HBbxIAtZD
orUKxdYoFmYpK3O9fUdSbSXsCZkJVo0JRUuy7xF8WWt5NOE23ORl6VOWEJ5VDYOGtQ2X4FXundJ8
pyPL5fHwFHHHorpMT7tyQYlYuiGFpZ60SNcCR9FgKRrXE2i3I9tLJIha8s3ajPE0v91SdgEYbyf/
Cmih5RkLhqMvpxHsUyUHr51J0LFYUqDcFdPbhEkuOoomgTsxuaTCFRzHVM2h2D8b8DPJ+l0JwKvj
adHCvlpR6Y1ZMAOWtpEFhKa/6wtZzze1UKoD0YSS7AijKsc6UfOukC+NAf9hX+PEMq3+a1jyCbJK
+zZ2CkMNHKnCB+wb5K9H+AW77aSPs/ugK3eGck0jgSFoTaxU0Ziz1VClW0YlSwvvC0rDxTs0+Y3h
kLOiM/a2mMMtqp58NdKPfs1nFnjqNr08YbW/yP42+fBYNmYJgwxIFR+EjX8cjhFuLP4X7k5FfkxW
Gl0l07SmqKv8i6mzLngRvCbK9xMUqI531w/JZeIS/93YFxdsKm4lnClOFRzQ2cohPflqH3qbp2wc
1/9sAzKIcXorg/SYI7eGMKeskS2i73cgXjbaw1CiNzSyDG0zLUFKy4QZsAYzpgd1KqqG09e5ODTy
toQ9oI8MiC09++MvPZhu9docUqzCYmbDC3y5W/UF/PY1J4lfm/2D4sk6SJZLI1QCzkV+QwrMVyQG
JIjBr7x7Vu4Qf0nrMCSohbWZFBxHZRSfEhtTVe+CzYnf5TrRJidoQGoAbRSOLeDaEL0vqGAtl5xY
9BjV2eRBpIJXU7gyMg2XB4IQ/MJlLNXL7OpGHBLccxnxii65z117yqvvBB1VaVvp8CTmSL30jpmT
MtIk4gNPBLURajb1uaN3TYwwWdBtZCQLE2YzBrfNiGM8QT3ZRhfZEvKjf907C7LnlJ9LJzfzzFWW
50rKRW0Z5x3WjfYytpNfibJ7Bs8XkXxvkVlz4nEAdcme5qqzXoeRovwxmaXfbndtWCLppncTc9Zr
N9Pj3xDYXVB8CUkbNzP9BEr4xd12p6rwc22vPeywkMssulnpLVsYiXE97CKPwpo4TP3FBOeSOnPi
t1YpV1k0JZuCayVuJk/0bJj1Rr+ZgowsxE/zBgYR7rW4H+5NAI8J0hVNi1U/ODE8/zKL9J+rJDvE
Jr9JPiD7cpYUmlu7yEPVsKMa8joFMfQeBAVw9gyVONWI4421oqjii2P89fOq2J1z7SQw3qx0ySnm
dHKFaGr2VNbFBdCnFZ6lHfXHW+GgQ68CpMGUkDxrXUY8r+98xsaAS7PBcNxAPdsvIRkjd8YvenNL
n+USw345U8Vk+M7QcwLsDnC1zrYdfyRog1w1ozKRF07yEt5ka9wxj8sBOeH9vUojVtBt+rb1eSbT
Ro6L8DRW4tzGi/RMaT/vMr0KL8N7/gfRcErNzICiEj4iE4q0rzpS/QknDwfZxEdp+vYz+0AIDs0r
5ACNV+xc5KYFqDPcpqQyFUmCxoROzTB3QOfMxVgiNay6O9V8/uvEthZxUCscc7BnNAvdfJ705NiW
Z3YNSGotf3TMeEdtMclRJ2256ZDG0A2MtT2nLyXO1g+iMyEj/BSHkJB+hukikqzQ/Vry+Ae7dsll
oEO0EktQZF5ovTycs+3BqtgRmwkovbJr1TAD353UqdboBWRuwdVL3mnxOgCSapq+Rr37lIBpvWDC
+lLDOi22H/2UPOcB6sQwsaPR9UktOq4V9QJOfwYr2+v9y2uSEpNf9cAF5WFSLymUuWLuR20ozjWB
/+o1mcDp7TxXtbQQc0L+9QrrK/UYFKjdv7L8+fqOg27WymeDPROUWNfOT6nIsq3/KxeOJhMOcIWd
i5R8puTQf3Z5h5FytIfi2JFwW6WNUydrgVfpl684MhTAHP7fGj5Ztn3uFufxM0xWwk3Inpv2RlEM
mEzTcMsrJXwFKTtjube3hz3W0ZS3irqcy8xd3QxJiHu9UUiNrB0YI/PjylBbxSqfcVYjpGfATXDD
+LYA1+nJEY1TMQe0JC4F6N2OrPrCehfod4RZXBHrM7pPe1gNJTmIAo/jQIf9kMTG58oFf90aeoQr
zfBS69VD65HR4RGdafhiMtkNNX/0vCx9lvSygUZMhXDHtVNdjHv/vkGuzeR+6LbPs44Qoyvc6WYR
PEMVO6DQKC9Hj7tb9ijOGpd8wx+gNTNOWA81AnTo8fG4PL+s24/6DgMCN525lqxDSrsAd2a977qP
+7Lqf/JJbNx3aHlSDZdjP7Bp5JF+ArBWg/4UddQyAtUeF61jMFi2Ea0jrJbKG7OqaShs2FIMSV+A
qw0UeCseD+1uO6A1RZRnu7bJzwU2okyAr0KrciOsDmJZ0GBi7Dm5BpETqyb6+jBhRVbQXOrxbZ84
5SweRzx2Qt7cD9tr3kaxoqnLxFTqLPBX7QbZISHIvoLKUIfIyuStd5kwkmWcqb7lQQvPZ1CQFzgM
ylu8LDGUli6hf9eyxxME+Z2X7hPTtu6PWa//nLn3bHWslH/VQQYnBnplpurxXK7535NUA/HcuytX
tHudWQkN/oMwt9ZpdVnlqfMITOIiONEkosbBIlqPKJdzSBFF21SIVn6TviCfSKYM7JnAuo/6wcOW
nBVJp63OiaDQa/QVUP6yC9WRF1OJySQbYFDTqU23ZWPSwVfbjjtk7cakzmo0/X2vy2q5srCj7j2V
VrlSXL5/D66Uy1NLhxc320OKjMktPOu0NCobfx7i6W/ehnmH6oAd57t5G8ND6phs3+u5bxXc7RWF
Co/VDh+Vikl8dbWx7QKq/q17yxLY1A4NxugMKH5jVSGJ9FCC597fky9VOYoNhL/bR2tr7UaKtf+9
pJDWKLZL0YI/A3pqnQAi+wGja2C6KTf8fIKpHM2hIYxxMVoQ166SvMKTGGQiTa7gCZxDED2nzZhl
1vaIpygYQ5+vVuvM4QsMJa+rpKfq2LwNtDzfeY9K6tb+9ncAzE4jTAxM+0fsz+RwUUW9Zvl1WXLJ
pFjYHl5tJUvQdRSq39Uv8FhTjJgVsJU21C4s2JM1wW5IXntTC+W4d9sSgWOF54H2XAAsml0jTR5P
SFPNmAdu80uAZQeSbEe2B+4/wE6AdMRrNHH9u2FKjNmFr8XSNi6w6HUXZ9pdNqasWla1VoFd440Q
FFGtmKqBFR8ALkY57dn1+q7u71ra0cQhmlDtNyrn218tQlFkJGDhMUqPFdC/2+kTPHUd4lUIcYY9
4+XQfa94Soim2kHgEyEBVISPseqUuWm83CRd1uz6A6+IR9O/BogaExsfpMZ6evh6ShmToNy+UIcD
vDIfvA4Oq1gKEqaVjt3Z7aWzfhRRLoqN8xNMCx1GeQQSXoQvhicLrfFgpkC8r/6DN4Fi4ZDT1uDa
RDQZhhkj/wEmrxv9jT1JhaDPsdoLc0M2/yzPusb9XTuazrUSDVnmNZdUSV5S/KERV+UcOpBfwT8+
eWnjNt1d9j5fV8GiyFuLfsa9useG65S4BC6Pspu8rmDVtQJvvze8Vmt6pmZrXUs6T5lGMSeRgfNv
cU4GV5O6oW/wZ7iUZu50TKYMHYu5qmDkByolzhL40BqfkVdQ11jMfny59AaITsPkyJTkXmTWFERM
JZoO1ac6KVa/loDBTpjd/HLtv5WdlCC9hKnvFAMWWtTJc5luWG6WekQW5MoJLP/eOlrgYFX/DarB
azEuLoyeyxIJnEju3fCONkfyeCYP3LzP0wJx4ISu48T+yMDooi9JixmxZ0vZpU+2a/3AQv+tCHrw
bj685bf3z64taNG/cnA4j+Nrg5ku2pmgREk6KOwXwkSEo5Eo2Yh/dvKPUGDDzJj/yzm1bJp9KtLR
SozQ4oEEGjFifihRDseh4CVzBGKKbc3vfCGCEZkYLaWsDXCC/7rYBahrgQvfeBgN/T0iRU2JfeQs
BJ5m6GTTLuwuaQ7XLcWITp3beZMRlStHmY/PiS8W56u5bxBV2RKaIGiLPklWWFNy+RD13TyG9ifc
Xc4iKmvsV6CyKRYJyboKEbVlvgJR3+um/0TtP36whjNFV/MB8Krx19GrrOkyYKdYH3OTWpKoPDVh
vadfnCnXREpdVTIj2/evgJMHUD/GxmleQd2DnlQmU2b1D2Psw3QDQLoPHoT+3NBaCJ6FMW7frnU7
KDVIlGTsrsq6vi8VHoMWBhOMcLZLjkmloM+KRHIsdaaXmkUKeKgxMTogx+tBL+EVLUBC8ISNbxaC
CkEm4rpdNGJeVzfbfVHnCjaZmJ3UczkJRrW7X1ePy38N+DlXyX5zGVZWH5U2/OHX5ujsMxMMIdbP
i9eRqp3HsGfG9IwboXlOtnibSm6HavcsR2BdGR7OFN+rEknpC3mm/xQgcyyHDlAxROe0yNMZP2te
o4LXxonz0+utCArehQhQcPdhCtNfSOVdYT60exJF+IIiPMi9k8WHS3xcdbzDb2C+MPZLinQH+Ku7
V2OAJqkVXmByzL6i7cj+UGozpWcEuyAWucFP4+azgEMgovuRdz1II8VoIDQEIiyWFcb9fdlrQPU3
mjnba2OPuIEozhWZNOtcKk/DFJBazkEtl0ZgFrV6328w89grpYjil1u/v1xRuvscdnq95/kB8nFe
rvrEn3iygRqvbo15npF8coFMHAPQYNllr02tbyjbhUZpJ7I6yBCF7mvyvseykxEL14jz0zq5dKiT
ErVgXA7q7/E7mCTiYgxdyjAz9ZMUDzSLU9yjUMBKPescuO+mf0v8/+PCzLqrPkrmJ/+7ZCjkKNEW
dPZ9k9ZCmIOxpOwp053Jk8seLkRcIG0SSZeaAuZAzOZ1FrLx5M09Hi+z5qx/xuTCCr+qUoBNtLoL
e1VHKZEjapdHp4u2Jt+0WVDjptJ/tBoy4ONXkqASq8etZwBR81wLZPVSAbQ1Ai/WIXRT/hlIJayk
/5SKp8ngQEscnqSnZbzUhjMlkTk8EIR6qlcy42Ib+dQkYQsTaMfBBawPfARL7VgWjaLy/DWiIXDd
73UI4SOwOPt4/Y1jhbyTDwxr038qWiKi1y7I3ucBTco/VTJeOw6jV60WzDorW7wj5wGQ/LoL4mee
Hm6Rzjxa9csuD4v5p+GucH4ZUeVunwHKJqIMzxH7QSKFxVCLiVMImeNKZcukb9wxVK4nURTLzp4S
3i95s7e04jd0Vly/g+qRlT2DCPeiMguWvdk+YVYQGKlTc6bN057WBbS4hbyUG/Ko4fCsmj5M0o0B
JN8MHiGsxsXzjjYcK62xdLN2c9q1pqemdPwprGf2Nd1XxvkT5lGh9N/mg/gemULoxKFBG4oKSCwn
sVFJmuCvXjRdjgKrsXX5rerSrBe952KqXDFGoB8D8hWGXrfUhMCMIBteTbi94mHZJWpY1ukHUgik
AP+zx3HtwHfEbvXPGBaDVpBdCtCelwc+LfA//TDFe+4vyErxUdFNVwBPUFhrTTxQl0gifnMR63Fd
yydm91Q86pAxcPVG1IN7nFH2BZFPTY967STGirkpio737xWsUd5C5kaSN9duNjG2W7MzCMUGPfMP
+V7pXgFf7tgsBMX0j8IiJxISmBCe00aHBVM6EljY3y3qcXh2Rm4ACMZHDi3jNI/VRHVnn2uNpFB0
E1UQDmPLeiIKO3Paf7khyUEFmCF+vH1vDq+oMl5UnAgPTLpunmVt6UXnE/hwuEwxWs+EYXy8oFna
nogSaS4yY4ylxEfeqqg6gx+yMfztQ3iMhDD5AiZgvolZg+kuY/8NIuztSTj53XQwkOev7LjM3AcV
P+nRmqpMHwz3WT1EbyvosoIomGOeS233ohC208cxpQ1FfE1EJxilcG3AVpgowjEPPJ1mZOdVTbdy
qvbGgl4ez9AU7ZXgiXoYcQG6SrC9cBC6oL67uxUBalxNReKdE0tziB2/0NJ06DMF6yaCut0+QdEQ
t0WkMXOu1vlfuBxvGyR3FkHVTxNus72fwdEaIF34OXYy7FAujiWChtDSAIjEXzsQ33og16FKU0e0
5KADSFORVFtA3pD/DtUGe50e3qHvcmLA5zX14CPjhyxclmP0iaIhcliYUbjZRc3n1sA3rI+LbY6g
3WCe7EqGJe94PgKcHhFlkahRWgi54WC6k3EbKcylL/zb9z4ODJWdRHQ2+GdncRuf//GZH1KTn1TM
9RWhgv70SDKwoxx7zJgbl4ut68xuisuvnBkNKaUmETdGcciAfIpxoQRXh5C+P7DftOYMm7e78D0l
JkQZzikJbNtqFB5SGr0k1cxJO5wD5s5Ukbzx9tg5Wtmk8vjIwXWyHPScTTOoCGWVQ5kNiRUbtyor
BWXb5JucxUxaympv596lA1JzjY7/YmPS+xuXIB6+rTbjlJNTzZ7SAtr9iqq6wQJTQRPNs87PMZ+w
+vRJqTq0PyKmn4x250zKUBNTGCBdFYJceWotqoBYNdAWS93lcIhzBgJSZG1lzhX8S/tiBkk/mrE3
GZ8ZoP5O62nN7Xr4ihKNRnF5loOPiw9OkQNYK5c05fpTeNp1c57fnXko1It8gu9nPM9yTPwobiJ0
45bnhtXCyXGq1OfIMQpqnyWzoWjBxtyg4GKS5B6aub7/1G9v98QyODDbkMutmYkmLRalsmN7JhvX
brbveoP5iY1paje1VtLHDXK72V7apUEvFQyz50NRKeP6wfs2KbCBhuTK9h3Fl26prKVAGNb2fzT0
Xe4MyD2RRH5+jhGuN2r4LSC48k37WPyHupHGQSFa5srIRAxnkLzu2U7FFtkdtUBfpAOmWOfcnb9G
EYwM/556rNi6cyjLANJ9JIsIQhYLp0a1bMqW3+LJRafGxi06vOGvmjT/2X9Xu0wuNGxKDR08IshB
dlYZsuWnBouM6jPq72ACl/GZHnXf1bz0sfy+KHXHyhiYEgq0iU+HKrSDBhG7YT7iughnVhfy4XoI
R2xLkak7xwBQmg1aPlBoFD31dQLA709YWTa2f+8Xzn3R4XTRjs/ahkpfxSsWm7zoA1qOCJEBGDiZ
arTo1qP8Mtire3EwWpCOfknSf0FpOEmbfmmngYyQKMKQQiuY/Vid85xVVXeIpvTdTrwOD8lcp2m/
VIZtcbw8t8GqgkSYKXX9tzl0ai2M6q8Y2KDoz4ZMHMnKxNatrjq1kIou/78CnBkpROQXVxY60gHt
6ZSynpzMPLVNqKptu04P14xC9MUAVgQY8FhgRbT8dD1e0U0BANbGrBLuua6v5JzM7T5DzuCfq5t/
SwsPaO45SXuioApFxbhnc2gjyVey7NMlm4hIdfuaJI7S8G0qjPRMI8sioNL1hRWiI+QxY+KBOeMv
f5I2NmYldujWSQLgsSALTImkkQGCPpLetlhq2ck0PkEIqJnJcbDUP0cCwTHnuoQTQV4EoyZb0kWO
Hy1WBEDTU47HGFnpoorzUXHdng6fUWP1QejA2FFKRiCEmPxIIabLOrA1MNOuPauBg1pABHOHcHuZ
6t8tiPrSiKCtut0jmTqlsQOueDo2waAh36d+bS0dC6UsIqO8AMuqCCw+tXQ7yQGALyuOCzIRlamA
BYsvaqMRbKcvVdyORewHa0Yv+3iIdimN989g/8Qfy6xjkpx2yF5kjuX4ug86EXmUH6z/3ntRgzlN
JANhnAHb8EC1kGWkncjb6KZpb4l26HMhqu3AgAVlNxZDpM1uTErEZqpfBZUw7EhdSeEfPT2y+I4x
SzbzIgow7LSeunZHaTmrDPUR2XPrnY8gHCV0V+gQIvJ6S2I6534uwaw0Z6kgWYIRVmhuqX5m1rD/
iMWHAVDmtXmMzuj2Xkijp50IpPiBndwu6eX9EbfKZCxGZnfuJLEsRb974vyFE2ghi50grbG9edAw
FKRKvFdzFSXtWYVHqU4eGXQq3hH1pMhyGeph1fAQZiLtQnSNDOjDwUMtDb5BmIjSR6HAEcCq0CSt
zsS2IdUxTlFOvXGTG8GvS8ExTw2lGoNxPCb0dST/4LFX7gV4LNaDTb+51oOn2g/zu7flzsjA/00s
9EOgpAFWI+kN8lrXccrkIChX7axRgz6kK1y3kGfuXdRArymYMPTbFSBPWPU9nc91HJn33uIG9gzH
CHlQLNtJeiS8lloLVxj362dfjO0fmgiMzTX/drOuoAkzKtJcO26t4ZzXFvpGu9uDzHzVAyXD4lKS
pHIlOUEsfrbTf2Ca6smZMYJd1MqTmCi2vj1OfTj+Tqh1yb1BGRCbf2+VjSBRpM3YfKtSFZZPjO9R
WylRLWS+YBfUoMamonHZ0hl5l45swj+vNbc6WOTyRCsJblHZbWtPGtdD3SzZAofF7WjSBbQu69AO
b3ZZES42OTSi8Q15BGkmY693FOhACnus64pYEZHzOdwxZpwOqVl1YgJqlN8R4dTgF42t5THWmzl0
fsHzYgTd5tAxuFzW89neD/l10S/tvRTmcRl2j/TVWfNsCVFou2JbjlzEmvdcXx9hX3/VhIqVSCI1
KGQdPcpgkTpKeK4RuheHpWX660mWrkMRbSdIVHn+GWNsJ7DoHMKyoNatmJ7ogqZNiFRg4028plam
w6LKCAKRGDV45Y1ae63yrdzmrwRE38aA1UnDjKF1mz7+W+kJBwA5dVhXLsdejM8f2DwvT88sNIc1
HV4C+eHRE4mWGeGuRKYItP6l4wYOLs7Ho15dAre9OV5dn4JuCn1n1QNwJWMNDlHevDQjYPEMEhIR
iP7C9T3ROXqh+JuG6OfEsY1SkBSoDga3Z3kOre8LgYMJsPo5N6BTSHWqnGrpOEsJV48U7JclxLAq
cIkVNKc4Wdf9wUl3a280EI02Z1ogLUT2oUhmcJbUt3yupE9PhIERpa08vcMMnWQ/odf5X0STne52
n9ywLyR6QX5/SJZoNvp7Mr6LQvAO+a/FVfjxFjDWZkVmV0HSifYNrIeo/JSeBP7/NljVbvl+UTXt
14i72FSwjlLWP2v0fVsIjMW+FgtTxyADlCjAosmVFiIyDDlY0le0oVNJzVuvg7FR6/Au5SXUB3Vu
nnlEOtXAX4V0CZ3yZcvwmG4PTI3PAjdGIuaY6uLkibL0jF4H+OxfoGauCszICm/EAr3F+lONKVbG
Umojt7X5Gk7A8JuSvwZlgo9/NEbiEEL8M+PcylrfgyvIeg7Hpfzrs5d7DZG3WmU8glwUnzLVL5ii
0P6WGxl/IFtfR8XE4UUoFOqZHrYHLuRm6UeXwrH9b1ptgOtgiYuKdDC7379xx2XveGxeWmhFiTE/
Veg/z89aey4jRDQ1scro7RTj8W25dqQMk+AwFFfoj8a8fJtp4z24Y+8mE1+EEWbw+/WdIIvRstNf
tedcjuNJLuIvdLk2Q3ID13Y2uBeinqdMZY3UybqnRRJpcIMsaq+zA3LjLV43O8uno2P400InO4hK
MwyMiTzouUJ9bSHvhAGjnPTw5I16Ds26+SNE70XTRzaMwyZAbO4qb2DVUOdQbHPKHI95q846pQWm
PQZoVDMZjaJJOorumzoPZRMG90jBu//dLjOCbHVH07nFQZXbr4l+62g+UNXAjVUdlGJs8niaByb1
XbuEhsD0x3OVz+8Dmqxo3D/0uy0bq6FguI0QAVLPIlX8vUvQ6D3/aJoKoETRhyIqIebMlT4ZtYSu
5NepMi0dEHfmnavVvNdWRJ38PNl9QjamXAcSm0rjx8ZmtBATopkRdYasWQmidIG8D0n0fsocYRg5
LiJa5jOWTsBdu4/qVfAzFM6m0PMmEqwQMzOYidG1ZoW3QNgFJP8flyrL23z3u/mgHVMwokfpAqHL
pU6s/g1ARvYSIrVz7sLM310p2BAWtSlAqUvj/ewPf8grWOGXCd+XFEn5Az0R5OES+OniybLiQ2DX
U7Z6Xhq9Hoz3HBM3qaBCCsZN4FO3Xi/5bpEAOeR6x2HRGc3Lv1hjM6gEEqU9M1+EqWxx999Vuy7c
8sQ+7K491zsiRa74gZjfdaWWmYt8QJZe0pjBKBu9Gd+nWTzlIRqrhivlspO2j2N2zI+hfRs2wzY7
1YejYNjWKkIN6sKOuT425bd/gW1e0IT3iMBC6YonGC6bw4w6/J7L9UwF2Nnl9/GssaGOObhAVKoc
97zJrY/zCjWCL+QkT6Mtbzd6J7SOzXeq50teBhLMZ6mVMYhRi7bkVfIElwalaTP87FEg+09j3SX5
raBNokEo+g5WJmAqgYIob4pQDTYNuVN8cxN9Gw3E3NlWZn1Yt45N0iCkJil0bC6x/gVc+gC6xL5k
awFrGvNpNeV8EdMW2eRpQI7GgS32QLVZX/qstjgO3JBm3bMHYp0+dQDGYvAG7MkZZkr3IdQT0QpV
tL0gc/7OVdEefYu4MkYsuxkhHArqwcnVacVdxgpY/H7TF2b3rgp2hWCFnyb01Whh7lQvlLGy4XBH
Lq/YqCQWWVoHKtIiepYVsAgf/g6opo9bqQtWe8ehWzZZWEVK1qpOxT800ReVtiu5ooNAzd4XdU8J
1kupIl9zMp+9A29JDLZyYQMR3J8U7YoZYvd6uupOs8cw6XVN7vPVCP1Bbf1aHvV+VZtkyMEfFwCE
hV2KiqrEC7HiNdh+d/BW5DzwRT3qvsCqdXSOhDtQcm34o+NYml5jqBVFPKLP7vFP3FcEqEy+iFeq
BPUnudN8biM6K5vBjXOfAf9++kBYMWcNqJzmf4uO7iwoY3KNOLcKph3McpNE4zXaUmKfYDHYOYeI
B55zoObSRqgN27LjFXuHrgRM9WuLggbvw0qoHIyMSJyJKCxrYDq0zsAe49rezRT0H1h7DU8fQt9c
iIcJD//wZqIWA+UgFfx4RFn2OJtRA07PpDlofChApLzNGgrOfk496IsX8YZNf6JMHxX2dtSECrHz
e2/u4tsO67MT6o8XRHYm4eB08tOYhy9U3EaPCLhGtnT1Q5kPMiK9RVjzpSkZbvaRG+RSv05HVkCX
Crhn6msnW4BKU2vzdoL3sOzUTwhshbyxDiESvO1urJO0rHpokaaURyjuDc9dJVrCjwMJtEMvW1j5
QMEtr69+4NnQmUHPqyoPYJBDuUcsaoty3U+DLZ/XJgfOfP2rkETg+TkXYo/rTALKmiTyiTfG/iSt
6eBENGfK1ExSp17ggUnEwrfCRZzlTsvc59A4NbN2ZRBBZe1XOEaWOBzpSfx3H8d7HjlC69oyvvLw
rj+zLQewG7WC+JqNgx4/vjEFNQ7VVRDIlManz3Niik6ABLb84XJVKRo7+Gifpigsdz9Ajp36kmDP
Jz02l2kv08GbSfRxcH8Pqnb0GbnOcxIVr1Pq42HuAhKtcmYHNEl6qmiwPCalG83gnbGIwAnhDdbH
jHOEEV7OG3NrA53VtVD90ScD2P+VJTk7gXJ0j8JGPHhUIW2gdOWquBoUm7ewoItaCV+8E3LDeNoV
7iONk/dPbDCwIZE6LkP2uDYR9hkxNbEUV21kXylQNVJpHMQ88MtQk7RQEZV2U6l0U2UVFplWlNwm
5XOaUJ2Gl9in0cCWDU55dXvGif2Xp7/pF7MJB0Ws0LGsuR3EA9EOIpLSQIojuLRIC5IvjbW0qVN9
ntK19JLJqYwHJsefLceADE6YThzANCyClPYKfZOllRxDActtUwCPAuZCH2OZQbMXraTC77Vwq4hY
6zZVWTmwWYL+o/iVlgXy7r4UbRjot635Vl0e8Z01UFPuvsUWbCUUzwcDyQDpzGBdsmxV37dBiM/8
fERyWCI3XptdGDv23K5gmpp0qoCzgxECMGPpmZXa0ks9D0TSE1ZlAWjJVu0BOYnzSnF3a2+qNzcZ
lr7ka9w1wfp9sT37J3NOlZPkI4MC0+RnyUlGx+IJ4yyJ1gBNTFStDULXyqLHSJN9O1YG9SRMLtqz
Ugrd9ch8Kg+kHKiqiW3wsYc4VZnSxmB7jUM/yEMAmHn+e73NhqyJ7fkOPcZ8VLSMgGQxMQ7kIXEU
Lilzm5mkNFQHWKi1MbfbNtEdO7GEiiXNRHuqteoWP+AGlvBKQGilMx01x/i6TPEhCaBnsjMfnoFs
/ZXAxMvzeNyd38kcO++UvHJ36zfsnmNtjwcT3Slk/gTnn3Mm8130GHTQ5ukWDkIhgFWsEbJs0fsD
pcaTS4Xr5ckDL5WqvXyTqlYQHcXH8Z9yws65/h0eYkDt8s6iNwr0tiWYGNJuyBp2zJfDqpMPTOIL
i1c+0PBrcjBuJPLetSdPPDRlJqhzPl/lonSCJEx6jFP2Gutp1HdSGQol1Q8NYtnMQw2wn5DHR9tH
0xrhICUMyRtEVZgl6glnLdXCadv0szO6ueodIUET1HH4dNpAxPwnDw2p2tJatEpPPnDdYdm2KUuW
Ul4AU8ZAYolzTdtgj30sQ6dGhzxFaNU9UCFD8Vk0hMRdGpFEvKn51PFxBk7Qe4UN7pZdW8jAj8lE
DztU7udiNBV2JPEbz892Kv1RqqIU+VY58zmhjnxF6p5LPh+P6cZ9lt8vMJOYAVlrCBxptPqtkNkK
EzZWOveY3oPHobtBYYs81pGnPnJ0rgHVdva50OrMNQtPs5lO7TEl29P6mMYX7ywxWKSLOr6/rMaO
83ok8MxH/HQvXgi//j9YZ6rQdEdWoKrpenFdzeOc1yfSQwix8rCjMejpGfbsO7Hfdvg/+mNigU7j
G+dvd97dKZwfTPpZhFUjUFF+jKuSifyvFCmuNDR5OmsXhbz3yyutTyqCBzuy5587S6Cp9dbJ8I6B
Lmlz0MqlKWBAZJTQBqlVXncTbCMljaQAtMlXSsBbX7BTZIGPQSao8QgrZXZD+AR9t0sCTT/NhZwk
/kVDtYwhvhVuyzAAvbfVIPaefChqx/wcpoGAxgdFydBeDPdWI7yHkMcEwUxqQeUQwO+RL4vyBtbS
ed6WkdBb+umAPdK70POxFJ5E9oI4Lj3Mx6r/sUcQE4ieK6VYmUdqa0VR2c0KW57+YVodlfzVoq9r
/Yt8HbHiUHqgEtuYlRL7AmEMVlywfzckuF3ULOTO8Ctpw4p3++HYGilE0H1woCDKmPDSK/s0sV8/
uSK6UoPtdZRFnfvn+fdvHCavVk+gGLmTnhD1JBVJMslZ+8rjkbXs4cusaqAeMEbXeZdE/cV8PBWJ
cWMZefwJoDbLBcvBSuZo7gUtG+pfW1KXSTozKf69Zc9oFItyouKbAgeKoQ6Q8bS+pUkwtxKwsmkQ
Z/l9Wa9jNPvOs5ZPsBY1svkW8bUpIJh6bLr4AdQiRsBQcfMc7SoWe788uIm5zdRkDpeB/vZEDkn5
Xlo6WQAg1jiait/xiDT8e/L4SGyYXwhd85la770IVE3iM6kSVm6dWoaapELH4lBobj/4PxClmuQp
74B8dwrRQkIYeGauFlWt/dL4SRvEtb8Aek5owKRz8y5knShRafRdlRAbR0ecdxRVbj62qXbDEf7N
TZ6gEfgHXuqBjSF80XdIqH6Ww3uRCO9U1Iz4CXMPz5LhQ3+jpGFaDCwM3Vzf+E+rsZM5BzIw5A8K
d7zKWyRiEi5smvcDiGiwDrEYEsNskVcNk7kDxMTRD3Qu4neZGmuVw+ajSJXofhrcFmN9xFRqMAI6
Xe3S06rynECiNfYpOfGaPddJWo1AB71TeXK3ErY487mZ6g9w6xXyC+Jc22MxM/0q88XZ50XVuMBr
s9s5zy50WON2GiAyBtuMUD5cdlQoLqk/UJk00Uizfpu9882AuM2s6Z/hrAqjPDC+6MOucsFMpccH
tJwB70sPcP5TCnCLT4n5pyGDMHa44GiZabXD+L5rVtLsrp7JsV/dnp5+/uTzoyArW3hakzmOLerD
i/04W4mCyp7s2HIZ7HmrasSWlpKv27va5bTnNUNjOGHCZf5J7MgrCnKzlyJbioBtQWD6QsHCbFEK
Skv2rFonqnP+IolfyWH3yYgloy4CAtisoMZM9iUWYx+U7YtBdkdP08uTXwdht26QUpfwHJUG98We
f7YUzspxgP55yL+4LwjU/LdT55mQgCJjdFWyQpW9tgv20AKgMJ4NwYmxmkuivYt86QmdRUKpLJet
6bvZ0+TEFhORpk9p3CdqbS7oCc6UtXb3lmnYOT1a7MPyFlmwI7DbC/jL7hJn5kR8va+wAm4F6QYd
NKtHpWtTCKkd1IvPYntof77NIlTA3AaRWONhaUYbINBfCW2BUGcXOvfkzsiu3+wNVfmMs+Rw/2Wg
BKIS/BuAiFAlEiFtMg/fr4cl8RCK4QcCtR4igumyZT8D3WQ0aYzlK+thwJR9c1AvK3IQtzumxV1O
VTsPU0c5BjMU3mujI1P+r04TEt1Z89WO9hJfzgz8rRp0w5EwYjT56iMKgFHPxrelPgb8oT7aGJDE
8NdClALLApxOy8M4uxfCYINiVto1MWrDGlRSj1WIYeW9d3iWKtswv+1PVgEfQZIwKmutRRMccghW
aGgrokwrRTMF9gboDNGyrH37VJ4CnRLv1E3GMdaL50GhempPrl4SavlQ3h80QgmdWkFfEoqta8OS
HhhD6HFBJSAdVrGTObCQTP5s5xc4lhftpzie+fejAQMZoY2Tx3K8JB83/r+lQ+DZLz4u5iUP7fV0
fpwgZ/TOyvhn6weVZoWn8JJfgGzlTrMp7TkjBtoV3pDwhJv7FLJ+KO2PM6m6dnwMoTanGMmlqJHs
Iwb+J/ENwubRLrh1djEVJlXdTNzM0+rrr7SlcpVP+Gqpkc3dXZB43h+zXVfEdn2+kNsPgpWQqBOt
2nFS8pOAgtMV/QPpsqM5kKLULjXmgSjugzXl3dvsXtAPPQo8GeW+WgBTNAv/76lHs9hEZuykFDwV
sNRHgYfzDbhicT0gN5ctsSkcAou7mRzqmwWyqYbeT4BwcygRuTNPYWGmJR3J94Ffr966M3uJanMK
tUtzcYmPGqOTMzGo793iL5dUhGYQrKZqcB4XxsPRGaJgkrrr+oIPKtgf5Het8XOHR52L4zbwby32
4XhxyJNL77dJ2HSs2imuVHMiWMsLMBD6/6FqJey7z9bemDLPNmp/t+2+zVbTdOmc4tR7DNSlhbyV
/Ogv0qpVHH7aivuJhmT2AtiaQ/n9lYSW6ruQshinQQ2eHIK5hLC6A6QGW1+Y0BRU1ku+ETAXmTj5
V289qu2UYeWFrJ5sOsFrMUlqOhTtcyY3DlbMjJuoEjPJ3pNxfPjFofIcaVAYt4M42e3eLN1jkWQs
dXA6EJmRsNT8Jvci6GoLpGSOcvgOFjxV4BkPbKMCMwRWTobZyfnQ0KIWrH5W7M/rp7nPpBKE/yfh
Kyt9YPKpONfEFnbUKEpldp8fly0bNxEKakqY6wL4CBVYc5DpjAXK7+RwYvgc8/uG3tVXwF2zTkNg
QyJriXv2XIl7bs/5+egZt4gzI6SF1EiDSaSGrqmbEb9fk7NyOZE9WR7bRm9cQGddQKvfDgdcSC3/
vANJw2dVObuU9xlB+JnLLUxETkHWnz76AROrGCdlJo//I3KXqdABqCc61KeoXyXAICgB7Z6YBGCe
NR9zvzLAn99fLRLgYtrdXp8v8j0dwVb5zDhuXDiGSNKpeyNPqfpCB0B3jiOLe6OMXZC5lTNFubY7
z30AyWx/B1CaWTxRtKN1ZEqsuurNRJEAWZjCVIxjmiYsUnBFEJ8iFp41PwmiowPeMeiXW4WJqH32
Vf4dMlIDgiC7rbyOyqiNd9Tna8+MMYLKsAYfN0Yo6mH8HsWXvOWFkRvW+TFBx5l7fJt1owUAOqS7
9OZ77yzSkFUEhvaie9/ue190bB+2AbqBp3mF8qEw9b5+QTKzMhtvkhGqvg/rlIgZd/E/p0+ZkN4W
4yj+aU/TeOByS83g/ZNhzN8od0N/uohumMSs/pnWR1fJ8QNDrcdA8ZTD10BIObkK/bUHj83+O8Y5
EX9L3f9gD0Kx/7+ug+wHByUwzTlfw1uZxp4S7J7g47hAI4VLUv2RwLFY6mPexRDeHVMySXeDGxYa
EunrNN6SlVBO6UdY/snaIp5pdmvPEI43tjqExMuTP4FR2rP1GypTTeDWKPPYzfH5jY8ofLM5O4Nr
um0MfRtbesz1TplBeBPa1tx7/+iPKKzkxTOpOCtp5oxgiIEZADWTmeJrt4aDnZIzqRvPeQoNA0Fx
6JbKY+3AcOR9N1kN4G5dqb1zVA+nztKpWIUbyjxGaqnE58At0rnZvA2cFnK61Tpni/kGtnFKY9cY
pr9PDAkpwXFcvYArJjDNahYhQMvwEaZEqisxvmn+RGpe0LWd5O5maeYV7bac+bI8Se+UWYycZb3v
W+22bN0rsQ54BW3ZtMrq7BOENtO7SaJqWZ3ulvTZeJVfo8ET69q/emreYvtxU2c19ZKjAr3lDP5G
xWINnMt+1vbFBMddYLXwo/o9A5Z/jldKuizdLM//eu2CJHbFkk+0oM5a1WaSj8C3/oxg1S9mO4n6
qMhYjQPfHd+KmD9Ov165oRESvXGRgcC0+VtZRnHNR//qduGCkqJco1fDxgMJPRLJtQQx0va9Ij8I
HdtWCgEnOyRQPj1UIPqaqx5hpDRezKEbLaj9LzuuRJ6xcmL42DmCuF09ZWewkFMBjTYXTH2Ot+fL
xNx7ow8OuEgNb2wbpzW5pR7TJKo/8hECjdw9Ywwm1Kq5kcw0eNBoVZP5NzHYXEBT79nfPWOpFYRL
jABo69B27l0iCOKg7KEkVbZ3KociR76yiJn8VoOt3hIPaHa3nHAv48nXbDDzcbNVO+abfcF+Mwo/
ngfRFuHZRcCFM405E3ZH4COTCuwUAJQj4gZUzeC7wVeY29cybxZVMnpTzvmLou7WngrtnLjRNNL3
0yHKyKkLK0qeFiZSqXTvbLwJv1WPp47JR1N0Q2U1HPMGs4erehmiIifYFT4gzvSkP9m1OrydqF12
N0n03Zl0LJdIdDKSs9VxSSQl7E/jh6cT5Xn5vPvDOSjdj6mT7/RbEecVpuU4Icfk/0GFwVSTL8jJ
1+aCZIiNK0bGass0A19pXT7gckFnozu/1JB1Achv+hmHKj2OvZ9g/rFDRvGCo4qTKJsLpC3OVddn
D+776VpC7yZLzEmjeLTyn22ACN/BMZ5vInSmmOT/YfN1SlJph6Fl81YF4UJ0FQr6p0C70sDgIj0H
eNKKMXXrxtg0OkWPwIVNnNrRsS5iUoNdbPsG34h7dcij2KkKGOznKOWNtgx78HiksDuUTfSeC5Md
nacMvZ3RNpRfVn65sk8frCbpDnQOwy2dhII0LmqNqu0wcdmZxNxmkZqZOELADkAkpCgN4NM34IeN
1lObj5ID7gIhEVxNGtmtPWlGRr4A/SKcO/o1N+8+8lGwA6onG8MC7CG7dEUwFNSYs0DPQ4I+nbxW
umUK5umarszvale/oC/+UGBrx/o8XsQ509OWus0Dae9AtGmhuxqeh2r/9tw+ngTkbj+wJP83lSX3
j7MZf4b8J48M7O1Fjd9hRtprSqUNqaFBykaTxawSDu0iqqiHCiYKUgJxSHN05eJspRIG8qyFcTCr
jM7tHT3uznEmeQCDWKTz3n30Rh7R+2acOvyyrb3dtGiiobVAbIotCGkpVamoPYq4RSeEe24pPLis
sNgY2VlnNerT2uLrfMhsJ40XWWX0KoSQB7cmuJgN9urzYzQIjZnVWZkC0t59dlVElm6P9CT7v9tn
0iDpTASCYzJTzpt2sEcdoPCqNXFqSjFObzMcv0mGvXQn5BkUf96fNKTy+cGIV7KyVMyanYVDrdAt
4vMhB7cE7dKygehXmvMOVcXD12GLRUKPrdGuM9CjcGe1XTPjmSU8ctMw2rOSFUZqbP6IFyoxNdUh
m13ZSHtfV9jVZdfQcq7Z37QIfbeS6NJaq+ww8ZJ2TH2ebzknHG/ncGutBSLVK1crcRmM9t7JxIh9
UCzy/vI4KPZ69jGEKSR5FDfWWGpOunfzutdZbEcLPdiHsPiHz+cEc/a6oHNoEMmJoe+yMKyyq47r
LGEhVWedVZsUR3DMf5SseKUJ1WV++hGuTXBkc/cBkh3IqST99Hn56Xl6ytzJoBpvK+cjkThpqw9H
KZtf6AdYyffr7z+zKaCmGb8axSZ7crrgXIlmTdnfgPJ9b/HpO9OPq3mH3jz06r2erMWW3LQi0j15
XiOB+epfzNhVbbZNgx35e4osrLdVNUDAZbTRDexQtj6i8/mYhDn/2Y25ZfHt+oR+GSmqpnpEV6zs
S+X5YiVOe9n8yiwxk2hK3XHCmM/3syHdK5hDOgvIr3BM1OlcNWscvkFhYOxfoECLnifA3Kiz/OsR
32fzCSNb5PWcqJXIXJnuTWLb/KTBTcuUEiTZa81oG1CKzyuqUkB51TOl2YFbR58n06GRWu0KFulM
g3A9q/L4hfplaG6vI1qa8HGw422w6VeGUduQEc73OVDOnD09ZvqBO0YQoR02k/MsX391dqYpR1xQ
17h3tw2Ey2jtkYZdJQU2XKWFfpQotChBZ8YxvterGXHVUTtNQSJIv1GCMDvNwYzBniw8JIwyKiMR
NCirU/4qq6gy8h0CWnmzY611HA9tLzHTFl9d+Z798Ks/lu77wVyWefKjY1YWiuaBxoRecLGoDzQm
77Uk7Zi6l5KFpwUltHZJyQabKo1nqSMe4W7JdbTwCbvcJxj2g4KMEPoej8wlhSYw5rzyBvxr8b39
2vYATAjhJu4M4GAVA4epP/pC7HvdVaUtM8gXj/MAtUviV4MEo12Zl1/st7zdR3jjvHk06+6ydVSJ
tKXdd8BvWo1v3Yi5F6rtBDqjeUp5owjawtrNGIU6A0a4fTBevP1mp+dv5l9GqAkxNOYcrr7EF+mT
CW66JMnkLeNqfGB4j0iaLhf8J1nP4dBwzHG9dz0GjvwjWMyaYmAWCuxt4RA12Fvh06FtAjXjSKFw
gjPngtdbLf8mFNivP7BVxWXMXxcItw9cWH8Jdv9Iz4Io9WeFEoZHUplHekQVIVinPKj3powLasR+
F5QC9WWSEeMicfdVfUQm9amePgcwwvw2gdh8wpwSZ8WkcJaCsUp89fvP3Px7X6mGYWrM0w/VUncd
fJoUk8PXQVFd0ThEzAujKcI9njd6UKwDC+BokmwbUQQsHoUYjQN+b7jHGJeiYfYLYqvLFTJV03lo
CM7GywOnkZkmPaPMswYJ1PFki4N1oTTMOKnDAEjYJxMgBhmeSUAREWLsAVOb9WkUnsERzYMjR3H0
EhVC5tY4biXpItgTvShmJDrSRa+O398xRq8H6lSZScFMk2G/6qiGbaK5Mr/dkzEew7jWUGMwPwwP
u37ffwUOsAPGuS0zbJIb2i8UzWudGWDgz+4bctTus9lN2Xs35SpNp57+rHSYeSoWH5Z4nxe43VmD
DenfRZIr3UjZScvX9zi9kPvPHMbsX/7Xc5rdJG16wTfjsbP4va1A6DZnUpcbUMam66nq4iVjWEjb
StJ26SEkSGcUvpESrtsfDZpgS623CFjXmeh4J0J3VVjSo934e3o5Idobx5KxH4054mbdzfZFI77g
i5X6GK5aX9o2KoLJOCaPADc4BeDP33Mzks/qRYBC5SAfHOuj7/GUwTroEdiNvDSdBzBsJPQ8E8SI
utxp9+TPCjGVoE+v3Zr6ya0Fuc9/BEyM7EnSXEKnbvN+3W2a3e8RIvKerRIf/oinlEJPsThphTCj
mncHE+9OjVSLzjQv61vNSsN4rfwMUh866U/ZxtydYZ5uCdzO94iEJ1o0IHJSB8zEIkGSsgZT64Zp
vzDhDw5b7SmXl7dF8GWvZ90GFeqN2GyLUXBmw2liN4YN3fOexzxkrmcvxgI8lPvmBAzrMUPezDbI
VY7PvYYQZMR35WkMSc6wut7K88Ngd8I9RWyZjrSKRoXUZMfJ3LRXRSETYQit8q9+gZgVhk2zcXpr
NzqcYm1BHDA8N4ZdKp33dH1FQpJ/ljXRR9qMdq+zALcN9jDvPx/6RcTSS8yrVJFhut3Y8GcjZqOy
jjyxSlayEf7Ill0Gu6mTknDVAhGCSZIB/N3fw0exwWsgR4jP74RItdjbeXr/p7qlw9GYiwWDpg0f
TQBMz437mkL6p4Zx5N8Kpeh2cItiOZPY8XizpFh1en6D3l8T2Mj8gD/YmzHV2ImxiA62XjKhsZw+
41+yBEZ5CNe/ng75yWBkQqzzs3xbSyf+OAu0OedIKvQzNvHZx+ovczs2v1C8cQuqmVrMNWIIJp4O
0IP6s+KZA9B4gfDD/yTyHHbVKetLV1x+oXsh4JefQikUFuBQFHf252hpnJhVZXH0uvA2YVxs+WOc
Okwd49hL5QKPiSBs6K9tEetKef4BNVnwyxiUxP+JXMR+qziw83C6KsTj3+4YsJ8ppecIsenj38d0
gxOGVSal1NsjacbQxM17t024anwSupH9QSI82Vs3zwsRqHi1PNO9uvx55j9BiCrcqJkDqs8E9PD+
mQzaDnft1z8m2gQF1g3I+3wnMhemnzV8UchoZ/8cqcklWhlxBTQX3GaBmJz2G1SwA9btw8Vo5Qvw
l2DbEDEQemS8TEbti88GPHrE+guqz+p4W3UVOHBsRTspg5pg1e1fT6mBIEZOPoU3g2CiRVLPV0jV
6y+2+AeRJv/ciLL5ZRBD8LWa8hc/uUKSaOhmCQPUnugdgpu4rb7QrvUwMRwh7WuhkBpX2ulyFaqQ
t9rf46yyoja/0K/TF/MQPMktFn4ZD2HPM3Jw63FUCBIUhlmoUBS7ItVhRDllFd/zdECrURRn0Ons
ayMadDFxIkR1Jn9jkQxO3PRGftpcLXOZUud7O6awOsq8HrIZlIkICGN6QmstAE4pJ8w4mOaIAFb1
mOuyP1q22EM4em0UJHujpQm4t/XJKZYFbZDX6aqFbQxBl0XeW89hlFcsrdfXM/Jhzo8GP4Tk7NK2
ArF1Uq36dmO5GpfB6RTqhyPxLD8Fn+Ei6oy9HBXOtUzDNPvEVk+srou8OKVIQSoH72d8j0AIN94y
b+f1zpF18uBZrsCrZU6jvHy3tNiiNpKV7MRbU3/71EwZmkc6Pfr+mke7cmpTTG56KLrnOoS8aZMz
YBChMQUf36RAPs6JciZ23yAAYxGbzDW4tWrvKFcWQjED61wgdEt2ksXwe/qdg4fIWAHREuQeP85g
a3Ir+5ZovB6tQmmcUeOBCJ4Z6BdHyCDEioxoJ26kDoVigMVQNBpJ0/xp93CFUCybKNoMIr8i1I4a
gfzHx29O3xqsi2GEJk6SkPL5kkcA38xTHkQ4oTYizXGJV7oVqBhGy9mGZfeDkAGiUtHC0Rk3dRGC
Xyf6Q41qvfNkCK8VPmtJtsflAylYtq5qgwe3VSNGl8PNJ6rdBZcJGN7MmsYz0F8FId6U4O3H7GKC
EbimKwo9h2F3FAcwYuJ2fR8o21TyCv0tMhNec5SHneDWRN7ZFN+2dBiaOQsUnZbWC2TFG4KR9y3O
bAUXWGs3Re9igy9q08gZ4y4ez7XZnj7GNgaMxIU5Lunmp8sjTxDxzncNnXXtO1EcToqM/v+oKNbE
2vc9WcN4OBQM1rvRF3D/YCGQ7Jy6DrpGWiznAv7FTBhTwznEjn0aSHVBM6eLFhnp+mP9OWgS4/tf
f9sWnm5wEYxoUaBaOR/ihH+mL6vGWg+GsKhpSpkvqn5k4l7KoxAJTINgVGjKEYC6MZ1Xjy8BuGZY
a2E+1JVX0GdACMSJbRzvtnhxvINAom9padC0ZXCfWVv4/Fg61RmU6q225Q3whpJRC+6J6CYEK3PA
Aw73USAUWZHHtDHgEgVw1QbTjF/qgWrlUskpnWTD6XJJ/xZunU+jynmnafHf+qkEYJ5qY/qRsXPs
FA4M1gm++QQTMdB3BRyinR8h2qmmLDoCS8Lkf/2nck/k6AssRkdIYvyeV7+AS9UsJqZ6ZkPxx7fL
IrOW6WEE2VKoiX5wHHEh3xTm3SiIF8ZgIy/wlRkmFjm4SyFJPGzGdvab8czr6xDFF2tgp9lkvaoY
cBtV6dgH9iN3dkgHipxpfA+DvoJ/fK3cxCY9x8baanqC4N1BTjjBbgwAEb7KUlr2ChMPHWwzJZCc
r0X5SS566c/fLnSKcBskeQ2yUE/STyOa7fzeMjHzY4eh9IlVoj+ESXDRwvNwZB3/WzmbCq/kDcUT
LaK1HSmXj5UkiVOJKLnHYtBM9cumMaCgbqm/mf3Si5Bdhc5T1l0tWOQ9tdV4JFerqO2VtUVYDCZd
xxjzgiaCnOnSaWHsBkvNqXKZcB/ruCqfxBNeFiwd38oIsCPSPxInoj9QUZel/gTSfhBYxXndw5nf
t26fPK+mp/TeQDt0w31SGbHX5iKX0BubAVuCapVH1flxUAXm4R+ZOKSJUVuzKxau5c29+39jNCly
3fV6BPZrdwpLestGtCl+sv0FGHYMRWnNSkoWSnGdKYDylEU3bODIK1t6rhbWjthDfNbHrnKhuB70
rONI+Fqdec2zm2Zn50UfeRMI5nvFkSJbXYYizg//T7UY2ZrV6+PngJ2A5jjkvFB6Pi+3boVG2WN7
4Bf+pwJxrdi0q2nfTXxkFHiJUDuuU/CuacsYoicfdADYgnt/XR6oBG29XzBcztUM+axBpCeAIgku
7mnhL7OOoHVZOKheKzgLCxn9sOXAOXTtINd02DAeTq2TnBIh6dexCSueAcjMB6oiOWBh9+YAjat6
JXlNuWSOG3c2lFQR9sXXkAZgyHGhUXD8f2GZEhRAGnAl7U8I6r8QZT/nN2err16TKaKDwjU/uSKu
DgsipVBc1N9n3FAyaK72pXd9nN+lp+bCuCcezfVegl/c+B4lnh6BmRaFJztKI8mtxJ//gjYtlL/O
bA1muMzlt/7qE4d4yxYSLgCHLbzuoK3HIjcre+5egWPgPy7E5dHrvftHhhxr807dgEwd6CSsTw+R
bA+PGNck24FgXOyAc5RCMA0Hh7qGyM/6bw2d4SZvXGnvC/jaM/8y0V3VAsdxy785zoTWLqj4EhpN
3lW28hu0dYkfMOs8cgzXMh6sxtkPpF5IeYtPWuOWz1DO5XApxlbuOMT9DUjHWmQLDxuzPxOSdH3g
KOk+Wq09otEA/bhBPTOK45Gm3o3ifJhv+dKMtWVUaPhDk6q+8aPsBicjYmILb0ix8Hm2VL2ipLvl
JJpEDThn6c8xjbEiItM3e8wkUz0no0Odzg6sYW/LHGqf/ojE2ilIxPYEmaOKfLKIKxLkp48fRm7X
EtFc1aRZuY7HB7kx80GzJurw5uFRLH+FcRvKY7O3jPeIsiNxfbcE1lQekpMDnVlzS2dAMHg8Xii+
RSOmXk9s+kA3AbI5J9WFWoNblGBc65uZ8cCQpnI4Es/98fbu7iBY/eOAgCegqjwriHXDcyGrBBcC
AHGQ0z2h1v7jY9aIC8VFhI5jDHAY2ixXkhv0RqyhTlOPvHsIN+L7W+fuaRf07vF5PRAvw+YS3Z9n
7RZ/lANJxet0Ukw+qojoPrY03k6ehhly5ay0lNwM6pygh4pl+yK8yzyS9RuXAUHlYlXtkmHWLMsr
HM3HJ4yIWQZfm98tXqdiz6lese0RGf7ntQreiSfTCfipu4oTO07rLV4X6TrXhTiTbPq7roSQtOtd
qyari29vDOeekIv9X0q2fqWeV5TLVGcpaZ1Mdr7GIOQQSwxJJGEHV515SFbt55VJDAi506/EJ6sX
XQgg9IeXhhzZke/zEY8RLCy82I6QfgYDBwJ21u+AktUhZP3QwfkHls3JfHUe0PYKJXZubcPcBxhS
8zJmeaV6A1GRrvhBNtBygf6pVmUMKl0NWboB2H9hIDfoV5sVdDCbnMDw1Tjt48Ew9d0bH3vZSMov
LAm4GGfFCOWK5QFjbaxcfCia5Xa7AvypGqMIYZE/Lk6zF/gBvre8Y4975Kw6lKdKOntZ21LLgw8O
VxwoKtYgsUbi18eCq75U72BAWFZpQ+q7UQNfoJ3PA8lSZsnUlKCF1/UaEejn5dFoUJB514K4IaM5
TVJeoPguEhhr6jkBF6XTBU9eXpE3k44Uz/Hd5WHTlW0MtctVJiH6US/W3ENDwYfS5ynckxDXtWAG
y19BHs1/PBLam8ZEUc7iSCWihM46Qd2+XtUhrdPjTnTG9/TQthVbfWznr2qjaVrureQhMi4Gluuw
gOEuZ44h+ieN3FFcqKjTfBLNZJ5MW/X+KTdgUOCMpSyQYElApiX/e/4vlt2c5tq6onYCDS5Pj3J7
faUyk6PtZpl7Npqysz8RfQ5eGcSLwmlM40duN6++6PxjvL7OcXCoxLHHPpDAC5JSKuuGStGDPxEd
u1/Dq6rpQMlS52i85oWx4FcoHxcbsFc7WJERjVqaheOy0h7EZk1PoAGFDgoclvTxL5Vh0G+8lVWw
I2OUbfj/3DKIn0QQfoVkSMrZ6Gha7WucBTBgsRqwi3x6wIkSZy4HJJEgNq1U72MYSN0ukRkCetTE
WqKbxprK+yALws+u/wMJsv8GuDr4QhZ2nPi9061tOyYmBAxEhetyFoxtHufhwlZqdwqsjOpFRg3q
j1Q3INPsnTte4Ftw3vtEOdgPF9nmTIGnQEMKNOQ2pFAn/1D0yXhFqOpFgMgcXwq+EbjUrc9u9nF1
NUxqEMuwCGcvKaijHmHumVXgNNaHbrYxoW1IMUt8HGbYYmfSqL4NnRTJ/QtusC1LOxq/PuFAEY1q
fycGcgZgExsrPNDwBATeMgn/6hX+cgyZt+BKJHRAeEoVLNoO0lC9n8WB4OxN1UKRZQHTlrzGbq5w
W06xzmvRD67mVGx5oYsxKJBATa9n3ghrsxBMVcWRDKpIEPLe4Ol5VZgyAB+/kiBDf5AlMQkzkIjt
zGTUII7lLhDuCC2t+yxtd4kQPUkwPZ+9ud3qXzshch7MOSx/w/dQ3y4YpQ63z1S9PonTC7ToTIXy
C5T8/9vRJElYPTPg5n5qmg6Jo+hZnGL2+sbeRgQCqj2NjFGbeQSAArpAMqPyI1aOAdpA1ME2Zbd4
iVIrCp+2q3ktNBj6bYINNbxxh3HsabE7kLgnjZBnGM463emZAy7tt7DXmt/fctVBz0Jrjwy3lY1Z
AYiQDlpl80ID9vDeyXqI89uTbNE4+RNHTNkeRTMG40uWPqiw/Ygbf+QRhSZ5C/JmKKrq3l6lGshf
cFcharD/TfSs/B8NsPBitKcrXTbP5Qik+gMjCAkujB+YPIrlEOcSrwUl91PCeliHIvuvpn+Q5DEi
YHWlziKwCmXNRFzTC1iukOTyBiomDBvVx5KjGN/58fBEMKxYIkBOECrN0kcehpoobZCzhHQYKHFF
u5k+jAn+cvj4AhoO/kziFsVN4FbCVZjnK/R/8XpzFPnnHyRltTPQay3HAvwbIR73M4gBWmjf7em9
XzzukHiAiq6dbIKvdi/1IY0DPTuPQikMp+VIj1H5OM/YUP+5VTe2OwFIsU5OVx7en5OtToIN9ZLc
CF3mdWO3ggT8Ew2VeYbSqOxii2TvLwoDCG09/jkzW2rPJmB8lfXhsqAjNPHwfFcgl7UuxpU23Y75
wVhzvo4ruXMpgtAPyvURvedFwpX+NW22tz0Lks9sMEWBIIxwMkCfbgSuhlR7+AEe1aiJJ78ZhZZN
mVwPcQr30+T2vGxIHybJYwAcWT9eZCb94JHqRly44MtZPLPf/PjIL0/HzqGi2xog7tCfADrzV9cP
Yh7ZFTj+6ych/Jgs7wdWj37QzOVQsxbUXVazJHP0w6uUzzF7Yc/wB+A/20VIBU6GQDCVtsi/fNDc
QZGKxmOiTzkuXtWfPyLkcVExqdCd8ch/U6DruRfKhs//qCQ0vH2p+wxmHrkBA0S3guBf716h3hp6
a+VeKlxXN5o/bPoWWfCMynLPqpLV5z7gKap/+MN8s4ur0SxR6qIqwDEGMQgiVmR1ELrZCZCWnnzk
D0T8bNLwiunJ2iuJ1bdP2aWrpcjjOkzSlumtwoMOctFSv0aF2lQNB+EEE5A6FBkUxGC2A8TBB0M5
QNFjPoS9DIq6sqpYynYASBHeAihKny0bLz1Qh8ILmm6vd7j9wphwcUGsDvWwD48TfEPqxQdGv/9E
v0XfKGe/hpAPK/1Aty+STNhx3Fd2P8phLba6CpPjl0QK3GsyczItsTUeuV3FM0f6YTxbUi6+s3P6
ttwgKUj5MblvQXHNMr3OT3MaeDkJq4kvGcAS93POjKhlOSzLhXFhxDyjffvtIWswXC6H/p8+cS0H
LmAVsKcWZd9Vu8DA+ggptJTgsvioKi37AR3DBdLLKuhwj+EEg2fRoA3JhPcUlx1KYSIK1UB7ycBC
QeMRWYgiOCeolw+jUS2E1jNTRTxHLiGpJle87Zc0po4uT3iP6cK5C8v+SBxYU4k8vQ7Nhzs8f0ql
bK2UvCg0aXN3uc0tLQnzmDfXcFL/Zjyehlrb+W0UO/QeuV9PuVAXe1ylsGgrbroDEZQfllqiPEqD
3U6cSt3YyTe0XOZ1GsU1MbGNSOPMuu9GuzCBUXB1XoaqClKvLPZXDog4nr5wcKrYooZ5X98BLu2X
bIL7l+RnmmBne6G525YwsU1UwkPk+1EIysnyUlovbUgjCB5lu/VNd9iLXF9s9TaSV1BBJXyAxrTZ
0HHF3LPlNlkRhP8ScFZ5B+3P/lQLqqv6WzNzlBSGCHeLMQ550w7kSH4SRWpR4e7fDGbstDSDHonb
3RcwcnPHhIQKrG7FqfyAaiVMeQ4UlPK2qiUWTD75Vp5i5YpC1kCfqdCrLhPGO0WValQUIAzj5mim
vqB4DbYM4I/UsOb4otmcs/nBMu98wrX/m252C6cM409wocO3VkN1bCJofQSaFbpgAYX4eq78xHN9
BNU9gPeGTIju9STK5nP9oQ79x/sZzN8k3dTXbqjtbllEs/szHW09eyvYRHQiauzcRCNpspujFc4y
QUc/7iWVEg7VpksOASh3Qg/7bnfzgpQ7gRt9bwFjg60vxHzS6+BXJWQyWeyVopW1W9e5XZ6F2nu7
SRRrncrE4zswHYAQzKwrUXzDGPRpbG9g1+OoQyyZRrJKIWYnwRmr7uBuAmDnBtXELnEFGgfB+Fhi
EVwLz/k7sUTBep171JBPadu0YnXBhKs7v0EjUk2tEzBIrNyHnFHcvd0PVUI6iuda1CC+7FA3PqCU
mbSC6kGIecZq46077Bt0C2Ss+DujJ7J9m0ICJjRY85oJQzIcbllW1PsWX7H3OWJ6razFhi0TpNjB
881vzN4hIYtCEPs1JwzxE6gse4BhN4xO7O60np35z9swG43QD2UNGUhpGC+iYL28ESpUdwRDNUM7
N8fNVg7dKdXdLZD+/ADOSlNoi5v9BifYzjyYNwxmVPfCFT/dvqvxX00lIGmXH99TmcweKzXSrymv
OQpAyuxrvyd42VNMoF7ki3tRAlZU2BvQPsaTPmI9W0JNPwEoIPfwwKC7b/gG9rDIAQJrDyTrFx4U
zz5U6o+rf+RjIfCgwXmI4HmcLrnXzm7+gV5/6QiW17vyByizjxAH74/eZsX94HwcFUg9OjMxoXxQ
MsVC4DRBmEl/f3c1uH22JF0fHMu0784Z3V+ZpOlokHFGmQxy3WqnuyabWHnl/QWGCneu5YLw1Cho
2Foo1zRCa9dCXFMDic9naQrQs4gpFxW2sqkVdydH/H04Rom1kK86Rvo3RyqWT6s++QpGntNxGEDr
cdglj5yqDoXsndEaUtiAG9wQ35fLwMboneOVm3wbuLge4tVwNUTUuG1aoRloBVgtRJK6LON6yfAe
A4VHFMP4pW89eE0gTWAlA0VAAPMzDJNOw4itWtb3LBIN3uWmVTtw5xD5qJqTPiSp9e5pBtrDNX8i
J/ZsrrvoOqSuWYEabMc9w7AFWV2YSRatonAhGTmH/1hTZVfbbd/MMB7PeZvGskRZRJVmQet1Rpag
YGXXgMq27QHkDA0Mh/mPsJoPWMQ7Q8I0jMEMujZ6OZWC6/zerHZ54TiquNQjNcBOLDEA8ZgtrksM
795mC0PCQp12w8zOtDgftNH1jnk6qPTUf4FoYB9ZGJ987nz+gH0o+HaFaNeyszGOGc11xOF4wXRr
ho9heohQYbMhKM7OJzrpsZAfMRTAl0lHzr3tMtl6lDAWB/jZfA7DxA0jZng/96HPFzK4PgRaVbxF
lKZJuiLV27z2TL/STrJA16bwmbZm0l4a86RsiYP59huGZTIlIIpNRA2+XPjL+8e4h2Hj4yZkanIc
Sr1YYXz1Bfv8+FIVJ7yI8GbQiEXjzsi/vVgEFd3evIM2T2R21SJoITs1AWeSyR67kBff4KZHyAGu
4TooVVjRj5feqfmhxeZxI6cAohVtHT39DrR+8IDaA43n1bzQJMk+RLLUqXp68NeVOdRZOR9K/Ndn
JSKZSHNIHtuYO+fLBoG+ZX1d+Vo7x4fUTf2PlGhD2zEV0VSKx8ewopAF9FVJmYj1/qNt+2+CMCrG
O9CAdtChCAcN7n/L2MKsc5LL8GUky6KOYtJRE1uSlDqert8hTxsLbAFhmyo9i4VsI4J34NaqbP52
4KwJKB4WqG1KByABsE+2FozUP8GoE5zCls+UqSsQgo0X9hGBF1mEjvWA/B8p/bkaaQMOQxyuD1u/
hL5XbEEvC/2OmHN7c0wU9jo9Mbc5HqpuC7wAsV94sUafIIOXdyWPdZ96ej7t+DlCX5vcWn1zPy6P
svDTrHrpVzM+R/M8IX82XhJVnBEkXLWLX0gHMXmQsP5xCuY4dgpclL8MofhCZroKUogsaAg+Q0J2
QtuLldbrn7+DqgFWLaPu/wqt5sXMCIZLI/YWlWMRrc7UyWBuAMLSeQrOV8KBJ3pbmQIr7kxMkli6
DU7CMIyaRYa1lIAq3THlQK8EsnP1tHKJE27Pxm8CqJlqQgGlFar+CrHz5GSvGa0ToVLeRyWMrBMW
Q1gGQTSBnAW3yZi4Mb2uMoCah00SN4gaYv1+Z5AaI4GvjNkPo13mNezYk9LcUeTGahWYlmGGtxbM
WN2j/6bR0Myp+W/Fu+T2pRd97DbHipR/HM74tXcOUfvATe5f+WetocrlfB2W6lb/s9gZt+BSq7jU
ll8tkd+ZPtmkUMbsbHxSOpBhopBH5GCqeyOusQKqilOYATLOvEGDsem8JKlV6uYRKwmfeH06EZI9
pfCZLM78a2RLHy73oD94SXhwuwW0dPqTFuFspvariDD6EaUTpmupx+JrSeNDKPylDAUg2a9kZi0e
ww2KzlyGYN04glrC555ArR2QPuoHkbuSdKkcByr8s6uYYXbQpt9Gd+o9vSk0fqZPo47x3JuRAcfA
jJ0b3dRghtf07o1VLxK4CQsRYOx/2OQr0rsFSfYgrzw2/WGDxNHyxgY2klSqMJGPpPl59WKDmT2P
mXgwd4KJ8pOpBpgX4vqfqRQGTChr3Q/+lb7FhX/NwTEUMOrcciVzw/tAL8VcqJKAlc9szYeMTvij
bv93bH5B3zyAQ2RdByjhNlqfSm4I6dqDnCZtrZdaXRi41EOgW9AcYp+UScpvRDqgdVxEfftQOGCi
GY8z2DJWrUPBc77RYINsI5KdU7cHm8PrCMxI5zh3DlpRt/AojiUMAr8xZJXLctE7FWZiRMgqL/W+
Q5VRJV06XCn7E0WB67dKHQbBuAK3IsoprC9BjH0hFb+cVyVL61yHM2/mth7p59hS/OwqKGmeHEt7
49OWnk8kAlB5Zr01BEYX+uahE1jssiBQq1ZkzKN0cLVgIJ2XItJS5f8KmErFEWtBCUJS00QBmDxK
0+gHpucxIwtJ265xD83+xNfeujl/7tyyhDG9k1sk0eDFj2bb5yhQirsOPWNpAoe/5Ky9pzErcPyt
oRJoZvWQtBgFGJVsLu5SR3XdEX4LT9a9wWhXhvfvs3+3X8TYV6JRCC5i2Re2/MKlJmk0qZOX7qHu
ek3Mo28iv0eF/8Xf0UaooWjFA2Q3k+24VgbkX8lsyxCSmOJ7n5XQKWFKMsbXRUPQwDNQhxlG7CPt
1NW3fs2Wr+GqetiuSMbMW93i2pUhFc5GAQ7NQ7qOlomGJrcScICGZAn99ik9AbDZ6AkYDZZ/hoo2
cDNmseqGGmbdnZ9CrkkayOOInY4VfMVTe50sVTGsm9Xk+44jbz6l/L1SQO4OqXc3aUxSoVvLplbW
Yn/OYBLn8pO5omCwjgEM5gz8D8an1REkhEp6yP/Huqp26zjrGzHnDiubC0Dk2H9KieCoVYVGl1ya
NED6PIs+9hBTg+fN3mSp4q4m5etmmjLYTTo0pDffQXoGg+zzEoXDQNRnQbVu3gnLRDVFd0GF32oB
Gz9bYszkN/T+izKuGA1n4h1+xBDh/NcL76WezbO4eeKcRuV7s8HCUqPZ/H9XHV0EGXqkj7o1vOZr
iorty5PzWe1H1v7ak3pLHo8NcasXDwhbQgbyJ6e6KuohWOLPfjgKWmMGHJvyMof7E+y5oHMGyp32
R+V+rxvJnXzfvgP3sSvc87sk0zfByWyxTFtCfiYvVpFUQQS+cob7H3xZ9fW1vJV60aiESsEQW9s2
gsKJSO7KJiVfnUoQVhcNO7PKTNHtkPOAUke+2hfVJw6YS/0oxB63v49FkTLY1XbjS/bL/r70oUXX
GsYTOpF+3d+Wsq8D1u5VRZVq8OADdtWufnbVe6qUteRo+Ni3LDK2X9B0UEzqM8IhSeNjqh+9e/cj
AmLNx33zWSlZeTchO4lITTXcZxVPIEVAC5MPJsISuEk/tXJcDLhHwXC3vV0KaQnBRFDWzuSASrv/
QVU6AEhV/UBYBz6h6OBY0gyhTfNm66lRDsztUDPqIH0m0JD9TJj1HV7X4+voOb34wP7ryq1+sXA9
e1W+aFgqJ55iuMRRHUVxsd/hGa28ILKO3tMc2L2FGUSEnHtgLYaB4LRpJ7g8n3MTjigI2dIRL97y
YEpAUu9xRf6EG1BLtGfyR32ylbjE25lAQnMkhBiEkz0hoD3M54NvNyxSucTWr7M/11Wl9p1kYTan
peUkHpg2biMUtsXl8tnCmMtF9Rl5sQ8QTGK9P52g5iW1eVMa2xUv6NGb9IyxeL2V0lOiaJzl30Jv
srrrSa5vFGHz5RLLNCi4IhmTnlyuUA7DrvJs+L2gh7PHoBqZR6X7faPJNRnmcQ3H0p0lTkjTwW7/
Gzs8VACkUHKJn07ZPh62OGHBpbgfkwuX2kIxeghWFBhDJlS7D3LaULYSP57vKoGZHpOHCiGqhYaq
FnCIZUwwFAb3lEvi3HdvRW7sHpQoYrj/S8buQe+g3Q69Q+edBpTsOzLZyTfkiqhXgW9pMKmHgRsa
Tm2bg5t5kJmcLdz//yfXdjgysKhaI30HqBcoXwHOsZfSAcrjWguZIlY8QhIZbDcMSx+U0/QE+2dV
qMPSx+e16OkcCjZlngvo8Qulw86KetKG4Tjl2NjAH8aHWsiA9c/bgmw1CUXgzDENDdKUol7c10Di
grlmBvq+W46cpaAz3mZEuCBwuC0Y2clPRUCA6+jfd2ntTcE/v2XJrpd4qW1CAR4wrv8QieyL6Vqv
wjzAz4nzGNGuNvqfKJP300HKlZme+bZZCezCUgDF6aNs+IKWpOkx2IxDzy2xivPQ7792VLY45qpI
0X6Rwd1JrFu9xrcPKj3zbruqOLLIqZxepdFXX9doB2pKC0agG/dWsjtShOhD4s8PkxdWUcTCxkzp
XszHNgNbaSOYvICTciIAkEAeuKJzgHbsgBnbQ/dRaQ7sXaeVNqbVG6v42N/sHS1wwrVdlV1gfVZM
xrXcPSHY0weEFlcwHApLBy9s4ZJsK/uAcVel56n/wWd9/NSxeb51qM+ffy60y56EZ9oHD+YTtnyx
PnfOnvUHs/Unp7YYgQqvyKqXH4v+z9XY0yTjKHwfVOgdyhYHjW+lSEdCAwwk4qD94Nd06u79Prnr
GqA0q9UmNPa3u0yWRW1Z4q2NlPczO1ifFkBYzxCliSc03PQTFb86l0Y7+bvy/CwF6T0SsXWArt62
w27qFoN2e2iTeYbHXEbnniYzOAK8zJf7ko7DyyBQalFWQoszAihErc3UlmOrWSi0ibQ5IdcJj4Zr
00GuOQNUbNlOgu3gOlo9RdbPEOpML9YrA/gq1Z5S+zDg5Ya4n4coQ6OfhkqjXNWKULN7ayQarlr8
GTYCBemCFp1DrvKiodOP4DV23FisPhSIIybx0KAY+Wy5sXfvo5Xew7CFWudL4wPXhT2vLZ0HxeRM
ct1EKs1ifiG/0vWnPCLzg8oHrKzCxxH0m6zeiBhzJAnNgtnU1R6xWWq4I6H90IrznFDft0B/iouq
xWP58pkA0IoUjmLrCUuBD/Yj31WBfKrG/yI/CmQznCELmucjpW38uAAGJDZ9YCfud1Fga9DmmDX9
SZ98eJR3QwgUgAu2O4ddMdTOdVT/NbYwTWpT+1fmWWtSIG7v1Jrg9Hwjl/OaIs3iNb6Y1IL5S9W9
np9bHyjHWPfSXY7jFEmQZMX5QtGkmFmv1MpjGudS7Hg/BCnvWwm41LBenkkS98hT3sR/iK+zyu0A
In3vfocceM3smra9QT8EB1e9GYdFaJpr92L3vSlygfRIGaxckeM3vd5IPvC8V3/pYPcE93rU+r6q
W8NY82bhA9PJQVLxwodlqOG9giYkmVdwrcy9cjBBrFVuKgrQRRfE9kaYGhDpWkzXW/FM6+7SSg1M
AO44A7Ky8SvJa4LdjLb2XiktRvg6O5M4e90E0bJ8GIrzCRL++fSn3ls1d9j9KAu/soJ9O9/OQfcE
tYmDNQ094WSrqUmo4M1dOcq1NcujGPDTGASEUOmsNZJHqq87WI/NFjs4KLgOlMFVfC3HW3ZwBeNa
I1vzsz2h60UQ49UIW0mzWFXQ252wRXzIuMKjRCp0b83gcaXbPT4i+wdmBRpZDUbxiNFnYnVxrGXB
tVC1Ya+PrTTZIwA3DE0s6ur6z5gfcHsFP36jOp0xT6JilV+azaMWT1YYVqgT72+8OXeM20VyHEza
LY1dtSMeI77DHTOEjzZK7nSxhpVCMynb6Sc9Poaxs+e3BeFdI9+wZocaooM4fhWB6ngnKPxI0OnP
ruWynPQLBcPJineYAbMFsvGpnjwvB1FFK5xvE7pb1IMSaEmRmLDdRclYo317nD1LTZzeyLPPmYLh
Qa7ojVPRJof0AuuQ5iOBbu+iMGBg+j2DGdLkaLuTdjpVUPAiUpAf4MoH3zeo6i6KqLCr3Y9M24n8
J2FUFmLpUkNKicPTuArNz7pSUdBCFmOVxnw3e9GK1Bgr6MpY4odvH+e3quW/y/2SaSBti5jF4Ia8
4GxanyoTjzp3fdo+uiWKPGDpo00MXdunBUhJNLYzA5kCCX81xts/sNo/HU272K4+KJnlrJ4t0jQn
DyNHtwVslmaQFvJs5X0i2jKaKX+Lt95cz1IzaCiVQwtaA+e/jteiBfw1uixxvFi/DgZj4oJBNQ8g
Ae+yg2pG0LD0nWWb7HH390M0K0ttIpf3DfX+x6cn2IihutD91JLgMXv7MkDyNzu4IXP6N1Zc8tb6
ctIH0RGcn+z4Zv4IT6/oKAbvbSitC4R2O6s07y/TvvAJTC2zmqX5qzBiH3f+ewwH6LTE6SSKBKXF
SOEgxAotu3qo623HJ1Kelix95noPi4bCPa6CvOoL4UiIGDi/gcGSrYL153Y2b8dUK/DnAdQ8xts6
muFIOvzyZ/kzTq1l1RE10bScFjDknw+pzYtMqZH4TnKJAabnuwJhS4Sn/kVqb/wy0x7dus5IXs5K
v3t8ZcBb2hdu4j+/4ARFs6czs1w5PGQjhCNzAZaqjA8pB5WecZ8WBjks1v6N+eXpaWZYriZ4/4Ko
4Y0bhZQbujy4s90pi4i/g2YFrtmHQuHPEbmn0mMXJ/7Zw4R9tFmGo1HNvKZXlhw8WS0WMHeLSok7
o6u381kqT89NoZExHAfDRozEr8OBHqkecTzA0PZbGxVi7KJffFpnLSaelwzDB1gJaUMDKLemSrdz
ekSYpiWI7IzqAyzuGb7ryZkZIwsZITJe6qhA/KK/8dffp4fdwvM80CuwlvCgMTIYIjSOvsd8Rlrn
/sDHTZM1ESVUMZCV4JyhcCGHokGbFCKFzZUJqhKBxgp7kUILFu/6H3/7iWQhdBTPf29KBrCne4+/
C33KajrlJG15ITxKldGvCHAqQc/DPhhGioGsXs8IJoZbJ0DI8mNaVd1Lj32pfHZDprHSKOw7M+wV
a/Flgct4M1N66bEsK8FOC4scOPhO7GVb3COL0nOpZYaeXxrij11NSVKbvQskMTLJ/5TG9uXbnySF
m9nPDlbsem8vRtZjWLpkX1bPFs3efBl6vb4CfKok+5brqXX8rlhcvUpJ5aEyjjhhS75LB+xWF+Mi
38V7m79OBlU/UnimkWpVw4JSqLjwWMKn6uKEfc3kLkvbLFVpeZ5yAiTm2K/QWYFD8QVdgdNQ3iuk
ppw5N8Aq4RPvTfjJ7oEerPeIEaY9nbLLPSdmmZqShiPxSi8UIOMIvaXX8A8OcDCv2q3Ui/0sumQo
EyWxKuWKZLo8o3SpxEymTmhmev4YaGkGhPwYFU9ctZD7I/sw/wK3tC6nVZAMZvtF+91lgXboFc5i
qQVryfzBxz+U5Wy11tEtU0+f0hgJn1jn0VgAcMPguXMg7Gx4MYwqN21XQ08zsKeKctGAwq57BxlD
mSPuPWpGehOi1Fn2lToGABa28LhY0xt1S5hn+oL2y60OffxBB0lv8uaXVwBHf8zn37PLDrwIfJNP
nTnOQf/RBiF1Of8tVBfZ53fl3/eVuGY5dd1Sz6iRIjnQd5fmJpRD2U3ykIo+Jr77QPfUn0wXQWOd
AEbqLiIusQ459q5qEwR6wJAiSk12+DWWU7SDPj9mZdewPIJkLCibu2lh3iYgEwW3MGctxrwtPa+6
F7pojnz1DNP2aG3BCLnMP6kPDw/hL38y24BAJlasvMukukgiL/7Fo7e6fXO3YlNwXBn/zBcxUCIH
UScOveIuhxESrvvftRI9YJas4D2VmzKEC03MLgKVg2myFdM76rWnVW4aYgbne2FVfPkmtedaFlIU
hGqj+ZW288l+sOftPU5ABgGyBN85lYcDAEyF9w7yMDr8waBY6g3ruyWMKAQjzhYM8j+MY7VjPIRq
2/ZJ1D7UR8uWHhQVUyHIxzL6xrDyOqR/8FFESN4DptMxDkMOqGSkABTKzqQS2gV8K6laRxegNJCM
2I7mETnMMKqbEmVkMUSycUHXzdpngu0rb/CuayRcE/as2EjzQFVdSARILXA/0bjOuGREVRGiie42
WEgKv8q3en6jkPpu9T31dSzQlTS65mCDvGdB0fbbfJWDvo9TOrsGzCScwdxFdiHm93ZKcZbiSnWx
kWyJ2+19B6Bd31xwIBbUeMnL5uMdmFpqbQEw0YZ1yTd9quJk2XBWhgfcwbjCBZJkHbFReu2tmU8u
ohW6tL29L79YvUYud75RgvEy4E/0fFSfiGUmwSPGzjYYWkbtxcLHQne6XagCp+Sh5vX4JPB/DAES
8lqw3OOMo6ans8NuAlG2jvBdJyMbviPy58A8P1bBwLKE/OQqr/S8n1K++WcnEFASVuIEUGMCWSfN
F+AXyOuuZGk08Rv+KuY66nRQ1A4yAUIyHStwFGuMA5oTfVqkVW/XdbWgR3+hG32dbHILzCJ5ZWLu
w/PqGE2RkG22VVGYcnreOUe4DpYlXB3I1wrQKxjBa/BtK4MxnVLTb4UxBuRGMoDaZkNS00Ya39LT
NYv9dWtSAKEGFyIlwxe2hRguc+yUzN5lbmFEAvrLBXbHMNT/72Mdyu4PunL8PxaIv3rgH7tBZ524
4ik/8YtUhQHgQuMt59KHj/yffzM6Uoxg4Lda8Bz+OGYJqvi3/SWQephB8Cx0a9PCAx6mN3noccxQ
za4u6BO8hjL8+/elrfU5XNENwoqGUHFyK61I/qL6CNz966XwbCeGtRiX238kccIHpyt7A2iMc/Bg
L8X4tbnQBiTm00QnIwLYZ14a5gtvsKypaFIslk8um9LrrxmR+deFWNCuUdmV7s1FEvHNP1aVimXj
69lv9/iLi5ArqXiUCt33lCf0uXsSNkcq6cx8qujjGiFqL2EpCmInd3zucwaH0N3MaXYFE+hIt63k
StsmjFDqEqKEx5k0hArFzBTiE01tTbyr3PlhS3+PNnDlatgidIjMNKmpmOujzvj8GL+tEBHgTu62
fOKrCX6Vfi7Dg5GPaS0BKqsJcK2CSGkzrDWLIVAH7Ohd+bWxEztcLABE5p2/DmR1lpNc6sROm3mY
cJsTYFu2/V94hShgpXviNf2ouT0a5oNrCsHNAWypVPvStiPciHLZB+u6d1aIFQg+GepDYPxHx3kW
92w38adGni4Wqralavomrpi8c5oFpCyiwfijJkyHRkQ6u619y+d7RknEiAQ0Hl1i9XXLRriimuX9
JluLGlVCqVFb35zGTU0uDCXX6E68oiuK9GCFNUxzh1/7ITzLCfOVUKM9pmQmF7VaZRsPoT3MiC3V
koBbK/n0rbqWw9hsqaODedRyAImz9ebpKViQ4GwSoV9cXkAHLfhE3XXVEzHsUh3fM5DnFrDWcSDL
d4pxtND7/V0akjw3MESl4WOgoFGZUoM+WfkL3lbUJ3PcLnRD9BU0pUZDS5/VZUDQTFeNmTZt+Cdd
CD2BaWApNiK3wvEHCA2R5p6WMQmOeyYg1Ve7axQD+PinVMZGn6TBmNkk8cpvHmCrNmRfepCVmmTw
jorRwBANn6Qg2jDbp4Ib3nketyBCVZLyfw2XBWe0gqIaL9d9TvdvVnIjQRpI259B01C15i0vJfF2
rVEJC5E7lAOHNAxrslg7KV7bUyhmgrkvcqszdCZq1jGTqPcQ1hQKstinq9GfnoFRfD7uLAVMh1jK
tdHyyNCVoMG/Ga+pDPWkCgq+8bkjN1weo1XmdXrVEcArYaJlqYlhLWsotqjLNsaGTM5AWTMhdDFB
qfggVdf1FerP1cQTBrpDJRU4RiLyB/wl8YSe55wZjCYx+IzXnBnoJPcIoUxKGePQrzmL97+gpxFW
R+qrUGdqdJWJE/oK99nZu+e+ka9mHYdTf/NaYpthVGeVk5jRw+7sMd1/Bk/9iBeW383vjQgAUCq8
ZqFfqqeeqq/E7D7Y7pb3iEQz0aKAfRN+R3pFtcAZv2Y30osxFJIHH+8N0NrIyHlcZOR7GXMztffB
wAj5JyesAPj4qclP/MEdApSIaMElA/UzG9JDbueKnQ12cRWs4u50xPp5r6pmflGEm9vhp8+2hRxa
7DUTinYppDxWFUe3+LkSwWrqm9l6b8WJY8WOjy8PiAOwkal5oQzjbOfkLYLhfWCvx2a/VFV8+ycp
/14jXi+X0kg99uW56epS3o0nHw+aRkTw3aYLZFu/PKDPnb262mnRTBVOqFp1XOTPJprzf8cQdXQP
sOeP1/mwnuaCf0f6szHxD7sDDbJ8J1pjnSy4A9hyZKnB8V5T/0Qq81AF3EwmbkP1aRf5jJJYKZUu
+ZzlKwyxOJ32V+j0QOl8WhdthNH7RSpDGtapRRf8hx6C6hv1GO6ENHpyeMx5L1rsrZvXjm3n6v1A
zcZNL82ZvICt2AWgw63gCyNi1+/J2zqjxpR6jFnbjFD5CtPumqtuvwcjbX/5acqe32Xnq2fkga0J
SaoYR2ZiGI4xYnak9fAVEUGN1akaDdAZoYhogpLfJYn09Xj8Fgq7O7In0IWDExrjoQYqSg8aEmjP
BTzQHl/+hdAnzlK2fUYaGhSpJy70k8AKpuu3bEjkKDuwHrZu4qQWbMwFa25rI5q683EwdBMAF8fP
owIShTXLzDb1UOfaYqUY2ZZSCxvcECRyvfbKicE5LLIeLQbhXfPanuJ8o9lITK3XE5hGAJxk4rw/
k4xWaupDfa0FdqPnvm5kL8NYgxZ0iQtVY6ii74vYmIFZQ6Z3GFS/Wvw8KMfxsW2Baceb9zyLxm6i
qbCwDTCHmu0MkLD775VKpZ2j40kJBRVgpXNT+0/mQO9OR3hIl9UjJyC4PQR4JlRttr/Tdy4cVT5z
fR1hQ2PsMSA/XteUqMJcjHLTmejMLC932BIhc+OYKqJtcGkT3pq7dDPIrosyVw1Sm2RvPCCJVVBx
OmJeCymOugfqAafYRHZIgAVqMNZs7xsj6D9zMLjFCEh5rWTqCkd+vqpLTTmkilBY+5cW7B42ehrC
eI+lOXyL6DybesoP1xuIkSSkLdDpy4Tj+x+zfbKtVyeO6Xq5WT9OEHaPfVZqGjLOlbw53RjacC9F
734rTUJg1yJrLpyBKGpC5lywpUWN6XwLx8G4izU2JmRBFuQ7b/JpkoFvlZuhPxDZ/j79jdN/YZFl
4Zr+/13aHtJASU/kxqF3rAmK/yb4Kc3GebVagGmsb+uohJMRVf06M1mOz33B24nLIFq2jLm0Ep0/
TOeOAK4ss3DI8L6bPdamZMjaoBOu6vj9qrHd5rtU5vVUnIfm1Yeed4ZpM16YD8DKGX/tKjhHxudi
5JPvXfuaSMbwOZXk76r/8bPv4X9KbEywRDBlbdVVihlCJrOHWfaYQqD/JOv1Q7ZZaNN6CHiyPYWK
6IhhbJeQGuRTE7WLmQCp3fccPdaFO2A+ozR+FcowiT9U2nstBrZY/ReBhOfUKehk/rGHQWlWxma8
EY9HN94d//7I6AE311apinY54RfirManGu6loAK2II8IKQ5Nw7l/bLsl6KQgZPq3vL4NSFOfte9S
1RLRWklHT4qRB++rN2U4gaNf+hr14qKnGEwbmZQp+0IdlqO7mpTQj9votfdw8ai6KALFLezxr8ku
I9DRmpS7hnm/zFI2zJxlll1vB0TSby/uZ2c7IEpmr422X8zQuJMkwEah8HOPkD44yUdqfpT1MXGa
YWWf3jO2/BzCwxXuMeVXoulQdhp171fHllf9PRXh7SJQ/ZXn7pHc2FjnOqwFUsjkyIOsVs37DHYn
B4fdvsUlqpq3xdM8CLpxeTAqcEcZRQCjyMLW6H5iBO/6EXL7yp0IDxAt6bDKymzNLhotT/RMieho
GJ2HkwDJUzZfljm2OYgtQrbqzlBV7xNLuBhuqmiMoV5uzp5Cp5rg5fOvWISX320ZAHwM2Ev2oNmL
w0f1qysBQAXsa8eZpZOBENde+mcC8q/qoHlVI+vxUTb3VUypOOQwGj1RuI8mONv+7St26MgQKeIX
HpZEA1zAaAAdigrw5LgLltDDAtOtjYmryG3iTMXAUuw85rrESumH18NJ79NW3MxRr7F7NGFhC5hh
sPb3/cY02pY+9xH37O6Dcm+3uNgnsegQKiHlh9TghehmL13yNSNHJRd0jSb3dcJ9/dHAOkcV+efT
USMQgZSRhZtQ6HSklGHd+EjCLYVPCTRj2AvpTsjFHwmKIeFchQFQYa3baYFcLob6ZKccQRIlk1IS
5UK7GY+l3jRNZ2fbvCyfbDoP1WRc5wAvW8/xz5vKX5keHE6DAyGTQ8qQLhVKM77Fy/twcdKTX79+
VjUe70HEyhrg6e3HTveuR38NbcIjT816NB8iZkTklQYulbqVmpYxjV1Slbb4y0Iy7Ztd4NPH2DE+
2DI2cDAE50R/6ichFfAayleiDneVCoREhYR/YGUCVvp2LL4ooEl+3WS/xWQcKz0KdoOk7jwfGDiJ
3S6gMZ9D3L0sva4mffh8v49ceCQ9sZoGKbt7IFZmI/AaBfmg/M+PfJHto21uKE/gvq8XQmdw8dYx
z0ccIYwxrNepq5qWM5o1A4Kp/7paOtXQYhzKF/wzeK8miBF+p7Lz+ssRMtBfWWzgw2D9qp1r6oN7
En+vLY4L/cP/NIsvX6137PM2DKzOMlYsBZGArD5WnOQPEAWBiolIxq5J99JVFnXAkLtnDldouNrL
gheP6fA3ucqGbcJKyPQX1NzY89RxbriXzOedy6KQask2HEdh9/qciDALtwYtPFFuZEco17dRWuTd
usdwbJ2WeFAsGLXWzF7N5s8KqRX7w9rqIiQ1dt9mEL3ePBMZeVBtRX2gZA/5LoY6e5lEsFlmTE90
KOEIdm1W/L6JQRyjLZAR+/a+ANeFBZHDcYeB0LPbNLfTZZ400Jk1U4S54p4luIJuSl0fvuneRMjd
YLCl5s7kckTpWkBnXgl9ZgPf/lX6Ne4BgjPjYV2Brjk+g8Pa1oFJlblyEQxz+e1rCJnr7KSJF8c+
fYso7XVkylzyToCgNnrzjLAoH2KOum0z3S1D0QO93EtllBDVcI9BnbSVLg4XJk51+oB8u6NNWIG4
uEMpmfoLH1pObEqDVBj+7QUHD9FmKbgr/z9zLwOf3L+B4VWs8uVLKv+SgmSji4XZEg1KmOk5kZjL
bSlLhDW4dntk1VM26CZYOASbLwT7VjFVrCvyxrIbWJgxqn70E4I0ajQEEYLw5YlHTeHlmhTfG/p9
QgQZM2Zsyzzi1y7h3NJhLB9JnW15HulV1b9rTrDIaIZK2PotZOzcubNTEmrZGhmR9UqfWoSkN+qg
ESddVKYdUyJzh5XrH9T1YIFkgmnd4moc2Bl9/2BCDQhB6JS5pQjVbYa7ra7h6wsImFYAxWZgpNKF
w1pfeFSTVZ1jetQ3+S82pSv3gz26LR0p0hgo4xm45gbUzHDUBUtRePMU4IsMVeIl+J4mJpvYY+F0
tP/U2Gcvg/DppPmOxamCocK8//FicNuHXcmIWRv+5NP+VlOH5K/aeo6bip88Di/zeddjntVo6jK9
KZSWZB2a16mYBeVE+7S4KiS2deNDRmuPX1Uf5cn2DqCMKSkAvVzy34+bnmVW29s5d7ZCfSPWb7SW
AgKl+nQ3FNdaCHtYDjCDXKiPR00aYI1XP+BYlbs8yO0Ocswc5bEDFeQd0Ji7L3wHM5QyUJiBjCQb
rdH9uh0kq10Qdu4CF8wCSlVW2vHDscw/JqgYIAhb4FtYO/rM3d+RIArHF4S5Adxp6Jbf2gGgRpIg
bsVCmeZUeitwza/i5EVyEfmTCrDotwtVKWpN4pLAikhEGNGN7QKhbSxJnYS3JMzg9s7TdS/+X1Rd
r1Rjz64BAb9wmFnNt8Ib7ywkXNx4zo1Vu7+wC55XcPEiAFceT1IZth6beK9/1oq7e9Z/2HAbdQwn
kXr4AT+MDxDl/grM++hCq/XqP5Q/D0qc5R7ubLC/UmC5YOBUoulOWa5Oa6jq19GM3D6Xlf3YHPj4
5HObpevnIAzGeV4Miqi4GLHYrNO578bzNdNqAar7kyf13QpvxEjKX3Ua3KFhizYy6aFSZa57kTSo
sF+slJGJxqitRjLb6I9lKlvlC3ELDanYAjVyTgVzEtyPX0huxukGOh2pQif29YbwWj6JlE2x7yry
K2kOTuyjYaVVpNmw7z4MFJOhs8Jlkad+ngXGuyeg3R8JN2L+AjOrbdEPH3nwDmSfdAmuTellgk4m
Oq+IpaNHo6YBXwhJZ3coNMBKvrR96uCscjVLLtXNa3I3jBZRw5MB/y2HDDmO+oIsmJIqO2ht8Qk7
qgnAPWpEQZ5OyoOH4IhWqCMWuRGTJghoTWcsPa5jeUTXkhuxhnuWdiShZDi3sin7cIxLyuI7oIH/
RC9i55RcSWu4rNcv8GEiJt6KqInLb2Ww9lSoc6rA00nOmDESLhleSuU9YiFA+NMgAn6wXy07BILf
s9/Dmy59zM6Be3vwmlsVgw/Ma7k9Q1NspjWoKeQgu+ZjKXIvFrVJPpkkD6YUmpGkq/f9scb7mpDf
y0YqVZW35TcWaH856IUmDgj6WLEG/WIeZJsiMhvRxDtdhHAoLjU7ilBOGTUaMLeI28GTPC18g8B1
wd4RjCULwPKaSG8rRJzhQZFgplvcuHk87Fr2BbPfMy0s4C/LcVj9XlRlPjLSfwlbHguPm1RX2MvP
52gaEMz75rGR5fducjCL4Pz4+3nX31B7F9y+8WmJt+MsBXvUyrAelhWENFOrtFX9TyB1V+cZpthb
h6vyT26Xqb5yItMa1hAVGIWp+SjpaViDjZfbaNs2VruoovqUqzifzXkTRJcHsQc0y8LgK6WfiBCZ
ZkhpRlO43LCCSe6n76b2AaRUWePnk5YKkAnW/OymFs9L5wYVFYjNVLKF1VF7Ud26e17EldyhBXAh
Sj8vQSJkwFKQmFJVw5KWFYrTsQ8fMiEPVFrbQgc55SV7ziHcNAQ2waNXeG8aDHOh01ZFFF7gGj15
hxB+I6ZXq2NhDNAu9VQ2YSk6FW9zLW5GLk0f+GZyC3wUHiy9xDROxhtY52rpJYdGIzMSeiqC8EAE
geGEdV4XOcu1AC6UpbRHEUg2N4v98naK9uYocEZbaXktIesxhc0z+vdmVHOXC+B0ItUeY7PAa5AV
mdkq2MXGhKDlhZd0AOc6OGwutPL6b+/TwgX31T/8Q2G+devU2CHuPZ5TgpuaQFnX7LIxbw7k1KEj
7Xnxg6/PEGx9Ht6mP81tHaE66pc5FYMuMPwaJCyQicpUgzQGUZXIIeda8JFp5ZUa5TfBNHftajWH
k7c4WIa25yXYmwXR6qGsdcg6p7UEk/lZkcuyf9R0gAm0ebk6HkU8uVX7OxZfrk24QTA9FUyZm/Fg
B3AK+ea7OrSZaRv6hRBr2WpNSJ+uCjKP4qUKZ1w8BK1LA7CWQG5WdwhsEUUy0cUrxBejHnOpzGqD
wUOcx4O9DkkpYZP6oPEke/3MhBWcvCtcG1ET4oO0S12yc+shCxjqfC37a0J44oCngZKIav3rEKc2
baHWAb2Fe8n8reNN8aCg3RLLOqIAKgzR5bPIFGTbwrw/T8fBlAjuoidDwx9kimm7hZaV/JVUzogt
DymJ2OyYFEWRV4kvOVrQrAsQdGMQ6GiN1JsDyEasCykvFPq7m1ochQT5cT+tNmkSVtchOYHa8iR2
N7Sjoxkyk2+rwDdemh2HHO87G+KJWt17S2frxFKf6Z43XpBL4AzfIXEXtsF/s3OsZyiDIMhNfJz3
iBlxZsi4sq19tgtescKVavKqcx+xA/u735IBTldTFW25ZWyd+ljGOYHOh3YwScMPTXF68s/a3yZ7
eae/ACt9bm1ISBJUewtj68Z6ZKZcvM56Eyz9Bo6Vwk60geqAFLv7M1ymJ6F0Bj5naeG9TjJgdV7I
ut1PFTTzuqAgsm5+C6XvkUgvp7ptE1QfdLBV5vdWWFwZO7Niv0akAzXzUZTW/5SPcSRCMMwhj1rs
IXRc3va0BwqoA/boENN9pr30YoMhYpM6/uCot0FB1U/OyKk/eMqGecnFothrqUKbQkSeLNu8xw1V
WazHADzwZMN061KFVH/Jr976IT5AT1WhXiUtfab+tlq09gzrwReqxG9XjuEMV0/mvHf7aa2E8g5+
ViesQmyDba1FvXc5AQG17xPq0rmSVVAuUglH3wSwlxMhCEw7g3kNdnngrOqgbbvpxN29jsXGVIU4
MQBH/t9mOvmV5BqmMa3mlgJQ8gtXf443e2rWKSeqmGpsfrIRF3CZ70dY5kojnvQJgkIc5P/aDhsD
tOgpZizPkYd10CfbBuqWdCGcwHiew4+3y6iUjEELoKQN09MZjC1d8TTlxjdWl3JW5yjJbRyF9+eR
+kWCgUbktl0yekDWWvcm0MtxLLrG6ElktUgSit5LLeIQ3YwVuYgVg8bFz9FY7rdKHolQ710ckni4
EITxibCaxDKsSAQs5ecIu3r9GWhC83rs0IazPFmP8XeCkCF/8JUlT+ROokWByc1wlgOzWIQiUHtr
3WZgtmp+LKqJrVORxb+YqLoSwnL+JutqHEPE8Ip2jdqu2PCJg8QjgZcZQECyC9IW5XwPP9oHNPb2
vSHVKXH/h5m89lxMyDecXp2Yz4F0eomKE7uEXEjeFYo4++p7lOV3BrwaROQCSt8DlHs5jJsk5aJv
EWbeSm9uGPugnMTouncfkvWbEEMh3eKUT83jrCpHn1vHdjZQCIc04/r99prbXPJiquWnD1hrAjDJ
w67PCqSkjC9Oo2t6EEBxoppdpsAxaTYRQFeWpKnFZkxmsAva7Wa28v25bzLKdC84WrnMSziRjcxS
PNAO2cvOgAbyAogRUt5+LKgusvhQw/JJigG5Vk+2Wi6TQn3VzCOI3xruPRtLBV2F061r89BMTPBb
kRwOMhirMK841hmGxMIykb31So68tqNP1Cvktwu0QF1ly7BITpUJk3tLzaTA0j+ukR6SQiwhEor7
TLHvCuKgCndGdYT+bt8wznxJ3TcPgEJiepwwaJyYJYnGg3ZUB09vM26oL0oY5QZu++fYpQmtWSVW
T/0Um3egBkwhWK8ZGsznOBMpN2qqadwHv7lMXZM6IB6Y7ydkM5KGCZZtWnmjTxBS+LNabx1GSN7A
s5fcM5Enq5PErCTCdr817PcHjLR/Bo8/8rTuORovtQarE8y0GvsIdTHoJi3D7BHJWq5RCNcxbHBW
cCHgntz6ngkUcv3LPK54pe+IrSXltTLR+AdtIdinV9EeD3rXG4wW7TaeCrbCcEtPptwIL2ivDqdA
DZd0IcjZClJlWCvQXs1f7tYvMeIn7kWPOKJTQg5oOwtJ+Me2vwz5wHCTXO/Pw+Mb1yuVVfdMPb4S
44/7eC+VgzpsOr9ZXUYXoI20LYIbz73/2q0Puvh2BMDzRfnwU3ruAF2v+iykkqHBlazd1SmKTUhW
qr98kAccZVfAw4oT8bw7ol7+yeNzsy5Bu/vT25zPipGub0DvNN+AoBtnN2j+1eVySmiCsx+oaVT2
4vsLCIHYrm4oW5VpTdR1wT9Gghv6yOp6swZ2Pf5/hZU2XQibw17oHYZH3XdI0lDPBBUpWRKUhsQG
c8Tgn4x2zmcrHXiX3U5iFit71bFX6GkESCQCaYOzr1aMCEigUby4ntSK+vQTqAuLy7vus72q08qW
qzKsH5Q9F3/w8DZpo0jND1vmbaTTItMtHlJvqe4Zv+0+QHX9YnviMer2mJB2GO34yj/MtzjeLiii
EIdVVURI29lsvHgYFih1VrjY96CnOBeHaxPdTeuL4jNB8WDXyoohT0i3wzlxeduKzcHRqpNjplQR
QJqrzjDP8+7GLM9PMJmuMtgCF5y6aukf9MCj6j0yQtEHwc3Cg1JoJg8D9SefmdElNDWl9sa8F7oj
uJG9zDsOXIgEVqcfH6JnSQZxi0IjnlTa8+SbvdoEnOyANld8QVvqIYn7c32pMAk9+LAx3JEFHpTP
8aFo9T8lBmiNckzWVimFD6Y7FS8SIRIZx33C4Za97ooWNk8EQdkf8KoPFtBr0MJHj/zHZHZ+4ANj
thy9XDPCetLiUpssn3Qg5XJcg8yGJBytBWR2xQ/yHWZKpd+ObRWET2o7wJznV0dtW8zRPP4KMGMl
RCrlAOXHBTNL2ZnyHDu6SEXB58/kdSYyDqpzuqICdfMRfRmFbt1PjVdgqBhsxolAF4GCS1SVx349
L2Lgr3nWoWTKDgLHJPx/UkYAlHQqAm/OoJk9YcFKWtVHVYXxQ7T9VWb6jNiGqZa8jSq5ZVNybJBH
a5limSYfNLZNYZLRIjtB9f2MB20tOgi1KYmhJ9cIsSFVYaTdReOi3vkclBElgpr/sSI9GyOy7UHz
hrM5yBqv2+JxOUb53wRsh/F422l8b4O6e/aO9wkKXgKxNZXuRZIUN7Ekxd6NTs9hSjhf2447QpJ6
NelxWu+9ApnCiO2YDv36Cn9t5BHYVTJCIimQW1ki3F2KFpwuWj97M29st7x9XwxlvoHdo2nISP8F
0O+RCt9h2p9u+LatQKGKHKaxircypdtPrTp9l7eH6xzHwWIXdyXHzEMijia/goqA3lBJVVO/oTB+
XVlCl2F76IR9CPZL6THzPsnsC1dM9Uv76VrJ5kZc1vhneULPqr6eexnFpoXkdTA+gW2678ihkWH/
uIbg9KFbcDqsrqDDXtKuEb776kMVx5XCax5an7aEijrwU69e2cKksHT+f/MdK1Ej+eULvOGQHKyx
pyyCVY42ZskfNz6nt7qsmhDG1XISlqpCeyBvGsBx9q37NuOmEEkbqOxZy1rf8EFfDeUWGsOBrVjZ
W+c54whEdJyTdUPRULg89HIv0LYalpzdbCkKNZHJyaj3gLj6PkdP4T2n/u/yY2R7TIpkNX32UvJZ
JEb3mKVlR8199yPXHTvIBRClUsr3ju0ZTFeZgFfaUDjZ4yN30+wh4dR7zXJPN/priMEbVqajE1C7
PzOStdf64aNiEcALwGhUH9e9anJAlR+mVODGN0/gfY74WWsuWqvsInVCtUjzT5NeY9Uq4VvsHPJ8
KMlFUwa3V3XMK7s8cRvvymjZzCIXonSPT688Fjgbr78eRm6+6zdpoUrLQDGE/BK4mE1yXoHmuIM8
y/solWGoTFCsWvEhyAq5AGq9AOUkjHgMyDTZ9UJTJ1mzntXXAULXgoRWeSNzoLLD1F9cte15Tk27
4qRPChwAqc0UArh7QaGfXTjcXax9DsRT81flCdd6Temj6ZbXalFDy0esrghZqpA6cC5YHfjToFXH
KPqZkUokH2lT82/0RnAsnRYEOi7BBGZynzwkz8Hv2UyOj5p14PvMH75K8+dCJOQBPnLeG2Gf0UV3
LjyFlqwmjYpETiBFWl0+ZE/CiovOSEwfx0tMfTsAY7WqCx/YZOS6M7YrEsmqGETAxYPaJItf+M1P
R8TokDEerGzpT+MX88YCVXHWl6+ynEpuOY5ox+IDNUbn8YyhZx2ZOpM2gPmb0iSdsYSsC5URuqox
Qy0KkxdjmggFXm6RlMTL6SEM7T09ecik+1caRy91IM16sL6auzi9e6gnZE2AvN8wmQK2ETpxTFHS
l99hgz1YY9o2J8TMiX3s4sSAaEiHfMbrWaKZ65IRq2NOqJwVyms3R8ajxfdvqz4RByX380bzCI6w
/0dP6XF2KNPKX3gc91QyY3uJ4pOlPhIrH7M/OIROQ2/ZWRbyeBOUt76jXmuQn7UGL6FDNBeCC5hd
0Eqoo9FT2J4Hkba4YqqQDeBqniYbfyoQNQuFNjRzI5/SxuanR8s7f7A70Vw534+HPyfIMWsFphji
/52+glhJjzoyQQeGMVjPgnhSwe1TsQqixEcoDr4rH17k/NGm1URZg+/qmAojAUgBdkWAEDzYMO4R
7JjOVGaq6BfQAHyoSFQ67oxgjEc6rinId/rAY4aoCMEdlFz3beVD2sFlA/bEnFd+OHkX0N9W+t1N
a+BlQ5OxxDmNg/ThT0tZBvJZw2pBVuIv7cAg8gcs3uWgoMW5Eyzx8+urROIP9yhR9sTfkOk+Miv6
T+CI85mRm+ofTRo2BkhG8q+4qEpc7kj+FJtFKzRqTB926U3oTftEA7jjobzNcs0jnJZciT+hJFwS
Y9E8+iVo9LnBPsMe2oaeuIigCvvZ9a5+tMumTfcsyqDlrFdXpYah0p7+ib1ZiFyzHBSnCoBulI13
AmV/VlZduEgGBR3A2ZCvvr0P1eflZboux0/TD5R63GNzqIpxO97pbY5Df0pgQtlkLZTrKQhe9x/z
3EwIYf/IW7dfPBecNTsO2/PBYxq19OM3rGleYGvLRNwWLNe84+F/fsnZBYwqGZG8B46zv4qydxaV
YC/7VEzpPU+I5HKgb85sRyqBRuWOXgwEPM47gk0IfHEVxieE64p7Q9n5lmYuGAhheB/mRo7FYQBW
iXTGUEAB60FND1FxngGXoDI5wAQIUuQz5/lnzc0bhOGwThI88UOU9FjW+dHENuD+12bvnIRAF7GO
CMicw/pD4yI78b6QMlWiz/N6f6wraK3+xaOClhOE+zV84ZBEHYr447KR3ExO/NiEaecfviJ7B4wU
7yzCUpmzN8e41bB4gwypCy3xHrikP2LkB1sdHIhVZ77ghZ3M0BN1QYTG3YqblUEsnmZbJNxqUVJA
s4SfFqw1UeF+C0HjWu2m8LZMoaZy3VWaA1n1OyGTMuTZXoL8Xzp5N17HgaqlATpupM8MT+zt3f5T
/4+RYP6JQ6IpzrvUpeUNRVWlXOiMwbGRDObzamOKoDcAyOlROIrlxFFx03vaBFSasUrL/A2gZweY
gB+xprQ75saFsUn3zUYoBuMVvR9hCO3BSPeBcNKXWL9SYtG+dMqTGQt6lnd/O2Vd47xnLNUO/IGw
MMqsSzodRO8m0udMidJXxwVdvlVdlh5rS+24twORiuo44RT8A1JvjxVp2OUcjLmFhgpOzBob7iWH
Yz5SYOpq/cN8nWl0YgTd6YiLuLIHZmHCFVCRszknIWgwDRaOijP8kDXS0XMnJqppU3P88tnMRgNS
7i01hRVLBdUSPAu1pm56nD77qHVhoJgfay/rZz7+HbzMbiy+EOflTPU6nawvyW7mhsIR020jKqZM
/5oIz298R3c3YU07XwGWxQcHtAGl5HQv5kpsxq7Z7+vWKSFhbznsK8fATVCtQDeXaMTYNfYIhXZv
Sl/btn1c/c4HLExU98M4CfLnw197o95dbaqj2zRimpd9ObYFcteEGhPJgVjr/Zk/BQcIHgIPr82U
sKnr16oyjHRqrGbZKBa6GKAqZq1WJGl+oIaBl2ZgTs67oowbh0qSO3uPuXSgjkwwLMNHVPYzgb0F
JDlz44W9dTPPibcQXLwkoJoTUkUEKvfC3cih0Xu+JGVhYGnVVxc50qV6P2u6+opbRQqsjFxWN+eP
XqLkwsRvVmtWgXdxtYFvNJzWTgRCSUJPEiTY5y7aY4WA9m4hmHmvztOtyi6khJCmTh8AuX6ihT5P
tECXEAYBK1ZvZJIllCUfcrRLE62luXBubrFGmXMcVDDqbedTk8OKExA/jdwIOMosIZC2SXv4Ld0F
r8waOK0kYqmVoQ/EbBOSYiNl+Fg8PqtHYyK7qRXiucI22/atlaFOqRF5Cka01M1XhQxvJ2cEOpIj
nAl6n9sySBtgpOAS/u+q/Qmesgc2h8TK10Vuz9PEwD4RDpjatJQAz03t3XJGVkJbUd5V61vFrKI4
dhLy06YdxWXMCZ3/0LSf/gKqBH2488G/DTFpb6+Fj7zcvheg/cSSMywypKozqajpgZnNIWLSiKjZ
fpcHLn1q2tSagjzLx6MCwn2bSeoE/sau9WGiibonggBAcS6QQpqz1dMdEjmVW5/OpT9k8NAPUlM7
jBuZoMIGCR7U+ZX1t5gCsW4ByI8OdwMIqXmKt5X5XkRK6a4QiH+6cCqYAJI4gQe2lZrDm9Dmsk3n
mbNopYPsoDXI5t0bwRrS/1k+G27WMtanl7YXJgIkoa6rbkIgf5dpH3W0FuP5bpssooAXgYJyMBcH
rYSM1HQdDDMvCuDNRCicEgcZQ56BHeQC/MbaMJrNYfnXWDz4E+ofl24GB3IgA328c7iMcAdIXCih
PBIXu6rDr5fplnd2FcGTEvUNjLHBzC2LooFDv745ArlzlxKn5F+o8Q05uY+qbuYV2yp39rr8LQV3
SmPLduo6y6O02rohvq72AKjGo9VfTURWOUstVwN/fSNPsCH5gWPkTwgfCCLoxu0qD50CQvJMwaoU
6ema3+ZzLb0NnuAF+vz6qu+Xp6k/Snx2zAjjTSX3VdCVTv/ypep5wrhtzlHE+J3NmX/xOnapGyLu
06aXMfWuaxmUDnVO84XpJOBFJVAfQyzuLcgoSETJAn10inJ4CdtCHky/3Kk1/coFOvmFcLG04H8B
vwFHQqHeF5y7+h9YGCEryIjlDGLzt2Uz4u6yL8UDUQTgZUrJzmZUOM1X9/WF+st2FtJ4FPGOZtU2
1iBDZ/ABm79nw8TXD/Od8jRIWXDdE/SialJPvbaRWyM77kLtlBSc+NXJqULOHazKDgQvRfLhnq+H
LBGbGzT6q9f2Y/AIcKXpRigzJpm4TZ4wcZeMpnWscbwf7lpATJleWkCRk/bjx4OyRshUwGeybvFe
A/sHpekVJPeskrjSbkUz+wbpAxV3/6po9hKrTMixPdir7RgEePV9Wxb/DrRlRt5+MtXFY90mRn7W
5RIEihnsrEn0V50IDkVOdSOXA69jS+E5VacfK0jUHXn0vcPyNDFY555DroMypb1OJVygFhIxeAz8
q8mooCe8Tv4wOwztAxsfy/oRkhEgpNxFf2ZYNOtahmxVNi7Mb1dfI/fw20KZesiOC33adnEtSjCJ
yHfi5k0pI5Z0QUe94t6ZjMpwfT5v8Y0MYg/KFwgZ3kQJPgdMF7nJynPTmQk7qAAJRrw54q/hefjM
XccPeB23EBt4togVqdFZw+W6wgx4syovZuKOdiXMp2iUJOUrJlfDFc1Ez8he1nOtBqX0T+bVq3+1
6/DSE0vHkkqCy78gOXer/J9CrT6mM9AN2ZwfmrBDrSMzFoySWzwirgYTw49CvBNIRvKfnaIl2OPD
hesaWk5Ag8gjotYf3J8a+sVKeFsQ/MBTy+c1oSYN4GuLSmIRB6tDnFf3/pmYzWX+x0sjowQhOi8+
8UTTwLJspMOqHIBoioeZXJVmbVgKgptHb1Diuy5f7Ef+pj8MmwirD1xfRrNibJzpAZpaEqVqIrlo
KasYE/XiQeLCMKrLi8QJqF22rjXnyG3kqjOudM8+PBj+aetUzLOpH8+6kf4DtiFl+027JbIy5hXY
/piE8Bwab4puRo9UtkO+xoiMB9j/cJv+cyj1VHNzBC3+4HOTvOqacxqe5Y9dbbtuFiGy/tByDxiB
Y+7GuYQ8/LYmm8ET+g6uUWN7LcWXhh/+b2/Y6BOKMDV0e6ploeYh3louqEK1aPtp7fMo+OHPiHPA
0ehyY87jz48ge4QMwgjl4rXHyE4q54UupTW/bOY05bK/HQW66CCu4N+yHGiaVSAs+ZX6Fpa6V6EO
fA7weoDjXlV3WU74XCSWVKukpbqHFFl79YzmiZm842IQoX2giWfrOiFKwNLjyb8K4jAI285WLMMu
nJpRfB5PniY4rKNVqiW0MT66RFWpaom44qmSQj106i2MfiUPEekw60VUAXrVHVkqsu6ckowGP1BE
C/cs/iNc1K6S5h6TQNAMSSBtqon9VEG/YdxJrfEYUMhl9UhUwelGrmFwfcr/OmeCWkLj0oXk6ogp
WAyv+YT26BG6ZAOXC2gz+gCxk6OgMYI8BjeYvBsLtc+CF7fs7Z5Q/VUgHEJ1IIqoeqS91ZPV+FY3
I+OlexYiKPIAFCBaLlf3T8If7Sr7b7aiq4A4Hl0Ck+p3cS3dDl7iYjiWwpdKrHylKYAUHQXJ7Ork
f22jH937HSYN9dQt3x2W4ZVAoN1qUcbZkfXGFWy47j3rVHWcQN4/zNSgh0ow48jK1AyEffOMB1Ek
RqjL75+KXsgzzVouV6Mu2P5xAgofgPeyH+621Koyn/9wwjBY449VKsBWAFptGSNcx2PCO0QEqDkN
I+bAtSjDaHs4Bb9k+f5R3ILXv8ZfiCatLqT8CQTmcU8u/Zi9f2aHDrVnnxvtG3D2mWYkTY0jfSgH
hCutYcEC6a6sLIbFg+0fySmwxCeEPzWDWPhTYn2s1QO1xaVdeeTYCNefb71WvutUFvSkwav1WtrJ
ty16qRirLUq094tns+P3wXFxG3BR+TdoSMqMEJ53Zc8n4Z8x7ObMcCdD+EgErs521rsvl475x2kO
t7bOI7v3+V4hc3K17WmQso2D8V9S2KpTuX8SJmWeMK+OtDBXvbDRpGgHt5UD7M162uTV7OUTYgWU
pi6MTI74rjLkC2z6f68fT0fSJSel+q27x1vw++XtGXx34uVz+qnjwm+tk2jrNc5K/ur7UOfsMAbK
N8ua47lD7ix/6xD6LIxsWcSCaBK04Q8QZEsQjXVh7dzD/QVVgY5OazclDGPV0NCsrO7pyOABUFJ+
EdYiAVzwxy21r5VYyR/1m2f6e7KDYkGKV6BK82KQDGoOiQ//fZ6SOsacznFywqTJx8IvgAIbl4/w
8SXNfzmKWPMyNuvIEKh31rfMQRgELFTzDuafHvGrD3jnT/rjUyXzE/oT11M56LP32ZGwl22/6pwj
2/TEdupuZ/WefW6RX3vvgZ1Ah22W6ex8vIJIs5yPc3JGxsrzC2EA6IVod2X9LFkNNvpPC2L8/jGf
YpwIZlGYo6fcyCY1r0uQL4Apo7vIMlQunrJiFDRSHyRX5S4v4TlD5WfPxtCJ3pmqfoezwox+xf5Q
OLrrV9a2uXvu5TqOUjqKj1wYReNnMw6qwk0unOpsv/ETqQMFQWhxPz8xa7CwiyfhbQK4xjcqrBz8
K3KegietuNmSiDTJkp1J4T6lU+BLl33a1g+t15R7FIfoti95Y15P6uPO/m66derrYv6dnsZJOM4Z
l2mM7+vwKszfL43huZ/ouogsveBM1UNj7/oAyr6u5YKZqYa14c0JRb5FzPudnQ1/OoL+t+IASGQb
rY4h5iuW+wa67R7FyyiAsON44nxnLQ+OTy1SXCkk8ZkcYF5UlRMcZYSjuBvpWaMPjxeMzylgY0/F
F1kKklf7w4VFmz/IhyT/q1q7L9PEdWt6pLqL/b3vNlQr9UXBy032PGShlWYE0or4qfyghKTrSLxl
HcMyavCN6K6P65IkEs9rmH3VF1geKA0Vku+jaBNGTygulD6vBYnC/rFO6NuJRAu1zdb+LSsHJTDb
AnjkF2SVVLPz1m4UOyTc3aVc0lhdY5uTgmKSBFSxws5pvD6BtUVqedqtKb9H5SYXDhngtgYVHed0
UibMNjfBfRhpB9l9agf10hSJz7Fa4vbZ19xeYCs3WsXiaNAw0Ng6OicLkLmAE0HNnWWXadQLAa9b
8fV/4AG2c+HOyZx8JLgjrlG11AU2p6E3EKl1s6aNQp1lE0x5btgQrySdLOmmHdwkiunusodgRl4j
W05gEhlEMKokhXSBu/08CiwuuR9pVyZY3zhUtTU24Pi80jL/28KYariLFQ7RYJLEmXOSDCrdBXoV
rJa+kT6lKbbk0XvxbjNfFaizg9lzRk3VxzOTL8j3yZNOfkNHCKfgKfiEv0u5W02pz7WJoDeU5MTi
F3XHxfVjEUKDHdcmJSu0kBGWySqUfjN+6OW46dYQ586FBE9ovDFLXOwxIhuoERiywzIypm5EKGdE
saJ1OZQhiuJInDxNZm7uKZumDWmumScjNjfzplcgjQ5Wgx255TYWPA1Qt5n8gf+LCESgpy4p050w
yhJY3+b6ieEDXGHlF+qJO2nWtq30HgrD7pUYbG8nvuEjQ47C1grK47whEekPyJ01bGnWUqThpSXg
y7HLHcGfc20dHubhDWFBg3sBe8toBKAZCgSkEzvv5T1Zmv8SysMnc8rBeFYlf55fvSc9RsqAi+wH
CuVdVMbV4drPYPTVkKLmpinTElX4qTgcsIA5nmapb5k+KyGuveSL0ma97XQzkKboUvMTL7FVnUp4
XfY+PKPN4Ug+iGQ0wB9AdYvBib4wVoO1JHN8zywQxcHQ7cfIFXvVIdCl9876Lvo4okTT+YnOkwL1
oyzhP7vx00Q9L+IokCxwcMvpxsCKU1k9yHev5nterB7iYWcS6zqXzKP67ePwZ/3EbD7EDUWOxNYp
u9vZkDQRA6lfHbUyECTNxN2RFRd2QUF4tLHz2pWjJeXdq16V6eusBiJCr048qz5q+uqyNtc8XnLY
SU3sE/mE4lBknCzjeksP2/3zPTlbYYNGv+P1cCJfEFFcGT085WRt8NpSuCsyBgbyZzyZG3tF4jQK
QkCknpDyDFuBCrI/dJJd3wz8w4y0ibe841MfPqn5sRxSRSAu/7FEhSLUdaLRHFBg0qTHkW+HQXvp
eS3hmg7wjvtXFURO2fZOPYb6yNOuv65rlFivrMUsl6B0m1jNoMKaczUaFbfPGqFbMMcP05CDN1df
aO2xZrsW0kXBPoJ0jxnP1HJA7fSwdI1QztBoPqmEqijpW+8Dwx1kar9s7lM/Gc3tJKWQ2EI2azHa
in9nInydWdz28BLW9kefFAbRDd8FAGqaauOC/EqqxwfJwqGs1WBeLsoLNmNKzg1S8JyxQkcw+GCY
znxu/ZZeuiBF/6xMHnxrV9VRbY0lf3dGC1fX6O/bNJ1Db8TWl/+naZYSXT6NV1JdF0qtkOs5k5m/
v0/hdT0hWgfrRcsdMmjIz9B15PXrPZHzfh5AZwG2DUqhXcbxfqMvQdTKodTiicwAx5AaKRl5Yo8E
vdnrqf1IHPiDljI8uUtwdjaiCRxelY3DXvULqssKRdJJHnxB8i31KbyQVaJ7/cgRatPe6ulCgr12
Ex64y2pl3stzYKReGPmjKfYjHrrX7FQyHHvIy8vX9m4jW73Z/kBzNPkVLNySSHoZe14dCo1pTjku
spy/x33gvIrHBWJgMFSFWaFG3S40++EFyA8kY6qVwf193nm6sjeGRL+NhX9s5a14crl9Nye91H8m
o1Y68pcaPo1wJPhHwEkLUWg+kksyBU+Kh4G5KHn4VDB8IKJdMz5RvRIW+1D1+yhTMbm7Jwi4HBmk
ITyfZUNafyvRmJRgZ2MDEMBNG6Pqyc/nJys+yLk7ZpkkS53mcVtATLJEw528xuV7MWjDBKbVOUAK
WJPt+ENmcS9m6bjWoazhifDPuX7y4Y4g1L7yy18N9lBW+TvYiXzqjRtHiybXp3BKfRrKjigC8uEH
TtLQ32wA5gWWwUrxpgMYnv5FOGubAmxNtUZM1/G+hxSvexIoCCiFUZdtY0WnIW4+sp8/tuTKyEWh
yBMbTzKWOCM2shXm562sGpN/ZeNvFG0+nUBvmN11ZsyZ0fES45vWm5F7zy50BYtrR9fsZhDwg+Vj
Pmp5h9waCnoRxzUDGtwbm5BkN82EO6XT3cufX3/16nNFBaqEr88kG2Bfh4oET8EaVqJa72UsQ90Q
ee77RMROpZb2X7ZjQmFWHUEfYTxaUxbzKG5EF5oLcASXbxxPbnAkVWT0xaQ+4laW9DApvSIOL3+I
c/n/ymQzH6WaUw34ge5rDeLA8+Vn7RAAQU88BFEy+3JVSo56uUEAl8Olom8mYKf/l46//NJmDMEz
i24d2JOocJBfoBoUs1164An3HLpLi1vydEhX9vWFa5EAoQUmVDRaFC+zUoFnB9oS6qf2wCr6pk7j
9suAxD3yhVAPfEz7BZ2DZpl9NdhUJt7AV3XgbhhWd8fOHU6sY518dhm2JGH9p57mZ3pfHgyehpyt
UZKbvx3b6Y/5glW9ARzfENd+tEI4qtvUQWrhTMqPypNCkNl9//ftYrH1U6f0LI+y2Axg2y+Zj78a
1t1XKudgybZkB93unDjfnp8bGW37eB8Mpe2PzcPTO4dqzAlsdVlgFm8qs3rYe54sNxSwB9vQSoeg
/Q1DsXM/drWbJJx4jMgN8mShtJaivHy4GRu32vN+wY54u397pvmJAobIBNgPcEB456lRq2yuoHrn
jAqBjm4IU2twZeXbA8mnhj1a1bZheI0BHEO2tb0VPb2kqQRxlItaIcEKPptfktpnoXfj/ZlRxh+8
72QdVClnI0DnS36Y28DsrBGN30jOMKnTUo5GPJfcIeKOwNRo4Jvkxqg69cc8HcLiF+/ZUaZrfgOG
DoVlKn7JWc3+cBjyMjRsvP2schX5j1enBBVEd9/rqZvg6ELbvZ2MGXtFuQyC7d5JNlqhpYAbjK8y
aMp/e3BmlnfRKwGsjENp51ZDVkzPgzItsg2syH7JpF5b8HYO1UYMvHwRWdyuUtE49N5Mjx5fTzw5
J1SiuiBvzufhA0uOVwyJIAgP71xiN7eZnFqC7+C1b5DkmY2KSsHiHC+ummgPw8DMNYYg8emwpz3T
CTQxrDNUgasO4xoHr0EpE2acQPtvWPmBrnOJ1fA1UmpWnFvQ6vYKgBYh4UVTyZUhjd6fcB9y6zcM
yZZ8WLk48ko0kJVFCVZShjFnBY8/2tRPr7e1N2eAzFv7ZCBPHZtympDKyMxO/RwRyw/+SVqBQrJl
A8Y3Xh/y6fP2tnqusvt+s/omAuV/odH/ueYjgHZknLRliAtC2aG3k/3USQjjSl+RdHMltndC/4Kx
oFCXXWfDF9Ycm8inwlMcSX5tKqw4GPnzltH+IkBKjk+GEzw/sVh1hzqEV9XS/IDiNM/iIzi6O6U6
MQWlogIpcUIJfux0VPHW3QlOxlW9VxEOtmhHSeeMdPPm/wzFNaHK/pTEDQI1+y7XrLeU/wJM1wv7
IagL+XEJ+GvOiiNA4a8ZW82gA4VaGdIUAvfeUv/nV7X9xOucxwvX02X0qW66+xDw+O0ctyGbzNf2
A8oxxijDXebCs/IuQTeOuIVxr/85aPPrbT4rec7CkrQ5/Xtb97UF6a8FTEULSPZcpfuJMAiFrfft
QbpwrYw9e2ZpKpkLyo6G+1U3HA+eOsKZ+WfORqt01ad3bSv7BxLQAEfcDfRcF5HsbBlS07vq2cWy
PFpxL8yiG8fjtV3L6Lh5FTShrBLZJZNpt9zM5ANZmyjcoLbBpI1RGMCtUkeRSCPVICfUYLaBLnNN
DCHpbzDf+RVaqhl54IGXcGdgAlNcNrWlXtBrQe6BhdE2BPTNhGmKgekjXeoZnn7rsq/5XrJi6u/E
UIhPDZYmjvjwq2xtbH3rMlbwk2L+tDkirAu4dsAYN1+DrUkg/3zZvClc66l2JEly1gOs/fgpbm3P
0fpBM3NKUnbxDqf8aOurcOPRYkNU+XAxWI9ai062nAxNnAemFbtrTsuN4Syjhg4Kcp+00tyRP7pB
kSkrnebF0i97XlNid8VBgKPFvXhXu+CEP3LnIGiklKPPwjfUChh7Vx8p3UYZo6SBuG/7gJmBRLvn
+LlpLY/OZ/1hl1zxrqglNuoSSqCjV6EafR5+DzkqQTof3PvqMcmrBwsXz3kwk2ijeVmqpaCuOGCf
UBUpHdzk/5Uf3P4smMC/ObzA7nqP1PxXPDkbfWHtpU6Rb5U1q/dasy20qwSZ/m6LGPD5f2uheI+/
qJUPC8qV9p4XBjjBeKkxIL8MBUK/1tdzZAKJwXWBC4i5Et//KxjqxsbPuHxD8xnyO3+lDlICtLc1
q1XblJGi5d6ceMlnxbLyd7KG7cV+5mSdIRKosmVjukUWMEOxm5ts3bjiZIDzZaZXV2SDGkCc2Utw
YTvRPgBqsxJX8r3gJ/vY5vDR3dy9aPzCmU3hEsJyDfcp8e8yswiOX2gZggZ+WIY15bFiab3R63Vn
TZFzoB4HQ+wVI9ow/H6YocyesBLrIFPh21loAYQU/7lBGKrfGtJK8nrNIrxCuATbkXBFNmmDMIx1
KiDKAk2zWUiavoZvIdzb1AWR6bnYc3zHj/xGSpInpnJL1naVvQzIL7HQbj/9hytk58pJjhGHSWnq
ovOPDgI9cU+hHrVHsIQsXGlaoJKz1646CggRP6IoeipcFdEmt6+02b6CZENhnRkMz+M3o3dxCY6q
AO6gduw/7rSy30E3Jgq5B8BwDlrKmw/VtOEVaLWpoH7H+8ltpi72MDy8uRd23LMSgp2pr4GArJy/
1xk63FyRqDY55aZRFlWVgzBjSRyCJ955OTXv27uH9HUgpJqSTgYBP+LWCYXQseZfRqW6DrabtCzt
dtV0LcOcZqjIdxHo7Xlg3xNZcgaEVfgFImr3Aa/SGG71XaRGU8keRNm/xHLo4OPm7w+iSNf7UgrF
pYZAEhmuMoC+NSPk7IDkAggENRJC5EobhiGQoVBxleJs9JZEBoDn6JunUO6qLNIrkfCkaVET1X9m
b0PgL/JfJgVbAZCvy/pLYAqu6TqeUlb3ksJxfcPTmLIOPu8b/1HUy2tciyghiN18BnBIkHJeoa3U
p262EIcmiPV9FuSL7kupwlZzvIYywM7jY1DQ8OLkSLP33j5U6lxAjVmZAJ8AmKTQZd3J0ss1rF2D
NlyLsR5ghYAoHAbuT0eLe5SLRxReTbV5bXFs091gq8FeYWLdjHQP0XnyCcGn3/9dsJUU8kM9mm1i
mNK0x86WGktEiGQc8RW+Hld8jmwDuZqoJlMDXxXQwUTTK3pDctXfDkcBb7pAZt41whUenNxYv+2B
FaKPOveJXgiHHe5Sr5PX8V3ZYixrXauwdHQp/WGbSHnbC0JqsZFsI/OosC/eMkjcrAxFkCNxJZf4
CkGwDyWycH5oCwuhkiT3myg+g1nHqYMjEgwhKUA0mRX+URLg8l6bbgW/rQ292PDkv6SF8J3wnXVj
Vt+OMwT+da3XfLhLYCePyqhIaKZANdVXIB+q33TTJWqE8nU0kREPPS1BVer+O1NAPGjb289vt2Db
DZPNKuN/fvZ7pUZFhCTbNOm93k9yMdXzPqyWa8wnUwi014Kjv68Z2lTh6xPB/1jCddamJEy2yPPy
zobPUirJoehikv4KAyaHXLpndg+v0FLIaV/W1r/CUVKCm2BxU4BrPv8nTVWWqveohuI1B7bjFH0a
D3qA4gqzjf3zNEOjzMUdhmlLMTbw3toB9Ghwzmob8ag8UeV5Bgi0ihbAjQuBnplQzQG+/Nbi1MFd
6yUHLbkKaQOlMcMf8y8oTH0J92Gx5B798eH89fT7v+vmZbKZRHWth6EASLvc4vCtLco1LLryL4Me
tbDT7INpsJ6BxLdr6p+WBDrH0nJSs+g5sxFeUlv+7jwkFDQ8mTs6tufFEFCyfR4bXZIuuPcYahu4
tw9zssvsl68Uo/LNi034weTlaEdAJJDmxTU+XJWo+8xgs+RntqmZKNUbVmoLaR+NPuBMYyx2dnfc
mXDP+hCDeQisN2S/HMxY4UB29uPb7nu9zO17tjqGxtkxbFFLTee0YGX9PFgKa2CAgzHANN1xUtIV
QmgF8BkzAUOsGtP3GQ1BaODLhD50fPANSAkk2yp3FMK6XT4wBNMK3LWY98eB8eQt3pKnNcXs8ftp
pHz8k6TW+134JS5se8wku2z5IlvuB2Oh9oE9MvuROEWF6kYYrPbzy2kaW+bsp7JK2dhEDOs99y1H
4Zc0NxxxLAiTyknY5XGD7qvBnhfB4tV9+UqZExjbtw7qZbZw7ejjZMhi1jdkkqWs3OU9H98eghDm
ivc9RBET5Q8NiIVdeIQSe6ca9D8Fy31v6fOacK1hjEk9lm85ITdM+6T+aSNWLKE3P7B+xgIQtlTa
M+SDEapM3X12ZOhu+t1stppKZZU3x9QAHH1DtAo74dRXNkobHaqNu4BDnpZvjiZpFMQ/wlHzRKEh
2xaFPsc4nWqNy35ooOEzZ4IwQC5jMKotWftMqWjBDURW9i4A55e8zkJfV1lAWWwL8PEFY2Wq7I7N
BuNrKa32sYvm5AReLYYLy9Hod/hCiXlUQyaPFGw10N4xUIlqPdh9rGTqs81fc76NyTSJyOsB5MIg
5JHRYkDh6MrbziYK2tciSSfjTRieWL/kPYd8Zz1cVkZLSqLoqvWtm4vRAAxHYaQstVLZJeoxy3Lk
RFpl6KU1PYechCQrC231Vll/EE2WuDglny5Hpgr7HnKxa5jsL94ocP2lismeyqh6o9+SZfe3MVVX
L/GyeIehlv4irzVHyFvM8hMU3nKjNsbopYHHz0K6+weihXNZJY1kTi+khZruQTUFWwASFoke/vdR
rWUISl+F+Q9VvNqi+0LOy+39tblmTSmlnZ8+BSzJTOO4zUQ2J9+Sz+2FmlUiZHIeGyUP5KvXf21O
iy8NAMNtgi1864iDn46BkDQxyCCgUgnX6vU90rS0Zpyoz2+TIarbvXYf4FB/kxp5OLGtgQ/3g41f
dLsmWha9/s1o/9qoyhLBKXTTirdZpFW9G1G8L8GSj056IAy9VmF0o4Zuqpiq3d9fyQfmRyMEwV9/
oYXFVFwdKssZI1Mx8qbZX5jL5/Wy5jNRh3yM0PkEJ43tZyRKHK43rc5TiheC9jCV5yxyO8zHgOEx
Smu8mteaHYEOyZfL6os/jTzlJ74wK5A99B8q+uYcUM3J1AqF8bIwZT73TEtgKEg1Bgja/hqHSc+O
8LV06f13e80xtXG3OH16rEo3BG749Z9ULKn9F+zs/nrY6hrPXI4ntexVKwWIjk6Z8DMJ3+Pg9hx5
oC0eWcisNj4Em+dNo8FpRinEzQW9+wIz2gzvfWH0I6HVa0GFajQFzDhv8ocyvK84KMEr+QsiuK0l
AKnQZNcFTwTxcvmrrDqC/Qk0vByigVQOH8Pi6YpgfHBL8jDCRZX3LnRWYkjx5z2dOyrcTx60nsur
N2BXTOnbwQqaPwz4LWB1BCwrT6bqsovv07wOwE81YaeA9jp6nkmgPtwp15VxkoFnBMTyhAjKUXD4
AXLd/G49snlkkvliCk/6sqSD31CY9jQJZ1MvJrz3YHSJDIXRqe/nuwZ7f3SnzH8W0GnYaqo5BNAf
qnKmMLXxWgMOTqpGyNFv0jlte8W502BeHhdt0nv0jTJsVPGpiptOhZzXEMQfdREnOC4mI3QONRQJ
FhcOm7jMPhl9CxGrdm5iRTT/a8MFUc8ZuKHh823RHsz8Tj8lgCpbrWlA5tSRRv3hwYrzFv5c+vc8
OipMQ/5u+UNFCQS0BuEmLgySr5h1kO0p0pMPCp80ck4+KB+c+Q8HwjoKekNnrApDIMyfH8XG0e4e
qCMW4F6cs4Afox5KNqxOxplMmMfYe2xoUL1iNvwVcsE07lbokr+10v9MzKjpifUG5wVS9keOcJ1N
ZQV0E5Hp+sFTwMJttc77+dOvtyGV7UK4V66clAtZWKeVFkfIWwot9yKE9qSlcf6cbGoTJzRmoBtt
IVtUDAVoNdappihqH9ftkvD50S6YupuOf3pKJApeus9cLY0Rvwxeo6EsJtaQrOCfJCaiPDsWR55+
uWdvfWhnON+l7JdoVsABv7kuXub+7JyPrcZgbfwFE98ssjbJeQpXRw4F2hWkV5IEvoAIB2x4pqTa
KWXiiUyEnrObcUVRtNi9u9ICZ+D3+sP3g+z9donApnoKvetrHg90oR+z/shmlcIjeOiGEHvtmve8
875kwv7EbNJcQbiwu2G7gz817BNOcd2U5egmjSZfx0duz/eOF5rGOL93mmauWsHxds3C9EodByu1
NRm57Q4vV0uQXNV/GaWReRfUEeDaRnOo1bf5jvHVUNKfjxysrDx484fxhTVUEVNZhjenRrgv8+9K
NCzpXXJ442jhvtDePGu/O9dkZw4OjPg9FcmQqjpL7e3KGNDF8JsLAdZdB/NIRY81iXX+Y+5KARe3
4v6adI/nzElqg3Pc/KqSdGy/vO5IOnPH6FBYCC1rOvSvyoXkItApEzp/SunbG/S5G/KYucrJQc6W
rOdPL9LOCQb544OZeCwOKE9gpUTsDnQIqvQWpnZFSLzRV/FGQGgGkzcNRVJp9EYQU056ewjuIGif
wye0LEYuQElcQ8Md0fnqG3LlcLuaFHI1A8u9s2vdhr+uT+8a4BiUB8/3c2HDBeI4fQ/aAua6XB9O
/ZVR5nZC0ZUdDK+yAe0eLvRYGx4p4jCZt/bY1DXJGeYmHgKuzJ+TQvMlsGpGFlMljYfPaZDN2Rwm
SwQWEdjLdM9Pj9oLi0fC+1hKVF34g/+KY3sIKx9Hxp/6vK3fQaFgmwDIDymd9XvDrCShZQp2cHys
RzG4kR9MWqgZ4z6434TkLB+3Jx7k1ZIgSw3dnBmO91XHU6JY1WiHrTbsvEt9ZmGqwD+FDe8V+8k1
syip8HJ9sNIpplevI/bfZWlLfzdisgrZcHA99/O3zkLWQKTrayKjlLfoW0vhDJuFFJgplL9Bg0Kj
5SbWkCd6z0aapJRJruRlkJETe4lXTj0sSsXZIbSYl9p0x/VuRqGp5MjoZpNttk5Ym+9SCt3SFD/o
8GidNCUnmD/PMS+lLog65XeSgcyu3NOYmlYK6nNBugKUQhA36TTGQKS/d+z0VKbPGMX8k0Qn4YjR
kN48QgFstLSqFCFxW3TWFRP3mogFj5M9uyi50tiX0s25uxfiH522ytJGXSH+DeFVphsqZkHPGssG
Cl800QjR1pBpVqFwvHICD6j+i1TQLWmdJBWsTxKqNs1y5Fn8BsYnfDEcq5hfnrsT097t4S09kTWv
0J9ptInw8G+FrMW6Pn+nwiJKZPC1IQ65aRpuREGizVyLxoGC/weHy4y1Id2O5UJYSeP8aHmPu13h
W8D9IWSwxqtfSkbW3rNSlQAEKfiTHA6ECqg0iQE1eYyDsEb2JT85B0pgfKk6CZX5yH3z6KW0BuOJ
0J3CEZ2+xuQ3SMwg/MHWvYW07yNCPqkUDR3JCXpohPB49qfk+g6iPQ1XCLpXBQX1C4ttbmZyCIEX
nF+LipkoFEu0frjQtkFhklgZWzzPI3K8d9DlpC9oyREL412zZmHg+Rj/BmJaSeNhRLJSPAwBKBQB
m4l12YjpnBxvgz4BI+di7unF5mLcN1XhtzjJf1FeSXOqpqMdZWKrTW7ca5i4O28FcmAwZTZI6/kh
RA1OPXSLDNyNDuBjyM3NCwanG+fLvI0zJxiM8NlWfwTInqd5E5AYHzZAJzkYTglT2nXczy6P8zdh
fHghTu+I7fqdJ9cmc4mZvM1Q3mjgJ/k6N2nlG+c6hdkFyv8hgyEz30nQCEEp2HrJJ+kIBDOA2NiZ
9waqIrvuqUJU0XAOgmIGB49EGBK4s+ZLqYKsxewUFVuSpzYdHhc4kx2KYmWg15cn0MVS4p4To2Hs
xVoLxew4pAE5i3ZfDGMx16jS5Pbt7ECI9tAQcfhoqLsq/+gf9Wx+BmQ+x6h0Iyi4tg3UVcG6DvPg
HZjhs3sEA3WX1ANUSTAAx3TvskmGEj4gsbkcsI5pUUYum94c91xLd/EfE2AQUHp5hco/sJW1ajpv
LzbHgF1uHOraeDls9bKB02ZdC/of64ODGgOF6vlzzRB1uIRQJ9YzsCgXulhm3jM6slv9Zj/O87zu
/czFVF8wnx0CloAGhtyF5HEWct+RTRc/SZA6IzbBz8T/b+mIGgnrQF/0r9B/ZxUAEkBjhtP29KqV
cvzrBBzNgRwzJuQtDcrtGmLK1IA5sC5J8XD4DmWKgJVRtQpYS9X0WBZKqmFEjhfduB3nd2O0quQU
trV1TVA2WF+XOrBTagYrau4gBABoZihdtoINgyXyQEuCidlOfxyittlbc2cC5WhOWSvM/LpBw51C
7rabwxBAcU8wI377mHndEfv5jnGPnLNr0KxFwTBVm+9tPYWBYEqQepxgfJ6pw3jkcW5MF98PH/8t
nm1duRfleGCP82NjaqIWIwiXVGuUElWpdzy80C4c0BwaeStvZD7kLfaf1WZwJYgnJblvSWrOEso1
K7Foj2vx066mHSUYBPu52iDLybZp7IGSLr9Tbk0lAawmsD9/isi2BHLALw2gna0e6i57H5w2qgT7
PkWnI1f3MNBW0U54nQ5Q1YGI6cajTXLax9LCUvJ0Pz64ayD9+iu/fUdjFH/fZLEI2sk+g1wrcRFt
uGc36Rad0oDnIriXCqbKG9M+rGXuMDRiObKuepLou59EjJRtGU78R5qqkDAPesbVvR2zeBk9lMAm
ScZH+oPTkC4vhth+M2mnyPb818MtFPn9S0B4grKhxlKPdGAvR9HaarO3H45/Uhx6zBxZQfx2iZzu
vtPQlFGRP6io9YE3Z34/wqUePLBFT2hDqYuwrTYM7fr3a0OpO1RnyILOxz3ak8akLOqhnEtLt81G
uAhTklECmxtkxgBEyeHu6fUIts2JtnHE5216Jbjq0T/BECK7bam2CQvk+Zz90EXuh3oKzcQU3fQC
dziUiMOrGAIt2+HJoTTVQaAMZwoCkvspPlwPi/5q9P9OPjGFcv99Pstt5IZXeRwONdX5G9bHlPAG
aVCkb6lRvubieDLKRK0NUPDWrs/RPcTTJ1ENIbv1WSFYtuLfCiuSqc7WE+gvTILIt/W8nwMWBylb
4O5pfJKzxy6WfztX2BnuELPt/D4ni/Fz3BW66UK4ggS67S1aVImQZUSiGPFerQpYT74fH6sfk7d4
zhdBbQnSW+IJX7xyFDmdcOE9/pVM/qu9XjOfzfm5IDerKYjjTkDM+ffkKKTLD23xYYXWWee8Kwwb
cLiWItdzhN4NY4jVMC+8vbbABs8hZMVVI1sB/Zj+qmT+BfR/r4PnTatBwHnh0JbtCI+U/euZPqXH
nvTcrBay8dp+wr5WQslInc0o9zZNEddOd4TtCH/cCavjyd5FuUY9dVwHfCxhghuKDPXPepoCxp1c
JigvffdJ/danVt3Z+h7kYw+DZh9xbDpCLjhS7b4yoRZg9VvpFFuz2wULYqtnYfmLN3X93N9ETYs5
T2IuPXK7mg65RaSOiXnvoVxpXpDc69++cP62NCzLl9cuQtiF8GMKBWUjjiOWxNbFr/GfSlbctfEN
iveyOaLZ/oZzkz1Js7TDDv8iBXmYQ1raGit0aSXM9a2qxQYuzpYWtO3iFhbxGO3ccyi7e7CsmdHG
8ydf9JJrX7R+qG6vFDfF01PT3TE6FLQY9HaYtkjfda39QWuAEF3bKZlKhA7nuotrIA2VQCoIX6ZI
gU3VpCzmcsy0FhA+UuQlotvlqamrqs5CM+/LdtB38H2N2Cb61YluH0eRgnEkazLflGfxomXnLWFK
RaK2BsfJKHmHZDW6ZDUParvokwifzS2WzWW9kGab21z06Sgxq3lvGwJcd0r56tMVlB9BQ1YjP9X5
KOEB8cvj5FSOgJbdFDJX3/mMRpn9SW09jICixX7Drav519YwsCA8MChM1JsNYb6zMktT3VU0+x3a
7+q0TTNRUxtNwKWhtxLMQpZix+e751vzJ2foUb43EWVeB2I+hYEiiGa8TsLjZfRQWEfNCPCFQZn3
oC5csJg9bVjXvKNLqXgR8Z9wzzWvqwSdcBrk0+RQJwwqEZccoAzjblCRlU+rManhvYZjNsEdHM0A
fERFM/qoQANhNURkvW8j5+Zu1iu1oUtn6Sylo4On38uBH9XP62F7Cdx25oS6WpPbxqFeZ8bxBnG3
U/3v9WMAIWoMykOaHFn5u65FEOkVwiwNsLDwS6KNUWHjDnBxb/cd39YpsShLckfSgjHQZnGYaK5r
jNgnkRYyLl8Yu9ZR4tNuiYaEIHVkoaTf6FZN3wgtzbv2PVaIFXUDh9hOYtIENM3mD/e/A/uoAae8
Sc9otpAiSqndwLVqW5Pk5dKN1hFvpNbOZV7eweot/yVgckRgCAtwzCZ4sAj9HDvnyBLWxuNnJYFv
2QemAYFi2nyyVv+XfEpOro2XyFaeiCjqng/x0LD6ToQ9oV4TF9ihTOOtBqlp1hu6HZKiM5TTeINc
fDKvnKnXI408HsrVnoRUgS5DsiRjYY0VPeFfJtF/yxNQg4aBGyo4Ci94UQXVSSPXDqtmR1uW3JMF
9I9JIvI2oAtywIXvNtXL9zV+8/Ec8yXWx+l+J0pTLZHOaecnijvGgZxyS+jgW60vmmE3qHhiOuDl
H0P92v/MfET57FuWR4Kl8fKwP03RwSel9jLayKGVLuy/O8J4E0IBWJPkZ7DDMBlqzee63sE4kwRp
tS/pJaz41T13qI9+O4idfeK3vd5LLzAtuLjrSWqArPr6oMLsPaLxPaw5pDrnHOou8QOQZM2iCkNe
iWtk3IR+QQ5Q/R+aFBIxecNo11GPRdHgfpMtjZlqsugxj35gYY1Un2cBKMRHzZ7y6tjoZ6DxqzI9
9MDpElZNV7xQw9KOmQzCGDH0vqYcQ8eTi/vzx+9ubiNoIiSZU+YgBgfaLwQnmfKZWCRw+5K4CRjC
ExXwXywj3cGr60x0IGUAFTWOyRjhD1Dkaw90GGPgYW8HCcKthnmE3xAhTSD966toCxRhDhE44nQG
vWZC6h+s/1HFi9iNRM5VrtrQ/zXZxXUoQwoBeXoVO25QyFoYdnH69ban0C2oc0uQ8mwIeE4T/ZwH
QzaS0nLq7WGogLiI1vX/Ks6UHVL4gZ8WQPk2QuKdma6nU1JfNWtEWnMAiI3kBwU1lepbLeb2+q8g
rJFALsqLt+6CC6cmG7RAoN3bfWh2jgMvIM1LxY41zzxuuu8839nsuMkXAQR4xKRR2ywSbBn6cS2V
mlJ0vVpygaf9KvFZKN0HPUFBXiU/aoQLCOrIwesHYhbQ0SNa5EXGe4SHO0qx4BaO+BTESak3Ed5p
uGHrKfiQ8LLwUq8xbWAkTMt2nMdHmwnLs6MIGkNP7jkqqBRsK6RzJZ87254Oxs36HxygvL5ySVON
sn6EghaQJ1CAVIpg0yy69cqmqRprItF1uWiWWml/qVoSjslrVaHOfdWupHFRMGLmAleaMxzEfGY1
xYMDzNzHUVNeaieBIqrI4+GC80I2UbggXiLPfjYllu3taU3YoeZrxQekAcnNlZba3di55HUgqmNm
eyNi2CoVw+IJ6jJM2bC39KGDH9+yKmuG+kSFQxacRZAOznnwOTHuPCw9QF0kpbCXD4bYEfTl89x8
8t8bHC2uMzopp3CAuw0FBfvTsjkaxrF/fo0dBtSVvwSswLy+BXE+zaH3IC+bK205+0rMP8d6mylk
5bhcKTlaIi2iHZhxRvGMEH6Rf+sPC8ZdMMh/mLrSUKvhbXCDSgU2v0tNp07OUg9qZcqFU5gqK4o6
dKJehS5oU3VUzo7q7Ji2EkoL8BFkmoncUviqCHwoRiQSGpicvaZExMApUUmOo8WmSff5e21q0IRq
73DFvjagL78vC7Bd+Cd8g95WXwMpQjq7tcLas5EIKNmc/k9Xe4PSF5gkpbyoucVA+fqxKI7/EH+k
RPwN9uYDJo/q7Z2tavdFwxkZg4DALWM5d4Wa/lD11w0hMTihMUPzXoHL1e3Ox/6TAS4APDcunBi2
SPxp8mQc+Ra0/3YRV6QUrkuLynD1sWBTsrWiWbpaINazMF6gSGh0qeqtRApIroKqZDnWqwB5Cyrz
M6tK3B9hLwIUYNYFzxz2FXqTbJ1ONDBncZr7uTtcXi4fuzaovdjp8QHG+id0n+WRLWJ9XV9/twmp
T7Au/S0E83SHeCXGShd4yWLAFWDtQPtZ/3tQWHa1PJPEBD5EaTP8kxmYA97EvmVyIGzRlOFub6S7
2jKVgwnS9tA72Aa+nin1UmYLbEk8G0N10ort9jdPWOOz7Psq+VQJbSIg+L47XQ+kl5D/nXhdi7Tb
Le9C6BNrHoSxpJaF70ni4wI2yrL/XS4XoISGOLNpvaSndcgWxdZhVCMRzXfNBx4m0w6AzueW2i7q
V8DqTYJ7887rdiVF/slFV4BVol0JKSOu4cEmPFti74eywF0MAsjVwC8miYIzP9UiXh5fPXGHchcu
QhZMX8FT16GwBfpj0/6xu0mloUtPHCmSpMvMFvY8sNL0xu7IpPMw30nVPykTFlDx77l/K26T3e1I
2AmzNyubyRdCzL/SctPUr2Ew36A9TvRCDB5aTmvox8gZTkq3vwQvz1M1B+lXnIiNZlDsV3/8bncB
S8lHb8zx2+bZDBA6LrOm8VydEGSIoYmm4fTHqDsRo2cs6gdP509C2nk5D2Fai1z2m1zSbcXVRXtm
rvCw4pmRXpDp1Ch70mGrv5uPzIqjGZsRqPoh7yHcWwtZpLA+gq3w6MiotvlAp5EuhKcYnjglse9n
c3+jqTnQmH2I2CGwdhxLgR1PtuGeb67Mfj3XNwcfhe0IMhHeBLs6GRAOoLpMzmPqcIhDvEbW2Wzo
S5wXwnuXVn/oE4JoIZ9uR38Ea9I/uQVVInAD6k+4XkRtbj1aWPL+OwwRiBT2sVtVHL/jQ6dR7K8A
wATsq1F/NvMKnSZcdZIKYSqpH3f4wJ9SaiHTgsMjEYU3ZIjKtod6VTJED+NvDMxXspWbRMHjcoOh
sbNAT1PZV/dgjP+/XL8NaBygc83E48hQ52joQH0fbMMFArdC9nVHzj//yK26TIfZ3LbHwbRT3ayI
KSnV+mJ0Mr+diqtQZ/VYTWc/Z6asslL0l1v+/avzK3MKntOOl4enow2dROi+dPvrW/ToIJrLfQQi
HbpGR0kmNRZinw/0FmReLOGmqNPWPvA7DAGn6uz/xnmD8cyEtjjf8h+Fki1eRErefwM+00oMAd4T
oJn2+wcKemDdVwXc9fE+7Htm1UzCgIOcZCQmq6dlpP8woVvhZUKxvAvj6BhVkvzAgClAQTk2veWo
RL69BZGyr1WMU4m9e9nW6GE+BXRiSSz4vttufDBqGCWZ6GqtMGAW7cTavJEoGZNHp1mDipTJZ8KF
a7mdIvaFf1q/nBcHdW4wm4eEgBAj0nF/MMEQXUSgYFo8mOBowZrKDo899JrltAZpndRQXIso6WQM
tGmjuhCBWaiHBp+SVvo4rBINDqZRdd4tir5LXMw1o1yvkTwF8hPiSOesxs3AXvk/zX2ysPfBYlDL
KZnvA+E5VQpWgxAk/t9wzMLXWKv8/M2bDV77173deGUcAonD76yienpHCNgrFjeXcqyZmhIvBLBG
Z3thoi3Vbrxv8tERLLbq/3p9d2daMHek5/+insiDTztIO++RJm9iOaUpiw/ibsanEtE0PNbHp6ml
zemsllNFsGQnfOmOsIxBBMvmdQK6S/SJhHQfJy4yXrxFenAaKmq4u1bAuqcxnzdh57zH/uUvyzjS
oxKItQ7cSQMkAa/f/inLYnz92UsID5Hg2QFpDPbJ4/NVbQW4zgpWw+Q5ZmTjPoGTHO2ABZYoM3HA
1rj+yQK9d8yjym25rN1+byjjUA32GdbVYol4iXDcgtgdkZXB597aoKlrhVmxujjVkmMiRN8NGDkt
O7SRfYXyrNVQlB8IOLYj4pBB0C8EI4JMaM98fhs+bZ2VnWVJZvegoc0URZZeNXy9kBeGLThSinuy
JiD/W+KuHYrF5LcevfjoqJRHAgHg3pPU8VEiBGkZ8LjecAlhTRunF3Xu45CrdUenNI235KNm4zV9
K0VnFtQbf0YVyu044BetdwCedS+y0zAxGxFbRzwdFozUdKIfqJC0XxSjK2ED7MNcV11Airwi2/yP
/6bCfQf0JcEPbFqJikgoBfMmbEUZyh0ZXxKRa+PItHi4BhoD+sQiKIIXka9GpODWQ9VyNIWXBV1Y
Cx3YS3UU50T1NYz34XOflYKJxtT/zya0NOCgOLc+BQdP+pLucHiW3P7dh0FAn2vkQ6Gu5ZVr9uXe
IaZGRFOQcCRDdqoNh7O70JojVwmrvs2EyVzCxu9ckjvy9v5K9mFIqH2JUBMq0fKomIoPOmUjikU/
QfVLe34oIF52k/poIMGOsh2Ujre8Z7HZ6rxbs0MGeElCP0t/zpHqfa7QmHPdcbj+hQ/bxB1tpr1b
CFo5tfsZUrHL0CXN/vPRl1MuWTrnaz/2iuStrHlUmVm85fR+a/1lLZYolaLtLmDbCWOxbKDVUEME
7D3ZcABsbmYn8nOgLs/ZJXoLEHP1Fc811e3D5E14xt9gNH9V3cn+94bkDzc8Ej5y88cQ17SO9Cku
UcEDVRMUBgM8t2I5G9SAMKNNCUp3WXbEk0VY4mY5vDID4u5y/jSrEXdkMcGacM/ln+nXPgnfKQAK
IcCZYNWziT9Uat0fT+4tXlkaShC6WqjIjC6bUA9bXD2jXYs2ri4yrUp6Gye9VoVZbZhHRHCuqkfC
2qU3uyIQ2rSO2OsMuS2Wr/7PMkN0q5bTOHZ2GK2fFlc89WxPTNvwO8mv0IaSrx5NohyjqicmCCiP
bwTbBc5GSuifYVk2smEjfXqJu1KbsZ64DUMy90P5lFTYyw/mJlBDpBxUas/EKX2A44ODN2SwTysx
74dHOzCfk0+j8bRSA0rE7uIxE0/1Pb/744w5eyHuybEtJLXV48evkkcN9OvoPB9T9Bj6VTecB+pr
0nPd1/T9wCg1Sc/i23iieLzeDonS4U+Apf9qYkb9rojlUgPaES6USvpCEVqIks2TZEZIFS5i7gD0
5rU2VhH5XC7vINgV9VD7+trxAUaRl0Oh4kPdX25Nd6FRMoOEQBjRZAGHqa16sWnJ4A4fSfvIxqcb
CED+aWp8SSeU2OKenVXF9hK1ug47ZNMH6EkEYmYSzjzZiUcSmtDZvkX3uL1PkH324BnPzHE38ih0
A2SJxm0x/pmzEsJvSp24glZQZmRY4KWHoE64ojzYjcqYihiWhS6AkqiTGaEkSrWMeifd1AZGuELu
zKPECqbWMvHkuf+3rm05Ienu4w8sV5Nh/5StTnUnzvHqtX/CjUs1yQrfhGWg6nVC+CSOrI1EgxaZ
FEJPeaaSO1136rfms/WPfARP1ZarNKHyFCzJHFzzW/FHLXllRMm9Jihfx3xxRs7UemAD/LXPkbwo
6TFyZGL4KZE1XrGzYZ+J7iVmrmF2p2OtYNX+yh7+blSKdZ2PUzV6XVttCXer/R+o/6btGtY8Gg8A
GyvwDA6ihatpYYtkSerQ0xwbBrv9X7HVBp8YqoJ7PymF4ZGSWRSPSAF6cH0Bmoumevk37inszcMs
dnjq4KKjm12rtD/8lhOXEGJg0rGNTud8YGEpDWjG9oZb/hFyArWdkjoP7IUMponinjwxAgSstdj6
bjDL2EgVp78UYeaVuFMCZmVzizagHkGe2l0BSzTlJ/V2lRgNc14aCfOfGWU6cnIKssGSE/c5LD1S
6pfozHZmLGijOeXrEMea/5RBSbyuBS8Lq4h9MivPhd66GOe/Doyp2foIqFmGCGBfR4Voq/WUiJEo
WuXaAxtBaLptYfVaqUdv5RecNb5TmLODUN8WSdOqjOe+pWFIPlUavW01pCQ3GUHBT4ou8ML9l/+n
x/K3+L9wy+9FTn+ry16/YcAv+aexq1+1T77AVGourA6JsnKNLAoDvjISYm/vVrKTgBhsALJrgMOO
fB5XCTT5n9WazR+tzhwXIRuO29kn6PMIVJUoM8AZ7g51EY4IMcWapWd58rs446uDiEb0TMGz+rm4
/s0XTjcfpzAYcbS8fHQ8y08jf/pXZOctYd3TsuoZ5zCgJvxLz1Xz0l/JMgaa2K1r+iFucU5AG/F2
SqfDS0jOGUxBtgdtHJ9pStu6Ny6wvaRTgbMmdfIf9+kssikdOWOTPPb5MmDweRo863WuqF+1w1s4
ThOXlMf5GvD6GcSvbDTkXribJE4x3ocgSebFRvM0STjO8xHIqOaOOaHV4gr4aDJ0Kiou/73fHWki
ZYXQ/ajO5WDKQ65iPJuz/RkyP4omoRgFRlyCVNk8ozDd9Qd119yYBY89KFOtyRW0nUBCQMC2y0Xr
zIsHG5xIkfcN4Eh9xzpsQk1zViLopuTDC3E/BpTnJPxGvn0INwyl0H2csEiYhreex1Jg0HipR98h
HxZcF188AkFtN7SNZ5CqRgnR9kZLj/tMDFoqvp7M7q1W7ywii6JvAUsSQJt4e6FsrKLybHZuDV11
/6hkjP4LRxri3vanDyef9JMTk7C+q+2sfBqmPSjx+/EkCp54QOjYvQM6DL20zgiDp8hgQSkcjdGy
7w3PXrFJOo3Yv2ngrxreHnQTNrm6QWMxnnkXd/9OAa+m75nPy47QYOTwUL82A1w+Ydn0XESPXVKZ
jij5iCpi+fpl8OKih8vN9OqLTuUyBIypCabL5XJVTUpie4VbOvQuUJOLgtFOeI+tjVdwbonqGy0G
tvMpsosn4p2xwMaUD5qhhv9AyR0shBL99lgi/xRnWQNr83NVsDtQGS3AKl+c0EtXLaaq1vpEvjna
rI4nXW5KYwXr6HPl2rv6aSvvklE6tMVE8EG19DmEHLhpd3R505lBN79iAaWR7zWFK5ddz8GtdCi/
pyAnjawTZ5V7yXJwp2NFiQ7SzRKbql9Y0LmyWTs4mghBWJ41IuR6gh3WgqlZTkwxHf7kWj6iAEjD
isx7D+NI3EMLAz9yf+URxEyyob85dLGPntx7azbEtDCV+ZiO7fByxyzMZTyUW0wypde/493p/2Y3
/0p3tctvCw2+5BtQryvcB3IlsPlTox0dAZOVPCbtJ8Wm3rlHlrzuuXAPWuYb4r9ajyQsshfv4Xhv
Xpackessrqqi8j7FzVsNAeD0WQRQJd6ZDH7vpQSwOW/U2jMJuIXj3Zq/dHyWVpL2aLoROdvkQASl
2gksQ8AKDJvyveJjO956P31LcL+n2JZkDlYaihH1xeDMGMljYf07ef3n8wbi2KQfQd+iq0cI7LmC
e4fIWfPCKiIwYZmvJTj7+qZA45PUEC1RFdiYE85j0QjEjBuN8Es9rv/et5kg9F6CKEPmuh321KcU
4pqgjsCfwLed94hZubaqFKmAcXc2K0xBwBhz78zSV4PHD76hqGOtgQXn5XimWGxMBo4u8UtfLP0c
Som7hcod6BGisaDvi1/QNrBDkzLBCalC6ktYQhYPqwU9INP9gosSGCdfa/MvoBJSJ998knmKp4On
Z8ZmIpFx/oeMeA7xBhC2FHk76SdH7Jfig6oqMpGQbWLS60d9sVwODcVPsF5nbT0P7ufmmEqdvWFs
SJ/683FGxz5+1G86mDgTB8mntWt/2mzyQneA9f5taxeYjcTHKUlUeNrhaf2fj7Pd7EmOANp7KvkR
O6iCsCjUqEowRQzcCnjho/Ln9AkNJsEYgHXsyQ07ThKTywcHSrAXgWNSUmMO4nRnTpCKAGLf6Omj
fbojT1Iloibmx2dxiEqWBpXT6phs3VeA+erhzoPg1Z2v3iwub+6zwPG67PYyzV95Po9Gj5w/SuzS
DOdqAOcXnsSTczU4F8JUSZgcvJfieYp4Gfx4u0fqqYJKJFSF5oZt0s6zh6fYDEfsP6ZYIHb+MzG5
tqzCVcnbgdSt4+r6g9H4UZgxeJdsSyccJqy5AduROi12EHMOwlLJEatf1wr7QZKlkGBf7ey4JqBi
6XYaxRYBhLGDOyIQFle0VQZkk+YxwYdknpUqOsN1z1Gq0f2lOgAylPAFk0zKEok2Juew+UX4eOnq
CXA2j1xdwcGN574hAdjsPlngRTQ3eOOHHHjIF2/jc1OkVjm6HHoWImSNg8N0kK/tcPbsArDLeSxH
0ku9DWdFq+H2egif3h0ZQrDg3iq6Ia8kAeOQilcrh36CfYpYkE6KAjpyCda3XZtCJlz83eRnt+HI
msJf+ORO0yYvnYu+HxRD/VUGrYSmT1wwB+skgQRNMIsXgI2PPqhN01rR53osVn8mHHS2Pv8FyJbf
7/8TfL2sO1eMu9jvFUu8m1ej6T1NionZMzVGUrPHHKchexqqFTIr62IygC3I/J5jrYTxCJHb4Ndn
zoUkjvATlyKM8/y1obgQNm+sKEZ5N+CblBKjoue5uz/pEL3LuRsZfJWtEcWQe6CqdkkKG156ZGh2
ICynioj7Q2HZ/brQmHt7QWwU0jUvIeRNwx8pdOh+ZSINZeORE7mtqiV3vW9czhPrThlfYLP3IHSP
ILUkROtikcMIfwlcBsjn6aLTf0WjmB8C3PorindukU5Vbim7N542AYL5dxKNT+hbJodflCBpBhFM
h0uToeAbanryXNmKyvzbwssaSi6vMkb3rkApGFogdoJ/01gPrgQQ7bPdAIwHNQNbKTyaGJSRoGCd
RWi4Ygqh8/O06Z1mVLSEbtmPcLKPbNT3KXS3NipN1qAimmqEP9HDTyFdZK1GskM6kgEto36oq83J
SSv6x9nWKlmaOGCW5dU/MK0KD08sEdC+WB/q6cuOwQ6eJllRTQTmkmJBmQBPTeQhBnkTE0WKG5W1
xIMgEd/FhUgvU/+LqiPsHs5Y8xvLy8MdOG8iE4j0VUqt3TdYFVzypxlLBro2QwIG6pEY6GtnGwis
2C7i2jJxG8RCJwBao+2LaVirkyJbpuDUh6RlPEeVuD9yY4FQysmO3UKVf8aV5fRwdykhDbX1Tjd3
Pjyr6C36vwzzrFwvVjTaMypMTdZVnRvPtjI4A6kPOkLY/S1gR4vGj/q30A8CL25Ql/5zACo/WfOQ
3uxEhfSz5gpkSI13TFgplzSYM1NEaHy7EEvrIDSNP11LTfGuL/0IPumOkNxepqR4tDnJ5p2zWusQ
8YoF6VTlTGmjcgJZh3dk90Prjol/lwDlMQSH0eMkICuFUqsPjBAv+dS69zIb0oXBcdO195qOLEOF
8VBkcfZObUopvHY3AyAOU3y8NNhymOn3ISmscd9OaM/a9EUd5C2AZoNqRyVSjxgix1YHzOj8D/SF
2nU2cWOqQck8BTwlsJUwiD/7MqtHh5bKB/5UxUocS+yDc8zqxbe4PiJ0//df7f4vKMLNAo5PoWiJ
n/N4E0+peGj4OKzaKhA6HMLrfo74itH9WA+UG7SPrPJ98Rk2OhDbF8jFqhvwqrjZTYTJOk9npJz/
GBQPU8QEZn/rv7xlmIWyRD3LOx4O8M2I0j4ow9OaMJFwD73wGzYclke367+7eHNdSRqeu8GI0ySN
spDNBh8/EJD8qRTEMAsS83n2+ZaY8rYvQSpRr5YvS/pSuYHqpwzntjAR2eY7jxCx+6IMKz25QtUt
V22L2yUz61tTM7fY0VFFArXcjyWzTVFlYsfc+d4Budk1F5tf86t6FdbNTJ/JtAAOR9coHrpLBIs4
MTFzspez8ejh58+x96Y5Zvyd2tsoadksZws6IiAjofzLx8dFBJpt5TnIW0ok84YjjDhA358YnYdq
hTGQdXksM1qfxP/yy9AVda736mysRryu8qmded+azt47MxmZlJrNsrXjgijIyvgWTF0xJ7IiEmNO
BKpeKsit8oju7JJGUbCQAEoHOtHsFRZ/J2/iBnQ9DSTv/kyzIj5YC7rZSnAq32jIy5mFATTcjJss
Ze6HICehGhcTNaHhDvYWmdbWwmAIJZZILVhOUzEHru7+FJafRKkj4KJDuI/keAzK1IGDOK+HCR9z
LXf+O3J554cjXXVXOaPNqzUAbFZczmL4BSd1rsa7xDZv/99y8r6lZ975MtuRsuk1pYQ2zM6ql+QD
R59Jo5UGTcaEEt0shFDcVy9iTK9Aj3RWVg4sebtk2Pix9KXjkbJYA8tOn8JwT3XYo1bJ8CBXAjYb
m2IicqnTmYshsxBmdxfon6Eey7v2zeYrLdAHyfkcjkeKYTTG5Y5fMYl5H9PaldLrrudNDvkqOGdA
hQ2r+BL70qtVfq75N9glYv8FWhytUIO2ar0EB7tt08auIUIcqHaqCx7TbKmWAOH4AYe4UHKCdHjb
kZYfGJlonlTl7Znnvb4vP8PR2zkOPDsUiMiNfRO9x7uLoyTWHoFeHDxjdRuUgvWbE6T8UXxu5Sjj
U9FOvoJglCkN8wXgX0iBA0hWPG++UX2mpGx54nwYabDpKPdNLnbzZWaC0uIvbudhb3Go8/vJX6bN
IKG3A2hUmP8KbiVuXR1OHfe/fXt9Jr22wAnzabSz2+o8MxmEVoOLztP0VY02IzonG6bqR+smP24J
vLH7A/ZGVZPTZLBB1hN0dhirwmUxlDAUR2GW2Nf0Z/ENuuE4nW+Iubh/ZNXQb/wd0hs7kjTMVQsF
Vb2Gpelh6YOoOehkeqFYzKayXJdhu089/+ZPLGtRm6EwKIUSz+X2CzFB0o/fSjGuKS0HH6DEbGrT
DBLCNEqVJlwG9rahKfCaasMGCDxfgmiTzPuL/n64izqgQ4GQ60MsuwX3OjlXJGdhI2tSrLKhHyFi
QQlQ5GHqKfYhlIf3mRD62ej8rpnbZ69RJkJyjYZuJ38IAm6DuR1JE962dFtvylFJ35YwHsF1jXZR
lQUUiJtFGxP1umIGF8ZHUbYONR+iU7r7Mnu/LBO9gjwtzmhKUIeCBbOFW6Dy+2DR+Bq/zYVbtiMH
maL+ADz4mBgs/JMyDNlCoJhmWS3pbY2aUUnDPXtR9DfVi5sy2CkUZtgaWAj5PcFd2AWY9QndtdpI
6fFrICSwIbIey9/TWR6LeAMUCsyKgsgTpaiPQ8IOxeSFv4lCscbVeyk6hNju+Y70ZMJlW22cbC3o
5ttWRkdzDaNPfQsc5ro6zZFtdgdZbjbduTweczrmWKsz7aSWb1h/RkrlE7VDJcelxaqA2J5I2uhf
YqcuOqp9UfVc7YcmtpeHSB6pN+naoKZhvJNC5NwgRKOfreCjdnac8XYIDE1HVzC3SwsP3vyj0uvf
UDPlUnWg4jxcoWPZwaWTjoXaIl7eqBTnr1KFHFY9tmwLHxkyxc0krvf6c5Dytj43JWZVZPt0Chaw
VERDhu5hoWaErh21fSJ8ZwTyg+kcCKkXQe70Hk+ihr5aA9Hq75dLdE8HUVX78Ycq66yJcF0rD2Wk
BKrQmo+6c+hZOWzP/SFMbAz9xcEJcHa2HzPWqFHSSkYOcteOMzfHmxPBUT5DXVRdV0LlKiaH1qR3
5T1hcEikE2DVwwzewD/es8k3T6qY9vNPYgOy6rwDtoIL6XD/+E70ntXqIs1GF4MG36sI7xtJgUSg
2D8khlmyHzoQhCCZdEj6UrpG1xuuWreOet0pyrmpIvN6GO1e6NZ9NXg7QxjwO2E9TvfH+e/ab7r8
liRww8EfBj2BkprBHKDO6BiSh7/L7h+Hpk/5lXYgf2DGT52+xUCxcCWwIkAfZoM/V+d+0dbTIZCG
B63CPnt/+gI3L98XMKFcEUN5hJPEEw+/CNtBl1NQYGyuY6JZDgs8U+1oTZVLE5aTWjOe9DDWv8GR
aMgEhh/7N69TCVn1pAxW6KPIoXGnJYR50WSvjvx/8uL2iUgOEU+BW9xNT19113nYBV6GwY0ibDV9
gfRZfQImzB8YJ6OHKoiZcIK+kK37X9GxS7CeCZwAJtlGkyCwtpU40Uy+iAuAh60UlADQb0M3ftLu
vPPDs7KZ4XQPLUAPfFzdea1uAfXQe2hZk/leaIpfOc4e6OecYrPP/ej/G0lTVTs/VA33SNLqoiEf
h4c5IzdJYALos9tcFvmB+f3cs8goBsV0aeP3ZDYbEBjxU4rSPtW/FfH2qexCbVgZbhz/E/Cu/mpg
OR+AxxK2jbU7d6kDr5oqtUC8KEXdyhqSDUt+vi/TqrbobaSRynlNUEpSgrcrVBCVK0KwYMV1ohC1
nYy5i4KNEavwfBnEakXO1dKKpGDJlCTK1GHOQnJnglni40t37kbVfdCawp7cncSlaZHpAhoYnmUi
qOVaI6JMojxLjOgGOYVs8dOkXfQ0hWyXiD2GfQRaFNSGOhq26ZKLbjKJ2yEDPW/iFXMDdErWSFo9
y7SQosAMGfbtT5S7eoMdLSsxYNXga4GyQd9hgLajtEqZLTljiWeleS2BfGVVVSHq3VoDve1Kr4Y3
n5WHf63ExpqQ99a0HzD6MlA/XS0fY5vmQnWJVWvPgJIRDtCSDKMaFJR/kQZTNHipcSyFgqcsA0/C
uvN+81uMokzFcw0D5sHzI/q35wPy+2+/CDllCW3CgQD5AjIOKzRAMQRuGG+n1IgpHMewMM+zIGaX
22HsslCVJ4OdrKTr1D7MPQcLoixPzsWLl0K+NinUKAqGL9YRZHDmYYXSQdeXYof/D/CRLMo7eqk/
zWMMbgRJdnMAo2P5enLuB8aFJnKk0ebKSpFMISMtEelbFjwmyOgfdEo35xe/r6WxK+pm33SZL3FD
a5p10iHfysOr6UYZ47cTwpCAcSj8dI9/4rAiKUvlqF/WG/D8fO9upymYzO7NADRXEubsPxJN7AUJ
BnmvU0uWMcSCP3TkIVbRWPqJPJCzsvQ/P915QXAptJ2iPXC1BugARsuxRN8wnpNqP8RpNoByhOHN
C+YKiwmbsQugSEpe7Te7f7+Jgiu68z7xLBxj2PURJaLhOKXO0tFu+nJefVMMrOXn4d7/Qsm1N71Y
Q+v1DoPZFGRvyl7NStgZ1dv3RIdh/IYHds/wY0iFY9rek0EejECvv3Jj2rFLXbMtAljJfwLrdpXp
hu119r+Kr/M22bfodZgWwx1WUemKy5TVrxBHQqYbLqrk2OW7pW6p2dFpaV7tN7or9IRaGLRR9Xxc
HUDmZbC3zlPXqQi5G5kaPEmjisq1O//i8U+dPWBffSlH6tNa1KCDTUBe6HWJohf6jodN8mvAFkfD
Au5IpR+6O57o5rmf4e/lbPAr3Y0X6vLYF8QwW9kq+EqSc8Hv/gHKK60QR2F0Yltfk3nRtcWOq2r1
r4PiYFK7FN+/DG7pDlQkzXJTfO12USlbCEsvwpOUf7tpgXvZZoK4lC9LYxuz9s1eBNrJfwRcq+t6
ce0n189PywdrtrQB5t2fXrijfs62ZvGuoFYau6g6uc7O14qOFt4yaebV/SBWi1duU/vXLbFOqLrN
/zC/sbOK8uxlS7AbOG3obtgdUWE28q/Oqidj0yxUCOpL/c857USSU13xtZeP6CzigHToFugdolLk
LVP0hmQ8UPKzAgDQ4etm1QAnYEuGjKHI/m55mix8fzohggF9IJxdZAwkKZ8RTMQxqZbrI7NaqGF3
ASpzSH5k2ilsKI3kAx96Kjn+iguxDn6aB+9Pz9dDe0cHgrVVmMFKsAHZkxP27MFFFHFpBzLhYFqU
kpHZLnTDjpf+6DdrZnytDNN9C4QTj5m6MX7ydVhDk0JRexrjdXQCmvVTlGwlttu5yUamcr6O8eVR
TQ1gYVJYNfjm3amTt5HzMRN5/wt9t2/tIz7YRBBjjt8z8ld9wtTNn6Phr6lyqnxZ71t8GwqvVaA2
60LSDdrXrru3DkBcA763Rfn9vBBianJi1qS9pPPH3oEzA8uO4D+gso/4+hBvlVG5K2cjbry2AvWi
wPwbJKHaflRpLJpMk0VRIMwOMJ6IiJDmzOadkFsYAWX/1z2XNiy4XMHUzlCUW5kxaCemDS44APRx
yHZGZFLpFtIvuQNZe92qIUOANbk1v3gAPwj+M0yAjJewqT61UHnjkyrve3zbgcEjFxxs7d63XqbV
upYicUWRwe4m1OWYXK2rfU6pQQKzGnMg6ojMv6Iq2JmexrVLjVhmVJbnOcWKRQJIfKMcX8eYTx+r
ZkMi2a+SIQirMhrZW2CA8VCwVS26qjhqbYLVPIg9TTBE5rxou+vTy9Q=
`protect end_protected
