`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13728)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aPkk/LZprZljgyNzZTGF6gcxBz
LkEl/7f+3dcASD/i/Kg9Z1eVUqTKbuNkFxjfcaU/n0d4gYLkqpfuAwkUMN5JdJT1E4iyUMGDRfX7
uODIPpIeibLVwaiBTYPwOaBMIRW+s33xcbIbgm7j1ZiFUBrmwmpRHLtpjQ5pQ35H5Wt1334gt5ZX
41s7WImrB3GZZogShjnMuW3Lnoejyyp6xEF1wXTott2aDCqLy2NFMXrwYQ0OI171sqr1Oy75rAS6
YZoKNi0uZiFyrhorIqTnvDpQL29BAbBmt2Xk7ypWcLGZnUCIiIrrf3JcfZqoEhREHmXn2nT9fhPS
uye95pfrbbUc3Z1mv59yFo1yJTZrevEsVZ/aChnXrsrzGecpxSpLK34A4wV3B3fQhF6yQhAUBPXg
V8RDfyS0IP7BDzRoO4AqE24Wk+0tykoHP7K37q8JREeFTFKqr6DvfBLSTRuShayOOKRnIqTVaFQz
Q5kH5ZyxZ/8Be7I4/SWUp+99IwrRyZIMPtIEf6JEZWw20X3ociH3B08av0Ugnn6sf7rxCN1cp8jz
ROg5YvJx8+vbXN52UqqmOCkemz4UfaRQ3AcdRfAVPln5/JExFHxPYSxeKsQstbV2dsdN8/L18E53
T31cmOVpdfadJaQq3Ck1pJz6N8GUJxxn4/budLQRarss8Uyu+cGQhXnOKA+gowipuH654yaVmCqF
RHhwvOqvuRaueMCjv8Xocy88D1Uadu6Cu5Ty7jrrj9BDBOsNvD2XbE3rvRCOO/pAE9JUMyLzUhPH
zjsii18UJVfapsexuIlCU3UoAAEhQa4krH8nfav8K94Aq+HaepDIZU+mu6x5ngykArKalc+DjOB9
2VbprvdLfeK2ByC8314SHcH+6nrZPg7Fl98qAnoW2M8TvQ/LD897ZNoCoBBmeFdhFJc3zqlrWJjs
YKnoS7n8gZlD0dA3CiJaujsKMsS4BjJYqR63gM2m2kHgvI5BUmLVU1/DD1RNNyel0LqcSrKKrKvK
fZNXKkTcO3u3rpS6E8ss9s6/Dg2WcJkyREg1a9e1knNkiPQ8PNVRHxhkpWoqT+1klj6WU510lXdl
7VVpbAM/HL+YZ491vPux7CnBW+X+jNYwuIlgTDOi0IHOXVFfIEYDm29aNtE9a/fb9dVgYdUp/omr
Uh+hxYM9mMoVLBV4TOgfCOJXGg7vqKVPZAQ9ur2Seiy8UvwzTeeJDX9lV1TRIKd+oIdaSfWB0Xet
r4z1sE8njEAd8u8/0vRGpKIgrine3yY/J/zDSPGu9T2Lqq+n6n/emY1nNponv61TJmSm8fsfy3SB
5jdse20RuGDhKN0b9yI5KMWKBSBhyQG21vuk2E7CTg8OlNomUU3BsWXYkQIJN5OUlcmOqHWPi+qF
OT8cC0wt/W3ZTrXJIyIE8BYp1yLzvQ+i72AWj2dy0EILUk/XjyiQ/uNobDWTuVNOk849zmZr+tD4
C8jHQvw7E2xdhjmsrt6l2yPdrLmlSD4QZwJUVyRU1ZJYwj2k+h11kRWEMgVo0xIY/KtgT7S/qChd
rZgbDBBJw/dMEAhnLeGWRWJc+7coyp9SJ4yxEZCl3RQncAsy8IDxFk7xQA870cOTI2HVYX3Ca1v7
gPNXmsQgOU9WthFecLq5vdf77l+DMR2B9bGi94TSNdPQSj8F9Wgkz6g/mVQ9NML1KrlBAmjJuHwY
0ecdft7K44RPs9NBH84HtSI1659Fw2UWsXzDyFVLeipHF3fphdWOEaQtPiUbpX98cK3WnssZxXZ8
++bSmybfIg5ypNE5Oy2zz3omD549OV6SsRhoeohMYT/WeTqBvdwc0Zm1CTbgrMFRVs19e/xdsUtk
Ho+2in0DM6oqi9xiXenkhVGCAJC0WATmQnhMnXV6csFV+F/7C0MapA9bGi/Luvemy23xm0eHBr9I
t8wCJOMuCCds6jpvtJbXCIY1Okrs8N5UuBp5Pqq7KJ/7jotpKFGz3xZ6kdtlwwAEiuJdf7KLJTpL
3R0PuRlKE9hGs3uVEQPRu6ojmmagJfotv+bBzQjVSeptvXkpt9aUSv08sDgn76k/tgLzXYYkY1NJ
qhrNQXFCNTXMI81MfR/YRdSTljuLhYk0z02AsreBLrndHok08sL6HsnjwRkTN3ORxZb2GIHAOK6X
DAgpcfJ6QzoAdrbPtD7I/65mn50m2rEYaGeknMKpEqoPVUt2dO4aas4h/a3rM5l6tdwVU/vrAoXM
FUtpQk23VHc6e5BCMgWe4jvcUNdAVQN49O+tslXFYtVOPev7xbz4USsSTUEMItlFCfqK3hh3stUT
9G5vmshTM9frrdX63qmUo6simx0e/uOYBK7FvzIBBKXLy2Dz+4juF7i5ZGBqt1Q3CJWnu/kdnOWt
i9xUcPuEpQdEflBpsdnpzUzpukQgTYJwcvNKwzxi01EAsFnrp1Dl3AvZ/HqI96IBmWo1G3lNDqW/
0SPDU/LOw0Cu40rd7pRCa3i5PcWuHR0TX44fafSKaT36G7DJLF0Byy4+MzVloCtrajQKl9hTBETF
G4gN4cApxB9Vfl/C7XoAM/p3FtI9+SfljhQfOMRourw6e55w8B19C0xrkEDHjTRrdJAJbPxvtrKm
GFQfym+IWOe5YTcyRlYGnopfjOWzCkA9z8ctQ4XeuJvP7RQM5m1VXAKlOYXCXGSRtH1M4gFnTolm
Fv1kS8wX6HdlALdGpuyMFpsCIQYEeLAV5wieZYMib/xlp7QrDuKd6cTf2QMbDo2u2ElZUVKtEUFc
aIEJRz1okshesxvAvhsZOyup2RmN8P/6gIt7jqvEZhYch7SOq3mifN5G1XJbQjXm5fJihrkb+Sr0
eoTjIEtHpe7dFLnHetZUIbeFvk6cRmwZoa2qx91K+0iN7EtNRKIk4hGcPt1V05v7JTVyYKZ23iFO
Qlmk0lHSwehXg6Gvxd/jsoOh6jRtGLh/rrVsiwmuzMbY+nxVQRxv9+HnVWWrpggyyT0DEqPLur1H
h2XcPu2pT3rViM2/980DA2It28ge2I7Daqpy3rnmuPmFn399VGJ3d71lrrJA3ig531LNxkDyVF20
hFmWZ9mIRbxzKSubHZNVPyZMywViWjv0VVbLyqIJfDdlQ5qMmfbSOONT/iyUTgvXd4yk890JxcpP
AdoT7J6DzVm42gfSz8zeO09Welv14/nySM21KyCcbH6PJiI6pwI79eBGpTWrM3Bf5gLZxGe8qz43
K+QhZl4t8BYTuAxV9mLfJ5jepz9kMd5jNjiPY22Sb8pShiYbWA1wY5llF26UywaQnZgklYL60ipB
DmCDSF+mquAL2Ji6CpEwV57ipEr81ghIvmn/QBa7fN4QFOKw1OZ5CgNrg/5Uwmy83+k1p2xyf2lq
OUUUh4KahBNmFjhdh701s2t9/bfy2+6rucZ+v74S3nPZXxEv7etSve9euwhWzOn9HTVdtaJPn5p6
TT11BNWefV5/MPHvXOTgvc4bEe3fZVrXVianInh0bPSdxLe+ONZS1OEnVbF9xdIzJuFx334ns7BX
2WTZJZv1wmsQg3sdJxAH1kYW+vbmELpTRFvRylC6pTaCKX6hPKGSEsjo/AyydY1rPOJlmOlALpIZ
eSQ8P6Fgha3ImPa2QXEj8a7pS/dNV4FwN8Hk8Ll+wSrazfbtzSDPR2ckcHha7Q5E3dL9n4eWLqL9
ZZ50tUp+qXt92Y3QaGuNlXywv4kCeAiYIb5aem8I1KEYGN7T0aQ7bPvPEbMkbwNbuGHTpVTOXmK7
qK4ghUc8O0vLTCZPI203WrWCRQtaArbPq5lHxq+8kTAHrxyWFDzk+YGWOeQ+fVyj8ymhqjGKcVjB
M34isJ3reO5hqQl1R8wZcx2aKmcETSqGpdnnKVXmQVQtwiBp8vR9lvqE95HFBSF2jnEB4sY2iD2T
3zPru/Na4jg6qDi/XEb8YErbxVeHbvITjoGoR6n9MlkndVk441PaD/3EQ0fwsGZJOWi+PD3rw8SG
lgJMtvZD9rJKvPaNrgorOm8q4lYTUzNsjHpcPU6IIYMepJVqagmppWMNJVClQQW8N7D7o5XmcwUU
W48HN9QIJkBvGSmnGyqhY5EIebiNVP8mgHiBU8hFcqtYa/zdlwbAPENZScqkLD1aD7t4ZKmaJCUV
UlQ+CyxuWQvE0QTwWfL01+qmD6kg0lbbgx9M5fXU9za0t2dCfBWuSL+fR5NYxiBCtdrtzK7LwntW
QTJvwnl7XUtF9G5BqDZTx/hvQLbjh3od8acN1Fhm5TayrRMMhQLeFOeLbZRgC51clxq3H78qmHuI
p8v/UhnfRTg5mhqgkiwX7/TNljcCXSUwp/GIGTDmpV/4KTE8y9OHz/vZuNaZsmE2mkDfd3g1v7C8
Ig3KCB/X3cxrkv8asbkiAbONMI59S2yOpI/QPRrBUVj/PU+yKs4LilOS+xzwMvNuBQH86MhXbc/9
EQncZMWiluY2Ac8tJxnaLvLbOoxRX6YD7/ykndg6hFmyd1I7PwanoAQobyV3f89pPtNA7O6flk70
KKBtvIkyrHFAMOcE7WqkrPl1VDubC/z2fg52G2semh/3Gmu2eQo+8E0w2YLTSPS8qCL7Xn67pOaP
SBUCj4Trj3XumrM0mohrre/E7wMqnK/fjgu+oYlBWy+Y2KAWRLnfrM/Q2lL5L7rTxtRhI/2vKvEg
EpSejlClWIJcpQRrv/tzmT9b//cnWAO/mYKZzzLSygSf8965EMXo/DpuArcDc52PEjYv9v1stfLA
phNM0ifUNsQuSAvKb4/DtvnO4OlY94nvvSrIt+Tj7Tb0a+X2Po2EzZjz0Lfrt3r6WBJhMWSRXU5f
apgdz9Elxjiv0zDZpbUFjSJsGhddw8X/mVQ7SDxP3NN3iFz8539YPQWiMyTQHAK530BPktOY5RIZ
R5rIR7Nszu6llo/zdHnQQV/A4t6b3jE/KMdTSWwpThBOGvsaDGdw9kRph3ZLC+qnHYGt7KmeKkcQ
KjS4OhoWEicaIro+cnmEgdsA2dVq4UpTNhtEM3kUc07jO4fK5y5evS+zVX1oIRyId8IS9iTt9dDt
x4LUcdTCoyBAqjEZ9KV0p5BWmf2bT7VVTqcfrXNo11ZQMwn2GfMFWiPoh1lBLO49T/j/mU5G58Vt
iBmZQykBG07b9yyWKqO2ivQLsHJcaZQ4QHPbi54Rj27p8XbjBkvI8MXyZz1tL97xwszr6OZ2gPOT
Y7mZnYOmBygLrm3jMBhKLq90phXvgq4R0qNDL8NqIR8QmAwBw8oHn9EtDxoqgXDcyc5Qj7xM4zGJ
H3y9TMF+q6mZfar7SZjLKuVxx8gz/+Xky32fH41O1mpVedzmrQNAUVZCxJdphONgFitx51EuGFnf
EodjYr/WO0JDqDq2q4H1rs4xvzV868UE2VlzMdFgAgsMVWIEQQRndrAYuxcfOEKi0uISiwv2jIcH
LbnoFfBdc7mklSZ3K92uZk9zdt31eptZID84XX+pP+Ow1Sqe7sDYlKA9KBqAeO0R31Q6m8fPqjSm
c9u4XL+/WbdE70dOJCB/nXSFYwZfkmgrPr3mHWD2NRFHSKLDFmO71ZwPjv8gSBxG2UwsOwlpvtC5
t/wwioNGWfG4PFbEhv8IlqjUbBTtIGMTh0eC1Hkycx/ZUsFiGXks6DCS/lkRF44DMI/eML2DYsMx
85prCZYHjzSuL/YyTZ6f+536CqMjHMmnnTmmmv1ZcwDiNEooGpsCiXz9rJUqYQiV6lTFRmed5Ez6
zcyzmPHFYOgnAX/RCC0iM/KDBG2a7V6+CiXM/Osrlnz5g3/9+jiMn8p8KHpDREoFsRJgfjDIXkuB
H+/1Y5YSq4dXLS/6sYQRQskvJZwUwSpzrYKRZHERqeBfAlkJAdig064tmW85ugJw4C5fmpsEBlhs
cN8EFubEqKBEFD1g7Uf3XZM9UW8pA8p9Pa5XLf4lQcoitjlmLlWdMZs7KhyFIxQUdZknaZ72kegY
cPYfgKB3P7oktDR9KX7HOjYBYzegO6032T2o3IRIN9WpHm+SFC3CrlG9Yh+3HTUUUPm1VivPIuD+
Kb18RpfLVz0F4FGv9Tqt6tWEeI3A33iarqXF543qgPzldHseue/a7vpUeorqqjO5S6SUc2OeiasT
KJFlHACx9fGUs8hWY4m4iI0qHNBmDw0PKI5Ufz6ycytI12sPP84eVf1ZGBwexHHiLUqRlRf0PO2F
w7aY4Oe2c3U7E2yVwy/VDH1bzkZNWtfh7aHFjEPplgKE7ZI5K4SUjF7SKk24TM1puDo3OybufTLm
xNVZ0oiTv2AiCszG56me+Q6TGQ3UwrhI3zPKLa5N3Pl73SY3RbR3YIz/UfajucQGtDn68egPGxlL
SBekFY79U5yBcS2rmFG/FbX0I2AEOkS/HwkKORehNZlTS/v3eRqrRCB4qE03+OnKJ4aUkNZjb3R4
HPtletXMGBNGMvuVPLHyvEAWGmSQ9aWm3TNf7GiBNaZrs+MecmDlA5dt0yJ/euruy0UkSq73J5Oa
kZp2zQcM7aaRBvN9p7TGbytUnb46H8S7RSq1YbqYgEbX25Tevx4w5wcBWFzylxKgonMzKMV3dume
7FBqf5CipehIfYppw91BX/CT+U/OzosbJiJgtL7JrGUESjZhpYdSWONPdaJeJ1pKAgt/xtJl8xQ8
Kyd55CwFaFKI9BCqV1kPoWTBHPiQTXGSXGv7Vd+diDhfRMBUjvk5TmrgvShCGjO4uMjbh4gvpKb8
Q5Pn3iXBC1etTW0hCOYEJ03DyG/c4L1BMVVS6DZQBTM5Ke9cY2G9c31NBK1SFrHn66jni/j3TPaQ
RNT3F+l8emtS0vQOPFvbkA38uS5x/ah+2ffa5W18kYcM6VQkXENIStXrue+AVJAvAKYwydeRMXxx
KS7D/E4jXxFsFLwM6FqazHVkHxN6JImkitWHOXA01VpD7WPT5fkWpD/JHLNQ0q2DKkEjA04dgea5
abEQ7l/339gvsLAZQJNfAqT8+5K9v/y0doNOq51ncufbLRW+XtkjXXbJZfqILo1dyRWmusMRhHVB
+84fd55+hLa4O8w/TdU/lFFL3EbUkr0nmHIjAHxsxV6058Xnp1zaFpihKtIEsJkled7uYGFEAog0
+Y0kg3fLPY9BHCeiKuBxi5W0FUxCyK1ylq4WTqBCTNIRzkjiU/T4dczCpSSez9EXgbLeW13VrTkA
8bXFIn6BagKdSWZgHw6TZBkxNecCOCsVRPInSLndUkfkKM4LqxtX6c4t8T35DSfUoL9/aBrot0mA
THWppmsBpPDxX0jSQ8/RG77Nfxy/TBUu2NWjTx2OsBMftAcQmXUBZIAI8h/YibowFRgdl2RhaAMb
QzBNBeNMghzcHvhmrm4BhQpnW++LKn3EC2Pj8VS5meqB0Ld3hl7gPf5e2hmhI/TbWpjIE8IdVOsZ
B1kkQn80sDhcsD3a11YL3bvQ8OHEu/KUG2JcFM1FsnFZXqN4urXwK1h9XIbIJmUvwYrlbv6xg3wi
R9f83ApndKXQqhDrLhXF8y9G+O6tdcAlUzEAOQgYt+oOQ5IRyKNVPM1zWRvm9BaeibQS6d9KKRJ7
+7P6a1kpK3QPxmpzFTbnsksadE/B2KfQ89LyXNHl99N9kD5nzuE6V2NWorpN6QzcXqMAyrl/APcA
Jo41kfL1Zfyc2PxeoCwYTd+q2KBsYzlcsptBte/f0MYofwBQb08vkvW0oAYtVKsR4f/caiB4bMD2
T+035hWmec1ro7wVvENwIv35OiZpLinkv12coKRxTeNLQiKfcZGrS/g9Tawv337Uma1EnTLUTiMw
ymzIiw1WOzkMAWWmog67rdp+20WrLxfYixgPfsOIZXb2renO8vgzkC6s9GmAMHQQsRUbIIu6lqst
OPK7fMT5uDQR4f3pKpal35si/r0hsoLXOKbKKP6mZkbnIOPSLFY5rflN6UDcoz132WYv2cjjnqoV
VKxnmtrbeZRP8h4SnyfVCka2CVrvrpFR6a3sU/kDfm9jS7qN+SLZDyRKbxnAOzfOzSIPeXNZDjrq
pP3U1M3DNpsuxVrOWgOYsSVB/4WH6SdEtOh+DZu+qDsayPM7ajtZlbVPg5XXN5gKTazpwKmPUibk
RsShBZN+yHRkLnebGF3SWFnO3ogkj9XGKnHbCE+GvGPB+ARqTiXwPQ3/y1nt7TLiPUxbX352NOf9
AItGgQufA9kGk+HB9RYYYM1vfw6KMQ0GyqmgxUKNH5AeysnikD85ux1qNotdJ8UYY8zb77f0Xjzd
SNAkUhqK/D7eQZ7z9w2ThQ9RwF057o2FafsHJN8ONaoTQQvdBLx7XRxJmKhPq0uSsoOmOGTQJauT
5MJ1Xv6OBq6eMpQ5PjCzG/Qvl2onXmbI9iNeoIwEN77GUn4vGlh6EZx6M/5wzqI5InXEJyTxCYC7
7pntbueQ3dbCW2OR6XVMa9KlXzMhqDqcX/QE7LU8Y63Cc2gnMKlcmfKfRhQxjZW7BvA+q/p4v63q
ITSNm4CDh18fb+3FcTCFyzb3sEthVMaFKrj1ds5d541YRA5vDN0LhGvM7Pu27NfDDvzhkKgAAAvX
JqYgwT5s+ij57NgernlMX9tvS8nnNoUXOE/226tDN3PMKgqa29s+akX2uBzb5zxhUy2RTBOmOAyU
uRC8+KSqdpfsn0IkOKcHF6d4BDplVf2bQOKnK5J6WTw9hTiken74L100l7BF8sNsKlCtPuS2IoPj
4N9nKznv6YTWubCqBNt6eMwvMDzYImuWK8j8QqveQY9JpX1pjsKLG9cn72zD0PjWRki6p8I9bjJ/
f/RuQEnM9wTE34EmVuVqDVg9J/VOAlUnq9R7wPS1el0gR6uV83AzSqkNkK99m6ja2q1DEcIguqL+
koiD0sGXm5GubAeZAzEkA1D0qbRiVPzFDB/ZpzQtTQwYUC7KiVbNzPfgmjCWNpwIUP3rcPH/ihD8
0V9IzKmHfjYBIFovJTlHs1gBSapUfh/KVsL/CzKcowPQP28MNzPXtDXTQAj9cylcIL5lq4VWPEXm
ggA5ubOzEr8YIqhCMD5AWTgPeVdSkWLjpRsWBIYtd1/+8BNYNSAO29/1rW8n5Y/I8+Prn/E1OV8/
c1rH28+L4xaJp+Dz91APcdS/tKBcYTB2ykoKbyErQIBjml47LscBnFiTTNLg+JrpTA+LCb8Fg1ET
nS1tgMnau3T3OR/fl9mAuytMldfUhqc+YE8z8PsUhPFBav6z8gnmZjQUv8kjXfhBUqtIw3Ra7PZv
F7UkEpLE5mFvJpfc3tnp4Y/TK8QuFPyS2wP0Zl/65Yu4uRzmTIuqn1vLOBGzmG6RCs3KzaSWnIJE
EfwHsNFSuKhJhgdJle9gQ+zCG6Nm+iv17rXMEelSkUd7ezhcqb3uf/hU051wCOJTMIENGyJKgKD4
WFQkF4vtRUS9bdAsrcDBR0kL+qC/zIANZVouMQnNrfVkOhaqzoTjMDSXgDdxkEE1MWk+JiN4caIY
eDq05xS3HcFZtuBjm/p+PlxOKle0z83Lm3saW+PUSYxC+PEsbNsW4OMbpsnfXa9mhMFvUlLyVXv6
sKFoSmW5wZ7+izGfrA5QjETtwHfzou6GTPSkNu9OjU2Inma5IB88OR7q26QmCqp5jk21EIViirZ5
9ryceOb5npPENCef1rBaGNc38KesLdUaab6TsMD7ISwWHNS6g798jqEbJzh5J7bMJqXufBgtIvq+
s47VoPFVOCdqdQ0nA53vlgCjqwzxTs0LDfJf/yK5ocDUfeCjAFZWs1IYE5TYW9ReqgmroC+brv21
U/yZar0+MWTkCT97s6FdWqnwJNLDRGWfNT9SJ4J6jXBggV1NvNAFMdYgaCcmgmAc9HuYj7laCi8C
ZDO8Z61AeJd/2tvtwWxsfhevJxC62aOMQtek9LRd2HvPhRfBHYP/+akTDeFDhUdHEDd+vsLsDjOT
sANXH8TOu8KpQbBN5Z9xL6WnaoIZgtWMWGO2vnxWs1wBqgDTT5ghmXeQDv5wDQuh08Wq9B9JbC/N
Fnw+idPl+EkEoeCUokGERsOoUwUaF1laRl+9xsCOjxHti/u2CIGEzI0nfrT4JsaKT6ECwX3L71yF
waDRABZ0iQ06zyKA/R5VgFF9K+q2A+DeCS9ZzD1sYFQ2SttD2yvyUf/wzi+Udj1jrKeVjLwr/3cX
MI8fn4vOyNqXnqlTCmfpdGOsllGEpwxVcvAAUzcF9Km18bomkYE4UOw+xc9wiZfEaPKG9QLNTCwx
jUVsx0XCNh2Bov2vrhEesHp8ImyXK9zPQ5skmS1YRSEAe05OJhFoj/aAiTSGiTSgVbOGBGfjRFvQ
BQvgSdiSkhr/kiFXHx4WxfSnXYhrZiCzbNdyDh1fnTx0sflMBVIfWC3t2xeHKN/SZzxdcC5dGYLr
3n2l256RdxiZyKIQ9luHpdr0nsqouWVMH2EBTEVdk5WrTLckBlxaI5RyVfU4aSPLce5BWQ15a1uu
rSU8xZhzPqbTrhGV1q1NErfYpTquAvf1j41Opax0VEOu+MQqG89dvniTvRa+Xe95/P+k1Tug8P/f
+dBTtyxnefrjI9RWedRNxd92hEA8FSrpkVZ8c3k1mnheRIchAkC7QeesspQv/ir4BEUzAZGYWmkh
ygwtwiqlemI8H9lio4oFfvYTz4htjWf2ZeaU8Rkez9MzMXvPimRkF3Ydivg7oYPu19aAtzls3df9
zBFXYk4bkW8HDSKhw2hsu832VVQVW7u+LQjq8rUBHiluUZFi0S/oCp5Tn5zcYakh0vrwUU5oRIkk
I9cqCK0cSP8a43PnP8Vu2TF7efTcikPzON4X/LLTbErrladjwMFWH6EAmCRhll4ZEtRbZpVA8+VQ
JW02DkOqQ/URv2nnxnx/Wd/RMG5a5CB20k9zxnfovy+uuKUPqu3OvLclCGN6lFwh8cZjh7CQR3YM
x2KEQ9bk8RpIr/EiLlJGdEj6W5NS4SuFk6BizEY1UH8lRJRkIvvXkxy1QsepqvrAhNzvhs/xTZ4v
Z3dWZUuvLFx8nCOz/0P07sTLH2JasRPVNf+WvgzQSQAyvWvVnFRl3W47iPc2yX31/s1NJXjMibje
C9KuESMqlAY7Tmr90HCX3eE8vrnLfonRu6xmecjFzOMfxW9K8JO75Fz0rFqY9u/AQyLldvm4P8Mh
0j+7nGiUSk04cK4STHVnXDxlK0iEc5OxV4h4yIAaewDeaCpu9ah+OO0LrmVVHkHRqOp0tDeNjvb+
H8cPDgUp6m9Vb2CMkR/QLXz1874cfrX/2p95JjlY0UkOVRPWdcUpV8H6tiavSP077blaAnmBFfYv
12WGBc73nWOMVJF35r6H6wIsIVVHhYXsOosZJA0XM2KjLVObqTsBgJJ8bnNofZ9s7ZYPJ7LlL/uO
PtKXTKu1VQZLGF63/bFSsLMIszUAGNpBOK+Fc/mDIYW/6Oy9FhwPa5ZZpLQ/S09fNV+Mha9Cscwv
uTP0snx4lV2b798SlqnTj6DXiQhrhh/Ya5lPQSdU8UyKN9EQ1jaP009H1lagrV7F+XZQHtTGgNVE
NGb/WBwCn4D4A9MKTNnX7p4T0x65/HZbyfOjOi2k3u83y7+53t4cVpl6EJvy8cSk0CDpz22oA8ZM
ZxjECrOvn8TgDA5aU3IJP7XHomdww9KEVy+X1+nD9kehc1GusbUoWSOZi2ili8GV6aAuxtuUllK2
2vtOmPPKRTKy0hS53do9DllCVVdhbgy+9aAF4hbzxrtanyjRyF1uQ/5ZbXM5ryFuK7jy1ot+BhaG
efCbtzyKJcCE1DXhiWbvrkpOfu8iJteXvvnxTPuh5fndE8SgYwK7UQr+KTyDmGPEB7ATaGBLEfIe
nmcNvvOBuigPHo9quPWGBW6RqEOurpKzio8Vns8R7HphGKCs6Dw5jetAHWlBbHOSug6k+YLYVJPk
nWJlumNlChVmgW75v1/ZzSa4uUyTyB9xtD4GR5X9cGEn3qYt26MF3CGCQpaR/lPom1Hzt32QaYsm
D5l7eLmqDckUXk9cKKifNmFqpQXWUr7OxWOghMuPF6qBNTQPvP2rUNgXQ7j3YsjU6i4iwooRxOrX
AlKBBoR7gOmQ5THSUXex/EOdpxQEqxR1QS4Y7RaaO8rDJJo/6T2w0OMS7L8CnkKU/1tA8dSc6Ti1
x8wTwAD0vJ3zpCeIhNuq0hOCfRKnNm5aYndyyMKKxy9UMEFiFBB3tbT/YO2thv2HEdHi5vSmNrRg
H9+MpRq2je2FWlCJX4VoqEUxSEX7ykPITvmoDBPmCmza6tcFiXwY7zwkkjIt81nfkXf0gZIFue4f
4DVJse3sJkqbk5ewUkLdViHEZcb06NIb2+5TCvz7h+ZW4mVvEh4xnoMaf2lao9jfT9JSkkpzlHMD
mRQhZd17Fffc7GgTuJ+CgoY/vyKgELW3/YacreFLauWO/Ux/W7j3DcUqf62kUQFnkD8DviigywMU
XF/441TYR+KS+7CDVtIsf+WGkk3OnkhPu9whYzCs4uMwiTiyucYpq6mJtuS/83AB7NUija5yxsib
vXN/N1poNLuiMoG8WJbewTwXuyVU4/sX7ESBVHT0pbRZxwDikpAN64HFIYAQh4kDDNPzFL12PNFr
BWAHGpkP7F639tH7JagGCWXjYEA0StubiYExN312JfQtrJVMlpcgKf/N7i6bY5D2aQVvzUC2Va0a
HI7vTD3UbhAyp3JLELyZObLX8gQ2ne3dQxW0v4zRhL5n2eGbzZqxBznjyFK/RtU3MeK+2CzJvy8c
HEKJQNAoz9hEfN6j+UehvKg5ObGsWnxbHeGp7HxbFx/nsnPWuLibFu5/rpDzcbtBGcdhMNCGS1yx
PVrm3130Q8gk800gyzo0eawHN4/u2UJQ3TtdLhfBQhd2cWWIVwgHj0+3L2XOUT9vc+n1yC3rtF6O
5FF8nGM4AIxmpHSo9OiZvNhRP2puiAv8L13Q2UoGxLwjWCneYkkhFSf2TXRUPIIa9YSjnUxTeJiJ
IBR5al/+ZESEScpPSSGlvwIlAS01nZNAH29AUaJKk/p3G9zqCIKAusNy1n+twdEaqDZFqQPeq+Nl
xzfJVtALhFr2YlV6GJgyH8/wJffS19/HQ/D4TWXHpGJprjvcI3ddg5c1UdvWD+ruH6SouplrH0dg
i1B1jfFVmImyv8BxKhJ/Z2S3QeBZzCR4YY2qDs/srtBO/Y33m0d+xUqYBNN9gzHvGFBchCXah/w6
fknvQ79XylAd0UKycUy3WAxr9OSGP6rwKa8CZJ1SEpbG9vc6M19Ad2nF+1T3hU7u56olq+nvNCNX
oGkSW1XjQqHDId9KL8cpxYBGV+C9zm/uZfTIaVjopf9YwPZRwf9QeT213qR69XRUvj7Im6SN8CeV
dnJwAadFdl275rs8FvgLjQhY772qZRm92qm1SwNPuBdV9Fot6t+3xCleUbmHXa7rFRFtE4QFANmc
GIzcNxZgH6cd7XEgw5U/TnYldilZNl0Xeu+ZipxTXLR2eDso/Un1/xD+W0u20QvwxYrbfT8JYNaC
TeYCEfxsnNtSc30kmmDAWweecg0OS3l9FLO1Wp7wwKnCvP3uQszXKp9AYumoJVbRohmUPuhbkLW1
nlfVyVxsezC/XhhN3YaULmYTCesBCgEgCNhcE8AEl7SldlH4N7hiAFQxf6zitQV+Bqp2KJaQsPTp
bOClOSST5DLHGXx4d/vI5fS4hjhl4uFw6YSI3fHJJ3LNskhhHzrjkqGxv2BqQAvDVV6NSwIpCbS+
kxjADkjTX+cE4JDy8BKyvZdCbAywkzEGLTzOT3ujH9QruZ1sJ7EBq4KyQjBjIQciefTCgUeyfhgh
ZxQtDIitkgGq4L3vXQ8TRcZyesApVoNLPweM/6yGN4MihNGx6fGUvi3BrbqG8yuHrtnUBFt/gyVS
oIm/qkdi4APtxgds/sav/lfSfeeylSEUMLueUSBckXbJ1ptkWr9tLrWnkd0QlunqXsYAglR0544b
U9jQeKYw3CklpI4nnkbL+vNFuVJD2KCBg7FyoUi9mTqGqWiWLUsQ1w5s+lA8bInzY/aFi6onM9vO
0JPEttBAicz9UIWJEr5oecCi+JcGUHrJlKMli+D1/Ngf6SO605s2xkrql9cus8khg98fP2Kpc2Vj
lGFaRun7S6vsUNwckdnT7Enj7wzWVlDjMHp9qF35Zpjz5AVSa8O13oAIAYn/mv25kEpu0wnT1g4i
YDtDqNiOHnIW3n1LPmTOscIyUh/4nFQpWu5osrDYT/YDqS3QOCa5j+Wa6d+Mli2vU2sdf6UUqBj0
LtApNx7zJsbFePvkJbGkSffuox4lUoO6IlS/8caZmBWsxDhLyB5KYuCJZiXawRqNHdOUWtb8FwRO
feipMe1kWizZBqDshEaQqAZQVXIdDEQBAnGnD5Ph3GIPXL0LrJK4jON7KsNODL5JguNuGMwxNuJI
gQ4nlrWWGCRtxoH23W5Ybht1XwLwJNW0l+aRd7IqnXaYmbt0sfsk6BIMiC6HbeamYlNxc+E6byVk
6pRHkiM5yf/V0GnHVgs0kDUJ1U2KMxZXOV1zERnU3Tm4zG+swczQbNhwFKt1kxEcqmeW4QGYh61n
5GOiEy/DJhg1x/Lwuz8yHNjrK9+w4GSdKu9bfFRHfStXjWjCG4m11Kr05sf7mwGAmiRsozQONo4c
zmIYDhWVZ1WXde0aRjEAba0oWlP0xRg/uOHPZlhxnjJ0NFwOWbvT/V8lwTPQmU/hcTUNgCbbPRtq
uS9ZiPAilwNZdUEYxTuZQJY2ZfZUZzW+QCC9w2qzlTA7Go8WziBbSoiQR4WL7Q4GVBrLDqELIdY6
AcfluTRmCFxULxc9lomdrD4xOknPI0lK3hJjY9mkGLZi/XJCoe4gSZJd8R11m1mg1eUvkqv13bP0
isYcsRjTCHctfGvmJfIiKYacabUvNgcxjQLriU2E3QSDafEtBLgDC3yey6lUtH3ygKXSBwWaxFKT
4Ltg5KgaK78Qs98GhDZg9yEYdo8KTz91T0jdezgoELvjCNGuNRLpmSWUM7szFEVq7STwhoqFB6u8
CtdbF2Qb6oCXcwnU6fKkpKdSfMGL6Hh0r9RTbeepILuUD7QK5vdS55XopLHhEvqByQpCufUGajeG
xFePttAzMTORM3HF8cbFln8TGK8iaWGkLNDqzQuKwPftuY7x8cCGZFVkecthkwSx2C8FDOI5uXR1
zH4HRGwdk9fpfnCVWgMdc1mgZdvNjojzYxroiXKkd88UZLVuGcFMEIdWzpEXs9XCF6WPebWz37e/
wD0jMmCWVuhUf2y8e9/rMgfQB47xHJJLepmhcJLXD5usjRb+O72q/xKXTNVvqjh36hOqrYTcwZH1
DbTVk4ALEhUcu2XayhpEGpFiCemNHEI3+OUc2K97tBS4rCWttw7SsiB58F+4bqCp1HjcpKOqU2xB
BX60stK11/lp9gAmcGoXdq3GZwG36aX7bKmLHlKQq2zh3bfaOleOyh1d3fzpE8x0BYz1ne2qWuh3
NQ1xFe3sM41gIz9nuuJ2Rukl1CXxuOHMcSd9dIhd8w8M85vSGVBQNe+qH0slILRkixZNkbq6vfsK
g2rEWY7g+0f037khOooYD8XHIjP+8wkRTynUXIVRnzxlix17AKmLEBLeodk6iWxbftyBWuu2xAe4
W6K25OpWSyH3ma1983crBe8i0GBRskWZv7vDXcqAIpV9Yuu/06uXJxNfN/ZKslF6fz7aifqRkwCA
QrF5WvL2IEOxEJmNHxN0kcU0iM58kGzELfKs2093jRbKRUSdNSTer9xSQqadxMwE210B9ojSnRHf
FDnCbNyWGGugDWDY5QOFLE2UDgXRA+03p5cQF8/zBRVtcvpGl4qvdjA5fURSCe9fqRLlKpAiAp7L
ACHgQ5/QnEUJS+lrU9Xvldte1vtKNjhCjos31eGWFyHztYALHbKHJU39JNN7Qo5MSKVa2sh+rP0C
Frv8xbYEmI2CzeWrnPwtzdkXVPdinpNFxb9pWCuzZGhp/syk1Hr9FnZ/Xc8sOyUxjyrJds4uqVgH
s25hKyLPJsCYNiLYUnJ9zr6mhb0tqbktjGzV4rjd6gHUZTfg/gqGkG8nH/r4961byR7g6JjqNCjG
iZpQWbTVl92JKoeZXyZoaF3agIAHIy8cMOUKCeogcXh3RMwUJlsSlRqb1FgNCBajqm8OjWyDWTEo
5BlgBpZ78IFjPxS6clrOuoGwLEBYKkfvQsDH0LLiBeuZM2VDMPnr7IAy4995U9ODzMhq+5faNJHE
L2VMcf0b381AWldYCeJcjGdQB98qwAnQGHH3PTvXg61q2gYxZyIiWEYm2I15SWkEEqATVZRnIuyh
zdjDufZu9V5KYI9j11xvyyj7dcr1jzXI4uMgZQC2r532EK03fvjf1UmF5HylzC07viniEsa9IYfa
VSFH2YF1bATADEl4eemABHCUdmJi79gNElEY8JSDOurya7ahvK6dEXNHGF6PwxaC0ZSaH+QoSahQ
aDY3Hanxc0yn5TymD8Ob5ITCeJMtEQUz+dTIdS294J7SqSVq5jbLaPwkqZwgrAaXMw7WgTWKFuaI
m3ENhe9xCe9uNIR/4eFxoM2WXDhfHZ9wrIesQB7apW7WhI2GqviNHX5GFHPbwqjnAXPurE7n66+z
DiPcuqp/xRVqnwf39FQOtIqh4S8PUCaZKC8yESGRGApWUcFZL3Du/euicm6tITLQV7z3VCTcE4V6
5S8T+EYpQsvOJx/LWnNhuFsM+xqvuJfXHZ+/LhjypfexYoqBJO+ytn0It6kzDk3PhvYmwl3gTlFv
5aeyU2+7y+V0Yj5bWkISqeOwkO+ZrEtyCA5lS/J8NYXM7wqimLCzG4igzPlKfdeNyYtyUb1/e38/
56Nvgqb+rku3OjBWwpNhNoH2UwspoEeZVJ5zFbIAIp4dAO6wojk+3d1vnh8vQno/aR4vXSJBuX0G
UsDHgKiT25O8dKauRjwfcRgOepZnNzNNBLRRqKqbc5KNzh8ZdnW5ItzIWmW/lLC0a705P/q28dd7
m7wrZ7W1utscAMA7PWhQbFNrXyPOFSBornyZ+Y6c0nmVWWa3LT/+4HhcmZ8Yo/IjEK18BBvt4mw/
Ro1EVx+tOzKvP9l1lyirutykCDqqoZKsP1boMkBoIxn/Jq8H9IAzisJMYqtkJ7VAA644TZhXkSAP
41pgQlcDFjCdT9ig9dOjVXNu1MOvYqv0lFQT6o+gd4aYkD2zx+ixRSI8ZOO7kdwhT+PIna4MHk0j
q13VoBCeuSp6Jrx0RQVjKlOD46uquCBYIF7kO/DRXWqGqGqITwexDI7XLjGowxdMpWmSXOLr4XoL
4wvUiGgQ2XN25MJc/sOoECMggOeh2kPJIGYye8PRFPLPmiHAH+ozKFzZ/g3OT5m6A3M1871NvueO
DX9+OIvC0EG1B+4VfMdmP9HY4ilVodvagP6G7osPS5Hs/bNGHa1w+q8SwtVoTQJntbuGXOhNuZv0
UHDU7mtC0DtFi/BqogskKreih+qs2YEl8N2G8pTK351mCOUrCMETDG7fsWn2kgf3O07qx0cZpqCv
e8tzNFQvBPM7qnJ6bmNuWuWev7QEp6r/2l4dDGfm15a1Vbp94XhokziyTmZ9VLwhHiF9O83t2spX
UKInT0yvn+asq8qrTpB4vp2AMiemo2WAfI5tWeMfLlD4RvhAGGK5JEtuCMXe64CQrmN4qCXlhPRm
B9RIsmVsGvn1GBJ2ktA1a6XNIyS43yU6buS2dZNwhn6d6BJulOMqguuaf5wOSNmD72m1D2Vsw3RN
K9J/uBLqqpuGSRAVenvdWgDpcjob1EvUC4CFqccPXgPYmOeLZc9UlaeyB+QnbJDhb5WLp6fG9BP2
GFbAjDTEXnM6Bm+Hm+j9jeqJcoivwioPrJJpn5/pEW/XStKiiyIaWdhhU5M0e9xG9BDGdjPv8Deo
3ouNHRrbnu4jyxIWEmjbgVziqZd1+lsALdniqnUi6vGc1uMbVV8yQ2c3O7p5jMdMLweVWg7ZPKuF
vKy6bGoXPdPJZcUCWy4vaQh+KE5HeidQbaEsacFPHd9Df7RiwpGELpuZl5qhB/CGu8jiQQ0Z9LXy
LCNcaQbczJ/dS08IAVwYzodrOyFqBBMkJCH4Z/1JrP3crtIEzuPE/AAxCWBqD+BQk6hV0+y9/Y2d
EwagRe1fDEHp7bQHv4r3QCtoesWuET3licPsa+xxP7TT5sz3OHjl4z0N8MJUmqTU
`protect end_protected
