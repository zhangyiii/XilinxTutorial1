`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47328)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMKRcNvzOG7grs/8lZMh3KNjoyD
IXsq0a+K7fwBVl18ZhYAY1e7ftc76HaRu/8rLjkxtE7Q2J9eFQSb2UtdMq6Y5VOj0vNMKtDPUUYQ
EapXijfXVqWDBMqI1nbHZOALvVCnYVQJDo2a2eEbg3LVp46PYehYmYWBNiTcT3fHf3km70lpX855
2eitSDl3fEbcoRRSxZE8Dd7GRlHBulzhkWO51Y2JKAmruWiveSfX9qxrc1J2+ns2jpzRnDbHsJzR
mH6NXg52JAzAA2Iz+0RIzyDWsYKD72UiQfEHpRNd9zHdKNpsy5rckzxGpo5ZuSYG6SC6j0QggC42
BJezzIXT+wIKKThjvv/jI1a+/VFfCYD6pzU8fCBBf3oPvXVjNKWzN4ebtRMisdR09CkJ7AOSj3Pd
t+iY+xsCZyQMM/TsdHfYDJNhZuohAtxFnA9wChQWflGRB6Xf99BhlN6gsevu9Hr8ffemU6tQxCXp
rjcOEw+TOB8t2UHDkKPFVkCX6RW8bY0bJkEA2KeuvZgVvITl4aGa60P30nSo3QN5B7/9A4lFBWlu
QmQMJhHAcrEvnKCP/tZfZ7vZ5wxObBFAuFyVU70IKOrfleKtR4AQyBlEkpvjSt+/Pj8XNxQqmGZs
QVMY2S/gjOopI3ABRCZ1ux1W7nBo1PhN0z3/H7vQ+Aq0KMICc2nwmi5CHXHoKqMjtpIsOgGc7KQx
qDmdEisg74KxHdljo3AgbXt2QR6T4gRkxfbMeome3wR/CNOPsgtcgA+cf32xZowz+agqZFwewTbg
lRzkz9HjLaktc9fzU8hWulUb4BmvF6NbHdzwMTLvW/kiQ1SWAZKD0Cmev1paj9/qI1VjQPX8+N0t
T+rFShPQAhSjB0QBqJ2iAh9TXJC2h8m0Imrxd5Y3uYWZ9EG2V0xi3GmbV9eww3963quXADHbLjUq
bCJ9488udjpodX5wvVH9sA9qSVYkj5LxCbqyKWZnvMJb+a7Dyr/Fy7QFb1ZgGOc+wTraAMDjVW4Z
VHvkaMkffzSZgFd+e7qvKzbslE0akMh3hKMgbdJgUCfBIggqz8xFmkLyPYpeOMvdr6RBqpHxiWbq
FJqrh6nyL95e84cUBdQiXCftgqZ/8fcZcq1skHoFa1Ps50vf3+Or24AO177LHyvNTMT/fwQA9Lgv
QS7/QbjAprc5BTPCuTgxVtRVYf5PJ+GUyazrkPR2s8XTfiU5I9YS0qmbgfeJdBXXTWQckffoIlAP
uFLKUeHB/hlwM/j09wvNrRKku7E5gnl32njgOZ7aHvgeYdOG9od5Crty2NZEOjNelmlzRkdj4gY7
nfKxWdEKov7h73KbN0EyTdQUVHBKCtWkHlA7QD3fTyXMcGC1Aa27S+jlvscd33xXE7jaSjq18dhB
d/nfFyi/oPWbeIx+xORSMpEce6wExHVXWRLD5p9Gqq9PLuiZjDojo1nAESmqiKph1EhvkjDNwi5a
WdnMGpdPyWZBi+TLiJdGK3vXbhfk/G+i7NDP9XfayHcfDrD/zd/C0sRs8FAB7UDF4ogo33PMPoXi
sq0MS910zI8M+8y545bkRIAg7TriOS680W5IxstqwdBAe7rZydTEsdo+gfiH5Nx1j6lpZJfNXwlM
UrbsuzUbEblYbLM6DegYq0kc9QBvuZdpN2kOfSDO71GZEWChUCvd5noiHGHlT2Qp29X9OLdgDBQn
APSNFip0ky155cne9+++iaR+x6UgpfrXE5tQq3YYHASfYdjSehuNsv0Pbg37gugk8rtMw9GTngdE
x3FNzOkfQQdEL1jt3gVprcZaJx2KcMGiAA7lgpdqpETO5t9fZzvH4rf8+NXKA9thE4iXXU6mS65U
krgb6pvJMLtvTPB5W85h0lEmPgKF3j0uwcfUgw9bVFnJ02R3clrAt8OUHUi0WuIV9D4yJuSmfbLU
zhlMV/Ur9J+A9XSNVlFBHLXrxzjnC/T98TLVguHiuv3ybmWqMk53VNE6b7HQDE+yve2V1EusTrNQ
2XaHxO/OIxs4AmM19xRFFfGROI2gpcvPfKGNAza7pwZJegt4QgBUv0vhZ5mKzq6mMrL1AeHeycCB
BaQW/kaZ+fT/JB1DWiXWsxLP3dJsZVxfJzvVD6nGx7sUqTpehC3LF/F/8Yzu3A2vNWyJvJQKeQwk
OntCFxdPgS5CnlaOOmADPf79Hc4P/OvBbuGbosmcbv3oGhcfqWe86/saZ3qTbsqF2LvQchhWT145
CFDMCk7ZhYxzG+gbinPMBf1dd9M5lTMrQ/qDk3uayyDZtBmfNp/SQltYX1WSBbGhNKrzNi3ejf3t
EO2dqcABPSX8rMTSNq17A8CvwnS0OQgiK5N5tMu6duupNjFrMZJtI2wOfHeZcGh4nk1CSJSb8Osi
YNNTyOEW92VQoiNQ7QTkyymi5xpzexvSdEeLx1/OVwHg+ZEsH4qTJxKsP1XPTESHAbvgeJfoQCLz
KeBZmZvF6lkjJjl8q12IJiBT96RbQF+XCOl4L4GRxSbXEi3U9iwO3vF8n0gurtGyhVQHXYaQ1/gR
92+RFCDYn5R+3gju65E0Yd7C3onh5f4uoSQaDv2O+vPSCfN1yCf/yUXZi5oK747SsqbOi3HhiWS4
lvQIDLVwDlKalIotk+itTv6ay0ewx1B95/bteGq2VZLUIEl6iykbH6lHK2mEByNEhTWxLrxLTY68
lS/35K3Y5ULcdNJyKdNUYx2n/QKT++1yG/PNDVGKkNnlQr/bW2vteZCqJqEJCvvlILvshrqoYPeF
2mK3a/HB3/XwlGs1k81GfI4fjgaiz7xQ1vecjhOApvXYIp5KOiqJBj4YUiuIe3DnhdKloRjjb459
PTVvyPHOIfKlJBXO+VwlpA7gkg7zfbR5IngA/zrtDheQiqQGH9VPA/K3AyFpcOluykd1yb+w92B1
WcH1zsyjSKEtcF3I2DqlULUBXDzUiSlMJUgTDmMbo3sdxhWQdIBkjuWGQkWU1TfiKjwY8sswcsqE
ZgLB1gya0thXgI+2+8tSr09byOQeFxZgeo9FysDysXa4t7y6kMUGSlAHhomJ1sAK05g8R7gN3LbG
uZed+J3NttniZeoChTgtEFM/eqkjY04Bcfh9qsJEt7IFZbnn6phXGj14BuSwtQ7emAwxbZn4nHCw
PQsHTZtH18ZAUDSWXc0x+0Uj5uDpWRrDEgOETaSRaZChjzWqT/ajoDMPGG+hikjzOidPt9/lPj9T
dTGyAcBuniXNpJcSKD8Dd1iUEW8HdP7KB1wAtRfcSOprthf7wm7ZsKW9bvHGZM6C4YStzpq44xfT
bRRQmi39VbtFfAT4vNb57WVZsFjonxnSKtW6+PefkGH0iQpBMqAmLeMWxFGgyvZdrwZbBSnDTq7V
2A7dYYtNEU76Mc+5Wg4BkzNjbGTBKUqvBnTLZqJ1AdmhX95dYsztVklv6n8cTTlIvrns776UWXMy
teHz574FliXf3IgvP/5/lYmpVYofn/zZSJJXhjQ+Bm72u/HLXJkxPUVNekecmz1hEaCRjm4KZQKE
x7OHvCLmp1Ibfzt4p0AXnOL6+KylXhG8DU73616qB7rT1wlYszZHidCiBH4Xq52ZJMQVP4Vx/YM1
BbJ1pOtF4UD/Tn8I9YqA5rDFUuTUQgJUsYee7YfZNfZBppAPDc6cOUiCP2iq1GvsJSVF+lQbrhmc
gukpbaJ1Gv/px0x4dCwiadvpclg3WDP5LCHLHbr4mdJB+OptGcWX3LtDXgEjtFee695MdwETWHXJ
O9Jm5KC6zMETxvfbfs9BLN9MDb2lQZMuEJJJwR3Z/6ph7sj6meULAEE1i6udUjvMIJT+YPwpZRTn
K5ge2LgKpJcnx8XWv1hNwoI/o4VV9vdbUWkfgdwwmfhqKfZseI1oGYbncC/Rz04vR7pl2I+5t53r
EdqTFmMxgwkyiOgLN5u82MSjNr8SOGD4T6S7Acmdc5BooT31htU1gQQk7dbZFyU2jb3b8nJhLgeP
JdRjbuOI6GaNmQEK79B1npbg426ivxfIi5OEI6e/r7h4hZaHYSMe6GYhljqWNuVCH4BeUO7d5HzV
b8KDbc7SH8deHQIqcYAnotAYLCrakP4LLA/fhoDauan71YLAEXkWU7C9Aq7k4KIIxueOw7rLMeKy
XzsULeIubJU4N86X73TbCLg5BHV7lsqmB91JtmDQH1UBubjRov11SkrKfcTMTJJIVIASdj4l/mnS
0q2NB3Dqc3mgf6gLmkqFuCApeUwpZZvp6zSX3H9R9RmIGCu+93dqA7eSBI5TUDhIfGScVBmeRQao
FoRpIgkZ7rTMQAdeqRv2qFIihkzEVhF8KFYnZsttO6O08jC9MPuWXjCx30uCUfQs1PUHmJCNv3//
lRdmvf6VLmd+DyQbIx5GMocQ/zfdxtbtD5CBIDmdoUOmClZT+SLuLBc1EHVQD4d4D8fY/KYKRByT
9u90B3wyVZ9xbpdQnkdjxSkUkOA2NpX0b26aUXkLiVQpTH2sAyICuqkz4rWF8ZSTnGs9DigffCPw
JjtGN7/Jn5SHVzA7eUmqdCGMZPYcfs8XjVyWXNpcKXqvksYndEyrrP9s9dKDY1UqNlPRWE2yiecS
RSPzevGyIc1y4zUDj1YBq0x7l/AMxbJxjUOqISkKD9ra/Zu+J821sYG9Q42em4352lMxmjAEsm4d
OC65AQ16shhdQdDQuCdc/dx+ZYrJlUFszsvAwtupU64hT+A+hhZwSL9pmFjCxFOGeOCt2EemNjPl
IFqHycD7/wSnVMLBW1gsl2sHQlTtUuFszZrLJmWoL7l+0g7MFhgNsVAnwdUjvymehaX3TkkI/W46
8V6oSRfA5iVVj+XhyupdGmyiWwIjxFu/ZHvFE9gCktxLxWDbVVbZJFcIFzdWLrHnRTMK5oePURy3
p5O3mJmRzAJlHPVKL44uXuJVM1+/nO2xcU3qQanZ52DgwGRvLfP7pnvrN6L/G/KNNQgY2gKYnyLP
5xYFcheIt/BmZDgvAi+rfxlHOeiT+DVet9TrK6Zni+fzee0fem5rZm7H7x9iFHHqUBd+aHz7hM+w
tAGFeDC7Hf6ej/AqzRikGpdCd1BL9sl7FbY9KpjQwMCNm9Z4+Jkva3M2tdY2mAMEADYwZjxhgJWz
c11mi/DSw3Mwq5X+15BnoDM/+YQoz5CfmzQS4LwgJwXMtm1LdgJTC4sU1aFOUYLGzOAXntxF9pzW
2AxIiZxSckfXJ34GKq+3YOKkR+43LP4Gjd8qC9LefBqKpGzCB309oQ5b0PnoFwK2SMmzCQT4+5El
Iuu3WvYfaKozhv5TSNy1prqGe3Tr3Fra0j2bi17NyWGnmLb3CwzF9+cBTdNGryiPbmsKJnosCz7t
On1LcZcnXtvUgZYtKbeTEAAISgU2ce+IYfXQXnq88qAvp0ywwg4W7KUkddTvueLqabme1FvLGWMu
aeAMFpaJyzlxyFALdYwChmg3qu9P264GGAlA/nKJqkJGDsSn02pZe9hcpRBUV1225g0gtEmo85Qz
SxgSk26w7SqNCMdwYOdN0jxYSaqVhzKKY/z72UlGi1Dd+jyJqFdVDDcWs0NswY7SIRV5c2/4fTcv
WQheDWOqZ+qEiVM4u8xIEK1nE7iZXfWPadeXdrTrx06WCU0hWqQI1gv1J1VmLTLP7N56Kys0Wbka
5rF0p8xlzP9rtp+LseNdHsmRLQi5d0Hwozz/K0ArFwJb9hYMUDL/ZU/mTwR+pOyC2rmKdVa5KBhq
MDGE5JnWICvPtj6wRhM+hqPkjI3NrFnH938MfKaIkgUGt9fjgXWW7YyWN2M27Iuaa8Ne/iJqiaOG
LKpaQcTFu3pJ4bnNrHSSEF/p5WHjv+VoL29+kDK/nvLjcUVWpHSA5t5M/a3zGQsGq5ZxZx9BKFFB
pU4Ce7dVskYZR9br0tYfem5WwFhNKhXT1a+CTfxbgysCneZxit7arH0wASyiF4AcuMfbHKMoLAv+
vuTcfgLHZNOe1c14pJV5/lx4wa5nmPQo9aRwU64GJg232ZYv1AMuzy80di612Dusfp9rzdhW5yS7
34RpcD2sU70IrZHTq84qamnu9J7EgUQuw1nybhmZAwC1FKxKJVgXPKouB8JJ3vO50ND01N2NQElR
ZriYIy3Fwv+3htcWXF/Zdj3f45cLw0l7V10rbJmG7I/7mrx5KMl48BEDFfxpNVE/EuQ4WrriHyew
1V18CQfH+Fg/ybs8IBdOv1SXsEBrtf7QSUI1+GibNg6OOXMT8P9Ki8ePdnmbCJ05nuADMOKvgvLV
+5Q9Q5Q+SrcAFHpw1fqKT4T+xbja5fgaShP15I3aBHi1bSG7i2Bk+NlEiuBGlKrq4PMRqMZAxax+
SWKRT5auiC3ef8U9oNuRZ6LH1pQEKXdqmlR0T84o89BsYHrJkekYZKbxQ9p6cbkcjzj0Sml52dGV
ACKauBw+tR+rcoAL9Z9DhSFh4Y5JwxGnjmMKdxlGg4y5b+PO9T+Ul2ZJ+KI37AyZXQjELpWLZBNt
nf9851j+WQs4wGT4jNdBaTtAUxlpxpm4A9e0TE9rDZ4o1ftQCcr7JvIpbcXvU1KgeH7b8UkXE0ze
qZkCdihCFabdaLX5peuEBo93u6g71YG9keLcLz7xMNGwVPwldrVc7Ixg2tS9PoO318nlKsxQTjQZ
IDcZMa7H+JPSVIqs0/M8545Q+VVJrWNJs6r19CBoCeaeVzlM+lidpqk2C2q3bdstdd/5ZVlOmXSV
TILFyHXFdWCcdI/d+fWG8TrkuAlVwJLxPRuHeWNcM2tcH2R7iTyBIyBn12Xt/h9b9Q9IrSS55nO9
cxcgAv3bxIOUIMYfzTan5GEa/z49ZV8EO8FhFI/AviP9zY8y/bQ/It7mJxjJtMqwlMeK9DdsswOh
vteb/07TM3wrRGUwknp7QW63VhSslLhOlInihwimv8QeyVGyG/6WAHW+G52gCQ79fOrWTmRkD7NK
qUgf7iIJMwzFBDJj3rmGPhbAopNb8lzvbcbdKx2ffqN0VLQ1lLMmtbPvWzX9X2iwZUjtbF4s3bKZ
z58WoikI3rC+MXkpuVv1WPaVsI/f+5+k5bCIyAq+iTmPCUEqwoRO+VrGk6mi3Z0KB21681VIlcIW
D9RN5NvnpttuoBoqweT1WZG2VK7EW1gH4pqidDEzpDKTAT+gykJubN5PKn4FogU4v3zvT6MdzuhW
dheK3CN0OBXZpVxgHTwyXVn12P1HQ58Yya0wsleH+1jv37iNaVBUtGmbGYuaoTDEUlGRMOuN51UH
795wuVlOpgFKFMWSXz06oIkZCeFn5NMycKJSF7Gj4HAz1sGkJj6jCdK4w1BALar2nWWu8/LzzdjH
LNtrv/DJE5xhRWVeRd2Dh9g0tvtyI78pJlc+I8IDVbWEi3i3gtMPrcBqAi1KHxBDvpkKJ//uBNuQ
pb6mg2NeBHjhcWxsPjisl6DXk0bMZ2Hxj7xemwjG8zyuiyltC46Nl6Mjbxt73/uwESloiSJYjnzC
2orTfzhQsIS9t/5gUd4jU5wEvjzqHOIRArPFewBWz+YGd2VvSkBvGQse8Zw3ujE7RvnyYBhsbWFC
WFfYMTiDW99hgBrp6QuoYtCfDYxTJMS64xfDtruC3lc4TcSM4vvrZwezkA0HEsZYawQfr4LkVecM
KRVpAISA6IrWO0B9QhKls4Do/rgzMkxH1p66hdFtfgBWWS+WMfXyPyV95KAevRASidG1aHk2IPCK
1s/LPHZr4HTJqoUoo61sSRDlgvp5+XGHRz/TdIb2MqX0iovBfMlbfiE/hXSWH+5fVAcujW0T5nui
2HYcBS0T6FJs3LCoYRPDgrZr5vjsT4ARYnLJ5dECSaV2nF0ExTYVaW2hrSrJgPizlCswN2vKJ21x
t9dePcxznrxawu9YuStY7SwnYnCLSIUFYm7P7QkLQufqf6kl/kex9szeW2GYyzy72uhZHPCHAd4G
DYhJTJsu90JtD/fUlPhiOMiTqycsefJiPl9GL27D3WK5gHZiuzDu/cMcuBGf+s3tUR+M1k8s8jHu
T6+22mj90rDRQcQ171ol87vBOEgLjhHwK07DiFgtixj0Fll7mzfGZhIWp6bqKb/NN6LR/7gJa8mX
FlSHUQxPYSCG+sQOjMir5BHZceQik4h0gpsHKmqLrv4f/E9y0s1M4Wz24OlJuKsk2UwVcDK7g2S7
Ym8nMiKWBVPPy7K9jqSAazswRWRkkjhfE+ZGboaC/y9yKuFRqQyguTy4JbpR1ESmnM3pkdRhbKn6
vRlr5jCIZsxZDz0s/N4+U5I1hBVaw9A/P5f2NCiKmshNRZ0506XwCo//ApA+NebfFFsVtRkrlKfk
bgFzHPpB0o6i5dLq2e4oFXpNM3kIM+iirO73exr7bwRIDZAukPp836ju7tVR7CALAVr+hZ8kbTR1
9aHmKSWhRs55wcMmxtFlVFFsZZZdXB/AXELOCugJBOeeuOUg9D6oLsTStOlrVQ7CUZugND3WM+Af
LqnLMO2BRD3GAb55nsu9FiRkLEn9vKsD1RzhW33a8uSnV+2Ii8GtpyvUL2mP8wtF7kWNTqisTYma
5udJ/Euqy6q7Bn8V7ykMjk10wBBD/LXWsAk5OXsB8axr9VhEAF9oyNwqOMoofWQHRLWwwMy5GLWH
fnzSdYfJPl047o2WkVXEdkjogY3f3VPzFMKsa0FF80iq7jFlPQnOy6AcJ6hRDjQFzOJCQ2K//w+5
L3HNnnr9o0cLUv8ppSHbvnBcCleG9VVwKnbFpYc/b+oxnflD61vk85f3/YKM1b9l+NdszNnR4u6b
bM3ikxZyDcilNRYWpyR8MQk1OuEabq6PNCbnVePDO7bUkmfJ0/RE/A2af71GzqQB/bJoPKAIKcJt
Eu9Bq7TLSVgBFZ7FnKZVl9jkYPrSyISNliBvj6goffKTZlv+8GmByuMmWGRHkfKxPhzWkNJULkOY
1HRJKzrk7keENxxDT2sQnPIWD5SimCpbZdOW1ZxyLd8BUK8cTPsg7qqt4Zz0PSnNEAARgFOKGHaa
Wmtp1qXVzbzfGDzRxji79w9lOqJYSAIHK9M4Y2bJdkllUZlZ+fADDuSQIqfooYpCxERt/Xw998XC
8sNcNo9KA+AcFkYJLFif9Kf9QrobAbput6WSVceqt7JkXSbC3J9AvAf+B1294cHLMpGrYAbrlX2h
Fyr/8RxefR/53IW8ik5Q9QW8YiRXUL21lPokeRyuqeAtRj50fhjFCyFFk9C95yKmKh0mgSDGo2OU
pKMM/HSjGsp1DBZ590GSPAWpjj86XNKCJaKisREzdJomHzxh2giwqdjro67daXfJFV67Np9ILkLq
XauOgl+PqeyhtpMMePi0skyjEg49HSKT7V6WIBwFNBVxtv/JQGUr/+7NkEEXaM5kb5MlDBJaVfWf
Kx4PBktJcGs0aouOHXLIV+PDk0K38CoLPp1Pi73WAx8eSdPuqN8scPZVTz7gjGacIhQFgFhHiEvM
zghNLUg5H7AF4clbLB3J97gdrX7pQ+dvAKrshrIVvJT/PNf5cDZ5bw/+VzqYHHReZF4MQiqmpFBX
UjXY4hQgqVX5Oa51hY/io40ELzjO4IlEnOF3LieHMPKKPOd3ZyomTA6WtvduMTAZp5tk+Kg7/S4C
ReOpyd7V/kycQtgEdg8X7ERpQ/0ItGG91C+YfnBjrSs8r6aA26aH4umtDp9YT3Ft0Cr6k8hYMxAZ
9nvpzK49T/D41GZzFlVJQxiqpDOvxdBaOh+k4oVPqyIAHJ00OLom6+7Q7gGm85l/9g3c+vbJQlc2
+9KW+g7TkllCB0xK7kB1PXcQkOpzPEQufSUrbG2smsKg0JVeCaZlRWE+qEJzW69L4D0LHVrP4OZp
3jGnfugcQhLf48lftnwBy7zfWL5vM2qKfp4RZ7lkrOqK1/J6vwJ58hBeC6TJvBv9GR45wn3YnPSy
amKMX3gpeqXgsdf4BPyGlTF9GFle8GCR9NHlm1WkhvgdJKFzRw5gw0sBtSzGob02jNX/lAF0dA9v
fg9qPKvVCqS59VrKcx44Ewi8tFYRemJ0AlvGOuIMR3B010qZXAbQuoD4Kz3CPwVhp0Xuxg3a26a0
ezwM6vJOpgmop3gApbbdipAyGngqC5ZxYw1VRX6lvTCt18uwZtmNG6EWp0ziII2nyDpEYKdBmgbU
mVbQVd2zHx7cPWSnAynFzKqY4GM26JXMhfyunlmstMtNrDeb9H9Q1tFZK0QmudXdSq0hlPbTBLWz
eo1erolnaUxf22PbT93PUwG/zk/z8oxcaN8sHpBDkJwp+qEsqWuTHCwN6Qqg1/vT0VlnivAQ1yhy
UjS0oCJ8CI2jepOkTIP1N3+1N1sZNFYDom/SNslNIbXHQnvYsuys4BplTaoE+kpEMwaimoIZt39U
uZ4YOrAhESnKxNV8gLH4BjLrGCGNtMWPopM+0bmB6m3hVpO7EAF0qUmDJBxf8VOPMHKHJ37VMEsx
rqn0b8pHTwP2XmWUBh7PioiB03OmCLq1Tqtri0hZWLrT1WqPG/8wXjyT8Nr3OnVfmAk+vbPY4uD6
r6bmdvOkMJVtltHezck2I1Qg+x50rJqYViagBhxGtp9hJxpIb5D6nZwDtDIKS++vJzxS3Q9hIUjS
dSFmn4Cs0s5SVD/PEibTim/A5KouXOQsC2iiAZxj/BFCIdyoNP5ldfI7sfOjakPlV2WXatf/3ePD
P39+EO+bwzk5qWglSAjZPBqsdM844fkhxXrj24/6CfDTwE9EN9JDECZLag0W2u/Acs9mRtvKisrG
n0Q7luGwnORbzQkZbKz3SweXFmELI9vA0ylDlLdCllR7EIWmAaLGuS7LkDMlvVPy05xREsZ2V36B
PgJb2LMjIFhMEsv4MTmJVvu996b5F24ZygqUnVUdujjM9imD5pjMLbH0K5+Bux0yfHyrn/YP/nzE
ej53u8ZkG470vNUCmfEIYNKd6o9C0ccU/kZn4UxDK8mRMQXomap5zgEBRQjes15mJcguHqnjfXkU
ieQX2dv/PK4oi/B6d+mUVHnCER1kpGqe+GAYlQDYt1XhZZ7q/QfbyaEPg53Jw0y93faKPxOt9/cz
cHpCf6j2HqNMxSEz5pba+5muT0XbO49bG9pqt6loJ58dqEwXfhQGR0tSac29TP7LafFnPvoqGcl+
5CR+muus82fly6RVCnV/P7iPu3bho8O5pC9rJh6Dkuwlja2VJdGpzJS9rNJyOE88mbEdr1pfCl7m
uDkUKDb0SWPhk86+aPelyy+HvnBUb4rAP32ixfgoulzhYaMAgntGfKHHangOpIT+JFikwrHhysOz
s6Qm2otfhDbdpFCcem2lRXXoC8JvbmtCFrxRhwMjfbFK5ITyGhZeLEF3/BZ4yTjJ8bDWEg/4hX+7
WCBi6O5b9VzVt9vEluiutFPWcVdgRjJWYFEc2pC+yVTPXoxgp4zj2FUmlyNXdZBB4NS5CH8cwFro
Nr9Cc9TcNf6u74IYJf5y4O8uV5YTDjJzl4guqdE1ZppjF59XDiYfyhL7JJJ6DdIzzp7A8rbtOb7M
cvdKc7gjN32RUWRWctgmhpeojOW9vtTabCnd9AZanE7gVWGDBc/Xp2gdluGoS3UNIuksnLSeT2Jo
cAvEhTTmIevDpuYbRqhu8GPFbJWSLn/r8+VQtmbiVvyIQS36Vtd8v+YjWq0GgQiKSduoxY9sWlxG
uK7TYeA7jONWyrUj2aLvk4FiZwPaKEcqMbMrC6x6r37ibfSIMu+uyak8rT82hQy1IZWhXZ3V6jTR
rSBGrg9Ym8/dE7XHFnU8FcyVmyW3UVWxwMcD9ObR3LCeJTWlWH4CBjITlAbfB74tBMqs25QTBHXh
zaZy0o6ofZzSCwirRuhTidI1eQKna3NdlvMMGnAzklbg3r+l/dHgE9pxaKBsEFdwAeHGL83jzeOi
b3Enb2SD1o0Q9n2lXplN24yuDkn5JDe/Dwmizp4yunhAALpL85JnGCadfVGIArmOC6KZN72/9MWJ
y7GOM2cneOexUtZPVxshhUKnh684/Pr4RPJFT/F6s1qmIAPFkgPNzgQEA3U7/OY3RrnH/cxT4JwM
SeggSy8UYZPRiJb+H/Pwufqt2OPNELU0qYDJ7rrlYWMUIy0n+QzTv8QClZaOiLU8tmpAgBG6NWdW
NfwdvCficUGBKkaNP0WWLrO5Okd0Isho24QRppdDX2FbCojc3bUZ5++0sofeD6VvJCkbcSd4YZP3
68kE6d5ANhD430hpo/XqAFcF3BporU0fTo5ks7NfVOQ8bBHHX/hduKIgVj+QzhbQiLzZswJUefpV
duwgMD03P5V7TQUC2/tvbf6ucIpa5nLejM/xHhrw27D1D/e8/03znELdUX+yxNOQX+SwZADaB4RF
bIFQ6+y/8h8Sb0U4jEPhfHMcaDpC+0eHDGdQq0gzz8lfh7JLke9e3lNp+gu2lpJV5a3J/Z7X5Wqz
cARudMxAUJtmsBnhSrKt4wQXnNWTuYN55/gQRei4V5iLzWIQ0JIz2A/xHeEOSBbMTCd9O2mJaUjh
K7XN0AV3eC4LzK9cWwL9iEMSfYfJQfckbVJOIc+PBelCKhpj7R2fbOTKgn2GQs3LHDD+jvWgh0vY
CEttNtNyCxVK3RQee/XQEOq57ci3gpoNAj3h4S3iWYRzoTM87nwP27dTI9W1bw8/D5868hdSbnk5
OqIj6ohNDSW3v0MRfeEeAHtPpa+tLA0zwO5MS0JQiY4Y+aFTO1ULT7WWodR4k+ms2IG+kiItaGCa
qiSPQ00k5GkPGK6w/l4iegCUrGR4ZmrD29vwc24TLfkEuo1UkUbFziz+2SDfWZ4BTo1O/uww2k12
/FkV6KfNQrvzn2Dk72zwEbhxMtn0EMVF/C8i1sjs2NoCzTSATBJcjgg7gTwjo1AASQWuB75zHXEx
cAB1zEaEh8IJ1tHYf908WsDbMNFyCrBNzwKTV2FctRO6Jqh3EmZsy4k7m0SjQam//zxw27SUibE9
RW5vGSTMW6cgtEz+CcCyiXK2eL+8vEgBT+/ky1qvAziwuTbZDs7vBEUbYH6K/K5TpstunSr+34z2
roLbfgHJQDBk6uXsNaXeKRihgMmwuW960SXO7AlD8bgG004clhyIbmyG/KPiqkkO1C8zGZ4ioPB9
haYsczMlFKHWtFGC8cnmhcYPavtspBa/JeABeeNphG8dygzGPgWaiRbUlN7mfn+RO4rUaTT7E1cl
wu1PfOqp2xq54ohHRuwvO1cK1yNhaC01sXoJwtNb2s2loOfLL2h0srF+OJit1zuxqROYz0JmR6Mt
VeKlB0XeQ4K8jkU3Oqim35EI/hW+MAmta5UbpILdldeYnSb74zNMXVI8DsweDAkDK7YnFJyYIwtu
nhOZqwasgYs6sZYLOU9WOaRiTP6LooR1qbop2zLnzbkTfaY027u3zoKevLp8wSuOSPEDl8yhicVb
cvwmM9+Ol05N/4hzpwl/5B7LYszz5Z9OdMgQ3bmFZ+LlLXqBpp+aEu+7fTCV7MwZ3Of3bHDaMMaE
Lfbqml01XATHbdXS3n768bW/6VfHDc3AwZ84Of1yYJvdh3VpR03g1fdGWwZI7FvlTgGayuA9cT8M
fvyliaubYsq9q1UTl7YDoBLhYW9oMHwEOO+e3ZOun5tapm3zPp+CD1b1gks/ukyy2m4AxNRKEmWy
qoeqN0tOTSIxVREndmoSw2iP9nzKLU3+psU6j0fxHt1Im/Ga4m03zvAGsLcATlJaVbX2o4ZobhAr
YmvMB569VYzHrLetVzNwUpuUvg7MOFqLEi366QRtxWJmULbAyDH6IgRRMf8ZHa0LqkpiMvf4FeCo
+W9w102KrpqPU/ymR9lJzKQgmFcKkvQ0Yacbv6aK816UoJT+PFp212Wij0cuX3gtIpPcvzvrGgdG
AJYeR5VgfwArFzin1CIawg9PDQy+2TPcKwUL3jUlTicNqjL94WmJt0C3guEZ0eFdZ5OgTT8qQFIO
QmD8VTb3JucrjMDQ7/fG3fVk+0CKNK0pX8IP3VoEaTKPdOgK1rkHfpUPkro1VbmydMkYO49xjZpV
fJpZs6+T33GIAa1d2MnQGgYWQC5c6QK1emrYdzeDbhRk/qCXbf3eP0mTWJ/0zz6mriBwLJWED+be
1Gm5y2cHbir/IoFMAcTQB6OrnH88MkJwsKzUMXyxf/OChEDwV3ApGowmN/EGq2IJtGI9YaZCswg+
G0tBwJXKsi/AIOYzZaOpPGFR5axpaS+Aclf3pJqGGiGTjipGqV0+qw9MUjNep3cPeQdzyfa5u7yi
KMMAXkmGU7ySpsW9QPuT0dkYnzbr8qlr2uGzd/VHBMXWpVwOI/fJ2+MeVUc5Z4mSISH8kZyoEnJW
n8/Fba3+mTbQFovIBbUOTjMgWOS97t+GCMt8JkYhgHGU3vUjTBOGUQFbXzA0O2qa/EX/d9SxyswC
7dCosIoaIk9vcjsuytsgxAf+ZmX05FstsJL6gi6GO227mbmlLS1kMnHEqX4HAfgyix1kGjvran7n
PiQulv1irBeNWTxbSd6MMR9l/RJHAae5wMXugbpVAmkr7UDU4Bx8Ag8mA/mqdFvhRuRTZ3Z9Qsfr
N5hcs4jdL9tCrkHBeoEp0BmaLu6ZTrUUcOkv5nop8C6a5N9NRw2E8IJgrumnC/FzSvY/qh0Z0KfG
SX8RvINv8QjlJGUhotkgM08/+okrkr2dnWPDHK0S0AaeTT7Gr7jppsagS/FSUbHegeZzBj9geYko
C+Yo3V/JlFxGE+k49g/ZqYzuNC+HiDL9vW/mGjA+xB7wyOEf13xlMqawRwtHi6xrTj4T7j2hfPqe
D7fOtmTYc1MxqMGGHSrCuIS8JrkAfA3yP3gdv/vi/ocZNa/xeOlr41kWyWrmDsGOGXf1JGBKxxGx
Kmw8KAzIdqx9UJvuzPC3HH4SSIuGqQ5sriXGdVMndUpO8taTTu+nfxy91bTXD7FNLeLPUKzlRGMj
nhQy38gFR4tCh7JhanSiSyxl9ThHTRVPkJPxWu5bvKygNjlHO0jDkZVPkqkpPvikgvPvfH1PLOTb
bDdfZ38FeEAqOCCAbZa7vYZzzNne+c7GgERdeeJYeEJUfCgAmJNLvlQeg49XQPKARfEzCNk+BYye
935AkGSd8zY7eM7mAyORg/jZKkzJvUoN+zNgi0R75ApgryFTAIPAXXdvrn1pycBEz3Fss1YY9mKJ
Wlx4rzdZVkNZvrVa+RHUVwv80bfnv5lsP+YCrkQ6k9Ehf2gVDD388F8RLYQqdjAv0o3Ff+RwXYlR
KyBYSezeEGWqhmqmlFHIt3BHGJKHBAx0+aroDU6+lsZLV4G4mWocR6rQYXZiU1SrnAC2xCyWX0CD
xauWkfCISNmOOpXmlchga9Yo56gedYMi11PimxZT4mWMeOrt26f/UX3J7KpxlS/U8ERDJRDeYSCk
1FEUM6MTM1mCeXWH0P0DYhed5xhbI3m80llRH6c+V2b3oQqMHxGG/8mEw/J1uVrIW6Yisf6ka5zz
HIjgab1VIy7eaUGNNK1iopB+9ne7a5BkANgxVbqMt46s55w5kE/uxhAz7bpeQH3qixv7HEH/utDu
ac869kjmGzlZFs7dap7rr8VhwnyCMjI/hNeISHlRdYP866PgzDvp8/XIu+HAggDi9M+vvzmHfp9h
u8Na+RRgGsawz6HFVy0PtDmLfp9C6ZLp2bnBDh3A/NN7sE9gOaJQovi6DyGdWGLokSFGv7sO8wQ6
h2ESeaTDpdGc7kgBD3GR3vqP67ty6IDQ5+15bIlnVJ5WzoWs9uEw7ukj10JJw2AhPCr6QC1UXkQl
HIDKxFwuHSpWz53Ciu9gHTeiZNFsxUFmF15iAfbKf9FNbuJWkk4ANNSzBx+s+R13+vjBPjIvl2kq
wvWwW+xNHKD1QQqPas3b+60OfMckB+KHU/2Ncn3ox6ss42j3IG8A6RRID/+6CH0BgnZoxeioD1rM
Pm81eA/z+3pKDHR3eF0UYnrjWr3wC/Pzc5/AWVU1KEPoitvQZXTr89uc6BkgwxjK0G2ZdDY44P3p
p9SJqiVl8xkhhr5vTQ4Z+a2ApZQZrTk9bq0yhMLXS5M3Ho4Xd8I77f4ncUBlhH+Ror1QGeKOWKgq
a/OS2WhNdyQsmYN3CBLvs9OLw3HI7IHYOI7CpiqcXjbfWoY4dFnN42EDAnxfjAPn4EBpVT9RuZ57
b+KdSs3OGRTHHDR2KV3N2Xt7L0Is4XiKIzeARiQs5qeRx/Uox70FWUEmX1iGJUo0Kl9NGv+n7fjD
S+0/sblm+g1plHJdIRiiJXqRSkI+F16n65o+p9fPgjYE68AmZJ4+BH6y9/EyEIS+1v16TepELBmR
NzziNVjHn9RWBRBACkbh/UOK67YgXkoqveKtFDn3F2sXeiHKATtwSEIqkSfaW1sAk42h6T9mA/Ma
NymwIg+N6G5H8N+9i55UMIdsYB6NDsu4Z+3Q5ls/Pi6hFAQKJwysfBmAuoHgJQv3EjiY8oPB+JUF
yIcYwhaMWxXIPqLxLcFb92MnnB1o8FEIaLYudCC54ZOfs24UoWwAX/7chNwsAEtYm1odH28pLbQb
NguazEyRn9nWDx0S3XIoOx10C6SkvjHOruzPbGEULNkqmIYId2A3VlLn3VY2zU7UfAV8EKACHGJY
s6simjsygU8qVrgwcIj/0nMMbObbpPfXYvN4cZ4jyhnfQLxyWHd16GFt2eZ+oths3brDZyPm6eh+
chX5cUDQrg+OV+HtG6fUMGm7tuQw6sFIOt67tHhGkaDR8W2dOCVtvWwpShNLXjqgfMUdq3Rni68X
aeb6XvR8p+vB+79+IsrveA+tROzPSV1jcSwP6Hm3/o/NeOPJ1bhRy/JzTCIJRcbxNA9eb1w9Xf/J
yqdZ2rYwboS7j22Cf1wC/EUjRFufkXT3KMhDKgGtfF8SWJtIt/5OmKZ/FFIJVlNsfgUiSXjwDT91
rp6iJEh+3K2SkOuq4AlLIU5fyu7Y/+XjUQNfioCzG/ZkVCn+w/7QKeBiXHdzynhQ37n0PEz5LcGC
0rEUdawpxWYM7GtAt9891FAB+HX7ys9VGyZWvax2RStXartmuZpdviaC7n4495/lQ+jf9/9bKTok
OGSCAiTrBYwPxOZIVcgJZSmIgUwNni/8eXUeOtKyikHliUd18qTtZRoUlPPlef27KlXpM4e5mBiO
LKX55SwJ6N5JEeZSAtNdUPAE3K323o0bEJXGJPzrCFHAjf2NmvpDmUmkeWUxwvuF45eGXpa2pwpc
LZ5O4L3hZ+RE7IguA9FGglD3/P6lNh38fkM4wVnaas3MK+ORHZBQguD7bRm7vbr9Oto0EeHSxuFx
YB3WiqUl6TH+nzG/nDx1JiH4P475ey3ZZL4qSHiXRsMG33rsHeiWuHrak1RlzNeMgwAU7UUBlHq7
qMjjUpVMbfoPfVkWVA+zmO4cYgIbyycGClJhyy8P8u4CQvOvKsHY77AYKM98O3w8a7ZqmV+Ob21t
7lcZpUNq79igV66vKy7EPJ3SD5TIm79vuLcEEvfPHNeC/49t7tM616hQhj8Cajp1S+poIIP9BrIz
ntM8OepgnDqPnSqzSui8YjwK4lSUFpl+MhVr9AmIQLB99vUedMR+wQRyw2DJUXAKdYaQUURZ0HjX
RFpvaZWFQrPZLn1MlziRIBi63lXa8WF/Lu7BEQObZngY4/ACB8N4C1l/SPkC0LhCQe+Ts/ixJC+M
7Q7ffrztZuh4icfTXqV93c//CBKtDMe1zfVoEz/+lzgqsr5Wb8xhG/te+a7znr71oJrejtLGFU4p
sTEHtqOuFTHjLkq5zpQfW/hJM1qqmon56E6cvvuvy+kw547+TPk2vXCnnNn4dmcRvGr2Bo4hwR6O
ks/DB3jzDzXQQn27poRUKkKI2wrgquUac2eglrSY0q7Ep/IhZU1tlADDzZ83otZiGRmYKwSBh4+F
hk3PwyUofK3GSMbBAYylq7EQdMhW1QLSQAmBeYho/O4R0UCW5+UZxHBEte6CSKXlv213PDGGHqo0
QPt3JZnlS+qk54cALdUDWPVYjiKF1zmw4LFzll1YiYPW7TrdaxaJb9WL011phhxSQ2sRJCOuDgmI
R5uUr5TfhEHiqOf34LOGe+3E1urGOyX8Hp5oJw+AuZbcLuZbOUY83H/heyYaju5hgPG5k5F8/IoO
XvJtObI+JDrb4NsCIVzieORfF7MUslSbw4JD7CCaAGvWamuYBu7ZF/hn6o7/66qlGNPRq1tMzggi
FvBhwhedf1FpCamDYMTfafqVFSDtYxRPjJAGbs8KwSNqrNtwkPzGNU8WxwCEw/Q9GxBIpRkd8obd
SRomxqfF5fDX3nY5/oABFQphZpXXpEWNvZ8o4fyvxK0gq6EgdVK6nZmm4p9W1t2YwEulEbZ/g5ps
zfqRyohLtW04P8q1+mIgvl8wKbxyJ0unx2ry06FcLLDQkjZye1Oi7I5IFjnmY1Gqto++Zu8v+Jp5
/mq20sJ+0DMLSPvuw/ajzHI8E4kDr1urz8NqtpN362/jF2wGeuupzLzyxziHq9Yrxv4a5G84kn1s
eL+4bncwsX5rvPLv+D3kSy8IwDElsxEnX5KsPuFimLThikI+3OctJnoT+kjofKhEJEUFpKR0IImV
x2TNKK4z7+TM28DMhXSApL0IbNgJ/JVQbrXaGhaQUiNrWK0WQe1JGt9Vp7KCxgnaaAGL8ISu7BYJ
qDUxh7vUBakCat9lgOlh7rmurtjO+cP5jUvuGe70AUG3ZaBH2usee0pH6SZ3hYHTgQXXMSk6+ay3
UYN4QVswJitdUO/lDre9PVdgp5tT3lfTV5KcjDqi4mA46BvOaeoh4UkQHIB7vlrfn73ytbjYnYmG
/EE/KPgD2ORKlY2zkJrZwY+JA7VtMB+PYnbQN7spYEgF9l+1xVVnldokh10BIfiYLE9G+vNEdwyz
RtVX06V5HKnKUkXU+nubLF4ZuWq7f5kElV8XpzE1ZlG6v2UcG97IEKMKGz/Dy06910ZG5pxwDz25
Q/TTltRQ0FGteVhh2gPb6Ep93DA5jLGFM2E8DQl/Eu9NvpHSWhPwPFISwzdunl/FyXRbJxvDpv68
9aNfCwN/55zPtjANdMecxpzzvNpYuw72D9cbvq4bzEYTG4hgIqQFEfFRc1whQzT1ZKAYbhr5vRpl
xbndu88H8J25vUw+5ie0Au3SkV7BtugzCuA6MgaVnrwiPLorn1XxVRRymxTqDbR+tdlO/KOdYbgF
xLd5r3VHDxBCT2vPVvvrV1pn1O9bhIA8TJw7S+/Dosf/+DcY5MI2EQ53d5x5xYTUOxEBTv45XgJf
E9NHVHyXOIIUjre1sxJMnCk/kAGz3SLO0RP89ZWdcRoxE7zgYY0CbuGTpYMOSv3e0/jV3kHR/+6l
Pe//vc+JRhKRh67mjT2l7Y0PWMg7GZ31ZI9beUM/NIm15i3SV4+AyISBSH4gOb2HfYbFj1NlIsMS
K/C4fW/EbQQw8/EecS6pIAij+QOtikdASSVs18br8pMTQgMtiVpHbnRsmlmuRn6fOhUaz5Cg+QN/
x9MAOLfRNeAsSRgS2CU8rFQm5CjPpR0h8sQJBv+7xMMHumK5XoHiv4UeFKgw15qzP43x168xuLPf
K8+dzqXMtgeA1PtSKsWeaIxafvOMlIo8sKTsSF87P+L9Pe3rdoWdtE6vk4cBVQovPHjvgCWbXHug
JfBWOv0f7aJqmBAVSFusBPCwwwU9oY/bbhdRNqDMmW/INSU2/9+o5Kcg8Sbi/36XkC7Rwo6yEcNX
n83r4CVuFlg59GCBMFn2b7Ugs9vUak7UF3Allaa2i6TTZLkICULXWezf5pufbLgbIZJaGb3zeB6D
kJ0PDXSAird2du1q2OkWFmsqNxA68DsgfYEajPleYOffDgthckQCmr/yDpE2iMhCHPAjtXxy5BZt
D0ZlT+fs7G3wBG7MKXJA3NdKCH7qEZpZvH0xggWWeYqjJM9TqRoULODW47N4nDbuHwjGHsqZ2vy6
io1u3DA3DKPqTKhUKO9ptgt21rFpYoCxbm3BLNwQAfCT2hdko0zwv6mDYfVAK6s+zJWf/DmWtSRP
wbvhARuRpNjN2aFlfqWaVzaAoye83OI1UvLaoVeSJfHLF9XEBTowi5dYP3LR/hIpOkeyGnKG5r6/
UZnBwjI2p6d/BHWu2rJxr6YX/Hrc3lQoikIKZ59msfJfQANN6RtkhqmsZb10gVtnWy03PvmNsQDm
ZBQ5v7wNcg1wf8SulVEcFoeL3xF0CpH7+nCwXnz3K2YPDji9sieFBYTdHg1g1loTOc/0HMh46sSV
+Cy6mBGgmdLmwif+d11k3j6XR+ECKTmLibJGco+Vz5vPXLc8EgSQhb088VlHdC2ZU3M6SlHhrvEt
OviC1ZMpGRQ8QJOTwlgSGQiSKipJeggpVFm12qjNJWQLywXrtJHxZlKMOMAAI0dsOilbyr6tOREm
DDhjVQgUGg0uyFJMvd2UrQZO4z4SMX4dMaYR/EBfIAjlMzbJrSxJV8gYraWsefGTADCbwaeTfLHT
LNnu+pdAxM6/HWLED1MTQMWq62JOgDrfK02uzFiOKNsB9dAK6I/fjYmPc5qolP5esO4f0GmCvQuq
AhlkVB8Re0xt/UHfT/09W/MkAtH8uA5daSo5VSQZmT1XuHZ1nxfolBSGguwlyiV5opDWO0Aaa4/4
G2w9CY+YIIWDESuHlkxxMLYNG/5KFWc5rE381Qy7AozK1oQ0o39ZMdyGAPi3ZxiCZBZEadmhixji
HUnYaXSGg/MOf8dhoRscaw/BEfWsrb8BhU1tuF/RPg2Vs9O6mxMHygO+5KAcGgkwFWmic34Gs3xG
AgwMH9e4TONzB/K01LKAA6d7+ZyfvhRrOKqu6n1XVfqsEO3/pn2YGGjv3YCzjC/KUbDtqWOsGdcN
EpsuYVHQnVN5lK/GieLHdMdOw1kO42WbOPQww6iabr7tcuVJgvdS4tzLAfcUma9z74xX4vTQVtvk
3EqAYVRypQg2MOeENz7ZX2rxpJlTHOA3wyrXIp81m6NQZBI/kGU9/6tZp5SX+WI/EjplRroaoQH8
uIFAaaOv7vSyj45fNXy5EXxR5A+U3euOPjJQYyfSSGcNFez4oojKxOU6MgePMtpPdZyojceW7e2v
MQxDY+2DGt1JhUNYcXHYX/sRLEVOd9llX5gDUSeLsp+ROlhDqlt/7Vtsv5cWZAyQqUnIpMvnPcB5
BDhN0/eM8QMvTMjprz9Q/R4EOElk3Z/g97rEOD89hNKA4EdX8xwDRguJHKod5pagKygNI79dzE5X
SB2gf83x/jV9mGYeKkrmdg+edd3EfL/CTGWkXmMNS53MBBtDlOZu+x5p9b03LMtkYN82WzR9ziwt
C4cYr1OOLHnpos0RX/g9WBQCOpZVM7SYo9IQgZziNUN4Qlt8zfVmIdQ5QPPyczegXk9K5hu9fTAi
GHmQ8FUMFrwNl2GtJflrKRQ04kSeJQRnYLSg+CNrr7TnmymSFM+bNBv0Y2/CmcRzlf7/eAhpzJgz
/kewthfBVi0amloqlh8cS2gQr8bO3+QyvsEADjRUoHf2q6S/K0Jy4lrQTa2BPmjntxb6LPtlAGyp
U/LOjLZCxcK7/UN4klfRSFhKHBBQiTacKp2qJUrwFJMHQxdv0lHa1ByWdwI4kdwNhy+nzmy/eH8V
AFhQhfUDA/ay0Q9XIDEStx68yp04ADAF8DFxK2tntn3BI9BhEAe4vhXqqt5+zRiwChzF63o/fTFJ
Ws1nIQhENWCQ7VPQE6+46YX6c3V4HU0FpCUoADtyqhzNWrc4oaD1s2SyLKpnaCm33W7RBVs5YPnJ
FP/03Xd0HaWGQ1/MBNm1/bYOSqkC/KCXw2DF4bBvG6v2ucYUdXnc2B8RNpkdBVQgRBfauDRQDj3E
E4OKh7P3rT0Aoma7gIPlud33WUmJYg73551XKeev7tiiT9I3PxODiUHjhteyAiHxOogqUDHqMVB8
/yF/619kEoSQVbumHNdUcmj7nEfNc66xVbMpFPX0KhqWXb+b8TGRkZm3bDLdO5aR2sByJRw7To2+
i74EftMmEgxhMmKp6qxoWW5AsmLZOpQp4nRroQCuT7w6Ndx2/z4LdtAKgLd8DGpcgIDUWziZX9f8
aJYK552gr28c/qZ9ZqO65nOojr7XTcMM5CwIkXKbg2eTRAgQeqkaNbkRj0WSulZK9wg7CVqj9evb
56lSU3RpcW3ePN3RbJdlfxKwfAYTqDTjni02y4NUK8nMwwbaUllToIJQPlO5zBjpaYlvY7EgDmHi
40RuSrrBEywwrXJqLitOeO93cCMD9NtBOGtO1cmRydbZLqcbK06s7HnOWTW1dDElUJ7hc5A2oxfj
iFctSPLNFQlV9PAZFshS6mRFtWIWwy5WaAY4KtGs2tcdXK+6C469cl944BioHiaUNk0uMCEVKJFJ
KmkzjVJmMxOt176r/cs+F1qsEYX5aLdJE4+rHFwHUB+BIvlE+jHHCdj4HC249i/mUko+yvLbiIQG
PafrFvJqBEytr3lpqOrxLkGo0Y32sYGzR/2ARCI6WI/hvuahxSEF8lLf8/DklYrjLEzZ69xrMD5I
1ykkm2KeOkV51R2mFSO1NyQBh/vRvt4GBi/Z8AnQbbZC0ddVysqRgrmNW5DocCC48usvvzQHrTOL
NweCxinfJtWaZAI3n+aCtwGdqoIs+06tvZ7Bt6prtvzv/WZwlQoV2ezCvaf9KEWvUdZJsbr3bX+F
p8bBWxXB9XEMK6S2bJEG+w/6dSljjN3aQP/g5TTvs37EMg+SIP+szZGTDiGyjARqdR7sWbkd013a
4jPbvK4nPYbS0dKJCVsAVpNHqdBazRwBu5aoiQX3BS6EsxudUPPPSF0TDEf5jhbq38TLO+11UZrm
gS8H98q2SDZrDBso5AkWXKz05nFDWruM1IDgcJJLQKUGfXqLX5gF0ZzAOY9kS66ShKUiYLJwRJss
GvuwJGN/OSAiHAlmb898TJSoazaAn3jefDljjktMaWPXh3R2rbUGPo+ol48Dl8xHLfndXLSkyjOP
NXj0yO52YjZIcQxgn/z7B2IdQf96QydD56bGUM+aF55WpZjHoeCYnDecxyf+muOvKIWfCa6959XH
ysF2FetaBShWp0lU2QjSau1mnFbT/YBc5JpAJ1CYdw/5HS0K9MoRZ6d748dzi0gx5ekJ8IsyHerF
hw8kbTkq0GHZrZSE8CGGKkz9EyNkh26Tak1+/oR6hDCmj+uAkNlsks1rwE02qunkOwhxbqQPazKn
Nie9tXJLKfFkRVRrruiZ1dHG7hWdyv8P0gQWaT/3Yw97GYbruCGr+MwB7Zz8DlUMeyaVrX7VZU0B
nNa/PZ+5dYdbuKT0ghkS5EBL1mB+HKaB60sEPhHBxUEi576aqsKnS9o2Vp7w5BegEkh1/Ox7Yq+I
lYksNo4zv8e0ER+0WE+3RrLexERLxNnWF92YKNfOXmsWH3hbmiEM6XQbmNvBLXE1nWvhwgqfg0q7
NbufSVoewYNvjT8k4QUQYXNZbW6dB09X2CRkuyUNgTj7PNMFcvVr0VSMYoPCa7eDh+q977hcv9Ob
0ftTErRFnHzA18Tc62k5YOwaZXkpSH7GKogvxnGqc0qmlX6dvYkUqHtm7ctPNE+rtNyYBImtsIJS
ikNzUlOmJIhoOgZvdc4VSpB+bHtWX+Ezp7VytXLXXfH1KQkU2XDbd0T3h7hDSe6WMUJuOoA76iVx
RVc0ZA2JLOZELsl51lsux9VKp/Qbci8ULRDL/GBPF4/qCPF5vaY+nf2vmQFnpJ62QwSUxVzsYw64
yMfecqpoiU+vcSPvmTqDPLcvi3oW5/DhhDtJSjJ3ZVNf3WYO3NB2QgqnmaD6j+sJLukAdgMjX/4b
DEp7HaM2dxznAthf5xn1iZa+XTgVh6jY/8mAQCvhtZuuhn7Vjrxq3JdmZKTCXGbEZeshWwIBqGeo
qagbsFr+Rpv7KBqzvVv8dt6sPVk6hwzTAxv/UISFnsLSQ+ljvTc231UozWhjlZE8j1XqituIAjLc
k5UY30FKMunw7WVsc+6Z1HaOrVKFcdfY4XtckTnzXC/pTNpzEPO1nPIVibEgWYoBtYnunVD6MhB7
w/F8tf0eGjhpzH8nLjKcm3GeIm3ejB4b7KnGLWyaWOEsR7bS8UIovCVv3AggO7MCEktP1G9kmN2l
29WGvMTBu2DenHHQU+pRMvm14C/IxR5gWDRfuHAXh6SF6zqQGTNc4HjSJ63HA8QOwSyuTTBXABZi
m/n2haopGjPQOQPYal/nzPv6ixNLeKF4kkL/MJT3klyChmtdajQJqbTH9H7JYio5RqGXOl/oawp6
d9l0Yp2lZw4rK+TzocU9vfolmJQQ7hFix3NgBYV5WaVhWph7vRvn1yGpJFKJC7V9jm4yG77AnfLs
+yw01IJ6mprN220y7JiL0K6hr4fCSbL/i9kUhzI99LeZYq4vCkBY5qyjVzXa5z7TtWbvdQgBS74z
LL8xNjSs9vQIuBMHsGok0jCX/gyWSM21rahgfmfTDnx0+fIgP4V8fcG7JAMIw3JAdUnWYEAulIAZ
nTEiuMfIBRWqUxCMiSxVCva5os9am82dqpWq7+1zrwO6ffEX0IP66GfpCyhfSomP7VwYDDOmNd6E
omnBMvTnrzuNUfbNbAmouC9xkarXo8l27TdwzF208+PtLO/whKhbr3T3kJ4pOIHibFbJvHA8K0Yu
/rYCE1Ia6c5ylAOLNwAggA5OECRZRgmHD5ek17eB4N2RlRaELpV7c98G/KmOUkp5+6gOpGz383XI
u3i3wajwaK1PzNB1dUbjBnE8RMFh44Ird+Y2hk/tlJZuVO8jTpCnIM9YTJBcF8w9f5FZYNd7l6ze
efqqjziBpeLcC9NmQAD1Ummp7Fmo+y9+P2i+nVorpslw4cIOS9yak9Tk5MYfrcz4peyIYuwuRwai
H3V1L/Asp7x6RUV2xRmB+hhCp8lavorTRBK/RgVqB/5aVyygzG/DPwAzNub2pN0G198jIqvGCax+
5KTJTq1syIl94B4e9dFjPNSqFvVAQARCIdF90VRWujpV4ipHhXi0BcYky4XQ5JjKaxgp9s1NWx8D
CFv80Sjh6N3KmvS6oCMfn/JYjR4oPa2CQ7J/t4IiekalxO8UlzfXPmiRkamHMx2p1JglVDDXCOF8
cBne5S9GPCP/MMISZIV9l7URBjzl2hQjnD6ckuA7BYwbx/AQS443h1bLpEc7yIQoVde7/5YrYLof
D0rGmMLUioUNywFef7VOjC4ASxzwIbqOtsv1lVTt5VMJR+hhrQoJMMp3uF7qC1Pb+ECfm/iCKR22
gHV172X0F4i6WOy4w2uxm8FO2CHm2ol/9+0nZIqnKqA+dvp+XLUincx22jox1RrZUczj8TgeDL7T
aEFT8xGYdn2fZgfJRWYtNd6dAEprMqAPXdE8vxalRoakh85cXDEOQ+SFXZcvpWmMdcAg0L5g6En8
RmSXzDkj/wmv24lcA+pPrygCMatqeeKfHvyDnBVB4aAfa/W0dmoDk1Sv4/4UT5a+Krjoi4laYzGe
2IPOlLbuvY7Wg4taaHYfEhM3zlaIMfK7sj11D5ukcD1H1eoz5xheTUl9KjX+Gu1vo/OyOUU4J8kM
o97w6od2quqOPpb8gjTLOClg0zWGDayoLSmZGOAiQLp2fjW74v6uzBUjY/pwIirWfNJ0IHBMjD+t
5HKuOpSJGG/biv4oGYdpF6SeHIz14OlYuYsm5d/jVBCbpF0kHTc3RWy+9YhILcfHafGtfFxVC3W1
k4/gQ9CtPpqmBlcoHVKUFV7c44o8BxAb/sybjOyS9u/EDd94ef0MMUqTebkLEHURsVHgOCI4U1R9
4EbXx0qo3F+hRcYcMct7Qqvf16VDGjXGL/HxUzYmRWnFkf8FV0WAOokXaZRABjoKcg6Q3HDGksnZ
BWZdJjScMU9cskp5Ee4aQSCtwTEgAhrv0RkRYrmpl4BKmucMWgiH4Goac9KoaPKVgCvz/XeWzDRY
Ruz3Sthsy4YbNX5iXXdv1bSBzoP39E91hmt2V8M2D3w9FHpLcpupK3LaymxIVolZLW2It4sqkLlP
6VK0r6C7BhbiOUnRVGkZc5oGaOYtBuKnPvst7Dp9HywqRCDQZ7fFnNz1atqBxcWbXglpSwRsa5F+
PLYOvSlJHXsEBFmvhT6CN/Zs8SXmodTR7ZVJIxJzfdfenMPCM/L7oLb8AmwoUBQs7agq0PegUdRf
1ceCCurA75znwbNvQRzTxao4NrS4O2ciWQlTtxU+s8wi+JD5PCiHhGMjl8nhcNbtLT7NQ5tdtU7l
kOSMfzC6m8TN//uGqIvIr93swClnm3Ffrkq/AOG2RLqAIQl/r1VGZnHDoJBPIuZJB5rKMyN0Fowh
Dar96g+Whk06GPbjv2mS4R6fvDhSkXjo2nFBdjeZbNwsa2wiJ7YxGcgjNi9hzk/xgw3tkH5Ns0Ud
FfFPzZO94Pg5p+uAq5lHBEc20UDeWjs5qQafyxgZMfqZqxWMcTWUbbKlEmV3gqd+zHChABKX4FDN
2WySgmTS8sUHnNtbzc1ceE3Dr5O7fn2upi6gCUQ6FAfhcWPQZi9je/yvUb3Up9t046YTH+EAu99g
9dMy6wjnVVtyqaD10nhrS8xRqkRfrwoJF6uVJqEQkKFxOkgeGFGtxA7avLTtT+ah2b4IMU+yg/b8
WCW7Xh7innbVapufm78grQwG06P4KeJCjvEMzkwHDmI0wBhB0iz+yVAr8MSxeWouEdes+eMeTnbR
AQ/lh1loNinSCuXzp4Jfg8AzGNkpDDi+YbPhEBzGZNm46c+kWzHN+C1mU/Vv4hWB+A6yGhz0XoAX
zVYRanGGxIl/D5Nt3lUbGOjgrqcD+U0ZOKtHt28me7LCdGq4XJkkrO6GcjXKEGjkG1Bi0c5bPEY0
EqS8GoBAeDeENaYdSNvEUAllFhgHurxm5n6ePbcR2JGUULPFeyyElvljkq/oL4yqYxjlDYbvDsK5
eKaEIdwIahDSVvl+quKGrnkMrkDQWyHM2cLcXKZTXjQzkhsFirPY6FHsacSIjGWa4PRlLTgZmvDA
o2iA7KZ1bikKAj2piB1Y9lDc2+1TpN8e1U6hpHX7c1Z/HSlK2xH53l+9nsZyJwW5XZVYcstzPRmg
lJYWeD1ISAlpRpeWMsie55C99dGDAEPGopYxTxEOSSoS1wBhcrfqtycLMLFqzq8UkwNfG61u5Nff
Bs6zEh1oBzTvZQ0AoXbFq9AMvTib6leL+8czeVtiISZnxnIsHt8EFWpjLLnMYJxreqAKHTDycHK+
hf/h2zS2VEk9vr0h4wn2t8ov7mxr34onjr42jjBrt8B10w1py7EQv73QySdchdU0uocTf6e89cgU
qDHCARI8sTqcsAAkOuzHYVLWxt0PsrMdhmzmfWIJHF1xioCRYomL0gitPhxB+7au3GV8rgcEkOsu
GT87KD+1UIki/HQ3Ve9G1ZfnwkM0SqDQfiKL8l9Ci+7hsgARXlI8QyvvAMGMH5StnMHfJJ2jt5JL
Curka4suJme2lOoy9k5UnpWHFUWOmjWUx6zly5nfbxYcG99enRTpuNPn3Qk2xX77HYiDmNOmsfeK
psVg4xNxELSkcYdxSa2LTKn7Wxb2UQZ+v/wqGCau8ZmhDP8UjTSIVlBHJC3dXAOVDXGj2l//IvP+
KSjEKiIG5QWWsfOzTwf0jfl4BfssP/DSkBVom2Giyozl4n73tbrgvpjGBGk3v4Oy7zRaRqiYdUHI
NJGrlDZOUGP/VOy/EpuekQUxZ70BdZzq0kRcsnenoYtbyIJZ/NpT5ycJmoUnFdEP18UzyidQG4uV
PqDCFgfSIwmikAj5ICayfwnnBsC6QfvBst89qysnFGQq/VaH+txLWsGOw7KftBy2ElP54MQFESHS
jNgx0yP4UHGRIyz8icBox4fUYZ5W5pmvfoHSJKsapXnN7yS1+wlRyj5Codn+4bv5o0MxqPdLdZNF
8CKemSzI0QnCLJ40WdN+KnEoACisWFUVOCKZV6Ul4YkhIjtiNRjjN63cGqFS7GkHxkq6dGSmbIcK
A5BWY/aPSTltW59eBjqYk8be/IYJnbB2lVFwmTKz6A4HV7siPbie4FRqbQ7iOm45MzBMgutjUSoZ
irAsRsQfGAamgYDJfi9MWzntYbwtmrj2PE+cgfPpz6yxS6rQpUu2IG13sG2v8ZXm/Lub8OkWJ/Kt
qTLhf1kXbFCkPlowI3ARXQofN4KVUpSLoERCi1s7U/SurlArScoV0uGH24H8LU1ezi3AR8gQPWuo
ykWdgwLnmMCDFG3zc+PBpkaxHsI6m07bwHvcqT9M2i56zld4PDr/2LwqKcLcfxhFB3uJ7tZjt4EJ
WpzGaTbkTX7mWszo5ZIXnojejEvqeUZV3P5sds/imiA5wu7Nrd5AV7omdhaall68M692iFJYcKrw
AgxFRpbH8Hx6xFkQWXYjkWtfGthAQZaNsRshrtKHz/rLcoJqGoL6bZtIINySBdfb9fNu9Z/UOFLR
b3TSTmLm6E1efVCqgKskCOVzMvmF+fyGCpR2cBQxbjQCPcfQsLo850nBhBGsC+mePQbSVfnJYbj/
Lxi6n2HRhY65IlDA4r5dzBX5rwm+rAHfhNHQS8Wj3GlQmX8+bAnGD8FJlSQwGOKrUwgyH+9QJQ3E
p3hZZxhQjqmgNo6slCp5lQEOEIzNg0TpPvqiboCqwFBfGWxk7Zxl9dFlZL0JjYpu6sZg4n7G48Jn
5eyUtQ/27SuNskf5/7aSeEUhQxwdKqGdzBb6QShcbLWHomWKBjBoqIcejmdqpBvuBgsT5X1b0QKg
5WTVmm2oLDya6aAt+vq8R2CJjvVmumvozV7630EzfO7BGGpqeaFWNh6Sz9N8MWY9b/wrv6t4tk4d
bCDNbEEb5uyXIPGTfngZpV+v3DGCs/eb09c1e4cVH8FtiitzlmEXx2uEqe+xZLT/zSsnfgbVnA91
GIQfKOfcpuaJkMjHDAeJeFJ2EHY/V6Gwg7XtL33H+eeuaR8Io04gcmMIEKB96llOpGAMsuMVmUFA
VNawBacQzGrS439Nj1EMcin8enfo55iQdIYEwq64TwmxOscTm1gSxZyOzXHTjrX1gy6EOfkpkpEb
sLIh0BI6aCIOuzFTFRcUrOvsbSAu1ElZ6PlKqQ6bXC1L9aN3JLlNkOhsmypWp48TwIkLXskl+27Q
+Ebx6qmfnUT93HaEXc49krrm36s4vgz+4a/1PejJH0FIbE8BbL/KtZKah2Oy/DUZCE6pyeQI4Qmj
bhEPdX0K7Tc6PKdc9KJi+8jkhxT4Jc4PS0HXIbh9rmdvKI08BfEBHMIaS6LP98m5doQksM9bpzNe
R8i1DKh7plarmLYgVEyTzQ8AyNntIrRjwZg0A50HWWzFroTx8R+QCY/Dj6TyplqOqDdo+CzGNMvm
TNsGOfPP7TSVGoO+U9371/uF/9xTTF/yDwQx4jTUlfrJJYd3B5dDPPvTOCNffPj1cXCck863ODR9
+0giME1o6aMqssdfzc/2UuqELyqGifXcjhqgZLGk2MNQR9P5IQXvSsR+MOBPWQaR6G7PBShhIE3u
l2glTo3fY7eUFj9ouju1yDNkT7yeFNGXBCO+PQ5072ft43SBSzb8ccIkD0zQ+NY7VYofqypS1Kl3
Sq7h+POqaGLul0G6SlcY6b+D0NF/9HwYjUWiGMtwOkhqrDxdWu6ghvSSH4oCFxgLLU2J3an6UsLV
PpnQRkzNed2vqcD87m+yQXoxSD5pssOvQd5l2LIBWSneHcskWBeGSJ09s2gQT4BCyfUQjA3HpqId
gLEt6UZ+WmYyZiH/OJg3j/a+hJf7iNmWOK6xIhY9G2YPkaapSQ0H+/Ivpkw5UJOPq4dh4gWyE3BB
6I8nXC2ljuKXQYrjHspyZYp0q59GvEcS16I9gf9dY66a5dfF3lgVtRbMffqvcM8X847qDCxMLM0i
6s5VPFYXOrEQzf4PF51i3+BrMxJ/qb+JMCbb1+o/dfNqStDfWOH0YXI8hnutEcW9V1AL75lr5IEE
sukYICML6D1Sfd58osXXYQ4VFW5e9UnjZmZpHk0DqBYfCGFRDZq1V2sf0bSuC3axF+zuG81yxmDm
uiatdP42tiQO6vhqQjk5CqFiHskP3W1ZpBpWEkWGMxdE1mRd0x9Sb852IzXOVda+O1HjOwWZvE7t
b6YN01zFTcMNRXPwo1VQ11qtap5/9gyqf4qMoZzexYAJE/6/cVRE/H1YelISLIFtuHK50bW0bfqe
80/tPLaZFy625t/2mmxxH1n3X11ng7I7VBU9I+XWGIUeeWc4SW6v10jZNTq1ne3LzxVSO0xpBMm3
CwwBELh0H3YTVoq+jROtmdH4LYTZcvoshIaKM52pw2KepSVBaSkNjb2III3dBX2ypzKzC+S23gAI
lwzQFtlygEKX3qz50A4jJV3GzBOBn4mc2H7buHe+Jchy8+mUwpnOTYtblCIr4WGjSz5K8EYkqn7U
XdE5BdO2ydbM3kc7cSnuZCk810IL1E+E7XZyKY0uHHb6sMRmwjHYZERecHeprFblMgYDew5cyv5n
5wcDagxUW6ZMGskPfVbjTTklOKBWR68JnFdrBNs/ii+3TeH/j0sa9wlx8ZVBys3gSE6vPT60WACO
NSHGyCLcdzHaHYNcdtsly8I3Py6GhFsFUNd6QEwI/MgPvHbXU2DXPIbBdqM0q7AIAgcgRyCrHIn7
YXIWKYkz0vDMbVbwqISa4ZoPnpP5zJORO2ANZnon3R4slsar/FrTTyypRHeRfdel4SHw/Uwy2D55
I/5WaZRfygsnBlgsowWqe0/OymmKMje++tNi8fcoRRPz7VeVxhYYbnC9+5KjX5Aq95ctGPkjpbwk
qSKvpU+ppD8xGjcsfmXRnZuUm2f1aC+hxTNXOGZmqUm5OVtRUC52cJCGXN3/yKeXQJo5x/iSotuq
A8VRrhfwtr9j6S8/g2EE7LFhhZ/agkKXSkuQjVGYkvYJR/iWJqrNr1UU/1SG5bOjTK8iWiRwRU6X
HfJG1LZmn9EVVsVNPAzdVUU+odktyIbUS/1Eg17lLgQ1seIW2Xhydsu7yn0uaNEeyzqBTidQc6jO
MWsIbIilhze3Yn/0tSHpwGQs8ZlJgIaojq1jvjIFSdAR/LdlMD/cmSEcxtU20gBKJ4avQDW7sMwy
e+6wB8+KExyTxWr8Qhk/Ch1GV8MiephGvL/Jp2MHliTQbEvhhD4twhtBtEh9QqsU09Fy9XmzaeS8
+yohUzzKkNFXzaY4+upUTrS+0VWIgy5KrcOHUUWy0EXcUetr59j8MDOcAVSmM/FyntAVeulEkHog
LOI7jplSWZcjh7BlNzOXWsRP29A63QwnFpznRaefzrMdR+YaP+Bsez92WDBe/RLu+jdULwzx2ZjF
hkVrOK+xHSmoPhgsQ0VDPOboMxPtWdwgdNFb5tVGBA3w7+d5KwNsDuysf8iYjM23A4/NEwm9jHH2
Lt2hjq3ynS7ZimVrxdtL4Kqij9ZEKqmFnlR8P4uDkuL17ocL43X0WN+HD9hhnOJX6Sjfb4HyvITv
ELsnc/aVteP/DCzSBHyy7JuEQPVQ17/QL/WmWhWoBjz+ir71ynEfK2MOMbOeYDHShWePXDiAYaOa
bvlo43Y+sO84TTUbXIpeSyIyElj4I5+LZ9Mx+uGX3VIr5hKnp/Hhdy1KFSD+r/2xujDiRjCiMpGH
992f+pPv7gAj1uXCsvZ+ZF8tTfl4qVTTPfCE6JfIlNXllzr2M8jISJZf2xUuqv3HATq+KcM1tnaz
qt21IwFM+nJrltQyN1PAsi8/LBr0FvT1lzPLf1I1INsHmdiDDw4ITVqhT7VlbMdpagroMHvLG3j/
DlvrQ7stEK4V3TY2HH5tO0uvEFBKzeaDbdCrRLQDjmlW9/8vVQqSP1uVX9a0ilZNBbYzqhVdecNA
af9M9q8uSYi7rKkOPp93n6LdJJePl15DzpcVXwxgUS47Zv+FYHfKPcMcMHt9I3e+nb3Nne0ordtM
OqO5HRPxgPtgcUpARheOz9kiKnNgTIQsUaLJl9cO6MfLVQ8s7vU07EH/bpOJYT7aIXWjrPNplTsN
FGFJaZUtFV/90iOItAYTktHJJKaE52B5YrDIMaQKpKd1lqfsF07InUpBTUA03GtUhp589CO/t0gr
hVbCAl3GVzJqEFpKmd/XIkCaevmyRy/LX6MVl45nSl1cOdP7Q5A4ktEl1yyBKbxawNCLruz+hq0X
xwfkUUg0E8mQWGi/LzePZoIWg83sdBKUgDjxZicXyXoyXEN2dNfERfGuFq9XX3W0xxqF4F6QX/CG
0yLpbuAChWzzRvygLriT542Danb5BGcwuP2DEIMql/cnXVtvXVz/0ClXpgoLAo7MiBpcPlE5IN07
wZ4cw+ConZh/FM2U5BcdS8lDiMjQHYLNMnUW7Uyc0xyReA+Mw9AqmpdfMyV+tftHtItzgIL2G3Uc
5QBlrevWaXIxJtZ+alC7QX+qiQr4EB49YFVW3mpmSGIxi5B+5pVyQgvnEpBsRu9wbMF+JNJuH0iD
CdT00JE3VFUDPM+99aWbHBQBEQyO0RUn7vuPoHyPd1zBRYWD/4QC8EPh157Lqr0XtFzMvVIDNZVH
kPokxYDzTHk7Zn/ZTNNvPjOamDudvfV9Q/DrRNPrEBKd/nA7uOYakglWkg9bb8GnS/OrDmPsOez4
VPk26M1e0h28Yc+Oo29Kk76Kx831ocBDiwNJAMdk59gDz3RnRM4+FUO0BldSuMTIxdsEwve7MYo7
rgn+BF9JStT/7PMPOUi6cnZH5gtlR/ily2c7G6h9pmQV/NgyYVIfMFOqhS9TVtvb1MpJANQ8YwJq
PrD/WhcXaUv+5emlJ/bvbe4Nv+72kN0vMqkdRqCq/EPEwpgqwXs4cF0BiLrm1ceIuwZeEbJphYWa
QEO9kh1lO3NYRT1t7/26RysKj9iwBZEDH1De5wG9LhnEzMLp3sLmhHmg+/Ex3KwRhXeRo1wpt6j0
qxAVsryp8bzlPoHEouon6gBG2upachWMX/X6ua4OiZyyxHvTm8oYPPIqrq+mpkoJcJr+bbCwTasb
T67FEou46gdPP44EULRFuc7yCqX6i46AOTWB/ESFFA/jygI7Apth+TWrNQVlMsAG/+jiB3N7bIqq
pskeG1WD7VDJEW9dTemL8XikQFuXkNM5Fn84tw+guzGNGhJs5HNPNMxteAC+iyGLQfrVo0M346+y
kQKohxVld0+D2rxCyA8G20v5PtVvnIxE88pbEN4w4vqYRClpgEekAlghwC8QCA6bO+34vTC9CmHw
od/YNj3dd4eYu9UMVCQtvrqso3A1+ae67ZwdqeYUhRtG477YR8omseWOv6qv8T4xiMrS4daEaFOB
CNfHWslVlFN/r7cpn9M8xdiPJQnj1ZADscE9xw+rlH4tT+w49GyMngwtju9ugjckQc4PwNVuLfb4
opAnUNlsEhTK0sq25k4edoY+/SfLMLyjm/RSMlq6C+ajjLdAnlalYDiojdI6kwUduHDdVXCJ6NSM
K7gFEwRHVDOo7RSVY37mw6/w3MJxEgRpOagq+TGjSbw1eIfsFQZoWkF0CiU1k2ikYt6f3A6R4aWh
FIHJcO/kBG3VC7starQrjmLMJSPXrt7as3pZzAhJ7b8KzP4/+1BPh0LuH3c2nc8MynqNWKhGHWKv
GI4qyYSlMGCnN+Dr7fmqOxJIKW41qWGD4LbNME8JZftICF/0bjEBlL/1micE36IpYhsTQcetHd+n
IxB+NLmT/x+Ftd+V2KNn56JslHPHaYqV7Gsj36Gngd/Lkz9j5sLOCsJKDlpJ4duZXmbSrk2KrZyw
UtUEhlMpswBEkpqmOI1Iy7oso4F31oNTihHBiI9wsXZLPovJicnJTU+ksCi406suoQijVq4WJPPU
+xaRuqSiGyXSUOJjP2tvYMwLeIF88c5YyaHYWwczLS7Xt5BlC3lw881BkIPzV3/6oYe8ZydN57KL
zCAMBnWd2IEET4UebVoUggVO40/MM2QFrm/Lsx77VlX3QFqxGKRLCa2WsI870V24HyX9oXRlwjXx
YBpjOvZgcU+g4PAqadiwUplctyhiHazyWJ2tSvGR/0zrn+rJngQ6U5kGw/Puh51MW1nT2Gdql1Hw
K8wJvBUOorqx99ylpybzsNMwO/XIA6tG9Ft8tA0TSTwuYPK3G8XetafegtqHIpxWhdFAkf4f2lmF
zCyrA9HrOZEl8wSVaozeXmOXzOc38NA4tYCsmJbxvl/2lH9alAmqZ1OOoUaDZ/b+lOhGeLdnouvR
ffHdB2aGE2Lng/szJ728pu/JhgLAiDwvVIev5LdCiSk3II8zDdcVG3/2loUeHx9ENdNp6OcvXZZK
uiUFciVA1j3dcZLpBLR9HUfsf8vtVCn371U/xBdI3kkCSfJ1Gepwl9QK8kECD5HOTBBnmW4ia7jT
rrFHteGdocEFiR7LLqXdAypBAyob9Cp779xJobCCwGwVeokOjgevmv9S484LqR70mNAYWx4FUWNw
8wJbmQxjnTHKuMNu+cvnFTc7ZpukhaWwFAG89PllvVuufxWuB2GuZ9iZQBSovDfkyekv9yVBEPt9
sL3bdNfnt2GFLla2pUqvlMx/d9XyWQD/CT0eul64eMuRn/P2m5aUXUvSqnEPMh8YfvvheKbI0CKB
M2TiHqQicoCQ+mKgxLHFnquijA2IYE+DxeBmlhMQH1pAmIHueTJ3NYHS3bX/H8gV9eVwEzxWhbbp
mExQhWJyd0US/KgIchbibOSyK7svx8W+7XrM4ucFwt+bH2LgGg4vx0z902HKbp/VsduKz69/l3SB
3Pu27gzcvbDuyu4HncGfuAZ5+bk8Q2W4ADZMmw+xQDaDNu9q8EyXwUiCgp4Dj3nnTfCbYVjpNN4N
ACZSD4N2ID2aV/CsztY92y6PG/Ua+m6QzDVr5GR7IrUeuD3l7RqsNFY8xZ+BjjuVDtLuLj5cuz9L
Zofvm9AXabxkzDNaVM5zSDDMlbYMVWd9+L53gKwybWuT0SMhfFJSQ1R+8wSvtEoYx2RPahGKrDtl
Qn4RW6SX1aO+mj814ZUisN2EqOfe0SajjiJ5c9ca2JxSNClwoY+WBjMF236mLj+Ibtul7j55vhlS
tx5eSMYm1jjQVMD84nDFkTKdcTgmgJc3drfgXfd1UIh2/Y0IX3s/jFS+Lxul5FMrlDUBQcdulMnX
WjWJoVb2C6brfjrJswM9qZOjDoOesZd0eFq7vjpXXz0QkyPPIaCnJJpOnAZP/tFXEhxLlTmCkDXJ
Z6Bnnfq+vA4YlPlXf+GZUZHt5uhvXG8hld4RZSbhIpT+OW3zUzcsICW1Ja8Gip03t9Bu8f12YUsc
g/OY6okQeaq56RvvabBUHTzxDh+ZNphf/DiK3vHBpnMngXoy3LU+wuwCOfeWpbFYHjZZA+ZK2LHf
QvtRCU3rMfU/btVxMZ7xD5NpNICpZJ/wGP0iyQ9gYPWJvUqwgzxjwQhZcvvb1ytoTaNY7c0u8tbJ
+iUgO/bYtdUGre0QwjsNKF2ode3gG6HRfRmsex05UB0tydhm/Rs7oQeEnEWVV8lWva+63qkCb/Nb
/rNeJH6MZL6NfEcVdgJCi+y7jxLI9JkAvDSDY6TbTCIb26AHe1Lpv2wF3HAc5L60A7nyr+2nisGx
07LljHT/BiUUw0m/0DR/FBNaiB1BR2Q1bnzY2ww03Ay8voi2tg9w1OpI2RE1ZP9a+wTjMnwI5kUT
wOQ3OV8U8RqEqJdNLTMzwT4Z56lqV5oHUCY86MHgH+rcp5gGGOYlWZKqwYwerHacwnH57H9xYyWi
6FPodSFVEckxO9BF3numfuE2bDlpqkoLHCTr1BvWSnt7guegQiBZ+Vu/FAT920qqhbJiinNeluzI
e70RCqoJto2vRfW9asnyZSfQlpSGY0NRaIgL4C4ek/Q5QeK5Wf+LRqz4EknpFlLyyps/Ui2ph0/9
UpXZSQFsRCRKhfHXHHfVZhSuh/8gMRhwxAMSm1oHwJm2awEHZxL1PZOlVLNtqxc8YvV8tgKO2hwZ
0XZIyupvHMiwC3jdaW7oyOs6cC/ZpJKvt83V7mTLWxq5rU2yTVnuUUz5T0lGVD05NvY5KNPqysfR
/IKR/CxYno1HKNWIYRSpeCclcr/0Hx6vqNpuUL/4ksYuX9CuZlQsnqEk24NfhTocAhPiuC3TRuD0
4eTCNF73unsyF88zr0TOeFlhAooqXzwcxFoVtfsEIdnDid5BgJHwlTN4DZdco5Glmo2SwSSdi3yl
toMjMkcwVuObl0wLx3N/1K1QlGNDdTAiuIDB+IsAUnS3gDe1olTvSNi+J+zuAXXeevb1f5d8X2XV
btPuKetYp88qGj0weWjZRIrXJN+Cz4DYU4vghs7BTdIdwcIuOF77rCZRVEODhI/nXyoyQ58bEm7c
j9HWvfMANUhx23qRSLxN1tKxyUSRRHo6T0v/UXXtQe6RULE/sLKHhUjx1UPPA4GfvHFixu3yriMP
5KH2G6bfEKcHIenlywrUTylbJB6culyj8uiH6Q0rF6NH/dVdWQn1DhNzzn7/zvQxf1nX/An5aXI3
2fofVav6OGLHi47RFLb12JVo/RzFTxhnxIdJUVXgiRC7w1qbPtZB1kbQjjkUXDaXItYCHDhK2048
+20fJyZFkGarU6o/k5inuiJ02gZfDa575f8zrGYmeS30ai2S1GdoraiVTrd+OVdYQoJy5+JLbwxB
sebLivpPQCSf2BOA66acT9BoFrp18VHiTEIVqDiY1icdwXDsYg8EfjBQeIRuT6QBv3uzl4QrGJZp
IWwGLoGc3TDP2KVMMFJ82y1RsjpYMQMfw/aTnQIY1wBhM+N/1brMxAn/5awO7H2/zAsIlw7HQib6
+/Rma4bu8u+HDvyub+H4NyYEdS1qyQ3dAdLuWooKZugGbu+tf4PIaMfPg3eQRvX7nTeKzb8Q4nGE
enK3GYWJw3SPbmC2i2YNZAVve0Y6WwATAfBxIOIC7tsK4lLSAuAoepCq7pgGQtdbTHTka0J+Eo5s
QXjIj/FrcnAhx/l6nhDAjAmqEXcIurp4qDH7VirGFKdY5bs7j1VtN3e7x5ziAhUIljnZCEpjejpP
dPOTpoywiG2vheI9/KaVbutuELPY8g6b7qlKxun9r4ZAjyOLE0z6oUa7YlqlAkh1YG1ozoDJC1yF
9J9eCko+02kM8wIXGYevi/y9D4pVXRzdr5s4NCPG4tse1yVtESJwShmu8z1Dct88cBO8nbVPsY+6
j/dFz+mKji2rpfrxnvojNyB+uKhAoikssxYtMIqNWBSf/E2T60ow69TyNQM4ih4IKWKp1XTbWMYx
bJSoNI6dCRI6UydpYxfBxV6/WYIj8drplg59VWeivGliReyricyn3nDH3PYy4naKHFJamj8jx5Z6
3LIG+rtEPk40dtFWH2qmIXlA9zjAydYXAL11rqU8LSBfdxYQXHD/zwsHiy5ijuSNR31JhwFZIsvf
0eM1sLFP7iMVeBuMV4srGYzOXEdEJ7aACi/NZjyZurRwvsHzlOUe00en7dXF7gSV7CMErSFKHsHP
ncOr1CJWn0s/mfhalg+yjO+LajSc5fBRGK+aIyvPkV+hEMHXs8MiSmg8Y8JYBSTc7i0PoHBZNFFV
wyNEWGuhAy7CLBQrl4RBVtpFy6k82JwRUXl4HqfgwVpi/5zf/2VPLwDrgA/++Saeqz3G3eSiobRe
Jl0YRWjov0/Fozzp/9VioiEZT1FbXuJRwH7KuqNyUEL4GszAV2BwgLVR1e5u5XJjMbCpw0Ogs+rt
PdBnIRZeRXFbDbGWjcIBHgElrqJrWsflv4N1eljP4b5WF0b0Nu/r5m8FIjcapeFX1o7ayOoHI0dx
bcoEPmnbhS+C0uJ3kAgzDx8oXkpT3Q4LQXOews9flakHYIBTDl/EN9rMBXpLUh7n7Cz7aaAKUGzq
rTzmjmldbWsgMuDetwqh9B1Veuo9XMCvZ6a7OWWLrxFR2aHpG1I9RUiVPxLopMT1AWGLDhOxlFxu
ZwfvOHFeOE5OVUO+QWzp1260rGRi+jaD4P7XtnjKJD+wznpm7FLwrGlLZX5Rqy7LyjBVz9XtQyFd
Iq4stsl+CkSrsdJGmzNq4uTAMpf8gkI8aJlwJTcwFuWFgPJT+oJilUWK5v2yGoSZN0lmffhVmNrV
T+yJ4/Ykv+uE6DI2lxWizkeNw7mL8ROgZFIrr/QWmjNqlu1TwLppqZ+jx5WF0US8SIbPFAfPPxs2
i5a0cpmPkWfHW9e2sgKg7/UHLu40PIrGNHR/hdE/YViqpa+VcOAtMkISiX0sxe0bOOBoSL3gL/x2
aZQFuALf2OG8maTXp8m3HmO4Et9HMuNFLtg/Wiyib7vuSFZ/IicnYxnGgXWmfYul+4p2JczaYWX2
4tglEFQSa1r2YcL0c0kAdkPmjhbnrwr3IRkZYKVAMdGhmbyn0Om7r3AzP56qrnUbBHi1/VBgN7f0
X8Ye5f5kGwoV3gloKEP4AmD/xBtJLrETjMRXJrw4v1YfshXbQ47tBzc9WYFzV8j6A4/pS0oIuzAt
OpFImMJawX44Q4+hh8MoeM7egqukkQPB3qQbGUEwVpg3B1/TvnGjovlMfwq5fZxPbSavIrEUpQSY
mbgUqLOrf7lAI7l35v2FliwlL7WDzGzfVKdt8ZFqHFEq6d2DTOid2OvDQnx0qOEUlWMF96lvHnog
aapTk7mZh89Xm5ZaAUnkAFHlpR/+ww+TWDwp2n3ImWWV+4PiuwW/N9f+yD2Fn4Q5E5+Ziw19xdXB
cxNsb0wU9G8OIbd0ZzNAbQ2PNstddwGAKYnwwNiL7nuLZPhf4GWpN6uPBIwENTOWu+ViB4vpeonV
BEsr7jEoQMKCidbRyQ0bT+HATdGeHlfoObqdXGxKW1sdCDFZHCFUG9QZ76OzHKaLmUvQUjH7BG/f
sTBIDOk6WWUATwpY76jmxrwJTTcR/cqnE2aUp/H7FUPApDdorf0+RNaKH6xOkJCCVepaVe+/hV+n
b+78VgKbk1lEc81VKmt63eP9KLs3XnpeuhEmzeA8AUkY6WGBetofBCHTrqBGDdyt+KBktb1O1GAW
/bOXAb5+LJY2aZgs6RdKzlREYl4y2GfCj8o8S4tGPbzt0lXUW5ysFwcS7T11VEYYLEybyByH5+B1
ghL2ET2BRKvLCBA289HIYys7NikRaZ5lsP1ZjwCVWoz+Y4XJ59zpyn0HgnPt0s9lKMtampMV+ZTq
Tyzyf/j76CMrBN6BWIiqq9iJtKKDhcVioxq6SvTiXlvgid0aCvv2N1ZYx2ZaXPxFG+3nMR83wPMZ
+MT7KLcWs0i41yWPrmwYhF01G8A3XSR/mX3ZT6HOelZDmCaJwKLe5hjfeDKOdYECAtNfOkMozFYs
CT+f6aSoL5BX4OMNEL2iFlRmN860rBMW4sShxa/5Pjn7oAnyxxae/0W0GODFRUM401LSq9rUhtl3
gqWHdTBB1vTRdtxjkXUau/e0622cVZns+ty2spNbzGrEyo38F5/qmetc5KWMLnuFzFUeFB9ggkBK
N08ubkxw1ORRrIL2qG98oFLz9QMRMUi0U6Pp6exlvifs/8xRIMYqEg8r4ggy2sQJ1wmyGhDvVznS
Fb6M+NPselfuhDHKJqGgBERKAoVt2JkBEhMwHqZAvNsQ2YLfCYFZdRzdlspwlchls2CwOqSlsc6o
GEMcST5m2vP2+ldeqXW8toIpVQHve9f3J4rqaHEYC2+t1GK6pZrxYL/SZNgeGaPsDFyYNH8iwb5V
UhDmM56Vv3ZIHISyTbp4IIZLFxZaN5L+Hao+qha3j8xmUL679o92fk2gBYhtiYvVdbL9j+f/Cvz1
RgHHG327JGz6hp7CIOh7RZWeceeGbHBjtLaQqoiODsl7mAy2YvC14cd8r6q0F8+f2/SSV4WvSzad
hevQ8+IcE71qIdP8d1d28HgXsHdWuGBivwDFy4znmbJyLGsCB/YBABFsIlRdzoc+gbEhSpzVPiNW
OnsHBXwtJ2V9fo33wHlGzTowfZ3E7u/7RIO7C2CcvNivoDBiUtY4eAHPKKcRdZdhojuVrLK2MhTx
JCZiIGJMOLVUK3smRUsY0/IZ50oaZvkowFVVvvkfD9Bp7IhBQ0pL8CuGBflJEEmMxA8wfTP8zukr
HGyM03Um6DDfHI65PjS4hlAMaga5GkzBG/84iOjJudsxk7FLckbmAeztbJRBCFnZEDCYm27UUXLG
Y7QBmFUh8ux2/kt7uNHdFHi298ChySFgbp6YrtmgYTCc+HoSl27op+1Gja1TRqYDXvo3/kVs1bjh
f9JI0qM0ZIT0yZuaqnZx4qbv4YBOfX3oFjmd1hKu+ssFgygxhtf+LKuFxAhRbk5GdVT3KGK4uV56
zt+QTTxdjqxyS/2rjs2baCIVPBmQulojOQzSdGIpCyuT+b3H5eXsGvxTC5Nt+2gasldkT2MejUKl
TM0Z31CSzv1E5Ko841iBXgxCX/c+f6yWWkylRohjUwvRLx5Assxro/H3KSeBjQcmkDFyvq4HPwjx
QhTsy+izdfCN55zyDsg0CjM2iqWhjCAmCD/8eSerRMPVNeZ5M4ZtLwqsRWACefGXhtylt4AbD9JE
db6+zZij45pACRA+GJsHUTJHFslhrN391NdQNBHlSfKjMPB4M8Av/iQ7XtKiZatigEcMgjJ26R9Z
SVna83KSGxEVnrMCS4GFG3XWqS19owIusxZFayWSiN5rmYZq6BkwJGOT9qahOqRsHyeoudXwFqLa
OdBPTeFnXFqUu+nHkR3VY4CMK6A5hJQVpp/JYUl67cBRQwibHacOjI22+ClQKsEa06R59FiI242V
aVtarTwGdNzENa3YWXnm+4c4saUZK1+JefJp9Oi0pt1mCYndyxMohcrORESGapJwhF6xhfk+ikdk
V+Y9o0s5alm1g7mEnI3Uioo8sNqHBdpAQavhG3UKJq00WHqXYB+PxARiDd9CBUPHOcG44CM5Odye
9dqxAL5u0slXu4NT5onjDKYSZVP9vG7GxX0gZF2qo1eRreJu24mSoW3LvV4i1ioaNzLYLl0hYmu4
PWilXYiQTg6vvsD0MxSQRPeezAxcWL06Ii66hG9XVfZ2ObGAKlX9ZCfqy5mtJAwGhhZikQ8jUZrH
z/jmA0dJVl+3UtiFOTATqzqZtjZJcGEGRh6Fe7zXIAcoQvShvCP/Cj38hNjIDIi/C2biC4M1b5D+
E9sAhAVAUWGIw43TF0XS9QSzobnkI3C9PY6JwVy3gakm2xoN5wbLdjKztUPeevGsMxtl0KfPjoxr
B29CwW6Qp3FJYZrrK7ePR7MsDayn9nRqBd3s72UAwbicEexRsUUybyJ0ZWD7pOLFpAayX+ElP2CU
mxFVBiXOf7SwVU0OxllPlpZHj4zKPySU5d3Dcku1VVTcl/mnRhUFrr91ZaYEUqJGCq6AOb7+ZRaZ
THhfZWercTpu9JT+g8oyKGUw4auZMUywwcjL773+67yPTO01jTtJkUWp0C5FuNjyCuIajfPWFsAc
+BylMLmnMafRN5uLtROU37Mt8tKYhfPn/T8l2YWEJ3Jlh6nTpgwheudRinyFPd6X9Un0v3RC3aeO
WfJ3Ns2ky1U8l/DpOPQyUCjNzItayhBy0j0JYhxzbEo5ViaXw8FiI8gkoZlunE12KppkznbNDICB
41Ex31GLglLQFh3p5Q0vXeSTsg3kDQOKZgXKVOl6e1dxJASXKHIhKEul6bn1RZPTinu1+s3YReRu
TOk0Q0cMNlK7Ss42ajI1OmZlK4ZmRpEWu4ubJyxGIJF9xY+1PJKMbaOllS5aFxH9Q9FHr6vrMwu7
tHnIOIU2SMYy6tm3lN0uz4KUz5BPaPosPlu0O3gHfNpldV7LH0yvD7gXINM1ArV39j99mZXjOtn3
ypg0/HcQ1xGHUw5ZU7/80b8kuAZ4XybzqPF7si4NUwdFhuu/8PFE+vnyhGd4Y3tqmozlM87sjban
7ufnFBJVKYugUsY3gtgwscTjyxYfQcI04r4ix1ItRAG+vuG6RKkDAm6d3dHoylgZ+1pdn+pSkP45
X8dCYcxhC+NuAI7n9IM2GtaArp1fEw3aN8lNJxOLg7aBCsuypxOPWtyEHinsprF+VUKPpdOK9wkN
gV2rStnwGPIZIH1S1LBvGYgfXwWJeEO0TdFfNz6VDaxwN9NQZz+Q+rPPbtwyh5Jds4p6YgBKVSx8
bM1YQzdw0PNV7r1ny13pdoNhvVEj/x9mkEib+9ltdIKRvD9McEEK3bHDeCtiiSTWm02Biwl6DdAM
7IT1t9Y7kUnz9s/9CMj2W0FODBs97BR3C+tuBGZ+VrKfUoZH8KcRK7NPA1fa+nEgosmLP1ZowWp2
JZcRU5RFPjrh8ALCDCUY3YXXkWIeXuekJfnGCvIHmqORcflMqgOphJxJQTNB2rdgCHNP4QZafmCr
ouSLBLsQo1NKo8YlMXLQZ9YPBfh04jnQWUU5rinYhYH5LaF7KhV/8ZkTvqcoT9NWLtjI7ClBw+tq
gYt3CgLJx+alhJiJsouSwLysLLSxhwxryW0LcVU6lwlB7B/2D4lsn6oKD1spxhlPsOTd1F9Zidgr
ZzzhLPvEaUt14wzktKKecwU2cSd1bBLJACq/uM2kJLgJpkzY1AqjcmyVLJrwpSViSRFabAfjdr70
yj8V2thBD3o2nHlYDKEYj9mp4c3AcqfZ3lGWj1c4Wt9e3xRwykvjZyxJtEp2ZNAUEvPzKxkmWwGy
yQdbtWSsIxJ8yhdHjLj/mVVxNoF3TPyzWhtXAaB4tNfueecAO8nL2vNy1a6sBZJpBGdIB3MLqO7Y
AH+Cf2NpvMKMrxYk+CMJHUSNLlWvcK3q7FR7vEmOA4NLK2nWwgvJ+wQFJ6t6lI6iTPs16H8fjyOs
bZyTAcuGTBypIeL6X8iCF4I5AHNKBUesTADsDtEDb8o8RuxGBQ43PU+ruq1AjrNbs4uzp+A9IjRv
ECHa6nmkhuirlDkL5ZpYe71fIkxZeOjI7yF9XO9buOLJbUSPSPdggGIrvYSlxQOVe/ciYjv2aXCW
IMbrGG2idCKuNxuKC4hyXuHHZXrBht0g0Jp1wurxBwzPfccAet69obeqaUBaJTUyLCqtqMAYU4C9
IvmJpHqEmf/nQNPKMw1qq9ZFm5xkx2u2WY7SQ2pY0SebH3CAiKCNB6YRh92CqOYM1SoZlwWgOPFj
aH3PJPP6fO3HPZVrHrIKD2NYRNx39WJvMwrFqewihNTct6YMU57g6Cc23nL1z/OasaCFq/0I4ENG
ovOY7LuBHXY/UvfZOdJ5DvBA5rIQ71kU3g9ghPE2k7KD0kIuebDiK1knm6X87uW2D384BuYCVfIy
4j/P5x+p6bMFdapVDBL5/AGSEDHPxowNVnkfuP1FavSdZkMcBnBRHpYWnm43ZpFZ14GXyoJvwf5Z
l+FhjUzQ9IFeRNU6icfw/C9pDaA1BoCnC6j/1JT4ztNQKqLpCHGJGE/7KNc891hRlku6bPD11FSa
ilvCy3NrarYWuKFFDggVBiHC9Xd/LUhMqKIfmC3N8EeQEShXgZkFTFAqDFVRNCH/H9B62e/OWBos
pha0BtVjNo8Yd4EMbVSs8eA9QSfY07d8UwgbBcOTLF+GMQY6fBCBBFsc+erOmD6Piagi0DZF+ONG
XnstMlezGW+r7lAXS33QVE+gpbLm2Wr9Bsur+WARjSmLKopNr+q6ncOMgt0WWtTKDhTRvTfnH2ts
m8av4Nq8CcCh0h+QqP3lyVDLOeE9vP7/hkxZf4XPshN6zWz/3FcClOItcE5FfNx0Jv9zRXTrWJYz
0tbadBa+hhifqCOp2qEGCSKg3GODb5V2nipFGDt+SPGYvL4UbwtxXN8tt8Z7bhqbKSzAOeSKSn7R
v/nVCoXBPuzemx/IQMDsQfR1l9bHQSB4Uh/Ez+yQwScu+cWFLhzEM1elETWfW4zNmc1xwW3yoTN9
NURPjMxZHmnDFD4oYaG1y9XCH9tw7GdmRCSo03StGVafWo0TcBT1vFngAO0x5wDKgWeWIOUo+KOm
Zr6wDlR9DqDhQEbvonQcYhxGJhacgVfodIUe3hVZFEsmgejz7ks/+qA6T/fpnU4S8iD+s9pLzwAg
nUgIOR7Dbi6CaL4AI5CluaRR5mW55LDpLm18EHzV1DztQ4T4S+ARjg1zAVajwq+XPumiM5j7fjYF
jkkuQNm1WoGxCyMVNehhnh2Vt/P8OlpCndB2TXC9MuRLAqhjZDWa2uEO0qX91y2n0+2gOk+t5IhA
hTR2mEwqxXav1hMYL9yE9Z4xxs8OPkoFCmn+5X+0HAZF7y8byKV2pQ/leVJpyEdfT5dCV0pNn1zF
f1gYiv03fAW75bgX359PQAq2fx1eX297evsj+ZYMi47Kmj6qRRDHecrxY3eEzuHzslMviZsP6JAh
Ui6enB3tPy0+3aAjF38gvHClLr1eQnosDmo7krTm0OECL38TL4K+C+qDD63rvKzj9ayKBPPoTotR
xwg62Y4dltc0QV/lG0LymF7R825Cs8JnfD92oEE6W5EC9AJ2CVjOrqATblfz9xyH/AFAeJwZ/1bn
aLo2og2QL733i0jbzUAMMuX+rJz1k0Bfbnv9BMRbks6ABUMr/iTCj6UUyFJzaydf+cYs2cnNHVs0
fCoizWYFcR5QFlNKhhnxYuYnRGJ7tiq+lHCl54BiO5RR4Vzykr/KHfyF7waeSCOx73d6ZjQ95OwE
I4jmQ4nVU/vv5y1rNHbwOt5LTxjZ8eryCP10eOMoTIlJdQOBSTTOZoeVY+JU6p8fEUtFXxnmiIm+
LyTHIZBrBx1G0jfpMLY69/CqdwQDz5C2+T3zU/ETd+7hAVoYxB0EfqH/xUvbPnuwcyloyZDILrMi
KTreXEfpMJWWEA16QLAtdPLbh0kVam8WkBBqrQuMNCz3W6TAHPBcnj0D2dVlEVl+On7hSs3IJlwr
m1CIAypgIZ+O7Z5quTCX+gUm40ZS7Quy3pjx5+mye3kVm3yJ8QAGvpEuIblkH9VpKnQFB4WOp4Sa
oq8KV6IXrPg1ehiwHTtaSGOE3ujTrN5AzmXjJH/JzJw/Wrro7vzT0uQMeY0FEczqKY1eUwLnx/5C
mcn/N+grDlGK9G3px8qmwGJBRJTFhthtlzSmztUTklBIiiShqblWg2eMkkZP8hO45X0mhuAdMYnl
J3kKJ7jOhgdDp2H4gjkE+fRBXDN6W9eEzH19zgGB05VLjRgEnEm0dABFV0TrFOKI34knByScB5U2
oT20rTCDbKYEQEz0IzaiYSNKOHxpFEIS6YiVWpoRIlbsurqETqp1lRwiXRzkLq0AvyAL6zcCM6ih
5ZbLVh5JHi8DJ066RQxoh0VC5loi3W0/ks6QzyaaefhxKz2ePcLZ4Q/YHLBrRn4RtkByr41aO4ql
FnLKn5/+T7ytU8lXKmJmAwuKjSPqwEaQ0SU/cJno384DvaOQBZq+gIflTfhZ+aAkY6TlpXo7dmPa
AOv7aWlv23j01w1MYrsEb5hO+DRrHN0wuJNG7mo7JPdd1xQPBcKxz4Te2qjyrR0f/RpXxrgjy7+U
exdlVKyQF7xuPA6bw58EYquMYYesKwkUQsBeSjSGW8BpdLMe4NmpC+DPo55frCYqBvYnWUybO93a
p2JOTXieEkdjBFKZ/2REHtuRhMtxJ4FwCFuTUTR25QQ1FN6u9/150DvTWUsHyUl32coZtzgBPnVy
5s5zxQdkavfTlUNEbgEm/XpShZuGu3IcJL27xSriRyGJarTNkoMWlpgPmYYmUzsDU6jnl5Uv0Dyf
mVnR3KaJU47XCEfD41r4xwoxZniWMaJE8c2zu+fPdrzcoNnyXGVemPvrmSxQ5NOvyz7NrXyUJmEI
f3iSOYmmnQAySgkCgpNwb5vBaqeLwe+t1Ig4ICWZpJOb01DMGpS2Dj8bfTsKfNvtxpPabv5qKPSw
kJfq9IufDS9dxXJRN+eDV9M16T1VlYy855XpIzVPoexsMTA6ejgRkeiG58OLfpNEisSguxfi2ORx
eH6yRGvAPbmAaqzANvRoA1FCmg2fRkCvaFwr5EnDxfV0N59wlj+bnybbmTszp4NxETwotLm5BcY6
fK7DVCANRzf2+BAWHd2ruDDmPIQNM2KOkPUJPsF4peoBFip+KdiUDZjQhZhav8d/uaS7K6PCABpz
Sg/dz3E/PgDSmISme0MWPLawbEBIWVweBS7G3eeB510tWLQ8yM+tJIce6LF+gbWEFQY0zTHQQk45
vc6yx+xZ3TexumNrbPtiqFKDALq/YvviO01evUMYR+37c8cbQ2Ddvr2ODEJ2OVVy46UDX7a4Wubd
DJO//UsujSHfMxCY8e81YOgZsDQ6E3bWY/04ZT9dEuFcEXKLZzKoqKXaEwj6nmWCy2WxX/sAchgo
faJrzSvUIIOl0Qc3cKpnqmKv9A7LiIcIu8HROid9WucNZo66p0WMFdVRP4V6uhQsY9zSIfXUWZzV
t+XYFXZDSc6/KFGGOiIk3/uNwDLW9IUHL6XnxzL+EdoGAkxWdtNhQH4vt/OUveR0bPDV7HbRKxTS
sSjV/qCgzF1dbYvxDMzOAvCNWYvs4BgKfKV3q1HPd5SR/FqKpkU707QY/9aHe+5310zspGH9VCO1
MkEvsyU6eaTxOfueYikwIPP1zOFJmSQQJg10UWytM965spepGMoWDh7co/am8DBTLsjuST/UJjf4
qH7bsf3uvjFD8j/4VXZtnpLOE/Ghf/IFQXHOn9zBx6/77259jpKF4JQ72l6j5M9UrUkA7fDEs1WK
KKPDAjVTcztNuRp4w6vtZfQzoRJjIThVSy39LZDgbuWaTYXLZ7bByCR/gHc8Rxo+07n/ZqYe3flT
pwhGOgJYei9D8jHhvGVrQ6skNGVGG86tUFqm0zu6tDk320I4FTSVjbaD2d8W9zuEMXJZmCHVm+OT
TMzLDcQ4i4HNmA3vXqsU7SKN0HSgWvahinJiG3mwx4+Sd4dlEaAg2VpOpbt7VM0ZLuXk50ZgkGn6
wuzSzK1dz1wIUCyx9Wr4Y9nWU8OJ+r1ROXPDYwG8dvZ5HL74uOSjtxfVEVL1iXq0dwuC9DtB+omx
WTrZFPQfUCmqLXyvHPTggLNdDohRh2qFaz+qkK3XBxRgqjmsyq2WfIY33xODQXW90UByBu+Hmcqg
LyUNrdeShtk2ouFd5Wb6Vwn9G5d5Jj1dT4x4mL4QN2J3I0gRi5GWXXX0U+NZtPetLXz2wEW39dEq
TU2vwx3l4SoQ3h4RjXcsPGk/3R/ENLcTp97cmJUWLJbefM7qqUHl6pJVnQxdC/QzccAwvmBToYOp
zkkYKppPn3ljTFS/+2H0uGntdkRNy78X+FCyuyPZeeFnOEM99+mygnce5OgYxQ8RqD16sUXIpFIQ
JI7ov6zI2WDULh2pdY9T5LYRHR8J0f+sLa4m6iMdHfVc4irulQeHjqWCpT79L8fo/ffVI/O9BRUt
DRC+tAzpHEvLMachi7B6ebQvebt2puI+FZHv3CGhXn/p/exSYHfizlC4KZWKJRkh1ebHCb37cmHs
2VssjElHgcuq4Wwm/+MbBDcy4iX7QlsSXM9Zp7ar44UwDADPFqNAlYg3Z9MguNOhQVg90m+01Q5O
whceNoAZcm4GLPALauHVyMDR3VktCK5R0vp6mzuq68OWr6KphT7mSSl1qEhVOevsDCr62t5PE0Q4
JIky03ex8iYjrwYbCjUKen8enJEVw65+1bL+sob+i0NYAUzWyBiKNJ9QDwcXT1Iyv+Va65bYVXHG
s0ZyoTGVo9hKR7L3k51DtjKqBjbGMs02x6e3IUhYNkGcpfdD2gi20rx9ThkShLkpAnOFVSjogfS0
TFjWyAsEb3emsc8hGDeKxzFLuuRPmpxI/5rVBCY65RACvbOnrdZfpGbRte6SFHmv6FS+mH713BMp
k63FCFHtCCEgMLYowzVpyrsbjIWMg0Ytk/gtBG3Z/IzX9jKKG8emTpY3hqssTeUKFO5K8HEcAASX
1XxaihdmnR54fXiYQBKH23N/76u8E1PoFZ80Zed+DUDz+d2pQ5tJsn3AIZAZBqBvvXSrd7ThXhq0
wteKujl77J1cYsFcQEc2F26X5ALU1V3H+AWwDGzdeAgRjO0bl+MvuRv0RBq/yhgM70z4eAPR2KDz
CbDWg4Ht0ldMTzOI9l7BMZycerjC90iS8oQd3lFnH2O9cWYXF3LWHl1fSFnAJE+ciswTMcEBvk78
0lb9beyc84AQaGKzE9X8PvZG98v6be+0cBOkBIV4sJwMZjv14oy1Gqyc8huqAKkdhbpstYL06r7e
qXPKVI70hpp8EORUjP7yplE0kVqs+AYnDoK4uUhUjy2KQXwRqhQSkAxhzzAVvo201KAjehCkRs3a
p3mtd6LVKE5cBGm5wrrtBP1G4UeawzJM/oryb1kSLyrDtsplD/HB8Tm6WcKeJzvXDqtg3K8IH6Ge
bVq86MpE2Ubl8MaUavu2g6V2HB235uVeptGqId2rnNRMa1fpteRGVesyV49/MfwEOzy/DtKRiPEP
3NAdDsPbUHW9XOFFIE+jkO4Zk+Y5O3ZMoEknLPMmIUqMGvVFS09AE4THoaqayuD950sT6fr9DRlN
Bmmoxj4G+QTuiuhQhN07OSodtA43LmiXQSl2VT3x4g8x8tAb2FghpejD+/ClneJSVPoak7T/trrf
WPgkSkK6rMBAl/lZRxV1Y4GaJteQDHn5lgh4WqaLLXquVlpi7N3oGX5qDmGBtraW65OLuw8VD0+6
65/9xmKdStfwGPWMMr1d3iTLhuw2g1Q9imzC/uqB1I+m74qb+Het0nauQSuv69cxgLtYa90esdXl
Iceb+5aikruLBxYTnwPAZU2YuUzbAv5FrPT1xJt7co+QPc0ZyJmpbuEyy3COSSEDPoWVtLwoD+7Q
fE4X5KxpAPMwoP7moyC5MRnzKdXFO+K8aQ5gc1xXYxdZm3aggHoKGYFavkphnad7RZXDL2Qujz1K
pPL95fhocKa3qQYaec5OtZDVAvVJVgG723BcyNcrlhM3FDbcjXsckMhdSpsC7Rpcc4uhEtIxv1Fd
4bu6JqpkwjDJF4uphPz130vhM63AFT/oARpYGIXeYht9Y9ERNluml8ey1dP4Y9HonL6t4Iw3yuR0
7h4OCdUTRZTyuNfl8FB6jGT42uRyaWkFmnbafhzO6DYg5CXdaBKCSnCR19+1auknOnx0I1B1l33O
z09h/XGy/h3/JVsr8m9VJu6xKu+iJc0KgS019y0Pq9HC4+fjo4HVD0H0d8ng5TcAGtQMBXtCpx31
Yd7tTnH0xlFxRXYCcBhZAVGwLiaH05E/Iqfh9djtFn/JkqauYTI8vimZqCz9eLxQrbeRzsxzAwSH
fYKzgzaE+7GlaEM3tjA4LQM55rAb2oNCsh6G70QapDat2kFVj1OUJGJSbdU7v4lQTqKvGBy/B4zJ
RyH4/uYa/ualV/hJlB9so6JhCRBoxWOtcpkHfvjFkS9DOzSfqoQ0/E+yhqU/aE6xsxk8KoTb/+Jp
/sLMmXc6Ws4rwieCnm7COjSK0Sfgmi5CrFO/SUfSz5N8G7wR2UOrFGUD2Ql6ASUpSIgRMXv0SCe0
3SYdve319nfWYuraL7YmhxTmgs3XOQDV3AnEBHNG9VS1YQe26YL7YYu1i4Jze21ifb2OVmMuUwhr
kjY55QZ5oIkxTjVHwtOfW72laELXk9FzZYVlz3O1fv73vCIXzFp9/oUMtJK8JwtrKNI4oJTTl7YV
MpVDj1VfDr0uxQ1QPH+rCJpw5dbzROExKlbRE2y5/zT6erJEURi+qE6XZ1pXsRwM8g3r1+udLH/+
BfWHoR10XrRZGjCaIKUl0k7tIIXD4Kt72faSODtH/6WadMxhTjG/ZbFP0hj6m8lE1x5D+75AyT6n
I15IRg4wHCmYukkC6TQCDpC4Yqn22TWp93TkQm6b0mM+prjlLuQY8OMBxZk3FUb5lQhCvPkxOjlp
Ahs9Jp4VDfIhLm17v30JPYAbQNCW9HSh1nLMwTKU+L89emrCFktvOdZX3p6d/Yu0FdL675y+CO5U
n8rJQ7jG+NmbaqqXkqghl0un+5Yzpi7M/gPbS2g52yBNUdPFb4RnikSG1+tFZThWCOJLQ0mx7Ej2
foSI//WcTLlhglB5pIjYouKQkD0vPa9X9IMiuVM+6yevdxIt7JsUztI5mTbowIPyZmXXhpGBTrdI
6YYZkftkg59qSSgQ5g3HWDIPrduc8gl9BLCM+SInNnyVQhLe1qBSt4+/+srbREzQE54glHLYqoug
xPkuDY6CM/iXeMDhZ8JWnJsIbrzLGWCW6vMxtsdbucg+YRToLKiSnSjpeeIwgIfN95B1oSqYha4H
xIvIX5nGLohGDomXNmQ1vAHc5rlNRXOKJjKN11b5hxDyTev9ZV8XeA5ATDEyS6VVT6VXVwiDkwLs
DpXty/alrIQde5mgiT4GLCCxpirHd4ld4KCV058WKTUriwgXgjNBcVdrS8ktvz08Rhj9aHYNITw0
4hwveJW+/2WCJEMiJ4hEwbvkR02ivr9Tqut8zV7mRm3qG7lBqAZVpKBibBhQTHTXKCCrlVUd0BbU
CQLuNErh8t9z2ezjxs6yxbB7pCCsMFLK/akgNi9J+kHyum6sG7WEBGLkuRBq06uagCzKaObGTvbc
jUKashOrfe4CfdXiz70+L2H0BSvm+EHjEXhYHkn2qcF6hfmYFMbbGIYSfezRg1ONPylv0bte+YA3
G07a9ECqOBYEZZLS4maXxlSsebVvuLNeQVN3PXo5mg2f1AMPpfzEypS1dFwKangZ8RFjNKdFQvPc
5luMNPOpC+C7xZ6eMxhYIm+O4HQ1448YrDfS8RUgH12Gg31lEACmXus+GYU0Aav7HTKd8S8JOD8m
jSRLcwend+lmxU8Ljqx/WkjZOdnY1YC8zagmwM7oyomUji8Gfw1XGfiXhbRRVHNqVVQGLykhub+l
IGcAIRe66mhKiFrmq8nKLj3M6USuSpiwv/nmuAem12V7uAp+DNdQe7cN6ynve9inoHsyHK82Kiz0
URcHwAQqto/rc0QxWjomsHdB8oSw939xpxxBNoosTMjD6j5Cm9YgyCQ3r6SOMb9mAdz03iYJUN/J
Gdm5OSpcksqzd6+eFcNfJGp10+736MTnZdXkWI93baZCzNcdWTYbqTxDwWfCL5nBPn/5ZebHKAzu
oKetHJz5KUXYwDnuOpg7yGtzQbuKBK0eYoJ54lybi/G+8E9KGg6FF7wHfZsNVlvoMVaCu///3Duu
J8wDBDsgUgcoGq8Z5FejFGnuk4fIwyG2KconbBPR56E1+Sw1g7xg6+2Kot6Iv/zsEbfUsp2AlJYp
Jb5jbL9z7N8OUL08kmYMRG0fuVMrlTVc0otH6LZkZykacUiBKANaLjeDQkPsG93b37hAsXgPl0Jt
qlOQWcCJ7NulgpU0tPjJ8qVsd1wS8IDi6akbd3CXpRcOWP/BFidPJeuHchdf5QPtx0bGyHqWPkEw
XncutiFPex+TI0J8R5x+7bxKoeyI/ATrIJXU2FJjQB5chcuwmumV7f3WM2mdic48hCRfjs7rDALG
hpofOsIF/PirLao6OhqKxeUhtN5bnHpoeypggq9fZM7ej78hLt/88wk7hql3ZG0XO1mJp02ZrGy+
cJqScnoZUU19smL3c1DeF3mUOsJvhKh8pJw2L92mBEjARcWNkEn2bkTc/631ytrWZrRM+pfehiVr
vnZ6d0YcPQxfpj1wpgVyprNT0KQgsNmaKGms8a/1rZFgKYxWtGIrO3fF++gWYZAQdCRYZIbBokgp
ZYuG7Dg+5iYXcrvx3Xurvp+zXP7YaHBZQb/iaV5CQAgubjxYXLU227hyaNCRqzCE1If6ryCS9ilx
0I3ADqWvER3RXpj2OwumFvSS7FcKhNHriHH9guX8xF6PnH8cUJG/YWqfta6NHKpbRU8pzBJWeEwB
dlY9ivGH0e76VlACoSGcX9G3j8xu5QHNQkaV9p0b4ZioZcgC9aWRraP5M3fbGbKxR0UM+Gql8i4v
+a30CuYIB6U5Jwxd+IS6rjgydBJrlsmiM0AbNuNsMqjHmLxUYqaxuyP6T28x2cUoXcTZyYLtRXDN
4ov33GULt+ZRsAGWOtquYzp7qyJSnv+e2h7cU9I6DmOgmm6isQevXUY/HJ+TnKcqLiLyhHp5a7+O
eohXE2moY6fGC/93/M/wWkpV1rdiJlil9MFSZnnAO3q4pqHimi2gAMJ7mdFrTXrlzpR4yQyYmtE9
xzLUecnCG00oT0gDAMM4nbbz9kfeuZH5vFzBMtMLzsc/gWGGq+ucxbtlsPTAMRZrFVYI1X8SDEZm
tDuGH+o5d62dMj3jsZXugc577DOZULjMZn7BA7ImAu2r4IiJA4pE87322Y9OO+BcfyMb/ggEn19H
+PLzk+t+GRgGXR/q8C1LeiaZMY6vBD99wCqA6kdYAiWd/Fh0G6KCBeRfzHMOHUfje182zUfyQaSx
8UeVggQkrVav6JxDvq1j7Y5NGidY4EW73XlObrAGRzlTQPQ03NE8Uzicb+Fheg/cAJLJoC797J6t
JTd4y2Fg8e480UIWznTgD9udY6KaIXIrg/h5ZkMfRQ/vXQPY6uJqMBa+RCA4/zO3jgouf5n0aMh8
MEVkUq51mI9gRjv3K8iuLgRvfjl085mobuEMeahfx6PQfQqOGw50S7U1reAIdOtM2WJeu2gyw6gf
13NEmfUxPvo7psQqJbdyzPtGMKo1ed9pwk3X1zPW4mgksZ8CYG8FeTDylcA9fpaslbRbTGJ5LDf0
LNaJ5fV89xdfndbodSBk5UMRgDjbt7M+yV0qLva4gql9vbEOl4Z5oTbibhzM/UWHZ0JOr82LWLPg
TQBtENjp6j1JPx4aM6gt4YeuORfOcia5WqWCAb6xCuZ5e8Wjqlm/gNYars7n4lYqPiPjiNRYcNED
5eJrmanNdz6kB+PvPjk4u3Dgp+UAI+IydMMGQX9cHEgoa6bD6CCmRR5U85zuxVRcFYK/b5PjL2pK
Mt+YqjFkG+2TnylFh8dbkYk4qZhf/l84zioJQFVkFWGXIQ32Ktt8POXEo5aaI5DrwLfIE02gmI5Q
57k7r9/YlAr5btZoKZCUwj6LSfmySildVBWlJ7SBoA2XuYrxN+AjY7V1KDtuzgIZon5Zpip5P425
qlOKLmnXYL7QOXzYPRLofcLHOEVzFYZ9FjQT5hL39tyGl+FCcoLasT2wOCVR+jP7Wm9EJhbLv9FQ
CzAEoykF+mNmy9102ZikbiCcANLlJfNhkb0EItX2tEVFNmEWzN7mP2d1MNn7LVKGw1dAZUQI9a1U
XgXJkRxtCbHTjITscV4DjDIJmWlweiMZiQbP/obcAWVh9JHkFAO11lrOlqb4lU0MjsbzBEEb/I6n
OocHdrZsw2ZpPVIwcY7K7A38Rk9/1vMJ4U1Hj4Z+cS458Es/+X+liBfvL6abYvDC6LQFKLv8SLh0
0CWE3X+nbpz4qPQkMpEjcBwsAqEBOmhRamQzGlZFjAHgVHjKTC6+jCDFz8drTER1rizYM7yjtbBW
hmg470fqaAqEoSg3bPtp7nR09NiBZ4Q68w737soFoy+W4gKYiYbSPL19J8wj35ZJ1KXhYLSeCarH
5L5fdAsKQHlhR3d//zNgYAIdCXcN0MZsCPWOK98ADxdgyOWpFbAt4fQgsm69hFWwrC1a8BdQU5/C
XaqZLxpbQ+Kxn9ERw4DuvQmuK5iMmVNDab0bZtCbILkLcwnTpbgXD2SJq5q9XFRxsCvIBIVO9Xlp
fHgKoOu5MsaFHzhbk/3li9R9P8d6xkgww0eqWXQdGyXPp/2esbIrMxGyp3hfp2gXLCGr83hVr25V
YcMXAsKodvJwCrQcIABTSlFtqjk6plQAsQnkwJMqxikkJ49rXqK8MY9a8mzuEh//HZklSPK3t/IL
X0Ho8clj0VIJ9N6xOJBWwE4sMZhcO63J6v9s3l8arcg1a1p/9pz2On+lriq1N/vAmtg76gsLPDNg
XK7k6BoFDAKLRBurTBUTHdyP4c0+lBFADNY0+d8J61eDmUxOg7PgRr+Vrmb1kRdsX7nh5u1xuyT/
C3+LB/uoFV5mB88N0Ovn86W8yM/zA6VWcsovQP/irVQzXlTwptE8bmduuif0ROSG94B0k1IQAWOf
5BN/Xcs/g9ORQkf1ittzG/CSHQwfvFK3GCqRkBuHKyKWwurgMM/JwIoXSjdnO6o3kCiYfp31xYHP
50nBVVQ2Elkg3z0aZdnBqg5pvcGYpzMay8Mpxxb8ruTFHLhHaUecMWITutH8sUmL9w7i/1eDgtzy
JhiW4PGV0exu5auRD/pzGkcqNzqgbipdoZMGJA0T5aUDIUh8sgyB3WQbB4zG97CtZS8gAFMhYEbT
62QzFc74YUksxqqM3VEKTGsEkDq75UFgeGXe1UxCuDw2KzV1LOYxOUeZUN7Utt4jQIkacKVdkcmr
BzpFC1708imHHR8YlrU9UkkWBaOprONbfur2ZfzZAj5e8ZfzW9ppynfiysslTIee2FWdMtv7xjJF
axM7eBt65ID9Cc9spguevxt07e2JLjc4ZqW/YlmC6GCdNV8GVMz9tm9erwTwOBFQJCqxZNSibnmj
bVvwUx+pikdsu0gl04296psZejXoXJWVplfBzjb6shK/ntaERUZV5Ob8GCle4XLODZL9mMqVVfHM
fWTgQJ8FD4Railt9chISFAzGVB5vPv4ZMCyhbEoGJZOCbpSAJQ+NFVLZZyo+7kUo5zQXPkMlLqyI
DfeyetBCwFC8kfWGt7OEvCyKbUDsPPj6VWmX3x/ng8ZCPfQTLw04gLDfyAJFncGsQ4enf6MwGm6C
JCZT6Tf9YhCviyryeGv6bftVtZs8K7gxOhMA+aTVs47UXv2fellmiHJf3oBTU3+TsRdr1F5FmnQh
KBtpYkFsX2a9ZjMNpFVD2aDUxRq5qwS6GKMtPliNe4XnWND2KpsakYkbpRq9FMlzimmWfkkLNNuy
pUViuwtMA0ZbZWrYOwyD2g2UUxgW5EJS/30gpobUQNGLdQXavOAWfRSXXS9bhA1Fwif/vmLiav7a
HwPy/fVLSO3uPVYLIdxh5p6SjGozzcLLQzE/boG/hTueTYX25BcUyAb1TWEJ1+/B9awyE1aFXCvA
EWuEfViChU9w2jsS76b2QVb04dQkg2RODnXTlfEqDC9fWmx39EwCyE/RyiURYVgvQq2xabKNGB2B
bPPWOpMlLmE7XS0TTjAWzT+6wFm08HbyoK67BiPEd/0aIDkJx+S6PYErTvK9oRF2SVH2uS/MFYTa
xEVs8WzjpjB175nSkibaLxmsWaFmzxS5clMZCVTY+GmJzXAu9XEmMXNRED0hwP/Afq299eFAB18I
ZINRg8YXiAIpMYQ91IQITuaitWPk7jlrcIpgPq+o3X/+mrZIHVxNclqTKi1nR4OTvn0cRXa1Hn+S
moMe0eDs0baJe31HEkzkN357odYvc8+v1Is10RZ/Jiaw9xATmB7aejDrvHJctWAZ2QqDMDZRR8lJ
O9JftRWDtYiWfxTdB7j4FXhshp916Xq+0cHGzTS/Bg2BxFByDGNlBCGmfhTWdXdhMrLO0H92y3hw
gJPDgTyMDRJXmNRRxAJ650kA/EXfjeLOBbj74GYzNvdqnQHuhK/8XH5E89mhWhVuCfM/hb2G9Ohf
w1PIjE06UU3axlPpNtplY1YknHmaX8rF9BGlZsi+KG/iEMSsspbgj6VCygWnMU5PRx3nPiyrW8YV
JG8gW1I4BmmdNZ8l/QrC102R2G8DZlmelprKM1a1C4GhVQ6QWI7v+8NAOWHoXfbdt3L+9TQPXbiu
6/Gu1sYapr5PZ2K0jO55fdZmq9kk5+IE/u2w0q9oqgdcvdla3phaP6tr4ncSEykK9XO5xowklhDU
4ViIzJYaILVpsJ8Tu+VLOSkLq/vU1fjQ0WFYKaH1fsFtS0kKY/FcEAotEyU2weX3TXIxnF6PVH4L
E679mXTdCnQvIwvMLC3z3UKOa4ZwogPa1/Up7D1RnwqgilKrL+c1/vb2IWg3hk4GQ7gLP9SzcIqi
e7Y/IffKO9lfAAUhOQUfI7hf1NhBqn86aluPT5idyQ3fkWeV/hfMnIOuBQM0sSpTzu/lBoLV2Qmd
jssnDtYrXoqiXnn93qH0XmIY2UIL9HWV1fQKz2szePLyR43p142uVhznz9+UYcxI8/qpEouNQoFF
MF49sCdsD6HAlaWoF9fdSyun//CgVODxcuakVs94JWPXLWtEJlPBHyvXHKFky2KW0a50wzdqYE2Q
+EDoUQEoxZ1ZSzHk0mGrgb3LiVl3uUbu2Lzrtyg+bTBnT1JQN3Uyv6Ep2Y9edJRqZI1/gNjwqY6Z
1quZX8DNUcHVGNZyxqQUMvyD4sVQxbWvE93iGmiwKxl1MODIvTarj6XzXiljAjBdMucIwpwlUpV+
0ocDHUSxewqhOet07bLXx+voaSx27Z5S77giNhqGFjLnJmIBbLtw9RU9lVOPyORytERF5VcR21Ot
pG0xFFoqHRt+eLppec4qIwueA6XNHvqQ9U0UOVRxwbGes83g3Rm/NlBEyOJ3972JFHCi+Zk/+Jsa
lr52KozebvVesnHqipuYxuLIpQUlF2EiXW8tuIDFjm0VNmrNqJkKIYdplD8FgkLD0MRZnPA/NGHH
2S+aGAC1ONOtYdfsx93eXhOeUb++Vu6C6Y89+Diz+JEg/GpDf2rSuibsS4Pcz+cBwaKRe7DyMQpY
KVrTh5oHcZ/K4gjwNcVoZoyUc/NS+g3tm1LgfUZYZDImlXvZt9TbYMHjWArQg/KYrP5YkUVwlp/O
pFP35e4wLknMRqb6EU34zpsGimADTwnud8VxOQjH9rFofUmrULPQ2aKHcSkvF0yifuXmrtXGExDC
fjQKLLY6iMxlEGb3hH6pcomrt5l7gNxMzwmAGEOynKn86lz+BJGXp5X/okHvqJqXD+7MwMldoF7f
B1Ag35EuSwrSBa5VSWe7bprVU+E43V0lgrVV1KZVwOY/Lpn2V6RW/ACmcf/9HD2K2OVEde+mbDbL
Wh+dGBfkm5tX+gL6TCMdGND3OUYbPZGF4jK9uGZDciRo2oH4QYpSXwp/GOGMu986LqVvAEJjCVdd
/+OxO6khjkx5OfLpTCWDw2UDWQXpPcaZPDfcAaAjx/dhuY3OiSGoArFUHh85aI/TD81MP713z29X
q5sEHEbRQbyTjrjzxe3qHXylWZ1OHqp1ZSYpKfYVH72TRNRZv8eGx71OkmeOkXJJoR/TMhtqfMie
lN0haRnTl9WNxO6ZXpJ9ugI1+Zl2t9VCFuhGKMhkDC8wniUgYuCRwKnBnvs00RG8itEL3LxucGox
+tF4CBXD1AE6NP5zsa83KM/c+RZXg+82xzJSEtq8tDubtQ2VIvlKgzz0QOt6MDsdBCq2IlnvD8wT
kitY/pJvS7jdTvgA/F1nBcW/Efj2CRQopDEGySFmumFHL1HU2rZRjVI2orbmLt/BCqfhn4Vv4PO9
NQ/GPzhz3Xooc/OZmeXTcmqmikd+QYoPT3AZCUKr4kCVzXIyu5p7BMzEP1ENjC47Wj47zK8Ldl1B
sGDi9HyPEaHdFwEmS69OS2T7rgzKPLYEuLN8z46HIwknT+n0FrL4dH0/cydOQCLA2ioTHbyPSWTS
QA9QNnEoeKK4cA3LKrEDcaU0Csjmp7DEjBgkB2YtA/m7HwfLiJSqWhZWzs6QFnIlE+BFaux/KmUk
CflFPsFXmJxPNFvc8OMBI+pk7HONP+/y8GdcXG3MuOc7Bneip+qfCYcQExKJJVwa/Oy6k3zZxg39
bvFWm3eSts2udsE1K3rhecXt2CcBTmU+N+XnzrZ3Jtc/PoTPFq8nXvK3HJk8pE4x1oUii47v462C
Tu2iJbrJlpFypTbpa8VYANvKpajjh4VxOqOEpTTDu7sUErPgpzU/gsl948JYr/u3NxLDo4YiN3lB
3vUXjUks/HD8BpkzM+gOBzhr4M1IC0b/6MkRhUA1vBLH5nB7vK9PHMiM+HrzShziv5ocsQUHWcmM
7sZvuvhukR808PD48W0euk/wIyAttX7DFxGUsKU1tKiuOIW1OyBY1K5T5sEDs310cFHJLpmvOkz5
TTjtCctXz0DuGVJx3H1jyzJc+YvvA6wVwPqjOlPWw5iNVYdq0iIGDQWhs2jd0BWBIQ1y3THRitUo
FabL9AGktO7KgOzWLEIpvUiaf2hl7eYuxpxatKeZNagT48wMUtMDGQbftpFP2JN0d07ui9GiN+Qn
QsGLoIQXOPT0XxGYOKsRDJnvUtro1+vGsi874aiAzfkORO9+17QJ6Ew5UQvycjDOaIdktw80RhKd
Qy5XIYOUROTO6xry0SEkaVnokvCq++Ow/dQAaPBZh1tIgV6GOYgSM0Ea7f9f/n6hFj3vzsXyR0n9
3itB49P/PPcHOqefQ/f5Kpq92jcFtMZWbPb5bDa05RMI7DQrus1MRS1SGVn8sVqEpCV6dblcEJz/
GMQ0heejlQZM0nZMSPGBLhmxkuQZneL9i26PrA6OORYBkObMB+tGV64f3VgYuDgB7nHSClHQtCbH
pocypheTifiR9crCrvP0360NdKxgsWCthTZ9xMG6DB4kvsbPR3AIUayC7WTGSKcLfQWpwq2/6It7
bM+nxZtZmuag7aRSsEc4LE4DNaAz6lEotfRrfK9HE+CEUN9qWqczoS517BGMVet3MDUQa0Bsy8/a
X+7QByTo0pjC9kGCAc/mxJr4E9iNt1bQgHb9DkoUs7ZoSPW7DRzAA/xksLNe5XP16K7LOrcSf1x9
Vz+gwdvkQmfDXGKo9cd60MUb077rhYnjxJ9eUNhUd1TZ2E42i/p3y2/3qBy3geOXsebGBiVxrBE9
V4YKTe3ih2HD6sFAdolHpBzmd2l9QMe+8Mu+HWD+1WHzBO3oQZ4unwQ1WlDSkjVakG7O1orn9DNm
4Wn07JXwwaHSZrM/Gn+ZK1khXM0Pw+VYpnGLJL+2S7QicXEeyzu7+Fp6c30tUj1HkleoH2X6FqG7
EEhDK2EMXGq/jP1KmYYrSIx7bIBXdVzkMdRxkhcqyNAfCcBPKC7+1+P/S0tdPDHFo+YCBvrEzUnZ
Wju8+n9UePItF+onBpbKfS3wxOracfzNl+gzPTL2BI2/ZE1YAnsMh6pWnSUHwZRCOL/JlPqSEyuU
Gt4cvsj6pPfIwG/x8E/Ec5xLVpeha9FQZsgbVIuiNxEDmQqUEA4K1ODazNeYyxl6lPfKsygaVNQi
BsbTl9eE6fQvTGBq4iIwLBeo6b1Fb/OKoMQu6kVF3Mrtsbpb9lo4ga42lg4CHUDCbzLg6ho0v/B9
ooqCjD3Z8GtRO4YiXBTqRJO+Xz3UaKBA5buHFuNeS2CcoNikmfhrhcRwDG4lt6eqRHzWK6YnqAIi
YcXJTmauBcPbhI4QOoNt8mKkCNKp/oa9VIfiDeeHq8P9ipN3udWFvB1x09vEdFCwJxTEpqzQEjnU
wwadsiaLIWv8e0yA1A1e7P+GhVoLiMVip3k0MF9Zn4bmmCJ/N/Y9dCAYW1qx67NMOZQf0bjL6Aje
LldWziAY7/myohUrHX8HqtKLYdJ9DEFbspdUoBvKxPMHQyfXzxaWI0wGOvpfeViJAab9PL7cqZp7
7aoJd0iic2HD7I83/6oXdqoJmb5K02tyKa0mCFqXyKzP/iTCAC+DLYw3Zrw80AFlqSHY00ytnsq8
2yqXpqiWglqwXciQq2+dGxbdSl/jfZ6cQOznkngNRqLhwgevFcvQuT6RWzQDZTq3K5pjOB3PxNDD
kx6QfpvOvljMVA14BU1I0arfNXXGsU1TFustW9zcktnZsP2k/U+6Y0DcNjxGMmXVjbaAzjuDWAp2
ieUwvwUsSp7BaIiPGZFH/k9N1ry8pCnQKZAg36s+TOu4yVKtS9KplTnse3jLDgLgcbiZc6rFVcwA
iE+Hv9fy0h3eQ7yzYxT6YQR8sUJejR4ww3b4xXXvBkn1kmkTODi38GHUXD0XsbANrMeGiZDcERoL
vuoYb68azvZ0RFHGprvSvfMGeO5gxXsSIlEfiTYpXYDCnyfpJ4aenEjT8Uml+FJwPwLS9ynG4BWe
y1eC8Z09F8QPngeWRERuPkmOArsAn+5JULF48PR4Jh3ZQETEHj0w01yf3y6C0Fx8ataXLiqlLAKa
9dCE3ZBYM3piSHi0J4bbaFGYftemE16TKk372KWAbCNdtEMfaUakHjh+WpGTZnO3O2HhVVg8DkMR
ZmWDhwVoNIp0n/3xfnYYbpOMngsV+01D4isCgxrO1axzR5xsjJY/5V7OGeejpfCdGso9XpYg8AG9
hVInuzt2P7sZ/67Lw6uHOiT3zIS05ysCGQTqZlKnjmxWkFFen0uREmSKFgdl433t+ytdNr0D+6SI
rGSN9c4ozadm+p7PyA/XMmfBh4hu4qfGsalunK9fSXI/4ZhUOhhmF0U9csak+3qRDeFJ0qZdbxpL
bdh94vEsL9fTaPfNxTgN1ozmXDI1s07hd5rrD+VOJtOF9aYKYVEEFdsQu0Ta+hLb5hMZz4r+egDx
+Dlp5wNbeMIAQEVtJM21KtH1NkUxKT9dmbBEtmg6sitTxt1mrfxLkzDockEu2YbPqyTdcQklMfmB
xsxZ3ySoFv93p5EA47lX0us4DgH01P3Jh56X/e4cKxI1SekznqP0KALWrhgeKgCHYJWyRGGXspjn
MIQQ1lXP2Nl6UYN/OKIr01GCxB9GHzPrLCGrGIcui/sR2qyhlDratUHJjH6nNu0N1Bz4qgSGV9tY
ksE3MDsUQUopNetTj25CQx2P13SvYZiBwbSyGDRD0cVfdOP9/22mOwe14z35yS2yVdOIm5RLcgaE
TOnPYFMvE3zZIlMPv87r+7Y+aTBYGKxA2YvskTAT8P9pDTHDVuqgz17j6UrTXvTRlugC3DU1LQUY
HYiXU8BHh8aPP/0XBpMKX+Z4aSSpbLbsCL8jvLgykAjDE9zwgQhLyIXBZwCI1MtGM5+N5zyi8ZwY
2Crar759HXSD0Kt4tynZri1lmlxUwhzoPqeuw2unQ69RW6LUq33PQxYG1Nlo8Cnr8/6X0dUeybdO
MSbUp28FsEIr9Pmnr1gjRHNUir26Dku09tzbsiwcM+Hg2Charj8W+B1ujXSx2IuwOPSt8OLeWie8
NOGG/F/S3363xn2owOPvN056GKATy/G83XGImnswSmiO1yKzrUnogJX+zOULUDY9/uM9eJDi35y2
2iJGnOrYXbP48N8ZRld9lQDY4q7dRUQReFgUiXkXe9fXXlkYZiauT+U2UvUEVjbuKydA6m6hJbs6
HliQAp7Y1iqKZ1pviphuNoJ7uVYRR9Nlf62+GQEY5eqlRHin6nySDHdTA7PfTjRFw42AMm1+0HTB
3Wiepyj8CMpuKmzyIORHO6adDLtXNm6JBw6gFTUBSGzbzcNf9zyxPuws855/YC0c//b0ROjk/zwv
F0NPsAbjG7NSGjLLfbAa7WTxBHY4Rar/RmnxxkTG0tJRU05xt1/DBSa9ejj0SY3ZwpHMG/sxZm6b
Pusto3Cese3AANMOb50o042bdRP1BKdBLnfRRUcdyfa1dpq59EAyeZQF+hBl5aG/JV6X3gntP8St
xwYvOaE+qGWx6KZ3VRVuceI4ct+ss3pqKEFSPWg5MU8McVzwFmnQgaKyPd9/fRR9waXl1rsD7+vD
YkvLcWqzDz1E519avjrsL/ROdPDiCyabodEzs1KghO74rcvtL10MtCiMxg1rK9FPV5Pem6ietKp9
f586BMyA2s1sALgrDiBicz89LuRpctj+KYy+fB9cvkZuV2mfxo2CPncjoEh7kAJdpW/cRqiMtvKB
ihIBK/NnHrS+25FmwpJIpCuZXRHxCuPXIJBhwhLtitUf1q+jDC5tiYf/p+onIsDW6CPE+e3khLqz
F6Jl8xpJ5EliZn+9gR6+uUJraA/qK2agOil29ll0BTlNPfkvH1o9HHe/nEWMI4UP4JLQqXSQZ2Vg
KCQwr6p5G0vWSbX0H1FiTX/ftPIIw9iVpqQOfJnLrlcubyJW9ovDrsFoKag/biPBwnLM9eAJklEr
bxFHLQUhj+xhaSmZnPr+OYrwnM3SOWcFR8hXxMbKi7baVSsCzZE2+iHi/Ak/G3YAljXSrG+U+5HG
RweRn1PjmShfi9ACNwZvPElRR+6O2DWzgaUdN2H1+HM0ECTm6cdg2PHKS4/jV4rluvF7ftlnAMeI
jf9ecm9BgoxPoXc+f1RCtLKjHEw40MjxZrQoj6PFHYap71xQt5m1znlLpz/3YgbG6LjdfnvLeX4/
otSeodaupnWmt8jwxEigOnK7D2J0UOEx7phaqUpFiuUkRkwQWZn0dcIy6YuhCOpcvuakqsb0+wdu
NDylBm90NghqKZpkdR5RTfIyEv0MKJJbmOSZ+GP4UWYPuZ7i8BhP5RZ0woL/LIHyxPJB50Bb1S2h
H8/ei1gzdkHLcuGTAz1HmqlXgx7flXx2MS9tWCDNqQ2V59RTmHmyyww8xIqBEXqyD8/+7gNhAybP
DGjNppM8Jc7KBR96TPU47oB3obIW0fa5CO9zUwkouzLjORB4yp3VXwrFkkP0h968PAsKleCjRN1Y
afA6N3KzVtNy3lfhwFA17Dz41Q+nXrstpPDBzF25tpvTRq5TgN70hJQCDlfsUzOTRZ7WzxXDSld0
o3tYWUMD2Rm1uLBDnODieJ5+I9pF2TzIuUFYXMs1i21wcsVrvFTDB8mSN+vie2z60rjwyHScqrqv
SlaUSJ/h5+AVvhtQzNufqaKXKobh61ucoJqYDGvw3wOnBaVrDBPiS2GCFcDCyX4Dgbt1sBQNx/D5
0OGbD7ZyWOSNsXu+hTrrYRFeFiGgSLZmmGOSb/guAhRGfy7uBfWidhaawqlPsRdEiv6/6aeuwREx
Xnig7RW7FcIt+WBa0BQHbma+dSFjNLiazTuPGbGwggulumAEoxADPpejvdk0wGPBF/K3qz4iyU3A
6HqKpnDTM/Pom6/W3Tq/zI3rAn46GipVR0WuurYpqtgxG/VrgFIZFS9ZvjvotdNxu7vFn6aqgb6y
8I1+0gZd+U8HHiuWSZwRvUmG
`protect end_protected
