`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40880)
`protect data_block
hTX64IeLyHzfa3tJyS5DfnCGfI2VwUPJSF+Bc54ckFyLzlKrnMrf9iUqLKuw/4pRY87b2ekOsuOE
qglA73Febmp5FecPXQV0goMKpdlZvbCdxkh8JfZSeaBfKU3DOYCnmK86vMyHOJlF55chej0UWfs8
QEilXD7g3TgcUnP4AYikfBkFDtiSq2WQanGt40mKpyGHP+6z79WzDgE/pnJUz5W6E/Z6es1ClwcX
UT6WLW4ZYolURbm7Q5feJY7OCWXNWwsEjOT3hPhCwhL3gV8qvs98QHnLPIjLjlPc0NCQrSEFuezO
Zrioarn9X+HJHL7JK17hpnNa/q/q7tS+JJW3b3+Npv+GjTmcNXsCC8D2Nmy+IIef2YwLuMC9LQmB
Jbo5bxZ0RJYoOvmEaEKmkgdhlBmjrt6zbFmKGizdRWmx1OTJSP1w7N26Y7dmM1B8h2bqyiN9Bx+G
KktAeD3c8hFCTHYhp2c5oSILjBy8ZC5lPCTFWn+TGJJER7wCHwQkNbOQeRe/A8C79M+WtiHY05Pt
faKeT/flB0FpA7gSM/rdcAS1DZ+zDRl5JOq1WpyTeQ+X5eac2hPkpbFjLarbqlW5cgDbTuHR360T
uH98ea8+A41j/oLHFMGIuM1IdFRRIY5PTZMbfZ4FanR940uJ2FyWZAS72HSkbLV8rL/AXYvYMKV6
bAjvH97bZJvbHJPLbiAGOmmM9Q8SHYyOBPE5uulzgryPydarZx/MvlE7lhfzGXV6IxCXf0bUzC4Q
QfhSeVVqVw/h3lUbP973E+M7TfW2ZG1bAXUgqlv26kQ1GZVbL1XyL5MoMC2aNzGdvN5NmQIgfo3Q
3TfUkP8gl5ZM2/58JF+2bCPEeBM81hCkpIP37xj0AFPpWXrJ7WFJMV6wVfVyE7tWAozNtnNazqk9
e0EOVZBCKJ4VET5a/K0PAY6LjyGQHWbTtKs3xcNRcct4wvJfaCAXub3fRDHHcfQOtmG+fr7SWkcp
NQapySevFTS1Czyj+oOlCKs/WeERDSlQUd5+m+POK5wLGX1vOyf99d0HgwESievFtCtMHSIr8OUR
Z3T8lH+1872mjN4q7Jt20fq26i6iQAeeCMrvL8gjtJkj7WAwL/znyaosbr7aPajs50TNHkDcEKLY
xtUJbQsf5cOcnOIUxI+0w1hWnnJHTh3ao7Yxevajjg+yAoaB0oj/RGX1nbB3G/poouuzV5Sp36dT
SAihHcB7cdjW20bscxv13+F2z9UqMKYvBctFIsqWJXmQNd9vp2QoXJB1ZT9WzDAJpbhdmOAebfOm
OVksObU/uptA+v5KcAxC992HH6mQfHrXb7aeoHHtxLeoUrI5VDe8/xDBXM91sygtZhizUtuKV3Hl
5qBcJxr3DaqsJFBL4R+w8no5+alt6E2/WK3dslEHr+XwkZu7yHhhi/bweHVQEevD1p6QFppSVWi/
sMCPuhnwnS7L6kCV/XgdinsRdY9hY6/KEZCrTFydrJtVckpPX3c/CvnOkSi39XRqV5wiLNBH1vuv
GNVsMs7OohtZlxqZb4n/RRs13DArMKJOkJxx3tjCv0iqtVL/5anlyoKyzP+plyROqmrwZpQbh9Bj
qG5r3WeSsUOtNk0TzerpEhI8BomS2JcO/Z9iQb0YuUzBxCuLW3TTmZ88kCsLtdlkogtWUAXd8TOi
OOx2R4sQTemlX0bSsSYFzBkIm38rGRIF+W9n894wcPBqbpvbzTZ2ln/JBq/UFSqOuYLB4Gt6QvlI
IiGSJgce7YmImM0aARb2Nc5HXBF5lY55LS2zBWEKwPfjjOAvqyy2ZHoxCVDxATnsJU8mqNP1/+W4
p1myaILY4iMVDBVx3gW2eA0TLApCFpSeZMUg47yQjTvQn8/2mefipPpsiTbPmel8jBGGK53CJ5N+
UxP/Y9xdQHVoKFLxCsgvGV3+fpfWmD6B/Bi1GHQQCEyo/MeIk5+h+3I+YN0RkWXwUkjdQIbTDDBR
gTCsfZcYIK27xf5XoTVRiVJ/xneSeHWoQ1oMyb4zT9kUV2OJoR8yCKhl39jY8TXmbt+NdVtUhaRs
lv5UbL5QHbkh9l4bsdUc5/HyDrUJE0/LQTBlP9t7xrgrJvYeo8C1x2jLpYli6b4fzMw7AJG/XGwS
cQsx5QsT2GzspT2QZgljQf0XP1K63lNruOsc0GwVtJzbDi1euPPsPuPRzxPhkmsvreStUSBH3syW
2RRHBygEgoMwKDpO9y4czyVyaNkObyEdULRrTFeZfVmgBDdqZhFjvaLd1cv3YlaImH0vqu6alHzF
Ex9LKEaVUbpTCcWM2k6b7FW055XLiid//kMosYUqL4BBN3+BwER8CbQxZEZcS0+jCZsXAlewgyFX
vrfJYXfC6BZ0jjDcNMkcPnHvQcOWdjbYK+UEnwXlpjJ64bn/ixzUnI66Lgmrvx++bt/ned2xFIks
BaiXXDsoumIJiBo9ItXCxT1AVfc3PSdddJaICl7TQMJhVUUuNIXP2T47ERQjBYnGIE6yHxFuA0IN
tNrG9McGIxv9nqCDSQgx1Gtex050cl3HSNohgYOwsi3S4epLx1UTNBcLRJRPcswtgpLQG1rq9JS5
vbMD7bP8pxCHs/sOL2+P0b5pnsocJyQ/YkewbS6zSrWPqs6OhJqMqVWztZN1GY99o3lM/OM1wziw
Ztdp48XbCt5KfEeq1SL/MB2f54IVKByEfb+dbFtVNczbxaFRV1EE7vH4RBPeP7ElYUexhWvBbhuN
2M3wTzHIfisQhVb3rDE1PXTxfTByzqgIzvmDdTTTF+9Rb2B6nNtF6/aiTSRBjt8r1G3x+m9SOMHF
dDNLIjJm2VRu82OFmHbikttWAICrktntXnndweu5cDRtA5qH3JO25UPBWA/Rr94Jr9nv7zu720ym
f5poRim+wMt+6U1FDtpg63u4HYa08pwwPzdgitGz4g2+qbg5zc9nxu/ELYkYyKxJjIPpkNe/roQD
Gzwc1fTbxzI3wE79jSJhxB9/gZHob+fPrQzKx5WiO4f3BD20oyvzvYKWR22zvXNFbx9Vww0w2nI5
lLX0kUoSIR95y+BoGvhCr2JaOdI44FaCgFgDgnrJVg2/3rbWS8cX5dxP8EKhFqb7D2U1J4hvuiAr
rbUtiP9xrf9BM/fmBd37BbRMT1A9QDaWA3+kkfO3/p+5AL2QG8IQRbHIUMMcBkjisGFlybtTtP9h
L0YRqFnEUc3vDfs02wO2/8q56qwRsCNqoL7WGFgm2QEWTkbmdaCaApBKVDygiL98KDbEA1AtDcsv
FKcP4OTOJekdqHMtrZjw5JapvCJjVyEDhWdmzoKj5ZuxlAc7jvXsgri23X2LW4Z8tPsUukQqIvDH
dcM1ycgMN8ydHl7TDyDAmC6o41dY+4eZ0uaXOBULOftkG91RI81C3f7I77Hlu3U1+6yc+UgP/JUV
gxbO1hYHWplEHaM7piRm7JSpmMqETTV5MJF5iQqz6kXDfaRMlk3fpsEb7C9rx8HohXf250Z91UMT
6+JK5CUYKSN50wC7Ar56H4q0hOxlmBgdjNpoxm2XetMUlQfNOtvee03vgNp5sIt7LBwqGGAHFAa5
wgPFoDUp7kiOc0eArmwKU9lHt8M9blAjQPPZY1Tl0uZ9EkxBkF+IZbBp7yd+v6Ck+IZQzWrvr9jY
qke+pVUXojhdqcBHQLg6JhdG5Ey58oCAv2nkpW1Fcp8fck/GOnCnVffAOzlh0vLnIVkl0CT06shP
aoSWpmSdAxgfx3ua9Dcjhk4BbmMUtbrNAGlxi5OGIuMFje548WYvUX3frtH2FaB57KcLDj54gAe6
eouAButANGrbU9cC1N2ukg6J/1+JSngNZMYLkxk+T8c8b26keuLZNSvvJ0Iw+87GGtmPto6pWqO1
oim6fcroD5Q4sqfsCvXS7s0iwx/Fo9QfrtZXT2CgzMTlZcExTwp9IWWWUnbK277CfFUc5esl1oKO
lWfwEALtaRV0ErOpAldQ3aCZOfDfqtFirU6QJI3AeYGHLc85ou08EUXOFj5P88lqz5x9e2Q9Nzm7
lXMm5uLQSxEV0Zv5iAV9CZM+o/c7Yu+5XBpzy+YZIoCBmHLIxAKFjc/S83+vrXrRVgIvrzfqfDBi
OezzusbFdvyHwYptzkfjjk5eLbB4//3iguo1nIkYmGnhrjJlEGnpToZDGt/SGVB0cPAmtKlFwTtn
nNitkB/aQFxirY7B2/OHj4RjF7jgi+czuGgXlBopNznIIwt3gUaAMosSHPvGCc0U4K4G+3WXfJrT
sDMDrjkN2uwA7N+EaqMijLQOZN7GBVn3HGZA/pnkmH1TLacvRfyCzZZ16nceSf33OHET1XGqKoAh
FIiG+crSGvYRJiGoCQZ80ENM1VQvxWR7nJL4dbZSP4PBn8arS0FAndbzyq88myXIZichPNXJOJQh
PShrnWCDKrbGZDk2SOKu6yJpDZgEP80wbpmxA/u1RqobUbjkEEr6+cBZvt1J+oMiV/n6+8j1ZuZP
p7B3T5o8tBSvIpmv8sbafUekgez1aESmHGImvPVvbi84uiBZBbvq3C9PHfNV/dHonZd7esNYGhBr
7vJ2lkbGhE8xZBXPXqAskGjbjdO8GWbsHZKe2tV4YoHXwrtA2a2UdyAjHpM4QMGRiqsWCBLebIpj
V+PWxY2A/aoYvDX6mBSaRA2oLyg3SYoucAit0NizHxbahk0tBjFoaMOz81hc9/xG0Bxp6bkdvHmN
FHlHQmC5UyMBqDyph6dPy1x3oOJeHKvM1w5l+a4YjLki81SZ5OwJF24k5RBikECyflassam26g7R
mcDqPWC8DqbKahvOoQYMHGLnVjsSjFhYTGYSnennIHGzsSADX36D2Zh9CfZWA3xu6rg2bl0VHDrz
YhHb3rrtuCZZOhrPbeGKutg2u5jZTGNNTpCE8FwG+G1sIUzGLK30+x0/gpxs3O1DWFBoVVo6PiPd
W/ivMX6r9oVjssLTlZQQOMxEc9tXVXOxZFdQHUqQfuSJ0GzdrEiSMd+bqJSiO3fuhk6f+VG2NNik
sypvjca618X3qZX5ev95OXGhpulTOy+4QN/4Gkm5dK3bSUp6psZMvCElRpscsN4sKrIKJkuLeMqv
gJnsvWwAP3vt/PJ2ViLLCE8iuId9nesCNNaauE6o/WIi28WKrhg0qRCj8C8BXiMfY/Xb+7gFXfy5
A6MesNmpwNlyAVpjjO79gQZYtZ4QwUsZr1xU0SkawGQesLrS4mApLmDrY2u9gZAEkwRowlkzLUI4
HVNUQUVAmcsiWQnc0zrIAxiPyVQGfcpUeRK8mEOiVZA+tHs0vtYEgSQ39zjlCtfeqLoF9UXekzlh
n+PDoDnZe1CqyoRK+rMRWIgKdXHEFXzmEyAoApAls3qhtKuDih913dDl783PLZbP4ZuFlCcaZNzV
RaNuOhJB29J5WA5BOY4aJDN4dON+UisY6MbNLMdfa05aD+1+5/9sqUfHKf6XZMUvvplUtPENV6SS
S+4cIdJzbme3E/IoWPGc2UobXGjqzLLXt53Sy4qc3siZrJKhlOO7FYFZs9/gTS797tvlLTrdqmhQ
uLtrAGkYlYNiUr6i6LhpVMFLotULzNCp8pWqXZ03/JQw+mTWsgCLp0mptWuRORGksmQdF7RROxl1
au0SA/mf1AX6LYLCN8/LfCflbft+ttnD/fTGCOJtt3xpwW3gYVBuIdD0DNKwTXZ6bFKJhPrQAAmQ
S1X3d9u4Fff6YHwzbap8HWX7dp7DeL/LZsXHILIPnYJKzrxSyYfwmMH8OamaxGuwt+49dBzBKdKQ
8uEaOkgP1xOB8EJniNmyEOUhIVSnEd3MrgvV0k6ADaF+yYBSp6JIdo/XMmabMM8hzCGT9mmfX6MG
9efTWzR2JIrhp9ft4xswQhQcvRetN4UBOQISNEScycCqhigH6NG2f7I3zs0R7ArxKEt9rZgvIQYw
fk228U5a52H++sqCLW17VPrbKe8CisQLVGIx+5kLuO7ZTV8Maekd5vtfeLNDXetP+u+N543r/DJW
qKNW1c2uFlZKxMySrJ45Nc4PZKYbY3o8rGX/tS1QOqIXoNc+DSoXa8+UsXWXhvWOgnv6k5jSDWe0
4IpsU668q/PFP/VYL005AaLh8FfQnChf0OcDDgY1ZXzuupXRfo/0Db2JcTjExcSMgnmKIJV+osSL
PrApL0IqGjHUnNtDGk5xgpl1Q6ZFhkWKyrYtG3jF86Iv7LVtLxX5M37w9YNAIuLJuRjZqKlpDG5R
InEHwlT8/1z+ahiElhmmgm+LIfJbieWcEeU+OsFdETqrBPYvJV6Xtzo7fon5DcZBX9CpNngvCFTu
dH64c4qNEae17wbEBFceRrCJPPukYUqQaL/uoqNmiUsymrmLGGNwYIMZlN63Y1vSNDGYBtG37Unt
LMchjgnEVMu5IFQbyb4dkr8woFBORLDw9iyVT0zjmxjWRchVegyF9FZAtkvaScSPAVZEgP42t02Y
Gq8M2Qk+3k1S7Jl4S7U1GtOxYNtM/Oc4xKfDfRTMZC1DdBlUxUIHOJjgW0zWz6KpmNKVuu5Qjk13
4MjCTkhBhYWSzt8ewoJavhN7uYQJ0zxVVyUQWMAzzdbjK5rHL2bPJCgGf7n0NemlDoJ9VauxhF/O
LwwT4LQ1JuaWbziuv1fGErN3U0EPrzRLBVg7hSqi0xL/4oKR1Qe9H4c5BONTP/dtTG+40SKJaAW+
mozY6SqqFzZEygvZb4LSOkGAMseSBwrXrBGIVA607nrSKfQqtcPhFzjcbLHJ1y7PSQxuasMj2fbK
DOyDS5OHv8sBYqE7vjD2mxgjwuJ8KwFCkRTSlx51+lJhOch2w+xE9oFTSAJJZqR0x3KlUSGtX0SR
0lPXeWduRnopsrXf4HeIQonIMEdJ3/Oxh/EHR3f84gDafgI22L07VP9MG4VlQ1gPR+1JsoD3EVmJ
GSIBv2DZaVY7ba3vgsVM02zsyskxbtugaXkXJlYJx80dHA+n4k/R93CYuel/F784RdexZsnitnEz
ZEBUkCg0K6f6OXwxqKY/ZNY/dnUdg9LSIv2zTF/GASEaQaTUG9VeEQ4BBSmdAHlfhr7LL+DUo220
LUiZuNjBhIh4xeD8oMtK0tMpTJe/CmbLd9yjMY66oIxNW/GdFP7iCRzE1shd65yFmpCEYwdd5a3S
TiS+MWSBWgi62mRl+lArGNBX0aU4xahNuvU8qP+0YBxhy9NEmhyRgKzBRppb09KGBbeLohbcaIpb
Fnvx6thOlqnJCXiv6aNEBIkkzEMFqA5bVuL5Zxw2hyIFKm60D7/24R3BJLqq6b75wXH2jii8S4QJ
+r72MvEh1AKAKOl80DwPoNes3UpiFs+n68nhmbKf1g7WunutV+Ux1VzsHgyOnQ+KQTvMKxi3pn4D
4ushWTDz4o6DK/PwoXhGTW+n9faf+3QHQgiTnoeJXv/gr8feamXZxRtcyHto6mpolSEV7DdIWnhB
LoEFwa+oMWWoNmim/GwtzALb7DrxcxKP0W//RapoklSwfROUDb5KF9O+CpJ7f+H3BKJXxYHMEdgd
qieYZk4R9J5IQVWdkL6gv2FzL0eik87gATG0T1HaatJHL35/D/V1vfFH08IVDwY3wXpLyX/NsBFi
L/cGX2vb2VD+SVwOiLZD7Y5u2K4H3RhCeDO/i6wpg1/3d0FD9oJ2iZIlOFnp5QaM+fDTqg/UrhCO
un/YTahwKwBnMNJSPGPyLfM5dJ356/YcFdhSQl7fap/F4DYGgFoON82ljaO5OfAmWv0ZwDi1c+kf
rumg/xtNPIsA4Z2X384Hhb/3L9JGK8KO+wnIqrdwItyzu5zPl9UusurfiwpVun+frixKH7jI9Hem
TquvvcAyg6YVurQ/rDjSP23RtEHof1ic5wYzakIKxEk3ShpByR09+nx9dXbJFjfbsNB9jDK+Tnj/
AHuH5fu25sxe51yf6Bnk35le9UFTKHPNp94kWxrDCUawaXeluhPLqX7MlsgsNzfoJraIakOCdfAV
8f80o7pBAd5SzcfwRaFWrmQIAKEAxIo8aa3MvIO0WR455wgn6rWlEtFRJPsyATWeTH7C/8xKMzow
iL4iXePTMM0iIoSiT+H+sx3GGCaoAkQUKn0rX5JCKQCqeMVka0HTI1oEjEoXF4GB5TAbv564Y7Dk
GRRI8ubjdk11vY2M4kJZuKnoeH+wIeDKiw/4EWOwo6rg2HOZJUexdFokRF0GEvAnBI7PyuQhgtAu
MoZ1jzd1z/vJiH5pCseJTns1TiZ5KXmcWVcCisaoKOY6FeW58lXiP/kzV4DPsuEkIFgX5EuXI+vj
4NoxwD1T+ab9wsE7WrDIJvbRdGEDd8W/jKONafAsmf1bpM2yGADLFwT09GYaXjapk5QkeWhQC957
HvslC3tIhZ+5Bwq2tOi6CB/9Nei3SUfx8aPP45jrCoRrw4FzAjyDSmzFJsThMOboDY+etH1K/Zcw
OjM010nD4g7FEkOi29faXtDGFLY2kzegzdinTrm471Z9QkwVOuctPg+NJL+HnyGXMCae854gOGZW
al6Mgo/B/+VSfgABH9dROq6W12Jgo0XLL2i1VSLCB0on3/JM27Nl9KcOS66vB4oQWE2Gv9GP9F/z
2JbkIVGyf9HStYtAdFGEuxCmM/3BtVlIUYEMkIPETlXu+18ypG9w+WDrDc7O6gLRi9/0LgDhkz+y
RoliIFN6xTn8IFpU0m2n/+iOO6tgEX9OOsBR48qsBLzLo9YfldOmkIlFaPWb6ejTC9+OXL8khkSK
fDg0T9nkWF1EZNRRbehXGn8kT68vuNJ207km5dYxbT96/g+qM2LOr5/daU8y/CYIKSoyf6Leh819
Spg3dAH0UhPuuveEupfG+uAITOAfmFqzgJ+921vc5hlPVjDgwDC58J0BewmVBwr4tO6gFl9LzmDn
BIdcMe5u3PrBZWz/JedMuA7QUp008KoKairWDT6Te31PpojRab4UEZMAwMOIB4vq3+cpMYBgsxGL
CZ9rIzXoixzpYm7tcH4K49EBuNOG2fEGWC3w7bNoTze+s17L+PrVcnAle5Lu8tCqIGUwEY01vCcD
fYYW2RoL3mB07DQMivgWckQMB7+nhGmCWdb32RDquGHDq3v03OMctr5hmZJ0E0csBlH//AVJUD1y
9Sf2WpFlrOMWp8vmcveYoyPTHTI7wPXRhEiSUcy6jf/CWeyfcFmvHKSYmxVKHH84g5EloDQFNH6G
N9oq1G2jelzHMoeew5D+tyEhye6oP5oNvi8bFNPtFrLFWWwkV0jx0kHLUfcs2rj064r2ourS0P9q
yPeGD+5BknLB92IsfPpmpBdAD3C7fHuvIFWKuLmwnz9everzreptP819nz+Vfbh7SLk0vWoAuQy+
MO+lUD+Nu+BgiCcG2w/49ODDznAfHZwvLvWorSTmS5bF8a7DgLsZHzriUl+LOj5sLG17m1GLI9xN
rKViIipRzAu7mFTHdo5rq6A9CLNfnDvQBBn00OsoOUA6wDJ1lu5vULG/LK20sP+f+70IrrsC+DIL
CW6W1GaSIn/Xsa3AmP3LWuwYw73/PJDgrw8djzc3GFIsLkUFAMnAYT4YVPex/+yw5k2ENjwd4MKY
KsYMeFuViUP30LdlrsrF6995gTm+qoYX4DOLKstt9K6IbyygwX8LQoM47J1L456/3ittDvYjJO0Y
pm4l7QEp1U9B7Ch6RG1MX2wfcBX5hhwWfTx4utL3Uxu5ucsQdPXchRvJb6x9qPWnSmMIfUnIHrvz
sYw7YZJM9czZwnV5T2M/mD92Nb6v7u9UP7EmsPMO0YTGeXtFDJ1+h15kXZYTxc/ZCMgoXYV/SVqv
sNJ8y9Lpj5mE8LHo2wdIlokajW9Aer/VKbZ8A8hZh9Lwhyp5JBeAFMbTzDM1kkPcNF941sQTIx48
1cFNhcEzY9OWR5E40SvuQSfx1B9r0f4ryhOvvoCeKC81zi+oJtPrrMpcOoIVGJ9sP0iyBQ5vfVR/
havNl7vkBDW+2/YrairDiEQWIjQKeCzvZKvywIhnS4vN2ZAX34zV9WGvnYVaiti8D8/9c66Nd/J4
RXpz1+5PE8MijvEgzdRLNWbzZ6Lni3Co5bAoxb3gKlqJlJjZjoKXNEC3U1bDC4dux705xmq+Os+B
BMaCEAWumcIrMagWolHXKKaZ7Ud54tw6sCT5oeEb67bOpxTfcjQ0rxb7J9JSV7uyufz+XVeD4YCL
sd2A05jNbVcDyO3Cm5anz+NvkhEAb390LVCqEx96aUXm19+HLxPSmQ6qtyP5/Iwi5nEQ5neCp57N
lim8bZYZlhN7Ef+DM++NEFqP0NJ2kg/9/GBWLOCjjcylW2pa1+oeu8jIafHsL70tHTKmN2WrOXcQ
IV8S+8jh9/5I7V0sB2Xg2FDNb5wwNpl1Ig0JqukPk/kjEMhBObTATQNFBvJ4PpuT1lJDTRHjZ4rx
jQ6sQk5uJzOUih9P5I2R2eSZDLHzlGfAxqobldqtHqyG2Ry+dzH1AIcYmV2/7dI+Sr+geAes+jKJ
TN67A/5WUsE5v9ZJ/5sQMOBwA++4X73EVyxZb9Yqn+UcDIiUYZv36RbnCwf9zJxiSt3Ili7Y4oht
YU7/WCDMA7uHiSZlda7xeT0k9UMDXjYfzE20Jp+fNofQF81WWV12tugKmHEpWGSQv381b/UgR5/r
GSvfoSlkKvr9YFE2Ygf2GhO54t9VIYqOK9hqmx/cjpFmI+hDU4e1G+JC+Kxi8/i9f2XiJr1yhj8o
a+Xbt61kWCmej/OU9NwPE0au6fgGwS0n8MNLXQ4CCX1vBcCxMpQBiIgadAsb4uRkoHR+BelrHMZ4
gfJCi2ZMAjouXJ+cnmmHLWLNeMa4mdQ24WcQRTWLj0NSXbSDf2nbyHDNh+zfF2IRKnsz7+lqTMG0
m4ldJ1PYmiF7imw/1zclZsBgJm8duiy3MhrZ+shBKbhFjkfCMlRO8lkMk1j1qUKf3Ca4VSD+h4Lj
VxaoQuzguQTf4w6sPl4qK8EPeP+WIi4AJgBpUHcnot+vrxbY3AEvSzSHXtt7lHEFCSNsq159TwXj
q4fn51of78mnrkshbAXiUA90cjPPfmHZm18b5vAkw5fNa4H3cZM8HC0E8o0iUTA3YTQ+Q9fluyXQ
Yv38YHfmg9jHh86UvIkKqsiToDJsBFZBzQCx6lywdjyUOiU8wyrYqTwYzdNixaXvmlcptvYJvclq
4sv8n7ty9OpE1VCgetAjrRYfP4QxCtVi9ZTeZbJd0mUD+BWGH7zhR6vw3hSSsLZswgmk/9KSlUB6
xuMR/MlAXviySI9l+9px5LjfQmjRH3tXm2/GzuqAmx8XrJmc0vFB+/VdYqv7EAEYEV5pZbV17XNE
+gev9nIx+39Rn0/7IpKkShqtWd8Z1AZHBzyPVEGEzzo23D8MAYDO5mBZd/xJAwK0zKtx2tg+PCIJ
gHh/14lBEAoe5v5TnIBnOo2QUpaOypxpOg3P9cKVGbPnjHXXcoLWS8ukZ2WRn9hPb3OzrnIaWDWN
Ow60qQ1xk0gGDHwKD5AQK0S0XOByYW7JMQflap1hEkX6CFxABvzD0NokFuubEOhB1JajFrmFIH8T
HNqyUp4s+Fv1iqD5u2eO+3V9YMqVt/XMzv8pHoSKSYp3aWJGAEQy628tMa6kCqNiOntTO7Gw8+sa
r2berlWT/iBzjjPFq5hC9aGWy7Fwz61EoU0DV2Q7hM5R5FEI20ajBFKOZHy8n/8FSJ2ZHtSwMRm2
dgxdmpo2HGdcRhnjxqQeUfYj+rC4zUDDL8vA+sg/jnXSziC4JTEfjqjd/6aaqapoIFfX09rKkDQq
IQ5OY/5aQdG5lJ/HiVn/X3a2UwXEcQkHmmKKOb3Eqf/vbgfHo220X21aEIQtbBVa0YSZYf1MquMf
uQotgDeHOH5z8EgMi+ZrlohXC76cUkcVyaphhVnsLtnT9rdjS7RDd3loRsPbNlJUbMXSOiEk2hzH
skjBPT6FBMNBBA/8fJL25vKcuXYstfY8/06qJkP0Aun3DSpvu87FLEDyiaGRAYnF0fuZ8F4gZeHN
z9Ue0ZAGZnvZD7+MI9zkJqSnSaOCsPVPluWJ4BqK/YxJVd5sJz0n2ktiiEkOy9zojYcX2/DP5cUF
NOGIuq9eA1URbTkjnPxeQBIEpuU5LEPt+gzUTc9eo5J2I9/6Nw6lsPjuFMYtyUpYmNvpF0oTYEvV
XCJXjwMoHWowG50KXeuhkpPSJqN6D54UM2SLyksDxyZas/JItNTYG6snyFJt6KZ0NuC1923PWLSI
+baJ2wV5afeDCC5X7f9QEzbQzG5dyFvLvMVsms0trNbMxVbvDq3tRzAtBQxfapYCA1cEJy40BvZi
zwiepdt0PXOEuf5UahxHAoFa+06muxd0LnCrL5oEO2oDuT4AhA0Es6n6bqtva6Aj2fW5RGpsnx+r
f6+sra7BAA0Zs5GqZuHNkXiWdV1O/WTgOFKXdUSK93O8sIWZT8/ZWXGrt8ps199x7doG/X6nhPwX
ledCFUZlPFBJ1bTAge9i8OhHaUHVtqWFbVEvM21pxUlOOTo2MOkooU9s1+nELng2hoTJEpAd3H2u
BsicWvDCf29ZSler57sY2wT/kqo3Bxe0quzOmFxPbDzbE3yNvE1UlSVMdbXdZUnuqCF/eP6DizOZ
4scwBvZqHUpav/PJsfJKBTE9vIiJjiede0iNvqPemYj0LGAxyvXJzescB7+WDv2DfygIfbFxGa7Q
19RKFsKEdtDQ1f3QEAbu5AJ6kEtgkQzGT2jKHS7ilS5QLZNnkG+wQ/fYuBk9JnFItnkdzAlLCVMZ
Kyrbpb1QtD2urZ2hS1FJhJiiWtaHNb1CO+tyN88qno+Yf7WaOJcKui+QSZZCZoP7yDBl023Qs5V3
wQDfBJGsrwkMzn++YXQ5DQMnUZZCFndY0vBVa6k988hzjQDbhFbejyZm2cehwCnDwhmI0t0cBaK5
hqz3SsRDT8MRt+7puLdrVFrZif+ywFrncwF08nykRMp/o+f3+izHVjYLBBY7MaHRtBg7fJPLqe+6
TLx7HtHenqLIiBxl/gOhJ4EijjOoq5gBhu60uqC1FcVzQm+/7JIY3zbDCPUJ1CD2QXoWr4Mcf4so
igZStc69BsO6x/FRk81OsqfqngVmLpw0jZUNyMfmvKhIjUMELdhFY3cR65WFqR3lYE7ze8n0JRn9
kMPgekv9Xxa6+KKrivfhyJ5f6Jl++i3y0ntCjyha2aSptPIyXFtBs2VpVFzU6IG3EZb/XxLFUFq+
VgQJxtF0szeqAFvcmFpSTak9hd+3bWRaVY4QXyZLX+qGrpdGPzqaQJEyTLxVpD+TDfOYBL6Ih15f
qv7Tkl2Vb9UL035dFbi/bnFqyUqFfaac1hxZ3EY0eZNt/qkO2HXLVuACvSglcDjlUI1RBlqDPdgJ
6eh9frG6mSRqn0VEq+LeSbTc6fCa9TiK9wLR6vu+kOBy/wMFvSsJn6n9a/0CKr0cVtBFVVwsCgtk
//w3gN1T0DzOVT7tahwSuHzLcWmwGJAPbTaDfQUgFOqPhTYjQhaEra+XSwZk7qYJYgmGZNflS+mT
Bp3coChQAL4P0NkU6bAuSNROHIqtb3clL++b5pc46I5OV49ktjqKKkU5uKc87G8at1Ebq/4MUYkI
8NTeI4au7s83DeQfiLlI1wLlhVO6w+WZy/clzWyFCBnsyD55kETLygoQ3edmPLLpKGRJd3aekXsy
acO/2/LroSF2ugDWLguIeyO6E6oWMGp0RDqvjNxrTcdxB+ZdmzaZtHPH6S4oGUBEK+pqNIReyatn
Xd3IkU6HynjS7D4JHZJ46CXAD/5D+ue4axl/o3ZnUP+0LyQBxxZT2xjmxFA7KY5o+u8iSbkdTSGc
k87eaaDZ0aERhitYCWHwLPDY3rD/qf5VoT6cg5uqRr5YLc3pfff3EkLNnmvLL9hv/FXrEgmSqNyV
7PpeKdkzZLInM8jlJQBMuUJBbY0qN5TPlerJ8B4qhFmh4ErFlKZogK+uVOkU+UZ76JlICed3Vy8U
rzqUF+zvKqtez9NG99uUWuy6xA9vutWAP2lwNWAmG7SUmAS7Nuu5W1OCM7m7HYDipthfk8vQhII1
Rts5MpBP4gDGTxvK3jTQmTUp5qeiKtZgXDZiDmJDYMEPDaIliO52BOzg852oxigIy7B3KhsZtUr/
ODQe486YHVUzBve+1luglvEwSFXikKN4yQ+lwJW/C3AUJK6wuxK6a3R6TI/Er5pNyzjMfF2u7OZA
h5RKoJrDTwavYvGYW83aQn2S8CR0HDAGUTrBg3e8H16DUNjbV8R58++1I2xasUZrMNIQ6cB10qck
qX/k8hmv7FX0sWpHxRp3w7SnjQy3sfZ3YdTpJyFaFWWkqH/cGdKTrTeYt9AGCz92WPT2epxl/MRP
4/P0YeThkVwaeSRgo98ZgSrxr5Na7PxE0bNHMly2SpG40CysU3cTmN8cVNx23Fg7vOu/bncFxwa+
l7Ux1WX2pPHKKW2cittxDPvqbu+X5zGPIwVQzTpJoU0NbWMnFjy9avGzEDq83d/fYtWGgiaEA3NN
ICU09JOpNAUXLqHcqWfJ7LE+hb2Qj/FmztncZf0u4Ea2QRvFSRYnAkz0KBmTm8GC1/YykF22vV3m
Oz5/hrw03fv2cyZ3rgRQt9Csi/clTCciTQeFO+un+BMMkILcaXUNEuq8KDZbaVRslA9oWJ5V/peO
5um+mxYDV2I6S5xpAHYkFXW6ZfGSpx3L37IqLyrui4eG2wu42VPytPseJUnMkSPo4wx2LnedXTmM
4R1ryA+rAqaldNCeJs7fNdw5RIoQnXWeP6pvCOIw6cO3GxJM2REOMf7WNF6RVRnjJ2L6nXwWhhfR
FP348zIRmaYp5CmIHKijGdTrB/tc564mxkm5c9OBU2mnId0TrMWuKSs+G0V8v+lporgSj2fXOZ3F
dMZZCKUXGdUWkQia7kdvAYlcxLkkuNdwXr5z6XnfuWiT/RD8FwwNaDaASBljkH/GQMyZU8ow6pyk
eNSMiZNBIy8fsV6urIuL+IQe58OirrgOXMRL4QJ6ipdkX4jt2oCaXEB5KpJ+VKItqGR8p9kdLxH7
0qf3j3o+9oSOJtRR+mBvu1YFxBRjsCCSClVEmskuD/vEmH5g7J/DOjmRGPaYeHMSNJmF+ecoomGG
LhDscwX1uQwxStsdaYxG9Hd2oDGg3RKRoBzCwcL0es7DsTrBzT+19tOmZ+/GJ9mLuMzemVG5udYC
Eq3EgiR24OUOVOa0gaewVG6pxfn3PWCWdfTqVOvOa3scWKRf4zc+jj8+tYFnc19UssG/tHyq+IqB
LwnlTSxFh+pP595ERh1aLm8kaX9HNd3NrfMcouLBEagyWkQGRCw0BzU9o1uicESadqOpmr7XyDlD
yeh88R2Mm+N8amSGJvrkBAjWlRDXWomAS1V9vg81fsZpEIh1nwyQpyLJP+YvNsXmc+4vnCdtPLaK
3Bj+3OoTGHnj7ga2Z1h5QALtmD9AF8TgRfvH8LLovVkrk2cOGsvnYhpVhYBc0bJoFhBfXpdny8bD
JGb8KfajtnZXsTRuIQNJViIx1NWAaUfVmir0rYuQICqEiXgvOT5u7pKrqASJrfkqSITrJgAvct/8
kbWtunCdY47kf63O/21OwMVzjJdLSuzjzmmoBJtZoY1kRlUqRXPy9hF5Py2uP+HxMrNerTQuzwHl
iVyHDbkek/4zatQW6KQqHE2FXRgUNhq16RxDeFbLYZgJ310sXTPoDfKXMl+hOLodjyruD0fMnqPF
dM7JpEF99DDy9AXsVSHTT3WcOter3BbyprdeA4A728iJoSX21q6mKdXA/0ggZVpNzpMMNSic3WmP
Dl5H1DIlTzqLhkIIQFiSg8x79A+2hg8FjnrpRDHrxEiumaKOl71JjjkRMqRAIBjeeGs7nkUI60MH
UGu53UCEq4ckpxhIeuwY0W6z2z6ejy7JLKTAknrqQpxpxEx7gqgqUOPghsy7Oer/Q0qY+CITkYt4
ImUFO2wEgobhJZcjg94tMl1MJAttB7qRSKXyEymxwsIEowcxqv+0jWpIC8wkExKJRAi28wvUWEPS
zu6UE9Zxp/sh7Gyd2t1jhBYAYePdTFaTejIUGholGFFAhjrCiVR5hnqxAwoGsWza3UZjaKEl01/4
rrKx/2HgSs8PD2mZPLHOq+MiDwDmz6gKhNMTbA98WiK8RfaijLSGRTeKxB1r0UiGqdDJCK2QQrix
TrVZQQUoPdu0yuYYYeKqxVkRPllYrcOxID7Gb48BtsdKpZdfl3SCaAC0i5bRloGmbXxemmSWkn78
ZZkiNvJTEuS7UZgNAk6NVzWsgtwz4a6PxuKmQxDrsSXQ9nTuhTFc+15jgftyA1Ni4E7k8vLyuztJ
mdt70jcUviYrUo0iSZCIYUF8dGgyasFdUvZT/4bIMmt+Eu9NIW7PmlmjrZFXm5Pu4WqJu2ANI6kL
stnoriREPsGMufZ3248xAMEUT3Hr0ludV+J7klAjpjUBFVW8rKLOuafw7AayEIbRVYSCkFy3oj5C
5GhIPDMQvM2hv62qHuiR04VpgTEFkejBbVJKS+1dsNMoAMKmATgkaRVjSlRTWQmMXIZzZA0ZD6AZ
PXiNhTBefRE1MT2mgcjjZyddlDAwdy7IIBU/x5nqRYhJzmPBPCaGYUTuHCYOiglF9RviAcQ7xwSi
00VrzivY57Lj3e1VghaxgHOSL9YrC9d0yQG3aZ7lASm/5JAMV1bCLCLXHqcfGNV+nte7Kvk3oozi
fU9szbWF2wwvzn404/wM7YrwaJVr95yK0bZmTtnb9sVVMdJpOHJVR60OWrsdjRfbJDftoyufgnjv
aeZA5CgO7GEzm7wshltD9CM4V06QkQBilZf0d7L9FhiJG8guppS8RUcMVDiSL0BCmIejcEIDaVh/
TU7TRAfeJIj4xkyDITfAlFBW8k1S14rx7u04myeugT9nqskCYjn/njHyBq1uQ7pni6sUDR7nLC6d
wxx7hjxMv4V8BNZYH05RtQJ37A8i1c8XxlF9twwr+vfiJNlOuG2bpPbK3tJtAo5PK0YTwtVxhJjx
BLBhsowQQG1xgXVY9JADFN4STZE/fD9S51GGu/Bfe1OCNLKU6qPVicXCMJ6WsS8QGgCy2wK7VAQG
8lgA8ScYlAZn3/HSyc6ph3MIEiUhJ3GuDnesBY7qPAGLsbGMlPgWTzEuGGYlN/xuQldfLMtckXIG
93+tR+Mej9k9LET9+MhzK76FZwqODYsFPeT44bX4DmoDBZy9A0q2z7771fjOu7HLdVO78H65EcAl
b8+DAFujp/QkQTz19ICP1sPqSdtyzrcKfUf0chJUratjfRcIlOJHNhw14jsvso25lUAIYqQXARGU
92F3q30VQ1xFC4KrKzV/Xu1H3C6gs9qQ37taM8xWTUl+VUREFN4phVqcz4ZSlKpgwS9o7prH/8Ki
qCnJEPmirCPGhAi+AfRUdBrYxj+X6hKmbgRji3Dtu3nloOnssZanpbC6YnBOPQTzJNn/T/zh2jdD
4C/YxCi3FBopN+QYwGRA5WaT43KSZCK9zD/XrsXKex7vluL//GbkLRMV+dShN3M1CXnMJOathw1k
TIMHLkc0ugq/vavpODIE12SsmQWyoPZDjJSuI+pmOmDb65ak8cCmV0GlvsjeN8NyrRh+tTqX4MxI
pkwIuPtDKiLUC6H6mJr9R31SCMzWIAunB7IBFJ6syNbnYmV3VENpqXGSlg1RpmwDr87Y2X5pbOPW
8zcmpz6qmJuvMMRjVCChuHj4IL+jJ2KiZ6b6R4PrJtEJvcf0LhJX39bqm+sUqVFHBK5hR/VZI9Vh
umy2KHdV2VOryqmV/xXcFKTLVjdJ5N8zN4q8mBEQmSe67raanheJYMD86kCKtwgiQmVnecikufzV
DgHXJkUbg9lEv2BonoKX5hSfF6LAUJa6BBf1ETOdovBktuQKXk82kV7ju90v+dZMfs2kAH8gK17v
8RqAfzH5KhGD7ZynHcJ3QUkhLYdnx5OG+OLgvEA/gh/kuyhBnHrlvn0OPai9kSHM8bveHrys0YMA
9hroZo+EQScinbQPuoBgH3QjZniKVaeN8/Qh+L13FJMwneF4YEZYW66GzAqWegNtIpyERKG4F5Hu
d3dphGiq6RWLN3WvlFhqdqAW3YWd3DwKfm8mEiyQ3Anlbo3zvAxxbOH+oohMNjzryfJNQoqKziQC
FOHwrvUY7lZAt7Q4fOHHJ1S7rtdGvkg2nLs5d8dizhF//1t8vFNcVHF7+eSaLAWhcDLsuhGDAsNG
Dz6H2yL99XjjAqOZ5mgeqWgli8W8sHcF+OT15ObiCZCPbjgf9gWn/Ol5S2dP2DA12hfofxVlTp3W
l7hA6EbDapGDjkTPYCsMlTrWRDXPN1ghY79LJMJ6f0VYojbHqyUHt30dKRu6EqEPVv3hg9YbNq1E
XemkfSOTzvGVBHk30efnu2k8LQHYyJ6B1IxTYSvG2B9gkMJNMlpgcdIcgcxhpJGJB08ToKWc2rjM
cwUiITc2YhcpheAK3/kiVa0dfUMbeASx+D1ZucGgT1UpdQ5c6V6IPHvh4WZNF3y3AzTa9BovGdPF
aYI1y5GeSIZU1OrJCi7v0JL6rSnaum43I8X9ZYr55qxCyWKo+72WoQ86b14+ycHZyDrCYL+vQxUc
1FC9sgUzLWsiw/YBQ9uWvZ54cINpEPO/uZHQMgc5haL94GnwH1ysyq6pPmnUKuLBGWTZsBTIjZQX
Hx3B6IHWl9ixAiI83QwLShkf8/ndTyRz35ItdqFLz3COVrwSp2mV5MKAtyHFZ0OIsbMo6Z59wl0d
AMoGA1SOi1XvMEC2dSvw7aZA7dB5/TAOq5rvHzjFtjHDBiPVYYyUyx/1Ex10bg3RMV6r+XhVzves
5oBy7BrT54zGvLoS/+NstyLOCSDHgTsnhdSGInRWpzOTqPcJ+Wh7ACa9eYag4lAbM4ea/MqeFhOA
uGsvP9pAN4m68K/7SGkNPQ6g6QDzFd/cGsRhDbDnRY3rwslOg0IzPS0Ur3Tv+dG/laBXO+Sp8cGR
CAJ7fX4dmRnBYK91wwih867TPjRG94s/rj4IXfd9vgj/Nigg67JvssmPmxdXUwqpEKCuet82fk3c
Snjihd4b5nuO7J+OpzgJbaS6CxG/4s9IdeshpCIwlnyqUgbEu835Cc/nGgxV0RIz2mFiuRLOvPof
KfkN/T1LSiYJPThX8zthfh93Ym85ZTSRuYdbnxuPMYrVBeB3A3SoDhcZrW/zm2K/IxJXSBogGqrf
6BCpaaIl5vHJNw935cb/Awk+Pq4oouN6jmCwVnBXQHFM9Cyi6IJvzM6tXuVDtc4rUJpTZVMGKAvs
M+E2etYOEJJLsCF5MbPZZaUheArTiLfBHPo2vRkBkeUMKOOjzMlx3dpWl2RykO9q6Bf/O5taqlsC
l1GiUl7HHWJGaOHXHhKx2OAchNFJOIeHITdFkw+kLCrTbxbc8YJ/oyQPUOEaoXL/ypTTcqW21jnv
VMCaPcMlaC4lCPiDGC2FF3mz9skQ1BBi3ecO/NMiZaj18a0wgu3d/lvRJAC6y87XobmbtagkaXNP
ZRD+nEiEuIc/rtggG1rfzD++v2ZdwQGCNJd9M956y4uHrPOfRulcMXnJTqYSnfncTa7MoZsYCOR4
MuDMPwSv/vcg1NHW4xR2e1j/1S1bk633X6FD4BzB17YX9qDzCv3BNBGU57QD9ejzKbs5O6J1cGmm
UicS2m04+6F93o4AXPkFJ16gzPeErVBWg4k7Bg0dGAos/3oXfmGaDcxcCDtYITl3bKn31FxzLvZ+
FiM1no1yM3iFwbq88GvtSTkdhrHDA0tDW6Hg6NiS18ONCO1aRO3eVNyU55Aepi2TYda54/wUAYbx
+JpT8vbFe/lDuYZ5wT3U2JgUd3vGUHsZcGPkVJRO40l6P/qDvxZ2+1qb07LDzR4vt/HHifqhTlNR
zvFwlgTYY4yHj5r7s2mkVWblRyJvp6xK0HNj2JdtWlgqeSaCX3h5ZOy/GEgqseAgNTDSwFXYg1jO
UmCpSF5Y48T/g+rvqiTKkn10ybq9iRzXbgk9bN7Q33u1nREvphnoYJZMD17jaQui3HTn9EpHIcfm
ODCStVfr/O4jlG6d44UCf9yMPS3aVqkw7cP3C5xoxPS0NHJ9lGGaG3EQBvriniGBGJU1R0gIfnhy
BJTaRzXMKAoTvF5AKiZnQSdRxbXvD6z4ujk7YuYikMzrQXDlKXlCHA3TDT26nXs9Fq1I+sKujyO8
b83RsMbsKhvnOC5VJm3UInMesCtBBKGYO1D/dlb6DwaXi2bY1EzWc62xh6D05N6YJFXjQXzaQaJn
PD7g2THOT1nA+asPekoHG8qcnxF8JT/mxgUMU9UHWdQdubPFhkMAfoXKevW4UrQC0JYzzlWLSJ/u
iyVe1Xt2c6yqPqmMcKGEaz6aZfB0b52D6YNfUPaf1x/l24bOkamTQVdLw54wyLo8d33BChXg0XrL
pPTxrgIJGk0g4o/vKF4A/K2Dm+6Ied5Y55PjsArmzYef/fWHXr5xe81Z6EVsfAFy64CYxJff5+ad
Sauv17kN3Lc7+taC4cnXwDg8mLnF00UhDn4fNn/8ytkwZGkl2mSGF10yBphqsPjcxDXM5T9G9CyG
DZCXF22KItsxel/RBCnMFxKjqC02n4aEZnEw4ZlqH3oFgJHZAs0i0FOg84K7zmVM9v5g8N3m+hv+
4/UBu94+o3bUqnVK9R7arqzierxQ5HVt49NFD18vbzkr9lSsxx50AsvIoS7TgwQOof9sY9J2e/1+
jZgmnNvbIRa6HjLHwOkMALBFJ9EvejmlMraGibT9YMELFEh5X+YYarbF/ox8jar5wb06psE8Dkdf
S/xPMHGk57TmI92V8ad0HuH7VTjJfaH/ZC54guvOY3ivBddxhjI7TgtQrrqUML4dPIDBBvWEBaet
kSqaiImPEdJdi/8yl3+xoJJY/BgEhVBkk3s0FzpwwmBrJFtGrQRzbH2AkqkjqCqQIpHUYRALhwNV
SrQT2TgJx+6dKv9VWqGpYxYZ/xj1u4g4zn19bV+Nuqt0JGa1tSEBZu5BUn9rDo0uaLOtKh58dLAa
0eqI/57QuBRD1bWKB3G2O7DkluhAgKLeUu/hPWt7Mrefvn93Mh/L1abEfLuBthKzrEDSM0wYjh3m
1OuW3ovA3uM1v06xDkzOqJAwDYufO9mbhdR509cIfsA7I7FcwzrorZiiip9WjUWNXatveaEe3HM5
yUjS4jElFOJnrd3tfsvDWbmJV1wpwT6K5Yn15tilnQ/uP2bzqS7sq/cykvzT7yXxPTLr0L/qM72N
ebte1y792sOcWdZkcoWVwcp0Aktfm4eiO6aPC/c+EegArnnQ/sxKDrDAFQsAJVLHjI3ooMecNFg4
f/9InmEvgKnzJ+41Pg7kVnagvB5s1t6H/Gv5f7VhzMchs9BNFrQyOKE3hamRjW6dJjYE5Rla9/+e
BHowHWblo0Thpp5pPwvLbS1Mmc7u8+u+8tjaO4NJjBOTEGzlaXAP4fnystB6XIhqnVNRjF/eAn3a
Ust9vSlwAGW1QOnvZcRiMI+vmCNnsou8kX/fWrtrOhEJ+Md4l9Pyr86I1ZJCK0w+8v2nGuj/awY+
i0/IWaUacoocInYOSJOkbdO9pI3Dtm5IeDefbBC149naDwc/4hz1oPaqi3A3TzIBPA/mlSpXrrMj
pMSu3558v8SnkCkU7OEJgb4ngCLuNYo0BkvjZrvJV4QjRSP1zbjxEiHi7j3j3pF0aFat69xSljCM
Eqta1N+WwQv8GzrlT9muWgxUSuHg3aP0wzY5v1fjhJKmUukcTn0oMNSZzuBwIuy0SDlDA6fOdix/
TFwL2BI+nZL4j4CeYGUhMW4CPp1r4eU5kroLua+mM+Isw4NfvUPpQaNtp9q7vU4rBijO0aGcbznw
efUgy3l33p88tB4eNtivUu0NjLDD++YqCqwLfVSK7+4eS4blGXuRmR3rM3CbfRcUl0ed/OuqxHaf
ftnP7gsyg76pu2+a4v1Qcc91SruoLoQsXQS2gOx4a2yBueOUKkzni1jTPlJMQBtyiFyicEUWLxWK
kiEQfWZMUZnAVX8haM+b+p0csZRwg47050ps6eWXFC1L/9nVpsZ1NNfD47B9MCrKZfl8Cpjl0nYi
VkymE2McUF0mOnwtoXkYaXr1tcbSeHMSrk8CjZ8hXXdUEqNaYz94VxDddUfK2cPOY1N7fk9GgKPp
yKYs2jIyAPwT7CYOSbGtLTONkNB2Ly/fdLpWRrhNM5NuX69z4lfTB7fT/9jpATuNvvAgy05iIUWi
0G66GIcvQfOA3DT1I4R9uLRh7Fo8ITgkvS9lJxOz+t/X0nfTqf6am+MIeKS6flbPngqvrrXQuysz
3tDtKyU8/CG9ypBfguvIFMwyGHwc/S/EZeuWlaFIBmzh2/UajDJQiDcBCdLml4ecmIHMVjPu8Uhb
KxPI/hCr1uZYwtwzdUr60WOSfv6ht5pb5UC/VrDfxDSZGPcwtHsljBBJl1wdO3FopQstwsBVQbdp
Utlnr/8fPqdt5eAjtNWDiFRRAcM8t0vBx1w+LIARs1RdKgR+lKqAo93dMC8+vezudUQKY7DdkMsX
AuVFO+2+UoduldKAOx4PG9wq/lmxQnQ7TF3CaM93UX879J9hjJPsxveY1tcuHZqvcuVZrlKn+7Mv
uQz6ggf4ZbmyFHMmMUwShbYb6hdiO9bt43Xkr9EOjYOysqW3CJeMuZJF4SdzaUukk/qEPeijUYox
1mEe3mAkd5/C+pBJwDyIPZ10GQrT33eYac+DwRB6+XzcRXlwILgHF+yD24uFju5Z5LYAvjLaZnog
IG7vgeoos177zOsiJia61uiVMr6sYYV2Dycgln0u4h4xcjCkR6/jYXd48kN1xAtHBN3rqY9soW4q
TYFEYLtpyB9woJk0xFaIuuBu5+6HvSDJL4h1Ja2MHc9YV9PgbyY7ryNLYA3ykc632UodXW8i2YGV
wG2WjeaXd3ooE1VKypDNV6ZUOMfSKMgTI/qpjy4WYwDfn81QW+mXplFrDmR+czONnLMx24GniVLD
yUCVgfw5ElbYfx2CT8/BNZ5C+T9nMHnres1GACXIIpQ/kREvR96FaKrsETKcHqOGM+lwP/s9QI5P
ZNtmHRbEbAPWuUEBiDgFBdBoqFBNJU43EYAabw8n+bTXnYzvIm0TAPxeCvOtRzLhK0WqgUAnyVH1
FyKmNDzoEiYtu1J0B3SHcbGyKevV5UUZu5b3kAtCLBSKzekRKYVMnG/60FyiGs69pMMIq6jZ6H/g
i03OfiuXvNWYL4OHiwcNch4CUJI+SJICT0dzOaUNQ37aMdkdWSjs3fZwXcO7V61Ry1lPZ/MFiFHt
maQ9QJZFkk6bvlxrh6LXbd63m00Osbt+DiXctg3CA43iB39DGtOuVpC1WQ4s1A+W1wliGEfDfux8
8CIfwfG6r5WJWU4jhqQqJHtZSWEN8+pbGZJ4BhziG+0FPRyvqxISmjuKKYw1JUDFKnE3EZC62VTz
BovQF/Hu8b14TVg3tJBGiNxeBMrnRL30fxBCyZI5kOVLUxQZVxdYAuCLOiUQVQkCU2jlRArXjZv+
GC3xd5JICzBGE8YxS1IP1uLQGKcChXrkD14tN+RNB3Eruyo0nLLCj+/uwxAu5JiHJ8Os2Fqej8/m
o1DLgGa5m5J/Wu+s0SDjWBfAUou03c92MKnwCp6bCPFJHdyr16DXEgI3FExo9O8MJFQUaqbrkezI
Etng8JKQEjZKDsP2jW/fZx1XayXkTFIfL32UUayhICTaZr9VF/+rAjXnMK764L3aHXiq9E5fjjbK
82OOR7Hl+c3Wd8FvOIVT37OzuFuFLmtbMRZ6qo+75o8Jv066yS7g2Ewh/msxPItWltAiG0cLkDvF
60meWNelI5j8HHhpd3V83iaD5GYYzLTm4nnNYl4PAGfYGQQ9OYzwjODfYf8aoRkK3+YBia8XG4dA
CqaRhkoKndMdrzPJ6PGiQsmvqHLlsvFOP+6wS+RwMvi8OMjVzZO/zjdKA+ABZNog58gtQ+F+G93X
eS4Dn+ITNwZ+w21SMhZSpf2NlZqK4KBLqzMmZ/A4Nxr1U1Y0yP2qQ2IcUr2gbWkr3p+7N6XBEq08
P3KGGANwO0HchFem65IzNHsrwAvB9gHI0K9sIJQNucW7sutNAJ1X3EKBUp9rhat6GEy+b+pYrAq4
If5KHOMNc9fv9VyHEDfIsjImO2xeeTtox+SgnACLl15aOG6bqhQ8KosfWVGhosiUaS4SaH7R1lXk
5alky70uVZRNF2k8bbS92g6S52J+1ZrooMSKTlADzAQjySXITCxD0Q20CrwQZsc0XkeoOIt/LVQ9
uuFY50Dgj+NeHCMD/Gp/zGNP26ViW2pXpVeo7dvUMr2blfVBNEhUac0z/jHgPTigQ/xxpuD1BaTo
66mynTco4eCS+ncGf93VbYDWGqqRNLKgjXHozL1/X0K4QgleRWcZnrIgMyuCabVBFsZMuX1dvb/D
iTS6xK4Kw9XyXTzbbTY9u6/xueXHIbisLJE1gymWnWHFHVc+bJ+YVNwyqaHHFVLXYpJrc+vaXXjZ
AADG66/V8GGKoPZr/yASM2e1e52j78uvTeUsoVPitbgNxMsrJaqEYycgf6LyiaS289sdDTn/Z+3k
4GAuAmVp0fkUSQ7Y6ZhuhUrfzptyt8LuqNdNzB7w8kKj7S6CUxwm0Gze1T5yLb2pM1ESHWWSy7Qc
AO2y0G2jPecYKv9bE4D9UDN/WTLxSd5AXt6ouW6rPzqjNmiVlscauffOtVt/hMDYVRunBbBT80Vu
GN+IYMRRVvOlohBBF/mJCfWupamxuvd2uE98uC+t7AXkewSZX45eGG0ceVKwmDkK8HgK/UXZJ6Zh
QptQ+JZUfYmJQTL/8YAlNWgirBW5QwqlvIZsLwcCDgnVAFMKuIm3XuwAnpO7138x7TQaXRsOCDgm
ltAJmKyQEhX2/LWTMSxIhHoHTWqcxqGHxygRYLxYGD5sq1iBltthmp5nFrL5n+vW9Z2ZjFVe+kEa
mkD66bofpkYS+IqOLj4ltTOjMadvSduE4aNGzXTxrUCqFgSLWccdB4aY0Zq3i10VHy+Z1BcviZdN
rrqCVcXO3ouqLhBSd5t886sNuzjHujgrWDud3sLjgqhzIwysjduCVlYKLe/q4hk4AaBiqahoy4Az
xbP46rRbbYz486m3EOEu9unAE3oYhqZzhr8olDG1mzmvZhzngS5QcYb72HEiC74Xr/iMowy2ve2P
iEp8/vMkR9lUDr+kWr1W6X/wEoFeMZQqijbIuSpGEiU1Al11rD2JTVQrybYBGeHw9XpnLSo2XXQE
XlXJ+1NwFTinoGIAxQDNaivAkXSEhGyQ40fOrrP7iEekUHUxlF3w0nEAOOPKL8RV71Q+i7Mii0mO
2h4+04dmZ94g40Vc5YaV4FJzL5QQocbkHydG5SbsVQynBgvRVu28K2Inz5+eeneiIXinmSc0Rr+l
A9y1+Omg5qdwbWM8L/tZFLiKR5ARRZfJ8CMyz1OqSsSN7WqcFBNLqvfCrgLIpGjqz/PlbbdU+S7I
KNkHPfnSYYX0hRI2ikniqRQ4vTRiQPkHmiUMkNAwIPxUpWp0igVUYz1z1rAPFgwZ45bu9nJUeHkg
3Q6ul0odPjzydk6GeoZYYzKYS17iL/O6Sq8fcc8CstOoyZLHknTuZ+gDfVzMltsuw6JScXAOOrN9
TQuWfWYUKy2IHNoW1i0hRUduiNEcqeNiWTtVDD9VIiLIxjv9MbOYisH2ICm0MJHwH/6Jqa6olvYM
zG6ZrETkzi9vyBeZJZXH4Dc/qEddyzT8lrlVbyFr7Wo2Zd2vjqK/YdSKl14zI+GJTFby0gFXfSl9
c2y/pjGSZR1VBQhGN/9v9kqm0Px9MBHDYGNp16sQEOBdbrEZtApcUH33spGWcfmgql5N28Qu8Xo6
rGml0tUIyePOKbQGN3ARRVXpi7RYPItaVZ7f/sBv/MsK6wTG9j+DX36JPlhA9BpkMxweiv6r0dK/
s+t5Zetey6ICkPgA+/V++ta8beS2cP1U6nxPjrOF+pjLHfa323456fdbLmTxeApMomm3V+/xJbK0
3kcGu/00fpsE1rMAmX6LzEoschDuHgw88lDFt5RhDEca4BZZkpKyrwignuUXRSY7JABIUEgEChGA
0nCaZ0vPiFR8NN0IwWEa249ow1GHsFGaidLuUb8FqAlnKLIq6pP1aisN/P/1gSccQClpIJ29P3bF
fkHdRKr1sboHV/oF3Ovm7EQC27fh5AF4hWx7qBTLVe/+p4+joz68cBhAMux6vF9JyIwXBxZyAHus
nVdZMagDD9OqGKYqYxCS+xnHb5K+Tgs6F102enHCa5pC+07TFN3wkpF3FIROczeVK66HuR9+GJyG
GAav4F9/1FX0lO5pospEGJvz1iTII7PFQtmE9717MeMrgQCSwvoOt4z8f+YwQIzLaY5B1vwGpL5x
VaVq/yR4XumJxsqTEoF1mPp20KORM1iB3SA/haGwhM8W2OFAeDhMqViGlKkt9tzNUEc3Xi3OU3FU
Owr3QBaQbFxc9JJEXG+R0bkhtWOCAXGmmt7wTY8ZwKAs/QUeXdDOdHN4Bp/HRQgMDHrX+QEHXE6T
2UFzACPDJ/M78u8WobiAiw2ulkoJCqaSLsVjK0+ceGdKBLMvxluz1QsqITXn+ySURugmdAz2Bq/q
PuxezLU2QL+a6k9M4bQZLkb8RGu3n9wzseMQFO7ul4rU8isfgp+OlzC80R6yIngrwPuA7yHokUpn
/qC+kNN0zAZxymmde7mBKg3Se/FLV+OxgSpyNM24HsIjapdpGKc6rhLZl6ql32oAgiIhrZEvYoKG
bbiyiNSFnbpYSL59pcCmLucDCaErh8H0Tr7+4/kiaD6kb3VKl3upA7dE/vclOF8Rai2VbJbdgLz4
se0k1JCZ4W4YVyI/nRUS+mmDblSfkv94hPOropHWK67mSI+HsuLKA3AO3mlaygjX18DUPghAc/E0
0auhAcPFatUheMm9RlUWDAdFHLHYfwg1ahdAMm4BdZtMM5+a/NN7MEDavevkeCajbeDrzaVPpFnW
+CZHc00sN9BFe7oQo7ftg95q/+H16NOCgs4sGcPe8eAVAniY7RRV+J+NX7iwuceVSThU4Y+glnoD
zyMAmDAy8Hng1Oc/t0jWURWIzAEeH7AzKqiBWHFjugimot7mdqoLRczt2D5WRcWS454h+QUDrqsN
KOfsj0xcfuPRuatyEOxiY8Xyi2AzcGitmGNM6ifx6tSKWHRqwE5sKB2t4OOUvC54Y8DQDPZJu2Bl
2gC0eT20KgMA+W9JIWfgcA8EQx30vyDh8Lgume+922/v6TcMUfsrteJIip+Zv/1fl8UDFyNGFmLN
59du0oCgRsaukk+7wxv5aR1tHuc9sCfBQuKkqjRsi5vT0uBdaGcZdfa59EbXUtho9vY5hqyx1JbU
H/MZZcu6LwhmWvFUVnOMeSvo00LTlbSh2S6p8rjArvmwpGj944ypXs1R13uuIG8qd/+2y/eS13TJ
i//jAeOJ0VR91oBM6tEg8E3K48VKAhdiyaOjXs5/5GOHU1EZa+cX4P0tTMyK/W8TTZO8tZiz0g/r
YfjeaTJkNLBwIiOet6VPa+D0MMoF4Br9IGTdvCKY6atTOMl5PzvvXQRJBLUq07yAZN4nAPXR10tJ
FHfzvus+x8vK2NYkT15zjMvW7GGIZqlFS6yB2AaR3JOfvJNm2VUT+PfgRE97NngamfYd7weVd7Ta
B7CeeEb6L2ZccAsWS0zYIeXq4jVVeQt9iii3y16E6TtKjrqqCdQASw+JJRgpczX8No0l1PXs7xoA
NraPEibLXiT4eVDFFqfWdrahopuqydsxSQj7R1G1sfL2rKkIKLpAsJE8ST4Lb8KD8hJ+HCSpgGsC
akgW0KgCG21aLhnn7ycVAoGr/QeUu9f8U1st7h6W+xVHZ8yl02ttpB4fM7C6zWRT+wUUiUAViLSn
i0cvpwDT0wkuhhLJm3WF0SiP3T46E9oqH+JtIOJSW6OvCt1jLvHF/DOzQfd9SxKmHNNeB7cdcs0t
rRa25W79dRBUVeB4VwYQ5h5BF6PTqy2DXDBxQCPE5/mhN1zRJ6ETzL5AuXpqnvBzfwF/0KtED8Pk
0KaF8IkKTlUjSQ4Otbfo07PgPfCDhTpLF7e0eYt1Gkx6KYvOhCfoPHI8e6jFz4QBM9aOn8lwQaX/
RUUnM/WpXRqf7k9MBOGPDzp9QIXzDThi9yXcA303TdadopXI52k386aEyi4KwpYh68jA6Vm5H3jk
+nFQdBvUpH+qkmnRVzTlDPIlEk2lXIQAnEEPVmu2b1JBcTae1TkRbrTdCLfUv2lFn61b8XyExb2V
g1yaKpRLzUEMpThMBxCAJtTWEZ9F9j9NBPxtLf4CYO0/sLqkY1vNpp/2GwMujcjEb/dA6+KgUwcE
7CITCKn01thtvhkAbqoMm4VMIiV18FqQnwH08NdK6m2gx5wRCHAsVZx6R58jRbCCbwKCy6shX3cp
FXGrE5yEcifXt+XpllgQySGS+7aOW1/o0X9Xr/vvoMawKXYYknKADDGZp6SDn2P5p1rCFwVt8ZrW
b9W5G6AmIX+AfS1iCEQwZfUWNYVg/moMyLUvkJH97uR2uhWCOtUI/excBWN+lxnnNhSXTv5V3DgI
OJItIInpK/V/b1n1HCL0UGSjRYxzF3DPkzfxvUKsteLr2cDlHYOR/dIl5pw/zLc4iqIGY+5Tfj6W
3j9aUQqJw+pYv0uWWszh2kbCkccx6zts20nhgHUerpkVpjYdHbeoMKI3fDT+3qWGEiZwLL+nRNLI
ibAKHrUfp2Z2VYfbysMJKHKAGMUsMDpa1L7plq5aKv3VDx5gfb+o1lN1L2Jtjfseu+HEJWYgrery
Hj2QLa3lblpg2vSB7rSQGD/a+BRq9Aeg5njDm/OMZBUnOHYgfO/zMItDVlrHJDdnABINif1oFW3h
HdfZQQxQW70Z3cAClSKyXvc6xlqQps8jg/aP2xuEsUNe9cWM/vekK/7Z3+9yvUeGILKWlNcD4Zti
HUBhqKE+d91gdTkN5Z0MEh4J1YFV5LbQ98Wik4PUY56rxlzcooguKINRtB+Qrmu55THIHEF6g80d
Aw6fa3ai6cxT164O9wXYxYx7/QkZCFGt9mW8zhbxmfqCc6y3Gw6wMLyF9UzIFfo1Hz1d24akPR3Y
CcgGj3RWHSWcMYbhzaA8jp8le33d+hexFDfYFY7OjKpalNcXNjEy/OzyH5uPn7oX9ZN+FcHqNhri
J56Nk5pUD2vF0+BtJWB9mS4898+1NFnR49NF+dhlY50KWsUTnjQuA3HXgXVzWROOr9pQc1Y9OBT7
b79J/H2VOcZioEJ1FIo3qobyXRWMKMEdX5xtjowqvPDcFaIiU+zR6Jmu/g6J+3ZOKIkeN9HWTWrP
QChkoGwzzkv+bv6wIErVJtLNj23Qa6KvNTVEYhRh7Qoud/+M4PELqpibqTKec7Dq4qlyyVzwJdKC
uc+E24U6fm1D+vU+vCc9jUswxKqBTH7X6KV961i39365CE1Q3lWgxiJ9oqlx3VVL2a8KRSf7PBTo
icdGRmkvrOEmeC7kBaNgLK5ACKO+Ship2uM3g9/Y7VLADqYALn89JRG9zk022ut0xNKM9rfhKFkU
ZB95XaVMH09QH8LStxyRYMWRHpQNWshbVXfAht/JgjYaC2XABjWnnXTMX/8jBkkuLxvOrNKpylDf
9oBvoxWgmg5JaqqZqCY8X3DOuIeBOQoazkWgwNayqhU1S/0TIHgWzEDdaC9SMoGHlqB0olSIxmM6
TmlLTpX5JN4Z2vyX5C3V4LQZpbnrQjVArA0UZGy7XU7Zmp4e/L1Pq9MClEbP8ykK47wRJUpVQByr
+FbR5183vflFYMjqisvwcfunlNP+1pQ3A9+cHBdZEWXSVPDdrJilLtZjxehWg1LMiP3ACmC2cVu5
tIe9rmEeBGXS5lPBMT6CItZqYRrXCpq88iCafSZ72mkNExQmkle+NvqXnTfDNPi51PFu3c2gD6KZ
ZSIbJdNH8zX3jmnyxfcKIG6CxiNe37RUzb9rGqfkY2dTtlnodef5mldGq03BPsx9WgFCpEm4W1Hh
ToTi3CkzOlncdAd/lNJqfKLnctqBfV8GEZRyZUEVIGVI/b/LvEcWd3VvKwlKY6MobXR7ApBqHR2m
7wG9fvDm1uZX8AaW+A25uDUwDqNN1sYaNd1Pa5wgLOG+br82rf1vZ/rP6ifSMBnyV0GX2V/B2+t/
YNfWNaqp1rBq12plqiZF8is89fypddNhYqy921nS8QlVWTvXk5idpz+yw/gqL6UDgRgn8lqPSo88
eczOKFkDFuixwgVUzB5IFJBm8il4XkMWc8P8M5JGKFVPL8GykMXiaBRaHf1/wqXMTJu22X8vO++r
B/KS1P6wCXzN6IFkRcI7UZ+pxF/oZozUYGPQtRIZ3CXYUIK3jNq9y0nOXM+6rtTNcWdWe7AQm16k
+9/ja95rmdSXR7xJnOORc8kIMGVQXN3tzRZsVGttF2eQNjSP+LlzneJsXvSgNVokMU9kEpYuw+4p
FbEV7NkYjUYP8iqXX4Gt7jDzsTnab5pCdrGmyaNEc0CnzDrFT+8GUHyGv8eH6EfXcVl/Kq0CH+dS
gbtI61425tNXIjx1CWhLks5W+v/v+e0jSOo221Vx8bSTpDoV0oOxR/7tUQVK5MHYg5ROIOsu4qEK
WzZcjunNAkzcrg2Dd5F+zRHUz3B3H+qGoMTDFheHPv50ZpLA3TkFgbyfzlgzCXKGHzMt/DI3nT1T
qBbltW/2xBlhDMkutpBd+1nd5nRs8CTuG+KEWECYx3BdtaGc47xmwzsZikuePqy670H1T5+Khla3
1jcRsdCKbimXBhbeCjpLlC+csx3RK/JvkC+8Q59Wwu92SZFNSZZJ7AmSdYM2NgKd2HoXEkAAByVu
ZXVJjdUlgFuxJMj429awjEGlkb2Nh+/36OYRhw6OXo/go/1fbuUQ/Ov4iLlsSj8R2lXkZsl+xBqw
oeGa2jcqexJMuJIy/Pjis5Us/DRPB9rGP9UYuHzQ7N05orfM4PHJ0pUUpLZn7M6W2xEkvbXrRMpH
rb8b0OhqaZ1KtZreechLYAJ/5ZI/kEspNdBaGAjo/v3EN6tXaVEK6FR7UN1DV1EJ0ptfI5DKNI/3
OZrLdH9KVaASlfF/h+sFFOa3lhVNMikIHcUOhRfp/+zEKx+1hR+Knb2ikv31Mm0BVyyYeuoJJEGL
RZaJVEQdPSrn4Zp2hjcrtFCqG4FvM2ChigxKfZuSvetht7SWDUnqh69NP8KzCMQIRIaLEvE2jf6s
wPOU2y6S92gUHeo8WIaJXATqTzaADJqji+iUK5/9aYT03HQJUKkIhOMLUYPTTvTx99YZUoERBsSy
HK7/tTXdvANKjtr3zSdU/PRKVSHG396lQ1v7rWf532m6k89233IPkhdU6F9JJxJenxnFpfH5++zv
hXx3k48vkUDp/Y0dGjqXWNPMDNTFvOOq2M1x0YZM+5+JrFOckjLEkW/nHcrWdn62y4xSb+tx8Tus
F3pOdP36bi88NxWXTerpuuUldlRW7YcYj2jZPP/2NKy1CuuoF6eu49EoRSERNi7JBv8P4ain2pZB
w0YQhHe61hkAdIwQOEyem+0lPgUBm/JSN7nQfwlsMcUwSHeY7nY8+bBt7QipvC27JprxEP+zb5yQ
f+lvXkG507mI+2jecTWmdiGwBoU3f/pKHw4q1i5ABU9vfn/nB6ml/RwjluO5N6+hqTTq/UseJHE7
yrcHASTEiseEMGjht0D3SbSxv1rX51xJNvIbPraGUQ0/lCDwJGDb51djp5vqdPvmbdKfwqxximKc
opETgsYL3EHQ3MVgenen/tbT4ITx5vvcy3dKdrARe2DV1Vq3EJgNKf/ES/bn7jzo+zs+niq8ZJ3e
LXSTxVkpL7htStKd1ItkQehX7WkjJn6fm0LmC/KArVn9D1uZgbECwb+Lz9AyzKWPSMjfvcRqbsHs
y72XaEWgYkGZS1QLmZIujvVPg2/UVqP+pqUpa5853EnkM6bLQ32HiQk2RcfiEpUe3prgxta7r8CP
ZHxfAG5iaJjpcXFEvqu79kK2dNoR008DKXA31mI5EA0nSc9CU1BYd7fmp/cH0/+q9BHrh8dZ2gO7
G7fGHLU8geo2aW7L11Dofn71CciZkWJcMtkEu0LlX3mXX+8D+FHgf8nRLAE1MCngATOlMcdCIWfD
hAd03bu/DO15Y9pnC2yQAm5xQpAgyKElTMHusOa/s2jCa4xe9ag9O8En3uX8QKYZdhhh+XIArBRH
sSZwl7YB4sFXfTYxnZEsRvbvlCEthOKK5gGxhU/9/exX9PHnYoXqDsYTsuLbQEzofvX/Zf0kyT7j
nx7Ji8lPvlLy5/zTXNULTFOAbdkJvVJLe/roNBSAg0eAO2tstc7vvshDCCy1PuegYhO73Hr+FX1o
e8gnofLWiknxg/k4sf9xt5Y7IFmmFQ26AaH7TFqJ98kZp8+Gh2ozFcrUYhNFNjDn1zsk0EST8W6w
MUEs3QLzyj2Hcuy2SiSS2nO5YmXiI1st466tv9xHXdDxtXa6IG9J5TD2Q6duFHXmrlulzP4D3iqs
EE63JuGaBZBj+J8PrsBDbGXufxoiy7iGKwTiqrx52S7/ceTcWS2E/6rtsQ0jq0uDMpBr3KbXrpyR
b4/cQ6Y2XyKuuZZth6dEI0OeaeVE5bOxdFUiaTeUd4D0cnxNOxBxwRHpXNRLGCpc2Ksk+7LvxMWM
2NDFD6366Sf67b7sR8bibAPXaNJZQrZWmxXeGrrTfeaO6KR9e05tzN6LXdx7lwXtisUHIxb1YZ9w
gpShjoFloGEC/LLjPyo1oFBQomlb4CA2xQkURNPFCyhWfcm66+23rLpw69I4SN1Xwn+b1CCcm3d/
C+r8J5vwbNhhsthSw9cibEczjkvy9H+a5o9pDHBIOBgMyBB/Bd6Uy9+gjQU/chCe74ZI2xx3s/hX
e6gx2mNQwUXF+bfVzZ76sPzlgtFPR4/NzutOgRnbKUGiTwHpV+VxB0AssXxNcJAGWtmX78Rnivbg
NPD1RIqBp/JMITyWrvM7yXZJSNgq0jhPn0UtCS5jIjBVnpMQ2mFCAcn1TireJE+G25DyIyBaWLtw
/BBrg1iYeAjMAgzsus3f6QaD218c5zG1AjGicZZbWjPdUKt8E59EArE9F8zJYk/I4qNnfoA9xQEl
lMsyfmFzCOyo7T9QSNPXPj7nmGW5orbvLb3CQ8ogLh+aeTFyfwV5ZQi6fsPA0zu8nCHAiUD1PT+g
/+LO+yuMIKbuXEGvtPnL8DT5980L/lb1IRaK8dhUUuJZ+56SlMPWRhdLadYzoAumxSkdJd9L7QrY
OPAetBSm/Gi4f5MeOegaMCb3aHbVeiAWjiXii2XkqAjiJFcGYunx3IGidn17kxPwkf+sbfwPKQHN
eLLuPKKIuXVWw868ydFvTSPpTxJ+meS0dMf99AQMcwP9Fe+st3Rcs1taLl8CjtGW0TlHVmLodoD0
hDikEsjcYt+/NB5KvL+exUsl2xK092OTaPxCOqZYqQF73njxcSkIWany0si/Nm4Jc+EXTLkFhTJ0
4ci/UD6kCpMsoAylnBTtVAwNLVQ6VHf4/wTKy0URmOmYy45a02SX8KgJYR4jfKf+jbZ2DFg5O2fF
evByBdWfIfBgQ96qnct6FB0m8OmmBEi3I9HJBieToQBDNKZUML2lmkas0TknTzz/Fs5tt6Z15zZe
dTpuRpFly9fvD5yFzl5ydOwrtwCEjXq2mpfcO8tY0kQw/VRX7GX2oqkk9FDJy6SItINl7BeVtmM/
f0xLyPODHFvaEJGcXQajcMO6kYJp0Ayi/I/zOegj4az8cpcs8R4nhes3gq49uoaPuSL6fM6u9pun
acCg2pEfkwiPNEFxI8AGksso/jFRlG4OVK7x5bBqtxOU+TGEwckBihW2bEmhGsnQnjDcg+QH3MyR
HlEJ2dicBhinbePTkq+TW4ePbotohVpvmtIcHmcCa6wnU4D4JrUMLqFlqWLTQ65ZgScpLlXsXDvK
bYdbcjYi0HILcMTg2MFvO4ohqnfOUYia9RUqi1lJSULsG9yH3PWeJ8Qd3V3Sun7IGYNxU4x5XFDi
jJ5bs1bVW6HYtZXpD2WxvC393rw6gYtANdjyY3UWZGZldqdHIsQYLfXWKtf/CbhmEWZcyRvFsk+c
wgrfUI3dJSRG7Y01MJAEbvvBjrD+tyuPtD/4YFbGBKqI0vsC50QSqTGq3KXZ85zK3p86XYhsrOFb
IdVytLxVZ2Id/TKYdZCOPBiWmK1SmUsEdi5B2mRqSQeyzOo31xPjWbV5ZLNUOaZXIl3LlzjYIsJO
EQgyn4IucAwZ5tG1YXuQZ6m9tICYHpOF1iG6OCjsHrKYVDz/v1MRreajy53sUpRM6KtcsOSr0Y05
3OPaAeNk/G257HWyBN9vY/w0kqGwNliNXlyNe4pPTgZL/kCsZ352Rcnk6/OJC5pw4pyhmgzk6cRI
JhiyT2tdE1EWazWDFFF6TdAgri//7fBRVFqsqVeavL6V36b2yDtFgWy6bJyQCX0dZ4AhlA3yn2tp
ctCKViMyopb2o7tuA6idoMsuq3gFdAkC1E1JNZTWo7HdQAWcuxZHduPo8dt/nNnYf4f4/Q6siBNq
T4Kr2HFM+k3+NwFTF7SDdF42Z51UfmMEe7n8YJqanwgoPBaTnJx0LZOONAb1HbXijX83Dd3z5UCL
a7GZ3gyQ/uWSGqw4/lYiYYqtzz+2uqdF5SdxGiH8lrD2GJMAm2GF+2JOCRY4gslEx/Gk9VCKoOn4
f+vDZ/KNPPS87OZ7P9nbch2I5w01qKHuZaKgAq5Jufs17ZFuLqPmtQzn2BhfRyPcr202Dw9WSYJZ
/9jLHzrwo6Wahw1zM9QhFcMpI4hw5kXw/EGspwJeNMByLl2pe+soPphaGE6h4vjOZrpI9PJbvURS
4MJrxottTf9F6ZfcP1Ki1jAWnMoqaMXrauUm+BpEudeugsVpZLh80K6w/m2gv1B9QS6m2Dy3vwYM
NvPVCgktbkpv/S3efai/EKRPd1ZdLvcVKcWgu+GEIws1TGq3sWynVlBMfCuQmjnC1gSV2aDV/qf2
0jvFWC8eL4vD3/PkQGsj7jotiqcoq4mXDJlnfLfAikKd0cQATeyTuSg1RFqTbMrZPf4hH8sTPBLW
D1TN485GczAOTdhLUWyGbAYPplRPQidcKxCvqFr2UTL0UkVYkKWPUn9z/KIG3507ZL/Qo86JuMx8
x1cRmJuSJViW2nZbqgN36RAo9s8/fdAoMKPjYAV4zMQYpk3nbYwIpTsjLqs7pKyqm0xPb/gzDaqQ
HQwbKNvEU6vskCcI87oH99E8KUAWNchnCEq+hohUPVp1gwwCKV2UL25QIGdGlNt0R4nzmB9LhCY8
anE1Xeg07sCUKOeVoRR9Zyq3IqAkkbmd+DLahWB/t0Xo5ZY9ToE6DxpqjlsF8C/pf7qAPmPhqO7V
TFNAdxpZEjiuC9Z4Cn0ifhf8tZm7ikTzppgRow886PlKP48+8OX4zf/7AHnvFOVkHfXkD2d0sd33
5+/z0Hq/hE3rgtS99lWh8Zj2zRzqS6pVW+A+AbnQ8Y2L8ICQZpj+onkFHY72bsxc86BsZNRt0MU/
1UpGDY2lPlhA7CtEmYkNBL87BA/QSMymllEXZiMK25qUV2DaSEHcLXgljw2e2v3lHxLactPzOKps
y5aAxc+/g2DH6oN9cyXCInlfjXW4U5LgA8F+qd7n72qfsTJgS+4eDW5MUJ0JewMU9Wb1tZWdh1rT
mZLztVKrduSnBdnAGhoMBAXpYSGkOFdKB6V4Odi3AhctKTcYLmsPrJM3NUI5gGYsoZpg2zZJhWzn
YJxuJ+fxcaVPVcdrp3cpuNytccXKXbm7GHMXVvNiXU2qYi6CAa8iL34ekmvtV9/Lp8yiisvWB3+q
OP/lgrWAqiEixX7A4ZYWXmX4WO2RBNmpR1QttbwiIqq5Gu/d2gA/pVWdYT7K0QBA5EaXTjVrR0Uz
0nHNJFhALcT9TOlsoSWVopPeoCGtI4BbeJgovALqPTk1/dx+C2PnHzjj7y2qVzl1hW7wasIuyTzq
wKbtaZ+W+jmFSwyIkei1FDLPNcUXX5Fq6kEJMfkkdEOpA0cNXf8d1kfLfoKKHnfnvXqeLRGqQfFh
7LoihH0QsQkF32QrPFoz8ByDNaKhvXkFmeFWmU56BkraARnyXhAUHauV2JCYuHzo8YXfRU0mUu+l
l721KStV6w4wBhASvQ0DU9inTI1qEHMNfBENCb3ehOzTAgHnLIvQifpxizpnOnM7bDPe2nUw50yb
zA1es0DTN+4+bha3JpV8NmlDw43yzco+psi7XnXg21l/NaeK1pHeeyHepvG98iIqlwjFDW3tACgR
XD/WZJqp4Uk6HzQF7uncu8quN0jxjMswKoBcJ9McvJWjbEexO7oocK07+cgxO9nePjumC05UuI2O
R273bA0Rg43F7MKXzAq7uNEE8ZRFzRKpHUsdoogmQ4ppbQZKHiTNVuSUlmra4ws97zXawzwtAaAW
PxfEyamyI2pNAToJnFi76MRU5KTdxO31nbSchUTlBGwluMBKyJR5AbIUzH+1RGQrMsOpRLC1YJcs
Rz1GcHjmYXb8oNrgjJqxXaz6ISXFqLb3NRlN+kQlMcGLVs9ZJSfnbZ9YvhHoAEPQpBy5eb8624Eu
wue8uffqdL7L9jRAjhO5cxdFjO89KIZjfE0o65rIeRaFF2QFJmNoM160mnU9P/GgpUKhjCnBq1hU
yEnk7tUr7ZNYNJfS8ntzz8tuN/s3eKPA2HuyPRsIkyrnS7myb161e4YVtmRPm2DyYXYdr2pdEmJC
5UiaQLLJJipvRoCLVABU9R/Xt6cqCW0JCOXsBK3KDTsagduvtVIdPQnAOksHO7eQExBWol4cDK2G
aE0I8uU2/zcc7dyNObwmIMk59PIUDgKtpulPPqi/+7UKMcBhuANmYAOhHBjQKpCOWgNnnoK07+BX
U0X6lLRDIV203ra/kRL98smr+3HQEqQz0wy2JAgED9s9d+PfRfGqZiwSvyCHmHNTzL4nJoT/d1rc
wvwTYn4PqEJBozr737Tv+i45u7mj+Bd18SBeZT5/43r3j8al2MVjk9GvLxFlBbjuO6GAg+/Ib2CF
DBq+DLxEn5kqRDSWX64WZmZgyESKEbAOOpcJ+zRc9ynhZtD54jqxNTsKdISbRYfx05yOKr6c1OJP
vPq8d6TM2OCpuf1pGNmnY9zXtHbt1famhZ+L0iYW/dKbHPUTDjwYfkK8muZ3BJTUVg97zYuf4b5K
QdS4CMlwXsrm2UnfI3Steg6MCZfOHIdksIMS163UEs/2yQ+h+24qr1+IILU988zRlKodgrEiXN7Y
jQ1xUAySUMuGBA2JaeOYi/NmZcF7JD5lDlsb9MikTH5DIEMfO9gb0sPiWzeJ87RNSGp3JnDGV+P4
VrH3WeP7JJrP1c+02SZ4K1C/PSPPU12gaZsjEY1Q9eLHfldZuB7aWU8uD16O52fSkr2LmSg+BFmq
kM+Frn7VpykA+2el8TcHkdlUs5cR3He/kOwqJ2JG4FbPPAWst/uLTsF2DhfiZD0v1f2WO3AZm9kC
sZ8JqXqGHRDOfV8zzIogUkLsm0q6HYBE/kRjHZs8esberrfjzq7NIzybTukKCBhl5HZdtDOO1AJJ
/O3bTn4RcEEEE3ZqBVePL6nCkFyrHVUNIqU3TG5/xT0cBk7PDd5tK7cSQkUYKv5TXY/rIiY9Ct0N
5KEkE+LX1Ww3taUCLxCy2cSkCuo0vGvqHJaPOgo7wOvdX0XM8xwS84lUmr71YdMCpHtVcAyZJ4BD
FDImT1ZeQdU08+osm5JUVS9l/e/xyUBVCMatoEHh8k1uCoKM93kIFv82DZvxjcqFtVugLRxffL2k
QzBbn9V4pvGBBJ6JuvX0k9msTFPzKoInxO2T9d0Xn35IgpIHj7O+iJJXbjwAcOZIusJ+aM8dMo6+
bW74LLMlMdg3gK0tmJsE288HthamyWwHmstFI2fa4BVMkYB7MEG3PM8ItAPkiHVjcXeEYf448G62
fqSyha7y69Bj1gvzAl60FJ5KurHyOtTGUGkMXIF1mmqNCYhhSZNECkj04XOgxh9fasuMijgBDpbM
JmVzolmDth6/5XFetii0kg/9ouQ17/bYtdyL9Cqp2v40gfSX/oq7pu5VnUGI5rY1hFHothLztQPF
pzt4Bi0s/sDSdMpqmMHoGJA74o3zTekhTRE1jNvkZ9Prg3FGpzQI7Doy6Y1qyQ/5bDo9D71NbCmN
JjbAOkxHrVoomi/3meajkikOKJKQ8/FsERkPDzGtrx7YtYtebO0lqESoGjuDyUVQ/tQd49hwX+F0
jrwrZUW5yJ8TTmafGUVLizNDC3ECFv8loUe8gaY0MmXiBgO3w1qI6hCgQgJyuvXwTQxmTZfzawCA
AsXgut8mLiAYLuE4cDNkWQ2TS+WAVb77ubH+m57YK0ArMC9bNPVwYFGkBL7TlddZ/inzwmfe60ws
P/D9on79S43emJTd/kDNL6nZyZyEnpIH7rSQAT8BQwCisD6dw+7FDLhuvr9OsaQW5XVtnjrxLaWs
LvXtMt/0n1Dzkvh5aOBgB9bcZR1WW6CtDpcRddVFG0A65pH/7SqK0Z5ib/Y+e1730+/2FOJu3Fhf
B7iefwXCUaeDNZhXJndfEXJlYEw+5PYXvHkmk6cLECDPKO5oZ7u+qS2BdcO8FgSCQhVTjhoLIC7U
viCTO+klMbu/kWkrr+Uo7k+3Hez+XGiSdH5niWbjk4z2Qo9uKOB6KebWiB0xO5Wk852IFzDF+DE0
vjXGBAHVSHHDx6eoaVOu0RWnivyYljld11JeND6X495FulciMXacpDf0WAthUEgeCyjVTIU+Zllo
qPEYdMWujdVeb9nehurqoxIP46WlXeE5oVzc2/hHvtLm+l2MIV+7r9pW+hxjoXjXKpGLuEXKfG1i
jibbd5xZUr1sYOHiZucseZrG4pD/sJhSwuqmcYZnVRQLCsU/Z+jLUmHOyKImJMCzN9OCwtOF5MiK
CpBoWTDH9NyNuoEq1AdlXxp15qL/vRFUR3k9PE7ilrM2LRko1qiPWc7V3sk/YVRIkcd11EEYzsKn
eXjI9jL7uyzk4yCmrFu1dqBwTqZfjnDLix6a2E7AeSjtuHFSveMT17Ppmd5dHzUg84VRy0pcBzAw
1sym9ysnSH/aA7xdqlZRkUvBSvvq65nsfUnaqGwjjq5g/jrI/5Y4g/bl9VSrlWyIeTRllxOuAP28
xW+XGa5Sarnplf443tlJ3cLcaB5a8aoSg+tyG6KP7F0ABVlIgmcfxhKm/O6z3nGxoLCdJE5zFVZ4
NU1TvM/HUmP0wMSolyz99M4BRsLhPa3cwuPP6RkhomqlhshyeB51CRF3XkLuijordHhUM/GGra0N
rloj8+Dp++HmPtAQ7XV28nh7sDykTtV04LqqPXbBJL/eKPwvra/Q1sCY3amuS/PSvTzQp/dMbJPs
FcmbqwxmBMVNNaZY+Acm8eFAD3JZ5VxRoYCjJoJERqxl8jUyS29YmIlxJ8DtHaW/wTtsziz1CI58
IIjHbD4FOe9rTMHVfcRNUY0+OrEZnn9+5emYGW3pJTzOQCTaVHPEXIDs4VXkuW0KYF4M6sLnQ1DC
6tla2Bf5xcVvaa4Q90wYUH7EAFmZNECSZG6glXzYv7YK8w7nx27xAlRyoz8DT5iUQcXix2y+0bnn
RflNUKEVpkAL1RYYXQWAUUUYrdeAncn12Pob0xnQ6VjWglTylQCCvg8jBAwm6ahSDBBDLaDUicvR
+dgMRgLFeTmPgCSmhxVS2yvFrQyN+TKZKR4io9TYA3PR01RmEbAhE10HP7XKXvKACaYrs0H/t0Pz
0sMT3iRyYtYA2Z110vEjuBTJCytKTqFHxYcY+E8dTNMXuYkuu3XgONbVfmDUXacuhtrJssx8jP6P
pMBjNcOx9otyuDOoyiOIoxvxCBxOBVVGQ80mIGB4ddme8hkxtdZXcu+L/TGT9XxELnnFEC4yJFXZ
XYZ8NiAVzSVTczjNJRYOIlO1NBZuUdKiCeM3uRh6iN8IJF6ZXy4hhQzbxmtZSpa8APmESv3g6i+S
TF7r7Sh+8Oih6w6ST75UiRthYfi4e/WdMbEj+rXbKPOzyKPvCmPBUs2GbZX5OBbt8H8RFngbGHqr
VD3ZMnPq1zKckI1A6J99caXrqfPKjuHHSZPRCt6+eJoj0/1lVOmrI8o5KnieLgMRIAHS9JTgvbRQ
PViIfLgnx3V4UdRIJ5OwPYtQ01o1erO7kLlVvf8Jd7eQrjpH+sSE68MlobcPEVmJqQ7ZHCD38XXL
umecwVuiQRsIXP5+DF8256F5LeAe/vDnj0i3C6EK3YaMQPqT4JBJP4QyJsxgUrMTrxcUl+fdpe9m
a3FrtqaVl9S4b7M7KNx5XoORnoespBokJ/g6SxP4lqaMsyPcJ+u8eom9s7I38eKs1gMAVANWF4I/
Td0CDr+4ABmbOdplmamLjyAMOLzQNtmbhvYM0N9CT5kW6+v5hA80qqahxa/OeDGX7+trJ79czv5Z
lYkUbGzsottZUUuKmlVOMllFSQZQ8+WUwQ3DcTXiYk583M4kfHMDaXfZYdm4gLWvanHXevd73g1H
89Ovzbw9ghVr+o/ckEnr4NSXHdit361wiHaPEgSC1q9QOu9zseUhp7SGreB2UCA4lqkgihyJHfSe
z9ZQWN1ZLmhPRSp7DyZYe6yQCklyjZFQ5lbEbnVi4lZMB2Twpl56CPZZ5pT0wt80pP+lSjUbgBIJ
OJqcN+82IBkQbJAGCeMRsZ2LoSyjBMYRwqZwUK29koolG89zDhgyHQnBXOhSYeHwN/6N3lzu2ABw
br/FQblVArJ6nBPKmzs2jCHf/WGsjBA5OOoLrSyniDyLkBnqsCtDsja4mjfdFauIqRSBuUU1tJlr
wjmmO1Kjzy6eCI7quObMrR9/pEUAyLDdzyiDXchoqkz2Ol74iyD1MwZRCRw/LAyTmF0SNL9LRHzN
JeVCzotVK3xdubPIhxyFdXS9wd+e2794dTwlb08Kp6x1GKv059Qr9Z7tUJ81RMVziyld32sdFeiY
Vv/K5b0E/ppUA9/OM5sJtMRcw+QA91N8syfOQfLev7YbsLqqfQ6HK0o3YREjqxwjT7wRgPc5m/Tl
0XWaMjXFWIrI6Fxrz6eRUsHCxNyeYoIGUqG8McxwETP6wBE+YxO7U1+ghIQx8ZGv3MZHm2XhmGXj
rxYgQ+rcNQH1sMcjw0GDgmq58NMqAgdeanttKR1j3ZlLDpi8N4I5o+HsCyBbALuEsewmOpWVeQoQ
APK9Ll3iStW1acWIhkUXdFMADkPETQuLCDahaUnVpKm3jaOk84JAOO7y0xKbajmXFxtQVB/08HEH
mrLw32CiHnASLNwNtMcKjmKWSSRFDchduHXu1Z82KnxBT7hfpIdgrdnx0cwrvK7lx7thbOLT2FDm
s5MPtIKaMK6sNe6SA+2/+pFOsbS0zbSPD8MtMW8gRDHYWE8FJsKymx4cJ10We3K+J/0UyiJ0V81Y
P32hYuC9yBR4Kbhj4uC7ZJdr+YsLkQYvByzxNb5TCdFoMHqBdMbttHRyY4xPGzT3pHzp9HcbsGxU
uT5wNlMm+UuEpHBNrJonwtDg+31p41lt+YUcFGA2NL2btnmLq/KUz3/0xksMjMKveD/qNFOXYq8y
jq8POh0vfADu4QNdYC/g545Nq7KeqBINz+SNmnITF/zN126H7GF4MTeZ0M+n9PiXZf4IQGWrd/IV
WZ3smaw0+7qXi+Ax0RbqbazxOIjz2F8E5ej7mRE6yb0tgzIA2l0EPhoo99CLnHtrqIGBWnSgNN4A
yQsAnkNikkRdkYRvr0jjiuffY74/3eFlo70W2MkwMsoBXKoYkIHq7srXgjr9G8jjXPtsrkz4guXJ
ddbvkAT82CoLsVAAaUjDdvsgUxb6of+GOp24gJi53Yyjxwhcpgni2viE6PQ5SnT3sFRhU8QHG8wI
KheOu1v32lU8G8VZsWegJ5MtDga0ZW3FnfgGM2l2QsEwqA/ubktJLSq5tVQ6jYd3ZHX0w38KEh8l
EHiLcr/5kmYnaQ1QwpNeljO3v0sOX0842TAn//8mpkRV/JLdqd4/Bw3o14+k58irrIxC7LVi9Drr
a9H/u30eigI/Dgquk7o48Jxwmf1Tz6vnqqGLL1I9JZj47tZPd7Vz8sxYy5MItOSiBB4usrh1Zibg
Mqq4+iQf+11dbBu4vtTy8HawjF9YPWv4yqdyz4DdwC8+jO6Vldoo1OKSoHx7N9Du2o6PWnRGoklC
V2DKh1Er45TGWtWspcRfa+IK5NOnACp7EttNimPHn/BfUe5jRE5hcFQFADh7t8OGSoXzKYeczwVx
nBfMryMAplEo7yFC8blxbucd+voY9IZfWJnDVPzh9tKORqSaaOA9xGy0oTJHSYIKSgXZ7EoRy4CL
+GTGQ3NbPqv+lMoyTU+xZ8p0+cjcqTS3hdtrXyc2KO4b/vQ3jKr9UQ+mwA83XIhuKtoXooRFUEgG
DRvKGxRV1G32Jg8hIIHbfWXQkyER1M8rMjP4D1OO69eLWx84AbXcAnznXFE02jJ4Klk9N2vC7Gh1
0R4fvPzks5Fczkt2J9Vmwcd55iASkQtWRxLHrXLIvVHkIp35govhqhnaz1sG+1nkQN2EMv1x7s1a
t2ShDeUC0nFEqxqc61vuMwmwjc93KNa9POTj+hWqAsXdad8xVuYnsDUp/XX6du3X0OJZk4jf/VLF
7WX/s/T2sHH/7YUkYY3VWPnQ4NHkSUuI5qg+GCfTRvuaOWlbxQrSNDOUTzaN+crSb3wx2SJT2PQ1
AAeXtv3V1da2U2tbjlyT7QgJEuwoeUyPH4MwlIEP3QT7puDQF5hVr8VhYWw+DYHLtoVJAWiAvrrB
795IKWVdCU2Lq9BxcTwndi2O6lUZ9Od/xrHHuaXpG1osvAyLRLW+g3Ufg3QJuemOttK77Eba9NNF
TD4zlKscfb6uHOA7qnc9Nokt7dB3tf2a4TlAbrhjIis4jVNxMzxt0CCs/8143g8kHf5EfksOzSl8
r35fLc1IB0FB/fjVLGZ3J5W5swtM9hy4d3JYaMM6cBPlYyHAs3/c0m2t6OBlRkElNvU1P3iMpUd2
fkqxubKqVlwKLAY2ipPzY+P89K0SsoXRGaqkLB3zpNMM76mqZ11YWZFPWdknQp2PQDoAVrNLvFRx
+GBW5WwLf9/9tjd6ib0YbSVSat0CS3Ii9s6Fjm3gCL38kll1wRwSPldmHe7/8N4SgbWEOO0p7gl3
ClU1O2u2dp9lCjIndbwknfyCIp3BdVu7fzt+EBMF6tHJeCW49eq8nkW8hnWTFVTWS3gs3ddiO09I
xpxOygt0JgJL1y+637l+62nbXyQCr52YNXiqqcuEHx1E9wMUKJtUu34a7GrEcgHEW2Mni5e4LnFA
wGMdF0TBVcgmdIIcl21sf1FxEBojJDQET3xdJqJEz2EAtWk5SM+7YynraA5IkqgrbdviXsGpFTBG
hPN5Y+UhPY3Xho+46HyITFRFlzLN9awsra93n1dOMSNxrNUJscE1XsDadROHQn1boS/NygL80m0i
9xuRCQH2FMvMRxjX5o6+RQxiBMhSJqKrQitxvpDAdp8crLhS9Paodm02Ebj9ddgNjR3AUZZZfbVv
NAxdCBpiU6YjgMDjnGn2cS7/DHO5zjUgFhxB/VU5YC4ZP/Xz0aZJhdtQJMAlKKSaijNGhCNk31yd
Yr6UFmD0zOQ+hc0iPOYydD7TCHvDRrgGzz+MkcuiArOfypi8SiMKkztVx1R4WtDz4/gyGAIuCcC1
MrzefaGHLlLhF/6dILS3oZuscfP6kbWk6bp8fNhCvsfV1SLmesYJN3haAHnlA7e/64Fzom1hRQ6J
JIoHihxDfqINWW81OnYDZ4l36/5BtkSgdvrEeEM1fJYmFruI6bNwI4BQP8uMP2ANPNHQJye6Y60X
yBhcS5v+SMajN4Q8/qlJnqOj47acpTCLHxgc1xNaIZ64OaBPDUvWlHnc8At37vUID/gLaqezz88e
Fu/fxbIWJewOCYUUW3c9V7ZSphhcsue7aXLt4z1TqpuetIAU1tYLQOy6ScIMCbnXv7drBggeYLfV
kcu+tJACBRFpTTn7UvjxNJuNVV9XaISWailfB9e6Vw780dd/yJtplMFTw+/eH63qskw+wU2dIw9T
6pd5WP0s+3875OkffzR+JfMccKbQ60otmZgWhXOwruxlgZyRmT1gPSVqXG7BGIBl42I05tlUb/Kf
HwIWm9FBKzN8NCMjVaAqfdgfAg1frPqhsV7xy4L7L7csi8jQQZC3C1elJo8O7b6h5a8P2RbGfJqd
ichWgSVIppjUucHqyW0mi+jwyBCitkyG04zujeEojDO9S7CUlyDaUCMqadT6dUdc6ea5BJfigoVV
aqQhx2xTiXRviZVlPe+cQs7WDCxsHpEvJ63qQajbOTBJs+Y3k+xBUOs7pTvfrEBQil4GbhlbE1gw
DM6PDpMTvFTThqObYirHCYHCuqnOKNQuoyet2ZaImu+/msR61JrqeQ66Xb2T37H1zwriI+S6rB2B
jPO0Mp+QkIPZeJQzy/YB30n5Hiv4WzrmgamXVRxC9gDFde49p1SB2uts+HozT0uDEF1uJD+kVYXl
jax5zhJtOyd78nD7U+L0VJg7cOS2jRoh8H6YYEkDvWzuAdnH9BiUy+mFIvkjk+4JNR2stPiFOgH6
AxBHqlAOjflc3BMHIO5KB2FQv8IADzupZM+nU/SFZ51+quAYd3KziZQMjDsytp+5J9pIlaRy00JH
op1NLqzwN6IUIG+GtVl2V+Vr9JeSydXVJBGW3hyTKHU6WDidd6l3nvRqzSqwebYsnrL7N77V1osM
EX7EUcka+omPDKBbsLi4ZpMx12j69fY1VOUO/bEFMrS5qT/JgsO1BSlEpQiSybLpjbDnKG7Q6zVU
vtujJvHnm4ludZZtkghi5HYkqUUjdnQu8FXVrxUhEBcMCfX69vVeUirXBYOwT1zJGJ0O57YNQJ/K
Z9CQSTmHECC7F27IiSfQ+copwq+U7kUr0/AZS3mOV7Nf7Sv9X0gTvxjJ3WsAEouC7U8qj1K1azxb
TRi56+G7yMFaHlx6fhFIDN0j8TzKFFJW0sskAVyUrvfsvPPaRqbKEjySHJxnlCFKz7dQ4huT3W8f
73IBW3xE4bJo8eFNGdpa9xV0POHSDl971PpT4YeWubHL/tUQuYEA13bhxNmUCVioKn/ma3QGntZU
W0+dxU5fhDFjfIFvwBVvwenGCJHquS0h3I+J/jy281ap6n1/vV0XJi/+kbQ1eFm/jxQP76FQajVR
hNlJverBxrctXiZUBd+CQYdLpB92B3TQuFSfYX23P7xHd9VPp80vjnh359zM5e+4LKrgcxJ38Dmh
3bwWaWnXqp41a3Njd7t1eeNUL3mIjPsFtf3cxOTgGhRhgzOtjKu4iwO/GhQxRIt3a38UDQlXKE+Z
KSHAhPtUTOHEoHALlcGeOqhuTgQP5ucdxsuT9Jw6Ao7HdEjZYfuxKOXocHKI8PQXJg3ny/2yLzQ4
glBn/JkFt0eRaozC6aa7FsKJOPy5sBoBmm9lkZqNrUnncwED0sbwtv+J36lC64XFupLHNc0B2K2c
xRu5sczHMu7O4Yv/A+o/0eUk2R1cM0zemrP3dTN8x/XZvpQukH7KbTF7s80g+q0rIWd5BHouaOSK
FTzwLZ+0ZZwH62V7mdYmyI2t/L8+2nqXWqwTPw1z1if8hb4oFSOaFh4Tq5cDc52F6R490oK9sSmz
KHs2qzpqXf6B/6Y4Xgp7Zeo72uA8IqBNAqltWUGu9RoG1G/dNXsHttk2fmRA7HoPdy+6ypgnJCac
Y3nGQi7epfonrNdQMhEtbFH+/d2ILRTaGUVaW8ey52zzMKKLk14xQdW2ArLP63I4tohgwwmh1jen
X+PXLmbyJ3dKquUj0BovsLBXnPZFbwvo2c4jTDXgQeSKLnu8Ni6eDdQ7IP8VxosyPcH8CnETGL6v
j8sjDjdp20twpBuqQDbSHGvHaUqBlXnbpAhuOMSo5zdEdu+VyMkRbQUNBuje5+qvoHaEIQuNeWck
3VJbnft0OsQikEGp8GFWjc5z0dpRb5E4y8nl5MR4hcRjS2aqFywUhJUHI4emxAncdVHKEFi9yGhe
omrQd+Thm2SpoGatb/lzTM9j2xo+4gl/BYY43zVRXWeGUMPuzy9Hx9TWQngJCQmxzfjAT2zK2l18
ECL2omoo7VO8jvc8IoiJmnDIreva2hOdDvZRfBb5+ylIaWnowYpsAHeOsZcS9ge3+PNr7ydgLAPq
VZEDyHnOp68Qf+/GXVxCu9DfsPJV4RKMi7yo9Se3oyOCjSSK9xsaDGF8lnGepQxG0poMqOZkCCrh
vcQn1GJ5q0xw6AtchDWme8Tc83IyQSaPGkFfvRwhQhmSezMXXsLvWVnAv3YXmO3Kg4fE9dZYRDDP
78hb1RjopoqOjzhF/l/ekVrKJbM7T1YMRA8NEw9s8VLTuNKUTABf7YsmDZeYSSUIQKwDqyUekMnH
QjGFq0JyXRvP9aQIzFrJN0wgoETJMhQs+jnXZ4hB2dYvEOsQzstgtW/1ne3Vt9+PfWgOHWeeBQrD
7+n22LJYCd2jkplQFXaCytPX04a/jaedzWkWrK23P0Bb0gI9Ju/X6oPS2VclOWtdZYayfzbfX0pk
XY+zXKNyp2qM+Bp6jeOucCItDwSdswSdDSCOR8efq/qD3CvblEo5FZLRg56i//O/hxrxtZBN+o/V
HOJm0cvOkQD2G8TLyR78MhpGMrL5FRvmxL/Wd3zUEzHKd6K7JX8vT/iX7PshDGu+AQvYv34Bz5OX
nmcsZmSvuTPIWv5Ka5mP08GWMkuh4OD1GINGCeBC8l+pFLzG1Je5U6prgBw+hkF/HtLNvRawTiG+
ZJnAutP9s6ccfNOlNGVd4SeVep9GLhle6eBS4ggd5vvT6CMEJnBdmrLwyk0Ts2Nxat4C+s/XN6D4
B1Lq79dar58uJob6YxvwyElHT5qJerheE05g0UfWwK1zx6v/DD6/c+lByMpViLFpwLa7Kmo5m/eN
sKjWfEzcX6xdgz0cLmQWV/+9Vf36uJIAkZCbOwdKihKaH2Xxmd5zHgv77Q2+9WXSvYSF8MoJXxGq
aHU/cgul5UolFHtpN6Gpat3CVbI3oj7GjHmZMNByCCjyc04A3glXWqW9ckVvdywJT0cTXJ9W3O1m
dNWC6Z3q48XiQtmFbl6xPFG2xN1+bWtlWj2xr/uch7/3wMpIZRyf+nHv+RU0AYqKzc7l3RSoiHu0
Fyd+45Bi6XIDxWfxjr79UuhfjSPQxkncO/HgfOvaI/7c++0uYlNuB1pndjDeC18GfpqU95NT3m0m
Dq9umDPIqg5ugSPRKs4rXkffvAKpQmgVM6WyD9x+o0H86T/GSAYm0Bdg0rlk6ShY48BUd6qtir/b
9KA/GAegcA6vAwhtwiIj00MRJ8DWY2yV3GfTs937uY0DBng0ozrzKgxe39hvsfc6pBl1OydNSj9k
Jyq6M5NleE4oJeVqVf1EQLYUBJUKkeSypeGoCbqUfUxhRQKkHaO0I6PVKjfcj1tm9gqsKnNprtzg
8pjUW3+wq518t3tsnXXBU1kV/RebhrWrk352LNqkgdARn/1rwmWP7t5Kg22lJM2nVr+J8fSaZ7rq
efGJndoHWEGp3/1wkWyIqa56+tuGiglHsJAdnqQ7DQ9sup54eFRX/gmaCCsX4gS1xaiCXOHsFNZt
RXueoolx92Db5wGuOPumz7Hz/d+yWmLXqjzJ2diliqFiSU5AZutjVz9Ai7LnTieMQ+mIyExpC34N
DPCzkGTakhXGMU62cvMPq32GQJIncd5nYtF0Tu+RlhK3fxUcY9CWEkhT+i784B9cmDqcrEGAPPJI
1NMj95sDlJATmQWW2sPfnLJGj64J8wJvzZexA0x3porqi1NqEK9YZX7zs1G4dsfxRAK1CZwfvdou
kGj6WUQQgwiAWL6w0S/TdLXhOaD8/2mxUUd5A0YlV4mrZ5AKRmjg52Q7d/3yojnm4neQsv/zBvhN
2BVnOuN20m8LKcWBnrYaY16bjoPrxt7kA0UooSx0KfEa6jfF+DoNsT3nLlZtiVNhYttfv7O3plUz
yAA4hxyILgrPD5y0K3JiuTI+zFHSMpqJdotE1bMy3RcG+TVybr58HaDipTTQI8LXyuQhUv8hbp83
vD3ITr2rXcucJ1vEY3sCDCPGCavG2yJx3uqPjp+BgLbDRqFRhujV1DTZyVvBMFlBUHl6zBvIV2Xt
sUxdL7p7IeRNg3mWbzwVIq6lg98kfWFwBiJp4ERbragIJgov8lenTbTzav1H+aH6z7XTN/oaM/U7
fIc1FANT/FKYI7Um4cGZPO5b0okyoD6lGrG+QU8P8YwndZbiOv+QXiLWVjROSryEMMrwacaVNigJ
td1dFPN7IkOeMOgPQdglW+KS2ClwlYhLljgjJ+HenYUJRW9eggm5epJf9w2dLwMRE2czKKhibMeg
HEknzOnFujsKKAhsQRmocEXjIFefW9n3eLuwvrgjccrolNs4tokEtlgwfZGSrBubEDWD0kAK1Uvl
4SCTy5AT9Wq3yj2MQM8dmt++er8OB8ni1zBvErlSi0sia7rVRu9h5YBDcIq8OEuk/8KuthBkYbSL
HOHfNF+H+dHxJv59Mtm+/OZaYkELh9J2tgqM3J0d2BeZ02FHR79miBxNk3kKAUzRP56R8A0LhAgC
4ROhfVUDxEcNS8AEKq5nyN2W5c5Xq1AQWbJzXHXJuoWNpvKJ6z/7ORFsADq+sOYAOXl7pWoslql8
Uoc/acagluxxtFKUcABW3uExKgDaAEKkPPO1tC70ITGTSxLWtwk0VzZb17TbTpuQXe0SZ996RPO9
RLza7cPGz+gMPJtN3hLuYKIHF4yUmgf/IqO7AGiztn6yuhxY4EbiNkCkUrQJIq68F3IH/eLITkFV
gV7AnBb8BO4LWEq3vx1Uj93uEp17dDbIBzja79V7y/yQl1fDCyXL8W+gcW9XJrii4PoXsntELhXB
blH9jUV8JBM93UNr4hF9MU3E6uW457xtolUzB27cMUiNS7PUcc39kI0NG5EqJBBHDYcP7kd7/J+2
EgXxkUmbNiDujihtkdmyqOtnDL928BXMcWusuYVmwppHXquKsKV/Wh7gnQDwDLJjQi4tIWL+RhjG
No5ozGum1cG7Th4VF/Dw7le9sIl9f/ZWqk6eUeJhhbxgh4EmyL+uaZ+V2GlRJy2Pex2i2xSYhL/l
b+mDaCWozINsM3Pz6zCPfCV6X/9bYHggk85SstiEfWPnj8Jb49GIH43PFwBChiJb+FgaL//9W5kQ
Adc2MHv1jo8R4QDPvp8i8gSzj9XnTB0n65xRgt0JYLusF85fCOwD8B5ydhSO+mDgLuH2133enwQL
fB78MnzQuSN0UM+zd165UG3R/usYCxd9vTW6GxQSxUi9lkuJ+2dDULB2iFNLxbOevl5oEbTGy2yQ
XHvqZcKIBeIV27evWQ5FKMLwAsLSdZx66wJ/kYkajNisumKTXZ3mhKRAiInKbtR6749lhRBygZOl
JjiLhfyAC6xYxD1skrvtn9tdb8nXGy0EZvVnR3T+vNSDKhGvIy4plBwslsmMw9LtO8bk6etKb3gJ
JrgBW0q30DmsYQ8Z4wo+BVRqFY2FjqzWKvbfQ+5n+4HEikYFpxWqmIw/RLWxkEKJekIH7nuOIWku
lmrfaRDA9PLZvIBOA8CyPMsv2UT/v3eCxE1MhiEoeYwKeD4R+ZdAloBecANzar3y4ceH2ObhQDID
Ow5CBFtRzuJYIOPCPFH+/E8HgzE0emw1yu+siOdL6gRiiQQZehczmwE4zxvzZmnS5n22QEZ95YFO
ojwuzbWHgsVJLBl4T2T7FEF4ld+79Bo8xsRDWU9W8wZ3Wzjvsylbrxj69FGcNmxxbgGXC8HF70Oc
p4Pu4YEQqMQoWK28w4c2/kPudiaDDl/val5cn3d/mezaufCkg3aEWaQomsx1nI2xntlzvwqPFLKj
NvpF7kVP9KCkoF05+Y1ajVL/7DbXM4u9gVS7g2Q15KG8s+3zV4PtkwbgAOwkjyKa+sETUiy8cHb5
yQOIgn6FfyZoxhuYZT+xWGEby+Gw3ZCZ2bnV3BtWrcNI4+jcTru9LYtKNsYePk1PQ50uc9I0Fxb9
TE9cCiAvarA8/f2xva9a2uCPeZ5BPa/mLsUB7aImctowbSsOT5fqc2AHCuYgTIj6YT8r6hAPhnIV
pmDOk+5McH2ZNDdW98gbqnQ6y2MNcRnqt4CanEugFDNTCIq+9OvmIa1/+UAcl1hZOmfBnUUz7LUw
FnEkT0xtYQjTBikIIpgWNqPt04tJZOUnrwDsDIj4tfkLGJ6hOWkqf9ex2HgQvLvyWTL4axi05tls
P340X9ELjmbqhtWK0tRAs/OhlpwYx30euIN5VcorzrqqD/c904ulBmU7EMgHlMcxT7c7jRwEEXv8
m5726SkXOPyPCgNWWVI0saZWO7UYzRVmBx6TZzM4SDoVvaF0Y/KkfxC/zVhQD3rmwf582KZ6xVQU
/XMKQn+hapIIGsfeykbN2RZ3WfsqWgcRj6fPQ0QPrTaIs8T/faOWSBYEbSPNHBfw2UarRwR/Ex2D
wpDMkxk0Rg2Zp+OvyxraCbfFIMYfjCsya5c/Vzaq1bFpZmvB7D0/LF4b/xhIKuswds7Iow4JTfy7
u0xS4zXuVgMm5xuJWI5seYvLnwSovHe5xB0T93zJE3phReKnc3oRS/m94Le90JnLHe2ZFcSHoJFP
Xzn/zYIRBGk17HkfvGt4BEc+9Y8nLkRnT1s2kwBeDw16qzsWczK9MKlQ7h+UYoVf1Lv2BZ1CNk/3
H/a+FOnwGoT/FOpCAZP4i5IxbzGnMdZ06T0lpKJU+qK7XgD1odsxs8LVmd30VcyjrSkbj65NkaPi
4CGREIgIxOZCEEO9HX9hx7figI2KDABd9X+NB643AzNPjamlA9EhNd5WsW9J17/ENleX528wJAk6
0KX3SN5MOYQJGGF7h4je3V/Xze9JniRK1NQYVy7KAa7aEZ0IUPMw4P+K2UwLg0GmmEqi7aktnoZY
cCo5sndPigKUDAOsH8x/S1p5jZs18H+h5jB+m1i2Y1JzA7stEPedQhjBTD10egqydlRuwPr1YJFL
yiLBkskObiBXPwu1xe5ES7uT+MTmeOOrMIP7ewo8ea+7TRrgbAyfTgRPHoj0D2joNjydwX7H87f9
Nr0RT52aH3ZZWo6DUrGf6wR9R5pPxerP94AZdmGyyPD6ygfoZrVc+rzA/Gn4mJc2osEbZiFIt8QG
Qc+Z5W1XSE4GuSUjmA4lfNfJbH24/VehiEBKZdaiquRakNlDhl9J6wsCSitealqCVd2eCJFhCT3E
BLx/qXkNS8k/61IOTzHooGi7viOAEb4FBafOymroPtn1AHf9oVrZ9ihI9rP6sfJAxnV4QKAjRdnX
Czm2RQiBZhX58Kygaib7GI264Rfo6aRHRehPiZrWgnDd0H4+cuL68eaZX6ZvjQF5kX86nTSXaqZS
SgzLZcnyYlEgskQiP3WZmkr0Vho1jWb19+WD+9w1VwWvurcoUrQNuPKTKI7eGvBVtEeR+OrlnyQQ
w9/76LfOa62cjCTJ1Sx/1rC+6WrW1ioQyoL5As/PUiAI02MkIs4pkvFkUsJyeJfWARfEWZKAxGoW
n41MrFouAfXy8/t7QTA+Ic7gxALh9ujPHG54vUpJ+Pnptu9GEO0mAgLU6JNJz5U+w1HBBiCXLTXv
AeTQL8UNuVH3UXBb6rHQdk7v4U/TA03LOKNa14GxvkfhwZAXASeZtNhJfjhTz49L4z7yQTEB/dIb
BLbyw1qFfb2eQzpcuu8ZaVZqzBdAc77+XoTaEF2n0NS9Jb2WOzyZDEFlD23W7b1wzFJ6L3k9PnlU
lyemK+NVq5JZQ2Vwhc95tka2vt7qr7hC1HGyCIUwCwINK2eNPcVBs3N5mXShnTmH7keIoZNSQm9Z
u6uWzNGjdwKBlrLVZK5hFuVA9nAOOakw1TMXJCs9MauwySmsaV/R0gw/GWGy7m4XGseh/plz7Pp3
wNITUY3vLvn0yYS4mJJu57cz0Ypz+kINrZmrZuCI44WO5zhfP9bY4eXFOAcQZEpRUyQwb3bP0Q4r
sfJXEYcRhMR6zV9uiWDQ5JFn3/3y0XR8KOoQTtGfEmWjuMuTl916UBbna6OaF5f3AdCGrpLzoaAk
9uzkrt9MrjaI7zuJ+Tq52C3gM7O/AVGF3H/HteXGTeWQacq682xvka+GcmoZ14LA6L9Xqb2Pyp8U
Dq0SWf4cIym5iNy1PzPSYpviLI4f0MQc4XjKnSomLvK7e6wW2D0mxTVroGrU+Ngzd7CD1VJtWAE1
uIKfub+u8LnpEZH4CrVBQvzVQwMp7m26ygJTXv0SbC1nMFqyHbPdwYEeO6xFWuMUHuzomQUBm6CD
Hol9vD94aZ39dYfh2/SB9t2n2cSK0zRGW1QB0kpcxEi3rzn0sZ6GQRZwmTxLEHa0RO3it7+3qO2y
B6mhxcer24AyrSxumvVP66HTERtRNxkYR6DK57Qo/Leq5mUmv35WuA5vYYJ4FqsGoJRNTc+Kdk3x
Nf6ptZO/BjcVvOJIlhoQ4J4xzevnZayLQTwgS6inXs70u2jE2PMl2etcz4EwZVKzqBxy4lDgBb3j
Z8Dnp+JQzFYq/GzcmvQWxLEhLQ/LRrBLPSTvZy9NYFHS+FCWoFO8+FsiIKQBjnSF07QrxtCVFH30
gv16sLBc5WZA3Pz37j2rJeemUDnaBi7ZYCt7ztTpvRFr45XTFyDyC12g57LDQP3gAduL2EGtO/yC
TPeH2VXdZV6urChCKkyz9oCvmK+TTqtqUvI86pLqu6IPWPJwirxy2t+hwZ+RY41e7lCr/zXwod3Z
DfwHpwrkgBElLchgDaHS7i2A3N+95Srl5iZxtnVA8BPUmg1aEYAMDHbfA+SBTAuT+RmdwWfwVhVm
C1oc9cVMUClUQkwMKTxMmWGDstdBYqQWB6HS+fhJ+cTsEWtblvPf3IxrRCg+VhDlYnOhHzYSgaSk
Y6NhuzWJzYYD5TjjAfrAw50HxQ+1XJdDQ2Uv8GOcN7HUt/14ACK+FVfx4ydgw4JTPfSJ3889blcK
qPzLWBuYPDcU+U9udgLMalmq0Fw7/8iok6egZKMZdKcV5BWn4GQSkgQAgc+cE1TbRj4lgKY/bzye
A0EVJK2QbUlJN8tR/5YQ/LXUwEI0tESHH+cyuvptwVijfYlUcaqM49abYI6rf4VLP8I0NS/mnQYk
M03pjeOafVaXHRYhOmeyi52j7Ml/aipk+/JLn2W+pjV5UzKSjNZFJbwsjPk2Z29Ac6tn6maUheh+
o9HAs76GeulMnnL05MOQQIBuLd8hMnm9Knvf/YeRdyUuWAYhFkuebTxd53jD5JeZXep3tNDCh6hp
XzDoo/NDAmrEAWz/f6w6Ab9ixGr1loaoiB4yS18ym3ypkEGJ4YRChjmtuNsGyBMebXPdt6Vgc2eK
pIuqHTKdef3Km5hYarFvT+wJAemGUFno9s1mUMNOYhJLrQ8DcD8OoLE32fh9RJc4IRIWs9gdM58D
cJA8RD7k8SpFPCKNvZ+KDJ+tfQuS4nkjVhevTRimgCOB3I/dAX7q8v5RI3bo50YljfpaMi3/m0Nl
9D/j/lamexm/y1vXdF+RBfFXHdmO93VLgF/QyVnlzUZbUMrVbOqnpLWIjpye35McommSrAXJ+Ibu
/Y0YCESxvzWncErFKILjCjvWRdPEozppWlI60i0QUfOKhgPhcgc40DCdXvCbaaU1YrBoJZJErsWa
SNqwK0oY6P56tIKbBN1u6xl7wPScWwmGZPGeu3vUAidVPnnlSWqmLAaDX6rG6XMlt886I+IvvO+G
4C9fNG+Js3Ac5APZJmHiHx3XObUah8/ulwhW6/VDTzYhNXpOpFTeRg8GTCy1jAObsNMjH908Vi2Y
4yRNhnPP7dOvqPm0b/fT1GhhkCl3knbtyQPn9+EEuWToCA6U/kItUX/zqRZKiCoEZmVEJ5V1ejUG
ybypYPzSN2oi4IQmvEasLQc6lmzPN8l0YB9TegCxSGYEmM8DrSz5Zjwbc3nVgvki6wQoIhoRQHgF
JA2TQN2iQTjZGvNH019FMj8hZfUxtJpYK/2AQYP+dlxGydEJKNxZpQ8LNg7sADvyBRbsGoFL1VOj
iLd9onbNybvk/DmeG+bfmRCx4e4WMw7K4qFwC/RY5ErqWPdnyvsQum+oCtzQyn9HNvU/SC+EITF2
DcbuSnteGhoELlpFu+G4v66/Mhv/MbyeeD5uBQ9GCiZ6ILZ2SrMH1eOoAdgdx/wIK1KTXmpT4Nsp
nfTi80BGPrHQ4IBZ85glDCyUYLmsmQRVCa2IAx710KukY6RlLpNoasTi5Bsf/dDR//r1aNdpnSfP
BTuOMgnziCIv7IU=
`protect end_protected
