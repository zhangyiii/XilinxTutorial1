`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11024)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aPkk/LZprZljgyNzZTGF6gcxBz
LkEl/7f+3dcASD/i/Kj5BrGQGPFMOaSER1KNI3/Xy6RfrRHeinXj1OOMbIk/XK3jgKYTEB4PSsmF
kBxAwdQHO5XLcGW2pxh8ugTvfgYrlkplKX6K63PDLwoObcbElxgs0dYjbCJlyPCXRKjmX6i9uJbY
o9V8g44g93Lh4YefdooX6xBFh3q5N2ufrIx7ZBMmeDwHM3pHXFGpSnPeaewhEVlo3ZZRAHMplCs7
HYczUOpHyELzFE6XAvTaAOZsfyv6SnaaJN7kS5RgkbuHh25B/+zMA0pgCEQ4TQiq1QE7u4X75q9p
yhfMKgFbZ9Q/BhToJfCMM5PYBZDpYS1uKtaYJqOJHpy9r2deMLa27mXn6SF7My9WhbaeKTDT+HdD
52JtvQIDr95WBS+OSfTl6Jtpqrn0I3VNTDaSa4fIpkU1Mgi+HZFoLjXvkkdmNEhynKBKVBf4nzfx
Rhlen3GsBpRFBmmj0xwQAdctFiGIQqvKcaTymqqpaYBk99lrROFC89thgHnZoVDcLzj9yYq2oJMJ
Ydvxb6cRkAcI9qYMnxIK1wAfxBlB0edB2HAwGWVqxVGvb/lE63FlTpztHC5fMpyuknaPa3mho3sP
J0N5ThVov7fQh0Ll9/uLeo88gmqgWlf6s/p8WvgDKF1BM2OSgZNrh99PXXeq76sYm5yhq+7jaoSl
pYnMVzIqWP7EJj+4QkfUKG2m/IaFWmIQcfGVheAYKk2VXYmJW0E3k80D6K41iSYRSqJ+pvl9ED+j
bbw2ZvJyKBTkfH7a9xNXhdHdQ0Osek2HkHMVQL4gx2G5cfuCgAV2IoJqB8ZIpSO4ykJDn2YlbCb7
bXYOCxuB3l9hbWrMt+Yy3lXhPSUWysP0Gl5LCpn2HfhADaL5NDDzLR9t/tAkxx3DNRcXlvPtI4If
nFHXm/iBulWTUCgyRrE6nfuTbmS+2e7QuiBcjfLwvStiGbzXaHRm7yoI8Xc5Ojc04M+TkyKTj6CT
NpoTw9RJomn7B+Ag28cKFrVvtAssNsOHbt/4i+DfDpGqLsSiE7gjTmWKk5YeE6BOngYrkSumDO2+
Gr5jzpncXFQJOucYsQbiq43cszv6bdLBrqtgZ3Ip3QP5pylxHTRD7BmGB6f5kKZeX1kNE/e5Pfxo
jDKoofnO8LF6MdpLr27dijNhbHxWSIB2F3uAaTaRah7j3t1tpGGkl441Fs4bFSd6CwPOZNn1YQLz
QltBsffaUG8MlVTTshYYwR/pGdVqN8g0aHj75XGOetVUhH0549Qoou3FhYpBMBoHUzdZBamB+4x/
Cvx96UNtiSjafRQ4dQ5Onkt+i2G72Nkq+3BuflvVCQ7WXgTRHHmjUV1KN3BkHWGWcZQzl+VQeVaj
5X3u4vAT3Lyyj72t1y3UoGAEZqvLwXgu47dlMkDYKz71T0Bt7g7PK3GphV/QA3FUUvP5h7yyD1z6
1OnDjwB1hlEol7AdpXCpkYepxvgeg6pQB3/YcVsODutWwvapnMKip9za8Bt0Dvf5s+K90Y4joc+x
TtrnQ2X9uSKUxz86+mH0A9n7Kbw36nckFAvx/Q6CYVo5oe7E6QjccdVVRecnLmdBSoktcvMckcdx
a0McoHfUvlAF70QPGQiz45aFoiaEknJ09BL/oqUP0QAJ2PYKOrdtvqwfYoxzQh0F+4aWLhJ65pmq
eoE9eyEHmdwZyiPFgaoGrJznQRQleUs3c4TphZEcz1t2KwVuITngodVS8EZoRvpuXXloz8DGfOUf
82t1QZhG0S5iV1OVPl33vLPyq2O3ms2AkoYvjaZph10tCYZRBFDo7vH/yrp/wQ+vG0CSZ6yUrGnw
5y/TJlNLmU1WWTkIGyYn7lP/akhWMx8KrsmFNpi3rIf3hOvmRx9eeX554Ga5zg/Yss9NFuNA1HT0
7/UZ1Xp/djj55Q1oT1PGPtU5Kt5jq0HOA9jKhjorTAnYScI48rRGmNKjVt3J+08Ahj6L0emFJkzD
NRywE3cBEZJ9Rp6CIwmUZcqFTfFrsIWwra7snDVOg8odXNAZRk4nURDZGsfHCBbgRQGzxN9a2JzX
NE6TjjgrTA/NlTKw++uLKfZGVGQgt431+wVTpgP3d+jGRgbiW5Y2fK/Godg/4dQVQS2wnfbZzBVb
S1FvWHW9L0wjr0opUhJLIV0PDTbe/YfqLqHzyQfR/xMr3D3ZXrEvUsznDEM0p/a41VOhLcpM4CtX
1pXF4drdvDxnQlTrQJmyRnT1y7z1rwmUWTXcMS8bvULgkFvyZAHgNd6xPP0YfnXt0nQJyhfeA7Mm
wx6AsuXRaLA7F1FzJ5h6pz6O8BqE97KBsxNYz5KBgGpzFbeZjbjc/EvD1hGfvJjmbApYUPbDbN55
WIF3Lm2VtgFFvTFG7R5ASfV27ZB4gQ6Tsto61GFBEfrySX3GRt0oCcXl0REwYXq1f/4BsQr/bUgI
SJokoNVDin1FwdvW0Lt1aTSDqZ2Ds4lFcfmlYwD+CARNIKDrw8wD3DRl4u3UT52o/q8AKROrcxTX
fCSYad1+M7tesle9SMaEFO+xAKJn8bz87D5vbiExjgfrV2ABhLGNcN+ueubrwRLQqC+4TITHP+OU
SN4oGjkoslywrOsG3xU4IvFP9xpiFuOTOId+X3+342xUklbrqUljjf5OwMp1UhOE0flSkYip7jEL
tAdzC22vnQuCIv3WSDwZNfP4PCFFVEGwMpUYcp2SbmlMoOpc2DtHQingSO4TjJncSHRppOZHPQVX
X02bi5Jkgu3s+5XJ+D3XgK/+XXPbqAbOEX1Pj/Jg754wGhHqKUXYTf205VjPPHf9ti9ixSHbIRr0
6y/TgktEq9GZ9DyHUQfhTRf66g9ywAsNnT3VOLt5XNJrzhfZWU8NOLVOm/uq1kMkIYIJ4z+2z1iA
sD3AcLmmmYaXsx78kw7WbQwu4QHvlVH2zSES7k81EXyKULFcyf/56Trd7DFbHEJ+z4p1fK+5Xw5K
jGlqoKaJfgC71rzOS7LUaqIZmOr1HOLvBrrtV/fX2XbsKxiSAfBCC/MQyvZ1oji49llkNV76KW4/
HnsTfX30VeDb5vkZ0hInX9bYPulGgZFDBfzTdqyh521SXAGwg993BkapjFzf3oTTsZOV7iJ6xv1H
RnU7G2DCB8+Tdl3zS7PmYdTFh3/ZDoACtLeCIvTfYMzIxUXWw9bjqOV/PJ+FB8+rWPJbmcwKEsmI
dTnEasv5fOe2Tp4BkEDLxR/d0Cvx/3vJERb9nIF0rh6i5beh3mG0AWxEr/MR/9r7WmJPGdkrGfl0
PgaDTN9R4c7FeL15Se3TqkpkgyyvPHMHbj0bDNj7BBAsQ2sTy4rB3CTmgSsM9xrzUf2NpLrT8DwY
AKK7ST5Wvp/Hee+F4HutTtcY9fwqkZJeisvvpgTRdFBkKXLtaxjt2PwupHlvnSK+bEF2Y2A+c0w4
68AJwBrVJwHaPI4Z6oXPL3apvjJB/08l9K44fcfRWM4ZExQ/v5GUvuzjE0ekH3euwAjlrhZ/rJR3
+qsuomyNNGbxUO7X7HmFYlBx6lhzMdM3c5cldbicg/Veyq4il+9kdU8cmelixdiiHnW2ZPNDhMRo
B9Q/g4pw8WLyoX3xquTeg/f6GQbWVeKohTUu8fAgIys5OdZbGI1y3R/TkHxPjCeoA9GmFESIuAU8
10oODXnvdklS+YcxyrsWLmwOWWRtY9x7jhCArPSdtXIxKvONnkZUYx02OZyV9UIQwj4B24Q0TJz+
JkFIXW6QO3g8PaAfoxHzOGRX40/QJXHJyuR/CgwmS2csOoxWVTA2l+lFYL7O+5g26hENzGL8g6eH
VD1bjXqip0NfJGK9oPKI7YFTxur0/4BQtun5PeiOFenBW+iJrf7CZ5RHhu90vxz5HDm8siUFuLuN
+m5qmVM8KsYKx9nrdiJcY2Bj5rmXsUNFRnxdgKvtsA1EVFidswPhpUTNxVX97/ciZF0UpQEo21TW
8RCN4TmWlawsu0Hgztts+wkVDhKA64SG5hBYvKPuJyI4ZrrGFdGjkynY2inm8twstc13Xhd8/GAx
t4XjLqRptHXnbvD8jvNcOo3lTSYTBbeCwGWMod3/rBCESNSMqHeaOgTVN6+QAJDQlUxtIDeauC/Z
+G2hzW0P5cxxq5V8N51N8z3wdf9QpIAzP5f2vRB8671cd0OJbaEMcsY49CuJe23VANX7ofNtI1Aq
535N/ygMxgxgmWu+4WD+lxxHVL7q+LZ95V34T8brBQ9LB0F+cSy+af7OIXIJT7Yp/Xj+RfU2mCnU
SuZs0jw8lYSem0sO7biScpmO4uTsGLChy4hGgkBbcItuq3rcV1J3Dqethdz0RoDCn+FeZD/NVUPy
RzFMyUC/ZSPnGX4+U0s7McWtIonTjTZqxh/OOcdLNz5WksYTT9vrH5N70gdj1Iga0thf+07nLnyV
LgUePx9Lpl0G45pxCzJheNudUyRTP45HINLNQGJm8Ap+Cv82YRSYumDKPtcyT2IGoQBNE5hNKZcL
bRRIilkOraxvplXcn1cVpezosZbRvkRmkWufnL6Ccn3itbxe0bs5DJNya7d+WMLsLvlTpWNmIekG
4ercaQR7i+UWSChJX/baGvMSr3j4/fU77mziSP7jj6OAo9qB6/DEGjwOGg79B2x6YKl0PBqHP/e8
WGJubozwZ7vszBmgn17MiBlGylIB6wLnshkBk9ecQ0oP2VXTA54hm7JVoEUaYkHMw6KDnm/MiXIq
50OblqGmN4xM66gGvCsVhCguZ9+0CKgQsYzWQ3N1wO8i4+pdxiQ1ifShEt4l6J4oV9TjtgoC2LBM
jVNEYU3dMYfrqsYPkzTP3RGG2qkKpoUgXZzgd/ZPGahMYwkUWR+QyGK/WZyemPRYAAsGNaAsfdOe
k4UWL39j2tt107TrVuiWLAADafQUUXn4MTOw/BbXsxZJehCSdQ1ZLpbdvjFMQuZ4RqvvmwPDv7uB
Pr8SacPPmXN1sjCoYHDEkxSzbtEQvqA3ObAzD2YQKok5xqlPe5+4V7JmYm1cfmm9VW8UI/GuhZx/
yTOk5r+DPWom5QdU9tktGTr6bSQXaIZuEg7riEFiulSFX0m5lEmsFc2BhT89mgOWyOIH1Xx7vx6g
AlCS/tC5ZrvWRREogD2wG/dnfEjEIIeXBlpbsqbqmHa9aD6E2YedeSGdB2Zt3sqY0BzuCh8PBkqo
e48A/mb3zkxEpuZGlOMxFRz3UjiAzd08stORLfNSus25soSWmu4doiZ2AyU4VXb4tr+diLSGm+5F
p+iOdEbI1fazKvl5ara7HQWy+Cw+BtZUWO0n2jbqoR1/ktASMxj1PtrJtxrovY5r0fcenLPGj7H3
CDQ1VEN4df+YZC1U/3hjOOKiIUfrnW+3hDK8pq8vdDUt1QqekYJOvloj4m0xqQf5glpS7blyduEP
G1/MYunp6QqycAV5q7o+5+X3KyF/PBUzNmwKbPIkuUseVNPW/ziffX9KWQi3VKUPTD1y7vZUWdEw
no0FdVfW++wa/jIMOeEe86aDa8HbStaiJOWCwOBEzU+36miX1grWc2xy8Xh3rJqa3DROj8RpOTN+
qOs0Wb/llVgEailuFsxv9Kp9iX+gvN8pmcRtVBFfimrA1IEMoePnHu7cawhqkoYeielBx71ddkMG
2vZPin/DRHupqFK2D45BQm9JmNL7fZ3Dy+HmJPU60lTQdv3REtsYiBiR4cCSG0o2PeoTvNQQxQw6
wzqx2Ffz3w1iPYuxiTAvNvcgbcF986I2SxlYZzir3yGYb7esqjrU6pdre/LWtr5tjUDj/s4Jg9bt
dZz/pD7C4dxzLvV6KSR3qvzmSCN2DARvQ1H6j/Fsf9LvLHMc6zVmDBA/XATiNdNuy/F0iS+L0Yym
/nbM0ePI9pabMxaNrIQNGSM4gExiAZqPz3+ws2R/gYkjbiZj0RXei/jk+o98tSQPHrhYZMFyd3aK
FCLi8OjPmIEMYZ+pYi3eQBskax1/TuOkMmes/8oQXv3xn56KF6tpMag15VSXJPnqg09zQyF/cgQ7
WMMKazdeMx6uK8vUvWKQmZ+4VKs5k3+ttuC3EDJsqJpUsPRLKl8wxHB6jBYaSDI4p4t+sz+J+enH
RcOCVePa7X1Z44oM+6OS1ikrA79/2SCz3VPHKvSoeaHcX0qsG5Y1ibJ9E4BQNOy8UDogbhcr1j1F
a02S5wasNFK/OARzTT1AEHZHiqrfdEp1BFF7Zi/JERXfmrLDvgtTMzAasudEwXo0jJ9w+k8Caxa9
ROzUVbiXj5SkR2wkLlePfN1w1dKTb7NT9fAb29B1G75Q0Tx4szS5AKlX5oLswjZ3tr1t3rctX1a8
s6c071+CDJrnC6fAo8deQ8pF1haDSQbv4glwCrSkcskagOU+6bHUOKSGy0MjF2tqZSGXjVt0wXgZ
uL9jSJlcM9coodPnZAeg4FLeDX8JNCPg828x2h+AgNNOKR979dbosJlLMvd65ic43rwQI2M9zgR4
uMzH+JwWkQeVRX6IpUq6nKLRT8zW+xJslhWiO11ATwYu3nGn0M19aoGkpPGKv4YqUtgwijBKBBxo
1Rx7Pbo6Uybiu5AB36K8jtQhPbVtsg0eFEFlCQQwJvkL+QKd9v3C+YN1s/ZtRfpuS0ml1e3L0b7m
ok03mgD5BP9PWzbaMxwZk76cf9O/yuxWYgU+tMtyfZvghBLZhEZEMH4moQNOXybXpeLQrrf86j2s
CU8bhCVZQiI3H3B3zpHsWAwJ6f0zLNTEZuuk7msVVYViDWSIxyEOMBwGwdmlwCgFBk8xS1ehu5LD
HRGNi7IJYk/DfHhNovt/WiRxLiJDpXgJtTGHY2VDk6qBuVeRVBXsj1gObb+DEb93CUfKpRmJb4zN
NhDxx7908QUSMBUUWqDhnTpGk6K5Yx0yShTWpwEfJSR/y3Devd3AYoE+E22EXEin5XLvJDwLxT6f
IoQXSy24C1u2tsjOCexOjZPbHPtgU6Qi0WdrJL/bGfyDz4cqWf+IEuzHrAcrJ9OLfogwlg45h1kQ
xuklZxx1UgpRpZjDvgB54A/aVTW/Jzm6ovDpdE52HCQjFKbGlWwpXJsEnQgp9t02aQRJydQSs8rA
3Ks33DmYHO97jAeheGqhTkpcQxTO3jsW+8yKOEVcFKLrelh8JVrq256Aeng39fTaa/sz5eBeUAhw
XzoAVh7Yl0ed4SR58pD0vtuvAbpV/4GI0VY7LkfDDd++CjAngjCs80Ugrn/90yp+FmAaGO9HK8xS
ZXoLf48JgZ5wkn4ElqFfCw5EB5gjPbJD3IvrXW/oa8sTxi5+Ppa3xzvJGooJ6AHaMs40M+qfPcnq
115FI810uR3uu4mON/YwrHw9Dgq89EYPO9dQJec4ZFoUKeq+jWrxmesE/Wy5oePkcdu1+dkN16tj
ktO74XB8vd9BgT2GrFqol9au2TM+QXba43Q2ybzrIKvkIT1nZ/ZskPqbo4v3TLrGRAhDVueq6IN9
25boz+PmCPMdH7yXnXp8NwKy14CJ8/NeGezq6pjAVG8VaDjApPNlw1tFXiLUbnyr3IjBUSvpB46j
Hw8WyBtH5eefquSAyDazFKiBZe8rnGIZakAvGedwhdj8MCtKQzwX4cLfQYD9Cags+tGAeRVLE7zX
B3sgwMz02R1zBqZE3fffDsuUk8QID/M7s8AjvdMeFQ8I+UvZ/jzMm9iYzflCVHUmII7putvI8QBP
PIRrmAYcvhhvNC9v2gDqizS5qER+mlDMNW1x82lXZRYwXzAKrYomQj315d1qcep/4+kwk5WgiI/X
giVK1EpdLwKUG3oK6SOeIUJItTR4sZpk5lPLndsmfOXb6BghU233Jj0elaybZ2wXRC6L/dx9YZqb
oDsROWikqE62prWzLjYrPxDpk9T7vyFH9oMQd4B207PFNWumMU3VoRcL1r9YmVgGFAltnO6xVEqS
wpVJeabmzU6ZakjTqa9qJgFaZAQZRNx0iZ36Kxg6a+X2Pl3YpI2JMRsUeQJgIBYkamVSD78AC/B0
FzA1NKU+stGCmHPbKWKEMfy3H/ShSnhEX5zxPN3nKDf7xrBFxU4GFOofwHttj34Hd9NpUo/FjQTy
8ouMB6wiRGjEy8jr37fBVButzyNwIyuCKQQ4WRUWH5D1zazYvOsvxI9ZakrJpyzDyEDJ4v7R65GA
0nZImhoQSJp97HkoMoJy5+gICwna7z3yJxx0jo7XiyN9WG6VHJGgGnimMK/hOu+6Yvk3CneOH4j+
VxkaeqIja46zDl2RlwjuHifu1zLPlExJtTo4SyoMHDOjj6uW/5GmCXRLAVPvIPwvaLqw2lCS/NA3
Z1/VGHdr2X2RbxCetqrUH1GHKoSkzLAiQFHOylgxlLnOgiPwX+YQl2vE+62ThpykNiMlcpyg+ZRR
T2636Nieso76Yc6t3VSXjQdTdsoFqajULGkbGEaEK17JIMnV5AqyMX5DrUn2TxedFw5ybUGz9rMz
z4T8YTNNfDZYTsNtKqopfa6+/TyAh1HOa6eKkNNToQ4kAISlHNBZWfMGDiFg5JgHtQWzvgZjxk4k
uccvkVVDLuOKTJUKBeHz/NRJitamP+f1FxmaTtG1tcSPfpuKB3b1h4E8Ubm0Et6Jus8ibJXBEwMW
sEgaIkfL7cR5o3Gg3VPNW12FbP9wDvPgH1Fv/IP3AFyLVviLrMGbZWvE/Cs6otVHC/i570AVTCT+
XNuujGagVN4e4R5NJm+ljvacQjgEcHc3VH5xPa1w8A46g7kl1LTJzsJdmJ1nV+piZWY0fIYH9Fmp
ETs2e/pfWFYfzdcNz1RotYdh5zkhKD1ubRFhfKd51LPXf1Qzqn6FbuM78BCV0LCfypIFIITJ3Mp+
Pp4OyvoJepW09YruhAn+siNdCC/OOSA6s8CIDuIGREg5RVTKuAZsa/XmcHiKq9NNqjd07y5CAyz6
jLtKRsm01IRd51o9B0l89jDPxyBnLXCKBPF3TgzDIGqR0A2cF8CCOhEgbHJCvEq30HY52PpDRxcR
gCVl5GH7qZSBga+psbyMNS4gj9UyZ+f9JLxlQ1XJRN6QSFFZ5b/p5plWxhNq3EimAI1Dp+EYtyzG
+jAFuq0sv06AxrKSg8HZBMcWSSTCp7SD52tcIOnS5Zpj8qvILuHCD2ZEBmn/5y6TuanHfHBN/ql1
G2GNK6Vt0gpeSnAUXgFJoSsjYWRl6cX7qRZtvXBeH4xOmMOJDQdkaev06p3T7r973PBqaA8aJ5GS
xHUkiNsoOUYPa1HrDZ6tp29Nv+jF2YnhLvdFrrkq/EGrcVM4Hp3gsx8npTw2CuzokanUBCAlb73k
r9qRlE+nwCcGksGaJp+jVwb4LGEnqh/WedkvWWvfni7ohczcmQgAZEfrQALzI1GmlksfinNABuD9
ZCy/04rVK9oyL+jC0WFNihv8GJKPo6MuzNlGVKZbDh0hAZfLJsFnfX1O3DYI0Hib0qTwltXADIL6
xZZY8Q6RYyVQW4dnuMmXCkdt1i/RRt0HG9rKUfbgmTkNXke6aS29Nd4tXfZw5R0GDTSYsyr6UEoh
KILTfKZWr11RYnNCQm7N4ZTHeC0X+ZgFnUdSyBP3lB/zgBXq7rvbrvtC8nNcZ4encj/kBRCsT5+F
AT8htxE8ZjfzijI4CRNy2wt5cGWYESIJHY5pU7nGTxWZ/cmXiuO8tOMDe/pNZMb8oyvA69VRiZ/x
HmEUiXy0WB3a4iCkl6+dtA/WWAuD1XqV+UZOfr1llUZ1cR2iL7SDceIhJBtHEC1tEAUAmp7o5p+m
LacrGWXZ0fGCaiT//xlpbY2McB9430BUAzW2x53w14ShZqsYgdmhLJA5IUmPvKz7s1s29JJTj5Qf
DMz11YaspGgsJmivbDxxBl4QQSvLIVdF6hD0AUTXMC54xpFRUpKh4wa78204APp2FITaZjGsOyxY
/JEkD9OTMJwK9JhTOFRrWcHyR7fsq+KxU8BHQVTDO5Qr5ES/vXsBLEifnNLM6VczYGBGyXn+8YLa
Ncc8dnBjM1u3TpVe3YDLVUg7kSDtJleVxC/W/jrevUhlpbOiTXTOb2HWG0WuP6O/PxII+hEetFRm
FFHI7y7JyGXZbWmEtTYJFX4qQqLewESYi9S0ufxBuulg+YLChzCgDK4WX5e+K0FjK333EUJ7Ba+I
pRv7vvyVO+2DKk8qa+lf3eTRz7GGEk5+OZiTDrOuS2lJGeyvSqkuuVUAqIG97nvLLz5uqX/FhugJ
w89gtjh5peEnk2WQxyVH4Xx1DZFMMIwMXxVrHxGqrfFCou3EVU/wdtYiF9AZyhtMi1gExp2aHRf6
CNXGEAdJtYCiDJX75vrjwQVmoffpLm2zPc6AjudCrODoUtzaE2v1l9UNQoQHMcU9Zj2gZgxuoMgg
76E+nXloH/2alkd3FsqQfUPzCtZls+zNmVaQ+anG66pbRjADaelTTscoYbEq3VFUSjYIUc9/Pjpd
vwxwYATAS8bb64NZu4FuIcF063kxiB1RCMXF6zQYIPro9pJszmFaqm0ZIu6WMN+DSe3XGAJ8K8pL
KJW5uTjjKb80h39jG2QQB8u6tW5vB8cSw/wTKTGTCCEMtITNQmtM+fN+M2w3O8JK0AWOjq5Nbfj8
a2Z0dKRds+WAZENzkkmXBLXEfceI93wyOB7cqnu1fzcQ2WpGFGE+V7A6K/wVLxQ5kbHg1xTipXL4
b83vwZwdIdM2xO2HSzRbQv6W5k6J77OoBbGyJ5ZIBQX4euZQ975IVqpQGkbpN/Nb8JdXMyM6M3qF
GNYgIE2guh5Ixto+E23pOa4j8+hqemQlE4pXwmnn3XZogZhTkgkgfj4K8wEvakIU5ovIXr4sTVi9
KGAXXlT221DmD9TX6FgkK+V5rvhv6OjNP+AyxPnqDNC6pIcHacUbJHoejngdHP+if3SaUMEt9epP
hREN22OjrOp3lR+n+DbGr5pffSy4vboy8esZvXmwGC3gnR60/nEdqwvKdJLz4scKu739PAJq/vXG
A8MMyXkhTqWDsUmUCgnhsUzgC6UjgZpDZ6XKK8NJ8T9KwszxJBq6QEwW6892T/R62Oqf6gD6sJVb
07FDYJDrGp/7Dht/pW281e+1mgqVwpM1jK4PfbQ3aWOMscX353fKpTlWNwAsFf+aWZa/4TlVwLdp
4cgfbJbNg/qfDhN5XD3nS5epc+tzBKzMYYpQn3/a0W3sZXP5CfnFJTv91yM1/eY2/vHzyExz9DY5
ns6jlCMoGB+koZsE1iwHsqPOGXJOQDkSdqS/zckW1VkIqhRS2zh6ZAeUJtCcyw63ccOrOf3US6d5
uksj8QhifGNi7deMNPAwsKelF3nOxYkTU057OzBlqbkl50IHfqFHdMPfckafP/CKxbKYNqGqLdiu
qD1XUT9Xqth0wLL1JNDPBgabI2plIcfhpZVVkn0xmnK55sNX27gLGMH69LQ/DwLuhfMPSnWdali8
BCe4UMZyUZBLGUqvmWOHRNkG/fgYfuPODkGMV1XMlQhHmxcNK9PyGQHoUcJkMTZjBN22Ha4CjATS
LJk0k+LG/anMk80PBCe53RgEndSZIh1ss7SaQlOB7JAHjFaYSncn5A1EPcyUz9PPVt92rqre8QTD
J8YvbA0KnrtcK3NHqefeZ8q1NMeK6shxLD1UIVFBG056a1dpOgFZXQgZFkIVAtZhgHw3j3gO8JpO
ykG3OJxsjYtQDS5G+Pdj4yYxUF0Hh+W0JqAP9DwMNlMfUG4Gheqm+s2+D8A07nZL6o+JMkgDXRTx
x85E3bUK5vtYoHhbfKU2ZOZ5PkLR8Qd6b+9GoncuL3YJ5vvSB+7iZBZprnoJMzWBekHkrFwRh8br
V/i9YZTnM1llsYiuMEgGHilPyS9ynKC0zRs+OT4I9JlKmBPs+2rm8JeHa/Jf+kh0MpA9kMOJJXHm
1FCAnIgwmET/7wJuhnqMGMJJ+4CO4MX8HPL+tdqHk+mt4oDt8uW3DCNPrgUpLq6GGznNnV8j8TN5
7KA16qf4xbYR+a8kP5Qx1eXP27T4IeVp04QH18rRmIj/Bqg49iOMy86OkbnuyLAwbtIZAYjB7yav
PNxNUhsvO3g711qc8GmNVuaUk8M98rZvk7DoG4FXFg1tih5Zxuavfpd53nQlVNBIJMBJszEGasZK
wxPp6oj/hfXZWaCOzZxPSmlnwOktG5GffUyJqXeWqub/0OavM9aCaX73pTQvduXO3KAey5toiY1E
DnhqftH256JUUPmzyvQGuXq+SS5AO3p/xc28vpK/K8+vM60cXoDMGeAqKlEsnxDW3jp9rYwHy5GT
2X2ES2GTsgS88WEDm0Ow56/cMXdIBh7wVvhe2n8WnDUdGW9W9cYbusJqo7rtLank2OIU5KNY8pER
xplTywe11O+GFwklLEh14lc4Yvhwn5ScVflBEqH2k+8MPEh+uowOtZ782+qh9H2UQdE9m7pZLLqS
2Pmctedn379c8N//L2/GD39OeaYG/rO/eRJy2R3uewZeGuFM3z0ZY6aoHmS3Rnvjtw1W1gCnxM/Q
ON0ZTvF1VEhU/klVSUn39yhSY6QWiUrCLjqdtUZ0+Qzq/vEl04tU8tg7rOEH1ZfUfqFxrLLIOmRY
ofbXP1iMcDwTyj8VChu3H/iIXhEGVPRMQcDCwchuDEcpHSYyCFaxgP/guC+JuXFb4qko011U4pDf
hbFpGcPprSXsRT0v7/pmeSpaOH3NCuoqx7GEvCsEWdEsBtCR+TdRUzo5DWAfMB5/f2O1Q6Dueq8k
RpQ2o34+euFigoAjoGVMKQtY7SOilN+eiPeXnlmIKZ/RSq3bx2ocz3bQxpmV8bNmlq75HKp2ZvT6
QpIBAA+QxarJxarPeIfxKycHuRaaaJ74tugoOEVqCIZzugBa5l3OHFbr40D2IasrsCP1EC/slET9
MycsnI2xh/wj+6aChSzIn9uht8uvMS8X76LRJrFGfWcjWGx+kcwh/ILpDDDUyvg8Z16BCaeG3a7r
Lqpt7hTzGrBgwP5zUI66AAvq6wYl2m8b2RA5n1pBxk9BaoyJv7CsYp862qa7yNmaC2JzXki+lPnk
OBoynL5HBaRYlZxr7xaBpothKx9eoHSalrv0mqmEq6uoqFz5s/0jIiNQXLEXMgRkleSbGcx36Xe8
krOPGLnNvS6A194Mx01Svu6Wfjebw4JtGv3LvqV9hKHUB73CppHPggPpeuq+Ak++TzIojZ6UMJXq
bP+uftl6+9wX0Ii8FlF8xrihYiVHAk7YtKPkmAWU6QUajgBiP2EpLQNXKJRmE1IdyUZ+j63ivD8t
Wz5VFGXm0TbQaMnLQtlLt/uxZEVx2spEFw15JwgFj3omYmFJl+Cfatl7+Z1HpdZkrfy3LIOy9dGH
YnCct/uWqvWeL7FAPALGu071wY1o04LuT443ySwwlxZIWWPnUfBQNl2NTqlxIkpOEUCY/9XEP9E4
zS8TGptDs0s/8gie6YZdCVqjaIID5WxH9nT11NouPBI9p2Ofhu4xKS5+nIpDnR3sm0aCMtM6DQ9T
LXkFEeItdXAdYtZ3eNrArRVGngLlsSC/TqX3MKSyMrqbmKUKtBXmralsfpiKE0UAu2XVRiuNUDRT
BCcTcSMe/A77Z5KMamjHYq/ZkIR8rx3yHI2O7eZjMwJN7bxi9PNHIcWS71wOKdF2oi32M5vSju4J
Eukb95r3gOlxTbL7EUEtpCeJQsC0Paw5FB5GlOpcft6vkwI9k59agEobHbBJ56YVukk0I8HGoz0f
CqStXTzyYHLIW2lysUx/Ql3TUkYkm3h0ydz0I51a+tVRZbK80fiOGJqIBo0YOAvIPj1yIaifb4ul
1493Vf86SeL4h2+ybyM1hrCYMGo/TNLarrv+U6QomxWV3azP/GozS4Is6KvmYO6l/Rs7J07KcRmL
3qA6AJbiMaLhmjgkc8u4gms8cTSEPOV0PJDnxqA6Y/v+1nNmu17gZi2NnjuUpnwBPLRKE0W0dYR3
P6+wR7Org7OsmSgZwAj+pf3xPQ3PR30B6QEljyJwa3klRkHHpuJy5m7EVTk+7oJWQllwb3QplvWt
PUcomRgrk1s/SENpysEsIL77iixVZo4Mudoh4QrJ7qZf4bCDpMhArHm7FyIIkRyoT7wgNhgUMi5d
e5MItzl4jhIwKZnM9G7XMbJw/LcGVP7adfq7txCru/j1zbd8la0YN0sLY24BtpXjgh4+EIDz18iF
v1EXp543WWLjDGBB7S6A4M5hoGR+hOUdoz9KimP4hobbxxHjqwjka0P6zkswVc6dNBAhFpBnPe8y
b+omYSjsoY6uPT2/9gXog/BB0/ux81rtCHNhz2qSzY46YtIWK2M/3SH+mRDuI/xrGrWBUrzbW+mX
RtVraOIqkMPXM9c2f9ZdvKkiP+kp6DIzOh9SV6XuPDD8TbZcGgxOhCoNGXKu74Yw+99zC7/YDY9d
RtEdrLbLpe93yzFDt7Ql+lq252BmPW+moXAUXj7/aU4r5AJd9gom6ZfvlsfmrZsWDtnLhdVTAPIC
IZGtWJ453fWmZNJ36/59WWGOcoJRtKYUwmwO9ZQy/jGWE5Ei3PxMLjd+82+nZB9oYp/I73YrVAXv
jZfQlKnmGJHvv4zWRxFM2B5rUgdJMFQ=
`protect end_protected
