`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13040)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9TaBM/i2ZgCPEH+TSdpehCfiyRo
8iKS9ghH4ejmyvQ0cS4siw9LjE8wW8PQ8NL1evZPv7m9zIUJ3PIOCa5oheS4QMo4ePr55Fyo5CEJ
PApvWmU+9E7t/s4OYsjhrJtcfhiPprrnSene56BJQIL7fWXqQEVoftAeFmo62sq7twNBb7RFIbAE
h9pZBid4hA8y8RJ9DQWKxoIAWLD5zyC44atCDjh3O9Z05HQA47OtW79l0KbjXUTF38g9pnKo/LJD
uYKHZsO2xWBtcgLAjnlNATNvgNNQbD4X2tiiAu737hxzIR+LOaTuQejZP40RAk46ZJ6mCDhSEfzh
T3EyL5IcG1OPpzcnJ75hILu8+MHkkghwOH+mCJxK4pHNBhCMOjq3OXJNh3o9q/m1hViMqwGkaiNa
t1x8gmCdbk6Vx2aaj4LMhKEMM1gdJpodfjgalHYZvFWYH8xZsViufWkZJ27BiyeqwCHOuGF2pU7l
+13NzbMu+az45WdnvF5DDTg7bRdeeeMB62la0oyhtlOPCVN0yIuQI/0/Oh7AvD5Twr3uYVeeopFR
JYo3vzCsxvNAqh94l2ymWQMWnUl8z4XvNyRuL+g3jnFIoeaFB5ygDunPIbTYD+Rd5sqSSU7y0K2D
uPrfdSGJCoEe4HySw0pKHfRaTXpIImzPHw3w4S65Ny1npq4pHveP/C5UfE1tC/hL/UtEEssTxbHO
Io2Hf4ceCEslwpUtJXJ4tAIfBNzajjX7vHwPZ2BMwPIllANw6LOiYKx5Ev/xZmK9D/xdcG08tIQo
ckf3LEBGOQZCpHni4uzMGY+ZF4LuIdJuBzDV+NqY00pXJ9+pFXKjfYC8p9Jnvme7Sft04Y8daQTV
q8nmiHj7q1j5chVTAVS66WKw0a691CKD7cIiuKx1p21t24nC7/doSU0+TWYsWPaXnF0RI4GlJ9d6
oO229cmF8bNhg9RhvRQxIlApslUHYiNtWPBBYQ4q7KitauLcRBfgdH0bQeL+arGwleuw2hvDOB+h
jgjY2cGBJWj9jFjsI0D8AEFh+uzf8w6zV+txHRijhuTQANAJACD/l8qCgDIOEn1AyudKcGB0Pbuo
P7IdJV3BL+K8i3C+Uditbgs75CxR0ulkAKSaJg7z3nhPvWC+MJn+3/I996kSVjYF2g7RWEVfBmtt
F01FnnsvFMiLU4gBvH1+vozqxGriUz7CaiK4s98r8jp+GXiJUEaMcXzmLur3fU0yLPYvpVZ/GPfn
9hFjoyR3w29RsPwVVwEtI6UIsdAjld3Exu1jyPd0YL2ii5zZsNnz1bmEMywUUL4TgUDp/mG49mGk
eRByMXH7/7NQr/hxCBCHfWHG5FAtaS7tjZjtzwB4S3RnifG/KqiOX8xp1IS6MlsqVgUzERTPd0Vm
JeNiNZ5dMnTUSxj/Df1L0m2lEM1jISt0f1X7t/fU3HzmqSXM4pk3rr0wNYEGx5W+/qpg+E3YpgiV
z/BPqnQGScNH9fVybB6oREl/zbiHt//MXDRUgGbkQg0RjqUiXwrdKeKLsLWdBlACPJ1ZeIXTkvKF
v4OZD/+N5zCobwmIHQKgM6FLtbFuvJJIxYY2MRvk+WE5yd0axiWBdhQ1XAjkGFAicxevGt8qyQGH
naaEnUlTLMtZfJ8xpDSVlCjJ5/gRbneFaOibVQuAoAXMfsBz1eWf7LYupd5vDa6OniJZSUQUIsA/
WMn19+scgcvzZJv7vO73MSY7rsE/6rSrugVVRg1XcSXi0C11kQI9yQYhJ97flr9s7bJA6hB2gabf
9RxywvBE+v4upm5uJ6GQgQBXsJ/G1Z8BakqdkzRJkn98oIXrLmXWGOLW5FsWQYt/yu86+/Vv27eR
5XAaLU5+zZljsxbpCh/dzMe9gqSyxRTeUz9fR9/3ARWHeNTirmgFsFE1nDlVp3Tx9tQ/O1Nt5mzk
qPT7ui7jsdGULcOV0l4uFPSt4yOTcbmJ8OJp4Tq8eL1Rsjv78ZIp/k/zIbH02w9IiwJxvSWRkEma
uSSFAzWGBIsxwhFQTv1WQGlsDKl1YX1sOjnwF1mZJ3IUg2tJTVR7aolIk6BYcYkxyGka+9b3txTq
sPck6royL+EhaUGkPe12hl3mF5jrYF7FGvmcD3hu8HE7CUNmDLYBFzoU53LmlC+O4y7kxsPphx13
J2T+GDWTh3aWQ7pA2IgNqpL47Xt9gw440OCtc5RHGGc6L/MxRprK3fRu4eI5yq12avhDsHAjjtsM
mPbXlN/sXYY02RRuFlIgArDXXqeNAgwzY94YfPZxq7cbIxIOhgPaC5pC+mMuKaV3mLRYCcqKZ6Qt
84g2/Ox7tWiuLN95isQXm6KByO8mL0TtbxTm/gfY9FZGwQKyneRKDK+5C6lOApZAcpyvIDWF20Ja
3EDMfMNx2MHlnsKtWIkD9OBZuGboGte78+RaQFrxnSE0zv3PT+ZNM1JzNNTAX0fIYvkbqyZH/hGC
QIOxd0/IXRUBaI5hFCCbQcTsud8eYolh9MiaglFP1AfhGs1tVIrQWL6EeMwbT3TULkEoAY0PLLL/
0T7S2IMHtu0+LCl0nwrEtTa5p2YDqxU4lfMmvQyz06hLexeqb769XEbD2R8TGlGfSdbtAapAWOZ3
1C/EIqBUeSTTHx9ewSdUC+YAqf1znK9S+XeOoOgyQWp5vIkjjndIWGDb7DYBjuKYkGvCgqHYYwXR
roqdQ1OWzzwkVPDjb13UAHjRqNI97emNzBAzvhjNzfYanV5H3lYlCI+xzOc2FgfZBrkqM9tyPWNl
Cbe+IaDGmKOdjHXceRGDJ/eB9zjLt38NDQ6RJnhvB9F7Gz/f/dlaIbqV9b8dzJARQ4ytVq1dr2gV
h0dYYuznPjIF+UuvV6RZuLysCbYRw2UvoteupLPfd0S7v8ShVUCVlTAOBZOnWd14pgtzSiZEr3gw
vb4ej2CEsF9IXvfXgthbdvAKrKA7JWLeVsNk2jjAv1J1VUfhdvzwDrzLI2YHwDudOZYR9qZqAtuJ
uXfj+MY3RIGhvch+eF/0CRpdNl2VlgcmEnECvZaiXzmSZ75Ktcg/vD2sgRzIY2BBbJlMMP0eDanE
26yvwwHKSINiRAYUXQnZ9boYMTP2loZAV4y9gLH/razgg49+NVzU+K769NTTHKmLkZvMl3709IIo
wLATJA9J/8Y65ikSmoI+AMEyUc6UZnB6OJD49UGEiOIthQyanYTGG/8Co/BaC78sI0jNOnve+jkg
nmyCFCcfNtAcfNVVmCsdApQdpsmK7mXw+60y+A4pfPloxvOPaBBIa4Q1ewJPgVg/2/RSY4/DxDmq
yeWWsp5ho0mtLbI8H2Put850y3aToTGpkhiWtjnZ5Elaqb4D2il8QOwWcVUaI63pLLSElEy4r4NE
ie6M/bmKzCjHyeXCX/Ws+ng7n8uTg+h4fKdPclmNpH4miBh/HI1dU9L8aH9CPmY9tzddrZhkY/4p
YE7llIB+PELINpE/Q75O/Zb2ZgMnln1Ii0r7SKzs9/R0wV913U4wl6r3O99tjO+w8cdz6CLyQmYk
8fI6NOgj6Divild9Tsn3WDanM+Hidtehv/YHL84HNYz/L3H2oRCfuC5/I3SdyphDgUiffwUA5liY
GeXYuuUGcMjsL8B9CqVcv19k2C6IDyGNSVjIrcEEID5bygidIaUGgyBTypLY/tlyVNU/lqmkw/5+
DdaSBGpIjmfo7e26FscwSDUXXod0RBWuN4ltYx4EsaSCv2n/t3dM4NvmXOGhb7BOTovBuRxyxRiQ
lpZGztnpp3zkDN5hBSgtdvIvyQDvcWI+stFjy3kVBzJElx/gwwfkgOLfAvy4mhDPTx0bFHJKCqd2
FVgKbdEwHx8xj5nWgex1W5zpaFBMgsg/ddfMHF81T4iyV0rr/qlOfrCFeRnZTbiyyvdSj63O5/35
l19a44KCH3KXltLR4uJfuZwV7u0lE3WKPAswHOCNKYVAdroSjU+OUdAMwRM1hV8IRmM0vm8UKLGS
AkDmz6AyMolEQfpuhCMHWbB2Eas2nBama1qQzNObKoozyjMGx3+EsgEWDgk+C5iA2CqVLmD+ijxG
125XAsYpcCn2TZFsiuP95giIlW51ssRruBz5oqislAAFnU1BAj+thr4Wi/V4T7akTqZqIiZex3lT
soR3ketSJKHfwh+T2qBitspRO2T9MDc3+0HbjEPNtQVTeqIqQlkt/PEbfemipWvqdgxelgMFKqfR
NrBMtxuENjn3O9sxX4KB3Dtnk/I0NYFTevWYd+QMZ+r0LAdhL476nW+p4AZQRHo8M/uuSooUFG+k
mQ8TSIg1ztkRiPyeFLqxFrFLqKxQWCl7Qk3Cam9pZSO/zklaX982og9eT/E3G2nzoVjJYEQglGgs
w9QuDsC+HcFIn5oXOilMmYow8QfL7UTN9WLqSznPmhatRPIr9xp8JECrRYBaGeLFPp2MWlJZVn/a
UyT3MkkZFVnTQCnkgOIp86RpXB9MjcS4Ov65ZEceolq+sao80h2+mwlWmdgbTE6kuDl8EerUCKWV
ssiZXDryacBmBOyT8cw86RQDOJ42FPB02v5uYvUOzNUHeTcTht7Senq7E/NzaGSNK+FiLabuHgIZ
84aiudGuMazSBx7eHfuOgL89vMV33Jm7pmizjT1GtTmA47Ahi0SvurUs/Bz1cbUFi+bSet1Mdi6R
qK0Dy86k+xU5HOEBwBZRKvmkDH++1x/9OsxH+ua13SLCrxULecDOknRi8xVBGDV6/SssNOSE0YoP
9nasac0N6NEXPTVrBTGorW/nkzroLb4FyrzdY9751QwGxhIBqE6KMpAiFQQRz+w5aj6o+h17sXJk
O5UWJepbOtBJTXaMjyrpFpx8UL8W2LbnCtg0NMnMQSLEu/a5pHRzgLq7s0KQkm/XnNXPcBfvMYnV
DIefI7advDafAh71hjQ0OlIDhHHUc23Y7WkAvqCubk6aCnLFZJNqfNk/3U2FV5auKpLMgiLdlAbo
/J4uloKATuv6oj5UFM0Lg4FNdCDv9rJbEf0FyDZqlx80ggqaRkgr6hAMQl9kqyRCOGu9kLeAHI44
WCRI4T6fRD0aKQ4Bf8H1HIfegMYw1GDbsRWVh8/SfOJ/UHtVGBYx3c7jvEtSPi+YU4G5qLP0Qe+b
okTvsrQcMnvlwmiaZEvlhEht5IAh8X4XguCvfZ1uw2E/+ZZDGpCWQDQujvcz+UiU6L2osBs8Cqi4
nM5wDRRV47ZF4HeBRsM6hsQkky+ROf4KizASkAuLeFxevDizgw2DvWMMShBwON/0GLwuDgllXyvW
45vD4IcKo36//8WfvbbZWWM8scw7X6oA7V6a4D5IjWJPrYi0WaCnuhzho8djvDXj92Q+S1q99Fi9
nEZpYlv6JDq7Reh/ChHNEZUPcn9SX5mmzunj2Mbf59SFM9UzexYYkxNX8sQIi6BOPM6AHU8lOZko
5hOOOUehnSyePAC0S/aS05NA+Inp4xs8JADBDTmP7tG/rYEMCu+AE7km+J9bofWOwxiqXVIoL8lq
mIkVzI8uTVfRi6OensUNh05L91g/DsxxMOXKMTsfDNCZT91u+cBJ/hLZ+2T3bKKEq+wn2nDPqlTt
H7iMCkWG1M3TYGZaUqXSOHJ9sp4sh4invPkxdYMAHmpBOASX4YCKypg8d975YMkBF7L6b3VIjTsb
bQb1uC3zyrAkt0OTyEvxlQFoCuH9lzq7o/9qdSJvgOzZJYixsEs/tehm6rnxHBAVqLEYFbVScDpu
J4didemMKN9ufhfbDM9mc/R+1fUWaRxdaP9b93Wt5Bp1tNYuEr14aB8BjYgEFDcgsof+hv3JkIFN
zDeU45m4v6w6n02fVc6EMuD6c58l2indi4+MLXPc1HfWtTIm+v9kpG1jnK8d3CnuNIAWcuUPuo9n
LoATlkb5PTnPgNe5qnE8QPDY4NNmCTdNtBbQQoftdii0wBgGmj18x9jbuRU/wf7y9KEsJkqt0XJ5
j+R5xUJ+lM8vP/lSqJHHfkaTO+E/5I9hnsu2EZggaIPRJ1jy2GaNqIThnYdwCmgt1WVvCL4UDisY
AQvFQuK4K1/xOd0PyUPr5FMkaa+aX9KAmaUPDbEP8MU1R8kfRmwnIbaIp85fS+Cf4oUe7LeWA9si
b3jXutg1mwgOWYJ6lG7tEZX9KX2T/CW/0hJTqHHk8Ot56sW9nxLQNLtetQX4SpaUlxxfGh7xj1wr
xMYAnicYe2mg1xG51Zmifn44OCjPrq5OCk/W84BROoOpBeQvTjK7V5z8cf05iJBXx6SCmC1zlaYP
U9OzA1l9UKa7SgTbzcOpvkW9SuGJWsXyZVdZDf8CrvWzxzvZzQ2SqQGEA86ycT7iaBE6x4AWZ5SK
H5FBm6JVtDxWV4z20cMcmOeadstXYy94z+q2rFgBzhLLh/q/t8MVgPpFoItZZR9UN86wN32sCbes
PIGFGZ4EGUrUWNjORtQaoy6Q/p9D7Gufe74QV874jnZAoXzZWgbvSokUsNCoZAKUChqnPW3x8RLJ
rpFqRdVGK/Ck56XCzgDAd2snJsigTkUq8SITH48ZP6/e98SJ/qPSLCDTStqW5yFYW89rFbc/RMVu
YVNg9MPOhwjaUI3g0GoOXvw6vHdO0B3MT4KWGJjbNYZpASNh3Fm+o+SyIqJeg5Oe8gQ0mjZxCBUB
ynvrMJa1CMNyi3asUVtMv6FzFixeZfI4hpnOeJ2y3eLNPxBt0KkQ+Z06lMf0xuxcMCmIXTgFD+Cs
MT21ZHiys+WCv7w/X4kypVckJTq1bM0LjUc/hybilI+XMHx9OxXomEIBEq2rpDmudIDFMNqwzcx4
1PL8r0cyBbq6711y0GJG9W7SytcucXY0c5sJV7bo0U9HSolsN5a1LKyYlaRyP1Av9bxNlyhITjNR
CWNBWTMqo2tetOK9tr5Fkle0NCTzX7hrta4EBy64/1SvxDl5ndeKgIbynRzPmXDTRBPrunq3LTE1
gon++w4LAFEBDLCe44dQvqZ0CfKdtdvBLu8/ZSC9mp3Pa3bpVyDnQ+VZJF8rr/R2WabXl4/dMHIr
B16zo+D3wxhq7SLr9mUDUB2tZsq2IZRyM21o6cwaOJUwAOAEz2uUtI7MmTohBksf/daUIyMm9qn8
6ItjKan5ynFFm5iqRjJJpujssGtSOwdd4eeEF2KpAFwwSVWZ1QGzunVhrhJR9v5EXmjUwUbQoxAc
MYGilop6PlZmUUFesDcJ5tnQlkihSMGA0PG+eNhzTM29tRFEAGpB53uNrpPqxCy0WAkIKX4LqUId
mw2J+p/+PRaoBUp7lRA1YQMg+kWSnrmaBFiS46kGEOd/z8lfQ8qaPj6sIwLEO6GCfuIfv4NSMBhC
HK+ISic7bHkgF7MyucHBhnAh4UVNtaMdmFmoMRHuXbY+z6R468FJfUQhl5AI3wvePwyNw5EPbF+0
SotCgBBM+ALPJ9MCgeWpGFfOqLoFSmgs6vN+7wO7k2u00661LofReXRzTc3nJzp7dcviaiVCVsme
P9NLq3Y0RqwMs+K8tHH46tFlkB20jx2AxGaZIrSRIhKns67FpwLlXPBldUHOZoK8ZU9mqbIhlRQd
ZXqo2VWIRDsUwbZ1xLN0Mq+8Qo6C6Q5bsLXnQTmiH29uabpQDyFS/LbszPg0BYqPGkADIba8yR54
FbLurMA/peZwWEEKWNIzY5q7WwgjyyDuPrSbfa98QS/tjGryQsb+wE35qFvrWqn//gEtfILOi9GU
8Fpj7bBgKlVPoLcVY5oZ48/Y56fqoMNI7x5xOP6qI5d57jVDwSj4x7ZnS5M7yuNJFilKqQvYFgQl
STrbA9wt1+Xv3zU04xOddJZTmVsdZ/Tk3TP+xtREB+kS0MAo52HJ3xMgEikyh1MLZjmpl8/zgKal
gLPUdu2E2DHQWRlDIwxu9uBPrWZAuEt5PLQHqQEBoCaPP1J91HUNKyd4uNjI1EbndihbexrCjXlS
KTJWxlJcOcqOLV5ebfcyjWNu4byyZuKAc+ezFw+Qobr0nuCxbF5HMG/s1KUqRc584uwWVQuwIcqr
nTxUOSZ/VvL5eaLO3/e2ZNyxXK8PqkaVsBCngG3AW+MUEGw8X4pUcCMdjND/HB2vyWlIe++JVI/2
LvQB7R8Jn12qfNz6GH9GqD0qd+Ruq1UFGMcGVweAhaUrmijrnvU2nkHcyKNy7ENXY1yEuGNa5QWF
oaFVFAPCuJP9iHewEleTKZK34ulv6V93C1rzeNZzmhcQRFAaLY+ilI6BZsM4eNOUI6Er32zSwzbh
kcTC8itLT50mJRsxTn3mESaHSixPZ2wVdoyc/N18PYGEE3RLhJiRbXVXh8qxwIaSY64HksI0XIZW
fnHA3JcIQC9paMrG77kfGz6nvwOm3G07yczr/3jBIx4ac/62oUqjdZNS/K/rxCpQbB0JrmJwsq6b
//xOaHHMmyvzmNoJE4BoRNYXY9uFTwNe/xBZMU2zJIl8gA9whNOe6L8gcoeuv0vStEYBHNv/d2sT
kcnF/7SXgSxZM09JCoXicrzIccqrtrlW3kYu8k0jduK+NO37fUp9db/df5ZoI5jjbQLDnHuCYIwI
Aak1BGchYqxnPokF1tr5qtMZSvz0vxp7QdQJFNoiK8xDYworKvE09uBs5/ZAAx1lVo5y92OUEpFR
9aTUyy7ruuAgu/4q5BUI9hUz8byBGzIrmn8vZzqkFt22U5lSz21W7XJKEHlttAsnAUsM9d2qISZa
Bs2Lr17k69wYmejPk/+MZGU4RNVriLDDtT0BPLKhNl2KVobNtYpxBhX8L93rAmzdOfZIr3MuMg9+
5UiYJxlaMF85gvsxRhcwG3YivVwmpACRf9mysYzW1i5MmuAIkOm1CLMdmSaVc6M+VqeMIi3p5W6N
OPscjiAVUNbmBT9R0K9vwPw8TMze2M5nRMi4s7QSwpzdrjs7cLe2/9ki5FrXx6YChaWq/rpibiAt
y+N6BicGaN3a5bdv8EtQ8+jj9ODj3wmOPSUEFXN/oKXcJvhHCNRHhigrsEkWSr/MSBwcv1lZe3dV
m34rNTq03JHV8R/+TbU3ru0DXW1FJIs4zdlFtd1zYDVf0GC8njNgKrOWek4obil+UV8vSM7D8ljr
MaMg3z9tDbDxMZMvydzGRpEr+Vsszy4nGiVBpBOJ417j7mhYUlFWI4Z6TKCw2Azz6PcZZyN8zyJe
NYebuQxArJkAQYFYnbzvPJepfe2rLhJeVn3LZdFOWdFo1l6Hcf5snRy3vjno7j/q0uX/k+V70j+v
UPI0t5vqKNi0lfVpRpi09pe5C9rBvef4c5Tbdtq0O8TpeklHdkd1JG8vEFx9ikB2NHwpQ9YIZOgh
X7qfFG0TMKuT1qkeg7wiMEPUtVDKm3TmX4+4+pvoM6Q8G/JuQyoqtbLAzg18UPSOaQWOV9svsaC3
rj5D1xR2hr1Fj9OALEny/tvllCQkollFrIgxPVRmV0AuYThWzolDnYbQ5P1y/1Otv2eDfFqhg9WX
5mq+TBKhFH5M7pMG/kB9gcLZ5M/Wix6MwoOUvPFpi7RSgsjwh1RGx2PcrUXfHSHAKSR/dtJ3vY2d
mIi6MUDAXVnDOEYsJHLzrH76DQkaWGDzXwp6m0ymCTkyNxIhCiah0Bs48gbdTxrlWCdXU1F7UTpg
7UCSREkDNblucysJjoEAvJI+HYJVNlwfyBJRFNIfIhi70h3/lskpYc6gzEOVm57z4U0tKPx9bGOQ
ivVDEx8Bq1pYabp9OZDXsTpVrz22wuFkhSRIK0xSmspDBOZTyb2b8TX8VFGCRxNU+d5EV3NB/35L
e2t5sLXyQQeJbBqTBOWi8BIu9Ai07EPFIyDKPyVKR4gNlRQmkGw7qW+HPMvK8R0DiKluyc7zNcW3
NWiPTXvGJ6dqk0Au+WZJBMmeRAEJIFdrP8Ut1zd54vQAS8irqQpQJ93d2T8rVYXkXIKZkAcCHySl
RRzLFfsGYp3Pc08+gf/qQSJ1DtcN99ssMsAuKsWzYhr6uaKyEuusiTIMsLtXdY8n0Jl0rYeEH7X2
5RSuXhlDkX+FBnt1UySQpQt9dCtAO5buLSKfBJ+D6pYOrCYksb+HLEBoBLm8smvHrOsJ6JQH/gDe
C8hVXqIVYMMIAUiMBgR0dbevqeL0Bpvf0IdY/lYQ5dp8qez9Op1n0/L3jaX7VUMqS8vuk+rYlb9/
Rs3VdlW8t41WmNzjOuMSOl+/np0wtBnh9Z6b3nSQs3eHSjPrLJdYaGGk2mQcGpzY5XHSI1w9tfH5
5meg2LOxPEdqPCDRnM6QDSLdIKRJYw+58mr3VFZbl9rX1xwv5Y8yz+HdFO/A0q8Y1Tzi1bTi50iZ
+atKaMF9n8L/n+irqGMmfSXD3NU9ruM5Xfu1m8jeU78YtPrxyZQjTUPQgiuboQIRokTO+OUD36H6
XRXUgpKokGts6xHX/LuEwzEFZM48uIFDb3K3WC5R/+Nd2AdGxqdnAyHJlMfMDXsBvUoAY4lM+Gxs
A5W+c9YqRbf/mQdsbJK/7ZxROw58pYTn7zsrNvl84wk30C2r5EwdyGcWaEWjuxV9ckn+RNKiha3w
mArxyF53Loydwdfr9CofdenvmtomCSQ6F6OoO2c7nmR7xR8/qIaVcX5nNvFP/vy+3z8xF5uGL6WO
lagC4dh4VAIvA0Ds+BwzxYwSr2AfYHMbnWYkz6mUIW6evqYkDZ6p6Cbh5JC/9cOBN0nrcnChdjMF
Zxtm/eCiNYMRFFctaS40W/UGVkgLuiHO5yk3YAOaenM3i3oea5nPr34eEMKZ8HVK3xIkyFf/+yML
92/Td4oNctc80aECyDe7lnq49K6wc5LOQU/On02mmmxqJOQE+pzJcGTwitAVRyjgQXB6YyWV/20c
I8oP/v3oZ/TxbGEOPquoPu5n68a1MDv+baiv/L1i8ER79tQAE8AzXU1xiaJ5nTOLlBIyXELff5Je
pZ9s5SpbzEuhyepqu2LYYKII4jvlXnhAa3ePmwOI/B+d82rl+vSVLdcp2bS0iR23hwhGS/OLhR5B
KJBSXWq5KWvr8yvLeT0KiFNfYG28oiSZqZZsUDizLagBZcHWhGqGjf/32b/1mAA0Xn/8ndJAYzSm
Z3FshxD20JonWtuLO9SB2itTkVUmZtDG5nLiQbbLDNUPbsHSXN9R2i3lF1CstL5M2sTHBz2MQExS
yzOm4fEor76ahAjJqjkMzFsfQmrJ8LePtChMMbz9nXvthIdl6ZI3avXeDRqdsJWY90tU18JtfVPG
YDWLpoyprOTDBfMP8OQA+4Bs6yk9wodfs7aKkH+bWE26If2L8E+dPeUNzbGJKfojy1ebArO1XmF8
TfG6lYlf5PTsert5dEhhax0Pp5cngzt7YVRDdDQQuWJG/QF5xSQJ+EHXRg4CDJ24P/FkT4jMowJY
h0N6BHeoQ8VHJmfX4pc32luYNPWIBURW09eHjn7djvSRIQ2xSl+2pWn9+RTH6qSJ4ymPPBm+tmHN
FCE8sS0KTQcmMXDp/HpP7J7l5kAXLLqPRPbWdBiJT9RvVVHrJ4/viCSDxI5sEQvOh3MVpVznT2k+
cxBUY9ivNu4BLje9Ej9dij9Do/2XZckXFKunJpzH0yw2UukQhjbHZGj+wAQDgIkmBIHcilXTXuZc
SPM80MPtdYM+4XJ7sZi03rVHVQ/9uWrWFr3bQ0E/FzSK/a9Xrt1zisW67OrpQaewdIMXRWzzgyW4
FxGtwTWGpiDrGbQJTquRUMwmQdtyAkixyt/kT4pcpSgaIiHf0xgKjrmtzcqNEgswecMa+itRagkz
iFzf5ottHzTzKsB4F0x+T4c8cX3EL9mIaHdavhuxuOgUoLBduBMSiubqxjpwVfS2SU353WDo9hQS
L55B1qa9Es6BAw/mjUHWnsI9k2T2Se78FORnY17AfW/d6TMs0TYKtGC5ieHQQzBCtKsssovUOSnC
KB1P7VGudofOvrJUn6rm/OtDRHf/0y7WU/T17BJvTGJ8RXYOOogtfdiFUhel0cJflwuRuTyE+pml
XGgkcrbd85jEUOycPqNKTCg6+xBCghfxc7UR4BAD7BFeBSWvSjFFaw5heCdtRTCq8E3xioBTd/xF
6qtAwtKaAipUH+OqtH/1TiGhpLL77tPhU+ZLKcrLavR5gt/ldmDh6xMwsQ2J6v+SmlgmXjjM5oRM
knOI6FG1Pbu6/imGguzi1JcNsuKqzIkHz0jwa9XgkNISD8TWHy09zi67jEN4sNSEd2S5JCf5+68Y
Aa6+1aom6R3xz7Vr5O0aJ99lssy7+EsTTeqaILazdJGFsjuRgN6Fk66jB8FIacCJRNdDmiA74p4Y
E8oRQOzQlt31oeMrtOmTUoYmdw2bmc/Ql6Kwn4Xv9GsmZa+L55By/Ug0WbEKZhhMhxRnUNlKKQnD
j17KRKKzQKyo2cBXqZGoftcnRt/zMHsVjXjFeWzBtQbdBgbrbGrd7x0Xs5QzzHMZ6K84SnP/lfDB
xtBGzHACtB1etGQljQF5RI/DXyisX9jaFp6wYrriqaAoOeJYreCTDaaqKhxRK2JlYFPhlNPFVc4I
jdz6ZpMo/j1tzeS7qZdCxCItt4lkt5UhvYb955epjzN5uXC7qjYueYz4JMq+QQ5VcmN2GhnVFxBY
0BnhyDCXmcoxR8U8xe3Zq2QcgzGBWFDHvNHzaI+SWiJpd+VW8V8xLKYlvb4UA+9/nPq7ImUqnhVd
nByhVYQH9QS9e/IGjykZR+fFwsxLSnyNFct1RPf1eNXi5WyavnRabDrJAL/6jLCAT65eR66tUUEU
/D1Gp8lWvpeArZI1GrrbQwlDfoviHICtCZJMF/NyBhRfq9e5aC2nLSeTLZAg350tyyro+aFz7VkS
VHY/WU/KuSEk/qBpRa7IZ6wC+vHqKQxUpyT70O8uFH9xNQN+gBGiSNv5kML7DEejiKBK/ruqpA7T
1rA/kZ3UU3OMtV0JdVTZDXbVFSD6jO7JKPMqJSji91wfKB0bKUfawSawfgxSzfBnfQ4Wz2y0sx3r
9kSxjzjTLGHH26h34Tx/ysNaIyTovp4HyaK/4QTK5oG2Awk3eAp50tFWwrJ0uOiQAuJ8P/rwxOYS
4niUSI072aonNZIJ4jDTaKfsU0waRd75T13uqI3IH2hyL3/DbXhJsF8nDad2rAprDbnYMyQKGeml
ZXWUIrhaTLpT45YfNJvJ/yOVOJxL3W/QDDnHt4h8AyNd80EnPQJy9l4ZObw7vXNk9K1Ce6KIVCHo
8zB3VZzI7vcPNj400pBXLbeIhuWQpzBfk+TizqFaukjS/s/Ul4DKgA4Fm3V1u4qkEP/YPrLGOa4x
Py8XSw3vIhwY5JXCwmh22XDco0NV1pNnpfqXq26U4RZuAMOf1elv1hApEPQyCEqmcUXEviedPYdF
mB/2uS1XhTaMn9wPdkXmicVHM7Ke/jukMTzbUCONUAYr7T7Oyg8ylLTCYj5OVdTGyhB8aVVD+kzl
PyHZmeo29PognHjgjIQWHNkCDhKMAMcbbSwYGoaLVRDr+kNWVdiNGIt1Vls5qP1voxuMYheuO8MX
X4At7MQqkZs3ctpNNTp5LTUwWIkY9z4wJ+w4WFKyrlkKe7OEzmWk9p9S2qhIps+HwuHIPdghXchy
C2fu2/XSFVyX/sL0KEXa/SXvZD2OJX6QxrlAa/xKmAxmzwBzgqSKMHXOr7uSPT8fUtiHmu0jJeGO
6Cqr8UMhK439VH5qKqUUDAcMK9xPJVvdkLKbvb9DSW1Z3CMZjMZMnFCKKU8yJ4BfXyaH+H2IFWA+
NrpO3xVVCsQUkFQ/fJtdH6vr+2lzFTurjKODorLAZBybfONOfehA4AHLm5YIycImPGsCUGR1Hdua
5Qpqi8qpmFwJ+qA5tk4Hzco8Xggt71EgMctVikhTY91JQLdOxBfrt9Fa6ygsdy9zaE7BJJJ/jHth
wb+RYBoN2/bjh4Lf2ddnvNzgsjhRIz764HQ+muVBQBKpFOmapGa5ZBHsTYPZ6aV5eY+KTN56HmXu
J14knnWFIqvG+3EvcQ/CEaHE8k4KypCr1GHKmr23XKPSRGMO7/IhcAf7tb035ZiZIsWgspgBLsvU
2FnqRayWFTeYGwStT68cKUYL7e6tlXVf4wBA1doL5TIIb85JtJB5kB9yl8RCDpsn+oZb6QNPUPsJ
Ej08iMCgVOZu0tIaFpHyHV3netEpywhjHJytXq2kKVav2GNgpoIjrSY1yE4=
`protect end_protected
