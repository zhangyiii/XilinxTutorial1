`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
d5VJXu82JfSwswDjhvbEU9He9tQ5/1Rw+4/2nB84LUuT0wfekcnbAADJNd0/JtXdeaCUlOw7Zwks
Bp1VvQeB3w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T1a12gH9+o/WCd/uq6lAozrIbwFwnflilDyEA/rZKRAxvRmKOSqBXtjVpxVSoEgX9El2BLPK+36k
Vd8y/iFx5HcwlteYeuYuGTvgQerRA9ycH4Qwt9s5DC83MaSGod9ecMMI8PPrmdJ+hCOX8sXwEsN9
IHAKBa7h08XDRsgW0os=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZE3CBd8eugZohbo93EvXvQkUxCnosHfYT2eG0uuvFgW4E1aUdxFin2hcHpeAodvxBTyPhYz4Lsqw
3nsUxnz9hTb8Lhj5XnlqKx2mVFP8Z35n8lJk21C09QHBGoSukklDPI8dbQUv/KxN+k1qsLBHfCBA
FWz2UAwKlgCaoOPe87s5MUwwDM1/P/D4+XgEQCRDz/7JDN7p8ZFVtltMEx51xjJOCvfGoEeTzG2k
908lkYgt+B4pvwsuFOHwC28xicC9lqwuIR+OiqTI+hvqIl3tijnK9dhEHXmlIo9PqdVp3p9K5niF
C0wKwI1gK4zk+Z+Qv31AV2g5KDXjXxSpUgHlpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1K/c2Exmx3hO4tktdfNX/hsUCqBDw6bH/vDRPja11f/SX2mhefMgy+yYp/XXIVeJlyTPI7AwLQ+m
jPsm9qUsxInkPzY00BDkxz+XjPmDvPZhWK1LaTfp3S2KuDInJ2AYP1AwgClVQtpRFpipBFYqQeNS
QrfV5V8iPYsCh6rtCZ0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z2R2Fz5uoP9gCKKJ4H8ByaZdL0II83JUVbmmEiqboGhJOssYqqghHZS4Xla1DO6PE/W7lUbFZBMN
taobe7WZ5vLL3z9KT5znQ5u/8vqZfQZBnNTCM9ij+NRl3PRmkUPrtcd6xURukGspBspXFvJDNTq6
HoC8rJF2dAK3E2hXtQ2qzFXYx2JspRBZw2ARE4ENjzYZSYK5AhF3nV89pEvyjDlChnkSNr7Ec2sz
zSK49rQXLtbokqxvvzCHRCEs+NoMqKlklN93OyjJFAIzYffS6GiGtNeycU755Cv+/fAQynybNWn5
4vdHnb+JcudvHzAJFK7/azTzKOJrOSm9uJYTZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5856)
`protect data_block
mvi3i3MBI7n8zvuunOT1BP00WZoIE32W1Yzbr3iOt/IzCp28BQXhRhb8VtZsZ2AzQjjhh4sOcRfV
iMWxiTyk5ZyZOY9vU5roLZT5k9siOZ3YHrZG6ir0s1EWzQ5xGohEA9TtBTCGOmxMLhR69KWv7W/3
S9rwQinTKP4JWaGJumzJ3o72C//EKUWRZgS7+t5YP/Ic5oe1f6GfaE7GJr+y+Rlg5JduSPEpENi/
0hlBMEWjqnlSm2er9hZ6G61OszyxZ25rtjYj/aeGGUrhu1MYzgjOruRRzgsCFLq0OTSqvne3XxkE
SN4LoA2V79p4KQJJxJ3An3a7G0F6zC0iErIOg9fYSSydgvFrKhEoVxxf/4CAlo3dp+RBRGcUxRt7
Slk2tHuBfrgmBp7ToMpH/TpxHfWUAB0ZW+5tDc94zSm1Sa1TGYOC5/aEPLpKSjLW29agqTNTn1Xv
fD6kP/HD6D01DUt5ErMAqsEAGbBVFywom30MKlzWVlUzDHivqEGGalpezfau04YGlf8s5bBFgwSk
APruVUti3qV1eH1YX0OspCt4taPYGqtwN+fWpUgrpHiqumaJRhxH6dSBbtXY/Exk3lNUTdNMoMz/
47tEQnH5ZNzO3wdLCxHpx69EYTfFMKmNBP5+QleT2zRK2ivcH8wd99qhHGCjI8dMI7rLu2BIgW7K
0cvtPml1p3fEj1Z6GANmqrjekuUQEJafUr4IhJm4ZY81ek2VuEja5PqV5JrxRzuDJ1TRuYyZlqDO
gAs6bJmNOjroELD+0CwiT4Dn9bwFKccvTHN8UxMRciozVPo90fRxVZTILmLvZJEjjkDPv27wvqmY
9Jb22KuNJcZtUSETAwKSTqVgHH3s1aeRpgxk7wgRpNlsz5fRhkBx3nXTxChW5z6XqjvsgBsa/T8+
gzXpD1jco9R1006/BNwWX8ryzWYWeLj9JFqSmPVdCvaNwKlOmeA7VWk5NxRnFs62weRcEmNUy964
kwtgdwW9Sjm/3nat/coy8d89f8MGz54m+2O6SdNHGonDGBgGolvY0DEy8HLwcVyIzcLyTmV/ezRR
SZNQgZGuxCISeXmroLEUeh4tvUj571iQbUkbNSJQD44QtTaXkw0ObhG5UQN9dGoRgEoBVoviY83W
HhawcrzkFIxQMDlU/Zy9fgsgJCwHSLy7s5dHo67keIpHZK25tZQOUGnh0r+L+j7PxyKtvRJ1b+wF
T0KhiErKNwGoZ2Nad3IF3enBM2UmwxPllDST10z7I2r2hPIBpdNMJKN5Z5jr1kbdpsr0KFoC4ubj
Grae0FBONNoLifK1m0C0QSc3rWOY6hbY9E3D11GsCWY6Th2FRKUuWOa35sQH6VGRVS5y22s32e9h
JRglPcTlWjNk2/LXeq0w3UZ/ddQWt37RR1r3wt7XDGMSTsf1N8c+U9RQGsm2gEgaoJz1zFWyA6a9
Vrshswu3rGQKj8lGsrezXB7Mcc2rKmuBrQOgoER5yZ3OvdUoRQWt09EA5Hnrvp8JHnaWQtiw4IE+
HW7K7YuAQ5MvhmBwMVqiCJGkcxRvXVupPRNgsrBGoSbez1D0o7+ovvYz7jQRbR+rwXY/OKQSPbcr
9VKsBWfAbYmjH1SVMU5JEBDpzfuYCLtdVLbdTpTyCsjVgWlfGix71FfQYacu6tyOMNaN7jntiiOw
81B0vWN+ClWTJ/mMyGg+RZTGlxW+/f+hNDuQyuppVL9MsOGkH++WHq4/rGIl0yTM8vmkfXtRoxxH
0Wn2usYGlBKXwifAamUrHSHC78zMBQN2ejZJmJfT5QOS3uz0T/qzaL0JaZgsUsEfIDWsizznT7fa
8hfbfpeFdUh9M07AbTcpPH2BSVbTMDgqbY+Dd4d6OgRo3T4FYDusA7mhEF0M6TxiewJ6Y6Hvbay7
2pM4JeeeaSN9JQkSXjUhYmV+oUN2rz7am62FA0PmdiR59N5h3MXlAgAN+ZQCBDRd0A0AbU0nbMwQ
f8WWa9KUOBPf1zwwCbsYDU7Kutz0c+aCbdi3Tx2yVYUIP0IVsaRg48Wj+H/HfbOGCggRgfDHUWH3
NdZ2mssbn9hRjX+dWbx4fkIBmrASOrWhBZ9ntY9Ymbra/zjh8B9Y+oCDhKVSma2WMsSpfpC5zo7m
5W7bny4StLQE58izMuFGCIDyCHy7M3HW/mQ3jlcbG3YNKQJGc1GDCEpD+hxEKAhPrL/sRHj/cEpo
P1oh3oPWlGq1iVKpA8YelMDNTtgn3B4DdYMIajGi7/Mv/eVkJA1W+39MgUtmARfrzqHync436/iH
Z+Qy7CyX/vBQOCjh8ITpXMLdg4S2pzroU7vzQCvcdtl10CnIaSWSMeyUT0qnD18LA7/efXMOCY/S
qx0I2qGxTf4E0/7sTJ9ZBqyFEB7muEnZeN1kNe1Kkc+Ax8i1wwhuqQYIeanFuXBF6NmQs+5tRCQR
2HsKfr+3MM1NVownFsluLSVgklxytz0aniMsjnpK4EZDn3dK/xzC+qBXToVHdnR/PC/u34uexsxC
1tJHqWbONo6YK3GKdyg2jGX8i6TFKq3hd52NikMUG2W2tjn5wmIyv1rz3F9olS16zH2ITkIOAGha
rJMFRWICaRM7YiTRjXVfXx75YJAtC9WoX/X6CXe6Nu59adC0rbvEAhRH1+5JUQ4TK5mMdyyfd5mN
UXeKpEoV517UzZO8hA9vXeRYcOi5aUA/GCDICmEZjZhPmFAkkeiD2N+bl3YLnME7j8opwas+sQ7h
cEMu8JtzWb5Z+cHTfPYs8xN9zKmezATNpgN2sTegXzIwlAJdy2iFz4jYADBnAD4wmD3WUiSTbhWj
iEWzkHl3flxNer9lb8qae2RAwOvVQo+b2tob00Y7FIZHt7WnUM8tcQ2zrwUy4wge5kNXY/uGaegs
dSUdRdyQ5XfKhXM6t9IPudr1OmP7FXmd+NJbukUptpCf8Pe2jXY6wkJOdyVikTRmHog3h6dR9VGD
u0eNJigHGYNWRgtsgHwVuw6O/GvT3lel7BTUAtEulVDtQwlzSa1qQl5ItkjLoIHOm9HiKptwry4E
BnBqwoYn+Es0OFRZrV5MMV5iJ+InpatUEjtfO+glYfCI2D2ji6qirrhDJbE91jFV4qlC+lJXsXMw
llqsQqUuITvydpEzBigC6Miqlo4droZ+rU93xnpkoQ2FNbyv6dPhGbz2DM60hJ/hjbOn5MFEGQfC
ahK8bW3dznl9I3d20xudPG6RgjGscOfL2goaWpesZen/kY6H6mxXtm357Q2//i2plUt+o5tUhlci
T8plqxPAGCV+0OIviF2ztKLe58Lt+4QP/wfCwvXMcgXza3EPDTJQ498+KSe89vfO5bL9gyURBmrI
AB8g4Ogmmtw+ymkh17nRWjNQjNqqLwYWZm3qHHuhbQ3B7L2bNsZ1CtLg1to8MrbRTp7ISim7GBPf
sQ9XFuzJW9qYEhyeDwicIpV7Rg/NTO4X2kYz5N8OTQu96SNMQYVG996bFiB8RHR+FhS51AjLHXgw
26E7wvqVthMqmRuYJjnEWse3zzBft+xdZs+LExzhHhGAOpgq7Hk/vCBRej2UlUwmEBSMYue0i79N
CRWfU/hGecEQ7Im6e468Yc5ce67mQb8ONddKX15aoJiQdqqi2LFDIi3JMLIu7OaAdPNeNum2HZMg
0N3+J30o4aMdQaJplhU59d28Aj7K9r5+Ov02RFtTTTx64Zxk5pxaGk2r/9+WY5izmjHwAGIlMZBM
RfjQrsDCdASrNGqvJmptBeqWlpaMeCPso9jwE2ZFX4XaMmS0S5FdxLqgRezeHS7B6ay7rVzIKm2a
dc8Dw494FZgVyHmdwrG+mDRg83gXCZELIfu20pHp6zjmlLrPO1nL9DjNwapyc5gqj1GulcU/UoNl
OrIJuZjaCX65nUJV1r4BSLI74LNmkxJ5s9QvkDewQ8xlAtTn40lXqThV7U5sM0Qu8pC8rWl3yThi
a5Wg+k+YbkeOW9zJSau1OeWIzc0fANOGC+g9TTz0yolMqDQZBzAyHpt6xV79cVvaHLGfMi1nLC4Z
ExZkqoccV3S3XniyF2R0VVuyNl1XKgjpnnDlndk5EN8CxZXIxJ/eK5202goE8FfBYiXjh+ZkxmuZ
3gQDW4rln4UUL7iwjPy7cyjb1wbDH2Kk3jFtRdJngtJzkplYhGLaC9pl9K8P/LQ5oF5D4GUUI5/L
w2FEktDHI4FOiaBDAO8j+473dX18zYn2y8pOkJ4xPSZ+fn4hcC9NqEg9A1hKOh867woNcZHnXbrR
C/B5AucKPzl2YI2LxUx5/I6jl3QqZGFNe/BSpOtv98VhN7KaZayWb9uu91V2+16N3xRWij6atUPK
Vcuhx+Jn1y+ZPmg2+oSlgWL31vYEP99K4p75dsIy0P7HhobYbSwTDOyzw6FOSkkdz3qb/G6hm12X
27sPzODJShn2+6C6vKUIHYrgzNH6Pvjzh9aG23Zxx+KfQ48gsn2AxFTgoG4N01r28EOcTzWsG58K
rSJxoaDcHJ6sdEOKEdh/MnrG8uRYOTysLlZ/oU4vqtyIyDy8uTgggqzdxxGwaCYRJ9z8HedMsbcq
UlwKiVicaeBP4Cgy0bUjeNmJSE56ywrtmcrWC4x3joCZFupdV7cfqU0+7xMz3hrBePHUf/48sJxh
Z3aJzYfHGPMpc+dt9jTBdRfSZoydYw0pgvLEzY6NIQmHtlI2i3pGmxSeaTiaoQNlVh69KclnRLCL
VAJrnJwn2F27M5E01huPWTxHkSzIoGMBcfvKIJ+VipuQRPrYyJSlvKUlbPB27zUtHajazMPWOe0J
QSyetIMcIvWp/oWDbQ8R7EHvVOVdeiP/cAWvvWX0Vg8BU91ywqfotPLz5Wv1AWIES6FU0TY876BL
M6z+wlvmaZ8KpY8hgQkh/HcuOp/tk6ab1r/6xWMPDFrnw9L5GgeJ3ofUxo92UgbLwO0OoUSgk1PN
9boebtQTyR25foBfqcKQz1r2m/Zlmxug5zvK+iOF33isIfzEO9PBX8Q9YEPc4pjv9zmLcnYRpNSn
8Xd9sxvRgK2LGcw0Jx+j1PWfo98sWwqpxnfJgfRLsoNM9301GTK7ESaKIb4YkPlnsDlA9KGfx0KG
nLD/fmjWyB37l4GzRNV1NWIFsvhgMI/7uA3Rb8NfyhYUWrEZVZXULptjhQslAMZHrpb2JeEmEBsd
EOptXcZOAfa2YOx4BY6/+re8VK0u7MDQWJpfFRwzFKMMFLL582cGtsziUAFDrK06vmf/C6bsEQcq
Hgv03Dgs9hVN/sg72DLon2kXhJxtMUC3+siXHG5xAaCLIzn6p4zojD7Naq/059JJ83+BPd7QUDVl
E9Oxxyc93Iygxo/Kjk8KMz3ZlAkbNowX3RP7QZkt1lkV3oTdz/vzx5w8mEEDFclKEroZAaJujYUx
LEH5IkdzD4YgpSstCCFNc0C2YngNHZWreXU0Lh9vhgnG+qRneP22rmJRGBrIjIHGWdCIWM+eJR7C
zQx2MiA9wAKKGAOuME8awmGhJ8dlY7M3cSiPrL4MBL3HN36cNw5Qq+c6CsdLdvYfCybU250w7Jfp
pNGfNeFno1AXhFY4Sh3huotWeyV9pz+exG1FUBuWC4MbbfPhZQ/9/sisKvmGopFsYnxu8b2d6Led
L8ds8qFGk+Ru2BPElaJX4x6ab3nOs4QqnDjzHTThqVKlYfiHSaungQXOIlGLWGLfpVNPrG/mZlxz
zoD8KBMVhlnFulAcWunlde1EvppK9tD5bsUtDLvcbO+m3TU+G2GGrr+QGN4R9wxIzTYsfD5FElsN
mTBIb9c+i/agnWogeWf44XGKZG7+1FFV5ApEEQyl8wF5yt/0ktyZEpvJA/PLSDlNjLqh0GpdzX9R
c+xisUiriK5gPs+wRHBp5Omnkv0LKWKYBjAElK7WJ7vfS2zL7HryLS8ExKpGrKHTnAVJjK01ob9K
yIfDQr+tXsb/fGeMK0BNqv4Atk/1l0cPCCxdGc5dyjOYsWwPbM2WjcrLIr2LE/egKvNtTBZg/1rX
8kU9IKORnhhHhVp3ZUXxIjzM3m1ZE4hGGBiATzsfEX7apcaxJP4/kWYKj78ymrDYULo7Fo6Q2Wu8
tzDFwl8OfKwF6SwNets2tZfe+qbfx+lf3RELmIVKyrw/XkGZ9E3IUdCagBNqgwzCnQgxQqJBY/Pg
9LHxqqJuL52/+9IyGflkLANkWCk51heRShu9ZdG/myh/vlfNqC7WETDgM2lCjTo3ttTtChY8SKgk
z/SiQ6KW0t/4mg6b6R2Sqn3rBRnsPqPt43pgRa4+lilVP6b5AIVM7YHU31YUk2FKr7gcyGIOzpG9
LP27JDRt23OMBgpt3MozIwF3xCQeOMTous0TPLA9yjl1wESsQNFG5jlKVzI0HKBHAjloDkJ1pbUd
nJn48dfnv6egFADmoT1RxJQrQ4ZK0epFSk5Vye2A7+ZnnafAX2dRe2u32nmwIATI27xUBtpDhxke
o3hFoz24ziIm1S/tFTbG/Y6M9ATb2uPYS5mr0S2j7/VD2wSibTZmWOax1O59utd7g1MsVRJUmcdK
db2hmBOog7LlnDWTVompsdYsjcA0gqu3Di5QRXbK0RUT7JfvVxuZQ1eK8syYdmkr+If+QGes6WRs
nuncSyqZjSCfylSsLXsYo4Dh1D55IssoCeiyC79NDp/sCUS/owU0U2TGIU/3r8c1pksqbz6l9fGe
vswdTZaDKEh1Py/uh3NHp0Ol9WKD5OPTrdbVMRnUrbhh7aJFfpsEw898vRcaHCvu0UBbQyjvMD3p
jtM24NlZTXtl4tzhL/K1d4WP2DWl1IRiEteBRhzp92iDq5355SRGtZ2CD9g2/y9WwpLSJW6GzYPl
yMbqW2r1H3WD3DXcG+UHqfmYWG/hzX/BnhHMjDh8B3rPrAXs4JpMJ175Rc3TX7SqZFHtpKRMP2Cd
0Yd4YfHzqunqh3OCfND652fNzqGu07EBNxpeQqGRz2yvjEff/YJSMvHVAkwLmU5BFTGlF+FSNmXf
zgPJeYUnkTB5lE4LqTvWHmoww6wMIUEoJvTFxZI7DUcLwClrnyVgQBXHbM2v1GQHY/LOPAw/VhvE
Ulf1x5UgJGYdxW8fdbAHciidlc8jaP9n4gAsYf4adaOtKB70zA/rDCCn2g4b5dg9561z2V+ztllO
o3hzqFnw/sKgfI92O7wZ6Rmq+ObtBH7wwN0xTSuPVSRqj7ian2S79A/4xprHEdrXRRMoQFeAvMXW
0ct3+m0DN+DnxjapswbjDnAHF2/kUukZax9KGEUclJDXyys/MST7icHUC64Ir5Lxvraim4V2d+4U
kuzitWDMiAXOCWmHQUsXQuwGTX4S1MnN3jzqJGMcQVKw4Yg6naJHa4jF4vvQp5ZyonJ6l1a+upfF
+P2Mc7w3e6DA2dupzUui81Dx+IQAHt40gUDInLGz2J1/EnVSDcktAYot70lAh2um/U6yhFaQCHIV
J9zMBWAs0Z06LcnLbG1yQ+1rgh2l7xybfkP8+mEbKvsREz6mvGhPq/aE9iTq2RGDDIYRpNnGJbzu
/VSlYfUhtueS690a0iC9JjCY0Eh/LSmLIrl8pVUSFRsNmXb3tgOBVofP48qsNbHAtmXxEZJ8DTkl
aGbJzgVeWQcFko33tgumffSyuRKBqT2rOSlPrwyrsCS50pkOyOUKQiB5LHR+zyDdRag/T6Flpnp6
eDlLkUifczOCRaD+EELiNnrd+y/kUr7HEeuFKSJZDdTmtx+lBCtGkA4Wd2eB7J7dlgKxY8Or3ssT
bik78x4IITprVx8JUkLmlWUaP42AVH6A+ubFPoE8ZsQD8uOiVuy3wYKf
`protect end_protected
