`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAJ2EREsR8/Dl3O0QnuXBDFaBCGVoF1rO0mFb6QDvILV17bNEoQpuATHk
MmorMp7ZyQ8JplfedtxcjTbvtvgSDTjOlfuqjCiW4+9WQalTZMXHrtq5Cwu+SjZKn/eFOE9IgvIY
KtdcRGr9csmIEauugaGrL7Rr4gx4YCX/iltG+2SGIJfixiy/CUcv0xuPnfhOS0WxkRw9tzX6BDFr
dctssfH2ukspaO7IQ/pdUFOUs0HEhMDAiPDZnY15r9MEUV74opq0gVU5cQc/kXIRTMzxIIxoUL3h
NJxhlJC21ShQZ+YZVMHbtVgx4CmD6E+fmS8TobhkK0ytdHYw24rRkWUi7ChFrJpfw9YCJie8+7+P
VciRtZWKqwP9cFNUh2PK64oqQIgSWCiHjYYok5kVCgywtfrJR8CTeMq2L8H9iPW99VW8Se8CmQ8D
9ESgna8szdPVMztbo44w6/koTVLkiq/2Jk1dfrq7Rs3AZhP2mec7HZzQ2BKBYXZDJOTEz6Vw43Xi
9owpZtDXsFxXGe8JiM3/K9TpEvrPuWtPtPVxUM1WCYHMlfY3ZmSbkfwDhmdE3Spl/uEi+Pvdw8vE
mhQqyVcUr88A2CK12lNH6al03O8xv/Lcya3PSdqRy11N+L3uOSh2Vik6j9JK81QoETdGPkbLqWnz
TXdvJytb3H37cYtNYfwcvZZK7JrCiQDbh+dwpW6VKnzyIetvZypkPt2ghp1vAXLPB1P5rl+SEjwW
cMWQBIpLNAfYjmlJ4Sr2qyJpaISrHOufRuuJPtf24e0abOCgB+fa7XZlGWl1aMyd6N3jJiUzpWls
ySgZPXQiB04poQO3/w9jCNw3Nvx5HnHh1TlaFB3nKIOdYFb0FOS00QwYs1dfyJpnBSDajT1NS6hR
LqJfKXA3oarsCpOV6kI8znsxQZRLMxyJKtkNdmw4vSWbCBwHhza+rsO92mCM0MXfAolP4LlOEd9O
Xk8FXJizqDYoerEyM+kZwFWilpEYz28hW4VbUyrIS+cy5z8cuL+CvzlaiWdcrEIVu65vWy+eLH1Z
QDZQsjgDL/PNAnlemFEuFNpIgRdikZ6YR2lJZ+E9qZ3t00z+ji/tKj1sY8VIw7CHVVzRFK28xrr/
zmxIQCSQ7WqZMmi1lmiPsEkGTjK2cXSl4TnCvOaclXshAwxYKKX4VQy14is4LVGws37i3yLlhgdE
oC/ASkWggJNUxffVbgvuozCDv1TJidUaCiibHEF/fBpyMzNqRxUay2EvvhW+2nlhtYDM1uek3kSS
ne5L0ujgbh+3Ee2UAHxWiMs3PZzNihJtGBKnhvZ91RCOsk8YK6+P1J+Hl77DY4YuansPRixefj3/
dkBaYnpFvAQpnOfIV9aipgPuGGe7yZLu1rRfxlIp3Lc6MI5W2mOPteFc2CSSaQoxFlN+jTByQnhO
Nju3CMsTlZ+KX151jvlPbgrw8Iq+m08QUZwqxIDky5MZwz0XampD6LHcGLZmThndYYVe7c7M3kti
eHkRrqrCP6VQjj2eFXwofnc9Vz4NuyCxLdAWvc5b5ARtd+3qqXZF073RcPjDYrwidiQYrrxYE4B5
mxrGC6dNlEbiJgPJOvjJHMgLJTdOITjMscDm7DIxYMUF4bZW8G3pWoL906zFeM+yaKWPCpk0dOyQ
WeIJ/S3xktDe0qgs4YUhfE0JbfhscFMGv67FD/tlSyGiKLe5KSmfB9cez8eLCIqLz/CXn/WG1oMo
OEJkKrnoqGZU8Niw3O8LgQBI5Y1zL0bMZ+vkfgIFP1LOZrByiBgC/7HpeTfU92GS4Hqz7vPYSTph
gilFl8xFHErDH3jGUM7hvjX1tqzFpXJR72v88hxC/f7UNCgbo5qIgV5xDDRLsCW1z0uS83HKpwPc
qO6ySJugICJdsJ0gvvLog4Z7lhsgudVFQsH7f+z8uioqP6xLN2TdcnP0SZaqv6dW3/JvNst23q/t
nIMRx4PAtPeWiYJKrdFyNm1w3TA0IrVdX9jRDSd/rER6I2Mx8lpzlDlI7xD+AB+QBmJFqMyTn0t8
IYAHRnvebxs494gs8vcQIl3tI0bELfdHXgHeQAcdT7v0US7zh8nGu4E6H8HjSPJ5TFLAFuzavrgB
B+qDuSK7chnnysWo1hmAVuSNggGdY0rNkeMMXmiCpgXpndQxKLEB0r89fZS2ufmiqpcjlcHXJKeT
zuZ5TblhWZfPB9wOjAXCSDU21ff8oh5vyGYYNfeX3St0eCKK8y0cIm9GtnZmoIj+Opz/g6OxDSDV
g0mYMZ5idoBdFV3xEZs0hx0PMUnQE2tHjDW3LFY4rQBVHFB7G6TmHhb/tlUvDd3f+kMEmlmRlZc+
0QBk1LzIb/Cqd7h5215Y5hDOAwKfNidU72K8cVJbjdWh0Dh98RtO1w/rtRtm6maMxRP2OUg7AZ3h
7jwV7PMgeSS0eu9gAOetYFQO8ISuaqNVbxHTNRVSSF4iRRfITjwNitVEaOk1lHz+tPYNBEKKx8D4
v9Jtx8FEtuvUWtLAWpIrSFOfs3EgePiJy5EUt+NyM+BfWAxF1HcSIGxQKTew75+cBJEMVy2SOlrG
6tots1e1chfsG/M6ajgvhIEsLrUU1892niRx7GJnBoCHfAleMHErnGqvyQVyn1cxk+5mfYVEIBV3
/DAcTSCxOreclihXx4t6p4K2KqDUwuCor1nAarh/2+Q6MtJDYECEcHWcoJ3TPLBknAqOZSJlzNG5
tWWj1mNAZqKYBbsZj0V12603phUnBqV20GlvaduYBcxhRdU2gCMad61SzPwo0aF/i0cdrlYAU/5Z
FWsFjaQR9IFiS2xDpElQ0L9MNqHpCRi8vNJqXp8QoWDpymLvRcOMasRvOmm0KCUOO0i8AQnk67pD
Xkzlf21ngBTqa5XNz4I4RuI76MeggVsf9AVHXb2cC5DHD89DeDYfkD9AFwEJG+TPdYIcQjpXJCjM
bBULG46QsBrssbiTYl5zXgNzXblT3sfZAg5HW3uL6nDOZy3AQaGVMxPBs1PHpE+jENFZ6VoqylIZ
LdUBGRYMZN8bTt6d7fGI+ryv8YUrdO6V24QHYbRx6X01xb62iG00fAKlnuCm0ZubzjYd6diIBHu5
e69mMZFrpXSCO2xKtDmfeisEpOa+6im4naPIAb2oOwWPCWl2Zcsrfvbd3QpSCBRVZ0ypJ8qFjXIV
qOlfj/nDcAXUQUw2lABCl1OlwjNknkIyrVGxLKMT8st7Wse6M8RejiQJVvaVzAUCO+u6+Z1d76cv
jkIV0vRULAnRzKGAOdzfIOKFaYo2jxI12cs73sMVHydPu4EyVFnx3m6u1314RnsNuWPe2cTAv/Wv
Iy8Zi0TqYCTO2WUYiK7UnDvwX9sEpV4yivOL5v8VoW5v92CDAFM6ZBzO21viaJ5tdxLoJlzaGTPz
b69DnLjFanDG0/aVc2TS80MXBYb3b3BPe7VcuGhMqC+u15CgnqajlsaHsjj/ZaqKJTXd3SaJ4D11
weQ5mm0N//OGVfn11cCtKDUhNuGhO/T+nnu4lmr9v1mWNfWah1SPJ41U10b/Luc6ZpDsSwZO5XKK
9Y9xgTbYlYz9s+bsdEpEGHlS+9e80fPEh0/Ra3DNj8aSIZ7/kWvHR/hbk4fTrrPymKnVbIb/QlVl
wXOTvkRmztq6jDBC2UrRbC/Smsa4kWLootHnYgg31s4E1OGARZnxbbXN+IEhIL4NgdBNwBmQG/Vr
OX2qLm9S1Aqo2RpSB5m+ZYaJU+7C/i4kUymlPgA56XFfzlmcjv3cVJwN/mAAtumt4ZiRxE3XsUr8
EBq2jU2IsxW0bNXXppQdeWYOboMfhi7Uzx2pBC54xj9E286ehZy1c2YWPWtZVbCsHJ2wRN4HnSbL
IxA+C0GF0HuXr3YgmOgqUkJtSmhpPnr14TAKSUJmQ9kir+G72GCnfHewLRDfxUeTYGU2soGsoRRT
N0wX6Pp6fynsbf+JkkzLKvF001rYoK4q5fVxXhK0GTn75WbcfjzonEWzz7LlkBedRCxvQet/GMAl
9vbOqvz7VaffVR7Y+9E8xmFnV9CAXkWcbbAMCcflvQJB3ztq2iPfOeIt06EZuEtJ+CilJZwLjqtV
/Aerf9WCF3bsB55F01sh/LWIixDhTzxYwjFD6DUZJ7Kx3UL553civjY8kMKMw/tvzRtvoHEexl7m
50UHmxKAWqaFTanIgV+QFBcHJ55DOVdmf6dsRp6ZL+Flt/Dnx+vnT4922wp5jRQev0E5bZ9ufYU4
HF56z+s/AX/ZQp25fDxj5qFDPOEv88DZnl5Rg87uIbBwO79KFGghboMJeVYca3o8rL/SBLUEu8AY
n1nvbifAFK0sFgv4g+Kj2smFUt7033x+3jgiv452w0iobqCxb33ZEWbIU+/6/0dJvyaWcSGpz0lA
0ROvDSmaRiQu7hlviBoZ/b1t0YdpXllRheYAa7zYAPAG+VE3VtuXDxUQLSrNY5c+YTL2Xi0vMDyD
Q6J9yqmi5UJ0sh9WPap2efsrh7n+gpg0avczV8Muj0H/uWwsSa/CdR9T9lthlYTW+e2boYQFcIyU
EHKVpf+zOqGO5aendkn00Mxue6gmC5aso3qN+w3U5szfmIeKKzfFSQ0bbcK2WXeQr9bLn0svLMxE
KBBdA4jb3uTwedwBaKfItKQOoDrKVEU2ywIcRtjixCPn9AtaOhMAFKv5M/UCJID/06gfaI/aP7JB
UvRbiefPaTD65IkJFJPZc6nxVmxDnJ35E2F3caa18cyesEka8Tlwn150jKyrVz9/hORWOPMmRz1t
+ovlpm3+KyoomCIjuPGJpjGRPj55VMheP613ut0qg2BJv8lYFz6Sg/c9D+CR0FT3hbM48uI90s7D
zh/2A+/CQNXvd5KiEZt9IsbaIyq7XlsvSixHoA8jhMoOes2pwVlj5EGKd1aWrpE8zTO93SkLcJnW
yoU1R656tCoRd9NM6+St8FjlJ0whzNxGYYk9a2eL6FA4mVGubpohB/Nct5fdh3BlePD/MSzGOfhE
M2Crz3xfN3ro+1gr9r81nYFdLGhjDVbXgiUj+LLLqnjY1sbIfKThtwF0rYrWxUut9CSvNaJRhQop
BS9BKn1wO9f/y1HbNO93AaP8Zu/3iItl/cCzoW16qlxoCME1MtKGmCR8g2xor/R3sjdFpUsuFEAh
zukyPAADqbOhqJaksu1ykGofqAG2gSf/wQS1Y4JAY5alGlhcjtif4yr8JHsPXQvQHtEloHJgC10j
tVySWWZT8Carpzte20uqIinX1VxlmEfmIWjS3NL1qH6cHhilUS1SmzjdsHswgft7991jF+6B5368
1Yms/9WwDqG5Fdj131VAjuu6+JrUBnBOW+G134MXM+u4YTqEGXbaWbMZXtVFcugc3LcU50F/7/tp
jbFokXtjWnuMvZ3wiqdH1/TcKDEgjrbUnsJVBdaQLwKVDBmhREyAhO742xC7B77Y4u4q8dKwPLw4
YgSvo2O1k98HA7rZAJSulLkhd000TLK3tmEXrHyqRCSzCrazL6fdCFPji1G9i8YOC8FfcpuxtvIj
pReDROBkeYqaEDQneGnI5ZdfKQPnVY/gg3CwNRyRsEQAvjPSbvU3ZbU6MltBP4W5y4nEf+Rt44K9
ijJNIXEo9SfB/4D93mNNPY22r3MRqMrl0DzWfIo6mt2dtSehGCPE0NVRawXYGoVQzpcK2zg0zPhy
G27zNvmG4HplavJrrOFQnfB5/r8vp67djTKXioFxI1kQoLVXFQMBP7IWHRiruYClZY3w7fuCj0gO
f2kkw3SP5UrQQu3c2amaT85nVJ/MoZHWe7KNDjVzPtyn8kgErtTE7GxdMuSnLQ0Y6A/QUWIqRjOQ
xY4I3QtdYu9k0PdK/IoFL6Rq1W5MZwth0mA6vB4AHmV0ZLBltsF9TYgDVV7iJSkw82ud7yKTjQ2N
Jqvp5760PX5RNhezw9CCBKD4Te0sF5hZlUidWGOprdLRSe0VjfZmdxMnHuLB7fthmI0cTe0OmOLI
/bCCpCpxSHSLFrkaJlwLaFvJX4WQgPIUdjhX2s3zPlCD3WDkAPE6WduRth3cN0sVGadqulOYHlao
jodgb6OYx9RgoXXyOene4oV0NqCMzVCJuKl3kO3F+wvVSF219srMfCftE2fxGXw5M2L4p01uLUwZ
MRSGnXf50P/Ijg+kHLMzWaz4fAlAgRFBWPQUKWp2GSfUpuhIwtIQTd8rWK3uot/qNyv5pscCDZYc
PS2qQgqf+UpDD2y5vfdaE3s/5CeTbj/y6KPsDf+naxqbnM6l1Zg5MbSMOnwXPglSrELGmWBgLL5v
Vzg0PDur4i6q7vrFoj5MVkYX2czNfHTDHp1ql+05n0HPTaJFUGYo14ur7hpvFfkEz3sDYAI2tde0
rVLSCD808K40HBJZdYOoYgc9yp8ONtxV8IGnT17wh1zq9ZNgegRn8uNe9g7I8aqEtEwWYjbA1Gi7
g+7DwVmMubyPTEBmYtvv6nnvZGokIdYwGhykNKupzErTUZqORsoHzZlM1R7u3vdUjxPVvsEJ5/5C
ALI1FB/9W06wV/9gc4k1aGSyihDm28epCIOZxkJyCwvNSw/DgnqikuOyD4DX1VnTjyxOxMLRO+Ds
KJNx7sriBWnuxqEXt5/Fgy8rpL3tLq+BZxGnr3vSHk5OjZB6OIEFoM/ujonJnVTDGyQP8YaBLbbG
5VDUw9CohsiKYiHyrzaN8Ulb2Rmsp4Why2RQrrZ7+gkwpQ0GwDHLnPJDyKb7bFvwt+4EVkvZ+trQ
Lv2yt7yDJweOsSqH7l7RedocVxcTSHTEGpWsXluBdWqUJtwLRDpvvF50c2o8DPPycVPrYEimk36s
tTguITztRnlD6Kf5RxySl1oePYJB7pGLqwXzxS2Bb2H3ZeTf15WJGvCsraGpH2tAUJcGc7MtpHQk
VXWRzBpLtRBGTnE82IfLIIW3BewSddyihkBUEH/Bl4In/15hDgN2HxdMsqRzHMY4r8ewx8lAl6WL
61BsIQnDJp8YcVF5sEdZwGAhHjf4cuIVcZXYIUcP65OoyJefyq24f9miEm1rl3gExyAVez6Fe5+q
hvdOWdjnBFnM+OoFmNkmFyMiBiRIFvZrQFKDJTTBLsp45I+J9ohGq9mrZtipguonyp7BD6KFP67V
nnxzXHq0L3gcZTR/K0HrE5iox6hoCu2/tX6/I5GZ8OgYZ3nZkrPtXnUX/I++5UkbmOi6b1BlTVai
bjsIM5irfo313XdQrhd1xspmrTIs2CLnAaN8mHVcX2tklA8jvtcRrhf1uVz9tDhmiNyYQxjpQsM4
a1uXJYQ+kn6FDGxjlw86JeQjhS0rzb1Nr5oDDI32YkjhLCegmYsuFKao5UfzVh2HOJ56NdlF5n+7
7KbJteUlxvnQakjj/y+Xu2bcl+yguqkXP2M0bXfRdWVbkFeTMg0j/lsD6SwQTQ0UVcf5+31CUB1c
+aVLK4RUSPXJkG7NVnNZdOg28a0CQhYszhbyTli7keKg5BNkhPmCkOun/L9INei8OdMDBS03/MB/
b7sisxwNvpdd9AUxJ3t4A+HQX18gxNS3gCp6TJH1Q0y6EuDeUNDtBoxtT/6P/G9QNEVeZh/IwQ0X
sTGCjq4k2392fELNjJ3arWOV4HG+iIU7QKmC0O192gJZsciuh0TWzv0iUuXDTxumclrIaMpvHW8W
7afRO6Qe8B/FhK0VjDj5gIs5IxBfwUdJ85LdOa9lEpQjGmxQuo5+tDFiXR2hqjY5et7cFvI7FNUJ
ZhTJOgSSeMZWHLWI6TlCrnnKZBIcPU/4J5QVnqa0m/U5a378UkPMFOE29DKRYMPCOKit0MEjyYjo
1knKOrUnWBkFAO9m59mYEvrG8+NmT78zj8A87GWr5+lH92zR9K0d88A/CpBvyjlk+Xu8xPvmzyiu
diwr8SWm+SOjkNf5hMh5t8WU8Pjp4XScfxIlXdsaGifSeGRLvJC40RZ1ENFOJL3E+q3fGAANDNFr
3uYqxrDlxvLve6D04SvToGL3UMVSDKC9DDsUWFmKA06yWiY+wDZdKkqdaOUOOxYtrjqF7tk3q408
vT9d6oidkgQYX1PwQV9r0FlRqYEPS/6artjQej0JYx2NW8J1lE7ZXolFuaXUF7e6OwCfUCfN6YZ/
tBzqOJBaMPyEeUlHbnsdfOECuPpaOOfapttAcvH9H4/rEg6upNmBJb/KsGPXBz0Z0izXMEbdBsEV
/XgrMhdCH5MN/Wpdtz5hdr22y8hiSSOzC7Blgb5zIcZHS9mf3gwqPRq7pEs7G0oEYmHQonLaG2Ml
dBQi27x9GyqmE9u+kENWLCbu1hNeAoh94jVF3jMBJzs1YDNeNxtDXqCvrTcIAUeE8bqi51atm8cO
bJzPqhytCwhqBKuSPi0EcgoZx5kgBI6y5UvaOmhQXmCPH/ehGJsrAMkgz3gEFX9lCt96HNTXbX2o
jZiK4/Zea4Tnxlbg6R6yLYi9C3ev2DigcQvbEysqUv6QVJandUmfKgKLVJC3n0k3VpgN77tRkmuZ
4EN7wGLlssK9LT7qXSYZDpm1ng0d3DcSHRp8WZNlm7oA10ZGXFWReRH0TadC5EJUyRyCfDphNfx1
NZY7UuLyqVQjcw4T6iaXLdz8bWSTuLq1iJrHOpRAKVEcayxI0G0x4gX2WETxjbbrCFuUCwEtc0sZ
ceGeAR0O8q2cPHvioZd80crbdCZkVAmrzQyu3dCJh/CqnfgeCkaJLL/p2ueIiV1AA+JlwvdoKaOj
ntX0hwm4KI6eEf4f3y654czI966RyiF3vqosslGNJBy7Z4aMeACAj4vZ8nre1HrCIoMYodm6r9h/
TnNNm+A4lSNUSvw2WQS5xnau8Lkn8C8WLRJc7FvMBzC3zGhsdLwfhbsOKOoN3uA2ip58G2CKAI5X
EogAZuDKFZ30BwwSpwkojEsoyaD1Fn4Jx2FBj+kiL5a6YOPyQ2968N0Q6uJNWPmA3MsrMl6Norcm
sRwDCauPmNrtfd6mfJa6ACByrySuFmCnJI74Ea06+JXUr4I/plapHMUchnAAew6Tmwi0MrEFq4Zu
XqEFjYVMj6Bu1YOrN06jvfbTn1/e24RblhDIjaTwIlmoptL/mm1DdBEqTJYXKbcoIbyN1eQV4Ej5
bDbgO9eSqdyadBoHBc+LFyNEJ+hQ8XtpT40ciMjCiYq4nraHvbgwaSMpFFPLtNRm9J9SNA8Y/JgN
+AFkSxvez9Lm5am7xR5rKlrvamVqFWoh9Nq7ml1ZZzvF5UJn3sP31ffm09Pbady4aMeimDo2gmp+
svP0qdo7SRyiyhEL6RWTscfolW9tTOIO1LYXxCoxWc1knVw3I5KbZImtlcZRVdB+JBe9yqyhHGt2
8FcYHXZP/670idLuVFEnsX1Bar76sRyKn7RROWBzlzxG2KWNgCVhxomsZJ09mngUD6JBuhwFSnij
bvyWh+CWsXmGg5ocueoasDeub9xCURgdqWeFIIlY+osgOdvT1oyRRNl6P1ldAsWnY4SanatiJqzj
kuhpPiV76c4pb8DUf8G8jiOjvNvCRgfkAnqWDNWZIWM8KiuRLbsXNpejMGTl4Zz1dgAh9vOjgGTz
aH5DsbDg777zG/rB0K8xxfQIVXVT3El9i3ygy2qdmf/kap4FE62XUJQKs+E2H2NVMEyjjlQiDYr7
CrRheTe/l4hbmxCljNOzimlqhBVmpmSjZ2tUOYyqtE29LL1pH3nWnSC5S+Y0oGHqXhMYX2MknQVX
6QlqnzX7ky7gYH4Jine+p4KM7A3xz68NYicz3ERuJNEc/lvZn7ZJe8idzZ/r9eKo1tXFRML/KcIE
0jzGJae5YwTRuAXKnlMVYhpfneB87RLXrK+FbtJMpuOc9yD1XR/pZ/dl21wQi6zEXzP3hfiZVPip
EC3PQzwqu5xCPiJa1OKjJ2Yu8mm9wsdkScWfo5mciB/fOqgVzNWQwhXd9covumlL7xzNus0i15qo
PG5c+8zjThmqa/MaRJc5WFpCwcIkZ+Vxwtvdgidc6VRRU7vVogCXai8MbG632U4AUYqeqmcotGbo
9J7jfD2BUQ+JFIoj9xAe8QyefgXRzMyWHprWXP93mJtWcpR4HvOd9ZOE5iGdDIC/xEXuK9hfBtHi
tc3DfAH55Zgt2ZWNu9gtiHmTXFUkiuSwhlWS/BTe5b1w0uAvoYYqbe8Rf0N+8eBXKtq6jZequFnn
sVzZZA9V6VNob1V3Zkx5wcU/+Tevlif40GqkdNxPNnI0LC8yQ4TctrOmpmlGYn9JAoWXrmC5x3Re
0v0RgxzB3U2/Dk5K+dCRj7gcFSbBtcOa0Zs7vemCedGcUCwiI9lkx+/Xh/xPDKO+ycs5k2wU2RYt
dTa4GZ+VoS7MLeZjoSQ8xkF9wY0CMfelc7KCJMn6y+sYdgLok1rwEY4iEeir8x/sUyhfkMvzf6Uu
fbX7BKoMJ1wnBD/Je4uMgQ+bNxTtlr2WeXvWC2JDYLfbqipCEyhOtjKbEKyQj2rLIkHkKnS07Uw8
jMEVvTTPqo2iItvBVTZgZ2SUUY5ExJVxRIA5jBV2LlGefOr0CC3qExF6TQzWRVXsODIDSf2KPvT7
PETff9zdPLWgbWk8tMqyOI/MiBT3aLaSfD7wRToPKKi9gCNZ6H5mwg6IxPtPfKFXshKhVbTx9fc6
XF8Fuuzdt4ESDDbf6BUdHc5api11ZNkW3xaiAg1nSSFVqPUrGTT/hcQeNHBrqt5wdmuhLZD8bqqd
fa8GsAN1rB1wbQpOgzAlE07aprqG3vTGK7ImR60CUvLDogI2I9Y14wBFaN8nWiPZCqD3a5Bec6Wd
J63tjoT5vmAicgg4gL2o7xY9aT4O9PhoLmu7GsX0wk5eDOY9PgAhu0LZKmnXzH2bSAurHeyDxRxR
LPTKnRxN30m+0uEZpMX96HOOo7Iiuqg9Uo6Zh5urWdvWlD1pGJkuNGllx6vuHeFrSDcO15ig89jB
5nBJg5LRCVPf0q3bCxaM3uL9uz5OM42qr8KefHoaF/2105LkvVXi7N8Ff8IFBkZS2MS8snIb5Onw
/hoyidqr7AvFi8u9JmPGPscphoOTw+JYo+DO2y45ohNqnJEB/79sfgckfLN5ayYvP+IKuZR66NpY
TGkmdfufmgkjx4HdF4tdn8edEi34vpp9K40uO1oP9ZJLXxeRJfHsHRDzoYRmsTnpSvMu5u7z/ka9
rafokX/WzN9WQ8E1JIz+Ql5WHXT6yO/XloSkVCP+l04PyvNNQWReDv0TuPafQ+YRqQQw+GK9yXIw
kIaafKnidVqsdRee9u8CrPAdI/fGFi8wp6JTlM+VSrlhcJgchlmwsN/MssX6qVd3LCsEv2iFMQ4D
Rg5QlsLzPl+uus0ObZtWTUqq6f7ah4p+1Jj19u+Ihj3NXiybpwwDV2+qYepPY2Iv0pKlbGjt8Fvy
yUHfdVybweqFS5VTFDbnqGSujCzO5Yb1fvybEzgRDAHEskupHt1uBNEs2WaI5iWw7nElVwTeiO4V
CnWzfcvJ+KIY2pIjXjO5r/P2i/zRxDvDrqf6/NmLkw1zVhsdwJ/rlXmOVnrJsfeV17jjk7tXt453
wNuS0padUFDfBubF+74ER7jB70YQ0XOiVkUUnVqks2zSwKXR+TYwWXNiA78Z2NaaIzRz6rLnj248
iJYjUpLSltljRGAY9TabX5SGTi4l0tDpXNBCcT51SykZKaXTTuo/lHpCxZerZeP1Punvxr6LMlqm
3pvQjVY3V8TL0Bi1vd4oHbBOrN5cZVpC8YemDo4UxOhX7hap7aZ0sLZVc0AJsS49Rv9QsvXgdv9N
nfMu3Oqvh5VSuDTj4p1cOKSr/kUQRKfj+BMAVZH4nIyd7os55Eyi5TFMgeJ64NeX0Ohpcn5AQPIP
eww/UVMCCHZpCeGuduzhvLXgRRiupKqbJtSAs3Aud4SpZgQtP8ilh1evmG6RRI19MrAGFvQFE8Xs
iFsFgeaF7CDqVhE7LEG/i/mWiE0xyada5aydKIkqzXESkz4k0X+Hwl1j/SKiUnIbfmA1dgAAOyuV
P6HS2DAjGn6CPisEDmXiUEaej0+iptP2EbGnbV2GbujX6AYm0c3UaTIzB8p5VuMmJcLJGQZU0NF8
CjP2WiBwq+3Cm3njY9dKYCKQaFsEKYtZgPu205dlnG8jPxaBAALpj6hEE8GjPWXuDgQDP4fPY3jv
O2vwkwbqb1KhmRcU0sHU13Goit9so0Z8ZaHPXudH9oveYzQWScmOUPANkTbJbRWPuLJZp8CRzhXi
f8DxPBzMgNz2gtyNEaNqY4S4dROc2cT7Udy0MbONobzBxe/EacoDsE4nsRhfcTktcA8TL7hdQ+FS
zRgqscxJoTAeMSh4KYZunwh71G5w4N9op0/DRRiMmfHuQMNe/+TZlSWhFm0W9qrkvNsJLzusKIBO
gelKZbnlhBtb2A9lmdcpsxzwsE+jkYU6eFXURjTHrIJQCHBd+xiqM0Q+6JOhuWo6vMHjGYx2S6YC
ro9XLjC92TzewANU+YPdkc1ySyMLG+UlqfefVG7g7Cp9OclnwGmm/nSVt/I4YCGCRLSn2v4ExVns
xFh/8/aLvKEzh4r0aVkhu0GnE4G59eCwBgH5jGkJGBS7/G2zDOYF60EEUz6uArBKqwTZ/xeULCFw
Np7iGosEku1o+OkOnEQHDfa4uQwjNhybRwio9J0HUggtWZY1WaU+0+BzfjwbbGqxTgV+7TZIG5jq
V8yx93jmYFv4DXne7E6M5egOYOPYtQ3eR7ZfuV5e4cIg9q2ydZYKeHaEfnlmby+yvyldHEhjYOJl
qpJcke7fAfGq0A2XTdXnSZL5BqyAUWdzLdWgtiL/0EmvjgSfYSr7MFiSh27arlnC+NA5xCF3czvB
pf51pgYonkkGUPfYjZIzCQw5dyUoEEiOg8+NWhsS6ff3Bx+Oyu4+q4ZjrMt51zhJvC8MGknx2IAW
uNyjnObLTkXGfH26ve2k/l8N2aFZC/REUjZBqaonApL8SWzWAqm8F9KKq2/xF5ceByHQ8vW01roO
E+uLzFGwkLA3vmItle8V2FcvyZAW5REPtW1HHlpDs5tTEB/MLp2H8ZPwrPIZprvUUr1X1JWWnAyq
y9daubZ1oxz1Tcfc1YzYMUWyK6fxdhGcGohvtkJ1vuakFpwh6Gmy3sUfbbjYOyVPorqsCnmJ6oaL
Ggw79GJ5noQVDjVRhS/XdCigA1DoQx/Gol/QjWCawhClH/YQa+3cXM0jr9jC4sLE3fbduNph5ZI+
2H4BdHeDDBlZOTYzdAUzWA5wnrs/nDNftsOzcSSZ93CXW53+KTaiMJdVSoctBu5ln4PUP+Pfromk
exIv6WYlooChrtmztdU9VAoR+VlRygedAvV2Zan4MRIr8X2NxwJ1cu13wtU8K6ITiRZt3YvZqnhI
q1wVNZGpVDF2GSXPmnX4QawMmSbVWHztvl+V691LIImMeY3nOVYfSCf7TPmwuDZIWotCvuyzLrx8
xJ/mzeV5Sh5Cwd/KgNKfXyRJmBzn5h4kSdl5DfYqw9Ud2mu8taMjJKqHtpIhMKBnnFHtG5b+19IQ
j353ulHcPzhf2qx0HVOoq+QN/Mat1tlSdDhH83Z2o7kxaIuuF0xWkRh2r05I80EetZ+0rbwjDlhc
31WOD5kQ+nua49gqqEQrx9Jobk9Q1V9ovKoDkWT4o9nGNxTAJYUWCLeptzuP855QFvFCieVWnUCN
2X7t81fjwZ4XTtS3bisA3oIbaf2mZmnhwl/FV079kLEPY07cRHdghBgGAzJ5R8eV1/ZvfHWJOY5L
RvJy8vwa/Y+MrCLsyQycYw4X6cpIEq1KYNu/nDL/q7f/Zey9XIpoyAjZbIf56QFdho4bBwmv1CoN
ZWeMDAlfGYVoP1gDV/41R7ibw7+zBeLbtHmT3DF0P1PIRX04IIgIFalGmZsHCSiAsAXZj+8kw0pT
kXxTzbU0ddAkh7KmJpN+Pw/oYnbULMfWwYlBwtgpFSKiuQOQBJ/i16sw8KrCjFJfs5KKQbCEv6cv
wEVntm5W8e+b3qAIHRbf3bH+HlmrwUOe9Fo8vS06sHzOKdRUhylx1A+8PYzDT6f2cae219ZEPHoA
25M8y5B/2K57iW9DwPB3hesR6L7V1q71XI7fBAzbENTh8tepZAaxDalMtoXvQF+2HBnBthok9Qm5
I2l3ajj4o3hmsat+H3+g0r2qt1vQGyrC46PJ2t7WMWvB0DwWeEQ=
`protect end_protected
