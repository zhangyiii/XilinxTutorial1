`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aPkk/LZprZljgyNzZTGF6gcxBz
LkEl/7f+3dcASD/i/KgBKq3OUZC517cIUJosom5xIrZP7ogbipLoucJRrZx4D/63Rac668WQR2tt
XvXehOwJ/AHEp9jRPsQutrYAu3FxtGUXHsjpDuvlEQWTsec5sqEPiTB0mY6D9KTNmi47dKqUZBs+
tiYcW3MN0wSJWz0yWRlxkDOwIe8+BZhC6+qQaKz3JYut2IWLtkVrNtVa7iVztyRq0IT2GGOk9SRF
zTZkv+gi8C2R/hrHkTCKcdU8xmWsQwsIv2Q1jCBEOLi6wOOosy71Lb5Ha1hxrI32m2Piyx4SnJPj
n0alaIYwa5EF4wS17Evgj6P25nPfldkUvpg11cL9XFhy7sgEDKefrr22sA0/VpWWLjshH6EftVjo
7Hf9nyRYEdVapyPoEuQtTc6tIvm79PMCT+E+SZwQKcnanExfZ6otWVGF96w0z9WQWco3ELpYCZ1J
+AdiwlLaM9oSfzThSi/jCqkjP0P0pl1PJTenRvHceFK3dUVi9AwxEnUSStNItyWSFwtpPhM8Z2be
Hv00vEG6vQXmfTimbRm1jCp+DuADtufxpcmxPkqMwMXKZZ0EoY+/Oqavo2fwwP2ryTV8RP/939vZ
N6JhMaktAxeu1pM3CnTA9YDhKlnNGvOzv5tTiJXC7gylsEhvN1KNnm/fDH1VyVaQcz3lAdMu5FNG
n/wc+JiSvRjuUY2CM/9JXsljSkRSk+1YrJClkyKsQLh8pWQmirP4fCWPXtz/GtXQiL2TdjrxMvOS
uKAPiN5GCbbv/3rIThnX0eVkxcqtSgccb+M+eEvEAaAHHdQdHc1a/KIsoofCKoNgXhQs/r5l3Hbt
Nwaxn8GrWsqeZlhezEfIm4h04cqMp3P+D263KmwjF0iCoAjhVA7O8D2FZroVsQEHPwrCZO2BdqKP
JESdF0BWIBuBbLP4uT6Nqvxm8OFIxkgz7s0KaohyhkPd8MS+5E14L49jF6VZhJl4RPPxUTXXRvPB
6bcmAfDovSDKyiRD++Uy2U/xTMgybhiAgywdOdnmaly9s520Py/KUqjdIO8Jw0WzoZAdG+AhSZy+
jOCZAtbs7UtsHmVqeyjy3n8Gd7kO4EgdiPLRJCxV4BqSpbqlaLlnxESaN7Og1mDdQb7nY9U6817F
G0tWKUi3rBtn4CJ4lUoTpOJzBqqp91W8wKUKfHjWa+RcOUwaRBJKTXvMEB+QyMlCcngxhRO8iFuA
vWmQ7ppu90QnuRRs6hLLCiaY9GdqtAca8q28LxLxBQDkmn/I62cvWM884VLSIRZSAK/DkQOgdVSF
qq6UnXQBlcfPPjYpCGL35Po+4jFDophkxI5hl0vx0+PoNINbMxW6Sgv611+Tj37V5ufsF5xmWaRf
NVYyCyY9WgE3yeMdzA5yowj9/PBFM2IYYQfZLdPMRAqMo/+KSQxdye4ZP9pn6fdXjo6H1aa2/HS6
Wk22Q4Y51bZyfbtsmDZZhulQvt0fVsj16NB+lbLHhsyISN2J1hR5j3zXUkHQw+ql57El5w9e9NaH
1kfTu4+orNjoeFouZo+xOStzfCb/2+r2JYQxVdYB2UX7gTh2+4RAVJDj7uju6bwwJ6iPKf51p8Bt
E5RoJPzGgy4O8FihSOQvXtffu30vBmmkZFx9Akuw1D3rpWYDmhZMNKVFV67D9OLvv6gSTyHvQMTD
lIbKIUcR0BZwgeOdXpduN6Dba6gKQnfnfE3oTl7MBW8fFknHrKLYAcFf7d3kDl2IA19vybGg941Y
0OV0i/wpGMxrWn2epjateQG+9qQbs8lc+Vioh5CIVlSVDw69DUshAaYcKURRj0SO0hd6y3qfdCTL
2RggY0OtrI/0JYVk6p1ETm71ZSlMonp56L/d4M6caj+JpMbuQswziTYJ7fXtQG0AAIe3F1RdlDmf
w2LbxXPsE8gvHjQI3JeZ5Me11+ei+90vUQm+1dFBUMggWSOzhohGWOP4DBRt3XA2RCjTXUDQXJsf
5tHKzjz1TzW2krB4lPB7d07vMNI7DPM0aZ3XztW7Jw+xkYElV7vMmKMz1nd0Az73O5smjneNpEMI
DLf58mcIyvWSw5eajT9CAIwVdkvbQxfGTKZGdGwHk2wJL8py2xoKQ8IZkBkDYQSL1+gUn8KcWlkw
Z8so7NHwQwJh6i1XUZUBnL9A+teyhOQla6pEdIzCANG0J+IkDrfT8UpLfPz4yQTQgsyLmvbPp6Qx
jFwsTQt8OXu2/7poCv0UKwYuA7AHVfZqPoV1yzAYEZL+xTSis8MMwVqpTxYIO21pPt4eI54Y0sMg
ylycsfNowCYSxKc+9IdlySefyorHA0V+aFYTABSq4UXFowM7wZRs/1VyZnKZJpAIjnlt3rD/d8y4
ximpTa+Uh2UCO+GfH9XMHIMVEGCwVsZ/MvNh/pTWNh0YKHnJqyjtrA/G+clmO30FP+P/kIBBqHGT
9HBg/npfwVV9+fn3CSAAZ/Kj/rGrpUF2be9znnqm1Y2jB5cku5UX3a6eXxkwVLfMuEuLfcvJzByZ
la9gH/VXAM3frasuugoGCFhZvNSCpjmAMmcixbrgFdUKjcigEw7aHRzElgs1eX2iToW7/jjnVU+9
Du/x7/3wLpmbn78PVWrHDYjoPgcw4SgIG0j07z35lcYyxQPx5Zwm2/m0FLzBwKlzspsQa9oBl599
Svg6e6D1WoE2Gc8hqXKMbRAvB4mD6fGPYzLvvv2Ccz8WEAg9eAuvktDLVHz6vbzSkqPAH0q4mboe
yi1gUNct+ecX5mOyS+gc5MiyIIWfW6oSczaaKIAelGYZls08qBF2XpwK34XzEj5O4mnVQP3kn1ko
fYdV5yiFVzbDHcFyG+phdxMqYCtQoqrQqX4tCpvVv4nq/vlLUtDaAySuRFh3HPM3nizMbglhIDVm
6N3giXlxHRJ4aK1lfULcA6M3jbEUwW5v4zkPQ0g8qsnMRJB80wWFXolObMOkLlOe8GuvU13rwM76
lpS8Jy4tq4A2e5/eaUXoZ5/0+uk1owrB/PUM7JUDtkZtD4UUAPOUlysbxJecDvCEd1+xjvK5gK5S
cnf8SrVOneQJQiJ5O/Nn6oQY6S/7jX06OVw4S91h1rV+4qubSaSi/1pdIUpWu3oHxb36TEmVJFUc
1iOkWnqtg5RlYrwhfeKAvrCbH/p4v+Dr5O6E0vIpMh1WBYD8tEjGgqsg0lZlo9V96PvPP5WextoF
PWCqMC3tQ39qT5I9dfEUtrMokdUP+yn/LNR54NFG22iU37cXN5AapRKtutJdPt3E0T6Tb1EVhE0f
kUllBhGSoW5rpjONyX9Xv0NNrAZ7n70liRkcrHgn19OhUNOoR1im5VoNq2mgotV0R7obyFnYTvxG
m9akp21ITeWhNaqyG+qm+uv+5wX0PzqSDUxejfKkqHXc8fATwXI1yUKUJ8LkhRW6gsYSJqmm4XHH
rhDk254i37tUpR1zgjnov5RUhDQdbEmiW1DNZgyGTeaIDP1O3qs14Lqx947N5g4iwKMCkaFBNWOw
ZyBZ/jAaMscMmifltLh1GRP6sO34mkLUlh+JmVoogMtDmQTYIvJECpk0dJjrFbCoGJQZNyhFKrOF
zmF6CEGsQfKtO6S04m5K6h1U19ilL8wlQkZgz7GodQ5VFzAb747RHq1vZDc1IC2aXwlpbNvXbBvy
VtkMUXAF577/v2QByJ5JDu321TcidCLN2b43f3DhtyR6Vz7Y5XRf8czEpFBypnF+HGNqSF5ssrIB
Api4fVrd3hmKZzqdzhE6NnfQKk5qymU/JXK0Q3GKGEvLhb4NyFMjTMT8+w/lOwwFa0kh+Gm1JIEe
80k47GOHirSUREWdh1EU06Frda5Sa2ruGCDxmSIOg7nj30s0hqs6ckF/helao4rm+xHZOFsyxwzD
w+l1WqEI23ptTykeYfOCyaBTMh97Hq4bQIsYGjHh4DRadOoyuwsSeFYueqCMs1PrlLMhzSoyohdK
OlWK/ubEnSp5fR/Vx02XlAiTRa2D8doqJEiDlDLrCDFESGPwL7tWy60V7XxQeu5tUsnxI4DUn4N3
B9fTV7srsSmZbEqqKucXn9lwKp9j6IkQAahMHeeTVLOjR5mhF/EVbhFGKMlW8U6ZJN9G3s0rMpAj
UvmK1tgOJWZWwLoCFM6hUc8QIyvkE8NenW3fGFbvAd7le2U1UnBbnZEsRyxlN7Z/vxAo+L+cf/uO
r4r2kt4b0XszZIMZ/SL2EaUNbUufmipggINQPXWAnn44zrYuO8y8VPALUI2w0vInK93ls1oh4fPG
HziXDiYRkpOC09JOqA7iaLs+hl/05OREcBiJjXmh54lJQ/rJk4uQO6H61FLUKxFjTeeiJebYE1nK
1WIiPe1lkybqvhKTPmX74Zk+nBoaxR9Q4nAOxfmzbJik9snEl6e+yDQEhDBarQvc4t8glluuzJIw
F+MkT4juCneslIIlWt5wL7e8MIii9UCuLIn+GfUjObQqliYFtiuxH9E/ito8FXDW6K3NlXvp6Wfc
JgoTNr9E+/c9xM/+mERmP6Sh8Nh2HRxiTpFfYLInhEj0LYo23y550pXFF2asFwy82y7gh4B9aICF
aKhyEWzBeOM5+1FSB6qVo5yD3Ujw0FVB7yuU4DiVygPyJHnULRlGnC0hZs4jG8bqPSvFGCiXsrBR
+y6lEiLujYIYN6FjG1QRdgDw9SGlTEmk/rlBruo+ub9LvDioCMx58UWQ69WmtUXaVsmawfOTe0gK
6M9rQHxSaTcynngzMZZqYNnUsMmhFSAAUNfpzv48JEM9T419iJ6rlVdTeC5pkN6QvmbgVHQ801XK
/xfn4EnAkcQbgcNLEPPb+Uz4TO71w7ucCLK7aO3GYDEwyS0yFERnghuvr2q9cdoAPHhloZoNCMqB
gEGd2Exou914q92VcSpu+pkX+xHuCj16Gcvy4PNo5aYeIpypoHTyubZS0hB5pUnmCCg9wBofCJ4D
ttv7qZ/AXHYD2e0jDxC+ncN/4qHiF2o9UAxNIXdlqXnrnbtUmVbklgfpMFLkh6Rir+IC7IYO05pE
eC5WIj1odLfT2QbTEGhZ0IhK8m6h469p8eXlK6tzSVnWxPAzPjTomDGpN9dftr0JbeXQj3JCaH5I
aXodpUbux3yAh0nTOOsEUHzmYOl2NnImGPf+xT0nSW/D9I3OCiQSgOAUzpR0edMvWCmTeTRGDqp/
ug+Qi+VRNrhnhQv3uCLgEnlLh8Ig0nXBZswsiIZseLAJ1HVZIHo15LKX1o4sJHWP93YtMDKgq2yv
Htfs5w/4XzzYpMjhh+FB6m3Vw/c9fE7PmYqpzPnf+66R2HUS9THmihsqsS72Y+t9AX9Q+5HCV4nc
lB/11G0UeO5AVN9IvjXzqkgQH1K/hlwwiXHoAWvcBdVA4oyvxjv8E8rrGx2J6zSbpBWCR5UQH70S
jy/X3NlDyeB6j9oxBeEjBWJZX7DJN7xKaXplxKjtkUuOBq9oqSiyrerMPF/R4jVAMYSeht2zSwa+
5PocX8X1dKl9TmTBjKmjH5wJFy3mrEM9ZelHd9XRQIZcOyE8QYPzxp0NYuXrlAww4sjoSIWqPW6L
gEHWL8Ngd6R7keFqq5SqPgtYFom2eQ2YAaCq6x4cw09HAKxAog9TkldwnExBMVXYcuybzTUEgIy9
HeNpV4BUbRoEqexgNHHLNKLcisI3KBM/3h8rlXwar/armCooAmsmZ21KcI2MIF3dbMpzMHhhYUWp
zVW0jbhyqqyTOFABw+a90YxIm/wY42xs6TFuwmGLu2+xX+Y/W7XBtoIbaJtpxFNALLmpuW0DZuF+
O+Kv1DW/Ur1ZDSSMKbEq2FaS43WlxWUlDBdk9Ac6m0JcZW8W1gnpmHBidwGp6qUMxz+utYI42EO/
xRvFZ0ekgNzu37MkkBTyNnHadMBWqVuTWm/rXbSDOSRonQvz+RO4ST1eQ2KYbS/47pv4HCgjdJbq
EvEJVa1wgX+r+dNd3WMwvd9xXN1zXoedUaHDc3Kp3mKFsBug0QW0xJGdGVyS33T4CnW6W1ngbwKB
Ncp7lI+IodcnTyZN5BelE+ZYiM2RvOjp7/xYWYsmpHvRCz+5+x0sTnE8IqPYM0fAtGZjWNOtf0FT
QWqxFcGxHrqwwqP9PEUzFr5JquWjKNYJkFj7X3KZXiUZ2yyCMNxj6WFOraF7AyZovgpZy51GjfC8
cSJ6Q0srEYZpeF9nRhwIuUqd8NQoMCMQSnbC9vGIxB+3593zZPc1F0zgV/rkjKgd8DcCjCZpED9w
XDEk3CqY8MGD4tEB9rEeHK3FGX9jrksS8qyorGgvL2HLEVQxAIz3qBH+NpPIc26TaP7tu10kYcZz
gwH6nDWdntelTTG4im/5Np53yf+qAYr+bWnv20djRe7qv8EXkB+j8kBbDNik9OuUlhjjXOXyeVj4
mzyx2QaeTk/w6/ogZW8YpnodVGAQN/kxU2GOqOmPQ56wRfwpE85BX0DC0FRK8GLs3BFg+8Bbxuhy
YK/XWr0KR6/0vzxT+roCcewwTkDiaZrhMOuZRN2S3p4x1t/5sLy01B3+muYY3aII3xHMGfJ2XqLw
KeD7vWgC7Mw4dfau4MRMvgO+zAiala9guqwrWnuO6HctgPYqL6QXhnIjncKUsuDfR8h7qViWnPSS
EMOBjnEtX7r2/A6G7/h7M2w8FFtmluESgzcsaZYXVRAg4RTaHhBuPSY3ZSWnzKZrZgTU6ERaeQag
BVL1Eq/Msq4S4uj4/HsrsHG5j7VZfUgQ3JayqXpcwd4M4mvRg1WkXAwUAqCEI0SHdOc7MztpcMUk
GS06j4SP2ZdXMlt+pBzQkDeVkrJs4I+7F04aAowMiX4qcCm2alSzruI9OcaVFnLwb6BS842Bi39I
x8fMoVx5XTRXNZVt6+qQt9LO4nOiCseHEk/wKcC7QYiAbyD3030+GRNny6Hm3KgsmrzT4W2RcwL3
dEfHaYALY87qGP+xjvb6oOdAZzVQaH5phmYp9c0wfb6ibyEcEwm1pxVDN4OS6Sb3xlA47tb0MWcv
a0lzdeMthgNhD/lj5qzZuxzEa4ztylIuj2itKAxv7dgiLmGCOkAprhsjdMIXCz36Dr3hg9+CNIV8
LMZXRKwhZXTpOfN0KFn7iYMCOVzAJouzZvfk8cuy4XrUiEVa+P9puuYDsL1Aa7qke1+H8mD38Nvm
y/a/cNYBTQ9W9TrvlZwp1mMuhScONw1go1GpXgpmqsdXZI+CBL8IBfr5+bWBSHu+P/BeF/UQhGv5
3zO3f27O9ZKC58p2VmUA7OFucgBjTvvM3j1y8hUt3PVIVnx9DUGIHwmFdtUAgAFmfbQOfxS9fi1g
9OE2MWQ+bEd8YoLnS21zVCPrSfx/VhT0N/WrozbLb/wKYSqCaLiLuD/sibvr2OWe8ee5IEh/jZZq
fh7Soy3MQD6ec/swph4MHh//pgqanKumJV/bN8oyqLC0Gy+4jxr21bmKrs/64l18j1Z5heuXAbOE
gB3XsTPcyay4cLNFaeR6Av/yZNawfOnQH8cxq47X3Edj2lN5lKAKc6m2V/h+dhXA6v1AbwdTDZ9w
02zuIUhSnIKWkhNfisSa6LJ4WWE9lkNwDLKgfpZIqV11qAWYAX7OVAk90bRkFfhgk6i/NWvkp6wx
SvrpNcevxs7LOA==
`protect end_protected
