`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52720)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aPkk/LZprZljgyNzZTGF6gcxBz
LkEl/7f+3dcASD/i/Kgp6ausNehiRTVNSFJQttPYKRUEkcK5Nd4Tj3+AjM/7ZbSaaQxH26DuGqXU
K6Q/BVcH7ZjyLPnqXWa2DKOdNrDULiF9N+Ihqa7VD58WpbepjHecVsh1pRFAIkHl0vLTKmkDGr0w
QKP7oBk+q09yRRZH3d3T2lvAmM5N9TzRGyBLPK3U6NdesqfrhKKB3TjTjZZ+0R/EgGADHTQhRf7p
/LeWcZUbhF0sw6FgRgsWWX9EwVxAj5wKI1OF8U4LzFjjSMKXwAKCqiLWjFyTQyvq+jPU3yvdOe1p
OVDIkPF0VmSkmmJ9n7PdePOSRdCFKkvvAKgDi8koy/tqNQSu5BwXC7IBMjZ7pvMFZt0/kzccuT7G
7j4a2Zu8ZTgZ3gcyaBAXbSeLfQfQNRauWLomphpb3og3gZVcSuPweqqhX47u3HDuJoVOSfzakMlt
AOfdffBzkoLwYBNYTCe/FZWKZdoGCK2nizDXdLyp8nKxLQzuAayx0ysORRj6m8egxIAHdbZ1436W
TBTDpdtlH9MlXPiAjeYQ7u9uKLv8npc3QuSUMvm18ky2I8O22ctDWLc2Z9Ipqm7RsmUQQRgWNja0
jDdFEglDRkK4R1Pt/yIy9nmyA50qJPLL4kUjN7m6c/QgjGz1glTkmUJsvLEsLumO789RIMUVpae0
/5sE9ftiiJY8wsnaInFx0dJ3oauEg1khQGoxYMqF6UF9fktgRMZmmIazR48pREaLT2lGmCyK6L8h
TGq/WUgtEAxelVbPoq2ObLXDdVL8Yjy9VomuFN42ttaWO9ZeyDmolkLbzvw3ivqdxeIJs6fznHNp
4WmLSefeZrCVh/IWBVXfeeNK6ZMTiwMhbfAnAi3crNvZeMMbBoCesdFH2d46E/zpmUouV6fAn+qO
APJlBBdB/s8F+lNlGxOklyPjV9bMMXtWYs6Npy+SVluMVPd8jHpdMOUV0yNl4AjVvx9roKxS13SR
OmcRPRCX5rCIm46L4gKCAFPUoo8goS1BzET5xDG6dA0gLkMM0lsqr4/sFhJv1e6ZwBlHG7SyjNYp
lBplNMw01VvcY5BtDEaLomWv0SH8rcr6sTKEeT/ZAD26TFMc5WZ8MT3pnkwboBM9JY2CNWKudOdo
XM4qgR6/S487XL9C1En1EEhW2UN+M5jEWTSr0TXzXGpb7ayYsqrAWeTiKpH7Ul0B2ibXCfcn0hDc
UgRvghuh/cpjS/9/o6c0lEQ/swyVrIBG3mGYTM+mNITlPpKhzyAWUXhbkTfcXhb+HqzUCSd3u6LA
hB2vKX6lji7AVt7skJWU+ccjtve/Q8yxzJbd1Jn/uAQrH6GnEvI8zgdS79NVm+JaVxA8/kHhbe10
R3kgTK7WRRMc7iUIWNxXVyrVNVUE6S9SuuOIxl9qWljbv62nZGE3nBG8machpMpeYR/3UDZgzNqW
5X6OJhU3eLU+iHekvCOlD3GIBj1Zw4+dAi33PUQs+4h8DtYS1smB9HgFg0P70Mc2yPHURYy3SW8x
6zXgL/w4rsRMe5ZQtIxHRog++glCsSi0yMl9U002QwLzP46xv6JU3hpqqHRvBIW4RNsFOeikbi5c
WRYpz/lEi8ZjAKTzXk34+yu1jQbN17W6llluTbe+PqV0SZGpN/KgC4fP/I9TlXLpSElu0RqbcXzu
feTqOt36OrE9zk31Os8mhS5jsqYt90F6wYHDRPjGwlWZmdDy5YajNFbOkekvk491auttm+YMxQF8
7P3AjmqysvXrqvXIC2Qt+WB8J0eNJ2E8aiXpeweeQj3f07UO/VUUh6bx88sS2SYVwsT+F3UBEv9I
GuJ5O37Hw8F89jMYc3EszOq5xXMEBYECBza1PHqze5FkUfj5RH/SQ70weX2AUyS0fb4eWVP0d/BJ
96dD26j/Nlr11lK52Jxx4p4FpiODg0SlR6mZXRwVPqe/mAEsgaYeR6CWbV4H7Ihco8A43qYHtc9/
naL+F6nZBxpvANslb0rwaZliB47j78JTyAFNSU2Czkinzd61wRBDaMcaByoQalEY25o6IVQfBQnL
MwdgzDLl6PqDnJQfSWCJEC6JlFefjswUja0PxK183tW7n3iuOaq+tNM8ZLR3EyUiv4HHwURKaHl9
oR4rqqQak7SqRVu3MGubGyp4ShcfM3PBsUTj5i+HOoYK5P9uW3W1OAtzjLK3w3djJ05iynbleVDe
cAh5HZdz7RF7rqkZtLxAl1GCvplBQkGahT9hM0hWijCfqYB3dv7pLmi47ZM1zf/+4Rz+s5n2Xdmk
V0ITKnJN2zZ/jo4A1UQf+8EmPY7JNwPGHcGOco1aiIHGuivDlt7OVgLXUZ0BDYPi2zKin0i11ar9
q17fEF4GUdEnkPXTuxXbXrB338OsOvTg4IZ/x1aRS3xqcp96SmoycfmP3xmgbeOlazLmDo2mt6dY
9nP9LT7ocm7IpMMUiMJltKpDY5Ez3/Vk58OzHjtukXf9ppP6gkk0zVBopJVlCw2vRoHy7jJO4HVC
pdvPQucLMe4HeeahjdPNKIScZkMyieF2BeNKFXG8TRnX0in0qDWkUDhrhIMAL8M2KxaFOlBzYaSB
etJzWipnreDi/jOCay2/UrVidvHINtSH5zU8ZpHTfw0+w8oXNqutdwnJgRYJuh5vc0zUOv91bRCZ
inko1GPOCzhhNqHzVLqMnPMKJwsUnJ/HKjBLyNK6/yFzM6IMQTtje15cBQJ6POm0KbMKh9wp4TS4
ku+6Jj9vj19XOi2GX2TlFvoo930vjYot+/NvZoA57YPFZWGzVF4jUa9q248hD9s+7GZTbCl9Dih7
0ZCVIkm7KsB9VL9BnKBZNkw+qqqBZbgQGCiTt8J5n7IHIBuLEnKIihlrb4icqeTaQP81TMljAoZK
lYMg+UYmK5te/t33DoO0lB5YcV19IIvc1qysHx3Di0xED2/l74tjsUzz3r/HYyNsw8pgDMApwcYZ
DyNHlkJ3sYuBfkPCF/uHRAqdHVtWWsJzp1d+FPuo2oJYMpBVCw9GECcFZa/hDOxu76h+i7XNRGcK
emjA7Vo6DIohLLfrafC+UXZxlnyGVZAWjJalvGrxq8Tp6Vk5A5eUmEs+jNuzEpXe8xr5TqI2w2AS
rzVOlL5SfVMDjtQVqnHq6gQbZbLAxwRtE2uuWIooJ7kpaagIgH19sfKHvg8X4t3H1lzElE4OwO1f
P+jAUVcuz3fxbu6x2Mh/kwPr0U1J4sLfFBCtmEGsqk8vn4vNqdgGkU4Ne7IJsVaUR34wr/ZVM0qq
pXRvAH8ET+0sWXIna3yRlDsPONMgCkDxPVBL0yIO82baxL5WIO+aGU3jUpVSt10TDV4ACvnhsAjR
Ia9Ejoq2NJZLe8Lo9o1BQUyG4iTo4Nw6Hn0CIGgnGN5DsvWZdvj6qWI0U+H/QC1AV0oxKpKzH/US
yWqmJjVr4MhZtzrRC+If2tPuIhwsSy/czfbFhLh7EkNwokr9FWIX34ZOevkz0NdgR4yZIYwkGmPg
3fXvUguYOWsoRD+unoPsFrKeTa6im6SH6X91g9mjNWPG95PGQ7w0AQm0oRJgztWTrbuZhIqmPzOH
MjNq5LA9nTn6obey5iEql/uXTgFZ8IHbfd+NeCaqQ6O6HgbPgPoIt0MpzsEDx5g7/NQgzpcQaLpH
CwGLsjED0cgCwTWeDDuk8ARgbdgClnNQ7KjuJ0EY4PBbwIGvYH1NfHtQumfUWlMk3LjUkW87ght/
2jVJ4HUXLFud22ByJLxq3WoA0szuyaOziStON9ZmmETvzWZsxtnUxZeRFHtufiAj9sCKxQzGxOjq
XJfr+pzCFPpv+KCbanFPJqo4iE1zdd3BzbR7+qxJivjXw/ZuernOX5DjmeXQqUB6bwevpRCfFLlp
vv9zKpMWszhtsVXTf++k/gXlCzSbUK4zfPIuCi/dtbfszSVuSj3UgO/281Sz19HqKZ1HoXEAO98B
VrSkR9ZjP0A1LvGgPhCY6awXeVk1I2Em1IG3GwxjQdjRa+uXMbOueLZl45OwsYrIVq9WNvIALNUy
gsBXEKjqDHYdwl6qEGHIhrPfBAPWTtB0fk0AgC84kgw7pwiD/kskrhaIHQy+NB3cpGhFmy5Ehq0z
n3SxjzgGXu81ak1yzlY+uCiVcm4l3/zKwdZ1TYVyivF9GAZ2JXRWei4XhblQxYw9pApoTVy5Hl9l
WA5q1dXSaSRcW0xXIIhsTVQFQZXVJANb5C9m0fv0FNhVV9Zo2S9hQruNDFso1z7VCyxkJn5nqnBe
mXtP7BTr0q2ooOyKZ2ok9014KlzznoX/miFld7F4y+q537j6WyV1IIsx4Qx4Wm+NICubDqFDbR7L
jtFg9hmfRS6VTMb93nydkpIqyeB8GtgyPHzkRm9W7wnqpRIuFvRwG5FJa9j5A6LOL+eOVxQToBiJ
/7rMZ3gINqX2W/6P5rJBdLG1ySy/Eujcs6GEyUUh0/8m1Zk3y9l8Ua09BbciWF5qa191RCLoz8cc
ur0mdJWhcbfPJUq5Y8ukacql2+CRqOHv1d/Lk390ak/t6gq7VkNn0pceu7XyWPs6Glbs8R6WANDy
wIEaaMe5AnNVWPsupbfG9EXGiv1/yhR4bKsX3ejZKRQWCDU4xp+UUyxL9TjxhqnwHhmE0J/OeeJN
uCj0avPiO4Bh0s3Wh6ztZnz5n0twgcSkFr6/cZ/egUg4UzEdhgEV/I5deBRLDCzqFVsDupkJI44J
L1kuOL+f9bzXKPj7FAFqpDOU54RhWDPa2MqAx06gEWdQkHVbkyONW1NDn/gxUHpCPbgM7R3I92E6
B7i6qt2WuoN6V4YRtIBsbx9oZna95LgPB/R4Ll0e5eOtpx8uF8ENa560h1DmIy5OwnDNxn387Sw/
gZ+bdV+mND1Sw8iY7G8/xcSSZoxnsv1JUdKljJ7BPITolPuvTk7Tw7uSSNvmvm5cOuZx0HrHfohb
JEOHqCQ41cSm68YY1hO3arCT0/X7Y+2722KVYivktw4/2hHRPo9klW1ZghJaakMvRqeHEkEZBSkz
l/YLLzWnbNnWI645r2FRwoPcWcPerrdcOKwy3drH4LlzpxfM4NH3SirI7I1WqFWZMhnlOY4MFLJ2
/b5B4qtVhZ2lvfsreeXliAl/x5bAVttpLYV9zl6VHEzn0TsUXc4Q0H9EGwzuiDfzTo7jwt4guX4b
YGbn1t7a+kcGHex/VErG6nun+ph4Nwh/xC/HRqqOrmcaSyVptOGiZF6AaHuN0KRJlDv/dEgDJ6op
e1r5DhmVtzfkblBM2TmvCgjb2rD5jc+FmbNbY1r9XFYhyyNOvOXndgYmjLksaT/MK2UxRROAumln
ZrINQjBycOI9sHdv6Psv3pPR2/eNGrYHHtF7ZOi5F9SPcqGLUax3Gwf/KIcjVgsZFn/lJCCMGbMH
hEbBF/atNJolU3fuUg7jjnp9pOPHPOQsotNzSn2J2AS5KP70jf7MpQmObNeZ4m6kzkmE3AazEshW
UdomFDYnbduML4+pBga+dgrHfF2M2hqmm7pSXuPdsIOrkIYp+4xDxgvYA/hterpWVikil5gEUpTL
VXZzHAyKTInq7RoMggN93Jii0Mi8gFpIVEQspo5hLm4RdHyVRzJu2Uzgg31sbzW5IaJ1NirlZmzh
pyYQ5LPyzEeh8TCc6qbfTsFLnB1ciWAPEk4GCWUfjIk1fyAh/hIyeOrkUohFi22Ys3fitU3Khn+4
7/YZnvP81JpXgHOGTYz+19x3lahQpmATexNLhpxv53dizju9AYwjL9xc1dnJlqghNoqXSQiyWh6Z
wp0IO9ZHuj+aW1lGx6wlT0C4BRd8DWDZ/R7w6ikgQgZQL3lkg/YzlzFe+RcA2K3fTZvysPKZhiHX
glD8Tv3gEX7wXyCzLgU/L8Yz3itBXPL5bLCzsRtNXTUIsdGYmomHqNwM4fmp1qij/BGSki98eCOy
wfFQpjsNu4AkruPQYMPH8JjzUwWJZlb+TFHhaEDWoFmpMBlKWYAjJ9Sduf3WOV0VAirVV9y7JIqO
IX7JvGg81FpKIwv3OTQpUNyiZXoe1SOhocrZQVRiXat3t2hlOdslHaCtUXKCdzDTcCOE6BxTcLs6
irHCyNfOxaSNA0jWu9boaJT8Kpml235pkjQBdQhmErHwNE7T1V+a14zk7YTNWYbDfwQP4Ya4FpmD
uJD07+Pi8ek+mVh4ZqB4hkW8/yVul75iP5usVYXXn2KXQ928mUlE/ExsIzZQX73Uz+HMCjPVeKiU
ZpY/BmbxA2X58V0LTc7q0C/9BEAna0DxNj/3gwmMnpyzHMF6PrVX7Bthhy5Tm1xmBPzld9MicQa9
6buu1QPh58epbyQzn15e2ky9Fe7FPmHN4b56wlfRsOMnDBDV0+JANXdakb30bDT2aXdUpxNIXpki
AthfL4mm3kk3/dGDitXOg6LzhX+d3G2aVyzsQuxXW/Z4zJldh3Yqj7GwcfvTqgiaa1DLtUlnnkp2
nzZX8axYVCldZC2saCgq3yr3axC0meFiJU9rFBUFbZVnuclyym20hhj0KMHjeSSgOgShJeyLtb+L
KCXsE5SlQnH7d/nosD0MDvt/65mDzdakMikumAU+I9Oi1grZQFklseepcCF+baNcjmllXQ6p7pnS
QfWqE408R+x9KSlueGl8+NBXW70Uo5qJlHVma6REfRhxFe7thWmBDLDQx9F8HgWgsj5r3g0vJ3kX
L5zR9+mVU9468gWzsPLiwhddZEGSDbXm81KcDryX7WnuXiJzz1JduBK91Ea7FYOBb9CkwbJuzfka
fickrPNKQ+bjrljd6zgBb5ldBxSKJWyHmNXF6tnGmHamY464Xtm5+Soj62cXIRPY19eeACWxR5gF
MajBYffynDjM+twdhDYiE+suXae6z7RYlpSG+DyS+/P28vg20wW2lcVwvsVl7TMkxKj+Jy8jojRn
CGSTx+nfkEW/34XVabFJDwEFmYolKB5Q+G9uqJz4cY4sb4JGN/75AIA0USxY6HKsGjGQQrnDwIo2
hvVW+1ICWFnykaYdw1iUz8kb+1SPaoiBW+NYjhQ2qOnKNKR4X54sEZirLcsRHd7PDjjcjPcmAxlq
dJFgcrbCSSDjIByNIoCJRhJ8NHT4yKQ4ENK0iVKwowPQdxSzBd1HIhRJrlnN6+o5UsMVyF1zHnMF
vmgWeT7sotnXuPIw/jOGQw+LZ+6uYJDpISJ5LmroevtUgXsu/HaTJG8Le45PbQ20Z+rsXj05bPyi
2qTKXKRf8ftb0n6jLAkQ0QGx+zPhuqEXL/nMFia5LexOMSJflJIR8OwVVtHbolB4pd8rzsGRq4Ef
O6IjDn64JRsBps1q+aHCMcOnzvWSkZHYhlc0eUP67G0M2f9SdqYvu23LmyxebOAA2+LmQX5Luwc7
HSC2kbrnLelqyE/tcDTAc5nXjh78k8P2Xs7Pto90Mqsmz95qJbUnVuTdzxs+lGDXrZHmSa7BGFKs
zmMgFyAHe3AgsKSboW7MqH79eo2RoEcPtCetA/3/+Z7oVaw16j0yfcwHbQOWauFIa6un26q0JRw3
Z0b8d6FqGGe/dmLv0LTKTsYcULsDHADWWpr1+fjB6nkmD8R445+0PTCzqVjvOazAZVkau/MtgTMK
MWh1fU0tXPzKt4mLhZWNrd0H+Wb6IiQSEyFbfsdbQo0QLWvnmRdLUp2bBIuXhD5tAciX4my51qgF
qbKtkR8f4e+dRex+RVO8ytdfI+u06hJGniCGe2LY7d2Pmd9LG5oZbA58d0NL3CQNag/3/bMdLw7f
MIjaKnJ7OqT+J2re2DlzkekpCaJ59ruTfcR5dzfU6SQrU3KOtwjtCa8zoK4JRzDHyKYWD4oBZH/l
joTAVS9TZRbwQVYLfZcpb6WB7d10lBX5HguXZgsLk9VT13JmX0UP33RJ+uMXvd196HnR/LUVY3vo
/HUNeqIVEswQjcY8LEEmcjO9gRDv2GuxHHonk35RyEBsXm4sTQoN1DD4ayVSBmkYJYi/4D3dov1B
bG9mqcmKJbXJRaTcck0O+9QQVAtliQ3HjCpg9tYCvvWZ4ExCG3titEnsM8G13oggvZ3WshHUTnsk
2PqYNOjqOuFx1+bokKwyacHEiZAYR1FNp2TlzeOq3x7mT6XCXITHkMEhAygn5KcDUwvLeK7oOa3V
oV69ChoMmATJi3DZw5NKjjQ3ShsE5pyW3ngBeHUyJTGCqBbMUijL580jsdo2XBMnRwgiqnRX6fIy
gzqtGXTgX4Boh566biDJ82X5HEULyHFJW7srTrXUmpNJaiXE4VojKx/yctCXRvppUW7b5NJq1G0f
inPQ6LxIcMkBwzpzlMPSShCkhPzQeyGoQ2zFSkb4yqiKtNFiloZWoo+I3SZWvm1iz3oAn5uFUoMF
Cq90bbR8+YBmVTknyQ2cNxh0rFdrEKC5RiwlLUctwm/RNSfdpYAd1A4u0LPQ/HD4572VJIwDFt65
t9vO2btZTPiSFcYoaFN0JueHrlEJgbp+m5nUZTyh5rXXowjcP3kL3r1QfqpVOEENOJ4/OgmTCaFX
C/5+5g6NgxKKumqVbCUk8ka1ogViQqentArO5Du2A1T3ZmrNFHV79T7K71eawA+0X1ridlmk1MFa
OrMJ3Pr+psmevmY/pCT9FQpi35h6FxX7uJG2b5U1Lgbyvi/nnvS/96p0eDEfh/rNHMRaCWYJFjTz
f499LXhk3lrT0jaf58EkkmC6hCWNHpMzQYUMTWnyYfz/DpYImc3KlLPxqWwdUWlDHF9X0AVqYGdZ
c8qyk3OhHb70eFOa47bhQvPpGfLOEfcMnN8ltRNtbWi+nFlatBsC6pVmzgFshReKPMVepR/NePE7
LZkMNRyA6JGHnMBKc9nfkWVJTeC5XdwpaEC7VcMtsWnIMMkhQ8MoFCtpFBr2dZeUeZrWDIjxmhPT
/tMBwJNYf1rJjuaVl7eQqX9MM11GuXtLn53tlHukgaShiyeM6e4Iz536Rm+c/8rQuu5BhetTmQoI
NrBnCR9wz4zxdGDPnXmu+ToYUPBSj9GASd5bWK7mfXvk2jnLYKUIjYZ76AfFrRt4WCa6oKn292Pl
68Xgy6JgmIGLEnnqsGwpxWCkmhmWnjdSbM4ZyIgU1wr1FeeKPq6F6rse680BG0yp2yyy+hYtzzVg
Qm5ZAIiQpIzteo1pGlPRKW0BAOVikWaS83IpiFftpWHs+doKSJvPX4+4psHRKzpubYxfgs0cxF89
CTY6r7KgrA5rbZkClwtHg64nFkNb8aSy0aw6KVwN6wJwNukAiLx0MmG6wqITwkfR3rBDTvYcbKgL
QObmmXj7euXpUaGUX0EFkMNk5mZHedrcTuJUb+XbyVqXJgG2UzibDqjsphtdacxC3DaxMr548W+a
dVuDziTYdcvwEdUplFqtoroYj1kb4VMfgViP8nmhRRnx81qF00B8zjdIEcpb7oDp5wus8xQtaR+H
Y31DLfzknWmynHNNaCeuuF8ApUVDZFN/1ffjHacmTlNKTdzY2xE99zFWFpUKEaKMx7PAcOuh570d
nE+FRFFjdYQFZBF9/7Gat58qF5DGActeIYXIWYb4+vKDNLHlj1n45UBMSHWE4YiGCf4pkTM8OiEP
+EPAk7xdMpzwdM+7PAFsfJJ0lyHkqJT4ZnEnGhkFy6osH6bVFejvGaH3vzhhYlvTabCsATYy5xlX
0hsSKzxO3qI7yHc4gYU76OHQtah8s8Bqhh2lubNMpYPpH71EULBa40Q7szNtPIbT+efDjpbm7ceJ
0TJyJKQXE43VQrZI1NIdiMOGIAD8qjIKdtRv8aGQ9AbOorWoCm3IzFLQWqfF3ON6ywNzUEr8zmZ8
JZPhdnvXyyldHDGh/WuZAZKX9a3NKnFcFVgN2qjLy8+52gwP7VeCj5SEFtUyzqfJ4ViS06I3JGpq
pxoF4IqFxB9BILa5eIlwTw499FP2IeD/cdGD4QIiWxciM7sxPrlZxCjRir2vBVffFR/Gox/oSnpt
Cth0nNDMWmHa6v4Rf5AfjeQuT71rxv4tCD03BctUBh0zLD1W/m+PV/bv16VX6x84a6yX6Ss7SzU3
3kMUn4NAJ4e3k+NtLkI4hFGWTR0pVA9Y/SwNZRarBeIx/Zf38gzI9wEfCZ1DebR5oakgApGuTzJA
XbShphpxR4ksCU2chy8e1Y1xvYtHP5hdkrxIkJ12Z8ZmgUYggG1+2Ai+3RhEyfrF/HK0AdLpUENA
FvcglwLizCMZimqq1H61wQzaXhHoMPlzMfLfT/DY+sgQK+8p8fxTGR61jcLUI4+1gFaNxUWYoQpW
luuxVqZ4Cd4+KjtynnC6iD5QQdhFVbHoau6E/n9ARFewoU9X1tWZGSGjhz1xgGgmW/XCZl4LRhQV
XSlLySuKCORvT5oaf7b6Qd9O0Cy9nm7ER+FngqlD71fPM9peNT6PN4kA0PZL8Ox1jAoNJjPeBvV6
g/xbmEjEsKJkKJ/WPb1KSu3Y/bxcmPIDjJzq5Q7qb/5OYAZWBct6ilA9fb1fBLmP16a4+euNj1ST
tvnRku0EBuHe1UKPdurKob3P8/RhjhRDsIBsmFfSJ7bLapAtvHGw6beT+mPiEaW+GM7wRfAG20zy
xh1aUIokR4+ud5nvrDuhuo0mJKPt2Ker+somEDsUvYu7VFnzoRHoo87y+ISi/ZiwQ7VOD2Mn9pfs
o/QSlRoZGgeEjxzKb/rHDtRfgBUqS6PZyDJxT0fPUKPGQnlJJijtDQIcfP34TjZxdPqpT6b1GC1b
+tInoVSCz/NlMU0wscJUW6Iwcj0gLN+l/Txe3MhtT5X4QBSTywBNiu/FFiMX0bwSlF56uTa/MBmz
hjpBDGsEyYVQgAsKaRKTIcD30IBTIeDru+msQ/I6h+X9WK0RFSX2GXXbYpr7Zboy4AULw9tvg3sl
3452dDWDsw5HNIjLHuHtSzWPRRzrItdIwwCgc9QJJ3By5sdDBkOcOUe3th64WC7Edj9cVUphRl8y
2mwL7fCmqGDVoChMEK72x2TQCihtoUu3m+iju/Q/3TtZ4XG8HIp4x7sDyA/IRw7apq63oytRAya2
cS90uj/0I4av9+aBQzspoTIdEagRcYzu67PjumjVH4HB6EeriBklG7xkWmLPwmwxSK+39/P1p6nv
dW8XMxAbuX3Y0lxYvb3kQys+0w6ESXuGWzdvzIVnNJYVT3e3O4vOv701SoWOB9pI2zxQeFGwefmA
lbJnyVMOHIZql0ZiWh/l723Ozv2R0TjRF95GIQm+9D8LFh6bYMrdGH0iPONZwDTGhYQJ+BkoW3ps
lg6z8XiBj16Aiw40teoEl1qDTCH4BLr3Y/n7eSE/7GiMivZW5g9MC7PrSBHp4r5FJVHJy/53VpZk
thznhUbwuweSoVpUP4EwthNfmb3SjXXC5Pe9LRwP1a7icPcuhPsZNRHdXTqDg14E+JwbjosLhhzO
QR3wNWrmP+J23dT6rKEkXViK8x+i7dLSHeySN4/mjcsR2pLrj75Oenq/bulIZbSEZh6sV0LYmZ0f
/JrdkqgSNLb4SY9gP+KWZJPKHbQ/I8YJ33M0Z7+lZTG3OL77tpJVW5+WcpJHWTicCtRo2IA4fzaj
UH7ByTCb4SA5rxVLTxdM9fY3b1719l53OXwFpFIymOlC/0fDeBDfIZgxwLPlkvt3Asv7+zeTqkXb
OqIe3y7eK96h7Xh/99/HFpQDnJspKBGTQCtqSZ5N7ik1z1Cnsg7+Nk2T+ZggaXQL9hlAerBFCiT4
5PQulGy+gyd3879ZSfN1RwWz1ZmC1S7YbEtXu1uCxsxNSuWyr/4jvk0dBuqNCGtSPANqj4CNrd8k
VsM45ITJbWV7QaGiF/x3gP5YR75PR/afbQgKULMvbRQyQJePT7bHeqop/JMd1IELRT7xtuD/9EzU
dUsFCap0cK6RVux9bGpD+GgfZFAApUIBEbJ4kZzbk04IYlhhwn1O3GVTQornqDNEr4Y5N6x1GrL9
Ln8rOZawxRhpXB2ZnLLLZtBftuLCf23SodtiHlZPiGJ+PMWk6Tj9L+BNXHjKANBK1ufGUbxPSueb
BG39bsfpHjmxuGVpST+IJNR5lJ2ont4/t7SS407ADEnS2y1LB3vB/SQu0AIxar3P1XRrr9TDFKQo
kqdnZPJ5gRpTpb3CEJFNy/tt2jq+DgZJQD3/EYjellPjsIFJwagGUiws6GaK7z8zbgMQX8UPMxtS
EGZUQ1fD7ktlVTtiPOVe22Gax2tx6PAlesLVGM89Y2CtWt8uZXlQdhmFZZ+Pse8be8sWjHRO2Y/B
84pb/MgcFnCCbtqYKfEVpjAJg63PWkkIa2xeaapUxJg5pjRxMrYMcLs3P9tda07PEg+G9ev7VEWi
iYzr97xalc0dqyAwDJ96p2S0QLdehBUSPtL13cdgED87rd7kZ67eWXcVa8CCIcg9Rwr4Ip9u354e
/zoUPa+xTCWhcnU3xR4R2XUDgk7kG7uZviWxM9I0DUw/wmH1ME+Suh28S4KQMSkPOoLLcVvrfr73
CeV1CgYd3l6gvWcsExpOUEXLxwOg2ujj5WO76cj13jOptXXkw4Fad+3g1bymwAg7TSvrM+11jIcm
gKvHtfQpdrhk9Xwcp0aFKIxQTZm67pHCK0QJ/EhUCW+jAtPrP53MGjGaoYCugz4HA0UkgUfI0MGo
FLtStmKIVHymS0nSlmk5UB4cVnOCDsUt6pYfe8aMWNnzRxcz+r7ZueIGnnCuiNPn2uAXTymBQWv0
zsNqk3huKbnN6VqgoMTmjHoeckjmE8srau+krMoHQOSO0DZdn2Unht7P5xKEggRkz4WIFISIz/qK
I9oIBAibPIaXDfB/CGE7mJEyGYtMkD2aA/HULDfA5xJ6YVC019saUANO1LMDrBXxE0qGSA7SY82Z
ApspcQahaRKdoln7ly2gRv7Y8JXaqyBoTA7ZpbbPtaZTABUXp99qYfpafm0mYwYVoUV+3sdlRKFV
Q4kr3z3bvR8eEk5qo2dloxy6NjL0RnMnO94jzUeDLckTWr4E5NlhA1Axyxex2PFcGHA1ua3hFhNc
06u8a4Gtea3hirT/5CEewQc8PMedAJZJL8g7ozmlvGu+1N+fQH1WBEwl32zaDini+kvWRDLpooXM
iyzUYigbzKVQmaQvAYmXOj2eh25RjYmvB/f/N3GzpDnIbKOws2cI6nYbdKh3WCHwxgIFOCTDvSBy
D16qMNzz1RnDq8LARGC5HLuIxvJyJnRjs5fkLj9r4de+n/fL2EsZLWZN8IMwRGe/B0/oQW/A7fpR
vaxmtFL+IqDzoOgSaDDzYi+LC1i3GD0IxOgbGrttR0t7Xsul0lRhL3OB7Y0hr8gYq57n9JsMDoLb
lB+3MnDNKFQ0BBfU43ttcFY/YW5GKfEjypwOaTW5K4ADAwH3VqetWvMWRASuzCZFjzq5H39QCkfy
GEsd6Mv8IhTpLBGvgbRkwSXxfJUjweR7YsWxJ+p7NDCApRwm+pa3ELKxsDAsSkFBoTlcZw3IiQe+
roV8KjyUOspgYjNXJ19GHtMwBXc/GCjgzRFFwTGT1/nRDGmrfnlOvYBoV44AncpeLHSAGxbxMLfL
zbDdiEVflXnPW97hPYlSCd5SpmF/Ez+ee8/pU1aOIfqzAwut6fLSjz75ItKBaB9W1YnY8tIIiTKo
h1VzdcJuwd0Wc1pgfljvaGxkSonNIOFaNvnPiSEL8PEsVAJAZ5p68992tKLjbcUT3yKXTKvVO8Zd
Iwop9qi9bx9aoZXL4eq/S+j5GaCzCeJC3aVJQIUouzJwSrsiiHQ/O9ZJsWDvDZZV5n4iV9H459dt
7gvLEM4H29Q38KQbxLGv4iDvzIHeCT5IR4KeFJ7BxajVYeHJqYv7HHFYGZcpWKyIuIXh5hbYmBDu
UIuMGmsbOmdl45E3X37c3TpzPiGHdDnsyUc698UP0yXNOckiE6QhZeSMVmf/X0WmsG1iaQ1yPWYG
IUIgcd67mz68hpQr4PIkejETvyj93mxr0f5wX8KaYox2mlD5UO9jgOYjFnXNb8ZD3PbqoONneMLT
OZf4T/C+dJM9h5PMBPGZVskzpWWvmoI9hlo8qhImcTHNqI10s6u4bav6LrVVkLagCGkVmcFN/ZZz
2wu9iNeans2tAkwsL3czb4stRNG3GJAvncw6M1L4RW9W5E3Tz04ShLrWapSCZw64tS8g2kC5mMQY
MxHUN+TH/OPgVQiflP3GWVvnMMY7dKVP9VpZB/xQB53KXtodqqMwEu/6xv/e9yw66bMVjsbzEJCw
GiIr8OtvyL4g9u+fb2X3KuD8uzxhsFGa+pGah9rbnPN50axFVd6/h+mqiqqD2t1BtTsRTlsO6hSl
CFAV2IOK4++4dIg76qtTLfwiQeF2rg+Jr2G981/pRDHXS4CsxNVhMV0EvboHiVxtLOcF22vglwi1
9PmuuBSufcAa2HWPYwhE+MRE0AVFqKbgzFVw1ZIKaT7NDvz8qXnaVZfrs3/9Pa3Fjpgcb0Bc+omA
KaHp0ukONa/5Z+Wwx3Q6gBCNh2XmKyIddQICZfrSwHZ6H52tW56LxF38dCveiSuuly2Y1rCzYjcj
QB8EPIVZJwyb7fkHdXfD9h9eYo8nBrB8TGt9H9B0pocrj1ZN7t7AjyFosgsn0hVi6V+t/dD5SWG6
fLpTEZeT5bZkQsSWYbQDttoGXrceiNn+bhIUklOUG9w1rAQFw2K/SSHO3/63w5UWlzklJs+JjxXZ
3DPM8oP12iJR9D+ze2E6OAuvsQJvn4RdcKx3WRlMN3+KXQm5SgqTRM+j8M4DM7pxLe1nCY5Eqn2O
sN8//9PolY3ZvuSqEcvVkyFwfsPm/HyH17RNaPtq2kLWtq5pdROtzQVnaunDw/kTmMKzNfyaMB1r
E00i+TlM3tWnjAxcw5HU2uxwkUm5D9UzUhDydXYH82xtIQeCqgQVIpkpDQnYbj8Y/MyWDon14P1R
QoojFMEj7hsPnRMIEyVzXULUpVFDbh1KwSFcoUlamg+Af+SPXFDGiNBYFxcgTuqQ1KDO5voizg7m
esxT9crvzaSNoq7mKSk8uto+Mzv8YKmqx8mOPqB4MbFPUQSq1VP97HoOvo0zc5mzV8oPg3v8xrAL
rEFn3Ns20evzGWcIQBlKCs+2psR1d/rEZK4pTL3yxHWHemyH0cWq5xircGobUe+wcwmmXF5b+DHx
4ONWtlCEtNIbgXszJ01hyHZVXGWNY68fGPekOUY/puiHHJrKgFPLXgw6t+fc6TSEAYB3QIrUeB0k
IJ2mkxclcjyrANHKIDs7+/bMkrPONoBr/6MoZhzdDwDqqxvzQolVQ+Y80yjdgGsV8thnPnNjc0xX
wnEQj3qIR8QxVNKviZg1UsKaB8VyZ0JFYEBQezGYE3dUvZrWMLb5L9cqzwREu+uVzun9RkPGsqr2
Fzv5lY0P73PpzyhuYwMX2oZBSS+sn1+WboHbmF6ShjS9EApGWDTrYl1x4PqOyU9cEMzvWWiNyWHz
RATQf494l+LN6Cvv09J/yTcM9oYhamfhn0GU0+OQgBL6F0z8p78DIeKcKdVNxcgqQSBC89cKxIPr
l4oMd26YaT2b7aX3xj8EAIwDybKDs/V+LBcVJeFZbHtttifqOGEDe2kU/4wAuoiL5CJ+h/sSKDQy
B26l5LHC/N8j0QUdIEQZw3Z9EEUH2r0R0NmDWS66mDfXXgPLBOLovgjKxTuq5aF9TqIMVtecDKHy
8lKjuxUsu3dL6dYZAmC9wmZNIroaWe1Ee2b9WCzQk2sK3jtbDlQXoLpuPRkXS0y9rmvY2p41bOwR
SITEXfQPJLeYoG9XCWZER2TD+FHyt1wtLrND5ZpdwykFYUssMrV79qOapFTs4U8+77APkQfazUw5
CbvC/RHi1Jw5Jie8EjP5INBkuBT1gezfUW4bCwu08W659AvjtI/njvJzTRMeuQCdf5+lUexx35jP
FnllaJ2OmqRx/ciGg+Kt4bAxEMSCGiCbYS/5gqx6zxmxjMM4YH90/VpvrkeXAUQaCkLQCs2yJ24W
5zpGwhWCXMvHOpAaW8SP78wshb8sS4cS6MGVwUNUMQse4NJrwGimjIunV6hCsqtaPVDJahEghijD
yrV9aypepQFPJNvkiVi4Lof6US5NRteBDDqTdhNIoYZ/ICe1owzqgKpNtjNC9UxigWBQWu75eYun
vfA5rImwzMEest04GOoSogg2EpTs1HLBpC+y/5BQ/IschNHapmUJAQ/wwp8equBZBFWXB6G9WszE
09sdy8bwqBgsSjf+vL7zzQ7tSoNhOfTPmxOpK8vpPJhZ2RryEUjLe13L8D8NlTzcs6X70qeoqzuF
6ZeFOxEDEB1AOVJypIDngPBRjQBI3beNnuljFnT1hKiLhGIz03RPzRUx+rNM92my5L+paG9QqjKH
N5GU6VTijhZ/43rWuEbGMulbKgLCN6HOSVuI5CtNFXo3lWjla6uyndD5W/CWmLWHPu/fFyiHH7qm
YRpR0rTW9GTIO8O0Aavc+EiYi5htnWM9vtrnsmtT9G5VAuIkQQ6nG6NxW8cHBOk5O2U9BuvGfhiX
B9ls5loPHVDI4pswjVyzz4J3N8Od7S9aQEUTZHHT/C0tlqyTYqeyjnGbgWc2fG/DEzy4+xXfUPx4
Q5PH8iJCqN7UTGPbkoyw7xmEXYs9lKsBqgHirc+sl20j1cKIuRI9ojn9MZUyk6zukG3K6sZMEnlH
3z+PyJPs9fsEeaY1YIZ0GHTSYZMrRZRcLmsFkpNzhyLufBuO0EPQfQtrp7S1ru/DOFMWR/f5ERK+
tccSn9pur2b6LNo1wGFk3MS5naHNUquxFOjXmlw7/jIKzLDtPRu1jhr7V85nephlflvKDxuXIVnH
bD96YZ4whhDFF7ClbpyCQx7e4bDFozt/wsWHcGhBSFRZVkyTfGO1i97k71iVqwe4elD5DwoEM9KI
4XtaIusRk1ScAVckaecHjAhtJ8yyLQ7b3OZooB12U4aFBnZPSdpgYLL/bC6KnBvmQNSxq/IyB4k3
qy23KJpskpP5ErPG9wkTyOjtaIUP5i83rwTu5ADgGyafrE5H0ejicqh/jF58UWzZqqRcEEsM3yNA
AGF3pCCW0IFCmFurBWZ2hbuXZBSEa2JZ8kFYQStK5NWlNIi+NtHwdF5wYHHlt4sqzQ2Hbr3JA9Eu
RpTGR/F5MG5FA5mDP804+CklMaeFiphsrhaAOvT8FS4+zk5SSgZAGx/iGsSFqdCaK4YGc05CDJJn
3LSfCjQRrDZE+LlBcSgphbUe/2rlZGl50SuvfpokafMhuATJconocys2MRsHcUHeTqZPHUdMZQ2h
qkRcWuYbX8xxe5Rr/JybxMx+f7RUU9f8HS9/1NnaRQWYpGsYdan4T/4T0XS/lJh48tTGsUCic3KN
FaosBkvIghqu0FPyadOqEQGLy4v1KVdm/gtymCiOxrPLCJa0tAbbDgvzmrRDDFMVw4IKisnsBaBi
VY6oHUEMo9z1QVRjcuvsZPuk7srt/6lYbXdAc2cDl9G8seERi/wkDziujYKHspHC+X//xBPejGaz
aAvANOeT++FM9EMW3u8z6BSLtglpqCH0ws0dlKPavWznHr7uQtg+sSe5hzGn2dqFLBszxdByCGLs
G+oeeSSmg6fJ7o6OKedb7vsjieCVwONNudAbhbGa1YOMxS1l0uoaQ7vVukP448Dp8Mmmwzt46NdV
TMoPIV/VDQVVxF/GIk5yXFKljchSuQVfsSMMJ5WaxU4sJctbKze88CmfwJ6IpRu4DOWe5MYRomlW
9MLkBcaYqhdLQwSN2SXmKKzdp1fzZabXSbxpfZJ24lPK2y7qEw9VvSLHSCFOHO2xpvp6MfTb64HP
tf79OL90IPmMeldxh2QIv3qregzbB7FcKFjyllwFPjo/0aW84ifQ4rZlv/q91SxjDsIlhxLg3fLg
Z+9TyS+8v7q9nXaDES2vm5jY8AsizZ5HNqjtepDqKJ8K0I1bewk/GduM4u5gnVCEjG8Ds2xKRdqn
zSxmwWlK/6bhGJnWDzdNYkWPwsQKj4lKQpaARgqen+v+lBN6wb7MLeG28pgZox4HO2w7Eng0ChZe
45bRjgs/IHHYuKnofFrp3UaoTerF64kGUgIoN9tjxVqkb8lXtv+MKOlG3HP3WJiZWEiqJLQ2AlaT
a1qyh971PEd1Q/AiE3w/jEQWoWo24ZehLQ+3RYifQexWImRtUfKyQU4jNM3q8Hk1CPULGxBRHPty
RISre7F2ghhTX8gIwKSPGe82SpYd8IkqBrOAuVPiwP0npaNEpbBDTdP5tYw+CHr4IkTCG5ZUmPRa
lQEliI4lEXVFZPj6Zjnh5OnAw5DUxKcYjhD8Ku2rGT+6hjm1t9eHFOcJXzLjuZoU8KmySISTngKp
Aje3idNLVp328mAqtUhdGK45/Jd2YoUEu6oQyHLCz8meGBYsTQjU+KkfYTT/oQBLcWGpOlTBHEKh
eiC2FbwQGns0REAURnhXKMKxiVd2VDNxcy1MLIbgOW7gwt4hYyJFL9JB/LZKZtVhY+4FdJ1Q94gb
roTdYnltsErdJv6+W/76U9LjOSuSKnYlILCBKFUcSFwnnsObx9ExpX1pmcVEPsixVdyYBz/UoTgj
IxNEMUvBOmcTTpeZAeNbU9P3mTRNE/ha0VmA4M2oehrcY4yUJqIqHTxtoBSKcODveGfKnJQPHW2x
pOZ59klFCjDER/4DJNcmYl93rwU8656Sn4vOLuvT5CoO/zDUkga6rYIcm2R5wN3NcEQvqQteHlBm
gTXRiSkyH0tIVd8/HW0jLCkxCQAnW9jt1NmW5L7hjf6fdcYvxeyWLLvWs3Z3DdbNe/xdRXMO5GRJ
aG7smF/1Kr2d2gpRFunMoto4FQJ01mdVyEKPpt/ZBd0SLugeM/DLiAqSKWNSVOknDtF9j2+5fsCl
6ZYx/H1K6LG2lml48ZZpFkQk5DNLFEJyk2MgYGcMqtdbU1FsopJKssNWYavA1bf7Z34KK74dNFgk
3po45F+B7QJnL2txbU25+yKgZdGW/Eb+lGnbSrdLGyahNNgZNzzdlgBCVOoubUVOhMrLQt3cGhM+
wSgTNPEXJem/U5x7ri3wmrfJXg7NE8UW1YisPymhSzNPzbvb/yF9pbEA9wx1WGRnKRSTFx0rTsuy
mccrpK1lGYRf5GRkyqPz0NCNu3Z9yAMKbYo/LK071DEI947/ju7zj+RLZSpZUdsjmDJ/qufa+5g9
kAIjfuJPvNOXHvLCJtY7p8+e7NRCkjRHR3akGxAFg9JsUp+f2Wv5fNzgIvx8zkzIPkUx9NVkUlvM
atPqjuYW92lN/mNwRZNFOGOQCGymY74X6TnxXhm0viL3pvrNh92icd3+dKGd0aGxPTOh25th2UwG
ReZ/9cFwedFyvFQzSGpU5Sa5oVFYWgSgrATS3Z2MsAXKa1fwpe8f4hNUIFWvkZac4eQ/dVcsvycs
YNDGt24HmmCKLJxMRS+pF8SrXGJihza58P0W0HPvl3WKByjmUjaiH39anAN30SOz66whF6hMx24g
iBc/o5MB+67VK+qiuiIu84FBd5v0Y8QF0wafCyziEeXHrMLuiVtVFzBrpwng0O5v0GLPnSxwDNge
e9Gooe/qYgk7+NLJ4qnXm13iPgqLLinK8+2aJ82TRpa+0ICaAzGL2aqckpcUOwdF97Zq6g2ltvYa
R4pynAWLJgkChiyyFMLVTqFRzfoYtClSiMDD8BFKrHtkYL6RZCkLrWhUUfmHB7TvJMGkEyE8SwRD
s63KeKD9wwS3wIdU6XjUL/WB2CI/9/Mn0Hjy6GSfVfY/WbYITYry3fozvz9g/OKxzEi1kCuBWsAQ
T3XFyZrPN7mNnYW8WUvyiy2GTKmVlNuYo02IVEAIrP7ORl7V92uI7JUk+YR7SVyOvoGxNDBnOC9d
QdL+FjTRx6uNeymXLh985MN4h8UQZGvLfQ8TU6PdAbRHDegrUH7T7ui66WMmdFnosX/YhbG/+Acq
CALcb+e0nwKNZDp+PxAWBkA05qSP+1luwz6ADLD7XBY9ztqDeAsBIr5qVuDn+jqMVhQPh51AIFoq
pMBvA0e72xpSN37wcadoNxpdMi06cs0NkwCWepsblfGrJdDURmflrNYaQMAYT0v4NZupFCjSV/x4
KEdGXTYBeMLgNwA7HEcYdSxvJaKi3kWqtnO2oQ1968IMfOpmaz9FZuu0PQbNHi3iz+XnPT+qNDQ8
oX9bzs3543J877TDro52+QQOgNXQGqGEpj625qYHDGbrjGmYnhtWrhVt4hEbUfqXj8kLCZocgzEZ
TQHvMQz4t2uK1PGmZrCjWABqEKZ34vbkxnAWx3un7Y0E5HravSwzmhi4GDA3skD6NlLAwUhF2Fjw
MGuYiZ3ROK4b3oPXJqSA2I9zDsyvGHzEMzMDnQgCD3DM2XstgZZQe8ib4Pg/cGi5ub14QcQMfhiz
P1SPag2rVKYCSz5WTU3SIB+I2lHMt5MZj1tFZOIi16veIpIvHY0ThY5ns0mJVPa+1CD4opQCghHI
3e2oW4C7yKX+GzLD+SEoG8w71gpuFir/awF04sUnJ5dmy1r36gj2yUhOwTIq7DI1RqNvWRbTi3vz
JlBO0z9bfpRi9j/GyBX+9rCIeSIMEBp9QA+J+vuz+HSrUK5GdmUWyZdhAJdvKBJLa29cka7BYT9y
gKKEC7k+Ze3I3ZQSZmBVbmBos+SvGPd4zYz9LHy9UEyiqHxkC2VJPIcELCAYxtDGhjQMH/P4HMOQ
mv+q1tCEBZjfQ2er09tA/bvWsHIXM0Zx9zgnr0J6/LjL4ARS4nO9YOWXpOL16AUMu/PkyXCaEWek
U5d5/OcQJlvPF2fQi+el+4b4rtJ5E9u7oY+EVhW7wZvzloAWYB3d9bvdAWt1MKfJLGwGU8svB5Po
HD8rao8ucpaZ4ojnDmGYH34oOnKd0UapAcoV42MWzxQ+MH63ELGbxyKEH8u+SW39qqAjmrn0aub5
2lna0SfCqENX6VQ0E6AIXwWOomFaMv0qI4kdHx8d9Y9yNrNQ1fgtQIFmriCiimvzAl+SzSb9zqz9
j+chRWWeH2m/2+v7EQZqHHlN2NFbvQlMYLVbps3raBXxz+mge4WLtTS3ofxjM+7gNW+0KKpbssqj
e0AJfrivfi2j6iFL8cBio5xJjKJ+AeTOTwz6q6NdDQl0TpvumceIKJvq74JJqLyVsQxYqAbot/uD
NJzObEoe2SRtCQQl8ETZPSfEspEBr33rWOw7Xo/wnkkmMG76gbgdNXIFBbzpV2lTKKICQiKj5xdj
kD86+4dbeW/VsH3LZZy4BAAOeqtnuQLdSE5pGAcHbC4mr3wAB05UxEnr7YO6PEq1tJJ/5YbQwBWg
QDkNfY/pBJL2qDnyf6aXx/2sdJmi5esnQlnVDoaZH+eU0GPnz81Vxa1VfsNa0LQVSbS229dMarhX
913YeOyvFN3RIee/GaJsrnpfpBDEOxVV5KnFgcBCAHjTEbUPs68l+vp+1BakBRWW9t/xBlo1o2vH
Gt9/d6Wk2AhaPqO9NNKQcKa7nUBp6Xtka+g0N23dJoDKmjQXc/ozVNodbxqM1wBBwLw7P2Mpse1H
6URuYQ59HijyynO+L7V6Y5edY46kkg21lEbdBqawX7BjdVZ2xorBsZOSeRDKoffL/GT2l+FT1Jph
jWQTS/OHN4sc5li7zIYruxBSnzdXplxfMXRjBJGBsNt0/sH8+jnVRKrpXHC2YYExNc4fJTRivQ/M
LnMzN651NBX5LQyz0wnSsD1o1OXp/gEgE8k8RWUJSVNxLIrI/Yy6Fjszg8tL94acgUp9voh+Ph7O
tSRC1iQH/tNGBmLEu9E1mM0rP6+a5JSoWcq83l4JA8bKOafaTk4y33i++o4Td002bt3mjIc7ScDl
nH3XYQT+4J64pM1N7os+tffNGksmdlq4A/qkebX1KzW9VY7BFzh7psKIAHm7xzS2PaonsW/J7reg
ybEOc3jSIPSH/mGWAD/9X+aeyLjRFy8mpkUW1NXOWAcCAtcrj8G2jxVrNgmdgDXbSMPtYTHv8yEb
8PjUx/0RC9Jjx7AV34IHAiRJsk02mqdsmFDs1OasuTU37tAusAOQDfQWsf2Nyc7tareAuMT2qwoi
r+9jZUCoYgCGKy3HN8alX8nofTdsPQTh7/KGeU0sJM7bBe1rGpJCzmTOElQhHcAG4Jk7JGXAtrEx
qVlSr73Q+UytWcL2Mu0CM5C5gwM6y0b9gIWlxkURvYrSnnD6NuWKK0O1a1eLPfUihXmimrys2viE
5wOe0AQk/iZU6lzGtuyRDU7G9wsfvkYkL11L1PrK+SImWjnhIgA2SopvIv5O9NOTxiGFuPJX2ViF
du3FsUHvs+6cYbbdCYLtzGnkcu/entWMIdct6W92JxqfQaYl5Z0WDSpjw1LZlusG+79jo5bU3G4q
gTjGTKIQ08+3/SzKD15iRqJzu8IUQ9+xuoYNqT/rOjn023jOgiCkOfmAYz08S6tANkpmGPe2UTxg
Yu4672TG6+pY5MZi8PZqQABe4cxQnyZHQZln1hM1WzlPTlKhCSgh0l3RumQFaT4b4zQbnNPmMSZR
cK+XM6pG4CdSZHJu8nxbuG3oZ9BW9bpuTc1dPeqiIwh+bdH56CkXDuFXvGzfuKjjjdkIVJw88zHv
51Hx1/Am852UYfJpMLLaezvdapJoUvNJjKxkJjPgkY6bh8AzptJrqDsl3MbtiTihEbFRW9zBXWkk
IG08tbrQgjTbwwfdZ5lZsDBsRm0a0xx0B7gnD24Iv9H8OVZGAVMQWUPv+tRBBlP6aey8eT07v2Bh
nLF5WCJWDwXSBdfaNTdYrEZpms2Z4LQ6Ifp+VYUIIy8BDbd4CYJeixjngsXIwLO2o/FKFEZw7Izs
I09/C9z3nOhdvMhiV3PVxA2wZ/PQNSvXaezlJeV/CJKa1UfhcsMNTUtcJ8uLq6Wrs3yZonWk0lCA
C3nqHK1ymEx3PfKYjkf3eB6MjIogT6Wf5arCTnKHoF4/ya7kM2Cj+H8jkG89uSfRzeG72px8Or1D
j5QIZYtne3k0YZ0sVT0W6zRMB+Oqo/5Kjznth0XsBkLd6rSwA/whc08cRersrBW5mE7KUUfTVq2f
brnwl+uVHngfz1oYtRNoMIr+fVo2iW5hp4YC7lRpqPWQtAa+szlK4Gn9cFofgXBJsfF92x5sa3sH
Srox4zkNtGoEHjagEtQtBWkt48cV5TsVdqp5lGkP++I1xGlB3WIQ8UbJ1yOn7J8Wu9hRgyci3xzY
mYwbzHLgREtiJCpK1r6ISKHtsmZC6u2MkI0koLF9JlV/ttZPihZyhm/L3DDRiHCwSRQz2lVV6yUb
Gu2ABES8K01ARACOTwApOD+jUWq0XOt/uZ69cxEBwHzyOTr8tWkUdl6Ry8Om5QWYId2XP6ULfEQO
aSHURmEHlk4T2TJsOP0VnI0Uwqmpi11UAF3PbCQUBQpj3PG1W3+zHugg1DvJSaXT7U9mSyxEqlZB
LtckWK/EakzUeNA6QXNdWQ+EevC6IHYLcKRUdKkj7oMzvc+MOb12U+nu4gUP+8ryvE5CMap3+zB/
MLKweSoyfmMe/5YV16OWjnqoX2qCjm364jVMaqBhJAnd/R4MEfM1lCa8Svnm/UeXEwqSo6FsNEYl
4Ugfi2HuGhXHWdkKAQPT7d2CiAOHOt7lq0m9Qxc3uqo09+FpyrfKlbwyvI9dmc8E67mhmH6SRVik
s3yBqCz/nPP1ePxN0NN9LFi4iY6afcKGmeiUd6rwwzH1hMb6g4atkjjTxWp9I8oR9bdzv05r8UXy
pIfta1YHjCvN1syqwRD4gcb52K2We38ycJeMGuJmF5Tkq6TtemYJd7p6arua15v+L3H6J3TdxgIL
0j6iMvB/AhSTIqZgnSrPUMqufd0zIQSdVDLSXBpFWxNl+AkHy22umobJYGgmwkQo0hX/PtOuDTrG
F+3Rznp/OFF+J7QxvqPnG5ou5yX7B7OrSTgK7Q0m3o1ISOVH5HCHNmIQl6EfAtL4q+/XPOQhwBTl
Ll/6DsQtEw5q6HSSi9hnlj+d8pY+c6hR0U4ISMl1HvASErIhdVi9L6LbsRm0SJRqAMXNiXxZCQMv
mYn1Ow08RHfAecAzmBvFhtL9iNWlGA6e3quBwxljYBBZyn6J98/fJMA0KUOTpRT6GwVFJbDS/XKa
tCvSSZovbVglYjtmTPy0xtT4DB5eUuoVsBnRGIwCkth87jS1GBovaeVloVHZp4QjEw08Wc4D0sBw
xOPauRoh0JsPfxyvKiaN9TOFnjYrDdXH/SUK2Iv1kxijOEbaMdYtQV0iHy/EOb8eZKx1afDkA/UL
CXR9f67NAnsmr8SfrEQ7YuYzguFInfRoI2MQwuZ9ExDgCsKPJCQM+9J/Cjun3qeTNiCrtFrrOt6L
51aJIn8Mnuds7sHEUgUue/Tgfl6pnNXDBf4hk7bolgfrGVil4S14eXoFG7mQEMgsqx/i4jBNApCH
rAaWOKx+H9tzgQi3pC5aKZ/fw2+CIiEGhjAQdlUwZRwS23BCRktCbeKRTB7zHz715S3sq52/Rvzf
9+DBZFqDxA/Q5Lt7s3G4MnOKZYJwyd0nVCij0lZn92aTUGTPvE85EnQjAl0xWelIona3O/V/T5Tu
TONnlu+CuXbhsfzcvE30YK7ZspEVFsAIZvwFtC+OqPVHBbnwhGBftS2Zb8dvmD37B8wairw60M2B
vx+4znjapkHVjD2fdjpgFNeBrg7sdbwUXRzeOI1RTtDwgEZ3Cd1tBi4AqOt4c8KV5gEto0OfY+Pk
+j5fRjoUd34siA6dpLK0uuU4uzL+M09zYXRWVQnEtsd1IjlgT6nH4u7Jtw38EUrgyZ00HQbuI8gn
j4h3V9J8/17qggWpZV1/KfL9xshbRYznKJx/gjTyuolkW1EPadmqWUuuZ0sc7JvpDyaxnElaZ9rn
3MKg8Y96D3RWAYWb4ujD3TxWCsjfYljiNGt7cB/dGjBK/q5CUHfubfXXOwVQrEpHfOCw3bgLiXKW
GeYzWZVx/GxAkkA3fr0rcvLD9B2VaWv12j8JzpHm3ifKANrn5zlrCZPTvZVHWXen70mqILQffJWv
jizHllJNAcur5lJS36Xcg/XRBmzeIJrwr6ZF1nkAINnuIY/+Up7HjOrTXk1tiUEE8qsNaiAwkmeO
apgvCEdvKJi1dl0M4+665Q3Nn57mS13sAf0fQfrXyc/AOxdPLNuncC15AytNDMKekwf1y3REqQhS
cfagKIgoAhBukYrv3RWZYWk84j5tqM08JitMMSFcbSqxpkapPmdzk1r8kAoMoXo4viea3KaIdjJ7
GPvXdkrt1sMbcXV58eqBF+2zTiflCHjM3aAhl5Oe70qXxocrXhQ4i8c+iEwaddr8PIsVmcySPszy
9tIDxgyX6Oko1CUa7e6usDLFrhdmxcGQOmy6QfnhXSCqZyo6mQcKlzE5JSlz9YA8GHQ2BNeXNs2H
R4Db+kFQXgR7iusJdHWxWOxSGmQABOO8B593PIndhtyCZ/fa0hsuHom4u1zSDyiW7U7xw2bNo5Qg
LrQOg4frwGhTr6pge4iBIHx/4cOBJMFZymIISuSu4MaeBHiOOyfSMnzF0WkjSjKxHp2+SDXVBBQ6
zbSyMLVphV8dmdTI2jvZ/Dzyiw5KLA9bGe8x/4lJfsRJ+zszB/lZu+l76FYimE3cTTwUrXr2XMXf
6twGa0/DHCTBH0wVe/laAAiGq7TRfj7gm2IfeBPv5AHXf9OvyNUM6Clr7d9Ofgdk35djyDlvICZz
zoKq3GK2ZPt86YtK4gH8VvWERHvourRI//X6Q/RGwwld+W46Ac99Rn5Mh1+9u1tKkCmwUu6qZiRm
xOFZjLuG4qrAG/L3ZqiCnh7+RZMkKURi3w7t5WJfaGKgBEL33QpRjTmAiRHnV0DQjRBWS+X9ZC9j
cYR51dgplaaErw1XfDVhWFMiMHWmoq95Wvzzc8gEys4vUPd6xmCTzhZtE1L5Vj++iho7d7u0qCvd
GlDpzyyum8yZE+QI0Vjp1VQezHpYDSHZUBUec1hR5po1tSy413sSzyWZXo0HZ+Swl9H1KIpJPWuQ
p7GorJ/2YrGjNYiQkMlZcHm1VV7XNNwPcUgW68m624csDSJlWIUgKwHNSjNaeesY0YGlc2iLZ08a
xNVPKbtqWpU0mV6UvU65cOXQ1GGEAWu+6AAa82F+EasOkYRzNqK58b0kwAabREAwAGd7CYXNDDso
gYeG7XVPOcQJJWXaA/cF0GelJBoM25mzT6/g0qpn35qJtjbPrc09Ve7hS4cdlaDCQRW3g4seF1nj
68Q2UhkFtTQdZGxZBaHluqei5OSKf55DpWORRagkeT2x3lHo3jnFbH4vX++QzGaqbLC6+wS4Jdzl
J5+0BfTF29WWh/2tH/+gCXgpekMlmKvlgx8lhYb2WAlTHnRooIMyBYCq8MxwVG7TKxzHDiOC2raF
44evV5hVw9Zv3v0bO18DQhbWLh39YF1SQkTtuTtavq3AMFwelEtZfucVMM8PE1e/laSUDzRLWP5i
CuQTcxGA8iu1h6lKUf64v45q9LG7K/IiWFFmYPvoPeLVEvjEhzf01fRXRVUKSqHiU2Z/7Ao5auii
tUMKuMZ1WCibl+bef99V5GVaZ4I9M6i518lu9ohoLNO/B681bp0zc1Ne9aTTzf+KcQBmtqVnL/4l
nFY6TgQGiMvYE119jFGBwwgrqmvfTAz1iLl8l7JvhP+WHAmLUvyxWEtMdXIFVeOjmK5xg/zPbpWs
jCM49fy9XlssR0PNXwyP9oBk5Mo5UEXDlXRCdfS4mUaFY1prKgMXV3ZJWN2CRz/WD7OBPN+x2PJp
Vf5IJsrICyFINoSIh1h7zw3O+mf5GrPUF2zjFU3u3gb9+kNqdi+2heA/XYrjlY9iV8Xd3k9oAwFW
2GLfKl7wbKvGxg+vtRe1/wmnpAq98OHp+JSLAeQF6zlgBRH7eGd/nQODsYsFxJuDFsvOi0ldO39+
M71wEQf2Y3Nb1CmQySIOdwCL/y2v35wdPUvB/iWiJB3wzEl2fmy8uNYvJR9Jp/odrvMJKkGMqiew
BStrZI6Ogisj7nfMY48SPrq/vnWG2BbvgoUd1UKMiR2YWTb+LRePgnkDAG5wvvwpPrtz9UkTjYfH
VqoaUrD2DEEdfRjy63KS4GJ+BZyAUnmVOsegBMFshO76Gw/BBmmCJJXV8BcKQcRdj5A4OWUy9gXP
pCaGlcZgUFuSB5VmQj9yejclOVaSDF4uOP3qKcqksl/9NXxRu9SdB2jentqymX7wZxZxUbhHklv9
hh9Hx7/wZuQhl3N0k92eQ7z8j3Momm+/4gAKjOHyp3wFK31+A0c20RjFZ1nozQjbYQwjSvNF6iYm
E2OHTKWed+4N3gaCeA6Y3/JGm+qwuD9uq5tn/sOmfgjZ1ZPPLxUZewPF8vR2YKpuugZL/vSM4m13
5UjVSS4EIjLUEHaE8qG/C5dvha7YYJgjMP6N6s9vcvVLG+Qwh/KCEgohhoTMXnvJ8Y/+hHS40T0S
/kZVkEIpVy9lKZsznEfdAsJwqRnoCS4E5X7W9tF2+wQ+1NVFx+s1tA1ri8BJlZUApMkCI00PalyQ
5qq8YSWdqrkpNK4ULCGuqStDsXqO99U9V5Oan83knDbxTa/br45gRjVZ8dei80F+mWJh6xSv6+FD
lyxmDiggPIoH2jC+wZvrfJepKV/VKogWMjgCw52AxX0E9B4Je5h7yJqKuALSUQvNiIkDNAoJdE/h
mcGazplRgy8kTqaebHnsp6uAUKD+QbPqBTWzspLk1HI204lbglznV2v9ON7pGPvEQZROXn39U8qs
rcHFcxMnJGrywc3Wyy9Bvt5xAv9tyhjKS5d/LZzoeJXcM8UZPcRou7XLRiHGaNO6DTuOg9NIwga0
4QaXiTBLPuhkX01A8+BQc6Sc4IcywauCMdq/nfbfQRvB/iBdHSpSh0u8j9VaOoIyS2ddoLMCbkgx
VzVA6bV7hg1xfLHPNcjf9CsAS2O+4tUwXObH/c/2XVyNf+cTT6jalx2TBWpyL4LYIvwgGxtsjK9N
TKN1JemBFiqizNZiaevdSsGhzXRTjq97NLM1zEFNdtYwf8Hkh2Ba8luUAGBAYH+0rL1gnIy4CpSz
i2FYSkLEUNxXPoqrgbr5cNpIDLK93j7+NcRmRt0ZayV+KADB0vAwxsYIRC8thFZFnirOa74ZY9pp
jCn11tNbNV311pmuHMbdkh5P0xIOc00jm/lI+BXEOxRt/hDqsPUUUEbdlb7kRyO9XrKpem3tOKpL
92pwS1EJ4mAY0N37N1+QLUISy6C6KpiE7cCIt3g+StMSq2tkxKAbKvchwU9R020H5DjYopcgItnU
fggR9cVzQF4dW17z/rDTtHIiUcU7NXTQm41oBuMbl820urPLl9Rz/rVwzIxYWe94dLIa4wh541mg
GNo0hsxnJgsUFypBG/T9cHcunTacuaBc0L00m+C/dqo7J/UzuwH4cYBGIfoB+Z6oEhaBD28gzHDR
2YBhydmk/jNmUcuzLr4GT7wpOV3xZl0oiyofrQpw0Fjcf1Lzs0eJnGSvDLXrPSpSRdUayUSPWdiw
VY3Y8EE19tLaMC+YjbMpVn+/bZX6Uk6KwZ+SwrsCc7eYb/t48lT3odprnqDLhQ1fXzwuzekoo30S
mUHgGXUIqaf8CYyJrEehnzkuQIibMfgmlYa9wIyS/P0S/a+Sf+ZfuJws4IHedictIzlZVGiunuZ1
xbX4s5Mp+RKsVQ7gCsKCMBLRdVvZCg2GEN7I2VOOb+IGQVM9/MsLXRncNowxKJoCcaMknusdc1Kf
Gx+do6QKg+PMHnuljIvGyADrkdpU1L793tiH4mVn/jNsSuDAZQwTrlOVy9RoLHh/WnkWJvyypR69
D659ExLGYHqiV75quWi/enGSC7pfMbLi88LpL2TbhLepXXbOamibh+dhalnQ045Xrcz6S/kAsYu0
f/0mWLjTpIqg1YsZ0MgtRShZmdQFRzLF+o1zZcMI8EPBAcynYyJpCUZ78SXbQxGnnJBcvOa3a1N0
zY/DQKLW7Tx3JUhplwNVFYd2P/Ou5kXLv1+vmOd1pq7rna8hxoSBVVctJoXqiFO69vO2AHANntyr
XU7uacTWy1AQ7YQf3fezEyQozcQ8RwhE20gw8M62TfiDaYt83uW7n/TlPppOjAeUpCcRaYa9XmxT
OKZBH0noPNO1mgzmdmRly/Q5sO/xqWZc8/sNuAOu3wEqw4KV0egc2T2ePPwh5KC+csw9xwuR+5xv
bhHgB3u5+2Y6W1BX7S2Hiz8yFZ9YO0F0VnlUkveobzVPhTnuWXkqJAiZCv2NmDvBLLP5Wev57EvN
rSOz7RIQWetct3dFuqlIDqYc6tdjubUSE9bIqKrwmp9c4WXCbCn9pNKDfrigYcHcnYzvgrrP4+0V
mtGenhsy1l42qvYSJlQ8doLU2P5ozRja7lSCwPq/cz0kuJhQxHSeiH/ONdvcFIlR2uN+SkvZEXID
cEo/K1141V3nVwviYzrke3wpKlf0Drrj4mkgpxWoQCNOjjwrdOMjPiYViS8GkmxyrmWacGykfKaw
Yn4NV0N+ckBKxYuCPwIdf+J3pKWt87/hPsiAjWLu+vBgNWJyEgR9ZwzOLQ0i15/+QwbiM6n+wYBg
TqbrDexaabv83RP1leSEeV6Z5Qq6F5Hpsa9PDjquuL6fQ51JtnKsYO31AtqeQmL40CR9glCdNxsg
wtb0V0n2ve8z90ZfcKgNytUBzVPuvklDjGN0PW/K9UWgg+blweaQfIWPy4JrnayQORWutKFxa1EL
Z26YS3zH5dtuxH2oSoAltFaEifRuI2E3ZRGngHl4fj/OZfCJqDM8jsFE+g7N2z5NFXZlGRq6/J/x
xea31a3SyZy0ts8LxK9UlrvCHUMAnCICFoPQhscfCHdVilInAn4IcgDsHA3cXNb9GhgOKkKIT2hY
dz4Cy7xLWg6vB/FS6KyZoYWPqZHXZa41LPnktnsRAI22VayYV+GCncVbmEyjyBfvBIOBWWyyi03o
jqJ3FcrWdgEDQvPSbs4vHV1RMCuUKYw570KGSlzW5S5hOu2nrhIlJucgyrH4GpWnN9oKaksFGzI5
VZembIgRNiYVHPj0r0gFQRqYbAfypz/xdmLSQ/kTeIRhbextEuG5zz+MbfDTZOraecBFgleAW10K
032RTUkH8jgiFF0lwmdFXLEMSk0JVqMxDKhzfchKONan97ir4YLMGJLBfsbKwH+rPAjyVfNoQDzd
0LtLxqNgZ41YeYor1WDmHd+nZ5LrJ8BigrSb1X7PMzYfuKKJNmUrgOXGwCKETPzayZTZoyzklxdS
vX2bZOOAP8+1rdLj3NpAOIMj+k/4lOsqYE45jxmVGnmsLivR2eJ+gG21zDBTOIqC8sPdrOQ7cE+L
q7cUTfnIbeNbq0T5vhRPYKeri4i+9vY79ZMogbhn2cy2KadlIdewNg/3i6Ox+SZLohsvWojA7Fmc
0V3fXbABI7NltsoNMc9vuV3SnN6XPJSat0Tr+5oWBZmty8Mb17ex88tW+FhLbyZOFP6yhGTqaw21
Vp+VpDLTMDJmNNvivYCLSuxK7SUbfX6bBkzOi3xY0MaELcJgIkNj9T0hfDC/5Le2X/E3M7Lyamx8
uizqnU+urn+4IWD97ZDXRsqXXMhnZmg/Sru1rLoNLZGSqmVh/HeTUnxn16h9SRFVnKPPqG4f8+gE
qCiaBGRX2Q07Q7vo+j9/Rj8x+rsQVGqR7FsnrT6kdhQhb5ne2IdA/8owFthNiTYG3cccJnJtOkSf
+y7tiYetnPTmPdiJP1aV8jIzwcuzkwRoU4Yih13smKdYqGQsDkTplV5wbUzevUuBppchbRzkyngM
PrJwz55jvQmIDfj6sGJFQNuqyDRn6yqwgf4Z1JChGntM/qct6xSCN0GCoRDnsoAQ2wa5StMnmB3u
k/FXwP9/4rg21iqXzLHPTSi81kIWyMKW6S3GE/afri9uUx5LBX/75+AJLdfXyOdQuBVlVs5lCgJi
QezJUNTHrZm/PT5JYFE58GIEH182yPgfr8tNy6nWTyfnSaswLS1lRzcOQKhHrJdVr00y6sKAZp23
A0DYvPDvIwFRgTqzYpcF9km2zQpPMaz53+6BYW69aXp5z4tEtaJdsIJo7DlXvzMYOHzoWZHB1PJx
ZBqq35j3vrn5olk4sHyee3KzMgowjr9hUytmdmvg3NTSQmytrMpAk2LvYP3gnF30dlX2nwYEDGWc
UKzuropOsz9jvmjZEezgPk4w2iz8tMNTxxA/l2rDSHoAbCZQiylP6GNbpIYU9wLUljXTRTE5Z24g
LAyGqW0mwGC88MV/rjFbn8nJfv3IUJd3eLjq8aTkbXCj3TL9GWHXUD+RdIYn1rl7hYh3vSdHnzwg
v6efR94TfWXM7dws6i/8Es/rmWCOq3tBCOoynXmj5/bPctrhaKuUZ+LZih+ZXaIEWMwIZJ2kDfQG
1bn72vcm2/S3A3UwL5slDafHB/ka6qi9h+HtgpJPVzH14AcsMicJKlUsRHMMzrHQbGREVGZG5kWB
AH4hKxplYLN7MG/Lx0+pBOrsD5NuVA7FDdT/9FbNVM2x/b4kfKaPzHzI4tD8asFdZuTY3g9apsTj
JJ7nUXF/zrCrsOrYIctSOLPgZOxq/JhAdukRXFz2cFM9D4LnZS46tzSVuPv1+wVj332qV/x4dvzK
D04v5YlST//M3TWOqAkVj2Qx4R/a0U1nC/rgU92H9rp7Lnyvbx0G6gqDrEHBKoTa4cCYHVCdPhcn
y1xOoBYT8zmhZN01TF9Dcuxy/lgnKdykG2Et4Ys7LHtWwZMt2TRquTpsoXkcQFjkgoxQfh3vq9V6
Q0MBvxpVEB9IZ0w2Ou5MdVUMeIEJB24NzIFUV+2060qwycqKLqkIhneg9+N1ggZfU5/t8J5SY7fh
tGOfYpBevc3pwclw9zkjXcX/lpMoqU3lRf2jQSC1COBgd856euHlMG7mIIcaDWphIB0pPFKMTdhv
kiuLJP58Xo4gTLta7j/+FOzvjlmxlJDO+0meetEl1P0Jko0JAbxODpHaOqLNWXb/JBDZI8nSOurm
x2rFATRRDranGDWB22FSE9muxa9TbDmgZfLMUtKZsKeKdi6ar8g6NnWGRqrJtaaFkSzCyPegqE82
Mmbb9WP6uFs+0MyHaZusfNKx3n2UDCaDeoEnCwB8iS1eSpl3xUlHmRlZu4vqr20QVxjpWXpVW5Mc
ubFQnaitwnPQ0DDRBzSMqKJPLIXR3Mb0zLEjSob6o8rJVBJRl/F6SZ5F4p2Ec+X2emdSkVL1oR12
ggRlQPGfcmnQ8PY9ho+iHxaF8szdkbBdU9TDATrVBFHrUnrFsNIP92IeyL3sLPimYWdaeQrsHpLB
zANY9gl1hf9gzdGM83rYKD+8wAzVHktgUJwAmDvxkF6bSQ97xKWJph85umATtUbyor60ajnBik2U
dyxjHFZ/vNSlkF1KQMVaCAIU5X+XycoH7p3S+CGypJdXchn+5FuPfeeiIvEc5Ob5IMMheTjwNR9C
T897xoyifQOSXnNprdc1xnP9maf/RQO+EsVhiFpCWIWJBcEV3qoAK25FXPHNck0J5RgpNNDP2LSg
5+J4duaM38htKYA9aqHAWDD1lSFrOmNmhntNYhqqrJv5RfIrJzDH4HL86sSFgMmOqjbZM4vqwY1D
0t4zY19nFHAzAZ/QwwKB5wZwQ5yXfWA/1WnbNelrJDdtUNZRPbdDzL4F8RtFdrofVMreW1eKNUjH
/oZL2naXUan9wfW/nGMnqVPI4C0p71ohRbunQAFg/ik8eRFP++HA2w1N82DsA8ZLdCz5VXTIlbFk
Eqif20R9+SmpNfYyHpnM7Dpd1KCJkIoEMDRLxkTvcd4t9dzEdPjd16Wt3v72lpfy+Sy7Xrl8b2Ko
D92gQO59MP6buMohTfN9wuRm1z9Iz49sVRMo7oslCy8/6rxP5v6AncXgplqbaqF2u7jenuNuy7Ae
ckcvN4j3+3ZPdhVg3y1uBvD7xg8Bkw0qRUGlfd9t5a2gsSnY8NfpifCwUf5F73bfPstj5SM9uVCx
sWWgA6uH/5FTynkL6II9iEohQ4huHS+Um/bfWbxtHVt6D2ns8+cn3F+jfL1rVZWvDyg6lcWgPXCF
IgNFe96QP6OBv/0FGoEid3rmuWyia3fVrVv9wtm0OMsNgbVpxBWn/nCOIDJUt5DuevTo1GeRJfsR
WzM/jEE5m0j3ebNdzIdzpqteGUndwoqasF77oSOnMV+BZN/0NrTt23bWMSrMnhbieolUgTCh64Oh
6wz2RYo+9CYRpK+WWOR+Hb3FJ2KoSTL8N5dkkPOF6OfdCXsf0XVr7UWwUuqWusGBlgSuxUHWTkMp
Nb84yG358CeRwyVc/0NT9YTzmd1f4VoXP9vYQq9MD1ZbESWgfnbuoGgC5rCJWskpR5khmNhLwbmE
1cUom3H0Ts23cfASTPk1Scj58xAdBA4tNSJMdVUjQr638hP9a+GYBBG20jNNnJSZFDvF/G/tNa/O
Q+oo9wqxZewCTG1hfW/h5FEBBnhyaCJJ/X87p7j6zWdGTQonp65vroky0Q39vssYuG7rpRy9lrEZ
waJqprDogVRcPcD8ZW9OaOucT3bQDv4Hpe8gAEk9O2l+8hntfLVStCfKzpvEBBH8LmFuazFgZPWV
Fm50WFSam0o0gTk4//0jC/xDEb9MJat9uhY1cWIACNR/WmR44tT4f9Inm+TOi2f01rrLecfc48fB
5SL3tsjw7VBQu7+Cx+NYN0V3Y0zTtn9z6oDCHHAzyplbXoK0FJNOezESAFTyomdUyFAVYS2MjnOI
CvqUJsvfQ3eovDZyeL2TteMxpXeapEHKu95xB4a5Abp/nC3Gm4NwDLgPYXr8sNq8gw5EeBwtEZ7T
gXEgaHaaZZl1/+v5lCc+YaYrasPBL0Es8lTjS0mjpugKVXlaD2l013WAHj3u+KWusvFkeyP/YYZs
S+jzjU2fhrzsctLg9HdKfkW578ac/xecE2bK+pIOiwxPoXrpV+JyNpXDvMXnM5ClEoDI3C0OxZTO
Cy060bCby8fd34Uwwmxa+WnX53VFaMl+hmbT2MpxFRAJnD/YT9PhQWGbvZHs6MQLCfabnF+O4vvg
H/GSaNWjiofYRIviy9bWfq4fc/ld6JIe6JYO+Bbn4TyHfaElrfg4BafRUMl+cUlFv0qCW8edLR9m
3o9aK66Xce+eVXRuGI660Ngw4QrxJ17noJFZELMkVr0hQf3TCNW1ZTCdhqPyiIbfexHTHAalGuNw
jUlzVHJ+7/PsfDIR+5G+5mrx8u0qm3ILjcKw/NB1oLo2d3MKa2IjF1zrwALNjNPzYGFf6B2NBKjn
v4AWTG2klvZrqvJ71krxezxoRke+QkpF1LRp9syh5srk5MOqEiT7SvQxlo4+ZM7OpQO82TM14mEN
cXySP35HlOA5d/wZkqFjrh14z58GvCOaqENQk+pcUPFDCHOJCKHQjbz5dJw3Jy6N86JTjDR2z6Mm
A5hbD+uftjfe5/PwTp7x9W71zlcTmDOUBedmLzffcXvSiFsnAQdmJiOUlGK1LZaZY/39/nE/IU4l
5ORzPjGPmq1Dh+ZTuaScR9q4huV9BFfFPsMxJQMOU4xcuyR+nbL+uDR9/QKyN2V8TEawZ9+ZFyIF
1E21D4mOVllR7/GrVlNUR6mEHB5WzKiJ4jtOjK96xIQVQtEwOIjubXQulk70GOwkIYp/xSJyLOSW
YbFyF6v7r+SKrnXUYXdXAwvq8ggAy4S70XEY/JL6WKyl6D8bkLTtL7bjtwqr2OWkWG0pREgLmG93
vjDgNiZW9+jByccQzoTgOxzfaxoRo1MjTgwSuAtpPrXvDV2hWMuba7fdmjTp8zgNsxJK0R8P0zpH
ucPBQuU/WpD43i+vHIUVdc7Uwlwb3I38s4oEvKA3R1QZCVkXLqL9eBTSeYJoCLBi1YHqcw5JIC2Q
3czoYZFqm0Ol6CaeLpOvUZeooAF1FNHXhfmPwB9pbqZGuu3vW8jzEABygSn6vpyQ42fBsWYoHECE
ltjJCA+T78r/Jo1JUzCpmAuDN7mss2HS/TDbdIg1ARxJjLyCBUykr0ND4HhWO5DkCI7uXHY0Pp0q
rEYnycSQssOZUC4JES+4pjnizZzP1Sv3rVGFqCSBKuHo4wBYggw0ehQc5XJkdbkp6qNn9SpAFX82
4Em4oJFNGNEwj0s/vFTMaw6uhayv2UP/vav3auMiuH3c3++nOY0rtDC18kr/vZ5eQVcqs7RnA4TO
wlP9H06eK8hz8stZzvub7FBDFU5KISwhQP+kHS13OqK5vRuOMT56MRF/+Fl9ct3e9ZmpX/4KVR5b
dmRjyKg994ZNs7u36gL2BRMIf45YzyGAMMp8ZsPGvMFp7ylHyerW1DcFnSisdmR6Y6HE0xlSGEqq
shNJSuZZ/6sOiUDW0gtX6hwXoWCWMwpLWE8cli9zMJsg7MtIj0HPV6j21gdf9V7E4JxxlbZa6Wqg
EpVDMqbIs5jW/k9pbNjPo6IEEsJM0I/Rl1YvQFiUxzix2YWaYVRb/448HmMKH1fDCllznna/WYJg
lO/EWrpdscNqTC07XeJKXWEl19V8wPF1icoK78kACSJt32M+ngaxd8AKFtFCF8upECowr+GblSp1
r9T0cIbdill4VX1PxXlgaz9RrMuiU/t/MjeDftnmlw87KVjcOpC3d6QefKzmibNCu8g8wHBRP9QR
mus8PgQ5ZmyJvMh7cUMbumd58FWBUju5aFkkixcJPosddr+qGE19BjwQc7S/6mjOZPEi0ODO9BmZ
+4FAJRKLAdsDdfEBgnWNBuF9L2Ern2SnGLrBAl6lk58yB2dDSC5xz8KYsljgGnrkCZZK9KIfGBto
0O8d0QS32P2pCQjylaesBiOWVebDJNnB4+dTugySwjQz9EeI7sU7HovTOVlHDpYccCuc3qJv9MWK
a6/YflONer4veDXWWtE0rstJUmNdZTM/advWl0/NMPjNfJuFIJaHV+Ddd/B1L70QfJ816trm/0vR
6BYRFqWvqHHO49VJ28b09FCXvDNpODY4OGwpjdDmUva9DFc4TrydcYhRh7K00zHaOySSl0g0Y/Ul
y0C33RPUCXqCXaMLtqycxcmFJ1Khyt4qFGd5mIWz9dTe6hpCok5oC085M4w2b0Eu78o/s6vtsZO7
OGVxbsYjEitOMDqBXtCDHLsI1GGPlcHw2Dfz797mIb4mb0rkVzXkLYLAZKIHJBkm2izwl/InsNfp
YAPXsezBH47cfoSContoOS9IIgZGTurTOhQ5oBWngNT4NuTtPdou9mbqK5OMV4AVApVdZUTWoNcW
VmaaAar5Hgv9wEEKvGR8W8BCC37pruEbCG+C0fEQ3R7aFD2dT8oxIJmV1k8rO88FyokvwuEHGmlU
ou46g3IehMxNG+yg25JmjfB6s5Vxh1jsyoxXbfqIlTnfS2/+HpTUTXSlk4odBq6PvrwRldPEVNYP
ztIeUHjy5zuoLzKOnNAb28SZ3pRsVhLyY7/KCxKSzaYJl882j7cdLvIvlCuhM4h+JpxL9u4VZfzW
BP6pb7E9bVHBf454uMObRmejolT25PW64PrWB6pOLrxFUrje2ZZkn23eRIAZ/qMI88yDRE3/pHdg
J5+R2FmS5/BibwU2GaGIVMiXa1FsSTGYL1Kn/QXaznAzkR6fMwSqnA3qbQHwckj0GmBlqgCiVy/F
LQzH4EXYLbMVD0yDylNymvL0RXbQsdA4k0L3UkRwvOkZ6rU8jGgIyeOuMF5LMXbzJwtJoUNJmRD4
JR5O9TO9Vcm4SOofKePQDIiEdypMmPzEcsNXM3bswH0OF90/2rSToqO9gkzNzitUH5J3+OO5WeZ1
ZIX/mLqcg+PiyR2soyA8dOypFGivNAJeORDAWhJS+pyJTyIlwI1FkutTCuI6BJEm/zbrr0H+dlHG
6t4lhQVEx2jKOftdvgtUtKO4dTOTFpc1hq2OocbJjFSI8Rj4PaBYwE4fqZxUc780Jf6Ekq5zXKkV
/Ga6Bg2YOnEAKfcvZZMiyQGpFyicTZ5JzoGrlXfPNaPeMO0h0fmgHRBepaZbipkUwAQyi8zd6Np3
4fGRWhfd25KD5zHGjWfaiUxdUs6W5i0hN9xJlYkpy5RujVEcQeKYDKG6+TXPOxfi0ZCVD+KqmiHK
oU6xZKtngwSmH79IptgFdkZyAHWGdB4lndYRYTyO3OUxVRRK3Q1Zzt0g90IVvyGLPnECG/LpJmyU
R/TrD/Qm1fuf1uaPuNfkKKnTpyPjlodqVfPX7Uv8kvyx+npuiXZDA+c9NeOQIVMSzQsi9/9Jk9qv
0LKhZOyoV/cjHf0uNljVZvcRQRbA4N8Y3t0tPKomc2Cco6vKEL0+W4fyK+sOx36sKeoXLJcnQyab
hOuzoMXZ1Ak7NswNY3Tv6CFB/Wt2RGGcRRbZVqVQfx/j4g9uabb+ZUP0tfvo37JAHjBxYNEs1KDK
O0foc7QaxudbnxikLVekmcxfFXqAEnYgTLX+OP6jIp/IJV8X6HlAobGuS+WGYaHrZL58LpVlKjke
eOzwoIq4JXVjsiL+qEBHkq1eQACx5PqtNsxFfasOWtdblQl8d48k8om+4+N5aqJx5fSecEB43Ry6
O04Dm0AH/T25uZ0DKPTOKG8ZBRnT017qPZMOQQWR+aG5XvnaluJ0lxZVI11nA9U+Yn2DPDjd2TGe
QiOuYzyMCYz8hxV3lB53jOWn9CIEOZwdKmcmAY7INqc/885vif4sDh/u0mZslFM2Na1zZpaIS/Ik
84ONFx+Kz6Egy/MnIg4NEabdhHCObdbyO0+7+954a83VaB31TilGG1Kshpi8SzqL71kbFfGNwqU0
r4or53+qd4pqLKyRuQu+agHFCYo1MzuICkvC0dp4s+5SW+FjCYUXIPj+OPfvkv9c9kNt4ja8F8cv
Enkekon5gqmiBOCZsQCXHDIGs8bXw0+8GKtXlai2mFKTSc9aN41yZP0qwiLLsj4UD67o22u81IPD
BKqTPGvj0nlYUrG6bU+WI0bxMXex4+7Xs3k9oRs9v0uM00p2js49yK4vBYHLwlHN10hipjAxiNK6
ttf0ZInKEig8G0+aCIJH/pBZ9xNamJjgsW7z06Xvb3KKgL3XmXfwWCHRI3en2DNQBMjisj0MPB4U
SQ1NY8nTFi2ugwmjw8jbDr4ZpSK1LvXniX0gk2tIJDIfw8fdbaSs06zVgJPZq7qRAzVyUN9bpJAw
lLCW53UgoRbo3vWsmP2gfzNuHkOmgaeFmBSZ35Fvz24qB7LP9d5R+HskbhLgcFKCuGwklwLpBdYV
jIzCLMYYPjUoT0V94OPq2YmCYgTSRNgy/vp4YntPSjMltnHgP/ubvP5gI9dhPrYJsIxQMv5/GwAP
Luihve6pCeX8c1JnoypnDeLuOSAfoC8PEs43y1AZyVR6AXnQKmbRL+7Z8M9NhjHNkB11qSoYwEeb
mdRNHKhgkAdvIuWxUlybw/5J24TyYmHF/4ZYL/Spb1QYGcCqGg78hr+W2iH7nDqmNGf/q8HdbtX2
Y/kPmQ0m/5uEkMFJ/51foi0xWuzN77zlKtHQD7RItqU4eJaBEZ4NdjHFyuqH6nVd5WS1I7be8LBk
O/WrNjMWV7CUqhDg5M3RG2P0ZgoY8QrjMULSPNgyayjLX55+uuYkkrmuEy6uQJaXwoGp2NV5nUBG
/WASU0aCElKQxyPwxrrCcn2w9b4UPnYlJWgUSPUzuWgu/RS2LkbAEB2KpHMR6gV80GxmaWzZn2QT
5DFxiwYM/hhq1KTnc5jedb6zjTycrfVQo0lyuMtqcbMi1DtAlYGB9i9+PMlo3ha4sRErPYKMNRzC
Nds2wL+Sa2rPP6jwkTHD9ukm6Aici6ElQFxeLqHuFw3YOHk8NFcc6+gPXpmK84tz4pNuuaPOJYZ2
DWxdBFRxlSb9MuXLub+53LOOIjFG0kznYFAQR/N3LqpSXlB+7nRuJeNU6ph4gbHHalfyVdhAQ442
A8Ka1msWTDFbRsophoEPOKW01d7KPA/jOSridQJsBsN1s1tAcYLBgzk/NF94DSA+8BhMbXNS0agy
etr7BNLS/YNmNPBZsXxVwgN+FMWDlxe/NbmtnkICpZNt7BcVQjrUnjFQpW+Ya0J58rusGGP9JJTh
6OqDggGJLdtvRsLxejHSjpSuaol+jeP/Vb7kZYm2g0dZVCowtDHXGbfd3rpCMkyQtXwTNeByhck6
rMAK3btt2iTgGWttBM3APQc1JUqU91y6mAJqyvM4hcv8btAmpHJJug9/jvY/udEXEDWBMVD9koCO
+b4uso6ru/fj7iZUfxWXEauo5emj9dCM1mUzFHQ8/7HuO2SvpOsB4TMNt9enuvcdfrCr0tHU1xsn
rbLUCK7OT/s5pHGEjRBPBFnzorzRcnenhD9xTSVqBKronYFm7uZ8DqDpeFviIXYCKlCz755IlwYP
ahig71PwLRdgDRkQDPBT+2yPast4wBDukOnk3ale0toODbiGiCyEZ5qyDum0eO2635oKGi1PmDNJ
0S3MIXRJ15VSm4NSci3XjXSrkule6I1j2kuNaZUq9SAIypKopgeGlydwVl9ibLcOOpdXwA0nrQ7I
HXiSknVyUK0PtITnDO8CnzdQzjMTr8suSr6E02tE40+xjyPjyCM5FrKNX7n5mBkZyk8fOUTVJPK8
8mNZ8DLcQRlQ1R6AutbsIfnGhnz3T3VwR3GujbTplEGhcPmOJxR8tr+6z/45wSi0Ns4IT2nJkRw9
H0sLBbwQ+kF++TCKy4Gvb0r2NL8u8xJ8bV37RwO00G3BBSUoRU/8lj4V9QVcBbdjksjbeSNySmT7
1KYB0FazMRd5GsyZvSjt5qcdjYLoUY4SGWD/i0Z4nb1DY0tRYSf2XQZV1wQ/peKYcgL/PpjaLKaE
PgMd0KA56U+1rjezEYnawnoRndIk0pP4oM7LfN6/RsJ8s7wWw8MQ+soMz6nfg+NeP9+g1ePnV8dc
+WkXrTUSOt0fwprhQd3eum5v5iX2+H2/4wpZwcqejK+mMP9KPRo08YtyjloQuJC7N39aglxABPnQ
QQQSy9/p6LhTYRTjVcgCUl4oPrLNv0RHhOcIUHiWAI8kng65D3xDFw5PJ/ykIowEHmn0bb2gSLuV
la+Aa5WdvwrxSF5RniIOq+Ax1ZCgTpN42KhXEjLJkpaCCttCMs5ZUqqtxEXvLK/6JSWD4Lqjhu97
fyueKm+TBpoQpK2P546wSSd6LmcdwQdUKaEzwZN5XnZ9Qjzn3wjSsoimQw2GnBHO6xahxt1sI6UX
WlaUXUENvp4h32SGBcrFQw1xvBS4JFm+YclV2CrpwsgXjIRZ9Q7AxabpegtSUYtCTtHff3olEdlu
RRNOP+KXA++REJeulg+PfTiNmkeKSqr1Hpk/nfmtSGouYr+GjSPgCtd4jRrkO1ycMYCPGEOEYxnO
29m/qMTauACgj22o/8wPwYLag8L1VPzAV6Dgo44rWyx+1XnrsryQpiZWl4QrJkHakPAl0MFeh26i
ye3T/SFHKFBJ38R+Fd8iqqhfBITdCIx6+cl1tg2v0J7++sh0Dx+YichFA5OmfoBoOcb7+M3iz0u1
PoyJCh/9DomQGq5j4i6gFXS1pPfTOUdXU3sT1ax737QnEj14cyqfo6/ChcwLRfCT1sPL/VUUyMAL
BPoSoYUQm+PloQccr9yLPZfQTCuKY7IHHo7+cf+b+/LZMXHot8GgC7/59c+E+xpGn2/IGP7Yv6h1
7cloO9tIZq8rsHwqOUlKkmx2vsKl5qd4iM43azOHfiRv+JFF4ctOG48tpCS1hFLAoBAg0+ZO41No
CTrp2OHyD7dLIZ0fmqyfEkDb897SzB67NaZ+l0tkxE6USsXFqzXctyqLxBU3zHxRnvTVmuzxoP8v
HnZJm+9JcTMBhLUd9FyUQnYI4XqiD0xYUhGKlVLFuYTMdwwIEvMK7j241A2TfgIVQswwHpN3btw6
FBzXvXtLAIwmVgU0wguqyvh3ONiozjhcRZh95F7Vd6SBmFfG8idybjTCEEJQ95U+es3xBUnLPSw8
n/+xd/Gs896kR6bOzcERbVezjLQnTUlpkC+ecZmsIXVs6nfNbDcqBSpuV96vNP6RejjWLJ1BP+8+
VzF/WZvkk3IqR9Vl0iZoQOPuLAOW8vqMTQutHTHDh7WhIlPJ8pK7g1M1lhJD7aRUcd8rZOTJfxcr
VckUCuOjsowhkN8H5CAz7z9GFaEpl/TTojo/jFI3U3iTjQLdoRQbR2YHNykVyj8qdR32p1t7flV2
EhLDC98IeEf/DOu15WFsksZMjJ7dt4Adr0uyCgzn2bF5PveRYvCC0CTtc5ZyeapUcfBljVFRrIhr
LGr0AEc3sHDy+zjQh844IqGMYMke3grb/qgQZQZGZtvd+hEoSFrsLaZ0R56LQZbovTD7v7Af21s4
CbWbHw4Z6CcGGO8k3v3xEab4RkTgA1kzsX1HpcltwSdV+g05mb9uAXWIQNy0BePAT0xD15KFeUuX
Xw0hAT7CYfdi/+yT2ExgBshlzUVvSyR7I1Bz7JT54ltfexdUzVFQ3n4hylOUcqgo6vHp6A1M3/KS
PdsQGBM7N09x986RW6DqR+UUerkprCq8ZVbOgdqU7yM0F9omgEyS6xxVk4y1xml7+k5dujUEQAVE
uqmYu6yn6N+gPeFev76kML6NSzw97ZEnuLETJ85CfvG0N+ykOhKF5hSPYDpPJ0dRXh10bSm2jWSm
BaPFsOJKbbzE85ot7h7i7UEm2x7urBoJHjOa+YH+DSp4X3Us1s0p3MD/8dM4+ApQX2jB9uqj/Gcq
BSBN2uk2ETY6VnvdBJ2xj8vcZTmUEJwA08GaXC5OqbEicyodzlkCdurGzbZN+nsRCmPDH1ROSMIO
YPxy6hHy3kV7jxh96D+/fL+HxBk4QmqNzvSoi2YgFUiXanMtqQd9PyPWZ9jOYsjei9MjZJyzI7Ov
PjJStDhiBtLJtpHo/PB94+P2FZTAe2220UCvcbZmhMozFibrnneLyg/VPU7ZMZiHHNoHRXNlLjSz
9ZLzUVy19rw3fWLByp4/opcKkR71JvzByu8zpv1IIqB3Be3Ts3WWWZp7nOVSCG5eTFZTUsZwAT1N
SflmxxgXdOsgVUBvv4Q6D2bSqp4jv9V+hALOW5xuQCQWbWEqHej4cVXyWZN5QYjLaRanYsDeA3wM
1rkoGR+aoMu8msf4N/3TVw5nSDE/XS/iYL6LFsiKL+q7mkYh5R/4vK8i6LPajkNJpr2RN592Sptv
hh8hv318cGO08o6rby2B5kohXkYc9XwGSPVIGgJ7jo3fK+brzSqPCzRdRtt9/w/vwU9LWW3IhKCz
cyoUx6h+yJjemBEB6aNb8fZUSNHR1IrInwS453yatGL9J6LdDQO3Owmq47R7VVzqe6fxMjBW9MkT
Eh/Dy4MlxHN/Cb5CghSsFjWcKnNz6saJtBJVWZ1ymuHohh2UytRyj8+mXEJgBnPy/8KGjBLzXJ5P
BDfQZ4vmKF++ZQJr1hkIWKhviep+Nye904UB3BvbyKdR5WMY2bG7crj0YN3A1p9tPgPyCufY7IuM
2fRPpmNUQiNC8w+5SHRZIGa9z9HyyATYWqIl3mpuarlEZaLxCxos713GbqR4ao1OTif/ZY28k0lr
QrqAy1t/GzmwosJrxi2bwm7KhhG/Gia5zV+IXyhMpg23GNfnd8QS3Wpvg51dDeqxT5O8mkl4mc51
Zgmi4/SHktJDSezkVZm8OsloHLXBPu2tKgynJWUWJAgNL+76IBpYWm0el4eUcGipo+BcWDPTnwFg
HhjuxjeuUdKiQnvK/Mvv2wY24LRSsONew94+0hZ/evu0fPEQxaCWh9eQzERAHmftfnPUKfbvM5fA
iSeLM4NAdSxas4GB+cL73C8BjT0u6h5abIDORu3aiChgJupeVRkT+Mg/wl1XtQes84Zhvub4MnQ+
8dA2Ob1YvvgX+1YgUDEPcadq6dfEulZSVBfUJa3wSXu+0wA1jL5nIhTM3OyFD6nvccnpILydFoX6
1IeC3K50kaRwxQSE4bZcymTK1teyO/JKSiS3/Qxydn33n3mO5N1iP3OECPPhjOPLzG1hDXLh0Xla
ht7rXy6jd3C18xm4Nb0h/0QzAzelTMLNRZL+qlrLI+bGZ4cZxholeT4FDYC3UtRlRLMcyvoRcdHX
C+e289N5uAP/EddvKtnZm8pyU0qswSOcm4jRmw7alqVwjYR4y9oxZeTjZ4eNCtzktoooHMDAK2S/
2xW5c/eRUNBghgYxZCiHFNOGU9OK9PtrdSA6t1I81WEgW0cL1SBr9B30cPzYu4WL6ms8i5i5Z7Tl
4EbBHHowJZ04CfXAD9oPm1+BCqhYSXQEikpJy4DUB3Q8KbRzer9BIsR7WxY7pkl9aZhzTVvYobXO
gAhrjX++PwPITxaxHyp7MJeQdcdP9rjSd/bKUV/CClRnTcFTAFkgJVCldrXgn9vyXko6bz4SAy+R
aC6jrCaP+Ze72qS4OIarU9193d4cvNdJ0oriSOkOBxFnywxmKr9eenmlqcCTHrr+BC4xblwqBCr+
H7Qa9AdYL7hDT1V1Eo5hn2RIO2vQ1KA2jTRUScm9GaGp6lgQahF9bi/kSrEXaBdimysQLlwtBxOJ
Ga9PqMKGKkbhQhdTSDiKCfjcQ883j2xGbsnhUB+U0enhYECsvetTHsaKxgtTmp4ypZnu1rUzf+DU
UMZMzRQv5Ym5tcthgC2ZoIVQAz6vDdnh+TYEWB3LKdn07YbrSmvezJmVFWe7WTmiWTacECQGVowj
3Ale0VKj66+xMGvLOslqd9gTxKODgKDFhOq35NCWTEPJ2II8hNA0PuTiqsCy191Ork4zLWX4V7fl
ifkQn6AWGlq32+7qElzOBSS/nfCI+S+T1P+CP842Zh6rsmwEhI5ONc5wn0M2Y4ew1n5u6WVY/6AI
LRWisAWIUHRJyheJVDyvSWBIaKNf2fnO5NYlKx9SY2yqmSJD95ed8rNGGZW+ESbjYbCyhHibFKL5
wtIkvlmlQKwBgjcek4bLyQuphdWeFJoeN/3HybHK9blOBOb3rIeloemz2Wsv2X4GMCiegCmhqf5v
8wY/CWIqUFLrzloSzWiWFgHI1IBRb3omkGVxoKEjXXDd5nf1LsRBRfDbe+1krILkJ3nl9GUsSksU
n0G0/J5tHNL14vhycmbd8Xlkq/UbkMIzWYe52RoiBh6F/rfBk2aKF33fxGqApy/G5cVi6/hvfAhf
YawPl/pk2btbDJGLbeNn0oPzA8LEmfa3VMAalx3Q5JsXy57WknNVDMNqblh8hzynGN3/oyVaxrV0
fXvK9r78bnzcvJRPrKFjCD/tC/2aBXfB4/znIpPDqk5yZQ27KQKz6UVQygrV7M+elMBwLPlG9AS+
2e6jzF0DByM9VRNOCFrun69xsl2IfB9dlMCDgTA8QjuhWlIAHYuOIr1uS0n+e8UchHOEPvYidT/p
Xz5pebW28a+NXHAp3mCwy16aZPX33h4Mj1MfHh61nfPI5zvg21vEvG/EFpYcdaYfz1NpMWuLE9Wq
lBA9r5t0Uu/RW9+CNa59BC532yApSGshu1F9tz6JxNNp1lnz2R7RablJ5BmeBcMKaPnBP8mRTzDQ
dmhhOJFfV9qiy8q7jU+Fpac1lA0kgicCKvmrNdWQQaul2RTFcRamGkFojKqEjXMcRLJ6XDFZ2wtS
YtUXnE7f0TPIZovLrhprnuBKbh14PUfwmJWpdwsxfBfGGQDKmHvuFzKgSVq7uvwi+49A5UnNkAEJ
WadcoFZZl33nmLS2XCXdiUzcOJFMKHKbcafMz2is5EBhstwsfpy4vfOYU9DZO3xMdyvMrNTKPXCz
ZSIBcxNQIjjmcSmV+/ymhJ18X+CbZVc1PGnh9g9B+J5QyjTUZmqNwooXhzR73LHKcwwjtWXCfLXs
0M77FJRZByEwctZhe6K/cppfP1hLPFVNQtToPbgFCl/tblNxWtizEqLJ612Dza8yT84JMM9f7ihO
4u85Urs2FUusnD1cuOJIfGsvHWpwkadovoJOSo4jvZ4lt81ARPAgrC50Y3Qk109EezNR3FwmO2kW
DA0tFvAK/9pi7V3wt3bDIGHoTvhSo5XKJRh5e6+9UZL2wb9iG0D78NAx9rzWQYrxrqxgcA+cVsqf
k5cMDoogWN5sV5xAhRTMeEpDCKMg6ekn1KHwkCvi4/cr/tMav+bg2B8hQ6QtTAUe7+d8loV8zS4w
oqH+jBJINTd9znlXWQwNrmCZddWbrJuXXmxzehYWs28ZzcNkFrDWdVjCm+xs/4MQ6Uuz6kJdQf+r
zBic39V+/5w+gFCZvoy0EvDI/5xJFhXP6k4hdjHUIib3HJghBwF3yHoJKI+J/HoHTbmb7SPdPvNF
H2zAnCp5VT0q0L2KfKp3FXK7XoTSiH1qqZyWZVUVC0JkNTrzM5ZHSaLYrAE2UJxp2KW2yyEr8AzV
I19aJYtMP1JkDaoAcB+3eXi6AQeWqvV7OhJ0I1z2gXdVLwz7kX/aZ5CCDSqOkyBO23n0e4O/cV+r
zunyrNc0+pOBHOxGh6XYAekhgcbEUm2LHJyfOOsBUWSgwdKARs8QJnUJ2FEclUodtENhNnw3rKXw
wJ0C0onsZ+Y4npNU6a0hB0OVDkNB0vtZdzS/pnBKzWnNGtV7h9P+t8RKnwPOnkh1ygDM5I4WhIBQ
OhXqeBYPTOx0wccwyekG9Fcdd/leFikbYdDs36cVWo4EUxBRK6WWcObd09ItcfXS81auFtKpDIxV
n0Cf7jqrEMnnN0WJ6E7uNvk3gV1ohPM832aYTSStNSt887mtlXl0LIRFG8xEyKnWcIGX7Q+gy8B9
YYqXrRmloMiHjIRg0XC+8h5LrX3aeTiy8ClKarU56lnB3TbjC8i7+slivdxrIxIFwppPIrUBkv2R
7F/Ltve7HF+7Lx0Y4jassnhDRvm43KqM3CvbPeA2bIiW67SEL+7Nb67AqkZDLKnR/3yNVg/4S6ii
+t92xaL4DYm7C2eDMfAClakhuKkE/Y1vDT4Xw9Zxzayi5Ifn5h1gCY1/sSdL7KY3WtZNuBagPwOy
ezViZqdNge+Mg12KilAbcRBKvDgzleTrykYG3Er0FqnDP9p5fMrussciWfSR3IPGJuWPVvPjUm37
RDKwlDkVi8fOSkV/TBRhGJVvuvbkuc4KhJRIqpuZs6QJUhMg8icD6mTYbjGII4vTRLXyjBOC5lB2
MF60Og+0/skShuMSJUNPXvy1Bs5i1dy1LWflNZuddZdr32Mf4LHderappPxWPyonQrayUVUrapUY
grsGvlwxRaY7pc4a1S+VvZm2UAtrEoHAAmmd5tMz2Z19GhiyG1SKMQMRXRIQk8IuX8UlX4L/zR/W
xj2CVDgiFFvtk13thk+v6Co8J136iL4aFdYrh7hq7euY2yTHl8Ru+DBIYQ85ZolrLvum4q7FIWaU
t7abuNTJ0RA4rlIMPAtdE9PScLQpxAXd5GbQuuSsyS1Qwia8hEMmbboTc/qMUPwx5K9LEN69Xaoe
holcQC7bH7Acq6Uk6Qu82KuE7l/Z5oxd220A1YTtBF06eCNTICxPdbXLLBLtPc9zT+eTk2n+fjxh
ge9U1nzLKTsrilla6u88IIfZSyGgHaogoJYj7Mqrk5il+HAFK9ifgDGokY/I2kl9H/NJSDjsBvcq
FwAkENoqCrmkUxQl6yYsoyUR0IpiYfiEy9pDaa+47gRYM+y91ANNNxwTFmrJ7yWgQM8Ok89puqxZ
f+7ERM3Ycr74yZOsjr5f4V9EIccCMiTt84gjmy6pQ99BXkm4pb+FYEA2+cwX+mt1kt8MQ+4QRuvn
cv6vpvZb6NR9aO8tADL74Y5o0P2E27JuIlhaUGs7nV3+ZowVhIuH1Sqb/XB/vtjsN6d0HnZJH2aI
NJiD4ZBYJVLxSk9PQCTP7SWR8OjjeC/AoJysIJ5Z2UAURc/fG8mnJBjZQWcHQlA1ZHIA76fM79mw
ZhObFLaEzdsWw7qQVuWF6z+gHh9h52CmXD4DJNQ0DiAhHUeYThq2G3b7+U/iURfVYQmRRRCW4KVk
QrD2Kn3IkgOfQRmaAzzMIW8tK9kYmIsF9nV4bObNHoXcMzGyT/txeh5Mubgqo22tNIUTUWKvls8r
wBPdCQc7v5xbB0LRtUTsrXVfA/iFLoRIs23nkYAWGXsodR7a72rTWwmObKswWk/TYT0Det7kCBAl
twzVuLy4vOEeS7J01ayuCxSBifV8SRjHAAIVdJSYND6QWUkLywGkXzRq59HOZNTFHpZnplmX7oJz
elRzlA4DD4zEbQlMLZAE7qaH3R/v+RC60Fsx6Zz07o1Or8mzo59MDPz3ao45Eea26BurXiHHAM/X
TCAO+5XcX5Kpcdb9PQ5j92TwmXxxhHx+dUpV92WwGAVfKfBlrgVWr/qf9lu159i5xLdrlbGyYugS
cmni2sPpJ4AD0HoH6QIfZzPLYPB7OCCqFyqsJnOBAPf/Nme7BOqRT+mYs+jz2dvbUoLoidIp8Ocj
nsFQXQ+233htEZOP4MD02BD+lgwIpHabBDxs68tT4NOucrxn4xKYGX5Z59JRDzTuoQXvuzp1Bm4G
nOEnBcwEwwf8+Prh/NBQtboCoIqeTUfnahii8bB8TjrtLgJAso8uFq3sDFLSup3gr5A1h9wcEISc
Mw1rLbcP1Ulfm7LSNda9HESnxTo4C0oYc7o6H3ljb9elbwjeNzv4ocBgXpxC3FsVS0/rtNc13FI+
IxIrdQRwG9qqMovjOl7uEPC28w4Mq+8P/izq4tJinFtd3vCAZ/lipjdDDp7aOID9Ml83xXv7u7U8
MPrYBg91B7OboKkaeoUV1+Kx1w3SjCry0sxUhycTl5qivT9YAZc9gdPP+dgmF2aJVrpScBImMaQU
U0rUEVd/c+nek6ANW+xh6mWBIBK9au9KZf3hB3nJMWKZOdoPvn2KEOw6QvyzysskUb763Y8/feRx
zeWXGmJzBTDWKgQa3bcfIHWWKb1TN6HJCaTka8HRo8fy3IvxVT/kMbG5A7wEY8oLL8lsFbBa1Z0n
1cVWsc/bJHwo2i5GAzXwFqkvUCuUhuFbwLYggTt5Grxqk/FR5FrLr2tv9IzYJw2qim14w9l+PEc0
C/PzC/hvn/UegIso7TOpaG3tnNf4WMR8lOjkgEx+9JZyL8A7CpG+UJIYLCap3i0FWOOG5ooovCGA
RmX3Awd0fT7qqm5/mckx/LI08EQsnqLMNXDROAMWe/WMwsby7zU15tgurbz6cRnar8+vInCxkhoF
ur5K3o95EeQq1vE2ZyKfeQc1b2+ph9rTyps7CB8Ta41g5Xvrmllf0A0a7RS5IMMLqVeG8oe6US6G
tSDPvvZ9SIGTWnbERUaHYgegV9Y1pu15gZOOibKbFsPljpkPQ09K9T3IKRF33tb1x8bATLgROV+Z
atZBmdJv5BOz7GlQlcaDaeJGEudSCfMc3VaYvTKIZdAAsekbKWqtbD80Cx4V2vCHsdXxTN99kAek
DZcSqAKhokHXDQKR1DCjOwP56gZuQYZVR82HOPoDw7Y4MA5Vd2qQGD7DpXAhPNkN512SlUYWr65t
y3/hnmcB+ujdyzA6DEdCI+f9yIJw515G6gs0w8Rav9VqmQlXQ/hLWitl6Ab0lmG55M3/VZK2Zykp
jT3B9GHjZuqqFP6u0uGjARRaZwKiWq6z21HoanL6T2Ww+L9jfnCAIuRV0369GybzFBAjbskS7GGY
+mic8Tjqkig1YcZhOqkcyYB3tuVkoSBl9OH/ENd16VwbSb3iISXLPPqQtdMkfiTOYZO/vZuaJ4Vr
hybyRQ1IQhNKZv2qjZ3tO2+TenlNg1fZZu11E+TPRIi/lteBKmjA4V2MUCuBpB5t1c1mDn446tV6
iBmg+JikDppzcay+YKSsiqBH5njQmaf8tZDMPtjd38lTNrMzgWjRixQ2u8M5myu867FEtDAXelgc
Gtjq5/GeUtBEX5v1OoPJ7xbyQKS13dQRK195xf4RSKy0ROnik58tb1ALRSHhQtomeWrOQ6MchdUg
Hcv2ZnYLUs1tr4x2jtYQ8Blg7RkAa2tcNLpy1AEbAZ2q86xqzuG1j1YqNsGz9XGraHvKZqv4NXyX
ygJrzlR76LFuXwlbQUxAvQzwqt99GsknsfVPaYptlDMK0WRMOxOoxX0wUuqS+Id4asbK187SF7Sy
wur69MyFLsZqq8vpZUyxB8gvdQEV0YH9oQqOUlfJGqW3pq93NLMmvLP9U+k/+hy+no+K+NX/wfIJ
Heyl18qizm4BxbbESnYPS7AsZN3TpQRYwg37IrmuA8W6iD764UY71TA36uj6hhSf+n+eRSoXEkEp
ghLBJUjXk1VUb7ZnV2Y5eOMgOlPclhF/fjDVUh8UaCX5OV6wPTzC3pZHDr0niBPe9zUiX4lh8NNL
ysOrIt7tkABflLBrX46vuqBaZP9lWpd234+1PUtnZKrvnT0hqR0bfFYkHmWYixsSWEjhkGHNSpC3
Jlm0OAhhV+abjmJpXJ4uSXS3due+3ohNrDhmYOwv3rpVsRQb7RfM//LpzxVntJzUzOnd4bTei7Kq
IiPH4/Mn9O0qAd4w0LcwVP3U8naPb6mlPWZ9/spb3aFcWruGsb/P12C3jBc2e8GIchu3q4uo3DOT
4EVQY13bPzht6qwmm5HUKrrppztyKyYxiEFl/eOXQgJ+EuC7OHim8dx64gAmSr6rGHYVXDnc5yYi
Q5WarPs3eTuZ6E2RgWsVAvujjgISd/oKqKqwx9yjB2t5wQbFboU76ttE2F4N8k+h/uorN8ZsPKM/
fpGPJn8ZPjfbkiV82RHmxfMDlRoyKT+GuWu01WNYhRRAy3PsjSCL/WBKN35Q+X3lqYK+LfmYptrL
9LFE5S8BsGismDhyhy3Go3LBte7xojVvcwBEAmLzvJws/zRAsFAmJnLQ6iGzuO0rMLjBIpzWs++E
32liEF1+AzfDogJ/XY1CLuz89AoTH9cIttzBRjdjf4nGUAasp3mTMCPn/qdvS9yFoSV8CvrAsUTN
cdrPWTp2koBCoHVOZereP8eGuLqiHnF95yeCWI1SLYh0clCFNQ9fvaZWBhs5xuqDUq6XMtJDIYgR
1R6H7aXW2nHpEMdwcKitvNzB5c5aCPfYc6oHUHu8x9gyRz0wn6OcGA6rXg/Q+Pab47+MPng3xyu3
9kvCr0vCKqsy4w7vTA0nWr+gKU8YFJqhAR47ncmYkcaTDHUD/nJeTmsrFLynnYB2zqAiOkGbAV1I
y2HVnWU/EKeN43KdOpcuVWwR+ghebmMg+PiqqwqvnqaWsO1TqFuVymv7BUNTGfT6vCC2gk/PxG4u
D5kfyxQAwcxJxkTuf5aybDc/h1+yfVPnDFAoc1prwz26gjY/4/2xyMO+mPBSosGiNZDmrm3t4ZYa
c0AXT2WCqFVh6TwPKqqjkqD64GoV1A04AH0O8bfXvc5OLpl1I6y6iB6izDQCuGzaq7wZ25AAaFuA
tGnGNWSVovcrChogKL618Di4uc9d9Esh1xd6EHm4UrKsIc++4EvTGBjPqeXOQAW5rX0uhWg+qZjy
oNALwNSwhJ1nZGeCvmFaLcWON0YpPQe3VRgJgOXNxMyXTcaFOMo+HVOZnEVIkP0k4ST9aRid3w4x
6OxflA8HgLUqWGVgIU+Ws/5WeI8O9V/ApGrXNyzFZ+dt4NLz5Iq3/w4Nvobx0WAi4d3lftxTaibQ
a5xqycLQAg9W7ftAu/9/PPF3aWPgZIH2DdbP39qF7SoP3F0z3RVxdsFdZWdkOrAmZZofpCBvUxfV
fLVazjf1JLkt3hMH4hmnsnwoyfa0/iauvxlfx2kkC3mscI5iDm/WGlyXdjmEpjTGC+k8JaEhA+UQ
zIIugcNW7RqnO3v90OnHMg6hIrUNLk/SBl0fx2HlTBASOpIqeOY733BHlTOsXGIh+PvYOduO4YBh
odNPNgOqCsOBsZEC5sA8xglrgcXbmQErqHHwMzcN1aA5+LEksO8uNT9aSkc59KHJHlr0q/mIeXas
r6VbuhFuoKUq6QYfYVKZk3g+WUWuvbJMYwr9ZOAblqGFXFsiMqt5uL1GOZ6ZR8yOmiD0Vv1qr0rC
sdFYRcKE0dJJYyViP8FSiimBRlPkJ7MUcfIZ9u+eGERr0ze+YmK8noJibU67l/QX3V9XoJM3T6rn
wKJ7+g8Mo6gOBSQlUFx8+VlWmNLjbP0bUEDZn3VHsvTYmOQslKvzEKJml6vdUlpTPFWuKxDRV+L2
Z/T2enxLEA1mUIjWDKvDk+I5Sb5yLt2qYUmEAgS/PKuhjPBOCdsO2C4huzjKKK0Q/jvwT//gn4Lr
FAsUvUbXNyAhqh7AFsm94U1o/aIKO766M9DPdddYb5pKFyMU3MDHx/NgD82omc0pVrlETUCE+h8L
yyhDhoENoecj8E5FvHCiO4N0OAUsfPe52YZGeigRnsqwRYiJ1Xloi9eRaBEOcxS+Z6a8qVgmD0ie
+TrPZllHwS2jd8FIeERmp1X3JtUiFwepv9lqJU+d7zMG0bjqxa0SW4zDeYfqph7EDe5qN0/GuxIT
FniDMnMN/AyDRdRCTOTy8NJuQEAqQnuIWPz/DZF486YdxfovpGC9g1Sf2JM82L0S9C5BGqUf8n2C
kHXOm5RTo3ZUiL34hj1nTs4RO44vzOg8lwG2AmGo9keKtYk+a1hweFsfXdfQ2Qteepdzzfx/gbH0
Sz1EZ6sXDv07M5lOSYFn+OpXq+Zh3UEEZlDtHOFeDqT52E8ri31pBQDKpukcjRURf5bLdnwmSwoP
1WTl/pg+Nh16qq3xsM1PDLgNHbw4JN4IL20uPPtk0cgbBm24YsDnEzAY7JgP/hPwMahD47jhKu8I
5CY/HfdSLb+8Ii8jNvSMAXc7zl8MVz4p+vdYv8KJHmcEe3sAQz7OVinTME9BlSi+asMDks8n+O4R
Zu8Tv0QAxKClp8PgmJDeL9s3DWg4xvEfyETTXgYk9sl1NVwifcONC7HO+qLTEuMJsIhdpUq7glGm
5XfVLZV2dQm/Dm2VJIjeGOYizx42XuNjJSfliWx9+K89lDEM4pOaH0sLr+k/dAS9x6PXlIT3OBEJ
pJ57us5WDXLzIg3oL43E3WmmVUc58GXZDpzoMC4XGRtmVloKpQJj9/hMeUOh1LiDaNbxNwBTfRTK
XKhMssHNOvnRg/+W3AR9HhOTOSa3qXeFF5pffCCHDf06Q5BN2Tpv4JBviZP+nw35a6V9JjRMDuZw
qi3R720enJMLfzfm8QVeG1s9AJcWIK4veddVRI/cL3Er3uO1WVdnxZmOrOkyAS/xUcKh+wPjCJ7q
ryFqOUNpCjjm4iEjOkOFZl6WvOUqQfvyOaVSOLOf7U4i0xYiKHZ0PTV/x3fUZDKxgk49y54vXeNa
XUmy5aLzEWjvRuiTNgT/Wqh0qcMZXm8UeoG0VdGy/h3pf3E5ydOBf+bzpyYNWIR7htuyEf2emnSo
fxxrZRUxnKdZ9VB4G7ceLMaxFVsIazUmh1fkWTfjuOA2/TtuPmhRzH1G/W79XC2eLVz8JHVWUyrD
58Smv9977Lk8+Ko/KpPuWayRaQ2X0wLvC9q7a5OD3rl/5Xp5eURRUyNLmrbqW0U/Opu1rP4ye72K
DQEA+cetzXxCzJ33/Y21sqfmosDs7E5MNJxkxObxIMNuzBQ/eAEpehXSWZwwO+trtIPodAHA9YF6
eLg4NszmSEWyzk4Q5OIbDIep/2ceX+PKy9FrizXh7ZJdhqWUFhXTkOA4x3xsYmoKZKrDUZbZWVBr
+U4nMJ+nDK4PwmRJmMFu68I6haN8DvvYMHa94Jv5f7EDO90mhvV2u58/DId/nSAFweK19aMnJj9K
6fT4xyiUeX27nz/YUKMPbPJV5EXqxLXxolQmdIBVKEtQ8XCAqeHvBtNg6ftkHRY+1GaQQMM4qiOS
58Fd9dFtBXPifKasgljQifLVZl415ZnUxXCyrT0TXA+AIqrl5aYLtryHQCzajTnEbDx0PO0wT59z
Y8wZlEXYWQW/d8dwVbLOHcBenH2rvKJh7zRYGHMFbwiDpfLu1q9dCosnPm+cosBRmQ8lc6BzONUD
17WUS2mXbqmh0djNFIpS4GqKCPuX+qbE+j4QuLC1AUJ3x11V0803JSXTQXqpoN8bJz51gyhcz8Fx
50K+tEiP3KdBwu12nTh5XKCtnN/5VCBR3UdoYLCwHxNDiakDq7dsPQlxRx/mXkRnmCR5dTjjGpSL
lzlfmaSUBHsJCMUJGyjqCFGrP4Mz0e9Xh24mx6cxUumcLxiMAbuCZi1mvyM1k6vOYAQjm956XuS2
tFFIlgVMAnSLClJi02cslmCEGqwKgHERr2GL2QH4R5cX+fN+0P1QRM3Sx4nl8lnpwcPKHMSon0ce
0WsgNoK69V6z6OAIscpRf/7eY5uzDrIKYP+iOebWco1cpZxqc7uyBLZHg6k3/VP8FOho7lezLLkw
XX3dbW1gcbP9eXdQPrXhNiOy+CGH31c/plbwSKnpUWHR3Le+x3VNO3pxDIETsUjy0/g5F0P+cCoj
3VnNU2v9xmh52/B9vQg8jnldnnaCMIc8bsiZqwWwrZkX0m055zWgUGgqafsO8dfgLNQio2gRgThv
HsnizaHpt/Z149aFZ+kVELZ4s9xvt7VWdccLtpsqa7PZY7Ewi2V20XEQv1Wk9dpWJa/R7NhcEUoD
8qatQv5dFniLXl3HHjr2utv6bd1x3NvK3D+eHaqlpvkx9ZwJArFrWVe28VTGyGcZ0lMlI3GP3ixY
3pkpuuktfWIrtjYSfLNo7xJjQ1B4isgCdtGImi5LokERmyH8W5BxuYe9oXmwGOBA2C4hsyvzuk24
OSZXHXvWWZuPbkiaUd6JsrED0KZu7OIabaVpJeqc55BEN/dy5wObf4KlTXDZMVpkug8UkPcxuj76
SyZDsZhWkll6/YOhpwFKFxVoHANZWGTLsIkC5vV8XH5r0MgYA6i5SP55gcMPkYsF2yEpi6zXK3Eg
MRPch5+ORhlLww4SQpMDqbeXGNCBHyThf2oZTwn2L9NhMq0ew1o06gNN4v7Umcm/xT+B9GwrmSGr
HraDWQNJ+BMmsOw79ShXAqHf0EhZbEvfEFmRGTk/H3Xq5B47LrqxGSA5wb1xfquGHplCSNbT8H5z
A1PLLaKu9BaonWpnVErzPI7hezYQgK5N5tILYATBeZrDxRx5DhWtvLdlJmafwJICwRBLGb9WvQUB
2+I1um4x8z/GX7v82vRvPj8wL2ROzDF07j2VA4lhWdQmb2ESINAIuAUl0DMhcbMdPd3gwiF2Qc93
Z86nVK5pjhArfVSY50zEGoKPyyBTpQ0jJ0JOf0NOGNRb9paSGD4IXN9Ek6rdS6UIwLvhv/+u2VYu
lZ30TOaTmECszimTRZvZeLJo2tQ6urxcdRiWLV4liWOKLwrEm/VvTdPCOmwC4VltBU4PVzOMAo76
l1743VzFebsbYJmeUyZGBmtmD/ds2YOLOKMooCSjfLo56lBB2YnPj8pRIFuRi6Ps4Y48tuRoO0Bk
53diBlqKGjOngVrRgCYjYj3IceLsLd0TAxqPn/UtknTWU5MfJIgSaR0oCS/UZSykQVxD9PVvP2/f
JBOFTso4+YGDyFnuqP/bip0GEofmq81VdQchmuAC30E0jd71lF8IlOuLg4tKtSBCU230//ZtGl9j
TmgZ9FTlpB90b4aGOtIhRrK47iZRrXa6kOTkkC4Gpz+ZUjKUsuL7j1hh5cCq7K0yYyRWDJxkxR10
YZDJQ6FTZQ1CqKWUdEVDAvIekxjPHqNcfWSTfSE+w4TZ52pF4Z9qj98GQoP1HqfYq9yerquEM18g
juRm6VnmSRoRdk5fHMVi6C+P0+CG5xX2cyI+0DImtbxSceEq9XERDN1GliZoa88ffLQK2T2Sb9hf
TVe/cFLhsCcxxHOS5hNSTXdXRArNG0sSGOk2Kwumpb5zAWKDcvTelFkmdoICdtQ0KGVeVuruWgUx
r1fb4ojMh/Js09QpPtOUCrj6TAvdzhnDgV9J7lCwcYCJCkGdj34IZSeOI8QuWfZWEWH8NZuG/eMG
gcJteD+HKUrtBUr8wt66yrXtUGwTd12Ey3IEHaMdbaA9d4R/suV8baTdU7TKUZIlp7jKr3SfF75X
78QR2PtWZyXMXJ9RxfT74nxXc+p4SH4CsmHgDqb5e3KnxfpOFXeZuZ7mEro0JKJUxWwUpgItnFPL
f3+vaI3eqDcn8nSdvgnSWWKjI/2g5iLChkaS0O94xXqs4dnuhLn8VCrs0JLvYscWg6JUATwXAfKJ
hFY8aIsen04Xjnobro0mSBSPNbsYx/v+LFoRNzPC2Uk/pQGD0aN5OuGmYUE+GralCluD1hpZvNC2
FmdP1RwpJMqJTEg7qj3CGHQ/Dgu3jwW6M5ricJL8ija4rDYHljSn1O1zGc4fkecJu0mLb5OzVKKp
s4qj5NLKCeZTpv4Iiz6ANYGRBe8tOBk8EWSFgOT3JSF0jgyrVSVLKAO/Hd6yzEAfgPtQ0weyVnjn
hue1K9daAfHMJihdDxyFwFAhHE0irW4+3J6bdi//DB07HNgzbrCYXyL7YZm1gJjlhTHVG4hYD3gk
aiE1m0SfPOxef/CYTiVX3ZtaeKoePKb6YwCc1V2teC7C6Sr2BUk+JO9DgKl1jh2uOWnv6fyNhZJr
NtTJuiY5JfZZlxNgZqg4LScLRPf6gVpnka/fJHjo10GLTVTrbKMsdVG0xaYuw/5SptcQ7UD5Mn7O
qaKi5fqKscIdKOnqRkuh5XPIrPuPsLgcKedtFpUJf5TV/0gC87Plab4G+bM3QOHike234bvqV6rT
eMuwfF7RzbqGYDu+duGmiJ99BT6XIKSAPb6KiNNmxFGr45+g/ZNUmXHY0faqJKu9O/+S7Cl4JoDz
1jeWVc/LIKZ3KARHt3bKAWofl1FcrsDCZckXmhIYRoipyo9HZZW6y9IFceAWqIrxgks4EC81UmEN
tSEH9WHLYh8JvqACOUOySS/oPP1SicQe2uf95WzQSj2ySm4L2QHVWu5dY4ig5PkDayT9uWhZnPDS
YHCz1ZVicgzHr8BF7OfCA/oIeTeV5zt95ApNLtK1CG+zOLifgh+E2KwCdQhFtJ2S5HL9YM1IKEVx
yMeEM8GxHuSmr+K7Rb2wJZXvx/2Za9olZni69/S6cm29V7iDMIMYsBy05O2K5si+0YuDkV1gUWWh
CVmjTyfcvouxjkvBqciecxgN0WqX+N1D55oU8gXFt2Lqm5JtL9Tv4EBbVvN91Zsz/0v5K00NNGKq
SSepyOcn+MGSpJzo1l6gz8thXw5w6SCkZObg9fnLknyh2G2giJugAWrtoVV+tpS0s6dOUFeKjbew
PfXrOupJ+mkO85RH2PlbjlilgjlVPzJ2L1EoIdAgyCj0F2RFQNoQ0+rl/PRpFjOzGXRruwGOgr3s
Y1mfnKutit5zlyZHv6SJaNB/AcPjc7/auyDGTT8NzmXv5NEGt/Ztv/8XovovzuXr7EaXd7o1ikLz
3JosknssC3pJwtX7MaE6cISYOjIAa5ezChC/xPr2NAmUPb0Ors3+Dra/Yr3wo4eLK9R/HtpVj18e
UFpHqwyfkMDQzA3WoycUviSm9LUJLLj7IEKe7rlA8ni+PjtUOR7ncb9yO5++LthiQvynB/PiBjDJ
K6QHqrZtYmAZa+RLwFpFR8kYOtcLjGVP5VsyuqSK3q0x4W/xxNIaWH5kIhBfuSzQjoekz3iTmSMk
fQcuCus6NZAUjTXRJ4VOQ94YO0yMBUxHK2QE/AFlaWuAKHKf5wqqY3q0P/3/i2J4FE5fgBxxQbJO
skDdMUEAbOhZALBNigdYlYr7JxM5dX4wouwaI15zVkwM4Z4irI7w9JhNHf49G0JL6BpUBEkCa7fj
8/J9m1jPHVf/PtEgFqpcFXyBKU6gp8MTAxqCSLbe4XpVefn4OBm+AnGpv67k66M46gD7MzvP2FLv
+KcmBsLnFDAXRJUAtJWAWGyeO08nIkCtc3msnFvj7UV6MqWAi8EgdEyxrkiYBmIgxVfq3tuZnRmn
v6wjFiPMs9pvzqmnZ1Twq5nIV4onpw+XaWlctBh3rbwU2ntas9Y1y+AWunoM2gZwYCirx2VIXJNM
o5tO2WMbWrJvtaSDKStmblC7aa26Whpiw6a+0WB/RV3nQgBt79AvDby3T5pHDmaFCJW7CB3ccZri
lZbdoneZEiTq++rukx9mgsS0QhmB43JW52RojcW77qlenU7SYn0ylY3L/cCNGL+98e4+4mrV3wmE
chF9oDMEUr9F49n6qRTpJd9hnXiQCyoUdMH9S2407lb47q3kq04WALRpiAFL+cOA+4TJctq+YALi
mC7NmU0+075bS/NCgH+9MNid+qf6jCGherMGyCVgfMh/orNIo0hJ50KgacYS4sLPz410EEhYbo/C
qDSfArsAB+d4W74fawtbFU+YOVU7naeZjlkZC+M9yWCwATKg3CSbI2Ifac95SnjVe9Ljl49ANeJD
gmoW6xDYDerdGsF8mD1Ge+6tHvhsGFG5U2Ru+HXV9C9sN6xE4btLGmlKYbyJcvJrJ805EzMEfnaz
V4TG9wB+xRPfyTOiekO1/q9dAXyoxOeFfYvHuTOaA+oPzFfaMm+Ul9c9du54urBv10vbPsBTif5n
zhs/g+tiCDozHduSviyw3urqqnj/VMxr/GEPVSjlpLVoQ18uy/NMyriAAv3c2pwQMPsXhj/B9Sn7
nKI+indHhzxNwjKNpm8fK/BGJEfdDsMOjX8YUVtiyluq6tIVERRxlZdnjGGhcQ2MYxCOG/zGFlJG
Va/ydx1lTqNlkHDHoWoDIh45rIWckTq3JUE/H+zKY/FcfKMbWue2FevXg1evOzx+tLg8w+Ey+Y77
ImUUQOcL1NdVSoFEJhJ9P8p3R5lFJXBIk4WZL01W3vY5n1QzufnPfy63zwBiXmBLYB/a8hl5wzpo
Wqqtjm8wpqh64FKsUI/DMcjiBkYrvHvHad48/oElwZEtGJ+XwwraPGriKELqzjGMfPjltg5u0WQQ
Yv7SasVJfK7tn0wg9pAHPiJeHq7bZlbbZiyxz2yu+HIhU9NpmNOjXUwJvxKkyNt9CYG8t2A2PaL6
3GvFgiOxeuUj3If+IgqZLgXScJ+on3+n+jXYAyIZAXtRmUo9s0Hd4wyqOgKvfQSbDUgTHMfOwVqs
I7AF9i73elTQG6W+ClXccPa/aJwm19yXwiKElTZxh7fT8oEJs6wYSC7m6DHlMV2fqJz5AjFn7gfP
buTKLcXCF7bLBX+AF7p2LlZ/YNvHtWCRrpQlWxYQqEqNRO0hc9yuq9FIO5w4rmdxssYFfQHNyKT+
z76RPRzx83JsI2JHMDYYqwqIWdVyuUJxGkwc4gkl/qeuJO0XnOBAzDASfAFAEZnedv0R+7VFUi2A
+k8fQV6aoklA2NIxFbzzmMEKZt7074rdQGjVS7IKw7wT21Lo8H2NRNO8pTlQXE4tblAxqOmFbVjt
cJn1hNQqxPYXJdsUvv+kahkn4eqsLxeBgwAxNdLdOcQe64UnO5i4nL24XKVpH88aBkHEtrGLS6jm
gFdMjyFcByga8LdqdEld8eVInV2DxCDRfvP3p9SfjgZEP/QAddf/3nM1VxEj9gygSmgYkOIcFtvy
EdEx9nf+vIxspMmtjqOsUJMSrUgSfL6SAXP8WB4eV4hXLannHnrz0bFlSO/3TwBURtARxGDQ+ReO
qiC+dblKkxODjOd8wwUlJOnxxcelFyFdaSKgstPbtrrmKC6BWD3L4lel3o0ix/atL4MMSyvdUOIk
sl8sAwuRns2GcKjCJe60GOFOcGU47062Fh/iOiDrTGAJuX6o4l8Knn/QAQ6Y6dXzcK5V7H8iMDmO
VGZtlUS0ZhoxtJd7RZFxCJnlzgmH4ras/f37bBlWHDBUoUVDUKCCMmJoQ4kzAC7nKMgQfpcrGab/
vVnItsCNa0WegK3978eZqmAYbu1P+E8jWC1BdgSbXsx4zaPe9Bay6CG+64vITOUvsCE6aXHu8nxD
5iePSfRqq2uox4o7xwaxug5XRsTNwkDGhh17XLhKogVHW7PL25fFtgHGsy4crgF1xYuD+yIftW3s
IC59qoLkn9TQUnhbrRX9J4jOJf2bZ0/qfIWz5ZjHuAADEWpX1mZ5b7SXq8QCyDZkk8NgghfGWcO0
W2kuQBq8MZFTg9+zrGUbgGmcJsNoN4iqSbK+8M8JNBFq9J35LvqayCPjaawSAeavqTcYAuXiMsaC
CI837Qm1OjgZolpmRkyDFzxL4/BG+SEUkhisic0g1EPxBnrvaH7OyylQAY2r0tkXE7VXEJTA28eZ
6gxXslJtgW0eBcL2hs7eRNK+lylSWWmIMbEUBgbHimJEzQrjY9ATJX+GJawg59w+2ZvJEqXNWRle
JJsir6YM4168aqr4D0Giq7apYtZ7u/jA/a0ZAU121FHZbjTcvqkj22Udaga8d3hCEjPflD28bMid
geCn1ZjXDQ6/5I9h7vIvedsUCHYiORqBqVTt+rnM2liMQYb+Kp1x6aa20XSJm3twvmAy9IZQ3aMY
+xjzm4949IvDjDVTHN3keW07aG2viLDDtq2HRN/p7hYiXp8nQFyjuQo6MolNMESkPGSK9rfR0Y4n
bmeCwSuE3SVEm+Jk7An9ZaCBbtGuAMUBt9hi5arb01KVn6DItp2smXzQrOvfMzl09jcnhO+aw96y
A3jSjXYkFCnADdPnKBYDYDlvaJblAYRtA9xzsf1ZaNPEWDfPJRw15Blg/+9ae9ShUaZQ1dR4fAo8
hDx3X2zStgKJytGScdkKvSq/f/kvUR9UwBbprDL3O3F/x7I6rzZrKo5w2NWxztsCYjqJPJJbnx/l
UL7BSI4lE/2YvewubjZiR5mpjl8QPcKhLQLRYWTkyvDjtXmST4ntjH8S3CJihxJUv9l+CkJTYNgg
VD2ue7j0lR90JdSrcCDzL6cBnB3/FgDniu4IxtPONaqDjG2Y/9PoA0rlLwSg3aPGDJINCOKjpCsc
fMk3zqSTAbTXXLaisRy/WQB4NGSeGHouBdhTor+Jme1Pp9yAb1a1dfGa73iZTej++e7bmdEGOrDj
5tBVRXRWs1V5PH3G22PzOLj/HbFiw6+c6nIyAnMEhCReTWOn+iXC9HabHPBmPFqcF0/qai8Sd3Ht
ho/5JV0dAOkorcMi03bBpp1slMe47xcpUCPHZjA0ib24ut+iAucnE7h1U+YupFGhEIdpECoYg1RP
f5XS3Gjc85XogYDalFl+++EYOCeajNwfOzr4OeepPirs2r4O5W1hQ6NfGP2o2WDgCe9k9hcz+F0s
IFVUBuKw3VXSt7vpH+dN7i5NWxwpLudQrUkUbp5sgf9FEbWeF9WDLWHnLJHp6dUzl7+NlW9lBQmX
Qhpup8nsxZKoKxThoQh7ZjhBldfk1eWvfJbV2dxPtljKC1Kgg5F45d/o/QKKun3FF3gGBMC/e2Uv
Ogj7MTa8swglv9A15fDy1ciRFlBPoqe50cQzhvvca/mqydeF6GpfR0QzE1Fb7kRIqRTOf7jvIFct
uMIe8ysBxN2aCS3wBuXi/isYgAKscFoD4J2XZEi5GlWGKri7FFeqPSz9JmqNeSvcv3SSe7owyp6V
muC7AyreOcgZrqYm/sv3BPq51OHwwblw1iPMqG07+rismz7cgTyrtmr6i1xYRP8RouPC48Gm0pu2
vIKPV0T+er7tmzjLBlQEcXOWvr59C6X2WHaRh3571FefvFyYTSzSDuKJ5UDE7U7zm3TSsIgvqLrX
DlyI780qGTts4RZ1JOv67gXpEr2IPS+7qRO3fkZ9s1vai9fSOIGRDtyOyvSpDlC+aSsQkhEf2ucK
3XUcv33H7bl5xoeub+AN720KZDUG2Yzhwr7+erwwbQ7nYghiaW3rBfiGzVo5UlqKeA88sTKiKHWh
14VURsmX0R2A/va8T6mnEJSJsHUJQdGnhSKnlzR2aHlzwOtNN0RiCIFiM4NykAiobtHqwkKz0iM6
wgGOD4PJcALLr2rHfCkAmAmcult9o0nhFrGwGvorsInPaBz3MaNILOmLRP45UIHR9MnVQUa3Bdpe
/xcfRM/38N+kh5rS+yZZXjNAjzFGFg9jvlBoqEPcFl2NDklb/5pbSg+1PSOXfhYR+KAX1CAFxmFf
trAna0t94Mm97c/6qglxK4OVdUvuPi+37pX8laDTlF35hoZKM6HEMymZ8YYvgsfL0UDi/KJFcv4O
k6vqDD2SEyN3c//y/f58SkHSMbhiY/BIHx9nCgqIMxCIFrd26t1b8ZwWETNIly5ZaC9J2R2jNeGM
QPwBwFTi0WHMr4zVJePKFGRItxnwxT4DavCC0ojaUf/3zaaNuUryP9XuJILlXq9j6TAkNzxyyzcg
RzfXP9fnvAYKzL31OaYD6/cxf96A5FAJgfBfpr1QXhOFggl1WxbSiigtqZ9vqNB3Kv0daGIfHZ1B
wJCv9KEat+b8oyADOIJcIm+NombvLYpEPsniFRJZE31Fyb2Zdp0Bc4kAtyJaM7YLgApTlWGbCRZT
jFw77Ee6zpzDQzo2mKQr/Lm021ynj/4xeiefQvqWsZ811k+b/81ziJKFgtnt2B6rEOqF+xLLQOns
Q7Apo8q0zNe+pwuaOSliWsBXPbsufmvEjLkGjGS4WI6sBlrm0ukxmAbyi/uUP0M50v5NAh8B87hK
ldBWc5gkEUkpm8DaZhhKGATMBHPVYZtTUU/BsIHjpf3WmN2wsAyJN7rFljDuobZSk0OqrndhiV0o
8RTPAPEFmwQrGBDr9FS4nDv8r2FNtayaOeaL9Rfu3b+/1WjjK67QbJqQVhJEGETEU8KAYl2L5bvh
CexbxxhyutBVP8lVeNm+RxosYYvsV+Cz6Mbela+aRN/ZViqLRVSlMXXeGuqsgDJlNWg7DG+2NwiI
0u5hCk9oOjbHegLIymOvbMR6DXEW7g/oR7tHQoRWqVEPkG+7K8uRjv3CmfWoWbKYXIBbNuy/YdCJ
RgrmjmD6DSTi1ES/KvlK4mQfjryPoo/YAC15nf9xVoqgVGGPiCJBUr0gPWv4JO1Fbh8WcsMcUZ7F
P1f3YTJ+IAlEVtSUFW1Ea4QLOzQIuWdFzqfqLIobKqMaLFV12F+sCH3XOIQVfMzYs4f6Z55rfKHa
xoFsivIkjAmKD0C8smfhuq9kgG1dgvSiKBnJtSQ7mkA5BPs4DzbdkrxNPUMQleIu6aWvzZLxglnf
1qbRtvsuRdThOx76lPbJChxkMFSSM6ia4usjdKZ5NPQvLqjDRlh2mRhtcgszqrSNDU5F4VXcA7Mj
yNZ093kM5nrnMn3RWtzj7efKY0ViM/FRgoG0pFvhImu54sCNlOkEzCHtEh8ExjiD/bj+RODrtEP5
KciZREGZ2BkYlbeRg6sA6vFDT52AIV8yqLM0gGQM522GRHZ4C/U8x2DeFGPyN3rbVYRSAYgG7kVB
F+rO2oJWQb9sVK/HQuF4vbD90ffD8AbMNhwGLyMj/I1gE14kg8ZDGpgZFSoejWYaeEZA/zS3fmPH
DsG2n0iac+Oc2x7tRlnMxlqaj3VaEq5v2y/toFjxVxOqYbttFS4TngZ9+tOR/7RS3/j1ksLrNlEE
wOQGMXS07/iEVElIwKRacY7ZxOQAYEhpO2M1BADNfT4x9gXNcaOT7lGGL90uzADI3AhSR9gXze3c
i4s5CsxySz7Jg1sojReSf6KGsFvFbAh6UHf5ELtdocH0QwZpnGXTq5Z3iRghmtNc+zKTYvKRpZGt
UQSuSHvCj92S49mP7wvvMnanmtev40sDmcINRQAsZWF2fENyV0zKr0wtb6vOujYHNjr454HNASRW
qO7veGl+mEazuy5cAPwRNY0us1eK1Jt9z6Nq9BYgmv2xmf5zD9bUlPLaY2+BfvP3Yakd+5jS8JO2
lnE0vFhOJWWE6MJBrev4msgAvij1LWV3dZfeR7Xapv+RlxGWRmWUmKvcH5mfGRdapx7dQ4lYr4Ih
JaF1pEFezH50WTL+8sP7/EjqQnjTwD0WS952sEYRbpjQuFC3+vd+pW90a+tZbLZs9N1guyH+IN7W
8/XxYs8kVeoF1wzZxf9/RyqM/xvYctDHv1F8HSE7ORdy7TRFcG2GCZ7KWUA+EW8VH6fgtEWBPZFL
x6LX7Zr5NHHfnRn02jXFoRniWApfkriM5SjVCeyp/7v0aZmJ7UBDNZDSIzZpM7TOxirOp/Ht++5c
IzRcfK0B28oRfnN53Rz6LDtn6Ax5v48xnu8i6BflP8CsXv7B6GKcLRW1Qg1GjnBQELnYSPlNgNcg
tYAJC2t7+uKQrDYEl5I2c3cDiYNoDQiIFqVfaKqgU7O3HJ/Qh9eo7B6E76eT1/MH70xY/IizuuwR
QNPuwPKoO3eV+gdmshDKIt/bYXUH0X2+ZAHh7xle18BXD/+saG1TbwOm28VBTxCmrzSB25/1KFq+
MX74hmmIHoxWYxnCW3Cy68idq2WO7HS/5bR4Wl6aSyHKydkDpXjnNIMwy+CfydNGsCCxONdGSJBj
DIoRxki7cIb0JvvoI/E68aFXEeDtC0eWQC7A/tyu1cuqXZHseGYgr0wcsimo5PlcjOq7MFX4IG+7
/QIJeXJEzucUdl1gVgCMZ9e4DAxnEperbwmIPDWGaSIEkvbYSySCrPsacUVhtLhlYw9/eWca6MTd
hvomXFqrNEPOw5inGlXcq7ThSA1eYPx0aU3w2K4I029IZ0KXQfOl2a2PfPiOgzhNwcqswzeSwYfZ
WNkZRoNWSU5dQ7M73iBW/aBIEBAMlBmyQszJL7QjnVtop/JQVDKhfQysfWyMa2bgGifvEq4rbMKu
JakO3GRKsPasw3B0QxT8DE8hdXKA5PLSxp3gXQxR18pZ9+F8sHVy6mT+l8FZuF3k01W/PnHikADz
JH2hkvifc5cpdKmqMw4adb8py3oAstiDyrbFp4kpGqgP4uWN97jkSE+vfDJqVZiUiglX9snvtowv
GEZKH2GY4P4jtGQ6XEtmVdks5RJKvr6wJ6cb5bm5yqIei+7rFbo/DYdcba7CgsWJ66i/+gI2euvo
fOlcAkaXNxlzcxUu3O7swhCSVlgkhmyorxZAfwA4KspDJUpv1jOgy/aH/VJuIVvcjOBgGVT7js5c
7yJXZugEFsOLh38XlJ2e3JuDXV8HFGwHx11Wv2DWN9aU72/y0BJVOTxiwkVk1iNp0OJdMSnx2Vut
X5m4TwB4CLMisnK0UnWXPxeIxepbVp7TDp42I3ZkwnJig3bdAJloAj9/DAM3V9raWHiv1gr2aKvl
yIGRwVikbeBoag5/O7vAifR4+WblIoNfDYncxBT9dtSZz25c2IHzISY/qABVn5+b7sVLmXrSxdgH
MDveaVUfKKcOWLo19lRMo7YBWc8URvAem+y/ihgEWUuPZzOsq0LLs3Z6OdYefSd3yvsXlzKxpRdz
LKjaOk31Hp62++MxwW+j7qUmx+j8jgsoPDhq708nz3HecWdEkhuKJp5hrjwLv35OUkF1b4h9sY0R
QvPJ1M1sSlFKVuSxv3qSAPpMmQcxIPcd+r9cwUyOoyAb0P9lCAz2ifg2ilkdai3twUizcFfiGzBK
nSZZm5Kv/gjhMfnXOyAm03ITAC1OfleZkKGsf1d2plqEK2WXoilZrCAJBUG4xjy3C0oo4SvueEEm
cBdOyXbQYla4aja30AHCJcq/Z82jVbQdbItYO1W+KNHFOu+dgfm5JYxQoYjKTaHG8V1ycj9phNeB
ge7K5p7a9Z1gRklyuM02PT3rvHUVPIql+K0V2finOwse/w0WjNpKysMAIPIbt3LB25WPfkMbXwAS
5JKcHMex+eA49CK1VU/MEOGgdU5npP627ujF4filhqM4njZDwYdIGSuRhcRrDkyZXu4RgCgnrtL6
T7yIzFA45ihAVPR/0Vt5lnkMI461+5Am9qq9khVZJXJrKbPELaUk2ZS+Ek5g6R4wCaBeFkhSPSph
p60HyzglyifBbLdDoDfv05LwOHYw7EAslUntIIq603XcHtXCGi5EXOBuE3axWbfdBPY4cmigRzl5
4HpCuTeG9P5MxHyvY2GDh+NZqiwRHOJTI0ids3YmkJAC5XukeFwLoNcEa9QaXpqlYycL3GeSk/cX
Tpd73/SGgK05ML8CkKUdtMK+cS0Vp9hjw0RIVEjq232PufpjRTSVCf4fiouABSrpbQ9iZPIU1bP2
FrFxe76O9r/9U0mZ1C9NBNgmF45frfjjS5twyNjgyTtXuSXXxVkBmVV7zKL1EvipsAbDTBjqxsaD
4D9M2Dc0rrnltjXmc7qdtmoFDcqfTzIxRjoOaRQ4yaTrY/JiVQwvf1w88ZcsDN5Yk9YVo2AXPt8Y
YeGK1KJ7+bkhZV9ZsmKrwXarJm3krArd+oUZiE9iWIXU1boMlC07PxPITU43L9lw7k8jsnJTwz3j
29j+727XddivU/a7Q21aR3tIAt7iBqiC6NVHlnBZDSmnthr711acYuMHyFKlgy6o0JsXdZrJp/l4
18quXzRgs4jjYuuq681A0qNZQdBOExhIJdyPIU+vFH7u3nGSzTDV6TgBTZ+/OjH6GmXg+QTBKiMA
Pz3W9sYZZql7QPfN+Wsj8ZhcF+d8G3PsrgsKgkyUBNsrJiT7kPdYnsG2yhGliH8KbxkItdb4xkHQ
3VE+yCoPVKjm4SyP2nhLG7ihzeRGtGh26GoXpzrVm/YwQDa5sjjLu0AwkRTyPJk0sKSOrNtwdxCG
IQfGktFOy4oFpzrOCDx7KxER8LaJWMRNQgSr4gPREc39/Rs8KfgtB/+BBYXb1LpVl0K9CdQs0n8S
YYObYMzAPAI0owsDYTUmFk9u2uabxPZKVhLXLfak4zPsqNdy+5qu7Kdrpmrw3APhpmRS4Qzg2E/R
5O6HuyBuRev5MXklRA63G8nEkdB02D/0MXZhp3gTPInoU/akf+q1FE1NNhBsVxa6ni5hPoe6qG03
OvI6aykskx8Oskx+nOYZ/SpW9ls4XJvBSZZkJ1w8xo2WmYhx/HToAQFAw0sQIT2hCmRinLRXCmkN
8zorNpq+s0PL6F+QokPXyFxyQ6w+DXpNqApyojqmfbtX/eSMKw9K18QqdPntlui/BoM87V4geJ6A
s/+LhhbkGjSuxHhc20q8W7A1WhdLWuCZsHj6T46FRD7ydBCU2takmf48OzoPhgyWB8sAxfX30yJi
YHbT3DKdpV61hrn0d24hwhxWjfAB+bFTAZmFwgEtlDDfhdP519X0fGuvsTEH88cctUiR08dRkbDc
I0s5xzr4fXBJF7jMQxHR0CCfedKBniXnq7NV6/oKjwdCKoFNS9mnTcUjSqu+0okcADJ4DiQ+aGil
pIovFc0RlqXucWRtGYKLmABpV5n0lVQ2961zeGFcqtyIAERag2YV/KfO8lNA0fOgJ+j9nBAuKjoX
iP7dXugtrAlz36E1McMvBg12WF44mth4IcntC5gaSXql5ZVMlplQGVV7S2mr6aVin62qGq1PBYB4
6BsKbYU+rJrS6U4HXAPcHB0T2TLMe10eoxwujp6CcXSnT9BvviriSIgcD8caBZpehz6bzYhmK/Go
HyYaNw8Ba/McT5b13PdxNAVACbVV1f5DgPn2cEyYvmg21KuTmk1kK41NUJPm/35ByWnrolyvND14
EZTZjxw7pPlnliT/E4qkOYsSiBKI1fendvbMZEQ+sB+zQPUOOJ+GqHL+5waF47bOP5/x6Pi/oUrN
zGeNb79gYHxT5DJA0mOPORnrq0B0II/Fas/gUR/xAV7dhObZ51DpcjVN6MF6HgHufK1g72lU3RXn
ceVxqKALx+1hFjDUq1/fx5Zd6P6/45ByLVIEh3Xjyizqdv15RF5+yh/LeSD2x6W96F9ytKwWr6ur
1giXHEFjeiedsJeYsY4Mp59oyPjSrczWxAN/uU+6glbGAVNZyBdcCAeIM5QZYHpubRFDhJ6BUobA
DiaPuyEqqs4mRuNrBOIfTvoWX+ToDlGeXhdKfM9gEQJcvHY3C6G57i10i9vLDJFha0Mbu0tkssB1
MxqeXmll/qygo1K8ab0vRItdsDAVh1jkpA14M5jSadQpTAPbRD+qiQGCJbMtxetdrvYMLYmeWpnh
M5CBb+8d1+QM/bOwJBQ0R0cayFj+4iVyNmNCp4/MJHsiAC24N+GAnFhHABYgwFCnfS2o6Aj+8tyK
tJelADu+nWo/r+swUQahzGI1UDz+DFCZ/GnWkGrs+Jr4eySNuuMJiGsgrxdReuEMZJyE2hENZgE3
++n4pp6ePb+Iv/E6FrAQ8Ayu83xEEegeav22OCC6WLPCgWUOg9MStac+VivEAIKkeyR8xjuzV9XL
S3DbxRFBmMC7wm0inkMu4zKaZBe1qUK8PJhv8hiHVQHmc+0G/tUAAE68gjziuepHq+RTTY2V2BlK
3nImvC82Q8bhlNi2OQGbZIlMrJqrvicNpcyomp75jgkrgybHrtfTmfpgKl0lHx6f6WGYHOPw6giY
YYQt23gj6einEkhPxot7XbZsJhtlC4JSV1OvUZbKN3+oFwhtCQSRg4Zmm5DUPAHrIfCfpna5X7bY
AJvoWByeZ2NQytaUMY9r5W6cCgtFJbzCXTylCtP2LM/DDPsl7EH5ix/hwxl1hF6UnljdcyTGUkhs
HiOmof9r0Kw5qruJYLCfLaOTumeCyJW+CW/N6+PifXgk+EfKzso6SbPEt0Akhiq1rKBJxxSQPed3
8apTTQJ8Q6cDo8+uZNHKGTRtWcmyl3uNNzAdTkUh5BfBc8UTDVR9OjcAHnIDc60zaT4VCVy/UTQ5
wBZTIHgzrbfWqMs6bsS9uIWcc3+Hn0NnaoYEZyB2EqNfDK8QKlzybg3q1hwhbv1B1t/gbpm2gud1
p+bxpBKE/VBlg4kEN8joe/IAdMBAimLhxN35z/dWnezfJA/IXHzygeK//w679uH9gJshcuseW04e
qwPtX9eMfCALxxVScdg7MfxBI+GIke3S7Hae1uDVYQVDE1ZszrlGhsNiiUsumw4pGeur+CuF64Fz
BlY7Du5XTNL56J1LsRysuqk3qurDcjJYjAbazmErKPEdC5Dr59uu8Hk2KB8chntBhZix1+79dkKl
zWysSNqaFjaFM8RCy6oGTdtdkE7sAvwG3xcssWw/GV955767BjELUn5XO0nKwxxxEKEVp6uX4C6m
qbWkFDVoLC6j1o1MsaY4lidKKp8yURrzVf3ThSa9qg0KPgMFWYALGtyOeaZmLG6+ECVHZ1XGK24B
/zyqYGrLcUQHY2E5igWfUpn/2TO48a6fzSX8mUswG2OhPrAARQ5hPTYqG4dadhlSeFFNFom4lJ2V
lUN9WZ5cnYrH8+rJ1DJCuCJDDHQYr9StWyTi8QmGk65CR1zgwpiTxOVKzMaLvVIOZyyjY+Eai7pW
STcL3++igkguJDtTAIfsiEOB2DjsuYgXVEMlhGUZpvD3j6GPE2/GIYKuxhvyRBRbYjguwMXOgN9o
yNfi5JGSvno6gD+l2hjl9OAOZq7uKIvdnfn/UmLMYh/uneQvfiAwnd2FEn4uvW84s1w0mCuufB2E
8q8frUVjvQIrG8HxlbfN0SBTFpoU0F0PytmFx5W0cd70LeOU21y7amlmOqelMkta8xcSjree+GnL
1fX8qE4I2qJuhuDXDQZno+aL0mnSn9Jtt2KCfLdwQDABYK6/WeykkTVgyNR8B7OjtbpQVtwS3yh0
NcXRFtU7Npn12LnyasnznxPEyeXiQr3JP0tr+3AMte9TAXJ0qehKEY2uhJHx3mfYFNhRT7FlyQo7
R+01aA9cZNLvY4nI5Aub5tZcJH/6IGcGXNGzHKVBOU8TExqiXB2bX0h7C70b3urWKWsWkKyP6FnQ
vNrQMuarlDLVJz53gHPXAlDFmzB1ZE0/jbHS6UqF8Kuwz7/nUwtmfcCBgUnS/hUTvUrtiZrKzgE+
tFdGffYUASH+ls9Xi1be5HSp6am8i32DNlx1uHhUFq1w2fTeKz0NK4eFJ64Kmg3FM1t28xmj14qc
EGWHOqrkVZpcqLp8V4eM3Q5BBhfnbGzCa9yIFGM9886lxUak3HqPq7F0fxUMCPbj7OyvSEZjQeWl
rWkG4ANmkAjA11en4Q18LedbfEba/rK4vIAldpXLzl3YXF/xRijQQmh/eP543y+1uC5QoagGX1y1
z3C00sLhjUg5CRd2/8eN7YV4GOgEOTJ2qZsNedt8m0tx+G8Xwo0XdBD8OZ4kZCrp9/e6b/f2Fr99
uRDzEAXXElNzgbsU/j04HBU9545JebFNYDf+kUvNwGoly5dJybcsfXWbmm4B4fV8wJd1RoSDIoqf
D7efVqtxGw5Vv4Q5o1hoBOfjjhEKiRqWwlpciS8n4ANqmGBVirAssSCgQpM26Q4tKoDWvaJOau/D
9xYlnjJ1b2pf4NmpUYyyOd+xtswX6WVUyjjsiaa7rfWjDyFBvKZg360xJqJFMTBRc5uxiD3ziDn6
1oY7codQ9Arm9noJb5TpTzBH58lIuwq4n2/HH4sq4dm/Ge25kly0LeyDtLRZgKtsuDfz8skVr6eV
hklpE3FTS4pwARKPPKmpkWeDGr6+r90coMbqf4yuj9MQltaGECwUetis1+1YjQA2sEcy137tlWDH
Im1IgjMjKw0vuhGgTpdCij9Ow8mJTLyfgCQ6gcgvISCFsS/lx0vUOPEhPxk7MHvwkxp1pSXKaSYv
KskBCgXmBdOqA0pU/XKX2Js7UsYcNzC8GVioHsRnsBdSaJTPwWMUuX0Pf8B17kIBul1XDqOSwjca
nWlDbLpS5ElU3VSe89eNe8yBPOsTG4qZf6Lcf/3hvNc4j7Hx8hp1V4eEAvPa+trbMAmcRe1JEUjk
jKRpzJWyaqLhm/PBBJ/YyQ00ajlRBjGKDmiU8QpDO3KPx/44gt5D467Zz3vCGIK4Atn18phs4uXh
xrZSU9TFmyl2QXMUdYMMEKeJIFsdAji+Mey6s0bzwDF+67fO83At6JPjUixtf45UhAB725viZp5H
IRbTFu4/Loa/qeKGNPuPQg4X7rPIbjWCbNNx8Y+8NrAFBWdgL47+mzNFWqkyGBnLhnH+w0IxTJ3o
FzOowt1hP4Rw+fgAX0QiaZ7BueoHaSpD41b4CECzyP60ayMrZR42m6aeItyaIoerx8lIU8bmKq2z
Cr+zNXUx8+5PLNa+TVds/2jgA+YHb/vPB6jt+mjZYvA+ftl8Q/mNmtzgOKbUTGSbfKepaCIYXcZP
PCNx9+VkebhG5l+BpxMo3da8661HDPu4mZOZGjnZAZ8symIGPW2D3YONq5HpbYcDwqek7w==
`protect end_protected
