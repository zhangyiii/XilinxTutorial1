`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 239168)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbB/zJnlY9bLi0AUFrGn2gHL2x2kzl
0IsX27FVgcMWfMlKehto8ZKyKhqi5agZner6MSOlTj+snUolYVF1edgOYJzeDaPUVVv6ZeSk8blm
TTIcMUd6qN+ChLfF6bwTUDsxBfd01+DxRJ651LVnE9rBXmMZXp24An5U2rljrmxpFK5tdp5eVmL2
D76GbGgA5pyjzQRqZAdwvK54EHSPt5ocp2yBmegKTx5jjQ93ddEPs2/KvOqvNG+5rZJ/kUbhXXxA
Xt8ZiILf19bJNV0f05taP1rlLzUFw08h5/T5C1SSbaBwmL0u5F4Kh7oQAZ9xOePD1uWJcsZCz6A6
JJ84Z+Avc0vbD/9wmDYUl9RzjBI90Nt9cKNRZPdLD4ed/q5QzKXv7bhuyi3wXLU6WoJfPUXUWcBw
KaeHxJrpVBHqdWbOaLAN9Q5mVyLzGzpIDYKjwvKWWR1ytPCUj8DPdmZpR0leYW4F2CWmlfvhIaja
gsQ7BzRssW5ElV+UPvNdaEa32ENdlsDF4qxLyrHtmwqEjTPY/PNlOVfnzmrD84PK3ytyzhc9DkAq
URLNsDrAWUcM8Mln66w9AAvhqctTXxIMexK/8qrLo/1RALkXyQpooJ3KxLTiwKfOk+weKFuSXOX8
6tBpZUTf3QtNjO+NXHc5SjaCxgcFNerMJ/u3xVowufmqIdeT95H9qLh8TJP3RVkl8+AT+pnXuHfw
G+BTk12O7CzIIp9W39uBtx6FK6IWEYkEe6JmDhMBR652klHh+VBEUm1PMGlpnopXNYCHeG3CSm3r
EoJm6Rws5Un7PG77rbf9HNSfq6QMLvG1n9dXoDb0L5ZfRu3x8Xqjf4qehESsvgXEzas1M+l2FtV/
6vZnTNsky/BzoCfarbapj9dzjyiVSqnxgltnlHY3SfRcVk8Nvl3HhNtE393YlTXstGgIgp/eHN9M
h+AweUc8DDYqeBdQaR0fsoIfFRTl+wWbFXCCUlCDasI2fZmZ8K7cf7r1KcxlG/FCIIBODwC7PWNb
+iG3IFVNAxhS1QWCNCtEq2bFCAbsbdglnkogL0AOXaw79yOThEr029tCQ9q6y8spgyy5Ad/v32R5
HdSE6snFdpdI9jRNTW8cvDUazb4nvzWqD27DgvQ775iyWuiBNFwUNdR9ihRExBEi/sXB4JWEqVqG
EVR1ofVEvQ6CBM9ESnFMZaQECAC7z52THHUx/UOUUSLJiYMbFxN8fyoKRq+Oom/RgxyTsruuNdL2
+rCwOOE8AEOMdDzde3F6OYX5NEBbq59vTgnalSiekr7bB4D5gkrkZBOfjh09yqdObHlQXKEUxeuD
g0cX7iTBiR7NsAlTyCyaIFsdeAN7ot7ErJFm47gyZP3arOTtQ9gKjdmUWljP2+Owve11aqNMjp+0
AxS0QYMSCBh6phR4RcaRRpvZT+zaqIV/YDWCOVj3mEYDlH9ekukn6Q7jNru7RZGcdTsZV1yEqsby
6cTrKGn2Y5Ho5F5cUGDIw9ynM4QzA7lfUPMws04Okmly9vNGIspcw7dxRGKAneLJpYD2NQ2Lm4cL
05V5YdAT9iiAQXTbQ91kPBe2OreE1UTAnKNlemMElEdgjhfwenSkeC/btuA4J2/I/ZdO+gBsxzNC
isZo+GBNAACOExgrlM6RKegSLlWBIW0ZbKKQQ1Dcvf+XTEe/sbcWG1EcmNL47g4C1twEwDyyDM0+
mnn6bD1aeyIuetRJtqRsGBjsxqtXMvpBoDiFkRYYFXadR/0UubWaJVqg96exep0hV8ZCYENPhJa/
M4vJAgkkjIPaUB9yG/oaQ02NK8kUd7LqOAptTv+fConkXKdtowS39xYtKtK5hVRMZ9rG3WafIiGG
upx54kNQlS05fXghJGMbGySgdvwG+8twSrr6sqk5XzxxjOXPl8geSheKFjTRJdbav9uJ5IlgU7wq
PgqS06l95a33gAUa1mMXXQsHeRSnWifapSnLTnJdWq+iraI3wJ+ws6lZstlLaBttIAatR0KXJI4w
2ggTRjVzgP3KzH6xDCEyDdxn4YENTNw5U/l7eFed2YSMiQKb91hVW7hgKO0NiA9zjQ/xbrqiOR16
ys0ImX2AThAgAywEdcnxJIcPbT1fvLtab6llQjNHU7Vw3eL03p25PLSsRL1yb7UiExpZRmbInIwf
E3eLA/alGqoohnbtvCLXIJR3c+Jhqpxl8pMdcTZaVCt78T10hWrh7v9sMxSpiSmTj0ja9p4pQ/sU
CEPADPUKEq9+8O1h5dY5If0U5Rg87PRGtxy3gYxFROoDt92SdRPxE7DoMWlGH2RPYuwEESHJWKSF
24P2JAIg4Yd7FTBw4D5isygHgpGS9BWKkqzmF2peRw55f3CLa1RW8mXdvJpvK5wress65l0U+e/0
DMKnK8NA5tM3wqg9bHAxbfhCFU9V8NrjAB5vSHMYXCYhxQ0SKWi2MSnJoSgEcLIPHtMutMNA43uD
9wBtBiAgfoacpzEmjHAaUAIXixGvSFgZlwvGZa5E9E/av3x+6DLJJaCBD70V9D/nVinK/keFyBk8
xpQPf5fVn4wabklruE43KuSs3uTbLBlf1WAy3jC00zv4hTPoL0BYtlaaWRcKLqItXctvolu1/Bsl
4AlKszQvlUR+cIMCAB/3IlFzrhzI9LLM3wvVGVSwExY3CocrDjyei3LFABlJnfEhn5ulzT6urMVY
x1CeMkpLNeeQROHq5FApuQ7EXRFTxod860DFmCRWzD0i8qcavb0101Awolj1M+2patGl7YhRT+WX
cMsfb+N1abTQb4xnhb7XlFcGj67bhEd+ZP69Vpbkf6RJe1d8fvyFE3UvgzUUFfrhl1yv5uDU+18y
OdoJvm6zyFV1Ofco7FL9IIhX0FHbvj6N1ZyNdxgzRBii9/9lBnR2OppKaevkq7u/XmHkPvN8vIzT
hRPUw4/jo4PkhEmrSruTpnWK2PFAbD9bUa/UoAPtomXV/Y0Qoi8tnk7DcdpDkQFu1TG0/0Y5L9w3
YkwzfXHDJ0r4UXRyyCpGVHYLn7YF/Qg55di5NBP82N3alOSyb/njDjZqH50zSSb1chA/R3r0fTVx
hv94DYJyNedSPrqaAbIUkzZ0tvdK+EbXpkgaF6FGxImAERB34Pe3htR6HQb9PCbCtkyNjIt8UEU/
6Z0AORk15EgloWa2Gzi5PLSNHHqYEOnfh7ksUifL0Lb8UvbtGLDr4CAGF8fjUbFsoVMp1jJil/Pc
buJ2K4vWN8DT34+7ovbqo9X3q3Socsr16pm86c32INwNS2ivOhfLPCsDR+A1x3fyjZN8/Qiwc8VY
UFg7BuCrW5OVECdU6Na5uwhW78uOwFYNTePn8pkavlORv9M/GIxiD2NwTAdLY05a1QyRTQzHXaVy
KP5aOAmS3C6n9ItLeL5WmYhsM5sVIh6l+gBPChjTtNcbni2TaZazZ3dfK4GjSA/4270X/CZihgln
nvc5j9L/CAdUwNG0AX3mSxqpzk47ZAc7Biiq8Adev3JlOWCfIRt687hvle+/0lFKITJuGrD79pbN
qsjs4ksSwP5nBztwQcsErvGB8JCrT5kizTELPTiwNHRl80b63qMDdfnlUWz4Uh+E7qFDHMYDGYJi
lrCRz6UU+eMKOVpVaS75nHqmv3joWxU4VlLDJ+8eWppB3HY4jPj0uYs+g7RojrT/aixiGMF/uS23
dPzUlAlrsf1zRJoXJKTlXV2GVcXNfTwxbpE/uFCN2AszAzHMrxSjYVNeVUUVcVghEmgzcEZm86VL
4fjD6hEu03vuY4bqCKL0EjfOk4PmM2kR+HTQkJyvrD7blbESRiy0wS0iUtESERtAqcjLsMrRv7d6
mgKiWO+g379tWMmR4eyjjVWzZhPOeOw5LWrEDI/MTtFeW3njAkNUZo2FQ4bVyGC5lrjlzxLnZqUu
oVYd0Lwo5v0TRUfU4YxxoM1yUDvygOrVd2Pxv//NT2gTMc7nNxTiAmnSpS1CSq38TgAACA6yGJcw
Rfqne7e32SlUPofjKvXNJU1wNcUhtoOusQqxOYFJWDaWjmrrvVqsgAKtn/cjzqBgaKYTm4YHhSTa
QPPIbOAu6uq59U27RVeRm6sGWirmtkbChAch+RSTcHaEygF99aAxLip2OeMhpnQWBMRiVOD9QZ5m
iRQtqIctlu6JNjgza+31mJzjkkwRoLcA26GNZB9sS0fb4y43QK+DOsOsINVCDMrGo4yRFd4k4Urd
I2BcdCGiM1WV7OpQz3Ag/JevNrpssk67BdH0syE0cMZ1/CxQWMcNwdDykneA8rVkyvCFixg/I3aq
1mx6Tka5IbbVgYXjvUZ67eIv6eBBstJ8v4HGykEKGxzM1mgPU/61qylJwILVTsVRSZJqtSHbjNtv
oJRyt/I/kbr35EXfxZhiqO76y5p8SfVlcJmiSPdRJrCt0Zo9oVckNjbBqdT3/SeD4A6WBTgqtrfF
caJ9QRDswlKsoAM4Ujj8oMJGt44R3+K5OcLQ8tA+meynzCVOk3KevYHodHca3YKVf1AWuv31j8NA
QCFUqk2GjoF+aMnrjLFT8CWH8ReQp8Q6qmDzyKdLo1oqp9qh6mS0KD3PgQySlBNc5HjXaKtHtzaW
/hVkUx+pAJLocin0jtCB8RAH5b/alm3tv9lkhRtCYSDgXw7OIck/sznor9Ovb9ignrXz8RHUWi6F
UO0I5HpfDbwlnC1Flg9QO8obAHIQPipe7RRPFrEgHKVW+OzwYa6/73JBuCGQaPAZTtMTd7ygwGmQ
jqXPSw8vCqZvb2X8gjzJoOqP9tUuagl/KI5zNDQXDrLJk6ap76M9x0OT4PkH38DlbVS1htK4zEdl
6ClTDzHwox0Hauh9Kyg2XZWHonm29O6dSfnZyVObFVfgjn3yInrIZv/ulBPCOfcTY3LWMMS0ql4G
O7bUEuxf/8NAWFN/U0mAfa0KmjD7Zc1P34tFVA0p/Gp+VS3EgxYZPw/KpoNwrYBH/vJ+ee92olkB
Mxennhm9Gqrqg5GjnYzxt4ezjWQzUHlF277aoVsL7B8RnynsNbQuDeQ3xoaOGZfEx2sqA6ZvTiI8
VNKf4u8kozDb3yC8UnpBOdAz2GY1yfuQtyQN7ZofJKPUHGNgfAisB1zrxBaNxIkkH8YBtt20qm8r
dEpPBeiHZVfQp+3AxWWNPppDzWmVHZ0aj/4MvIoqAtAvaApNtCjowOWKdRwlcZd9CyUxDP6I0MPO
bRpSwzxIBHxuDVPE4uqaUHJtRqSbTosywhNr1wdX0fFrefj6C9n01Y3SMvB+BOFXF7o0dLZE/e9u
NJ5wg0fH0Ga18dCSRsTYqptTX1As50zYXdjHPCJe3CrRtyLdLQwKChHageMkSYOSVBeRX4Stq8o0
qYO//h+mKrSjtB00vIi1kO9x1KYgqebXSOm0AZko8JupD95S4SJio+7iHDIMIzGF+QRBn5PZjg/q
B0oeYH/8e9n6ahy5sj5wLeB7H9eAIrq4mCVm50VgdVPqXCpt+9T/DJ9xuFDHZ6HVfm4qJTqOyJ6k
kQau09qHiQYhLSDwNGC5bQuHWK2gsEWRyKd2vyjsBQElZpVwq82pC+mmoWyqPXupxMb8g01k2K9F
xHcH72Ss9dpxagVbsxwi8Q2layxsOnhSFTqr3NCGxYxfilMllbUQuf7y8uRKNoUZKCbgun0rnMmD
SaBEQAR91I2/iZwJ+rK4k/twAttCY7EXOV++StSqHniyRgftCladYO0UZmJlosb1SbWfc1X4kxxx
CSMUIdQnAdNehwCMuCjy7XIzvU4lzhatauZ1jtHbKQ+rKoDhAdwecs3k0TZ347pOWlsKPmHVQMom
hRYgXztTH1F22MdQ4TIeFHKGfEn3VBiL8Q5pBXsgkE+RIYI44hIrWVMDoP0ia+m/0uVZ2dylsjkN
qhWUpsggBlrV+5d3EqhBSFJ+1NkhUYZsH3HXuxJcDIfd5BXo+WusLuxn7uhL/W+eTlkid8sVWvLJ
r/DDhjePpIC60UP84ne7sV6XdBN/VWEdLRx1Ij6OBBgXB+Ut7J7pP5oFEBxGpzuBXy2+RWAxrXf8
R/p/OgohciVoERdAOcmLeAK8zrk6cQD2tYhocP/Z1rK5oMop20/kr3fGlsjBhqwrm32Xc0LD8nNN
SBruJefvGEmwlNNIVSyx8+ZHvnzER+vice57/9/xqGvm3ZX7l3X+eoxmZHImc4CYv7my+CP+tiN4
tmuRg7CajvYigr+BAEfngt5uB2myTF+37KbonNQpAWBnrzC/5nDrKEIhrJ1CdnhkT2VK5z90A53/
QFUrGZF+gR5PjByZbHNef/43VkbH7mRyd8jLboQy8g2yvGipLjc/ZA8Y49RfNCL9ntzO54EHG+mJ
v6vLXZmJTBEURo8a4jqSf0qwL5e4UcrqgOZW8P2jAVk8XleMcBMb35RAsyrhoGYzQ9rhzebsokg+
TBl5gkjHLKRAKouZMMI0/NMoiLqsnFOUHsuQ/UPgZZjHIAPvEnEiKJDp90skBuxOgBNEJ+8SxJlb
9R9holvZUvymZXR7U9EY00+MX9z9NL2npvqqTpHCo0+nM0lwYZQukJKgC4lzCbHZ9wYg8QAU7bXH
a4hE8PTNi64tYjS8IeaKDAssvhij8mGAwQ0R+DYdHGEXHoeq2N7XSeI4KG1A0w3/3c1/xYpMd33f
ArzFj4hfWngMiwafWiPMADc36hB8/Nys7FFPBOfb9IPJLM6P9G9AwrtUflj2FEi86tc9hNrb3B/n
Sciaf/FtqFMo8Vunxea02M8RUr/lai9jI+JpZJe1jcBnVfiiFIQ755B/6zl4w3A10ByN8IH08UIS
EQAlBBYKr1zo+GoPJrILErZBItG1x+oc15Qp4egZuSYhhEGu95ZDMK7fjDhzwDwFAnWy/RcYQ3fq
eKo0vR7XFOzwfREHgKNtAbS1jz+sJlUs/vEV45p9mQdWGqLgxazMtd80fXIGmol1EEYhQvCSq+L7
d4PM4qcFsoJltTUnmIkVXr2sgAU+QUlQVXUxFnzn5uBPVHBGfhN3Zzw17BmfT/6ycAqcPJaF/w/x
gc0s7EUgRj4jXYvsgRikt1w8M2yS+Kd4pWCKmtt2PyfZqmzriiPK5cQI7rD08nZgKU49oqiV07Xx
oK+0Ckd81pH8GoWXzWTyQKbXdcs934i93Ms1RAmlSprHFFLCJQnBNwKVbS91PIwuvSz/D/f6mITM
YOiePX0XLSsjDMONcNY6shziDx+1rUFJz5Gz8is7erbvymbxa5A9SyczcG37Fx26tHY24H2vBnwS
V1BeDaGExzsEyeOdBbZK2uRnjExibut1qXxaM1/l0Mnw2lUiuHBBWSO/R6/2APttiHxp8eNjGbIf
SnnVfZzKt+hPP5gmNn5zDDn8w18JuM+bdtFiwW4INnQypOrVNnUmZ038C3WGryUvC2KV51DiNa8Z
c9zL/hbxljWNCZlhiFOk2R1JNlaQjK6v8EgYwn1HLBb4iZDG3C5aew87cEQoemmou/ucGTGi0N/N
Q/chUOFxq1J92tQMQzzg2U2HERlMGe0kYvLVUU00YNvEfZUE8io2I/HhDt1oaZwiSwLGz41L9J2y
euYLzuNjSNAjxK4hvMyXsOCDPCe2m3zWTE/nCpU5W4wv9V8KFUDbvUpKHFjyuZATVbTbp2+FcJ9b
7rZ/xMYjp+LwBue3+FDt4uhD4Zi16TS4melWyYKS7g9/XR5Gck3JmbcCYTOm3JpEr6A8F4X/kTaF
y3nqUhlb4Trqpe6PdLmHztLLgjUrq7RuLeeG2b5/434RB/sM20Q3vbVNWJLPRruH6/boGWcHhdeN
ULfPaM1Y/8xSnCfoL/NTbS2ZEj5e57Z1KcKe0KqFoyWi1gkIWxBB3lRGvfg3WViamMO/BkapUzG2
q/+ZbIJRC19wiy/+0P9/zjFE3FYS920Sq04gT8zl/+gWSQ7t24FQoBFy4qFTFsKq4sar8fFs95xb
5O3G9rPOR1xtGOomkGgoYlK/XJh0Otb8Zy1wX84YNWKHq4dROTwlpaa1Jc6Px1rpl0p0AGPonic9
NE8buJeALsS3Mc37O2F7BUswTKlf3SX5ykQ3KRPQWBcGwOvS+b7RI6FoOHH4upbTX2PSVaWJFw4y
ybJKKpxHyR7EJ2SKLIiGag+gdP4Zb7BZDUnyRlfdrw2ItOixLy5ve5ZzO3yMlJLnQDcSNCv5Bx6s
+9baFuq8jltR+Kd+y0OORjejPi2Cv0Ihby/LIVDgd4iL7v6tYlrhPFCKwmDXMt82n6SriUJq6Pkn
pTbd3O5YpRJfKMCFlbf2sze6pGz+WM4eKweDoRBt4aWfnEJDPEcj30HlAi++Vgt6ZlNpGyDwJRlY
qkBCUfMFfvZ6dwojG3um93VJdSFM8MG7ecYIMjc1qnvRCC+1CuK6XHoTD2bsTOeD/0pk5qTsMWOL
jdawq4ETHirdTtYomyHJPpsl6GwV0vEFO79+RBysGLR9uVjR+YHJCxDs3izIPf4bh5pgTVmCaAPN
+wp3tjhsQsfR0a0fRei8hrYMMwnf2+IzQ1xRMAnYnkg8ZxGNG2ZjBL3xVVBcOrmx7xMAG95EevT1
SiJrTjkAGprs8C9IrBdmKjDCB7D3lSYf9GLDvBZ8PU+GPg6lfslvT/Njxldf3Cs0gWW4D4+HdJ4f
ihfA4eeTgx7GiKLtSjQwBGxj+ZLD5UNffsHLpWA3Ojpx9o/U0Pm2i4RT72m5WCv88+GAWBgQr8Zl
8cRWv5vNx5fakS+wG3La55Q1UCVIOqJRKTmsGApaAuewR0bUPVgomHTU7BEIWIpLXU4niGTifv2I
uxitSHWgOOIYi98V16I0KAv4qx8lud7FIgBo/PwlKnyFr5tEpiibtiUipj/ZVzRvgwNO0dZzcUFb
J9ZXs08Rpkbh4PUe+jjjuGavaV/K03hYfXi+oP+ip+b+2ohMZI7gyAPKUpq9MYjUOT8AlsYzjW4C
FdC9pfb3XJ9ztw4SYLRXXuzOgzT7uy11O4xWI+lg1b9hnxoEs/MP69cm6rNPmSvFyZ9EJ925f6Pw
dZ9OesluRubQOQjq63/eQHsNuf8kJghkVkQEsDvEE0wQcxSYa/ovlKOJqJUIxubkLNjpgm8Wuawk
Qmy0CS4mt95X5/IYJ7EFHQSx8hg91FlajpfTSx7A9IwjVtf2twu8L4JfC6nHsk5GsQ/t+Yvs7BRG
aTDxPp0KOd7mQOt29YYFyksY+d/rHtO/IRssYAfhr9j03Q/XE31BjZcyq7A1yku1I+xreGLDYfpt
v1zhxz/F3Wpp+qtmoZGUgLg2F0TQH2qyQbi/vQT+zR8dtyBzv7pXpUAmaR+LIi0nYgDNmpzUSrx5
H8UexAQXpetmwclpi2YGdNdgAr4qkLo1gs6lb6SUoz9aAslrJ8hYJvOuFJf41US9gU+5dvdz4zUG
2lGGY59e6wcrcstQVSNxULbKjcJJCqtSIwkZ+UOuke2MmuliOaEz5pP+G/Ci87h3+LVpHpfWVQCh
AeCqlYc1xpMKb2U3R3gT9TJ76MW/PkcFyOv+JYCdERzbJTA61DCmbwF77GqnRoH7ZE42UYBX6gcT
SyUMwpjwsHofwqHp6oG5k00rvp0/UMusvuqRSqAnQXoQdTkhAwnjpITgUAZuI9ItUkoiHs/1mLbl
zDClxlHSg7rIrXuh9WSyY44vp4upmyRrHj2thjNnfwavREym7iqTvZDw1lOG0tYwrYznNh3ie7bU
oFP6TmbFvyhx09ZnzP/ZZewSYTgnwzWM7qbB6NIiZRoOCaP64dJVBQU14MGqxrXYU7UaJSDdHuZY
7u55CJWZCmN0FbK1qtbpX+5sf7oPczZRv2yrkjmfkLyYQ3bxsc2v0hNdbZDxFTka3kK4x6Dypuqs
wG3mHL7+sxwC61oaiDeFkaDEVt6ojBEvDEAtegNtu0oelOeK2E1g9Qi/LvaoAHz1Hxiq/fTuF+Ue
ic8h9J/rWRxmgsElxDzbqxVTj4QJAE1C4YFvXXfXj5C0Ywy8rElvFC3HykanGDAAf2cE2MTx6n16
1Mj3A80Q8UYxMXv5PDtavav7diIHMq+YjwI2sBjU4iEWcaQZPQ+murtVZC/5n1NRGjTJjxlF3XlE
dO56V5cMWsxD+g4bnrx8k43hgKqVb+TQLG9oljfzT8Jk/tzIbgyIdKctr/puwXA8nR2I+WhUFAXd
H516tKVADPmY5eEp649ZuAp6/k3cM5pcoPy8nVHcyfWZZUE7Jg6rsfKlN25uYKaUfuxmu/fcJ3p6
DlNVkvQKv3P5mHKkyCNf27R/D+HKzjIA4YF8a80IY2sbMEmK0C82R23+SV31dy1BChkCHEyFyHqb
Y7JtQNIM1li9x1gHrO8L+LgY/Io2PpR8kN3rLSx4/KO0z5PgixVk6DjvamoVxoOr5bKBcFPBDeHN
4FAFRhNpX2bxf7kSGJzhIpY6oTIiWrN7RnmJAMIcIIz+SmC0YCguPWF0BLDRVjJjo9Z7S2slVFHZ
5ZF39j2zzcpStA3oxqPPKRhg+or6iWKu8hGi6Nfp9zHfdbKmwIQHUJ1zZX8SEcl2aoY8NLLe9MwS
ArcTo3jxCLC9IagLmGYhvh3xbNQVgJNr/jVDHv9/JJQkRvrt5V8XQgSdySvoMSBf0QMyuAvBBdnc
arllgkvQpgNIn5jO6T9Xy2VP57jmgiUa0YvMdPBFl0y3yH2B8ss+4JfVeS3V/CSTuBW9hhnmNVe9
YE/dA6P6OJ9djtxCg8my6hrr6Qb4t7qqZtmyHsENETwujnU86UmdyPl85h4l6x+yVG1Nsx52BVhN
/EWCDaV4tUGHNz/EzwuJCsstjPwj7hVJ5E36PHzTGAAw4fG/78Cz5FcyWCT2N2NB4SiT6j+Qs3nj
5y2ETRSzymR90uhUFNyusCsy2YpKlOwTx0PfBSlcWEdnTjrWuOk/BNnbtFM5T50sVWAm5R9ejJWH
v2razv3cPgtviop3SUR/X57QedrdRDv5tcEO92RqlU3fUECSJNiutaEBaTnUgps/gdqK6lVpOvRh
WIz3k9NX8mvMJ/uH015aN9DRQHn2Bj6FEk3vczq+tsv6NqndW/4sYuGnefFDt7h5G5rugZTBlckv
CKz5KQ89/K4Aomz6Kp4X6TgvtYlk1kGh0pOM49e3Z86ru2/I3fBMLM4dg9axLNq8rUJCd7UX0/kd
oPvgOPJCy8olCWU3DmJjFvH9QXGuHQEBPNEKn2FBrC+49Uql7pBGSWzgeVLR09yxdx2Z9ezUAmHS
MpY/kWkGlkRFaiBD/M3Jvpp6r31EPADJndOQouyYCMz2b7KQ6T7MxjmUyb808O9rtypSU8yGbw7B
ilXyIT24plkNfdq6YYmu7Iiaa6VNG4Zpy1+lWm0ywO1C/IoStuW+VgWZcRj4S4oFRphnKxNm2aU3
McJQ67YXLg4w29B34vNwTnPU8c6Y7uUpvLVzQlA2A7/9ly0Ch68yvw8iG4rPcHi1hObyZjQeb4ko
qkF9FCYSCrorMWtz02CUfK8sf7Ow9d671RVg423VPOKy83Dpntr0gWxZt7PDTmbytSCm/AjhTdn0
h4l5KvADvyd8LlFT8VQxpzm9XENIC1eGZ7lcRehL5oyS+DR549PFrP6rre6SF9/ykzevNkzSA5Au
fQS/dF9g1WmQXLjsb51gUFdiPjregwYmIscxk9DBFP+YkgkvTfDVkAgQStKbNKvkJ5C3u+jLUpB9
Xwy/gZI0JEHDRKlSBicZg7AF0QVBt2e/13Uqr1fPD991DHKuLCjtI9SEDCEpLe6MFjA+yugOzyiq
4VCKtpV2MDWCBgsNA6fqWoEi+6vFoZxQZs9GopQu6/7w/domWYsSDBUYczt8YZ/kzhF2Bd+N6kr1
b5FBys9oyHB9yFGzYUIrzx1PYA/4Ki2rBWVKp7y3E9XAp/vG4XZW00mKd6M1EiGJNio5f8fZMWSg
OVpRyfI66RsDb0TaKAV4RNkW59JJRwejFSc0tYx6a0STRSKsYtnkuq/fw8l6UG77//nZddvbJVUQ
v8aW4cTbbSWs5fk0I2Q2asxJP5vfaeDbv8iijrTYAPvsFbUKMxzBlVRqwCi30CejnQThshlEmBKb
pmCI+oJqnqgDVYgUdyR4ePpuFkJbfrsw6dIVM5X3ZNXbXyvQX+mcjCdFUeMhe0QqcxJtskHVluiK
f9LRygHl/WC1H+c4iCyoSz3dWNAZ882Qgd6D3MlUiZXbESQHwSgjHtewpRdczmKoJso6OCOaXcgI
0DluAfzaAFNqoKPu/KsSGPL1QSAaTzOCfutKNpb4RZf+uMK8XXY4U/LvL+vuTGVZ8UCX9xD2eZnp
MqJsox75qwDOn+IwfcCCmP7QFtpmNtkSmhPB44kRBt0+9DbilZt6pwahBZ90kvMRsLE+ioXckc0M
Bz6JubF9dW//JxaKSGyaai9nv+3/XCzlJik/iTgGSxsqzb+KfnSQVS6wBfZMjtn1LE9pdiTEAmJe
++Umq8VriBCLbmhsNdKww/9Vf5P83PBTg/CHfMupdNLg8QKCfrI9xewa6AFx9tc/jtXfzVsrWvoD
nBWrvJYKOevqsfgc+lOCGDLubR+225lhgQ6QNh685YmMCnzFQkbA+NTSev9rLo8LGdsgmBtrO/zc
h8kLz5Ty3ulGqszEuCdCOsACz68SeznWfrgihF+3yuKolzaojPD3DgPYHa+7xBYJihxvidOuy/Nf
OAbQ0q/4fbuHanFIowi0deZTowxZ3B0YulwyQsGzsShLHk6rAyYB2QN+ngc4ZVCmqKxhs7txEh4u
atGm5zGTeujrA9SEHrS01wp/R1+VVynUZNQYYBwUiRNKpcWAapjGCiv29Lo3Yfa8DmGLNNF4Gq70
MlT3Gviq+e33lv8Q4gHBsrg8b18oUScYKyAsA0ta4tEl3y461ltgbpTKRZISWZyehpG6YGUTJsrM
VukJAzZ0UkCACqjO9ghJS3kyLpnPPkK3dNsCX3oNb2Fqr1/TqGyopHPtT3XMT5aYxe6t6B+0miAP
d03+dJhmQVZNXUUJz0dcXNSo2vqS2pZf08GmleT+TBfQvf16QUa1qTj7FQWH2mykwheVYAxpFkg/
Q+CX6/iWgYSF2KNsmP2sm/aQLYFiNBCI6uBT6d5EcW4/Oc7uI4tkC4NcNDCR9v726aFtAHfu82HE
c0hSyOkpKYxPS2ZfrEJXFELCWarZ7dQHfBpmvvyfy+lkziNZ+mtNYQjLHwu+0RgwM5IzdubqeAGK
Zn82HMZAmnI+vXydG+WaYSRs346IvxxAycP6SRYeUE4HRoduyje2gQfBTF4iu7uLkWstbnzepVhs
AutN4JCUdndAXV9IDoEXshi+0NrKlJb/Ugl9l6/BcqZYRlp5RJZzTXC5z+dqQgYLOJ2on+YlCTU9
ikuNp4ld4N66OB3u8u3epRPjT9fzAhmhTB0eQPDsds5ZL8yaSQTUBCNxX9FzXiZU6iu/ZGwiNlAR
uMGvAe8EnA+ts0vFZg/qiHNDG1SVm1Yc2FHBfiIaLLYFOT84938HdeNvto0extxp3DQNgDKfmWjn
s/jAP7IOReQ7bCe+UfolYPBKSWM6vyukedSPAnLVWJw8ZETRJiKRp8ZY+ZPm5yNWYS7OynisZ1gn
yHBXl78/Uivsv3NMh6TQ+f4Prz6FPaW30SrZBMG2uo1W7KIfFmRpLMVzcrQ7XEdIripdTK+hH/W1
ulFCCHr03jLBOsCH4uKMRXENY7YRmS20FAMZ/SyXbCL+6MFpp84jaGVi/vh+06QCkPiymRXc9Ava
itZ6w6sEo57ZiDLiNs9SUlGYOFqc/5GGMutdKZDoTjF7smwALyMoIVEP0jsmooHKgYbdud3gNtHb
eEEVmn31Wz65QE4eshiDzcuPYMbUngZIlC5hsIhGqAHmNh/Hgr95bnSk9g0732i6uHkGsKavOh67
DBxaybkyKs0cFHXwonCeovSBROXKd6sCTgmzxlKawJw1JW7jVd518mKdXo8bMDh+cKASjUv+D5my
e4EvmtbeO8NsmGC8+TGNsrS/RlewDMWTleWJshiet0nmDe/3BPMcmKHN5Jd/uOYtlUf45iJhxqGD
WldWFxKNvd1hHwptPMyhdTSD7z3FxHgR61DBb7WGRTrT5cKVwoIrlw3SdlRriCbjsF+bhfmmaYis
4MMC3ZHvJ86CFc8npB8B2kNSpVtlw+L4rihMsk8irX+jisMwg74Sa1/a+1nk3HcQhmDQ8smwCJEP
uq7yG41PzzORGrwC9l1KGx7H51QNTSnykKzXXrpwHOTwRwJM9vZ9eqjOz5CmkZ8gGRv7yX6i+NIK
9xxnZFZqmxsufVw5TMIJhVT/va5VpgLG5/lOP84wp2+zxpCbxeQDztiDAFrNqb3zii26s/VBqpTw
m32e4nzstkRIrfEDJs6T+x5WjlkxhW51Os66YS6G4PoAj50edoKVMLY3k8AQyhkfbyq3GGOijZ7w
r2J9RsKnRykymjBOCmA/B65QrsjMxJQVK2XJppsdzNRqIEs15Z6yZYUWtKrQeYqm7GrXJViRUhuK
Y5n5HNeZh9Nkk2N7D30nCOjigKuusd1UjorldbT07SHo8LvP7/dybTq2cYfSEPYTO7D3vqfOG+1R
qGsMJ0X5v7rGDGQ0pJK5jTgDPvtHqHHSsKwk7tlljxatbYOMC4WKuktds5zSgzKiEce1IXnYCKSJ
VZGIYW4dP5Evalk07NZCHJ3/+H2dV5m8yiWQ5XJwYRoSzlY2tvAZ6wuiD6sJDJX2xS6xLHMx4AZN
2mA4+ihsR43jWdTaJ/WRzBTozMtGGmd8sWzvFZT4MwH6pmy+9pJJG3CaA1A6wZpa7i3fqd0tIQ1z
AkJwZCENlvLZtYE+X+udPAk3b5TPZzT+s91ZxQEcaGwExxsZbPa5hbvhSjJPsCwb9AAr/+ucnw/2
K0EQMlTMyEa1JgFm23n9RyZtNhj3rods/oqp26fe3vjHtppe28f7ttGtg3HI1l7jQ/hEgqlefbhg
xYb4JU3eGKoyR9P9yJGbWRNLanVcV27DmkzVZ52YeTsoXQ2VesuMJ8Ml9ifTgimkTA6zGfqb2AVW
0GCKTIa6tDkjMxum8Hh9KbMBcClx1HRy8bDb2PU1nme4TVcCJQQspTWaFz2+xMeBXt0yn5fA5iIp
K5IcNY5dTRRVKUHQ6/XRuZvIzvs4bDH9KDNFiwrNiWy34m0I8vccYi++caPTCMPiRN5vJDt02W64
CrNTJteEXYzJGBn/Ye8BYQ5gacPB6qPzTMi6Vj8CPUcRMH7xuNuSxCqsqRp3j4kD5cpZRVUHUVHp
7qfyULKBsRbb1TDLQVPkdU+WoalajuHKNXRS2DYHPb81QeS0oM4PQ9xrx1xsWvO7kppDjn961b+c
UEC7mB9YqE3emc4NthMLUZidABH82vZ3W+gjQ8V7Vyb6VntM4rFKhUxpDlDVuNr3lIQFCw1N0CR7
MvTGAlJGq6qYICJjxbmveuM6QHGvYUVy9IwNkLFKexZN8dMYPT+kOEReZkFD9Z7R2ZpAZqreLAKK
c8sg/7tyYLcG7JLvAvjzZoB3HpJDtuTKbSzCinRezZfzgNq040M5inrSbetdmuMl2HKblc4UR0c8
hZ5AdgDg3bw0E4f6Io5ctUJsRAkrjqPdycCEsKF8w9rOveThGiuUxfu+cZsdYKM1E0AsXZ83tC1M
/loWVT3mOl5Y2b4C3oUsdYxuAk4nz4SI/kqsjWtF2yAor55xZpdr0TGGa3WgyA4VzKuG/8nzuQDU
al47gg5SSfY44l1ZiobmdYk0JwxuupjJzFwh0xzb83hjCW7aItiGaucakfAjvWbo7rsjrEzqB0Y4
02KuIuyTS9GycWKvIRA7hEDW+s8edQcSCbW+B1ReyvDgU9MrovpaDUM7MasHMIoJsMQMEIbuhRy6
UeDKDRih8WObHYcIAQdM7lQkYQH7JhJ3a6CE1AO93Ap44irJAu0tBddcyGrLXHnOi3wTrHnmU5op
kwvWDBHOxGe1DH92/G0V1M0w7rMUnPf8PzFYzXPCNogEXuxUgdwNSi3S9jE9l7d4ZVzw18Rc7sWK
Vo6RgcQm31tsM+13bpX/RM04WmKncwxkPP3zMkTofyvXx+w2o52mLn6Jy4cvYs0qevHjSLGXJiyr
arvkzCjZckBg4/5vFuYk4ZVpEPyky37ZLiTlEzIyo0PCqTK9Q5quZL1RINKvSns+47C8CLa0JvrB
Ozuz3JKz5kZKaN7GxQDScxxJS6TlS0IJQaXg21D1+E5yZ2yigbMvspG4k2ZaerglieK34ULRvRvE
szhehFl/P8ISNYIpNs5Kelt+WMQjVXboZTSheeYGOByAocpx84FBfNr/TL/m082xtjqJZTb8b5DV
nSIIxgLhviT/nRrjrkhw15n4E9DcFXljFfZiGW4CfXEvyGNheeufMMnLYKNT3aaZdjWSrON/U+pc
l4p2W3RfUnBEXz5U52UR1pKGQfza48XK59nSsafDSlSBTwOKEFkwN+3tOzr9CvK/sR6Qa6WESK09
iijdcDkTVLSD38zFH2D6/ml8s2hUF4WN3HR3xP83wHufG1zfCJzrcUDjrGOfLG4NS5IVgCINdOXh
r9sYKt65WcQ3knLkn4oCCfjnPBKjePXAKW1R2L7RjLLl4Is+0CMs8iYnrgEGGIUkJ/Pf3Tz1d7kq
XbUrV8gETQvQvbocP3nPtcfoa5MvChc9KF/28CthsTwB0acNZLXiqwmyQJFtS5i1Ncu/81NNJqi1
HA3jr8wxq8LSlfnhymwUils+Ou6n27IfGdn2LMYLEmSopPvTHVWsag9Eh/OvaUj+tynYbsvecrkF
fg5MFnWwisyUd2HWgrqcAqlnm+DWRR4PQfmkDbzsF7snROniDTXk94vwnyphLvHrlazA2LpAJ+PH
KXSoOMAfeh3Hw5vqPuj+oRqkEka6wuNk3Z2QrMLfc7tv17N2xTDdj2OBBy9kUR5p103ZDujAXk1p
QLZPBhOV+5q27ASIQYTAeBQTRNPAkmwH/yMvewVsscuHjsVN7TvKw6X5ltVp+x1vy0GRtUGcFJe3
6MuxVuriR/CgDWSg34PAhut12vICSyrCyNJY72ozZPcbdwSXEAqflhYseckeTWF8ehhjGgRkaAAQ
LVq7kz5F/J8v6jitanf36prwyCvMkjlaLkgr9rbL/+2ngaUf7i4aOAjY3uNBVloN68s5S010DhLw
sOboBSk+VHiljk2obhf54yWhBiCLuLlHY+7BVBvlOKAi+srV8aec9929rQtN6BUbiNPU6c4eEGSG
S8uigVNkN0orsJwWZNVuK3s8X7MVCS3arCXJez7r2VyL9FHvFMDFDU2sKl3D6TL1Bj9BnBsoYJLx
zTyTADSOOXvv/ngGsxPQY35bCzMzUIo1naqlPVzlfpiGXxzzH3Vfd2RYqypVtJ4tf4lHnTjV9G2a
Dn3d1q8bR48j4fZI6JWMfe+sT6fBQbyAJRyGPZSVJi5QXw0Y7p2sz774Tl1QK+B1dWh76lw5k1DO
G/qH4psod8oqkicv6NIp0C2eyVQfZS/Ckia/UL30lQZh/rrD8pnEfp74dSTpIkwuvLrObxMBNHDG
Xh2pCw7Yb6jUTaV1qcmqk8kbqyqIw7pS5KrH/7FZWo2YYTHjkzLX3IcHCjB7IUd2qPRE4ZouGxHn
HFfmUmeQ7LentAbvofMYRoQ/aUWJuoSV+7CkPBddwo710hLJhSdiDUReqJ1t+l1ndxZe5NrqMdi5
u605RtAEDrovR5pvzRXfZdn5B2EjmwePUomkxqXc2CeYWKv/EvWyxPbFKLLFZCyQFbQaIX34+iw+
xweJVf/2HUAANCjDYNw66VZyxrjqevrjis7QB3UOpfc3s9CvClRuWfKg+D+8PI3lmwFyH++Wi0zU
zHJ3yUGudbNK1Y6Mg91I+aexVuXTFFdUO3SuBo/3dIGoeem8xC5sNy9WGMnBX5zVGdypUpSZuiRx
+ny19N2RJMxmF5rQfqH/k5KDL66kTFXhMQhkVpPsxf7lryLaop/IMNk/09ZZLI/cFDHMtPro4e57
KzeDUWYj3MeL+uy6IMaq3ZwMVQNaj+/fJTRVCr81MkECbzM/QAZ+GufeYEfoKr6f/Rj8cw0Ir6Bp
7fAzIU4i/ODN/kU/leCGog8xRzy4VPjbP1ZnubsH0y8+0/d0DWjseoOx60t/mMuWf4h49E+93bWC
dfmdWE1EFJFnXyVs15Ubab1HzXpWiKpLaeH6rVII5vPHNgYl0Ns14AdlBgK1OCOiNjoFADLy2JSF
gJyBy08bAvj9uHUAn6Dk9UjUnAKY0oVQ3xXgfnK++DPic472sgbrbfZq7x5epzQBCL/1MV0Lw2X+
6eSUxNNZ8m9Fw1074peYNLanANy3ZIzOaOWE19AkY4nsqKJAkGQ4BGbE88M/ra1FkyUfhhRLkmv3
hDvDTyUKp6CcOjqjM32OqiDHJDkWwkBUxyGpoSFTjgRR1Wz09m0gI7so2hahOawCjT95urnmddq2
t6K59onYxByKR4W44zNry3jI0XvR3cT4ZK34iPFMksH7hgrL4IjxFUX2FBKm6diEdCmZ/+hapAec
OsHAPi8dEHSdZO+MGgo0tm+azKhzWCA2DZfGkTOpbpJBdALG4PUm2EMjw98AUA7U3ugDiiQIKZG/
2hdrpXxv6SwgZeA3buRpQkhMLKCEPyqjev8c9fslnNEAN1mQlM3dbr86ZXkO4E0JDvSeG/U9QR0D
TjfiQqJcJxpdyrRGiyOer1mGW+TihKljiwKrVSGCT9+52MqKdvP/26Mo6QC8wCC//rUGrpstCe2O
RIS7ddwpHBe6c9vCMfQ33yzCPeU5qOBz4kVZxqNkLlrLB9ieLuH5UNAJc4nGSHnhhpBXtINVWv/d
9QNJTKbXdmvNzFkMswc+n6UeKjcH/4lwNJtNsluNHCA6lqyT80dc3/YZryJ3AzVe/8cvxr47adD/
xeZOJDRII2gFCIHdcSKmN80N54YgR8kRlg5ETRZTInPfxik0GZewVo43WU68hU3LIZrRZZL3yGcQ
d5zrsm17qwS8DPh+CbQZ2d0JcccaGbmtivIcc9kVkJJwIdpFPXtoV4lMI1hQXFiNjswBZzxhzpXe
ka2KW8kVFzUkOsVA2KXhq/GegSv7KjHvk13Aj31+CW8Hziq5k9cClcQAdI/uOewl3kH4zYdqPB4f
E2ofk5bir9wTNHoPsxJGQLEbf9YtTYWbRkd0TkBB+rfagERXiDiloC2XfHri0n7AJVCaw8Mc04ub
uSMySzy7KcFTUxzpuz5K5JIxhc/JWuDyyxmzFvtXKDVRsDIyVrn3jNg5JrcxZo5EvusTd2p5ZUP7
EM0BG9T3uQqwVbY1jKkLtLAdmvqEsi1hbPgwvjF0O9VUJB0pPe+oIYRGylqyc+qzYK9iBzayK8/D
ZeXl9Kcgy/L2uO6ULsw+YITUJ/DspjztYTw+YRav9/CCxMyMz441BblrMJQZOJz8/3+HXFLr2SiC
ZjFEyXjfbzCsiRkRFwPXUX/Cgm4P2/DG1P+IBAOAfDajcdLKNxY/ydVE/93DfBBkuaJTYPBRaV7T
x4k38GNX8yP0LZTnIeMZv5pC1nJ/0iYjlV5SqAjHQSihJjLmJ2FvcZdyBR/0j8IphiA3+jF9Iv1D
wziyv9Uh1R9mYSQNVS5a5qei/nzm/fvgOP7KaAHdKjUwj/zYYhMqoEWd6bMiFIRUOpsnNS2uV9Q0
qC3tSB7dqPyeM8vtvVWlyyLdRChVPEoU5ztaLePmH/6jtj/HB/Fi1Y81c/V2fFuwqxFZ6XBUq1C8
EMXekVNAMJGPDQQgxdOZTaTOMu7NrCRUGsFdiWyYzO9tZ/a54MVxITNLE6cjk2ZOoAzd3TvxlBk2
CfzT7Csm9MetKOeDRYo7zLjbO6pSFGnUxyxafqeYtq/n1VZNMily2lFeP54u46MxjfTp9prwlqsy
oBxu3P1c1kccwVqgFsLv9PlFoYu7r67oZ/74zS3MjTFx/M1vruVQJw4ESY617sIV4XnbYifVX1iL
DrQP7mx69ULTxArpKG5n90i6C7TDeSELIClYs3dhzoLhIbYsGhoMZLIutG1IDV1rZst1wTRfsv9E
yfozgkX+4X1G/Iw47x+cqXa4UugMi/JJ656NcSc0llWcoUvZpfinNMCHCNVvsQRECYjIfrLroN6n
pRzABoS1Zm9PJg7ctZeyXyO+4EbTD9vMuppU4z5NxdeE+rsxFu+Cbnb7AIot27k5DeaFlopI2SKf
ZQ2qFaKiA4EiUI4eAVDHdNBPwQ2Oq9dptC2icq4md5WcJ2317BlRzaSdTSIhzAv6uXu0JGq0nqTz
mMELZjcnCAOlfq9gi0iUTQL2SimqGSTFoO1ScRq8CxMA45sVCBw1zy9fYWk5l6fU95yx8TakRu9w
j5HwdLq2oBHVzTNaDFpAgF1wP1HTl1w3f8VD7UZBFcmRlmVnwyT2oWghEora3/OcKN7/7eN5MydD
8k/xZeuD28BxcNpmADO+9fyghxP5PgVoqFh44a+uv95r8CjdepRqJbzT2G2RBqFGC2Whe7WPUyX8
W0M14jkyynuE1nQZysVGxgaqwbnQtbcqLbCgxvK5krspdMzQurKbuzJNTvid2xY7HaN1u18dAs3P
zZQAKwuQi/G09VFnECcG7TmrlertxC4DHbHJsPfWY/wxPwMXNJSwfnf/wpx1n4CEhMPkz97t/Dx5
TPuETzpFSABs+fVFT2Hjr37uCk0KcK3vnvOGZcVMk6rhXnoDufihlBLD4Hfic4lDwzaffzbqDLZB
j7PvuQBfJmmrnFFjXmNTYnAZ9Y3XFRNUtaWcGVV7rDDKFXLHKwu4AJJfpp1qIHPpI1Ix2dY3vK5M
WJDMrLyMEkyAOFbudVtEaVgQIGD0ROFquCFNKPC2FaCGiuujfWsbQVDpSWeptdeGNGH8WMGMIC/a
aJguO/ivIQo1Vr62lMorIotS0uULOP4+vTISREuSEAGsXr2yKkXmIHzxAcR6L8Gx4J7FtgvMEO4S
HDUj/ad1IEZYdMDGVKCwvNkLUqpFRK5vd3YNg1VnOBOmtbXGn7x4uxGhUEuxkiLFC9+LG1VRY172
l7jzvQ+B3D3WTeoJBu0eFkHjd3URMbncUVu0ysHM0A/B1VMEouy8n9ucIS1ngpP1kZy4Prhm5V+/
+eTH2n8UqgI8DADiLpozY9sckkFdtYmAe6w1XrokotkxNtlZTUChZcMyerBCYmEDES/N8B7qpBSl
7qvrzj57ZQnTMZ76LeSOetckw7+dvx4tsdbT/Lj9FMPLy8o4HDFEg2IAnWiNIUvKWTZBdrezOnGe
oX6rbORd/OGXxCJRe4mz9cwsyvc/wwaepk8dSr7CmQ6wFCzwgSyJkeahjzsdac+s/b23YYvVotjh
qrMEtKdhIRdLjTFaNdShGYAy0ROd91Lf7l9QuUAoNGZIkY7DH1U/CAQXPmtAKb8BOotfAuvZigeI
SBrILo5G3S3c8rE5RMUfo08auvqKe91YwRYVrjV5nRbxBICaG3pSCbUSxf1wjoBKidlxVwpBQbOw
1EyjOBROmCTxfbFj550bOg2w4a92LhLCK1rb9nlwqmO4xtJAQYFs3QeUqbJmemRmrh60bIvPuaz5
yzdmBHy55SidiZF93c3MgReQHRAfSNo9aRAdTnAQGDUdnlOYH3VKSYKKmEK9RZWMlyDY0YjVl0v4
TX1X34gxcNpwL/BY/SKZOSwcY7e0DRpkd/zm2CkeVdfLKcFD9DTUYb4/oZvFzXKPwXVoZZq2c8kr
VnxtIt4Z/rLiV+iXXXppPGvWWKOQHdWg4Ht0FQzv55BT8VGTFsNoCdrX73eWORKkeLJL++rLYHGl
IO0/fV5GxcOFOh9YHGYymCeNefhJv2JFAhT2dxaJjoQ+Of7ivqqjZWPlMvgVhSgoFsX1l8hrvQ6q
oBNgyo7yQI6adlgs5L1C++rc24emvThb/v1RmIglsIg0jEZ4uPPUKJXYKthLuXNL+X6J2GItTOkm
uCU/k/zOn359oN0KBcHBcccOnEHWUWlgx8cnSWP9pWQC7YLPn+/Wtrxqnlp2OotcJzd9K1Li8Ghb
+ybyY3yxq3TBb5fhLAFIaQaiI4Ge+kv+7eUbprHL2tO8OhQ7opJL/YCLMCf4H1gJaKSJhJaSJ1q8
fsG3aQTIfA0QodA3z7uLH/ocMJ6byUYKglb0bvFmIVo5xs1WN8nsV8KnGdMQ/5OGex07y1eSHqiD
Yp/gIHyNFURijCi2aGPChb9Gdv86uaVpETmVTMpy8tbrHLm5JhYGonbCIbKF0z/25YmJfH4KVWmH
YfOD+DdCD4PkGqabUYnAFowL1r5LpdX1l8GrMZQS+CZQv1DSTgRS31WdsRHKrS2FGTd1cZGB8mvZ
8scDJT5WE9XIEpTsEPOgHLmjEaRvqCDsLKwVKI/V8cs81H+hkl0lWmwFs1iFr5UoNmKKcuuyNh1e
FiHYBjlWxhPLhgC2Uryh9sONjm/iVFMjWIjhuCq4+z1KwWhm98AOX9DkbX+M61mRKv4xLpdejWyk
rQ/ZufhIWVc/cRxbB7m+S7rbTSN3mXqsY/Q3CdBDnIogjlnQSQBVnYPFzHe96RWJlS3C00vcm/QY
hH3SYXwKQrBp7dBUOdNxqSKs7wLuZfZeExIwRwZo5SUVQiSe76O7fHsQDt6v71IzZ+2+rQ7Mn+v8
gyDt3QOv9pkJl4ocLB4dACYg2Ryq+x33BkeSPyIC6YOdZ7TFnfMT1hQQJ0Ch/wbz/BPLBYyaYCc5
c23nF+BBenFsKQR9cRE6Q8pybGo7gBzF6oIUtMFU/NouTp06UYofzi4Qxtp9dT5CORir8o3E7LwZ
N4LrBwCNTVXoUfWvRYp4eOJrbmM6vW20MggIl1ufp4Dtc/xmNjQ4LT1q8PmdWmU9x0OSoJ7doFoM
d3elbEF9gpt1TIhaTiYC7TQoyNrcte5i3HrB+vNoHNeLQ4mT+gDvMNru5NdxDuqb1FcVlwo/JpNR
NjUCY12gAPzvj5ip1vQnXJ/rIttjwbNhbhuOue7K9kj2cV9jNIbgyMqbiHiavikt2aqTVXrJAt0b
ihXunjyPGUj/ApaKCEmHApik886mH4mSHscP0/PI6k4K3cdKAF1mtSrF/Cr8Mo7WXXw00Osb82Al
ia6LYVExPaeWr5o971fsAz3txfC36egzQvdSqf3YXH3p2UezGOLRQl6Llc4gFQQGaoR1/PVFK8qE
pV5I4OTqPvveF84Hu86sawfVbHw4Wzv1MiJlx9dteAUuu4j5vsg4xcJYFPD3yU9NBlaSAkHYjNMO
knxea1j2AV/GulKw5UpAUNfNUs2ub6m5Rx69ssiZ+IaMahom/QNFh5cVS5CfUhFWcoKz+S7Vh1sb
2CTVRqV2g8ba19xs+DadA6FqFXRhPRL0RBolop5cPUFO/oRx6oASwX5fUGiJjzlaUjFarerNL5Sd
4S51ig5SXn/S5BgnmoD0OjzO0wQ7ViRefXVe14SgItjdq/DqbIIYpTUfs2HNMUA6XZCD52J4x3PV
AW5UoP5t5ebm6I1C5egqmQwc+AMjxH13vAJ3McQDJh5j1lYfndEeCaMhi/Ogz1eLaQF1TTvBECn+
9dsfxfmH+JbBw2zA3sbAH821YFWp9yO5Ohg4gTH8p7+Hzl3aWQx5oJH+bWQG6dM6JvDNADz33FNF
eOhcJW5LNGp7rF9avN1IKltklJ/VhP+H/MDeVw1Huo8L9oPk8xWB8PGa2b4VwSDj6glyxsofveAB
1Bceq68ykGowbtPUIiPT1oUaaiD4ZLqgk6WqQZvDkiqbkLWM8HJai60kb7FwFXjMFROb6xdEHFfl
60TdJOLNPwmxtshUAbmb8DEDs4mqkVCucRKxVswWyGFSp3d+TCWlKcepI+azeiHxlj943j0HYrbm
A+m6cdZspXJlrEo6WZea1L5VHpIzsqPVTXlWxA2rGQlS2R6g3R5YJWdc4EE3P7BAdyDz/9B8bvPQ
lqC23+J1tkaRSMxp2NFX4NokIDu7qa35oHQlF7xrfA3oNUHVXP3CvteNdGTjVcFL9YRxB49edn4p
0vQDlx1n6+xqcd1WnX+24Csf7rAbq8t2ZwQkkYXwnL/QFB/3fEHhHIHDP52Kexh43oYX8qU09RbT
2eqSJbGZ/58++4jh1iBbm56U13933p73kDV7LT7gz/pOoJ/5CkarE8Mslu879YxgyOyyUXKxS3P2
aCGAUs1+EEvf5fk3D8uml/59aWY4TiXQ6hhJNRGm6slbuXK7Qd96/oefT/AqIWtnVDqc9+OnBxDG
c2P9Xr9/rtkcG+WgfOtNlk56ld24XpS/4aJWrJVaTdFZl/pk1+l+6z2fxp8oZN5NiBDcyY5eMkQE
Hh9XdcBJ6NAuvTHz83AuVW7qFfaK2yt+fXDOBd18MDPP4kQ7DHQNh2X7xojP1eiyGWfpfq0S2Hy9
V7c6nAPmo6EAdWSgbzeyHuIqob6OEU/8bbsEv3hv9wT+evJCz2KOC3z2Di4NbSatKNhH573LIkCr
45+dAcr/Qhl/QiG+Ex4iBaPuWDZ3s1jp44j3L43HlQsn0x1oJTJ3MnZA/KQzsnHIZtUIh16O/JkQ
+u3ji5WIkBYrRapHKyFhrtOPGwwUzaMmioopD8VbTlW8YiTCPKMUAWUywp6oeh+EhBOP7Bb2wZJ9
ZYw/qhcUC3CVTqhnub6tCPPNc0fSzLwZndsQok0D2r6kSXU6f4kze1bLrYw9pa2MUDIR9yWVAbGd
+0jBpmR6a49BhTan6V2AcrO0rttfaxBK4qVnfyUgdCI6NK+FrZ54b+gw44O/0MQRzd+FgZZuyRDK
W3fo7khbvauIPixOq1jKTeWRe3t8KqP+FCGiqtUAWxDEDdID8OebYbBXwZwnphE+v/IUCYuDm2oA
4i48A+TdkKNbN3+V9nO8wrdVzmkibhJTD9zM1C1cPvETvoQuiJPU9AsV1LO7odD4HCCzNU6QTfr9
c4QF7ujlaXHf1YVseE/H8sIQCy9mwCxmQ4V+8b2yS6vmRm736vYiDbcsnYa4qTTIV5Wzt7cLOYcv
UqtGx6rOjHpvjQ6ZsKNPxPUE4lHnL/UHE11LOlRNLnHcxx648gZ0tXrtk/T7t3wTjUExgvRDpiAA
bohqTBWwVgUhMqLB7UyzMRs4SZd1PskMobMsm6EDG0dfP0nczWp9aR8HCCjLHYtRMQLr426iJiD1
QPAJSeV0zDGKUehIB8GZzvRSik4I3SDzsQsIRsOS8xFXoZii1+5r/WHQtYiEqGeKIwAJ+87qjvL8
K1bu9f8sfdK85EXTuVtUfV3JuvvEDQz7RtaU0RkfSgyNyaAidJFzsvmZU/saaIV/KGa2aUrRl8ME
DpmSikr4ETjwYdqzF2T4LjyYsz4T+Uaj0EGIOh48AouHONGvmsm+vTyW5fyodzvEq7rxdnvrRlRy
vlznhyMrNOaWuiq/MesFR+nE5jyej4i93SBbpqdIHqADLEIe6Qm+V4o8XyCYqQl+NSwpUeyyswww
v6B+JrTmFAXGv5bcT3881hEmhztVlLah/1NC+jtEH+wEvP5tI7qRhQGCmQ8v6D5wknmjuWDGxdrl
NyvkrPxikTYxeUUOw34CZ5gI5MkDlw6bfxT5i4NtC8sMjp0x1HU/a8HeSmVB4NEy566wJxdUn+Hf
5wft+QvUfQwPXGzbK4Muapl6shkDVAVrs+WVxLIZAjtYlE4iRKE5dAbC3x2hJeBOyh16QvYJXAC+
DiHpaF/btPZBDDaxnrtNtlZjTM7LWjp24c61nl4UajwaZmFxzhyvZD8qLVwjN0a+/r4lxTInDMqc
k8CzEdZpW6AKh9R1B0OWbPqMg/KaQn+FCcpUdR5bfDY5YRY1C0o5fs01BttcxcViH8U2Ta48aA5I
F8N4gIszajB/D895AdBHIMI7H5RsU+Wh0/XcsHx9aHMiGS3s4xNd9nxLiEI6KGMUuuXolXjmCla2
1XWy4kPYTpitZE3Yiz62TL+HvVawVFYjiWu5L746JKARrYMN2y1T5lSxPYrv1MS0Z98DcXUVRdBC
o1+MbjofD5YuxrJTrdGsuqPR35qNYs2izXwu1iun/aQ+xAk3tg166Fw+pBIu1HcG9EdETaNHrz9c
SZVVz+OFKdOJ0Hzlh/fB/xBeh5nVQn6nS4xd7sUkkUr2EJXrBJj8UudHHRSH8tlnUvxH4d45S7nd
zimZp6a7UDftS2VS4npfCgukVx302bNxPLBExwFbRf2/rb8mCq1AEG6GGIjed4Tk6TrI2n+K75va
BaCS/oNFUYTUbOclw1zmJPGq+X6TJ4xx9J/DQfUatTinxFaxzp4oeyMckkTnIHeelHeRZATYwkZB
yfML3FWd1Q7fM10kifZKUXzhPZJg6ZgdTViapa36zUkJNivwdav+WISQrlcmbNXqUt3vbxSCPpUJ
rE+z8A9epF/nu4v+2lEDeHnTKIo0kKU38oSoMvle2PT29Qp4F1sXWLAM3yk79nf6TkQOpxqWxf33
FjnYDR6Zw1I0GQKtcGyEM1gIZusp8D5VYl2zy4veVx5HnI6shJcRmrOYWrIhtVOyBupF+kNtCaE5
c3cY1Ap5JrE1Wsin5yOX9YY1DlMrl/s8L8+b35AdVBG3BPhCqImq4e/8div8CEVhe+N4/6boiyTo
LSOZQ9eql/sTo/ZSC0/GVGQm9HzD04Wgv/C5quSVxqMJ0mYwVvZrkhlmoK0+ekBsPTcMuIPv+u9g
CHzJLdAK79QFC9DTBcfacXXFkch8wbTFniV7d3D1/HyVTuUMsAv/sfyQs0G+BDfXMyvYThr8qMxw
M18yHqSLpHaBKQkJBBW642EUeVkVSqj8OVOLAk5518m9fZ4GBpI4VlQ640g2+dDhzLBrjFLxR8Fm
H+L5AGUibT03KJ/AdI5Kq0APxSJ841kU4qikY1HkQTx4wPzK1HoSz/1pd5IqFv8Y556L4tcJH6sX
sqWPzm21jyphY8DK7JCRiMm+ICReBe+dzGdr9nWa6DxN/VIzSr/RtDFt+cktCPSLDHlg19w5JU2N
hCWnlM6jag+otu57NCi6yCdPKhS00L9ng2hFqIVbOY43UWFRIoNhrta47aboi+ALUpu605HcSn8d
ntYKc5yD2OxONYKNG6fOhY15SYXh4soX/rnNYW2vWMM1IHyYuhLZzlbHzxFowTYhJ78NgCRQuQwH
tHzd/fV1JXPQL0xZXmthGrjD95hK0CIRosarj9mY8GQhXaDnjAi2zfcf7IWpLdB0AZvvc+UxB9vf
ZaxlooFCWanDCua2+NBDTBBYF8vZpRpCeR/JjltcXU61h9W9Rkr2T1zt6RpPAQQhkhvV7AbIiTFJ
iLX10X2hUh03pTnjOrbkRr1WQ8/GT8Z8gVtd/KcWK0gImB4XBGnLres9dkwYAvBG92p8ss3stF8s
JZA8N9xP4HkcWVO8w6J47ddXHNoWbzKjsHcr3qXTYIaG90/xy/NdyoVD1PUudFl+btfjycM0USxl
ZT3LiL8+7ocvEol0HmT4iXmb+yKekGaLn1jAX2nGx06Hq/XkS4x6fcukCUShp6+fTZrxXsKaEa2S
drbExpl0PzTuVP4hunwpNKcvUcdVf5PzC/77msHoQ8ba6riac2dZrpZGpn5vZ5f0qAsQ+8VsVOvy
KW8XshPge0uP/YQMN/Z2/dmJ/ClT4ocAslw0kNxL8Jsh//PxVNlp5mdLQA0FY0wJaWXZXjB9Jb2F
z5RSz9eZwbLt12p1f1dEgQPXyqrWJQ8BDYhE56ONEX1zOq9l+yMus9QTYAK8nnuaqNQhXX0yoBbU
di995NfdoiCc+awnyWf5MwPhKP41Y2pdbwrxSWQwK/wk1MKW+WJaG70VkzbqpxJTKMQqiYZYF+aR
Z7r/k9ASVJgwk1KuAJqosKjjLyG92usvvLVuLIREfe006FuLyQ+L7d2A6Uml9D+m/GJy5srS+7et
cpx5eQwoT7ZzKJQJwYrb0KWYe2AKsF2ms8tyb0WlbsmtpsoCDtJJYLe2Dag7dwjKHqB6VLt7d5Lp
HefMwc4epYWbnE0ZCmW3coy/wYtogaXW0uEdqb6qguvIrL3JSqebWHqgJbedM8EZi2FGUsMs9CG/
yGl9Y3GiNIJK4HDNReYZ7bo9vic7Wn7kzE5Qpg4q16TjajWMFj9TRSgM4j1mJra8KYEzOSs/HwZd
G6lQ7WPn290jL22ji0zRv6iS6tcrGsp4AQM0c8rdRGHnyx7T3zDTKoaqy9iB9vIXzlcu0qivRrjO
YDfEqfrEUIZlsWpOSLgdMP6QSY84Yu78Giggrxgv0d8kcqGRYCuHTCI669i2btaChvZp/y8RloF8
CKRwpg78ACa3wv/gzLDHyi+cb0I+JZc82885wgNQF8DZflfzEzF+6m1EbIsT08iWcxayMLN6UUFS
3K4wpPfZJfH0XVY94L2lux4O57mf7/17g4dc502Cxytzt+i1n6loNxfzO8ffz8OD1lOQL7zt1A+v
4S+5TYIYuWWDokB7RKB7vvxwKND2pwEfI9cL/KhwfdPNTAthUziywdRi4FsgcAnf+dNe97/VOBlF
JoyYz2HgQbx32OUnIQa7M9sbHHjIGCpcFZjetNWweq8sWpFWL59JMgl+vrSWeqRnYOd/UAclfad4
WmjCtYm35EY8XiMa06gjEGapIirPTQVNNYnV7akVzBpdO94DxqtwGp+bfsyiVe3HEN3Jx6gHSsO3
CWuagxPh27n3CnvxxXKGWQEzimX3NfVIM+s/nYsRclol2R5d6aCz9ltSMWpb1bgDA4tWmXT6W+m5
sJOywN9xa51AQENulKNPXivdDt/XZz6Qm17D1MyyeYgYO4kc0GK6HVSp/r2jyUm/SfM6+IX/sSQ+
+cUup17pkGAl98U7/wpDPQaJavj4LXgCYJ/BrOw+1dcyqdM310c0ycVSAGq2PO9HjXiKlkjse+4K
5OD7GUuU2Cz7ZAIT9geGfKElLPC0pSb4RGM+k6EMUXxZrN4hVu7Y9Hs4gj1CrgRCVcHwzN5d/a2n
KBGsOQv/9BsNRg57QS5TmZYxifwQma6kROyDEC6qrdHwRAPW7W/k6Gx53K921Zy0boyC6bJ6tx3o
mAOR5zcjSQANb0MlgkTzeWBLwoNxzbWwRcYT95MEyDv/MDqEMEYQ+fP5I9bsPCK4Qre13yB+hqwH
XJ6nHvVszhNvnkGjOsHIrMR1Bgv/1H9qAlHGrNSeZe11vMdTCzanB8J/WFZ79EANEqKbdxulg9Gl
2EOKKLbTf2W9zT2YLzLbdJlsN0eoV2uBAwFRcAwQdg7NjCCCc7FMg3tObg9WSl9EKu3h3nzE1+E2
7H7oQAAhY4h6E+lBMqV29IMizyY6Ii8cQGfg3Zii93Eq2FUYKuI8BQeaIE9EtijEkvu1CVJ6svgz
lC8pth7ymbChRNY5S0PG3/2FyGW9HgZ2GcGz3heylJuRIdJZDzjjnBL+Cj1F0dvO1Gm4vFeS6pWC
iGRZh2bdZ1sEyJRmHxXFSzsR8AaN5h25U85g+dCZFIi1xTjnIXlkUgbtjuURa0QYMJ3Jn6k9DlTS
5e0eQekAO7VFC5VEjf51q9IgioC5KwVD9YZu8l9X4s4jsm6rJYEG7QUXbX3vZNCJFAyKmFGC3Quw
Al2izx2WqT2pjrG4vhRKelmwTcvY8PAuDL32Dzv83nvyHKiTQ75OgNYakZmVWlZXFyOzqPr7QNwm
Saq2plg9oQx8RuRKa3Am8kdQIhuFWxxqtUBmFzee7GAXYa7rU+wG7toyQfQl2zkR5DuWgSdzUAMu
eyFrVSMlsFqzPPuSDwzGQEtNBa3u+Tj7zO2aZdeEIpsFgPpr0WXNyNdwmQAXWwqyX9LV3Nil5mW8
SK+Y5Inx9vCf1qU6RKUVQBxpfWj/mC/YYa24+u5Xv+mUuT2BwJ5ZJCALhKYgmsNgpI/Bx7rNZnm4
MW4Xf0YNOQ1aQeQmagQooS6CBzcbpCw4ln1/A/UUQIl1fxj0gyHSc/ukExSK8LFmqKAMV53xdESY
Ebv6J5oDRWLTDVflTiaT4gpq1R2gqdjVdlL/UbRlhzc6MmQQSxsm7Z4BL6uSViLxbC+MfjYBqoVL
4LwQ7US/vPqKFSCjG0O0TMCaEXfG01VDd6vOB95qjdik69jFsRovKdKFxspYTWRdCUb6PlA3KtHS
KAi7n8NUXYenXh9ENQ4GCtE6s7RtQ+SHez5JI0MvN82t6nB2+vzwl8OQlct4wcR6iBdP4ljpe1KG
RhzC0P70MGK4ys1+zJHsPSaaixSQhwgt0QaWSMPfShE3nwaxuqY0vzY6xXgwxSRFzbLgff+YYGqz
pQrPX9NjW9ObrrHRTOAa9FPhuuxYq+563is/vCZztZ6rvvR+wMnoVheHWqgRIWs7ZvbSJrgcbDr6
qSmbsQqcSO54wOeBL/C+4OTJe3dj612ThWaTylOphbdwrQOYhOKVIFmf5gBANXvk4lQbNlYDXfZ5
xSORtXDK9eGFyQIvTv+w+DVQWuC8/lfnK3+8S+37aIGE0txyjO/ZBreU8+gpQIhrBX2ZNwEvZzu4
KdLUvAe5SEwKC5N9eZSyK5ntN756AYOx0dWuuC88g/NLcr+UmklwP3Hz+DT1w0b9f6yXTOgdHbOv
nNu+9YmHFZfOtbtNQl17tij4u/XmICC+dmJPjgM/zM5w8IDQ7rmDFQd16ZIcgkPOLBZwmB8giVGj
ClVm/GH6dZT2TnLN6GNfsb2XbNZQEttZMYevYHKWewt20TcCmqp4L+Nrox/ButoLfrO2MtfapTzG
u3FSwipKOdu3sXurz8X2pufkfn74W7D3hbKsK9phnyhqOR4EYgGT0IgbrpQ+xQaAHJdFNEqyx04l
1Yd3QidgFsfxp4KRX2B1mxbZkBQJNV2LGVNQbmr6A3luiYC/F5/KTUnuoqonf6HHR6pjJPbLMuZu
quOR5/LwQlkEkowKz5CQBWMyRLn1zIE76i9a+B2sGCHyLmDnZfEP45ofFL+JolAlS1ROXh9A5Q9B
edZM8RPRWxHI5hqfxtfzJykX0ITA3A0Ctz18LI6Telk1azrQNVixwDtdWRf3gnGJ1LLJe7/g+00H
f1BF2vxWCEx741p1W1iMzLMlNtD5X8IU3sjZc33b+woze7fPm70xsE44H5r0d+6g8qRMWz3zZS6H
VkN0f/2gWkSszUvCRdgN0TFC82/r3i5hD3kEDYpF5jWQUpvVA2LyAXhKPus7rGlJUw8KCz6WAlgR
xJJvQB/LjP92f+vMEXj0GEAnydJZi62NVXzAZqAyypBlX3Cbs4mUuaXoaSo5gMX0bbCJWICYIobE
3K7+BaFQeFUBpeb553TKZoW5E7PeRuVJjgvsD83ifujI0Y8vM33j+dcJ6KS2Btzp909ik1SjeQYX
+5P4Pb5JTqMLMPBufYO/YDt0NZGgEqis7KQ8Kw+Av13WB8//mSV+rPxU0PCZujpD5dA0ApnrrCVZ
p23VNQMXWqz+cCNKVoIN+xWT0/lYz3dTLBwg9R5x9C0U8BO2N8N2MMIPNSLx05tzSW+cDmsRA37I
Gf4TnaMjHKzuSpFdNPWMIieaiQIRqCt+PHT++OE+R4VJHT+lsa12vNaV66mcCd9Yqv3h8n9Azu9U
wEs7FpQxajXQP7TmHBIkMkOKxFRDDoL8K1eQrxzXYA5Au0gPETVMDh25LZqmmO3t/THFgWunXSXQ
GjuhN5EsAVDoiSen5mAbw5rvSZCfN99LN9J73pQkcx8usn7gH2sNeeODr21mVUUwOs6rvu+ZqR0k
yRXW59oSzuoN0Kzag+ddbm7CxzM4ca2Wanok9ziulV2r19zlLnMTR2JCHqe/+xkYZ0cIra7L9dVt
z1rxv2MgBtNVc4xfKKGaJs2gjE6tU2iGC9lprFvViSQZDB7SRSfWfSl2CRaacR6ZHoeJS+3CLPGk
Pjyze+pmB/BTH58DkKSutXZFjtmiSnIUVe7DGaAHzSTm8pjf4YXOGSx8o6jyIQBo8/iYwssXNCRS
UWS1cucEeQ6A3GoMhaLjzJhRq2HiH6WI9vdbNuANr08riVVIY8HDYDQ1sOzGV3Txcd8EPuV5w7ja
MyeQhHUC4Tf3rJHEteXUKwtliq15nOD55vyLLixY+gtzOjl9KK/PVUSjXa6kNTJGFP3Ns4xt2I7K
h05toa3aZBoAaEdM3+5otb8URVGobVnGEfwTINHiFHgP5zMPIopeFHE6d2PtDc+SP4RtKcXU5EZ1
eyq8FdSu5I6uep8B/A1HtbvZldkwlDf4HmgqNJq6V8k045IJuw5WNvxt5CbnefhCJKTBVi2uIoj9
A1S2WIRfcSsPpE+So5y4SFeZH6JYLIWzxt9/CzsuNqagyFvWuEBVqwdEWscygZ5tWfU8vSfg4VoX
Or6v0+f1KLIMShumq5ZZZdZ6WMEWQhuQAlJ9bHF8b2zzIC3pd6OjD90fc2kd6Z4bmQMfk0pRYa6t
oIsubjudFohmDFuzEQ8IV6jw4tU8Sjf1Dyn+q31nomRI2aBDCdKRFssV7eFyuLvxssABgxHBySwf
2wc/RyPI+hB+bq1yQWfe6jVMj6QqNSWLYKFHf2wTUck9u/FZxs7SjPXbFg4XfDCRw4KB8ggwXzZQ
qmyL98aGLDB83Ge/CcZ6GMjXBbPNp2N7sXkxdm2GnKOdjj24pdGdIUaSOmBKS+ZpJSo6ZNa2fnVQ
qEEPVJGcDkvVF0kJuZAy4EX85K156NplFWfBQz5QbM6isCv4qxL2isByCGzZIRblLNPR/6ovGyEl
hapihOlrDiR8ZZM17ekuwqcS6GgCUEXRc32ivRLEWTXqvBRfSo7S3PPI+E/rDY5ROcT5gyoIWp4t
Omwn+NZH5Hx5ahQ9Lrc+00JlrxlDgiBiW+xis7+1tpyRdAfTOz27lO757N6MOdAaavAr6b72tKgJ
NMXOhGvgBXNjSKrEX+yHv8We+DcFUkYS0m1MyIidnL1QTbAeb+uron8nT6e7m6YL5+i+0H64XUeM
usUBC0gyXbxuB4EU46G0RonBmtDJt63daqs5p1jo48FzBxHKIomlUnSzt6SbPsNhJt7tTsDgyQ8L
x0JR7mU9VRqf+W9Yv5MQbUHHw2kARSK36dfaqT7QRVS1OTK0GK7g31xOy+KZNjGpxkfaZ9J5n/Kf
OGyi7Zmmt//oed6apr2A04kThLHzU+NK4E4WUMC1vOxcaXHYIq1vTq7/Cn2JetgLbwtUlo9H/dg2
V5tJwG/gEFPLZxbLoEXIF9LYZ39g6TAwhDdGYp1ob5gCKGsJ4Ci1UcusCX6MTQFjqeQD3OqkfxR4
NcOLI8z9fFa0kDKdi2XrKWfL1+/aHJ8/VdReQBcO/4ve9Kl3AZF/NOXnIpQar/BUz/vFk9ZiEgZK
8MHdYoUJzdhuZ22w7IeDgL5GT2ZVbdxg5aGiu3v5GHcjsn1Xx74lnqSvlBZ3NXYTXRuRXns04nNT
V+9GLyKT0SD8OHvNLBHDUAHx2WotNovSxyHGkADagAjE5zBaZTbpxf9VhKK/yl19jStkTAWRqupe
gLqPLQ2WR7mxMrZYmG2ybc9M2e9TixAETIk0IYhgVTKLbj8rlKksRuZ6I4sNg3FuxhU4CYHs3324
ifDyqQKP/3k3KS2EZBOC9GvKl84PRUMo3O0drKqVL+LJk+Wh+FihAaa9TOU4+/QE+dFydhTZ2/Qt
bfb4BFStD4EvMUwuIoeStshxllY+R0J5Otwhqan//yOsp3NzdgqIhLfjnfQhu6rAPEMw3LEfD+ky
Na8gTSwM9VpGdmQDMkQTTdsuAqYxAV9sVCW88uEet3TAgCzYB3YrPv4B4UaF4CuqVV8LGiN2Yc5O
1DOvTq1ucnMlJ/j7A8NaeKazHl+RA5PbxLxJVhPwrqX9v+dwPW9JDHxat/vj48myjjIG3ikLZAYH
i9SxQqdgq0ReW4CtTdQJdmuzWwZuD5ggWvfcqIndcDUoV2DSwfHCsqQ0mEimPUmRW9g1KzO2Kc2O
TQKO7Ujah/eBldQGmgOD+2KYWHQl5ibss0Gi4FHGdy4m6txqmIhCOKp1Yez79Crvpqla+QQ77nVk
AYM9eUP3TkEzeMus6yl0u0hxYWeRJb/CyBnm/7TpZiTZEfJqoI/zeSzWw2H2+fojF7flIilAljKo
tW4v3Ev9LgDY1P76+M7p/M5bRPYGXczU7wwLCmHalpAbrNkRky7vSECC+osIDa3RromvcwTT57tV
IhA7fReWh4WhNM1SvLDryPdWmZdfhihrWqoWbIcL+i0PB3/BtZ1LK9Xh67catHYDjCuWVIojSMlw
9fLz5j9ym6dMluLonw1nKJq6zd6GaXVVMR/2v3Kz/k1aYeyY2TbZp5NKzky8MoGDLolSgQ/klV+D
tkmkfvgvqQVXtNR63cU33EbTHQbdyHPyA5BA/RZAcdsk1AqVr67hrAjg3FMJZqedGlX+W2sg9pK1
JPoAQiTDhVMjRc8SwcDLlVh7w9GnCHbx5KM/AZoRabE5lclFUzalsyLKWwMYKIkQEycZczhQsh6x
nxCiK67aZeYznN42bux+Jf2822psvIl976Oy3oi3TTFFd85yOVZ5+kHbuwXaKV3veKHZ+ZG05tj/
qyNfBEzsFeeNfs6ZDNK3nwllWV+iptjU+UDij7rN0wByw+uzgRlf0hi5YE/jVMI+rUzY1bPTtQ2L
QB7MDxZs7rUQ300FrLb6/c4d31pQB+RKS3v/1CTXV3l0CtqagmY5J2CYcDFW4GzebvcX2ZZ62BuM
386NWMiF6rkugwGpyQ2jbRt6gFlC8KNMq6yPhK3C3/f0b+DhHVhdacD1QE+94eq7AeNR71D+YRiv
TRUfMK89Us6DtMsL/55N97EjOwlgQoUSPgoGe45sJEjZfc+7O8uiUT3RiFg4DqEnXO4RhbjY5RPW
Wvu3xQOZLGcDJFUtxqQDM4ijoY+lXI2lQNvzxBl1XGZKGPodcffpTa1eP9GOUUgozcokGTjUK1Ep
ymfdrwWXXzepGykV8aLJzXuS9sigSRKeEP5KtVgsnQi3a+QSLf84Y2QLARbnvXpDxTPzb7pILP8b
MOE/DhBV7f63ZM2+CrGb0iISlL/jjZhVyWir6rcjc/F3g4Nj8V3YUEsQqLKSiSQjfk/p/EJGNki4
D4IVdNLnnYCcp84piO8TEcFRslY9M0Rn58Y1/0LOd2kf9vqeSiXfvgWT+nk8CZju8dbMuqPzwqZf
09OLqMoWmkF4fSiMxENryoabQfB3LU4i9qbUkXnO40WKwUpIDQbcEt7QPtmc6GDs173ovgTrCAQ7
9iedcaN0g7btbbxv0lFV3gxS8ZdPl3159WNx804OBHCdXVwwqwA1Rz67Y3vOcw7S8qkfpxlghToO
iFLX70GslvuOJz/iiaiGG7UNDsVG9H9QkLOjMljHunMY3lhJMzheghpYVJNX00aLtEQ9sCz0KZ3c
bFClQ0l8K5bD8a9eoiuX6kCuI1XqvgqCGI6p8hEoj6+Nsbpn9v9Ys0rnSuoqa5QXptde7QsK9abr
yZYK8MOcXk7jpur0MbR6q8esMypporHS0NiZLSQr3aPUqawPL0C1Kl0yhT0S+v9Yy3aH/bW03AbE
A6Dklq97mOYkkupq4vwpIyVrJmjrP6dEWjoSOu9WJ/hxcsJ5ZVgFUDak4hrjqdAtQy9Dzos4QwgG
XvyDdLWiQVunZAYDHRfTAMoaIAev6XREt3R6Nvt/hht3nx3mQeo2Q6crXrGjOQzZvEiuhIv9Ljqa
QoCmDxcgcAO6xwDrUg9uB7QNMaZ4zLIWYQcz6+el7QHHla6mHy196KfuydNWgOFsRiLbfL8xJCbI
ZRgDuybdBVTnFQiK7i+V5QThICOGyHi0VRDH+0MQr/m4LKDLXL1yzcDyPeRnIQSRgKhKKnA9Ec4D
jdvb4KqzbAJcGLM8lQdfud/jRZrH5UQh64FZcIzYpx7kMZnbfB/jwb/JgMg4KkQ1BqeWmoKVvQag
Fq2IxBiplGAwa2GORbSnG8+B+0D/KiBWgCyjazoiLZ0gTGrzJpUBcpH/V5doST5RIXQ1+DSlxQTg
FIUE2cW1KDx4c+vMZH5q/RP4HgwzrICEfUdJudk9auRTTsRrvFcOrDP13ojPfn6RNEh/Kyx0Xu5o
iGRTPMgco5wmRdzlAdrSmmgwBVnWwtxvnlQH8MihrKhgBN4FCXuLfj3sBwJL4UqF7zA4KDkNmhOB
F2U1BV8HwEoMnb+llWuo1Gxy9vhNkNNo0JinYGwsEotEN16NM6jZ8DJev/bkOkyCywdiaDmLO15J
ZjfzghVHlfLYr0KLU4DNhg8AWvr5AzKS3w7XoCF7HrWmJ3F7ID0ILZjfKSamxyA8klQjpFLYMe8v
9ytrLQVNj9EAYj641jD5PS9M5FRFcdj050VkJEJUpi/yQfKYUOi84+CyI/sewvPfNiB1Hp7V4gBS
ejXlYn9vpA6LsPpA/GXYVxnWNeoBjHY+PqIIm9TS46KJeasACcTrB6IDK3xd6OTFgy1mNK8r6OVu
T3xLC3LPC6tvonBjwGEA6GMpSFJSZYluC6WtzCaOMlcMV4AEyjrCf0kbBypljTnUvF23oIZwJPXK
rpX0YW3mmVUmv+4BALPrv1KGv5aazgY78BwLNYmN4Utx5sGTC5B3xuG03XtqHPuZUDSt+u1ZOM57
hMx97nQVXQyGZEtsIXeVgQGXlegQPgRZfZCeWg+dLK18rva9IM3836eykrOpFrU1iUDbsU4oKwYA
bP8zQ4ivkisBtnHql8MJHAWw8r+yAWxANG3M2lfBytEwdqFnap1me97iuX4DO3F/W3zh4PaM/uVO
tSCvAt5/ZVRwxulzDZgOPWecb0CDggS2tVSIlKasTrtAQ6ux3zwtbKRJ0ZMohEQ2vGkof1tVwQ6X
upOHQCi3goea+9l8Nn5PEJ1ntJjHZOsIt8BdssYoDPpF4YLuJGdlgwLZS/PNzoE9XsGX8rdyusAk
a5CjPJMj+0fwjr5lzCw+SKeSB9JtFTQQTWspzn3c9DXFBduZFmZW0WM1098DrEtkG6Ffu5Ln27ST
eKWNV6U6WkWlEHlcPRb6nyzfn0mMd0ygeuaXRKAN25RNBZx8kj0MOHsDczHz4/HwHKYE7sYQ5c9U
lCjLlkJ0q9AQr7Z7lkvCDN4aiW8qqeEaeGiTVuOwPHKY1+/BjqT+fcu9N0pnSTAXSCxz6ORImyg2
sYNKksSK8tNRjy78Qd98GHmgSTbULHyG7fpSTLGCnysEs0VCbLHUVdgU7uaL1uhuPBtbU4VYQFte
ynsmcIYUYvtyJQwB/h90TVnKBN0BkRb/wHiw2ffouDM7WOjpORQ8toJ+j2wQjNGk4ph6aVxNjkF2
zSJbXewLZQolbzgYvaWNoYZcQImLDUYLG53aJ3xAxza0lie5GB3fiTpxedeRiWrSTHLdMmO1Ri8R
WXeNXvHtstzPC0v6n5uKSEDQ056nuvUydfAfakAuQDk5qBVp+W+h8n0O+l5CTecqr6EsaduaHJyq
mvSq8s2QfJCGIfB4SSnvjoDnfXS5S+lvJCfq69Ofd+pWeKrBzcyoEva2uoRZGUFOxcFMgo7Gn/hQ
KLQRqrBZ0/9Jm0DjLCY2cMcU6GTEq8NNwusWWKA1lZC3U0G4h5iHpgnBrJBfQKxe2YeCpV40HYKh
ucGvB9Nd75pOekfgqtKnmhLKX8GARh0pxzR6kHyw3Mq4bRwXq8hsQR2kkjuZzEY39Or5OA0oIyLS
sR7/l5xqCAYWLyKFa97qteAbv/L7UlAxiMsWsSmmw4CEXHv7wKTFJIOxIWWufbuE+cjE2btXMlgU
ddalVVmHe+Dt2beLwjt4nrfmoevm/qzZT+f/ub1If8zGKKH59gSHjAlq+Bjea2IoK4N/zI++upE2
0hyI0ml8/Og+odS9rNAjcuw+eAxvdtiXKykJ4gZFLsDW2q4pzijAWxSnJ5Gn0hi1SH9fzgGujYJs
sjH+plNtLBsJMG7fguMfyBKahdLXYsh4QcfnLmqr4co4/Ue+8xzqum78ZDI/OZ0VBwX1E0UA8H9o
ynKmwNYXmgEWGX+Vgk1lTW/zbRmASs20y6JwF/OfHcx03gsPDkZ8lX4AvbqosGXYRgUkYKxnWAdX
RFRM1N10zgQJoLDy2ZXnj0aaQ7rQHVuLD9YEiHV1C3xTqovIF5+JCN+J5aDvIyCSfdbcYq6c25HI
uWY9AfjOBaZFwamYaPxkSwymraAUwQoLhxYJ9kf2XY0o0SiB8vTaOgt1Wc74GjltkXZY2kachM6D
yL8xDUepdzYyoQoX7rCtTrESmMw6fYbQj9RyvW4yBpVrhGKMopkgAwm2JWV/4o8/CRGL9dByHk2H
utM36abhn5WvErSdf5NTSlVsQViGsMedG74CEwdahHpgLr4LFFzK5LVF2x6566zbs/sb1g2vW0w+
V32sCF9yDHEHNSMxrMTfOfQ+z74w4xfyMorDxRci61uD8chKklMv38Z7khf5O3P7I4DfiWcTyRi5
zj8abKYg/nGg4IF/cncZVdsCdWKL0b/9wkKgezRCaiVcg4VIHDf2UKyz8+Cy0VKD4OGMA10xQux4
dNw0WTnLFdqhyJ+/CR6f5X1ZqE9xt/5+Twof2zNGk69tDE1UNmR16B1uYFPKpvq94UkcOnQpDv2L
IChits2FtUMyXPnXx+3bHTvbCl+h4qLe6z8T/DAWXxaFoOCSVuwGMz64Zj+ybOFGvXTfCcqFQ29I
5McIX5ZIF/rvbZpFlj1SFZbF37v7n/wK29qqRzZoyXwqn65NWo/nWt41yPRQ6zS2fx5JlzvOQvCQ
I4eNsvuz4GCljUItWNAnXiNkfvR8vwJdPcVnBGo3bo6Q9qONgZR+gdPWa8tpsH6PwKDZAyeICInQ
DU3jS4IxziVARUsNEFNXhFPSMNWL5/FRALtWN8SNOEjIJxJcABBwqT31vSvN8xe8cs4+Nct2lbDM
LL1+1rs15Z2G+wwBkTldFptt3Wy+/NeLit5klyEPtiDh5EY5eMlBvfEU0ey3yJPf/WW+PmAeC8yY
dpXSPFUO/LPrwF+dxTsz+1C66g7JgJi7o0V4GCp5seDGWAucaCbLisHLxkuD8LgKhdtlMJLzr9Fv
Kce5DD4sZQor2Ghz08hZNq5sO7pzkKnK2zuYJWDZXEPRNZTNzew9oOGRcTwOczKYBnEjF/2vF4oi
uvcXxqw+tVZPUoUBAj0W21E+ZDgDF5DNLMKLImJGDlLqmGg2z2hAynVoIhuQOy67M8K4rkAzNCqL
StHO+JGX7ihRmNswjTihPBeKjghsT1eEPue6oNkLFwY4+OG08g+eJEP+78MKtNLVr+GxKE592TPv
PeVc1+owTQzRoMeQ02idfsOT4SWxO37WhRTnJv7tYDmHHZZqgi8R3AAJkiCvP0G1jB3FaKqbGcJA
5uMMmPb7d4rRjwuMH9AkNSAhLNJjOs5Cyv8nV9YcJkcb9VGtyTKEUxLykTXHOgGsYYYZ3UiMEjd8
wr3j9D/ddgL/kgms9oa6ONRB/NShGhAkFbbRJDthEKstpVW3sql4snXwMwX00RUCnFRnN6Xwxe4Q
OGVGdN/PFtHa7fmhDnAaL7QLIZ5AJunInjJOiPLGXq61GdMAQFDKtuZjYX0MjMmG65vBhWv63fcH
EAx9TFoYwrsuf9rBQvjfFiUnWa9wbzu91bKBlcCUmjaLWOP1llAXVFx0nVWyxfWGv6Vm3qr+WOFw
yRtAbKvitSttFgDoKim/55kxkW4Et4dwTjirkPh+gto/lX+aO2QdLm5MsTL2+PX03zVOVFMyxeOO
28Y2SDcyiIlbBxjbU9xq+RwsoF7KJN/dL3O9Mw7w9U0NfL7iZMVOSLbZrcFMGzHPB68bBaKFBQdp
bnmceRgh+6ia+l27Igjr8jWJKH7uMS+t8OKU803LnGDoB81TUZw4O3KUyuLyeWd38t2vVfQOgjvr
roVkELaztiWK73e73u3yKjP6Rn7pmeNN4/puQDwQKizD2MDspYk59eh7/JzRnqk3nUHXgjLRYpw6
oWgKPqEeqckWq5ctDXsF1yrI/M+cytv7TSV9SZjbWOUFAt8iQ4eDn166QnJj6bIb6lMZeMZ7/pS4
zQOZkyZMbJOaAFqFde8CAEyGeBLvgAJj7s0hyq/x7olFNAIVG92ZF6uZsiKOmCAtcb1KkQhCzM24
d5Ncu02NjvBpa6ZJcW0mMybdECbqbuEHFHY2bXYLvVW5XEE+M4e3+FgjBlTz9hHHRZIoM28sV1bW
r3PR4dHVtgZG+jMlpDTiHLYSVgmdqhdyY9vTHdEy4Zhp9Fe87vTAbNnpCNoKS0ApdSr8wK7iC6ZI
rKY8M+8zaSRBaDJ0jGm3k2YidNPQZgmqoE+NUrpa34hrOZ5BYfyiudN9N8cTb1mT3I0ID9QqK6Va
lV59az85KScR1eDIN3INiwiiFz6zRqZxhN6g3okTW+riaLZiHvLMmbci9oAvOUX5lw3DRvKwEK2Q
qJ/iXq17b+45Io4LP/koWZdaf0mPDZzU1lyujy9G8T/YbSyU2EFjrPCgGvm8ERTX/oKRiW/zzHec
PKnT56adOkbgscyTGEsFkVwNKR/dI4vlSwiMlEvLGcELyNhPskYNTpmotboF/mLvlorOf5Msw80a
ZFtpk7luogOWM6Ff1zqivKGmR7zDkvepWwdDIp7BOKYiNe9HiCozwRmLk4fOuykzkoyDg413L9Ux
j+8d0XFDDie4YToqoe3VWt45XZ74n3gDgRassmsvVkULG5WGq4ndhait/Is8Ve8muMedC8flk/7y
aGtoFr2DmMxUOMxh8oDqc9++fOceE9ga5YukI7DXxlY/SWkGhkdpYnFwRFaOcDB0LCrC4FksO5Cc
rlwAwgHDLzFA8VaVE2B3R6eANzOST9tF+zXUJP7RF86orLw5lqZirLo6IKzR9WymU3q5WhLJ7Yev
2FrvT8kNVkFhWPjjPctOhiTE1u2WA1BzKKzkJiiG4jGWiPnoDqh7Pn7HufKa4oKSUCEkBFpSKKwt
7NxwTVC+ShkX3DJEAKKi01uyDJ2hodKONQnVoaNu1SLJGEB6tYUvPCvoj1KIemnsiz9w0PpYmmVh
D3xoulCs0ucFK4Nf4lX5a8+DfWaPBD5yIp/eyosS0EDDVg2h8i8hbyjPMdEqhX6RfZgi9xx09bGZ
4R9nkCni7mEizeLUIqqX+LIcbX9FMLnNZ5oxZulqOeH1P+0TyUkjxRwnCtRblAv5Rq63eIeyXId0
kFYYMqnwx3+f1L44vcubXaGYGCNryEwtQaREIJV219pmRtQa/n4xMKBMXU7Kc8fG8/j3g9M5h7OB
9SQ3Mfg7ZST2L1KOkZRUkLbF8BUYbyUJQwz4BTE4t78nizuaBiyghK31qQNCJKK2ODZVoCOc0ZF/
nSeEEs370utQdeJoBuHuHrTPE6Lp/aKu6NzfKe6jKvMiaFnlgUZyMNuRHQWOiDncmTP0aEzLpjD1
rIRMzvJMZcOu7wes71qaSoQtYYvM63/gKBiQnmBbCh9CfSk5wcjtkw9cEcVTjTpGyo/H8uOvuhcL
1Iia+RYe9H9FSnwOMfi5LMwiodk7mmwN7Uwgvsfj7QKGXg/iwzUTFcwKiihku5H0N67E50DZ0eNA
PRX/wzAAH6Ui+Jj/EP9SwgYOdTO+vvpzbOgZTGElZg2XdNZPIIXZ37TJUc2Y7R+DK5bp1W5UjM+X
C0xaqOcWsVHokci41JUfLMdOXPpVeYV+/lKmzb1C06MUiJI13PxTnGNlcE8E0sAhUlG4uSPofY9n
a0epi2OEPPhoyHEozwi74Y7GxAeJ9TCvmsk6NDqTye8agre0cDcxKBo+mQbtai4Y8n5yuqzpxaxv
mv3q+tFqtRuQwFM4eGuuiaCrM1LLhBfKpgCvyIYI8BirLEezViMBJEuCx3vg5AdMX1YIuClYb1qr
4jWyOZThw7HG56HIwDNvG120/Qqd1pniV/ts4l0iq1G8RWzHPKKcB57FoxfAgAqbO+++rYpXjVRj
Krez4YyPrAA6x4Zuk+wn7ypleN4DmWIWdKEHGZ+cdWO8+oVjEeKcSxPtGvvOMEeZMc/xcMQrv+RM
Uhew6188CoHzFWC6uo56/rn67F4rdcyn6yHbuO3S2972ZzeqY+w6vzSY79q/yXU79qjrk7RRuHE7
Gw4wq1repQ6IXGiXkleCcXHxAugJCeHmZLkwrQn9NMtNuDJ6ZHUCLl0Jx2lreMHYYb7MPFktZJu6
OAgdCro0gHPoTrKAye95c1ezEPjivFXgGNNjHenvbg6X+m3dDau4ety9mt21pkGktdR69mm+Qm+4
GFhXC+mpAJGN6CizJqjfs0zwebKpSodTs0UjrBv3Xb5z9ZqYNL+h+gFiGP3e+ue/rqttwXm/QVZ+
zoCKlamrNWy0xwfIxiavUcgyPj9QWJHhwHDo9xNtC7WRAgZ/dHWjvT/hNXbQ+3/N6/090FZCxSGY
hWFsXwM9joc7GF++mb/JBTJtZThnYPmGmRdgCjxpbx6zy50OGwCh9iuc8ACdM4eD48iu/qU/nWkO
8AOllv6ADtegN30lh+l6aKlE6pW8Hc5hGosgsWtVkJ5xleENfBfX6iwyDVaMbqiyUJxMiym/AQuX
uAbRTXMA9RAAU0eN0rzeS3Tck3s/1lxs8FZ1bW6M8wLOIFwYKgOB+rnInX4zN7FreoB2wXWCz1R7
/j8qRnwbkI1ls8gdcYA4mA7gfReHI9E9VQnp8t0Q8HD4YsYqh2zNidyvNkyczr+RFu+/xSsC8Ve9
9u3kdYTluCjSvndAVH4jgJ7R8rhOGRaQ+oxczp9XNUXPp+wMlZz69hHBC70Vap8oN5FINXIl2Ty6
NsY8+RTEqUmnJasgRx+7VvSnIXAoqRoVEQQkVhCoxPBb+4JotIzP1hricpqi0yFyoc/zgOExPF5t
9szEvo/ETdo+l+CFrPa3hh/7PbKYHVzAwZ/EGwVABubd68SFUnGd9q+FQMvJ5wkGmIhV9vdA6E2A
vnf6t8neAZBEAIfIPnzr+w2buUrm0Bucvpg6u0QsDZVa8Oj6vm0u+LbmIF7j2o9+N1P0sD/7fT9/
dvZB6jcSKx11+fogSz1MFPzksdHJMPneVC6X/fxr8SaDdzkGu0/COHI0Y10IGfw9XcAeqfCcg/py
YIBMreS0MttNvPdy4XMXh8sSP9gr2aSEjBrfvn3BdS5wOQlxxmB5Dc0Dt9JBR3b0/2hlbSKcQkAB
IMkYE5bdhZ9mN1UlxErsh68OYIaCwQ0aCrWSjQqR00jYb3g7BLDYtJGDAHcfAdfCd/YKRaJ2sBdV
ZFvc/uXU4ui1WDnRChX70fmElgTDSLnPSmc3m8DbRbdiVETmjZJAXCAsAnKmEkXKyNXuga3IXWmD
6f0WtxNqMG1Xyakcyohk0RWBiOXzxDvEut3zU9UxR25CcgTt23Yq63WL4rlxIO7L4B17IqXruzLS
gXmOMcQSD/auzAUq1WNHO8emzlXYjFeGyuyD7U32eNxR/siNopShfhdYDvJ9/J7B9HUfgl0HePFw
TuublUo7/gPes07FEJrFbjT+GHY2Yrbd6lUH6/Pyy9HQDtoyIYJMVT536dEmTtjnMpwI+TQQ1WnE
D0CEc95eWzIdZKpcFFlnx3+twH6XK7WT5CJL12BdQjCwvmabgjW1W4dm3TdfMt05zMVHNPfBeoFM
Ws3xHYP/O13zgzig1QRzVxl/DhJUb3azyQfw0b+XWJigPH6GTyALdvSzYy1kTwz8qqS+avwA35yH
BgPmbdll5P+aNTkPdamVWHMCvWFDsHuYuvT9ewmJcIGpux59SA1VcDOPn2yMjCfQ+QVQrUjspSPx
/QYVYO8HVHu09U6JjhHla/vMfV0FxcHV31kvQ7GdFblLK95TOU2jzn65/ZNfq5d+g1V285ZJmLrL
fpfADEeY78SULZIBAoSX+SlXjOouK03LL/d2gY2upaxpsXo1igVbwYFIvkjWHvig2yUrgG2jSIm1
Cx6Wc5JPUILRjI8pFMVxGNJHEFV3dMsw5/cHuwT1UsI27ZJ91tJz2fdQXZ05Jjw0j4YPDgzA5Jt7
3PwQvjp+Oh4bEmVR60Zaiya+kpEODBZuaxxlRQBe586ltnItRarL/JQC5Zeh7n3LnQpyKw63q8ZL
QOPEJNOlf/VCkm3Ird+6DI7x/+vQaVtgVvG2w2LN/O6YwXkXtRsO+jSe4DQWPMMumqFVN9YqnepH
kbV8kcNs2CdKc228aycgW/VHCTefuyruGfiL0jrSU6b43TVe+h71eKYGSuSfNtC9/v8Jx4pkLcHr
UIO1o1stGHKaiFZZtYynXER2NkY/th5hgWGX5d1DPSTHT1rBer8LFSHPeDceLvTfJ0u/Be5WwGR9
TCPeEHpUhhWf0T/a9QVzcF02MH91OjFa0zfmkm3NCN7Qp8xdL3G1g4nLci6zbaovN9zyxBX4vWbN
NADX981BrwtIEWj1/vNfnHL6pLq/jmciyqJaY/HNYBEB/KcsBA3bEVhMxnNcydIjxtDdWl936l/5
cy/Krupg6+ThPbNkMo2NKjA3K8Fk9CMRahX0FCmxmVejrGnkouuYn8bpQmUgqcApb5G360DnQT90
9GciyZZs/QYzZjlEfVsfQegbrfPz8cSnJD17/Odm6yvYgiNIN0n82l35gM+d5GWCO5BumztGIUBr
H2siCzmAnNfWV+y1RAnMquLGtb9UgC3NVxZCmEJm/UTGYYbqquxGpCG3SXQ5n+LUP6KwLW+xBUbg
sl29GhKHqylxOqpKgbnkjv9gj+Vz50kbi/kbWKGTMpzMIeoMfLfp00Lckk5qoCNI9tbwDtNTXTm6
n3e4grtknIlekdieRTvsDz5zAQscj0ThHyPPZc9LKBwS0h7O9CB5Ebylzmhsmxi0z3TYs2vwFnCE
gj7fUYpGVTebZOiPmHE2JqUlfqCDt4PZfedegOq9Jk9q5BDx+230zxyMJNVjjA5ejUO9a38MIa/v
mqguqekoJyCvJC/IiPHYJn1LhWR+X7dZLT0JgpFhYdjxP1xGQpMUHOBbtev5ZtX6RpA9Ta3hDFQa
fJY2X5Xz8TM24kB5tE1XQoSRgNYSbOAOgGaQY0lTEb5llWmVsBR2w3IR/imVqW33IIor7PfZrTWU
m8SwAZVyUMRYB1s9MGDoP8efE7xGre+hQCu5xfY5Gws92WUUWsWlS+brjr/NOgPGu2N8xNgP5CvT
O1wAgwaqMqBeWvcXdZgCwFFcP5S6VllhQ6QkTxLxtnXcml5Veh7eGvc4VG+SAFOFzubXxqnTDctL
BCOffmJ2LrG2wpHMQLVpY7TJwnWJ+HcdFOepHjscDkjRvd8PwGF0IyH3rBJO6DAOnuLoCZXBf6Rf
KecixoKlm2xN71LDQqS5ucsH5VhxK3Sikm5yr2W6eu1grNItjxpI5sE79sJIAxh/gDeTWP3GpfXS
YzrwFrc/otUqaHuxSkS/DV4ZeEVTsCanLVSLB9T4rVm1psUWzHy1f4N/jzLaqc06PT21amHxeVL4
CmI28CR0nyud6aReNGbVQ5s6lXCl3eLtVHOaC7npIxj0HgAcgn8ZWwPmYQOZQZy/P7DCoBQmBoaI
/sfVGNxAhNoG06EJiqhA0A6QxEUxuCIlhvAUetH4vOLNQjHMSK6MwUXzBPPM7qkqqYMicEMnN5JY
JlFf67ZF4TZTz9Q8VVzxBhmoCyx07t5dUkh6PYSlQ8fB8eecD6QrPUpSlqFsf5UExl/PHfBeDDZP
J1bT1XxELvqTwuOCApvchAF1zSVbti7puFI2M8ch6K3oOUQWdwAUBJ0Eip1NgNRjlU5+rJLdOUU7
Exv8IhkF925QEdcysrhppxpxIILbm2s5u8bgTT/sxDUDt6yTa/vvxdWovbFB+AWInucybBUTzz8D
knghTDud4kGZu3ql2CEyxKIwpsrVjXlvTmmDMBi5YFA9+cR3kVGxeLuQ1TuzIf6lNkLrovXei4iM
J8gvBnstHLENoQuyCkfQmzS6VAcU+C0Rf4N3KSQU8ece7Qxeef1TGymylUQK3LpGGwHupl+X24WG
W0HmEqGgxFJNVQk/vnvglNmHV8lg/ZpS1xcAPppfs3b5Xi9KCD1C+NT+oDJI3zOwTKVCerl/0t1d
5YmF1GcuPD12Zh1tQ43X7zDNrfX6wNr1QB/tLmj+JWEBqgzQmFOEPvyRQBHlVrU4swXPe3r28Lsy
MGdg1dKDhBGXGpcrkOwZsJf5tImvN9A0LQZENzJeFjOIhH0OOeAWsXZoeTk4i4yR3p1Ssdw//X23
7C/yWX1qqQy+3zEIdsABRB9cZ5wy0GxIXvrjlbgnqFXbV8JsZSqVqE9XhP2kiXPlC/MlJFMA+ZFd
tuYsB/UrofOjsGhYk9R1kNo4wCJoCCXIBbKorTVuZ59sIyb+JQgVwvgAKm31WlUQhuFaB6/GZK7R
YOoltdLTEs2W+CNCcd3+XyaKcGI1FuHmi+6g6QzSBOjvZtb/H6wVqm03Z9I/oxEeDZOBkJjx1yRF
q7NHCiieQ++Q6608cCbUGtOeHE22PfFgZ0Dtdnb3yXYR1CxLdEpAk0XNVQSgbpIEhnq6FuwdBroz
LnZbd8AlSjN7cJ9sEUtMxmIQ6plGpA/2Tx8lMeoMpAmRkgeZg+5PzTsXt3dHK5xS8SWvIyRe+h6r
3zWl9Zt4NuPAFtdr73MieDba4cke1Dbkw1TSTDtAKe8liSqfxxOyvDdVfTEYsqNZ3Bm+PEzg9B6g
j+wcTJHkvg5ruGOnp3vdtDgp1l2ruGQ7OPRHgftuAhYJhgWv0SLXzUjbSyyH6VCCXCqLP1c1oJ7S
NCmFuIBuVBMSfFISmNhSU/oKrLVh3+tsyiTUG0uinWqoJOdz1Q5cVUwV/PG6XlWLEF6ivjLnxoLY
gRrmyz5fc9k4hJuA89voMjMhgD+inSZ8qujosJgLEb26GucqEC54baBGXNL+0Ng25XnknLLL1Uqd
znt/PzPBuefxCAh/SPEGOxP/Rw/x42yAC9KBPD/DqtaqkmXWsJPRuRlBaNmfmnHJmA4WCbLnZY7M
9MOI4LQFqsM8tRLe9/GwNHwqhjpGyjZ2bUCCc1sNRgKW+gNUbmiLb6m4H4fvdhoj6yBxzHk4fRPW
9C6pGxkTljAcp4iH1RROiBe6FQyFAQ2RMngUGTH72J/jenMZlFI2qT3wXPn10iz0vwBIZNMbDa15
I/PrrL5j/gVZZHmN6Ji0G/dT0PXAKiFxDtOUnvGKF9drnSyvXlAavHd4VTCkZ+IsODwr+6wuK/kQ
e8rHJIkwbAx5lF8eMyoo2LHECE9xQFsVQMsUBMKtn7Fax9jyCaVK5AdrIMrXc/hS2mr5jLqfQXPE
9uXu2LCvRkWE21DUoleoK7yl9RLSMWNnRl3pNSwg2YCVZ7Y+A647TQf2u0XjVp0s4+HzFukveXRF
3O6lAzVhY70dYNrRQLtsBQRiYziVM5/o6v7rShR1THefOc5AC/W8DLXChQIXO99sTbIP6KU9/RFq
0FEgxTIJqOsSXZF16aQ4y+FNmHZaeDigGiECkNovNV6at4zUqXSXO48L6N8CxNXDNHfL1kFZQJwl
Vb0Dp2we9a095BlxoM+yA4ucAbb5czD4tqofjWiX0TwyvUBHEkdGfdr7ZJu4oIJTPEYygcILFL5S
pQ0MH4jYlsSskTC/LTwAt0lkGnSg83Bn0RxFhR8Y6Ffdgy78Xi4ZZcbqUx2VGm24wpR5cL2RMo7f
/xWmBRgEKC8/yRzpipqT2ZhiSMdQ0EySqyIslfrNDu7J6pQl+Eyru3iIDD7ppmD4uJi5Vsq8u6T0
11fv3s96LELYxp2QYFG8NB7WMGxkew+OV6UG6lOfiuc3lK3vChVW4YEp14O9bhU+WgTQ24ZAcjl8
YcOQBVCURirnRp3KoA2Z5J+dNlP+OIkeN5q/+ERHFk8Th1yADEwqsGh9g5kvCGMxWdByB2apoBAE
HWaeeFuFjTB7XMu/0rELLlAjTEte7M5u75mga5z11YNYVM+Rd5I0TvykrlXlehXVXAwMV4VWPhNi
IieQ2tYjrADJ6Zf4D2SyPRNjIBH7ImY4DlWm4IQo+HrMisYJ+ZWZ7XkbtTtY53dNzJgD5uU7LuIz
2t5rkptHOdvePNt7ohpDVjHu6oGLfKLEH7CbJh+ruwWSwv4uFA6SXMdImG8Iu9vN1HWsoNdkoYhJ
7WJLz8EYvg0w1qf9pw7pZ+pefXAO1FYmtP5mD1oO50KS/z3qWHEAW32z+QuGA0pgSHCyapai4C7B
igtVTyxLJ9rrDE11RlGX/ol7Q7kooJDSWsj9FwKOSpBRbNvVnvKXDC3hTr4v2sLCTt76XKsD0IDC
IwrtZapdBBPHh4UPrGF4Vk8o3Jh++NOs0MLIWgPk2RMTwV9Eo51XXTbUT/4/okQWh93mvCx2AR+4
UIOe+xQJHyALa76ibV8FNTew8RsybLwTp290r57VALKffc/A3kKzHLs4ybRIVv51nXNwU1g7AMD2
RfpuzDgU9iMCq6j8WLt5kYi7JJDgAgN0nxrmmwt5RvPNaslA5c2JHA9yIQDSU2eFZs3fnGNRvig5
blQu3ujOTdrDR0T7nB+q28A72l4mq4gnL9nRz002uFQ4sa9lBPHw9WL1J9VzhqfJQVUQKI9ZitKO
puqfVOL5lpRz+zAhWRPcft14H48ZM//h9+YRRxcsYMGm7xVXa8cb4WgyVSBgmgDH3DeBOVjPfvMp
qrWtVoFpPB/tkBRUr4WFY8upnl/+mLhbYhn8/s4q/TC3FzbNu++PDL3AXfkDarStXc6uPDc1vh8I
mPGY82G8f6NCHj6iWBREYdU6l6F7acT/ROYM60Q7ryej228r43QsZnP9IZ24UwU9uk9M+e137/TK
RJzkMiOlDVZ3CWhzrG6O6BiTqZASQazrLhzuyI8JXjn9QeosWw2axrOboZzcF2AewDjyCUuM8xS7
W7m/tSEQ9r2TI/x8ywj3ImIce5eNDPfioWV48NMBRrH7tKUyFeuq8+9X4G3QtCHR6cKkNx+YI6mG
KIq+s92LvP4V9uNX5FxWc2tUH6o4GiIIqHCf7vGomc9jWNj013OrZR6uEJvI1FC7w/1JBhKviine
iC1u7kuNIatT9s88Qf8s9sRYljprkYhD9094XFawecRk9O9H9YPivn/6nvzT3usfLI0880TM9uFb
xRIceHDcASdStKNJMS/MKxW4UGi6+fw24Idx8aHKFohuUnlu9Wy8fmkk/RcjsqlKamGXiK5jWJPL
mcqU72v+DANp49z522RdW/N2pLfd9O9vT/XpRNiWBXMr6HUwgpcra3QFNLKfTQ0umrtdXDmHMyB+
gimf4oIy/KICVdI5xyBrugBPBmdusx1v+6QzPexmFpzjW9oqeqGq6mm9+OspD4KOvi9RBySum+nV
Ik9eGxQYJaO9APdSkgV8aurhPUicl2Au33sqOJX3RGaC+Z5jEgfs1WJgzn1e2SR5X5vg4Cu8rZWG
tFtN2/0Dtz7ZpYv0E3mKQq2CYkvvzQCxqapuvSSdf/5IvoH3ckzlQp4iaLtdQJdclQACTIsW9IZT
e70GCqItrv7wJnLZ966H6YDvS+1SvhrTDd+AK4LJn+/UjasQssPT+7ws5uYS7eqcizqHGTuGMSNp
EdPlNBr0Zl6tO3EKKN4O7KPsOD/5aaQ/Wf73zfD3a5B2xHpVxxVRqb2d4pYwIDxxmy5YEFOehaHX
Vpyph7wW8YCuNxgE1sbUiXts4CrtmJP12z3Qf2WCPevrbNWEdLppux7YVgf01ZT1NONYGNiLzpFQ
ZVkew8ef1DfR2JT3pOAv4BhtYngt459MXXp3oDLtLjbp9X7t+6DT3/SUZBrAFe9EqAU32afn8uoI
kbXw8X8UEENeAaxAEbPEd0WFkevDVlH89Luc7Ox9azqHvS6Qb36p+9UhNsYezw65E9uctAkgwMAB
N0JS66LbkBXLeS6gagjP6eUvdbbmY+Ue6iXFjV3sfyBbLQDa7NZB5YPVrkrf93eU/k3P5DPvNzZ8
LGPCKfk00ih501gJgUCwa5bUQdxqbo4wN4wfF4qc6rEPQdo61659mib1ykKJoETIequsbFflr/+t
7xn5F6GS6xvcmkQgbTPXL1Z+N0rDRWUOAlaN17AihlsKlhhHwdtQBTmEw5rQ3vAdVVSqurCpzTfP
ICNG3SJsQscZjVYxZx+Zpgq2wDC188ulrA3JCTGxZCv3kf8Hg+8esyGbejWEO3+YgakzwHK8/Qdr
shWWtHP8bGVSA70JRda5FKztjaZjmOU5+AoBZ+IDnMbgV6EcfZNU5F0yXEf0pkKcSu0XK5pc8leT
VHJ4U92FaOk5NK1M29ecfEgQrJmHJeGNmkqyv8yjI5l0tM1HY7I5SPUZe76iaFtzNE7C+5AKnyH0
Gys7pAQ8JaTaZGzMBc9GFnfHiAGIoaB+Gvry6Ws+QvilE0LfMnJ8CQUzGpcYXM6QLHsxGjqmkRvi
25Jz86NDARocvSHNv+jcb4plyuOXQdw1CpCaab9oSqKKTNg4uS61NJo9IdJGJ5VEnsuwrC7ojcDP
MivqHtVmErOtpTSU+RBMsv5OD/Td2yNXBlBq9NkRxPDb/oeFY4OOJpv/0Jr9Jj/ARBYxaj/Hd+PW
7JJS3C6qGV3awjzJmRN48ao4+alMWY5e33RcmkasYipvTxAjYhQ04OtL1axlL3XKdAjgCaGSbZrB
9NlizCRAr4MZicy2GgwK4vccvZRCbk9N0WWmlhBgX6j69yQbRzLQsSSPfxWLjWLDv9t7uWppcCLp
mrdvFPSeTuMrIjy4p04k3DvoSCGuzgrF6OykMOazI6N8mksA9xy3LCqoRpuc+nZ9M0enSXbyeBwR
xG5d+pgIXecu2tW/boIe1fQ3INwOhXTEeXaFBGuGIhCuiEnn+zxXCO9dHO9tj5/qPGWJQkoeag90
/kj/LymiUZ2Apiyssn15k/hdPZ4xr2ueHVzFCmKQIqAHX9jm44ZPeVG3OHyq38ae7tyfVueGpikm
BMaxMUhTDJjsJUKcbep4bCKdChLGjZ1VTtDeEt5qGasWBVaVjFJe35J0Fp6+10NVXQg1OETiZNwN
c65EeAkdFJpT9s8JOyo96p+/yFw9d8Gy3/IQidmX6V6aWpH1IGQzNHBZdSdloht/Q7SsJSnL5UmJ
UFcV2e+cXbg9mrgnyiWtkL1VS41PSMyXSAwFpny2z0cu9456hKPZnpLzgS0A9zvk0YGOhcZFMRG2
+w69shbOt1E0bVHWcIuobOFvgDq7aGHj5XQpqpRuIE/aZUG+QT+5tyzgesmLsTfdvO0ArspUoYPJ
z+7viOfPjsxzpthJ/P69En7c9c4Z2+f/YpSsCH+4AQxVl+ms6IwtmS0PvV1OoiWCe/x52dPnlhIG
HDs2qR0F/cjm6PN9DrE605Jr6p9LGZsC3jQXbb2yidIHjFQyMPxxEUpAYujxy65SDhix9dJo6YI+
QZxkBV9UQRZW3UOgWm6WBqF+Zwl/b8Kr6GIWK5P4lWg9X/m6P/n1Gh1Qwb/ogoHmNopIILREolBC
DCFb8HW6pDFyZ1Bxi63aEf60mVv1+lNVA1RCB7VlGQCyaIuWu09R7vOo33MC8oBA28cw2SDD32nf
4Y9vyIdSlAgh+LsYel0/5GUAQc1CWOPTzAYcAQ6rammPqbkUylUdMLnhiGmAnNSrEpXB6oJ54tSj
hwZoNYKDm93GHxmGfdIh8CfhSFWYBTxvxxlWqbvHoG3tm9EjzB9v7/L4IkD2w48xP1ZFkXgutL7W
lkn9Gt4CQ2iKxMuklOkDUOAVlmN9TkdnZ8FqvcUKjZTe/X59qjelSg3YB+3IQFiYqtieVS2OFAJg
5a0sd9adrNYIvAzPE2FU8seM8K5t4oYVfO2PjxDvseu9lsAK9eiI4lJVKmbYUXE7lZsIwfzPofZ3
Qz/8NETfNThW44dqa647mjcaCpsPFHlXDuYbOWPTAqU/3R5pvxv3PD67Z2TlNGR38kJEGJYg9ngg
04rtlSEOVdx7tuZZqKK0LN51gqCgm5XLV+1+nYDOTuQeg2j0aUE0fcgyGe2zIod48WzZqeGWIqVl
PT4AlcgZHzupHESo/ABkQ/MbjGtHjp489jH4D4bbbP+1L0e73+ARdOe//7b1lR5w2T+uIHpYYVxH
EA+Qx14S5w9cMnOGJm2pf5J+CqpziYFfU/CiiXcdX3RXAZZylmh9h50iV8EH4p595khpEkFIvVWq
++5BbUZSVjLxoy6jfaJ1aiBf/rGD+RJUN9OsAul2xBLL8wALP1VNrKC3udmQ6rNRrNEPtSRiHJAc
Ao6W0VTRx2i4TYbYWVTWOFBKrT4Wr5XNgTkKqKPemECUk3rHDmCA+nRpsRVfvEwzq5M2l8UpwmA9
pw3pskLCvq1IqNANpXSdmV40XECJ4EZceyora2KHvx9SBNLLlsan/b8I2T+MdqzuiGBoqtRltoRY
xaE53aiyS+7GAJGG6JYdo19YBZ5Rh+NNQTkhDKkKQlgT13ZMdm1dS1gQiQewZqBIykvT/eOFpU93
vdfXQOpKyxF+COAQ9lh9QtorgN1AF2VaFI25aAZ70kXroWNqNaFXy6rlZRKbBwaoIQIojI0yj9mV
czcp/P8QNu615kvFmfbdElLlaSCpM0ycuCu6TtCD+BSbmPxgzjMePLAMhhwQ0E3fgtvUGiGhxNYA
tPB0phg+nSHuROhu0mPhJnobrMEemqwGq/p4VWV+out5ozQGeR1EtxStgvDr4WPGpSct2GKJFDh6
S155ncSl6O4ROWzbzJqgfYNcF5K+p+1cdV/dpgOX1hAh3mRpNQ1ChgnvzoFdkZBHgVNhdDTimSPS
10p53qWuYV4Ax4+cdfwzndG+Vinlqq30VHVDr5nIF4883/mwqrtzV0yL2kyQ6OquLLjnrxn2hBHZ
DlraygwENnog3Qg2c9grTpDkb0qvHsYJHidBpgOsEjO6+j0yiXuMgd7IIXd85X0+DmriqirMuUhN
+cSg0njCkDtVT5gy2dpgncAnt1cSYwQwoyiqP44C3hSrHmO408sv170lKyqTSQxEp6CEy36heaXE
6KOAAkUkQSABvyJVu2L/SX3M5e9D/lHP8f6VMC6wMfVGie9NPBNmhwJ7rVAJ767slSZZ0aCzAhgT
G8pqccwMoszRNqzu34GL1Q8oIWq345Y0PiaNmRPkOTtrfcCzpw5RmNkv3ppRddlG0dOGJeY+NnrW
lOt3acgwualyS5U4Uwzl+qEff/nUH90knkcMacss9bGgmo3rG2hpGZzzqD7BDdelUdbFpfQiQLcS
k0vb0Uwn3BtodapPUVkKMOEk2Us7pHBQ48/eOWJuWtGEdPEKHa+aCedwvIsjUoOrp7gAznX0YObp
Tze4sgzqxm4AX0UgfEOCjEqhsJCfwmpCWlDL/7cN6yISQ9nxQxq7JQiu0ykGRsV2eJwEb58bz+XA
ZmFYRpCD6SH8ds/Z0s2SThEEvsYam+hc+Spnb5vCJ/7pV/0JpzYqfSeBXNqWHVjCB3ph5Oil332C
jbixKYmzRAACzTwhjlv7s/E37uorfz2faapkUkRPWxBsvaPi+vvzFM0uSgtsTHUKQuSHw3zs2Vsw
qxgY2olgUEEwTnxF2gmjpU8ygbGpsvWKZfIa+esSWRwAC4EgczouFBALctM+wWTxMoh+Tn5eZ22b
x6WsQVeXj06M3H3kUgigDfZaP8gLwYbu6a+A/D99e0/eozuMqIgn1w7iPdJoNZNSwbugsaZv8IFE
Iz/46SdPh/3MQmoMf8gJXeLKnRhFvDc0VWCB85CcRbAK8lU9tfP6wZgMog0t1C2Q8KDNrjm4XDHI
Ea+mfnI2KJul8mTTbj/fPsne7wwULGk8fQl7B93bZBxzjUkar1Qh9mkjE+HivKd9KxOeDCJr5qqJ
QHEQsE5ndJXPPY7F+Eha31BKnJW2ia7r+NRuYJAa0FFckmTTqB5Od0oqMKYQneOWQgdeSmA3OTJq
gWCglFwd6dA0s5GT9e4WV/kfZP271IGxbGY0JcipDPLKYP/+tCRLXFJxoxBDMvsYeFwHs0bgsl8Z
mSK22z6Y0hC7Jdvat0iotXs8+N8uy5mmqfPokNHdp55o875d85g6OukAs+pPwozuAAKaSReaTK4V
7QipLqa8jaoubHtiVtRt9+VMmS0JRL6l3MBF3/evOMG8voEjaifJSxfdIzY/wNmrjXv9fmPrPREr
sf8jXlhaBDhPdDAkxe4I4MJgSh9fxkaXTueJpO0yTzyiTfrBbJhB5pS7v4UvuqXXp8qf0fxPiv4L
Q55wRBlTexfgf7Yg/gNil3yn8cDBeHaEIw3VxiIgawr+9HafHiY3mk41QOyK7HgVrwQmgI31IT+O
jsyAWAJnh+YB7Txi3ZRJGZ9ubm2n8P1bZbM18gxzgyQgouexHIrWt/DX1NZVEtGio6ya5YmfTL7n
Zx9YPuAZn+txG5vAgysb8uIUnW9p1vEQm0b5+1S7pF7XGHxYfGzhHhf686dF8RdMxNdjPi425fFW
dMJkYjpKatCqZCGBu5ECV89h4bRWDTdYVI7jlxmUY3KMSx5rzrxH189wT+FKI1bIgyNfYKiVlgCw
yBmRMZu7/sJFUgplYIvHrD+H1G40n0FTOow+riTFQhrSS5hsw9w5HCc2khsBidLxiNAhOFR5PJSu
GaAmYC+633g6DZ1rAE2OgQoJs1B+Q5IOJ4Im2fi6GO4bXOJqz+ng1Wtieoj4kgRaW+14tZhagN/X
xjg+540/8WipD34stF+VpwxT5UVWvImfG0vOIvlNLW9j2WTT22jm6NpKGAF2vhKd6AJiT0wBQzAQ
0kWPUvuP0i9vbLmzPXeUZFDGUEW21s7O77vwVh3FCBJU+44GFboiN9qu2rKHJd+xYOGAPpPID8Sg
5v9QFucAPh2SgxgGYwR+LNrKFVYB+k8UvDpYQGD3h0SnC+53PalQhchKaluAUX+lQ6CJyNFhAV2K
4mXRdc/c3QdLImPqIc8PiTSi0v9p63DnxP5+Pwn+Nx2p38UBKysMnb0b0M6iL8xD/HiJrO+8gtd5
CLYPtpzidELsy1CYGcN1t5Mhr5qm9keLIeegGuzyr2d7juKyaPojrsI4pEGa3gevURi9k46cjj0a
LOVswtKq6CNVxDBbNav/DYD/bxd9JC41gct4lZUfzvQOTvy6LIJt7wZMWOJu0XoPXp6GBrAuPZfN
nJU9MaqSE5H/oRyxO/OjJ7zIcPLKORVp9zbFMcvR79DoirTBoIJD8zsknqBb8ZtybBO9302s3TGR
GxNca0ARnvRd7ZBh2ilctEodvi5toVHLM7r1Q/b4RyjSnw+uGvLb9lksRxDmoit5kE73ZNLXrPAJ
QcCEM9OSuTkS0QLvhENxzHD+TbHNuTHdK8dai1FR7bhW53m1w2RcamqY1vgMu6G5h7e4WSjulNrq
7bPHIyPLyfeFex1iDmuMxwLek+qjhMtfRa9nuTOK921J+gkEsz+T2N8l5mE9qtZcLWZoP3Lq2kAw
7wgt6v4ez/iobD9T5ODxP2ZSOa5I0o8fs/FpvVz3RrmP0E1k3zA2a06gjcWh1UDPOub1tw7ZFzZx
B9h9N5AyQ+j72LuffOqeQqyt69LT9iknlUd9Q3yCcYKv5wc2BWe1tQ2n0fTfvImChop/UTHHh76C
IIsmoUqBdieYSPOg9/BZOziiC3SCJ2EIF/MBUlBwEaEdxDP8WZJ2zUsqs9/NhcwW/lVRfET/qSeH
prRbP4KYCEsBsaCHcVSKj7vAVJ7v3WWvlj8WHkKFiYXaPoZzkmBzyYUlvQ1eLlRqeGy2WkrgR/KD
pl/6Ed/oWVWdRjG+k5YO1vTVxVfQzHEwTz0aO4VCBBYLO81vr+PTPh2K8Lr73koB6I97Dpz7DS5S
IwawtSLe1jMSdsKNCqa4I8lMAClW4WEuBmdUfX1E2ulBIqQekEyqh14NM4t8Um1BcOGb2DmDaPF1
nz8mq4NTe0UfPKMlj/sQYhWdxOuOXbO8cSZ5A8MMVZ5kI+RYTqPskB/8qSI4lMnoB3vHKKMbAl64
CYX5hG2JGHmbTbsbXHjvnLFSqYxJ4kJ+jlZ0+lf+BkJ6hZJYkRyFC6kd/XlqzUpVuWsj+IGd6zXh
i05KFQ7jHac5Te1+aaLhoPpbQngjljiOehjZAVbwK4ByqElNGZVznG687UK3MnI/m1VPrAUY9C7m
+u6IFHbEsjjnbzaXmsRhP+twl8UvNNde/qak0/GlclWzS2uxvrm0WU5xWoNxdgLbWkIKPbSv0nts
tkJRuZ6EzQtYrnh6gELmkLCb/xf4jBkdEoMtnGStua7mjacyeWINy2vuPv8FOKkqgIcJc1/WqOq5
skXKppGETG6eijv2/qSyieUP4DQNzTrJ1528IFjNv7FBBoptreNgQk1zo+8UdCf15fCnPZH00vTG
vv0rmmkQo4vTqx2125nXTNriYwfDjyqhbkA5Vh0YSN1A6yZRK6A8eWluzWo6g6uaxsXWhI8Wmr/p
fivSqpWIDmws6qfx1KWbcaxo5otre50e//t4v02UubYoCTu6qvXzIyBS9LT6qVUxZ/5/+xVwiYMa
aIydOCGe+B5kFKl7PVI2meih3gUNMTOprSSt9liWNUbk3z98Z4UCp9MKXlrs1FL0fEPQ2oMqTHil
+BbSq7TkJxGEd4Cy3x3oQ5G5DJqBKrN33cMljJG9bmlTQkXbUsDy8rtsuWDsHQNbpll4epnJ1/RM
FCQQs6T2sMfe1L5vNatZM2D5TK3AxQaJEtTmn/JTnDLmlPgi8cStNQN5cfFVfpdZtzVQYt61N4Zo
7xsXuDBihewHSfQVC39Udntla74aWcghD6lvliXWoIOdxWvf6rkueWz8EO8XZX6pTE+0Da0IN3va
Garoaq1aB1rA4U+AZIdHaKVT2urKeN/m45TU8VZHFpQFQvrXUtXHekaWNJiLFHj63/CkUF1CJK3W
zX84QVweyvimNUEZ1E8FyODPwuje7KJqvSnRYwY0ptR7cMDy8wcM2hEAP0CMQAYFHHtSORx5Iev1
HdJRp0+zsskGkCmnXJAm3VGvmpH5yxAc8SzHFYB1dD1qH8bFz6wqrg1aumrTstLprr7TtAeMRYU/
oxdZoe9uHoJB9EOZfTcXUP6W4I9rYNRiiBw+nm9UADRRxsoM7SKv8S6prA6GRId1CC3GK09rURxw
9Mp/rLiK9J2tT41FsvHsRAsen221p5OtqQteYLvyu0B10AeP07JQBOKVOigaZxISpGR4Skbcctcz
jpPvvf53oWjctdcUUSRS+mmCsmMXSElW5cl3AfGQMPqPA0PRcnOtEiiAoOFO8dp7hK+vq2r9t+OA
TOow00+AiqHBFs389oV6Pfw6JS38pcv5IohKfZ/RPmiORVuaXQVA4tfmMX7DzSHvD+iFBRHlZXbO
1UTckhlKF89Iofcfp2ldRArmO+5EdR87HP/w2dehj4CqcPSFjI3j91wMXS47GE/bxIQ3UQwA72yu
+4zJHfgpCIypll0wgru6IoigUKZ+m/INA5XiGBc87glYwmbP6Lfw8WdVVmZW0JdbYckXfh03+q9d
3OsFsBDFViC5ZFogxRPZgp9S5qENIlkBEOWadPY0H+uU+IP+hPf/3OHm9PBjJM1QsgwSDrhvjkLQ
q/l34bvEAXQQBngFfVfbDthAMgMDktkStqmPQMLqxOKi+EpTzipRf68iMquOGmas9fruR6Q3QpmQ
FtyN4N43mpr7ZmENcnQgT82HFBSblMOWrH+8VntFCZYYGnySy5/5k3ZVH17LPRFm36Fdm+eaWNCE
Wyae7rTuzSl/iVTba7aea9OCQADe2/4ndeQQFVQGrlGo9+IAkAwQeUhYA//8yBIrLLp1iBhOQiME
Ww/leRkbjJTAxxaW112TzUP1Jg+bunQ14AzOSgihl19WvwKta9e0yTi4VVKQYjNE3RJqxq2ic4s0
xqG6spAV1IBLZcLf8l8+pTWyTi9vHO7wnlMkVO4NbVfye82Wk3zW5m+vIgP9eN31rhTpgYYrL2s6
GjZrLRQqSGi5fKaa64OsaQTuNo+BKtk5dDyVjn6uaYhieivOV0Q03zNsQEFfRbp/Lg77+8AFbKhN
8bUGPwEsBrn6V2LkhRFaHhOJuiq0dgda3mOIxK4IeMlGIUVNffdjTpCPsLj5eHF3KBnP2QgI+VnY
AzlAByAT69NtIlziw77LuyMz4UUTt1TM0LNa4s89jkbaLJcpuS4thrMS/JYBUOITawFIge0z+whx
xCkAWK1GXXGaT/GzAXmzuYCJOqMk8pAS0hc87FxUp69sDxFr4g34qXYGJ2NMPF+QcenOm17rjBNh
JU3lr0K4rAaaRGXyyfuATfTQJ2Kn8y4kiTWiv2Jj3UOM8yAcXUbKPQvSCQZjCPiFQ1qJC6R5OEHt
XlXKGfTeoe6HfPVxsUOZ8nNWifjYSpH2DqD9/E1TVsZeP1EBlx3zfQmEqhp2QkWtu5Vc94tPKTVR
ox9WMmX+Yudg0Hy3FVbiRtBcujIwdQKmHEveLvqJFp2tuqAyho+DeWSsIXPkjj7FKIjwmunFqzfg
R/Nwe5O3J9YAJuwbOVCqh0U4Kw+eh3EKH8QM7DGgaOHPvYMEfrJCeKWtWIliG0Xw+v47UrhcTPj6
2zQEqC/SdcFQrx+PyBDO27omrYM0QsVrVVdSHiZpuM4JTfdRbqGWxi7UcPW6Q0ijC6SrJyPEd7zo
yvdTw0crY7neJS8K4NBTSydAe35cd4518Pdr5atxm6ORBRE+4EGe40XSnmz3SJmW0e6e9bBzobbZ
mJn9Q8dPuo6tVOWoueNitIilxy2MecVtH+mzYn1ribA5YXJyutadrWJYh8L8Ra28HmMV+mZwGsIf
PCleEy9A1iHLPlh0OStmSz0ZRT1DyuY2Wd6O0390ExpdcWRJa6LgH1swcJCeExojm0StR0DjKON6
c0Gt7kiAijE1uP8K1dW/VSGTRJKsA222xVa95vjbV/YJaosE7Hz88PpPylHfWbHbVvPXcBj8TseG
4h0PfKyc4Bw28vWO8jFb69/eh1ZC8pizKiWpmqJzwCxU2bqEtCl5mej80HF6KjLG1is06MKZ9P2x
qZMSNkDBKn7S0xe+ANAUwtLwS3AtFwNraHMl2KYLKMDIwVEQEeY5wnOPzP4noDCcTGf7rPynRQZM
0GKq/1FSCZAFtwuwhT7LXxapvvG0JrKWSQPwsZqVWaAYEiwapE62A+w7LncVe8vnmdWEXqQD4BZy
sUfoJvn+kwxviGa24U7sVqg5RMYWSeImh/OOLxtFC2xpL9q532zX15/eDw5g8yeje3Q74iHtlo4z
KW31ARpgdnvKgIcV+onHRVekpdhQeFmM7JZH+kqa6E5s6VwQJ070Np2xMWokVa08UYVy2bn4Pkmf
4ifUv7JKa/pyUMhaDVlbXyzG1AWVODaVxIWFHni4JRHuo3iVP5fv05W/0jPKMZ9PoHxFoNujWUMB
MTShAoR447STYWILWsb9b8y9l3bi0lzed3J8xRban8i8X9cskLZLVIqtwqSU/6G7HfkRQXDEg2aB
OGO/9uAJ8qKeCPIkUqoANF8DiAPR/PcC5SmDV0yrUSgZGdKILQqZQwoDgWhkjbhpWmbX3cP1u4Ux
Xp8AjqvSUhGCkLP2i/ktcr38wo0TJJQ6ZBRNB7Fg/TTSY2/BMvWjBi+qu5mBmb9OvfjmVZ+DtMhQ
7GJi7eDSLD/RVnlvuGGh9p9skchKH5hqffrXwfLQOmACCQg20dkR25mGvIqabiMgbZ0x1UE68cJe
ueejOTJ+cYoCNJqBHkTLb0i10r6dEErHa2mCJmWcUVJklV9O2JKKDnWFODMnhNQTnIwS6d+FdT4a
vQ+XQe/FdL6zzKTIyLuBoOogpNyMTCHvZ0X+mByLBSco7AG2QlsG3Y20dGl4F48CpALFsB+0P2rt
iGlzN0nPK6ZPXXAI0LAKg8fUnj2VW1RvmmRcOPN+Ym5Gs4zu+aosQ44kxZN3VA9j9LXEneKix288
m5KJghXgxibwQn6S6Pf59X8gaBW8M827aVVIxX8+D1vMFj/5oDRkYaxjKhfLgrUkgeKD8pwvmffe
cPHGfX8nRy+4maRppZCRcujtJfvKvLH4RhiSTrnHhtvbxBTt4C/iXT4YP5DEI4mrzobCGdeUnIrV
0qEBLluH1xh7tNbnLiY6Qkk4AbtgzMlNb8v39LQhEdQgGaTzUUdzQGDynmPM6fVBA18q7orKCW5W
6mVQKgthcAY9KtvDZ2zmggdbD9L5rCJNClzSTY/ZRsrqAb3HDSFmuydHUnbsSzIBnu0AGsbuVGHi
0PtWvrq7NHRWMReojijrglNTdGhft9jF6LN/omuh9ufY7pXZ63sNP5aA1NSPUFTvQG6FP8bL/BF5
13zeJGUQjmGB38mdUHaApElER7BgdDHuNcnj0nF/J7F2nXmjdlWSKaah1zOH5UBEeieq5UQcxe6+
MVGcn1k6RDpVWcM3PV7fQsPRz7Il1YwgA+ZOc9ip9pwAbojBzpnZn86bhdxBIToOuv1EM/fzfatn
jCpDPNh/acggSxZelK+qSwIr4XcZX/zstU1hCbjfqoSNdXUXQY2duOspnTPkFCb49rWY1jy0ocA+
lk9d46eSb8nvb1f/jqbDjcP7/QpucNibvQ3YIPm1NwB6MX3jx9lSUZ9DxsKRsmuOjy5e7qdJh9DB
pRKrjpKRefr7sW6g6qAskcmzumY1hn2+n0JdcC/aN4Xua1ADAIXhazSPBY8LTmfgqll2zmltZszz
SVEf6bTHsoBBj8VzTYGbqVxqTuEQKhtbUxuj70uhY3/0lQPItPwqW6TUvAkPJq7iR10DNac/1ir5
Z/3F5GW9J3SknoUE4hiWZP8hnFebhuz8E+vv4nPgKTgbAPL9WlXI3xGByVJLddZG6qvT9mP2n7IN
ZSOlxYFkHmuXZIC9uMsAeOzTIqi8st/PgqzA4CNZ+FkdBtbiNfgiSAkY3ATuzHzB8BrikPN5HbhH
os8ElLq8vQ07UoZtTVy/OSZYmDMWJiwQ3v1Ju6RZp9jB6weQ6rCPASEUt+dCUUsCTJ4PVpfzKtSh
TEf6CY09O3qgac6HhmY7EGJv+oFV8mDj6fLbK/d0Eutl+3sy27jV3bIkrreT74J2jJ2SNxQ3qFOI
ooYDhz997kC03QNL/05awmQtUGpv+MTuZg52gsDBldRQcBANLsvpoY7k/hwK9IU+n2PZyy/PdGja
PPtVHxZ/U7buryRbiNoRSJdnuM3+icpjKxuqx/LgNx4tGWLezw1y/2lC9R+Q7qxjV6CrlUaArpVR
6knYrYLS+uNvOFsM+XWN5i2mr95gHhKOEOMfiOrVYY+jykbJUH8o3wKzd7Wek5mJDvTAyzAmK7HF
/yG5QYNQVfLJbb/cc5HeLWT3mn+arLhRgV1XxUgIU05wSUMaOlr6yXsXsvi03r5gHhNuxQOgd+d/
sYfxKuyk5b4YjXj6nZqrbqvGDD9LfUR2Ng9PkYvm5O/KNgiyJk/DAIDHLFoBxmBfd9BDSTQYVEiY
X4Zo/XkK204GA9iUrldDiBA2e+HvCbGCGVB9qZeWsUhkXhwQJwh8rR+kOKmlGQ5CMUO1flG9ILYx
Zx8m3vOBQiRfMNyrsdthTQKYTH4EOpjsoELdvCieJz6bgOncKcRuyogkAqvuoxrHZmChVFrzxCxk
mSRNzJaVvu+gxCEcHxP/9nDw8H4fgqwcNPRskAXPjb9hAQVQgJ+JKNPTlNd5FAy4lUYRHRIHbbuV
kpehgCUzzlHs19X7yFFldMEdlQ1QPDS9PyXQhtXo+lE6/vt6DkuMeXF04gglBYlA7VrsMPS95q76
0WYKviAhnxoHWijxc9iVCQVBfPhR41YkY8mwcVOkGZTQVe0hlW1mP0NrILOCphnD7q77OlUKQas1
tY+Ge5BK5cZLRORGvcdgd8W9YDqgmKWtT9Fd7ZamXXhNVerqGdBg9wJb390ZMpo6L2YXZP5qjguL
pE7+Edpmheb3b1IrQR1KXvtQm1CmijfKyJCe/aD6C9KN0mG2v2eDWVQcowsw3cBwhhqIM4K4Up1i
0b2TCt2waXQEgrW8tO4diPyxG4jV6HaJKn9Z28zS7Arqsx5jqtIER6BzpkZ5wRRsSeEQzbWKtTmF
JuIfU5CKd8QdyZ5eV8vxBMxcFrcYhZvynzMcR0dvDss2p7EAHS5PylGVoV4fUgMO9+7GBCf8mB2u
z65QEYf2tEuYEtWaEEewoy49mW3dWaPuVy7Ut043nj4HZvb/eeughAblaqxA4EcU+5bkZFUyobPX
uUw2pIbRlABFrK1yjRWB8PF9Uxqbnge+nJbHInwuKWiHSNvyh/lVTw7JvMHNJrFZ2kRHKquiO+Ax
iTYp1BBPxV+qjT6Dim1kloWovZkxGK7QHv30XZxUglbA4oHniTgA8VeIetq7zx8FdI2gnwK0gajc
3Igjfat7rKLK7Hrlm9tny6GQ634CMW8Gr9XyJ/7NpzoaxEXeNGsDYtxYej0gwtEkseqQQHCeIV4B
p7DdPGK0Q5JsdqxexbPUKJZTDPsBFi/1NLZ9SrajHH3mkUELdXCXAKXXlxOaYAYWea2yHCkkoGKK
TmY9Bf8dz6mF0sw4VQG8nXPVieIAbaN2rg1J0T6efExrM3UMFPL2E4qE9gTwK6Y0Mk2pu93FeUSP
a+p/JKMU3YhsH93f0dvQwZGNZYE9x0VHQIKsl/+elCnY9VKs69vRDPXX0NVwoRTsrwqzmzk35kyx
Bj1A6XYPH1eHUyqPg6aVs4Ws5wjuNJv7LI/4uLSWJOX2xscE8ZPyPURoToD1BQ0X//YCrcsj1WgL
sNRUB1qxJGZrirKb5WPXv3GxzCXkf62tBEEwzsBuijCPx0j4Eni8BK7u5h54X/C2an4WdYQHU1XY
QJLHhPb8tipvzTqmQ5kchtQZAmimZ140Kl7I93KzSKCj9gGqmv78AYaFOF9C8NSrXiBD2hIZNrkQ
1Zc13V/TzPAc9D+eeG/w0xNea2TWJLq8KoppQW37dOz9gOYmtjFyJiA5hLNviaOtOhChffFHXyPe
/6nUm2vCw33NWfikY0noy454ja83NJLcesaNu/z7vtxWdWFIILowpB6W0FB5A01UjhMIQ8nZzEav
/HQ9LoFAyiRZan0WietQbIhFBeoftC26dEc4WlrXuzlvbtQSrmSrOaV9fDYxFocn1rWY5xlMFAXM
eouSVatzsBEIfBWeVpfdFHr4/0Sv3emZ2NcvleAu4+CTJeDJ8M0jTJlijcsDpd1CHZ4rY3lOZLQt
I6C7bygjbKyZv9re0oDg+r9kaN+HUgK+jRMqt0j+guh8LXcOd/46za6FqP84zKE2wymDeq5Uqg4z
dqTBvWWXiPsy0tmICoEFz6EIVGcN0FAFWef5V6fvklreMDA4yyBX8MaweCtHiDX4qTXN7tjcZF+G
A5mvEM5YH2BBq5q2JmfRipje3VFbqTjiSd5G0fb6aMAsf1Koju1Dcp1BOWi4OfkD+IQ8hEaWNkEC
FIJiYR3+tRKAoaUYw59tjq9ZOI0wwvuBLdDmkZKzgnQsAGNCsv1lZcv9LKOOQb+E001/fmSPcSJP
ylfaXNokpysaLssnwY+DS2YUvAzFw+RtoYyHqWxlSS01EBTPzlWrxHvateNxdZXx0+5AkUS6x+Vo
mZY14/gExO4DIwXjJHfvK0emVSCxcPrXbsauLFurICy4tpaCDhBfOa+0ZdVCly0AG7n4co4j1mYl
pOMEV4JQwf/GeOewTjcIOrPcy0j6uDBXp+q3qOxEX3epjtJ+7vAqyxJJQ4ExPcQVxkqGYM95bQUJ
GQv55HLtVVEWNSAzpoRU09i1YWdb9BZ2Ymh2nYmoDcRPo/DUTm5AuAUBgVNZ4OktGt57LJXReQS8
45hbI3Px/pz/LLy5Fi3iHTf3OYz2269otlj4QLeTI/iXBcOycuxsdHQiNQLeNyinTY8Qtoq3SMrA
BFXRnppVlmJ3GVGwS2R5kCrA9xuBOk4MsXaISnHejj+oko/bc93TtnSmWKeHL+rTNR98/gshbNNB
qayZp8UAYkXY3jR+7BRaC3BA7sSlyFzfZAi0/Ww515kqQFNjyG3xFlvpW6RAIdsDGolr1T47fV26
Jh9V9ZOxJyRN+K2JldN6X5+9lWWiP7xXZnJLjq+WgOCedrhasvQk4PaZZKYqibT+vrt/6sod3a50
wJB466RHAMBo34FtVBvztNkU3a0w6lgWluBHRcjQYwkz33t+My+Wm/xctFbEDxWHGgRtW8ey2lZe
HCae8zY0bkVGJPHRu4SeHNdke2sg0iBK+r9v7EQPfupm4KzlLghoQNqYgPi59OBRZGXCURrJ+pbk
UboojybeC/pcrTLPn2zEaCBeqcPF7rjKZS+uNFP1z3czSw+UoQiQ8UWmFKJqedrIRpEnVS0RwbKX
u7g/rK6vXlcWJQ4PHaNvW5yMwRl8aYzAK4oyE1FF/h45Ey+bGoUTYGeJ7YSFccaAPvKpIu+d8o2+
CpRXUvt4gOkcJSkk6zpGeMpmz2PMUTclCYbteWFlHJpKh5Uq9uPfbxidssg+dAeIKb3lL5f53NwP
wg5a9LTWMS22wgC8WdxinaEJespqtWv52uzBUyQJDlb1zbDVDpBEBsINFeD9NcxprHAQW8cxZfQV
qQUkciiGwrMMkfzmJcFhaFU38TVIwuuszDQGL7UyMv37zVlOCBtnMFrgslX6t/AwJ2FJdMwzsg1+
OXaTOavVjsQICTf9+0pwvpzUH0JYXc4DxNDmcZM/s7oiM8BiTJJgjEpcI1IGYwlBxiswQkIbl0Gn
xOJLbTOhkPRS5v2qaWn0LNDle7Ee9CYsVAlYw4qtEQvU3cM2sCesaNPEk6EL4VpnuyOrAn5sZnhc
ytHvS+EsNM0plCHBmiMeEuh3uQifmg9c+raYuI2oL+KBy4sf1cm2X0xx+Whp3UyjogshfIsreDiG
vQ+p7UbFj/2t+b+fQwuV95W3yODKN65JRNUUmBI3KHWD/bT1KeickZDQEQfPCJADZq+J93UqskPB
qYXkvj21uzcGVRPDp5pfwuopKlKu1xd/TCtDGJcqyKOU7UOiRcWIjT7ep5UGc45geqybn2erRB2t
nFJS0EdnyeR9DojypJnICLbAXB2aISS1JCbe9OmyD6CCH4D8l4594Rf5FwBBRI+RLy2uKhDR2p+h
yKcvENoSyWRjlhW13Hv5zkj3VVVxFRMaYvJwDJ+w4nvV/+Hc+k6rGzLc2iBVsCKWXiE4YzjlXZUZ
MqLRa+Dj6FbAXTLbgvHbmAtC06NLlLj3h6PzuaPbkLvBWMBJFwEjslftwgf5ycxIlq61oe9HhJhC
8ZFoGa8MCNmlzCGxkKl+pWxzpjtuBVEXKpe6YXZH1Th8UIhLGkClhkisYauB0YImWfPEqK2rUb2o
oIYklHfcbfAadSg7JUrMtGCNTG4No0sy0YqoxK3bJTSkRL2Zk2d+Ad2lic/LXQCldPPPZa//iYel
FZv6OrtwL36Vgjeaf0T0UovJWtAe6MOavsJpUUOlSyg7HpefUdVsqqrp3NIMvpa9/td5XvJPXlrp
ErYnHAbgxcJriVTbRrnUohom8Lub8a/bhWB1+SMr7dOVsm4x1zfGBYfExiGxFPRpHZ3i06LQLEft
pCQOp/Mmp1HjXMEUkxC8u5HgC1a0ySoEuF75Ls2CGoia+jf2AS80JOv2F1L3+djC8gyRkK2Vi6Eh
m9pO2mbi2fJFCTMl4P8tkYygvShLIozmNZT/Yhjj7/coYf6bMXdBxN/2b6wLpsXqXEzY+W1yTwD0
27ce0hV9kVgkrXXMXQBUB4nhZRvTeVpGbLIzSNnkAM6Z3gTHDBtEO+2QPtgfgL44JgUHEF6hbH6f
V5Qu9/a2mDsTU1RodY4VcWgLBPi/ZnEWRzd6+bVzHWmdo9S0qTm57lkbu6uV043d7I5+oRWBiltU
adCd2Mz8Ecbrr5pTEvWOrvJZD8eHaVWtphLACyEEr3kBqY49TIjOTXSpmCaFWlFmwYXPACVQC95F
G8PJxzOX6sKjZqU4LGKfHtY66b0dNQ3EVlF7R5qyDruxiAwvpZ/79D8u3fxLG82BA+1t2RV20AIj
2c2VSe1cxmE+CEVQp4bdQiuIEByPmkBRwhm+UyMjB8CLE4YMFXDecyGQ6FpRekjMZLFXJDbTtzCN
SXoX61h1KRa9p51phbZlpLmOvRDZ9q1aEpdhuaBJs8stauPNnIMPod0rpz2JH18VK9TZpxZTwEqe
1+5IC4gVADwr8uiAh8/KtwOtMPJ9uzMJ0+RYahdwg6wJ81ykhu0/17Mo3mrnoLC+oRcv8xsPt+L2
PnCpdzYGmlYDPQ05GDuFUuq2ZFTYIrhmfB6Qh4Def7zIqNMisrc1w89sHeAK1oFLVlIi3JmQXysb
v38FYpgJPHr6Clj+2SvFxDsYH+EI+0ehAV/y7A5fwaxURhxCrujtu8MQxSIJou79/+y1DwhpUdrQ
UiiOPjNsepnUah21DGDQAuzh9LQEgNK5KbOxtxsP88OejZQE8E2v2IlQtFS5BIzdYz8ng9Vb1S3C
y6Ub5ky2GTih+aNrFvvQXajs8bbLO65ZLEHmbV97JVp5DQzhFuhXWQsXAYMDC9zn5FTXU9lWd9jk
oFAlsythRAw09hfTIO5ZZKIzla0wz4UkITxTj3odS30neJ+Ly5Cdb5EdNjcsCG5fV2pjnLFGdJaz
dCbUVtcZN3gNNcGd7Emvr0k4XktFuLBFD95ze6UMco6faTB5SF9RHR2IdwSYszDoGh9jMNcEu/Kl
C9sH20Wek/6APxWEul4jgtXg+68rGXVa/dX6YDcCAeRI/eYi3kCw8vzL5oqDREfYhSPPI66Z7zAi
oJeXIW4yEARq4ESvCZYTMP4d6tsdqMVLwBID+H0ZweUtoKdBll8T0mdHeGfuhV5rRg+c7ry8lovm
CmfyOYKn/vNmhAperFcLTacqwkdpxYfPLBolOYL/2h8nJjeaXjMGUvdC2r1iVVN5WH/MokLIAxEH
/KFAfxEQwZrc6+GXS5lSWYoqxTTjUAhl+KtcJ1ASMGGrGr2+OMsjrCSMvj5uAEksUbWKT9/co2IR
6pD/5fQStYZRuAeK/BQ6ZQID9nROi8eC4OjkBid7cQL7qyGIC3WqYNaKQ90qhjRnrWKQGV+s0D+0
6Pna4xtTPmPYKUfBiILbvSdIiip53EjY2vSN3U2v0HQIQ/CdwzIwk0a4HZ97pAUrK2l/nvwdSJMX
XfIEDKXN8uCbvaEbU0zzDDbQAXthJctIiIgu8B9bPjzRqCxlVw2RaDYs8egd/Q+ZD4Mo+okuA5RB
YUZdxnGRq6Eaxo+8dIwntJmmsaeN0uyz6fVyBR7tLLgj/+6xPuHlzIKtifRjMWp8GQxRHl3qkP0P
WeiZjBNzaEwE4Xc/8FjQwLYIi5cKpf7iBFZJ9V7gG0fsicEoNW9kJVGzkdaOEXkCqsNX9Zx1UDVk
EqRt9H+PDVCeO7U7ObmVSKlcGeNbGj63IMSEtXsR99/qtCt6dM+oEW5OmncJa5FRl1T3F96Jjrr5
Z3Sw0vzPpNcIyUBdF7HH8xPxW29V7qBf18CxuvkoCvsq/aYS1KHhp3yo4UJT+5+hrKn+UiogbLjN
vFEugjs+yECaxX9v2uxFWQkGlApJ0Aa5InMQ7bfgd1F+58YnRlNrTwMthAKOxI/lMC1rikrH+vLg
y4nIjLHybHWuEeWwNs06x0h2NU2OBXb8se1wEs8yg9KhsQF8qo7HbsXOE+RDVGjNsZq1MJ4lnsHU
dC8gFIaBFWnULBWitZVmHaxDx7v0/GmKEIs0Jm/kw5QrK+5Jt8UEBR/unL5n2en3zfGK0mBOjVbO
dLa/pAyjtXls9qzfszJAH+xx0pHK+64bEuOCdfcUF61DoCy0s6dMNLsl8u0/u8y1uEeDiF4oXSqE
6tOM2VpmL7PSO4pUcPeAqZHVUk+4qNuiLn8ubqogJebscqO78kv+xWAzxIr5jPpShhZpK9H6Je4C
lwl/aW0Y17l/ElRxGYQwRPi/WJGTPCTwp0L68zWORXoIcd3PsVWZ3/KIOIcZJ2vp82VPMiRoDaR7
/UwR1+Fza+CyNHyAaAAlmL5ClMgdQ+dXQVWpfCieNqyncLia/yq2vxXUIMqL5FyS90Cawkb1Vvr8
Gun340HMjwfF2RoddWrieWKJslHGtQ45EYO6954ChFThDI+FmJatyvwuuCTKgR4FdPtb0mtyreV7
ixfrTad+f57m1qRv+X2Tm0z0Th5KulexL/YVwCsrRbwAPtaJxaamZIbRwqKCXdPq3tEgTpcLFc7r
IyM1RJxL0CG8xNMs15kdJdm8/FrJGRx17W5Al6GhEo6mjVz70DqAdTmg63O5dbjXHZESusxfgsEG
4c3fAF1MLxnf/CMmINFown7X7WfRpiMxa1FHqW7eZqyqtLEdgvMZSimmGNXWgdBYuj9UNfqYKIZv
hgA9YPZnwMiXTWe0RVCADV9sauAbATGEdscMdwejvHMRLgTinwE+KpRc8IdWxjk8swHYQZSsrW99
JiwbG0Zx6Lf7sHIHkNDt7dyMeT7iaaPUdHPlDiifiJho0hrA3uO57+vGamwkKZVWq6FmmL13a6hs
pHiLyawHwUInDK0QOF4b7a0qdQFEtPhKNHLXQTkOITtc87zZd/hITgH2RcQvZfGwrLSBANhZTSi+
PuDox+k7FmS/va/f7R7PSrWaChWFas+Qn2QEtT4Q1R8r2lIYdLVVFE49132d+sturX+BocSgaR0i
Mp1CMFYKo/afdGBRVl992OvMIXbre194PS55ybYyoKVFh+2nnoPQjuaxX+iD4N0SZhYausMAXykx
hyo2O5GCE7Um7G2F0X3nJcloGULIgeGBKOfZUlkY/B12DYHkCD+GbBwhv/pqrSIU0bwTjIEUrgqi
E3NuERSBLDyCIUc83hzt6lTjml4xw5E941nL0tRGTS2vTVZgehO2lk1s6TuW7PzoA+GdHquwFNPd
7RL/STuOzkbhlw/rHnQ0JFMPj9/DQrI51f+LyrIaXZ4M0ZaeG6WAZp+kjBur5ZpRioKSdU5fyJW/
449Zq2G95+k+fOaFidj5qE+XTSxBGVqtOGVZNSLOw19nqfYBXBzAztfYhvBrj4WvJTWw1jW8W+pI
vaHDkMywlAuheRJzrSUmm3lzKA2SqQhbOIS2MGdLsTVdhrH2gSDkR3RN+8ZRYneopYE6tiZq/O2u
7RMvs/FsfzRPRmgTqpQRJkixRORYONmQs/32g2KidS4KPfCU1fDCxAxDqsgFr7J+9Xfw7WCkoszA
+MqavQywmOh2nVyDZTUO74zxGNooA3zBmtkryFMhH68FQM1m3qujVnjXypB45uLcu+BH+z52l3mk
Fz36cRJQ659TQGuIa7VRIeekkWdXFa+n/t5YNeI23w5Pyr7Fj9FH5ddI2xMPtYt60YDt69fBksK6
aozOAy9bwYg+WAT126IyzS5ZVlNuqMoGTrREFHlofGJDaXe3m1Q5i2MWZMSJPOUIQf6aOl4K1S/Z
XClHngTuGJLW2O5SmRD2Mj4LPXNN4GrF0LzGnbOu/onQXk7uWTPWBBSSkgtyxO6etqY1NL76tB6k
dpII0s70GyDC+9fDdgO04bm5CTy1Yw7dAdKoYS7fR2teQUjoOKo6haE5DwboA9Tnxq8/Gh+CMWml
CkgT1iWdbdJYuwjiAdmr6lK24F9tO4m1qQC/8cfNw5SjvIO2SRCfytw3Ek9e1FJxXgs86B/gjiqY
lZa3Ys06898yx6v3bOOszbEm22ySIxa3zkV5gsLI/SYlcOWYry3zgP8rhCikU5GBpsrIS595KJE3
7hlAsYFGJqKff8CxXVZDNIeDmCTnEzQqxwykToc62+XGwMuHO8/CnAdJc95xKX1DFF9+jZQLOkvK
XW27caWFNgkAzWWYbdq3Owh+sYphQ5TAEinJX8UkEZ7SRUBVXh6D4Jnj4DDDdX8wDkfq+VyiV34u
JaDqoGdBUMAvyxYv0SGknm6QTXuYVRZPsPKHLhOk6EVdgzCReVFLcHuXzwEKcmkGBYLa0Gre6v7s
SZoL0K52r/kbWCRJ8wXe9Y7vUWtI0hpVAQsbyhIltxg3BtQn9eOioRQjBNQVgCsd7vzBs25jbjz/
b1upAMrEpANy9S5qPsAmYUtq1Sw2MrS3ox03nQBmxLgCbx3umdLh3Z05P13KbxluFa34+8XJTQvU
63jcgLgSDECTH8DQPUgD7Lx/7r9ishllWlCo/QnAOxyUj6mUslAjnDoAqNlFMox/1bGuIjWugvU5
1DSXHBV/XRFDjqbISEtM/tgzMvHvZ7l2F+Ue75iNlAa+cGRZ7F5lL9+1gzPFSYskH15wgVf8Lnfp
yvHvrW20Oa7r0v9vJKj6EOECK2PdIkpcIBqHJj806rKLeHG5mMd8CEYPtlXZz3i5tUq18ifjTwKg
jDFJGxbU+RuMCpmnuaQPgTKpDRuTJblE0d7twMGjoHg5HDJn7gbuvWywTf+atzhppU2uZlzp2dYd
e2Lr39DN3UpHY6s4gBpFJ0L1Fl7V4zMIus2a7whsWAYsk2fcXOhCTP8EZF0btOQSVWJqGoAq1d49
RTD9+CSimu4R8G4mtPlLeDOqQqtIcTrDMW2aXw9R9stBM63CaqJDzTlalEBRijUSP1irhtwmbAsT
4fd/tC6utK21y28N8ITmu1oN8ULWp54VchucTwZg4yqkx74YQ4e1OAvoz/WsH1WQKkwqnjQqxnfQ
JoHU60hRz4FkJ471cQeCvfBEVMJCBs3cp3syhZbZ28Bp/UB9hiCf/9qd7eYUBrgL9fHPIsy213Hx
TZ/D5SSKmo1kEe44HH5rmtzo143ysk3qoaeTR1g0okZiVo/CFbGiXcTUH2x6pM1QPXi5MgDDVC6A
6Yx3LmyvtNMRd1F2e2/JwFAsV4/dBUv7qKqMluqyZhElEM5UJJtde/3Ujc9RYeOuNyQo1LncLWCk
yNx9ujo2nLr1wG8ysa8Ze+GIbvLtvuiLKadie31p1DuZrZWEy6IK2pW3F1IcQKMkQ7Ui4L8+lBvV
oNe3pUCVOORq+vmhIduQa3DzK64EU57z0rZwzYDq/HC//8GtEMnILoSuppn1BVnT8kabibS/DNPa
5FH4JEB3Oldov8K7vbUHSmdvBrxkD7CSr1EI4tc0MYogUlxmZNkisO/5Xj/gn5PJ4x/o2xun9SIo
OV01mfCha4Mhk6ELcQDp1noxxJQHQkMgo0Fy7dKLX/FvlhifRbc+19s89DyLCC85Zg5eMCl23m6u
3q/Tr9bexDRokXYEpfyOQd3cMDvyOh1kzPbXSyPa/SO/WCTu5eu7A2CH1HNtUbyTaNXvzpbZsoL5
8mpgr5RTDB43Tju+Wt/EA2v9mM05RCdd7RinFI4AcLSmUHVRTpWG+jruXyzKzZDwK8NbBjwBbVjw
RbN1Q1TRwMioamziP1gmz84ir2XkpCTIaLIsBtZQtWirU1k/9Y/Iv0uWRF6yu60siVE6+SJLDoxI
8CZguP+y2nvJqqGPB0XkQWdtv5SDgCwkCxkWFiUdD+z5TFAUjKoXjbTV3zmyXfQ5w/P/3NePSBnr
AsGls2Cn/i6Yl66oBrhRH8WdBNfgIi1/LqFdJMKnGQYYb+n8oWZXRrwPV+FuB97LdHLNgzS0cSlB
bPaQZvgLYpPsiggdObqPCNopzPGUw9mZ58sIcGYcsIq+uIPJRGTvfFh2zr98nhbwkEe8/tmSOx15
UBseJf9nYSX5/9pqLM0O+kOltQQQBBD3n7511sXzIZ9HtTYgE1oPr/Cebu4VRaAJlpm0eCOawTn+
fgVU6z0PvCDPbgy5XINn14MwQl6xNkdaUTUTanW/Ja4t9XozIr1oUag3AaEEw3jTgu+tggRHPj9x
eQPoBWh6hncEbwHxGPut7wHQevP/NjfZBZr+2Vh5TZMGupVM4HZPZExnZvt7gpGhq+SKApnWRdD5
Yl2Hayj4DysKfEBya6GAXBsEmcTnHp4UUcdwv2BC80AIfI7GWRNCbR07dDp10tfoFIot8YTTk2l4
9bogVubW2TN5timbGhAJl8cr+kCzWBZjgByS757v3A2XzhJGwDK6QW/JNkEApfzTP16sVMj94jG3
t5GqrN8Xrxi8bWdqY2XbtoDSSOClpTtZGY2b9no6NQZCA+OhrBVNJ3JXJHvTf0NXudBeoT1I3GAN
GZXS/d99uHWi/JpxL2jXDaHQRVx1AdU1123oRaQgrCPCY54VKBdJpdAi2lg0K5z/60xJ33Pkz3Zn
R4lg5HPfXLxfRVJ4+YX63gYS5azuF5Afw3vGFxE5PTLGSMORiWaNjCE5K8V3n14thBJ7cTjzMeMW
iJmRTh8HkLLKyGF0yz0cgVMYZloVRqBPRYJc+vZUcR2FMvXS3qxZxc064fQ4K2KRfV0WODeJaU7m
XrfPGq2JUD/FVYcWWBIIfPSkf8s3abxnBJLuCFF4307xVcl8+mdvnKorkNrLeBdTUNjGM7MRELL/
iWhQc+ZvJtJpDX9mE8GScBozl2rc1+ytTiWnHppJOP3wGOFY6HHE3hLw3fjmVRgRPcjN08bHZfXZ
CbgW9WUNdkI3JIt+SA/PU3j3Fy0Xcycg5KMFVHME5wCDcpiYnjkgrooxebUW/j5M+W0b88wo7Aw2
JFH+JnJE7vGdbGi5pINqgYpRjr5kZG97vbZdcT9qwP5CuEn9ltrRgGWrgr/E89d1LXLuWIC97jhU
Dh5gwKrf3YiCIOcf7X/r7PUftUlv3027wLiJT1WnQGB691Rkk7OqTil0M78W0cimE2JCZvmkC8o/
vBkr24Fffpt0NZI94D8NEg1OeOgxzump6k5O5a71rOmkzzEV7WfPYXA2uUdK5md8XY0lPwSv9FPE
yKPmRlEYk2pbTZBV1b9eFth3X2Xtk8rBM4zPu3BWHh3IG9JMYB6i/EzVxcLsB/TyTX9zozP+kBcd
uD19ezJy9qczGiK1JzZp/1yauzbRGV/hZAQoKwJMHmhLwje6xcts3sRPiUwdG2E0jZ6+ZrVqejPX
Pm2j31oZFy5gF3e6b6yVp7DKjdZsow5qoEk95urnGiAY6FoA9Y+Uds7+u0edKGbMPpLF748Uotxq
ZpBvvdbWhnjRtIlSO5fw00LRHu8NlXnmL/tf16QQycuCi6qREQTTn3XxGWn4sHRpOKwDcL5USyQV
WjcD0IHszI/hEDrpyF8jKTkejSAO3K6fU1Nd50nkCSxPHe+sPiVECPqrkgJZX6YX6XKIlp64KUTz
AMBJ1azBICRJUe+0jQr9O5us3ONk6eEh2twZEnIeona/AjMCBFx1Z73m+L7ogr6JLwWbMWl9RcTg
AyOiVwUyshuNUGTiZ9BngqdbzlhlQiemrg3uMYwmJXSeOh9tikXDB9vXmUwbRpzwB7EjP33xsoo3
O9bRqYADFtKVbwfbznZ9NAshSYKGy8Ged0dAjHAIuC1eag6sENJXWNnMESS6rVIYIZeupjdUO1UG
s/OJP8TBQUnPLFnWTX4WXxbPIISuXJb4DaDyvNxxYevN4aMcs5n8tPP1emG0OZyMami+vOtqgwUz
WbIYs6LDWGKr4KTFBaTSSGIWAMmRIJBhPe2NPqrjZnIQH3jmgE1UtmH/y/GraaoxD9+aohADpyYn
8oxVKBw0wIOyvT4exu8CcxxIq1WTqdK5TT8cN1Nt4lR1c1SRM4lovKlfgXIbl8baQw/JPg4pxNBJ
RRxwYmN4ZHKyoRH3I8ZuECilqLCcke3CSOhsc9gr9/kcvi83xTP/9fdHteMm9PCvWn/+VRzHLjrd
lqMbvvj5X5E28xMKAGppAvGFOc0QkOqJ6n8Hz95e1DKFsX6CRuKnJITGGpjS9fvhjUHjSyCP781r
Ol/ccADqx+NT+fZpZ+VxRkVwTrvEXMH2HinN7EqmNdGJWY1RyTKlREdVRFQtYz9xBSGkgfW1MGDm
Zq2CixTvx096wER3pU4ga1hELkrMw3IucpkYW3Z8UZbSY64ehdpjH4QZfxrq8KwZ4e+AzC471nri
bjr4fuiNcrc7SmQX6FOON3zGH2Ab6MVCi2XaEbE+nQsLyOJ/Q1Cmcs61gw/2Xa/1N9gCy2pEmiH+
YJEqnugo2e2Ne7CZGUmaOm4DF9If/y5YKrDi92nuPFYHAy8ob4HSHjNyHXfWA+fNVvXOpU2F7oIb
zxJypZjScE5fV127ZnKqlT199J3pHq4Cjlg9zDG8V4BiznrOxs+bT6pzehk7C6sTxNBw86+JAvR2
r/ASijC8/bNE86hMR948G8nG3t2KdKS1Eh9SWw4ozLFRIEce4sdFcHPeBeRfCOS0aiPTMTLOor/k
KwGT/nrwfKQ//YWG7vnQk53FqgoVWlq4xFfQL/ZcaWGdEcIQpenTpimMO42LzQbGumIjvREbwRIM
McsKblKIhGVaR+GQMjXcmMXMCrhumyWHjsWoIervxlFrs5jeS0O+IYX9SbTOdIeNyqSWx9uE0RDo
RP9I2QiI4qtQxjhyoZMhs+Lsk1kBBsznWUqZyC1rgV5yqk/lvYK2OUobSmy9G0EPKcnfGHE3hWy3
Pqku0d6sctDW31tN9aHzH8ka6lUBCP6z8lg4BNaI3RNvaBb4+spZK2wgnpU5xFyT9jS0XTP2gWIw
xjtTG62lWifZlgJjRumctbN/m6OTTRHcShd1yLtSlwgti+Dyg2+QoOOFrcf1c5+psjle0+R7kgTi
yCtMNUY5qW6uqldoZRBWNsDwVMdSo/URmLRi/RZli9CRQ+f9G2vWhXG5WkSqK7UjVJ3UmwkPcoxk
7D1Tay5JS+mpQswivphiCSVHPpy+rPlhJ1iKJ4wBfD+37fn4WrtY+KEVmga2DjtH+xVNqxHeUDdd
8siuwgUMUa9GOgvfszPA6vsl+7kpypIKtOdOw8Bp3mDTPVX9x9AzY6YWLLmQXwDxVT0et/+/GPAy
76dMQmVgFyP4aFAdHjLdhkNMAByB+SAdBHFBsKVBtlm2vy7Gj0XSKtLFGIRz8YhK2TOr8qTXZk+3
gqh/4yZ3hYJ/fOEOL6QKRPk8hsR8sR74N0+txvz7vwc3mBge/Do/0tGlBFvJACnaUlH/foqsLlZ9
AiGcLVsHtzfDs633vrzK+9RSZPg7YkZ7zs9fMaDxVAR5ofqD8aucQYv9IohoJy9A3RuKWW39EATH
n+mUemcGLq+DHUeOptPkoRb08A6K7DYZZ1FydizaK2MzknuSn5ZaCLI6mFvdggbi+3r7LebtAgu0
inC8yqcoMmY7OyV7G13XyaDrE8Ro3YIlqpQ2JPWflvNqRwOXYX8l+iI1ZYRhprLiOkXjNDAZFLuO
m1g/jIIAOSnSa/4svquSRdz4huQ8n9ScAnCbgBbAopKqlpHDdQhYENwrbJARHgebG0FiFbJgk69d
crOAl/26LBEytm3VD1RIzl65J3g33ZvGAkTLGnMZVGBnv182wNdX76TjSSzM/wFMJHKCrEjF0oAX
wiB2sHPMiCOhj29jWOSeXVDwYNWj7y3S51LHnYn5RbuBGhMocwKpDtgQGNs6Atbb2d1e6gRCiPIf
QTwwHDZGe3Imyw2dVVrEb3heeuqVokfE0cCkLYjUUadIBlQYW4ajA+NKP+HLZKlreekSu5+Ut4fJ
kF0ABQTiNnzxIUfu34FiIqyppfLvBFVzmvI873fGGNlpas18jfwQ9GFDkwDovdHmLRSVInP+xwxh
5h2mJoJhqt2qizf7FcuvmrHnJygHjfAUFGX8eDMW6GmRys/FfI1DSOmMkR5Jdaw3d0QbfqJbNXU6
HEeUX0hgcJqqwZJvSShSbFPw+afShTcC1aC2RwIKOyKYJd0bAMVeMdtowGWQw5FOXQc1GuS8Lpu/
bWdJElt/G/BLbtf1W+Tb9qlsUq+XFUvFgsu+uI8jw3Ln69t1rGHEcEi+l2SA1qQFkWz6QmsHc0Bh
00FUnQzGQZlLiB0/AWpnE8BbJvIucEOr/dSMQb0yuQzOUeN7nqSbRCqXwUYpdGJ3bXUt/ve8TnMe
pARLn/A/rN+saPLZpBX0heDPiQqbZRHBS5B+hlur26qI6V1Jx4irUrD1gwFHjHdMhUMecs6REhsv
m+Q9O0Rn5yaVvJ6ovvo4zy8C7+AdKpDLEEPV9D6y7B98+kj+PYhRc7MpXdN0CFQGtpE4RkUPjF4g
KsnGHOIL+p+CkrW3BCKbhUP5xjXWuyd9YsB0VPZ8gYpbZWw6WcsMzPV74uq+LdvxWz60QpUYQAA4
fagoohz0ttTjKTQtL85+BQqpXe5ssbAdN9crYMYKNyRIgD9inJntl9M4fjtz9W0O4pGmWGnPtOqd
0NTYRHjhXeM9jW1k+/AmhfqRfQK0hhdftYSj73nIcCsavvOUzbPGeQBoy0zcRY6IffgAPtWXKEmr
fY88Q9tzXcVI31+eRzK3Y7fDVI26jBlPsHdaNvEvzyMHtTft9aBmjfR23yxbI7VUZqOyxLwLZL6G
A2S6ZTimIM6qya/02NMe7Vk+aSXlcKlQs8/8pUj+yacDpzGjElDhHev45pauAL1A1k6jDKcmeCNd
VKPsFs9PqYWAgqybFLIaLs/T3TDTVbeAibatFoE5ZZvIvy4CwXIRRwdaptgLsAyaR1f5ybaI7DqP
r2dzE8rhCt+Lcc06t2Cy+2nngt/ZWa+JUEdIbUqhyy1RU2uYpsEA2QYXuijVxJaf92F1UBCP0pga
NrKM6sHKSTc+DTAPMujlCnfF5fy8/3jSeXLje5ibTqcWDqj5Q/jmmDD3W3xYKG/IwPkZxMeVS299
McgwNr6yirn9u1nB3E0JCGAE1na9Ci/VSwEXFO5hOcMHbObodkqLG8Qujtc5zWmgSHlcrYcWq81U
KCGRRWMNaCU+d358iWPpqlzA1KkoUiTx5vPzH9tFMLkppem/hVa40f69i8vG/zzwFpPFjZ1BwKxZ
84wtyvo65sz8ldOoNpJfH3IQL23oPkbsF9hbnA7v0z5iUOQL1wOFzMmMlYEndMG6/+7W++H7idSK
s1VCBXs5y0blPy2OaAcK3XROivkbCNSlwUDGsIR4I677BegPHEhJldL6hLwldkRcl57BURB7j20q
Y3j+UHKuMVU3wSx1gNXBSml4cuPP6/GGfOjQrJr7nhcJ9E0YWs3j7FzL6S4fY+2ST4McQqHbxJcC
ThtbmkdlE7CTYMIJB7scQ6qinhLVo4V8SpDxb4+TBLhxmRdcHerxUCQVXBBcAH3yKcMW+Bukbvf3
TbTfH/SOCe9VU/QPRKGVKv5/elrYdoCYHtYSHExvfDkonKdIILyKyeiUGS/Q4iI/NmZ6n3yrBA7J
ppXWbuDVFUkuyOsGFjwKPkfpJcGeUcwgDxQQuQ94uMJp3ch/1a1ExCaSUoBoTU5WnuwCntNm0wtB
z0ZvSvCaqtonkPPcp5D1Mqm9/+LY65/VgSfLcAH1kWngB50qliiU4DlpOAY0XJ9xHKWnFq6Au3pJ
aA+2RtFCYHCxGIf4LbVQ7U/x/yyd6jduWWLsfv59DpdhgJevAcZWvECbkv68Vj2rQB+UQ1qOjLv0
jsNOBxu7ZKkkL/RwFeo/zK6P5Lp6U/3Q1jyiecibB97LEAH4PXtfUDHk7zaAF1ib1uEig4waIFy5
Ap8IH1Z3Opkl95T6b/NQVTQ/ALj3UoDIVdlgJvMSElqBqAfm7Y+vHYwaWme7jEEHymBV29kCgnwj
9H8JqIcRC/77EULKz7c+UXnFD8xpwVLHv1P6C0iOCSwcxlsI2SE1s2Sbum0ChXgwMLz31KISrWq+
dLiv19la3WJ6HwH4WK/y/BTJUo4BA5Vsa33UnDJtd5uj5l5PSwjkZzPmUIIuE8w1gGyIGK7a3Hw/
jcb2USEKe94VrAbxGH5lEzESrtGeys2RoVqprfFY5MheMOOCI9/jSXWLuq6X/tsrjhTS8mz/UQaT
B/D0L32leuQaWmnQY+PelRHJRO97AIqHl4WUzEvi623f1Oa+kYedY7lt58vmLLkn4xx2ylRtBaZp
gIY3qn58rau1HdMIJWBarsxtlNXFjYLC9dtVBe/mGndHzNS/OeYhwRdYj9MrLlhHXM7Y66nhzd+Z
WNSCc84O4J4I6KdVXa9XvyRCV/b739AUCcUmmJNMCfjM2/fDbS3uSEmrK/7fnGmckyW8dZUN2NB9
pOybPr82xAcxeKyeXoBoo4GSYVuMybrlA/NxNySuykNpOO8ZvPFU+wxCnJs2jC1k+XBqgtQopGs2
YvqUpufq+Bl199I9Np2MC4erJZ0Dy0yuoCVl+X5ae2UKtETmiezz5heM0W3GW75ZE99XxNX0KCTD
yt1YUFkTLsP0x6t6xUncdjRg/x10NO8FMtqhkPk3QHXpBmBXmS0gXfvRfCwEAtgrS5F9RFIn2bE8
xxZnkZEh0whD9HosJGujAfLk3mUWu31zu1St+Erj3AjV0Prrvxo+iFNObfYAe77UR6IN45tg9Fg2
wxMWfQX4xSNP6m41k58nCEYm7Y8rgThtpuf0Fr7YbBdL5XxbVwzHMBf7uOsIrfcBSqpfjTqhlbTB
9mqiKvoyB9xgeu7XZ/yR9SZC94KJj7IuILtmJTcyGpZe/v2ShdBWAcmVk4DNTS5+u1U46/lCI9WD
UsH/RD9JQdrWy6u28NpIOZDZCMvRAeCdfak7VhhYbBPkrVpkYZcMYtCxEirB23ne8WWLrP3g3D5B
yO45X68M2IzX0WN7WUe/QlID3FokvdU2HU6OFbtu/WQsfW0UBJ2po9X0hkzsVNZxvCs2d61ktzSL
s4EtdPgCpchSfEmaKJcGVda+MjWLTlQuGNMlO087MMGn6wv0sqfLFyCfS6rNe0qoPp1tR2U5sww4
97LEgyKNuFkVaeiEqYRi5N4kvTCpVDY71KbnpDeHYLgZVXQqs2t79MYf14ShdLa1D33RJq/Ey7BV
y2cM/bOmfIHnX0oufMFMyiNNWHOa1eJKvGs5DCZzAVss8iTpuEl4a0LHHUUARgYCI31SnvDf4AOx
hnGVhh+Cx1tpkAM8U0rY1vVXbLOr1g94msfh6Xge0IPv3fUEV4NCELgI3Ckqtm/KshVAyyGMmsuu
cnnlxyRYSERgviHd5ytENbAIxZ8CGMIZJRHl2g3APhAtFPGDspkTkohA4XS6d63VIdl1feqFskd5
MBQ5LOdQSQBVEBJ7ZJigknqbfhrlj6ehc6iaMBBfJBIJorzBKPbhmJuFERPiN5S4TeSA1xRHKR8k
aM9hlrFeUCcyCV+SSLeSQzSe4mdeXLIbcB8EP+6KG6EuXJ6LxAROJVR0xxwpPBkroOsvYiXNg5V/
dxMei441vOEegTaXRYW6/1k5hmrLfja8Q9aKrnufuw8oGDSJ+lE7MCkumlAyMmiwd37aZco9CZsg
F6nmdtQiWI0K9NwsKbmVjRSnej0kaHDQ+7yRY5PMfZsXJWxuFZ5fqE9d+SYWZjFLYkdKiT4PkFEi
lLkofXhG/rRFO2vAOce/e4vWL1brmMEQFlC1kWyB8K1jHCC1egRk2DH6HORFUIUArhXEKkKhAJo6
a1DY7B7VgxrU0Y/REry0jHLZhLhtgf8C+iN7opDaa+gzeY9zzsMhjkMxZcM/50QsMvTRZywPQ5xu
FynvbLaTwcyD1y9WmXisyY7M70lq2D9S+vTHwW27NDt2tpWDnMb7QMw3ZomWnwN5kf/hHLKC2zcs
TJBPtvhx/hsjmNq6UmOtMuy6o7D7qaxdTsFat04dgE7YSd5Q4gK9zkSRTgGtPwv0q4/zzgejIlqD
s0h7hYA5gqecK6yqYQMbEeKwVYHcyTC0k//XxWo8MlPfg2kClohI33F1XXV8KUCOXYQWCoRE2NK+
2E/yY8WcCxLOOX0+xkhOHPl5o7vXNCFYX4XaqsTBKC+pDxNHnvqMp05I5saz5IZv/VGZwwgJLGyL
GinyZR4YxbVuCyHyXiV4MCbfeSb+Vk6ZtMjfQWhcsaHgct+z9lGEznKL7dL3cpe0/Fp8Eu4ivrbc
3qspxJyC7EhSP3zfgFO1Nkntj/UiFJV2aqAPp7jHKlCfg3YWvAZjbdHW5Pi2YtynRs7yyk+LJhm6
EknXD4wLUWQl7ArLTjmVdFBXXmedYl/8CytvWmsnoAEDTq0gAHGNct5LJPrjJHAiZOb+vkwMLxUn
cE+JMhmSkgrNfEQ1QwCIlSQQQD7bFc77CY+PEuO2JW3BRqC5PQ9kAViFj6k8KcG32U+kXZko/gRf
RXEicgJyJV0RNg3Ki/iKr+1oDn1G6xgkH6vfjG8p3hEevsX5ycpjsXPK2RaU96RVeM+7Jy3esJNy
8R8dpDR46f3EJDcpBMd0ZKbT3m/07aGtQk8v+PtiRT8iQl4rUdsnoyDtRoBcfA430YMtzEUb0XPx
c2JcLEqpuhcniU6hw5fktJjDxH7voL8on4CUjXZ1UCifNv+uaKv4a0m0D6Ln2iRi/h1+3omuLGch
978eShPyyYseeBB5Dn4kxIwnmTNukP/ZS1f9EP/AcRRu11msFG2FA3VHYIysZKurdnyyYCVe6mj6
KahfYpWAHc+MMZP/HXI0zyBHgRig0++bdss4oKIemkn+aJ5BUj72+kfmv+zft2taSlf45+rIQShz
NEYXyzj90t2oz57Eam0sBkbQ9vNzmGFuOcwYVOKhle7XRAR7dzZjHCWCNrYrkqNo1CsXqT32Twa/
QyMkEwmTp8n1xIvgoZaf1s5fNUPwYBa0xBhKBuej2LW5PpLAtZ2cZIOVSR6S8wUC5kBsK4IUou0R
06hcVPdy5KR6HuzWuevJJ2M0mRNKAvNVgED7e4uMnGw8938wlBeZqpgmQjEFFQGV96kdSjUaS6KT
MOVagH/dSPw2SiSdGA6PypQL8R3cDebiWVTJqZFtavd4PZ6sJr7sdT58VcCjjW/yxLu9EcUWa8wr
nshaeYnYU6eEu843Khy9vKin2to8Fa5Ar78wql0amDsvO40Y1EJ0omBhadZyNLHKRhRgJK62ivmv
sITdcGo7ZDUIRl0YkTYr9YwiDbDkfy6LSFTLgjQ46esDVk8CliNZ5Mjvo+xkZlOlLR31xqdJopKB
WYTS97jecXp+mVeZtBR5dKJIAKokip0lW+utbNtwfP4py8eJFvxJIbiF3WHFMjCdiGwgP4e8rAO3
oJcafCu3V8MIG1CmXN44RsCc40Bwxmn2Dec4vxjEkmymIa1ZN1A2SJhHUzgyURp6anZZM7FuGviN
T/is2ql7VS+cQaokCj1xSfiuZ80ZnnGnLGZlh67tyWy+fNfIe9xPg205ZaJ4tFQsRR3ch5D5f5Yf
XxlbC7qskQr9/is4JPWj9oe3NNOMCODXyZ9ZEu+CVlrC7qIfuB1yayiR8uq3PyzBl5EbqcztLmOE
8Plcf+oCy6kr77FlcHKSB0AWGk/5sFmY+3qptr6mM7kka1sj6W7qlIAvyn+Nv0xHcosr/1+Yv+2U
i1MV/OLeKESLLqzrJqfjWiThUk7/dKTYqsatIvm2wPxVs1ISveBu6+7lqEpHyffF06DPnlEq5tGU
1FJP84GQTKhFTkQMZ7w43pe0uvQhTcNzbp1wjuJv6hdxkaj7nML7N2Ye+3XMQVr58oy4Fi/f/Duj
/gbEBhooYKvhvR+DNIP48WkzEMwu9qscFpoTQVyYw35FPmnG0v/zHtZUCzsMJRJAIgOR6wEIF0Zw
j1kMS393XNCbTt/iQJHS5T0T80fzunXNlKylCNF0fktsYKcypz4AIhAhC1fJjFWzj7QYSzorqu2g
nxCImveHMpFBW0fdNKR6jluM6/DSe9lt8I+QLQijtJ7ryo2hhUJLRCW+VpqoLZ55b6B0EZKvZV43
Dc8UxplSspAigbO236ZMD/r6YIEcrQMXBxk461dwJrbU36SjoR0pj/HkmrysNhqBdbQ8O7CPDnT3
2oSmeuSP2TuCNWi8IQakVGyQFMjGHfzQaQcJkrmwtL7UBoqAayMi8se4C10t4rDZCeXFQykMPHg+
kMdNyykRLgS7LSKCexZ7S8IWSZ5WfAfZfIhlJogyJA4I6RwtttBkq/lGjztuQdeFUPfBkLfkskqy
H0sFR6QNrH0ZPt68qDtI2rfASA69xEx0X7tROrn3tN7HhO6ZLbvTgrSnDpkTRRs6afSe3lTp0xzN
Uqi6D8Whgly9RMajZMhH9IUPuo1N+atgtINZRCIzuO7/Ja1lTCc6oJsPfI7LD4EnGMz+GE+C3LX8
FQv6pGbD9F9zNvHOw2YokssguvNAj8mpSFUYYRkGxoWOUtI/rOSLYD+nTI0gWItprwbozY0AXTvP
Yye5adyHBRDrWDrzmXDs1Ig48iLuW+KedE8KJhyXax+Cjrq+Z6ye0BfIsGkm0vQP+xW5B7uzwax0
1U2a9sOsStnBWJaBGaAOMNaVSspfr+/ch5uSxlJ43juBNi2sskpk40KKpDCY6peobwnRAAoGoNUd
1Goy4OH4kCOgbbFrWs9fV+jTDA79j5y5/fvo6RareplEGENxmT9Vzy1kJhO+ghg2oo6W1aL6hv7H
oZUQ9O/Au0iFq3wLEgkmkEBxv9g+OJW85ekqgkzPu7oxpiKTd+vrCKV7DpCVhlG2lq3iPY4n47h4
6sYHjtSpqx75aWvcWWUExeIX6i47GSxWhXVcLdF22WoiK1k731nQZhNu4nVgFi0kwFyZhMBBSlT9
93WbsBt8MEYaIYp6uL4Q6zxJnkSEnBjVmWQUhu3mV3iURFlvUhHAua9cfG0AjOoUAkm8r5X4dvEl
ecPw1m4btaCFMj94j2XowESML5kxbWrQiWv2p5Qbu0hM64a4heQELLIYXN7WDaNQXtuqAVtwyIlu
jHoD+TO4YZV3fTY6tX9pgBzKXO8kkffSLA+SVSwpJokT85KHfEsmQNOXkxHC+NWe01g2M3QieJxj
r5UcgzFFefFCIpmwg3XbfjXaU4Xd80P7hEvPLB1ofefug0tueW/VnC1dtvBRHF2qJaow9RJP38d4
12ZAbnDq53lIPbHRrWs0n8Oo3YQy74gFyPYYv7ervTumms44SXDAd9tb48XIuZSQXxReDvYoAfPU
HgCmjF3FAiGNCPg/OXtb2NHsMiqlQR371L9UqNv6RTZ3t2Vxg8mD46GGoXANIYytqYHs6OgG/7Lh
MBKVj9oRr2TQvKKwXg4rsX4Z5fLBOneZBCEdYVdlhosg0PquEms91fISKC3Sf6EcQUd8EjhKjNNa
RCCs/DETpEplZe6Jnmk6SgQ9eQSd9d2Qj8JW5Vuv53S410O9WmmdhSBvi24pjyrGHc6pojKZZ6v/
8emsyw3H0XaV/j/pjTZ3Rw3LHOozXtJ6ZeDfN+YHsbb3G97fOxwbLw8X6XKNBRp6gavxelLfU9nm
nW39D5QbROdC/0OVwdwJyL6x0qNfsuWQW3EL/uLE0+Unx0YsSD8kI4njM7IjGlWB2xcClM4AxRfu
kkxDEa+C0+mAKf2S2kmbwGeANWPEfrLNDEhKKQBu3OzUJc7AWIU4+EkjzVF1VuusCh+eMVxngujE
0VinRNtdsvzomLn+eHG3uWur916pKc7gDeukCCYozrEn2LyBL8YY34XSkEDYWm194lk1XIP0pr5m
u2vkjqFh1J3WBKgu3DceMihHRDPFU3gmW3XL3s/qtjsF3BhdFLipVIAWCe1WjbcAsrUz1JPmDhSr
eVkWxin8GDMk6Wr/q/L4xUpS+pkAwMeUdZ36sn6Ui4cqqp2iXBbgBG1MPuQZlPQiijPukrwU4EYh
1KctGTuPaXwcZhNGnuMBY0/3UyFUoBTLrw7c5JN1jW2+2GzPFNzsnWSrlbXeXoX0OKQbZWwwFcT+
PswffLvbNF2Zd0D8voiJlLsDUZGMGe3oVYk5OFfT8M/fU/yoEygPvpIPYTaI0Tl+KP6xLSldGFpq
hSZjD9H/9M2iWUJyvSAZ4scD+Vwz5KT2Xa4pEzOSKWux5v2F+uS1zjxpAJobJCvH1/7OSPThMg5P
3mJqro9NVPcTQM/zIeO4zU5yKWPuj+owneu571iad4wKEMm+y8n1HhTf1/3VDOu2d3uS+afIV+aE
ji30GHI8d3jWU/jjT7gDcpJsKZ9cGOOVSBHZ+NXtZM/8kjqHRUgcCYlXkWasIEE073tUiHvsiNNw
F+KNWRcydxIWK3dSLvef3rXa1J612JoFPvMqhqa8R6GiTy6HQq+hf0D4UOWzCAax8L9iH/2Bgpvr
3/PaOTR0uPUrEgof7lZ5QuEMwoWyV4I/7CxxD8NQ7ae5TwoQYTINmdEvA7kwUdiw9B9NsiENuivo
t0kpvA5e8GiPfNVTCPXUpXuA3BojIePpf9PNCd2mL2F4RHIJGuzrQ8t+NM0TGryrr3iIQT0SlY98
Ul5qLjMOmi42TpqXBRiqas+7X2HKntr3TSEsiVWwq15JY//DdgjrBOKfyl0gp22UDfOwQECdOVGt
M4v6ohS8hYvl/2xCNA1yFsw6FqE3PSFpWbrxrx6iFDiuXkFN4kypatXf8lIJzK0a/19JsTwL+HE0
pJFeOdL/SwrS+ZUROq0fvDGXtOr7XK4mVVOUivn7XSUgchQJv8y8lh5bIxGsErC4iA/ZvlDM8eT2
DTLxdXyzXM40PDxgjnHFSojCMd1sKrpyBToG2P4M0A+voO+9uv4qYVKMG9pkDgpQDdaZVU8arxbs
JrX7Uzqm/tmYcC2qeKUns8DLQsNq0KyqpwysjsJv7wVXxt+CjwppCqAXRukY3nJgpIqeVg0LTc9/
qgYCh26VspU40vLiTPGoaVZm77Qqtn+O2ts8Zl9sp2ZZ0oe8zLXjR0axY1B0dP79v8Htl6oNKvj/
xqq+lZPuu6WgXbhO1FmsiH/3QeAv2gX8JHs2G1rU+8LRw7SOizXJt1MI4mo+E9sofLhrRAmSDXQS
uB7NSPiTEGKbG6J7n4WCyEekrvnObuUzr0DWled19BKemOgLiLLhCM9CIDSd3GWNtgy6xdZI2kM+
iEEsnVGpHUMSyUJUAc836V5JOh0pToPeIrA3xZLEuA50H4sn7AYsjDQN3Qxf9ZFqrVql3Qf/prfP
NRdLdiuxSItakqdLtBga7bIaPAz+E6pNH9K34t5GWrqPaORZvr9NFuOvDzQ6rBdOF0y4P64m3xsu
9Q6/b15aSocRq2uU7wL+Lzju1Py7YGbGflxMRry3Iqc4SZ29c0oF1I9SxNL1uOqmmjjofWlTm5Xs
/gVYzJcaJkabMzA6WOAGiN2s+tDGmTwLeOBU3u8U3RC5/kuyQChBaahYxxdGY8WMB6mV9T7Y7V47
/ZdK7AJGzfaa6BYbGRxyK3Ys8+cxknSgI713c2iT4/kPAZQhWaBPZLkO+TKWrs0fB60WhsDH4ESy
3QU9g7OE//QVBAlk4TUOwOKoCNcTJsKTajO1UZs/rLQYkAPoec3EeSpriXTOmZyA6TJxECJeBq4F
Crz/gDQ9MN4WbTZ9Ap9A+zMOvIop2iHDeV3H61nhh0GGRTl8bYmSEfetuUxqC/E2oJQ4zLLz4ofM
DgJ6rny67eUXAvqdxNXuXNiy80+c2sDWRo2PLOvi/kGjF4XxWmiFlisVwcHv1wQso6iEKBue/hKL
7s2XtUGhOhJws6SS7srwyLskbd/JydYcRRqHkaY3+Llgqg0EmRC779fvi/abfIBpr/R4SnsOJl8x
2wmbYwfA0mhaJcofOsQf88PyxXalMDe7SXXcPB086cYq0CAD3x99Fa1PGWuWLeVOdtKqR6dBrbCU
NrpX5UgvR8dXPt6C9+mTaT1raW4CKD9shWhvFkly73Q4bkGuHojmQQ8Td+by6o+BE3qBpUal/qNX
dU3sRbyDAjWt/7egANRApmHYmKTKsJsfR+JXElSrxvvZvey5eE6LtLEBZN2Sg+jpP2Uvhfr0Bkzf
0YcZGpH2hW2qV8QZMGFwBmN6bkjUUKDWuTXYUu9DauXCFvhI8F3QXmZyCkw4Ipt6EqWiz9wPpy0Z
CFT7GjTBuElrpulCOq4Sb4/HxGiRTpLKwcJOllfbYSIBxh+4lDVYWg4ax6OcFMcSHpMiCnD6frWI
VanGrPCQzH7mg2mT5QPPtRStgBS/34QKSrn+b1jL3SNSXSn9nOhp29NSUF/kjAi8EcqRhyCPgk51
MpPWcheTc35m+ZHjrvXTj8ZBegguxD71vssGEJTGnyzwg3+ka6ReKjdoWgDa3415iZ6r+LIXrnzZ
xHnc5oAv2MZBwG8gt9a/xLmdrvdhcfnAcJbN3KHQC0wl2BmhPiHiweF3GbcNQlGp5Ib4u1MiZXTw
IBKNISM2BeLcXeODNQ8b/D8cHXWMM7xamoDtmwiUK0Dp95/Oyy6eHwAYtaoP+mch5FNLa00tbj9L
xeIx/hRcv99NTAMnll96WyFEcl7eIxTkP7e0UmFk6qeDjdxn9VAmIqTcVj7/XpEsacNfK02V9pup
9I/h5qzwaoX5hD9upVGk8P8Lw3L9jA3oJoThAl2K2Uf4x55cwspREmX+1WpgJd7+sWOu5GUSIZex
/z8X+LXOW1dvKvLC9Vap9AFCtzkDd0E3s0BNTVoqi2hKnDJyuKZptMptLXhEL+oaBOZmifErW4Ww
4eAUUbmdGIeJS21S8nw6JPeo0iiga2XKls6vIA4vxBrh5SNANCBdkqhUPLSSM2rnfA8leogxqwGZ
nm4D/ibGXlKypHQ+oYjLVl9LLHAqMQtPgqh1E9BH73X2PY0CUse0F166kS7eQMq76Peb+8wHYk1b
faUiC1a+hCDEL3gr5C45G4wPYbzURDeyCu2VzbT5Rpvl27oAcrW+WhdoAtCiIedna7k4zCWlq0Dt
mP/o43niaFP9oaevfT4IFz/8pbp2BGBsDiMqM+rzoQhKzgyBCNxEWG87WUlsU8NNarWiL+eclpz7
b4Hmw+YvChiTWVsAe9oYukBzUC0T88H4fOmNoCXkfTd2Smxcpr3oZ4s22n9DMoSDgQi++YcXxyZJ
wbrRChysRSUyaOwloGa3Du4QHuREAeiaroUGa2/fpA4XhzNLavkTsnHLXm4IjU48Jw9sxdKbC7mT
IbaMKC4J7PEkfNA8lG1B+m9ECEvWP3b4eFA89CUc3RlFK/UNc867JpuFWYcR+4dnqhc7piPAv2jc
WoBMm+FTLZRbehddRLQ5JlxHXXfkdq5s2OR2/JhwxNDgSAEY6xWjq1WQvhJxHHbI49Iz9I4JRd6W
gU/yWLXr6SfrUO4eu4sIMD+5YLL0FUw7UODSuCPInrfzeh1UiMTJo1ez3KUxyfPZWBa8gSzll10t
W/uOO5b2qsD3lwE5fJxTBTxb51pUy3tLIqrJ3GCBQm67LHWyLeJUSj40DpsZoD1dWS11BPTAKRMZ
o0af5tq8ON6S+9D9s4mVhvOiLewIlzMrxzxep43np003AerRhOzaw3XdI2tx1ggvrSUiTTPS6MAL
j7EiXrnpJjE5a2MhfedukXnqfZherCIjkb8XRBudzDeiD6q9BEspCyZfwgWDnbQ6wqWq6TCKGdz/
795vhDVxgavTGBSaXN0NS7XI026MLEYQ0a0i6DAI1msfEuHd9cgrEHu7IHKpQFzmjBp1KqtLDVo8
NGkpAZQGsWdy0+opohEU/Fm5C+tKgd+oTXPBECMMA2O6jEpQ0AtICw2AdVaehMopM2876z53tnoS
hFdRnYBHQhTToUsuy9dvbShLodC6DqQ3b2Q1CILUbOOuoH/oFcQCP27FQXxZm0FlTQMKP7NyEtSp
J2LUkdkO2afATM/PjTW2ZGRPky68poaEdPqgN+P3uUJu8UMGavaJd/YNiys4gXC9h+g/VsGd+FqW
VBjla2Zmpj+DaVKFdyiNYXUOv+RK2WWKxfKUNZM7uLhK85++fMTpRCa7VhRK9ZesDnYDjY4t5Osj
2bkFHy4/8jTQiJq0A6cqvtC2eyk1iYhGtK/gSnZrGwOJ4z5zFtX5rIo926c4F71WI4xGJq4hQg7D
W15mqYYUrU5UligjE0bdY6w0lpnyZzadACDcLapcpsfeCSVBltx/uAWJklsRXZT8XvSfktGMWBrI
j45fuSrTOeAwUZKZOKrmcQmbzCK1xMbt+pLEX3MRNpms3TlTaREjkhxxzITSwitEhlzTFHYAUl87
lSYN7QbRZqjBIkPuE3v5smaSd/YZsbvblDANOZq/usRNxZmJ73GCoMxPUz3LmVokc+z7CQlOldC8
+WhiBcGa4C540IPFvmyHDBZYXCeVX6ELKOn5Nnr5QCqFQmDiSwE02RtgrRaSuV8VL/G2sSvEuHuO
AWDlghEOeTohwMDkn3zGfONka6yw+7WYHM2mNw2Pd+DP5I7uFSjZKU0/uymsxywmHcaC+4qttJUm
fYgFdtujmiEProsXiQtkxQZwkuP7BlN7QDDNHJeEfAsNly8MbKAK2JvmQMIYHyA/BE+c8VfylbX8
aZcajhUiHXnlNS3RMr8gqFuuG3PZd/d2XOmdvbT9UN5BVnuUjWIyRTpv506RVm+Hmt6HeJXEc1oK
xd87izuk3xi1PEnhFrL0DMmgzFyHrQwIxcR4dbF2i4mplVb4G4t6Lnswgivt5k1IXO0RO9PnQBVk
VDqc9xENjf1ZvqFO0hJo+g6VkxLC21MucOb5y++6BCIb3yQLDxK0VAtdMe2hL8jYHJCOibov3T/j
keAxdW+Il7ZJDtFZmEKDWCM+MsuLN7LhzIj1aX27ekMT+zdlHYokt1V0UIle6nO4phLT+He2/p/y
PbjFiUttk6N9W3Q7jhRqXmQvrPGTTRgf9Erfbqkvv1ao1MXAQe5Kz+f/JCr85Wn78f/uORw9fuAS
w75xycqXRXBUJ4kKP0oG4KrAn6QvmgBwvQJUgotqsvlGl0ArXejd3G5rdtJ8EKlbyc8w6sqi3Xal
RQgpS/yBr44OAKh2lczB+1PFw+acnA5Y2tEomXfNCWDi03D81UC4+XTsEZE7sQx6vKsbIBpyWPnP
JXVKJGhdgCsqlR6Pn8O/0FEs3Iq5o6SRfYdOP7kBkL8QB8aSEeuKH3jLuiu519LxYvadAH5CmpbZ
tL4KtoUVFEMQnAqqrgf/B5bO8YNmV8beyVt+D6Czf7cWA5DCZX+BU8BjG7CJ4Dox2FDnatVV6C26
/THW7O/09jQ3aZHZ/R769n6mXD2u7J++aK3bAK3/FY+qlHjDDzHj50Z7LnRZ82uw4xfgE1Is2hCZ
3WTc235LksTqS6or54bKeYdcOQ/XCIG2Bcj9p39g6Nypgw+ykXtdukUieS4Vf1stwOOJEfN5y1n6
V6sTay0uGfFZ5DHlzC3NuQ+Si5QxNLvuWYXNPyDlq2H+7+rCAfRpEHa2ZwLKQU+wzhCSamzkTQcb
kq3OWc2dCpmuh2vrlShXMfpaYcqp1YXhj6rVfd3ozg2/8b2kl5tKcnFcKCSxUR6xSHAtwATZ+Ihq
KcHdOGL4+ozkEzXCXTtDGpC2QJzUS8fDCcMTpUBVmsn/Goy0wYMAVcgvk2XvkyTueSYekmaZVEst
UXayE1EiL9oQop/0JA30TK8fOCNoxeQONH1CfJDxgb5jB6tzk0muvAwAmk047Wb8+GvMd47ViFNc
A7k6PEBNSZXMJQlL7L0M2sG4q5Dhh6OXsNhQnutkcP/RZoSQTolQwPQ4gNTQZUORFpzbLBWDehbw
ed5zIMke+fzbU/5Vy549eiC/c/cknaWyqw7fW5YP+IsOrrBP2Znhb9+EaJSqj9KpQBAyjsb8Vb5s
/OG+xJjynL8eFBtamirckaOWWwnqellH5BvCxeUylpR44QmopSf5timC0j2O5oyTj5gkS8rhxVm+
oLrXYsv3Ms0OEDX2fvdjQ/npfgtYYn24r+tfenDs7p+9Cozvdocyn0/DB/xoxbLMPZ3xbm5WMcnv
UQKuAmJ0NKPofTgfr5dFwIQ+/UJxAuogrQXden8rOgel5dDza5tkavvIYYtYDSqCABJP6kVB+xks
biKSmVeDHYZU9cH1CNUGqV1eks+Lk5aswwtU0PIoeMNMsEfDYebw449rBDc3zHaHAbX8irL0yGtc
o0Obx55NSqCNpgbvTswCoW++uullgkU7Wfxe1yR0ifD49BojhgdMt+QZTMztFYYBZv0x8VGjbS4E
FAw3dMG0rou7Ol4o7zp//ZpLQtNLx+E21uLCuj9EadHnQxz5SiX7mhPtkwcmtUUSpZyyZkvBWYdj
5xLhX9cpOyr0KD3EDU6ejmrc31IlVYN3Xp/4y76bX2jedQMTQOEcDStfe3Du3JQt7a2to99ygkgG
yi4ee9SsSLeKzWPDY9nk3K+qn3PQL3JKgju8VWog7EEPIE/yP1gjOJcw1s2SiPqhMEXAkhMo2byc
qHxlbBxGzyywleDZnvWJ6GIpmmWr46rcEHlq1sNedm8cQ+I5k3VihMa1M7q7rYbETpVHbBtxkO+L
EzcPDg0EByjjkNubXyg8CNSIp4msQRjYWRgLWzURa25pPXh1mDVymMoI/wmCrUTDLRQEIC5+YhwJ
2AHh+kVeuuXx8nXfZ+B8kJoZg7BszEg+ZPhKAu7XXoRQfOEEODc70rbCYfYjDid450UMyJgaSUpd
AGZufC7QsJS9ekuEr5WVfYN+Wl1c6jB6eIhhbcnMlLD8DeuYcg/PkDDi8vt7JRyF9OCgVr5vfs8a
HrH7sdMQKXu+P+bl0cLrKp9+yN51si5wrkHlwMC8Q42cN+1BLkBeDyJecjFU70XLmhFnpugdnPWd
CIHdPOE9WoOhGxvSzfLeG5nvXDnLMnD199O4xgGKKYH1KOxh8me2lghIfqjo/UNojAWtVVXiagpm
C+ostB7KWMz1Jt5gSaNA+E3p2VRzgBaJdwkO5YVTE/FnESnyMCm23oLZicuK62UDHGNO99ejCKa6
VvbeBhAMiOgF2OASU+KzvDokEKWSLxqq+5rI2vxRQV84JGSvKBfy6VmLlzM409bJjqMWGWPMynXQ
RfZ+QX/Rm1YFd2EvVlEFpNYF0ENxaIFLzqRYS697onAEYF+zifJQ4L5okJbT0b1zot0qIx99tu2b
qM/B8ltcUpKkBpBf3KYFmPVq0MeZW2WdS8yZiSSK2aIchphQ/tRW6MRSGXUdzqYWAZcZjwuVovYM
kswNaI0mRtcN+EUg4tfP2+jIxqF3WtjWMw8IzgoD9pQN1OB420TZ9HFQmeoqx1amh4LXTNCsK8VG
1OdfrDe9tyRMOoauF5xH4LqJnJ4+4xX/jaNUyWMrAzVh0pTuQ0QN0SygiyHpVxAKVeIluPeMnfAz
n/bChgV3U1vS8KkmnZ7db4YQWnI8obPQf47CapgzOw2Rb0EtX6oXymn6XCQ0mt2SYVn+6u1c5Rvh
nGxEsljRU442enRW8S8+alaKf3eRyLyt3otLa3DwqFnRcldDWkz+Q8oqoPAwg646RwBa9daYqaSK
fFw3gviRnPK716G3Zes7M/2fXToV7uekmvtTTaATCQK+GtWQksVq/eWCGio2J2rDowcgG26llqM1
u/lAVmltQQURBFMQgPOM4e3xwdQc7uUqVi5LxNxBopkC6fMWDO3ymrIvDfu5x/0Nzh0G2Kt3W5X1
499FubikftzebobaKtOb2kKJA1O2OpAAVwIB5nqPXmiwAtf36h3rp4R5Y1tvagRioA05XxeaXpbN
KWWygXWsU9kW9fKHjJODC9YnL7EXsZYDVbo6p/J9CdbPo9ksgJYDCL2/8Ww93Psy0wbYb972X/co
h2E3SEJC9cGvkFiy5OEgAB66gP5b87br2HCCK39YVwXQNPxeceJkRDeRPKbbjzPs6QYmhCQNDDtY
c8bjoIiBEK4PZDI1iCpnWAQAvd4sRR7QQ+ciJLFDuQ0hBXItRpp3wbAShxAC2M5kDMXKH+opOPUd
dtFDzw3LdliP9CCTa+h8sRBOgg/QFBV+xFDASGy4dSIEy6tMmwZafAtfR9ohdZYiKbZvReTLP+73
6TBX+d9wMj8lqDyiy+MWPjuKPVB921AVAyIPDGLHU4kpNwCtxyZXnI+RtGhZWqFvsUVjWSyqONnH
R47G6FFILSBEHnnMreaiDFeEYcA5NvQ1JWZbPiGZRQxJmspTgGfqEMn1+qpuPZHdfCK5TKKgc+QC
xXkwa4iE243QEDSngKrhJK2Svib+J4s4ZUpidLycu22hYDDr4zuVuSYftZy1E4qwKAvjr3fa7dT2
xULQ4bcX+kYIes3ckqkcak3ZTc3H7ErvNGe0b0Jtl5R7GmjANZxJt8FLXVU2tR606c66ysboHOtb
WrDc6jrHgFWpFTZE73k/XT0zfg5Mf9vDZ1DLEGYv+kzVhvzdtloqLgGqUoHZTRaKK0i+NSMeGzTF
Itu3JgHjem43K11XL/MgboFost0XKNoJvN301sfc6xqhBhYxQbZVp3p2Q3OJTKwVORm/TU3Ho8+q
GEY+yu/R1RJfYtYNrLpWI46aPLoCGmRZ7lWTkjg4bjxm+lhxRVVT5A4yzfTf3hAnpgG0HtlfwaWY
H0/lTulnvThtk84PZZD8anOE+JUhoErhwJuzkwOsaiF70xdQyTKteicMI01V9k8TlhPqMPxgSuWF
9y4LZzRLaXPvf7+0buvpIBvjFbjHjSWHCl+3nrWCHimzzyNjO082sH6/xAJjFdilsTuDwtedwzjz
IJvoZsIE2QDelNdLgZ1Y8kZ/smieDxrhzJjBiIS4znYo2sPHL2AGRmvUwpvoRZyT9vSgDXm2vYXM
H9fDt2T3NKafcwZQ6VnnWSHpB9G7YFZBFfxVxVP0mXqnSjsum0edP4FP9fdFbDIEocvO95NWqebB
cQUGTALfA9QOtD7IX2Iwvffe1XO6yn6RrayB/Pv6IpEOa+TkNg5dbVdoL0k4UQgyg6Gu+ZHBCqXz
EbQfpoDVfBjnMEuwqVeifRUmWeGWoWZN99OUJTGpHlyQxZY6+NEU5BFfLOqUi82USVP66KnY8yJK
HOr+aRbAhukrjS4+lT3gLIGv0MXj4EyUwLxC/jyFfZiAv7wIckQ8T/NNi5KW2etaDdj8X9mFWHj9
bt35aTxd+7rKCt1jq/yidOaworYh3nZlGjZno4fARyDHCRRWl+D58Io/GC5/btWMvitar4oTb88W
NGXQUH9YVSpqqWjjeSl5exnL97ifhl4bM8066Hmj05cO1aS3jZw1qgWW8vXcOw7jAKNiaHN8P1zL
HorbrgkEZmSY4DyNcoPJ4ugfOJKn+m4/LY0vGOzUDPRct0Y1vY45jMRP1dbBNwFJt3BGWpRycyqR
chzJZnSoHpTat/V+UjdueiGg4JYSW9eDzyrl7dXuw86KnAzzcWcAOxJVQ4EvZViJpM8VSFChwnt0
XfkPggT1OcpXH2euCIBIlL9YBy4FRXZl5IfBukaMHDPKvIcHzGnAxB20xhzQr2dxPREoBlh25pHu
5RaAsPyjYdbGj9Thf4kEf/ma9gFlZH5LghNcFA1qPuPifhUQtBPfbFnr/nFcgH0Ww+3cjelEXlJO
KeP97G//TE+m/kSbNyaxTvIlJ74C5Mivk3+D/MbP54XkUtSimi5xRTaLYmzXnODh/bCP7/mShUyr
+sX6mZDCjfqtTsVbiePIr+3KdhMD3/WbJn/SJ4JD+2UJDJpA4kv4lrBVNMy5zoVU7WD90EWNkKzQ
lo6WyD8NRAnjSK2HQXnhOSITYhazWHvRvZ+Z3TKP4kuNBzh3rB4GUMhtmHWCxwTSOg8LCi/ELu+h
7+oGYk+IggN4boRalK9HUtDtjI6c6aYmDnsr6gPDxfcOW3YhLE9v6O613gSoqaJQHungRCUSGB4+
bWL0/NRvHqbIbfEzqU/Dj5RH3wcRHmQMfFpkz0nmQ4Tv22aaZNBPF7Jv7OUWtFufj4z+YWdMwaHt
JL9aDIm8HnGDzF0WpkXLoiKBVA25Q+OLfZ6c5+jnMt9RPCxo9K8u/S2wjRDusP5K8vDgY2hrVYMX
/6zg6uwoyVT1bFY2bhts9MiaPgEjZvPUNd5H5BoLSlSzY2hZgU4wmxQ829vI4jAjtNNkamt1zun+
BSMhiuFWT7rk4JnB0DyU1UhVL23mwajluQQZ2Brz6BK2WX4s6dZejZCkZKVYvLroYZAt4dNXwmyT
9PiPBXWk2EXYpmbFMqZKorASt43FNr6+C0akPa/NN3ULoBk+ipJzFlneWlCojXMxbvgOZclzcrmu
urefteSe09tE03uZFvuBVVYW1gk5NQTkarL9wuX3ZUDDyMVlOsSHMQQtXFk50TaBY1xdM5iFhE5U
0xcKKnArmYgA0rYsJsb6Fg2WGG702YUupLFkmZJPTsx2htdCiJpuTzX6vest2p+HuYfl7Um6CoKa
5eio2d5vi8ObNPWqWCqSspeZH0jOHdvpK+8B0/CD0MxevuEmu/Ip3I0AzXinfND+zCUZTo1AMEpk
OE42uCeSZT6weAmj3bmhJChu8INSZx+N3Br57t+TGvyHel2+u/gxAIYoy1hl2fbKiBpmcz6XKSS8
qe/0Z0crJwRpIE2P/OJH4aCDxtWpxPZ3MstefnAsOkrRR6wmRQYDRzJSX18jFdViI5MUQ3Q7HF78
xI67RddiY9QlgCMO9ohaqvwHBrRSODeYopgQG8yDXPi2PZT6IDNf6SZrtW2mzUwFPLSTCp8Cx8ZX
a/c0Y+j5Dtdm7fw/yIZ16sLXlxOkAHbsK2RbyiTqJiz2D/+W2YmPovYctw2EHDoev/rgMRZ8vXDy
bgNBvMuvlGHryYNFAw1dn2GN6kS5bwXrsLGMYsSDT4zZFY5yXMB7ZS1yyuc7h9MJcYv6MMZMt0kH
F57LRpesqnKdf1P/tzuIkHAl+NZK5v5PhT9S1MVLDxmiFWBjjrRGMN2pFCHKvzmSnwaew35JUSmW
Uzqw/AEcwaIxIiusJUGQ1k+d+bMhe57Jq8MlW/FLmv+ce3s/X1ccG0IFAMA+5hgEUtfsDny9LqMp
GyTYcKY7PT2djsfsrRWXIchg43jRtn+3r53Q45NUqXM96rYpbLkUUAsdW2jtX62rJjBxNRlR9YuV
Z/KZNU5seLF4gcJRGMTuZtiTlXndnYTm5Bg1acmUtjD2AKK8C/ijy3MxINaQUeveHSU6v6pS1g3x
CpwYe6bZ7f6tZZ00oDmRJiqFLEaK05VeF4Ab9L81hvwqYHGnXPXrfZDcsukH3pxpRl6mmlriEwHU
ybI2k3lQuSFv2nnsge6oktgDLD12TvKFxzCCLFhC640tKC/3nTxDZc20/SzMuwpMdjLSpw2syuOf
O3AKgn/LeD7O0AKqkXDQc0v/S8eDHMrdH3HRd4xUm/OlPjWeekH4yHRJ7oktaMG8NNz+NFLyAIIf
ozeA3WOFH9FB0DqGlZmUwv+qj938hFWiDXPpjK5+51775t8dV6bknhn3pU2B6JuJ51rkX4A6Kpqq
Zgv3gyiADapRKxCvdlpqV01YYdTcBUBmZqNtk9ncAwBa+PPW7geDXPl95F0dGDK0dnMfhUom2XDM
0IyWQw85mgvh5O7vzMpPACat1F9uiBw+Jw4CstUF4f90W1DBXL7+6vFvuR7E6KifbKa5awSiQfmH
R38La+PLCNuMrwTr4U4875p/uHWh9AndkDQLD2parFUGjEanJ8irz5isHF66zr5pHW1M2V/9iQYe
Q75gsQsXzAxpQSW5wKQbsc1m5WFKxcjsEybJHLEPBwU2D8gTmJrbSKY4uDlkNLOhvOt7We454SjO
umnRYKKoNB17ZDNaC0i9u07FVprjIync+i7DvvC0/e86weI8SSkGSGDdTiSkTTF0oiIjC7oG2ah0
3zlkiGFhht4JP9q8tnDNI5I5rHJGES3a+BwVp8nl3iShsaQK5YsbC0HfGQj6jrok2LeClHOPjOuD
qhrAlfNAREAEYs+Bsk1boBrW5jySiFMoOvY4J5RFy1lhyrs1nPyFgjPbe2hwchZqo+5G9JuGa7Zo
qqXvqT3+0pIuwdktoVwx9H7T2nEt6SDMjWy7ifHN8FWatSvq4Mz8RwmF+pCuxsiLPWMg7GrHCdvc
jgdtAVudNWuUqDovhK+qA/6IsKWAEm3X6CKvEIZTs5qXNMmBSrT5qSWc1UcRqPRm5sJGqQp4TeSW
hJGbRY/rY//PQyzSShI0PXKzefersqE4HCf0w0WR7OdZNeUnGeZzGOlGRPkV84pQwwKyNYGgs4Up
8qwpoN+k6cqnwI27vvQp3xFASz5XJ/Ylan09JgJJqJI4ZY21H3AoPX+eREVirpZlylvfXcj2691G
nnM6qQ2dii3p7XG1MX4T6xAmgSLDI1qGG/6sm4JYYqkgJOfChpTbD4iTtXgE487uscsbICXBAFEw
ftqS542k5x0LBv07ATxwQZC01Uzoc0Q9XSeK+xCQgXhMs4cqk+ZwWNbzzwHpww0G4Nvb16/kkZ2U
hbPzWfg9vYzwQJzUvI+BeWQ65nW2yif+s2rC21Iy8v2MfRRAwYQie3NsaGHSDUYVM88OlG6XZHG9
UwL55/5dLExtzJXdYVwh/xX4vXAiWe9bJC5ZA9W7xgChwoPMCTZ8bR5Ea1pJTd8jmiprPuL5nQH4
ufKl6HUxSYFyQLwbgDne657xsE+Hilqvskwr5hqKkfnnexKavTJ+VQW6u4SFhYtS3dyNyRlS09UX
5dSPOSv8SK8ssNtDg6Eq1Yt8BIysehxKYsESE5z/CcvSijteLdaF/M9i6d8eVI/bLGRxahLzvBN1
FNerPMopbLOlq1MfE8ZgFHXPaz0k8KSPTeZSYxqRApFCxv6DRducClcuMM50w1P6FowbmiSjy7DT
kf4iguYqDltUCGLpLDevnlc/6UsEDiQe1mLXBIXl6F6ua4GqyeCwmtbjoTMonLSIOZLIWHlXbEsp
Rt0Txr0F0YGdiLU/ftptNJN5TM9rCtRXsVpanWquzU5pWhc+bw1Igna0KZuCr/llkmGUgQWze+2C
MaPzuLD6gbtT45K+9OiDORI/qFNFR0ZPXCme5xdxlsv7KVGr9BbtXGGiPkj7yJB4K0qZ18fC1AIp
MeJXXWXLP2hCZuk77JBaTJ4ue4bM2YUGKL6O2gCv48BaR0Ba5oqvQz/+du71unHVY0Ow+DvcxW/n
tGMMY9RI60zwroD1HOBnyS0VYSAd1znAj99jkjr0QtTd4QH1Fp91tWaMKXnVBwUd1SAFsln6Aj8O
qGGbxGeB6Y24Y7BHJgLR5A3EdhMn/za7HhzMAXEZ/VHO5asMd2sKurty0jGOcTSJZHpvf/Mdrcap
a42puMC2bKUL3Hep8MzKknfhFt23SSzIyV++6BK73H7nQPss2jUhtNEo9HdA8+i7mDjG2UUwfNxw
j8KPCajlHUjMuAQFXdVs0RDHbWLO9+ryQpmF34MKj9LN6bQRAWjHtqESRD1GQk5B6Im2132YJvgm
9nXGrmQohsu9WXBSjQdg+3J3vXySWXfmnDsJ9rF0IN8UPsCXyEEIHW5SaWyZBRMkENPb6cy0X8iQ
RRZKug2Yg+r3IuypEU39E/qYLNO4yKF9sMPFDTOe+IgQJJGfCAa0UrrhsVlImeVesmZoiT6UkYsQ
so3fCMv2O240qMBfmup4IHquSPm6K6lJo1dSfD6xvzY1tBXXfdb9B0nAhhiwbun1iJDKF3z7uJN+
0+5Q7djtgRmqp/4qTY45QBzrZEexFESH/cPcDIFkALQ6YvrZ6unqRmBDqf4mcimjXhrOE7hpnS5r
8moYds8s+sqHKwit/gsY5w5TXQR8GzNWKRXSF8xr0/eEr8gPMq+qDyd0Ng9KocDzy9zZUBGlJFFb
8v9xtdguYpa7TPQrqubraxwf3lKq7MhcLk2OYEeMAD60AHVUBJ+eSP65SoS4nkRGD95hWCJMDxQS
xTdHQxxKwvucyZZnKDrXHfCdWXkbEgftASRdUaftOSPuDhIBiTf5SVHhjWobNhXWWNjtt9C02cZI
lhEX067Fj7OH/Ey+WJq+8OnXjGfirOH9sGrDm5JJsYEZUYkRnRJ12Gbl427UTWyeQ46Nq4pVY+mz
o/W55UIRV/HPKqCQlLRnEDfYCaUoNKEibNnTrHRr9W7wo2ap3jWkpk5p90HKC/yJzjCnta+gU24W
US0HC0reDctQlSJmPY5vdyMMuhsPXsfP2/vqCl9+CHBswW1gtIJwyQ2MpUg3DW/TOKLH8BWjYuuf
zbgB6Nog2OcPiwC4bYmuujN8Y31qb3PFE6rqBJj1Co+4Z+c8Ih6wUm19CP7vNG1Hh1G4toSQyaBl
KnH+xq2KKY9xS4kfRnXc5kaqp7pcaWDJBUhGIehaNuVXvpvD2VHSWIlcispumidNXquKfdq9BDPy
rwF3zxwS2dBulP1zZk0PCDXla/2n8SQyTXmqZRFe8OsvQYAx85P9r96FaISnvtcSZiPWnLpwutGy
/sHO/QngIuGhC0wSsbF8vCwQMYwyZvi1hW9MsWi1+L6yOdVczb5KdNzELVLv6yfMELMPC5wuzBDR
rHHInCPrDspcrQghm54Hho0LwoUQBRkpVNhPLSi/n8EYrswOXJY3FFIkXDi0SKvvSolN0dhnX27P
GIExDO5lMuz5zt9WifR+V+i4fLVNZD4HtADQlgKVV3PfJFob+BYr6DYswBjO0dgxdJSNvhjaA7x0
vb1ZWo8xmr6gRsNoIIGfSd0ROtmvTCJUbRw6Kx67JRBRo8AdHfJSCPVpk/PaaRyTiIwCelGrdVOK
5QxGBctHt1Dmnw/dWHtu1Ij/huvtax8+5ePqF26kgzjV0aNyNJNctxgxnwhljsnp1B9+YgqZK9HE
8LYVWGwXemCGR9LFGBoAqIbRUNI1q8irrywrB/ghzj7+VtkxTDYd729ERW7iWSJR2aqMOvLnQpGy
4PqcneN6sRTt9oL7X0CSk7ado8aiIMToo64N/3mVf6NALvCpF1gkiVVYOM/G9wjDJ82zTD7Y8YSu
dGwD+n20+Fxl8GzRyR0ehd82KCJj5fHMeiPjiYRRjQMgZ2PImdKon7qke3pUaPzHFAboC6ziFOCs
MJL2oGVg8SRYcU+wF6LX0lIIAqTFUF/jvPPDAkHhJNT8Me9aBirRi9+CBCygGwPwhSZsckVzSk9f
npBZt/A2YeR+FR2FeOp/NvJdAOm8gqRjX/kpAMq37Q2ip/cHbB+kQF4zzOX9ncUnycF2IlGmxSMN
pyYXkNqU8bPvhm9KXnL+zJKCnJsFlXJcSqPgGCpWWK3Q4x+AY+1AQ4AvRTCKlg92Jp4L+Meg8246
rqBE3NRXur266K/2ICQgK1P02WVVjFFy498n5EbqnD0p0RB1tAdP0CabKvLiF3H669zoCq+JPhix
DK0hL99s4hO45Lnd9RNaxOff1KRSWiRyC1TCg+hXG5KgDsweiaOCOFMlmBiRi5PyBD1M47mwrjT4
ZeeHMWuh6quw8c3DzfQxfy4kUr6lXgf7j96etJgeJIJTOoZohA6rvmeViK38j/3Pgz7FGg/Y0kyV
v47gDyC9yxPffpedBn8X7ok13KyK1n8dlmJSoexfC1ilsOyB/luK7pTcfTbVSCJBeKeUYZf+x1Y2
dXjj2UEXQskiEO9OcH2REejDElweSMou+tWnfUUuwf9oOrZAFvImYKzZjkpqaZQPCBe/VgG5HLV9
n/ernEIV0HZOvYy5qzxncRHzuMiSqkDb/zjR1Yw6Y81sUOmIATw4Bl7MGGg8c2pB/TbZCQaVdB1Y
runfIVAspMIfkKFDG1xMAHFYFFWDm+XduczdWBwh+RFEa4uS4r6X73OSPmByrbs+hBPm6GCPpIT9
HRdqAXuzIy3dA6mBWNe9WeJRVL7q31R2eW73NhFz4gv5fzGLNBhCozMyubXjHCZf/IQQ5FwgyfkS
27934ziNQiBMnVKIRrafWwov5zdGLAMzxq9FPh0dT/jeoDMs3YiqSqZLG80WmmLJ/Co+j7AZ/wj7
H1pr5KZPWuXd9Kda3eJFlhU8yIL3Z24F2meUnkKoN8sAybk5RFmb8gIbxWqYSvZSJndr+2gRs5BR
pm6VKXK2TlRglhz0udfKXjcXMu/b8eubhzd3Q9LRBscAftk52n5C9ITUoe6tNVI/7ViIutQ7hp9o
txXshqTxSCO0Whgui+llW3hUPOZco243Cf7BS8nqeET3tYunGw1h256IZflWgIhsareLAKkzzfgW
aoYwq6fjlkB+piNvsf1BrWMsVhIkhjeL0z1cQURQRWwTvB5pja6FVRTUPuWxRXtKloIFsVrx9tJU
4BxLKnfLx5MxXgRV0f9qL4T5HPMveKqUTzsjOtfxtdTFLIPk255n2YEUKPAdpThEbUgyTF6n4OuR
E1RBbKK7aDpk6azIV8zvhArjuCfcB3ZMucaQC2GuZp0/ExZrKy4iBYRY5Sc0fCJgZprYCUqxTXj0
z6s9i1QKsFhoBXWOncjgLsoCYxWTNwr0GQMq8Kuj7FpxewE73aLBnCsQUbCSZxKStzWrK1eHtWfO
NuWAYAlQs1UPykVWHa5ZeVFmmt//nU64wj1Gz+lwWTEF7rT4ZHLe763s9OCWcjvpqTuSRo9hkcn7
QnbN2be2wbGK1mv8Z3dmDHBEgbe7bQAZNC4f021ShybWUnWzoDL8aFzEi9IUjCdSuJL5rb7IZWnm
HaKCluot0/LcplasnyL4OlWzTr5YKgI1NSyIdUCQMuwCzATHjMrE4bs8ahv49PBQyfSQ9UkWji2C
UxyESHQVWUo74J/DoTNAurqwluujz2ehBQ7iy0As2K2kPdyeAXVUy0OUHoqZIwc/RfhR663MqEp2
aj+G9VjPuwurUgtc3LottWWOJErGdf3Ifr5K5uPeuqaCmjrFhXFQUmSgEj/rCbvFbfofiT+7lFfn
BXTCndFI8QhvgNdDJU3CZjPSNRu05z5FjUi0ot5RIX30l8hU65opcBeUPIW0HfL5CzxyhGfOXCD4
zpsZ1m39wI2dU4U/YsPyIwTRv1XuD4JHsIWhiXmndWsoO/q+n3DnIV8hcM1D48Y5RgG0HTTC9HaJ
30xqK1NmYceQHkS8UgraQMAxtf3QFWboLr7vUC6ff7nslbRk5Rz2r3247GZoB19vAWir0hgbLf20
/v4KjwF/hEqrD4itNPKXVKqlBcNd6jUwoqzaKO1ndgkNSQhXVZic4htl3vvuSOIMcOjItONaaqaM
Jtx4/9EaO7zatJf4fwsbuaMPVkGr6apJUp7XsZR0126jU9xK/LtnVk3aQJp4RSMHQ5BZ4z0vluE+
r/E+BuLpmxrE7Iez6qSEpjwYDBNOhJDjbY8wEZSKgKpV8fu6RNmAJDaePMI2iDP5YGBzz9Bghs9U
E++Ld2nlvb0zrBrzyMZND5AFkDy/2dWcW66JqSPZzuypRv6yTjFhKfEN7fDXrVBnAudq3OQ6/3j8
pq0e6TtmbiBP1tVGmJE2M1OAyNQ/kSBWecqEg92ORbjXku9zT2joviT+8M85H+ZLiO+bziPi8YJw
9HDPwCT05vVut1WwUSouKPu632paNxNVDmHi4E2gaoHdIyvnoTlls0gd6Y6BQo9RPNLdg6LAJ63a
bkDIwHiSfZ/CuiEak2yEwWmXHos02ENZ94UQFtVKL4npV/MPjApUYJPC+6CVaX8ayF2s6aRyo5bO
Z1CPtPbsv1ulgofJE8YjyoluH55KDXYoZ2h7iUSQT051YfH3jLuqkpseBm5nGHBnYE1pzo0AgS6S
76XWF+okpxizY/7zsXkyABAK9o62BAIPJe0usSw2hsa4Hy52WER+/CoTNmv16qMeTuCJQO7pepIj
g9n5AhIm/h2dLCp5tGlZ4orwc3gTTW/XHyDdFvH+948RDUC4nmrrgyZyzguj+LmoeE+tYOsrdm7B
ROAUYqlxHUQKzsXW6z/q17jwHgbO3mzXwTwDaVtfqj15oi22ZWC1ClxsPxQmSFXLjrHx5zy/cKsN
PTHOuWqAJM6GyvrmlErf9/Z7VAW6Go9hW0NZFlZXU0qYnCdk9PkLevA/K3RIj8+7Mai38BqceBKh
FOOhHlc6NX2zlPzI+oFj67yxjIdmJJZHKWVUbuilsYh2nd+KtSnGJGDbXBIDVfHaaFID2vyr+khE
4Cg82sKdZ7ha6U/xpnutpM0JXiR956lb29BoppOVvL6FgionhEsK1V5yweVollnVgSDVg1h4Tfak
uIYVzRN0xvAisVnaWdKMerPoVV1AH17PWplZyXcDzB/wtLatgjTs/YFBa7jgL5WzglMRe8pLg5OP
KEYj/OHiPxbVPt2bb0eZNTlT314R33pFx8IS0+4rYvwnQvV6oI5tAjvfNlq0dBxICrGfItm0D9Hi
5W2d2CMXp86C+X9vcK0u3Vjj2S5dnsmaiYt/dop24tGXspxyBvLapCKNjTJDLCJPIABelNecPBe8
oLWAfHilgYXkeycFgX3jUmweG7thaAuS7zBB13OF6ITBK9plt14+0TuReJOdFBrD4J/4PI0S97C6
X/dtwjvcbhQET7o+jj3k9HrPyVY+c+FhmqMlFQCCslHhPrpot7SOe6i4pADlrx2W4s5DKNU4GoZF
hVADu9y/J1Lwgf0Qgpk0+OAchFWvmBD5CqU9tQy4V+K033gNDEUjzGi07KCLsE9wBpGwtJdXY15H
1BqNv0dHvui4PY5ldGc1y9knTC45UqBdcbUSbhnQVBpTZuMaCrUmsTZZaCoGuy48ZXnIHfeBpSdJ
WTKrbZwQjUj8YFWaML526RzBF+EjhCA59nlT37Mk7PNOiB/d+cLwkwfrpo4x+tFLMsxJyRbNuOSV
shwSLaMpl2JQAHeZj4QaVuPA/py7MH5A4tDVpPHjh8OnQOZAUqm+PtTT20ThcWIRFwMKdfgaw4Ie
0gueNrLJxk3Ocn1aFunyGb0J/8ft6cRkXBKLlNeSwMDtUkh5/MJb4mpDcyHjBJGk1hOLFbbfrVLK
J3372HWPLpAW9v55oNIOIidumHTMBkADHHncBMS4BfxOXJP7GSB7+XylvKIzTwE6Sxj+me/B37cu
G/a+nT+HfG4QkMMJ1nsh6e65k5fuiCHsg/n+ALNAMi4lfAey1HE2aJt0D3q5di4dSoa0rsVTt12C
EFK+Xh8q2GqvJs2etpAwV2Cv9Gx+c08DnTVHSrAL2nRrlxKSl+B+VWUHl9ZKyIHtdoNBeBKUxl9H
Qxe4gar4wwiUEiVUczDMJHOvWTuNyCeeLoax0Exf7I09zEHt75JiKZAt88zPaRnYx3C6kPsAzLkF
KPecsqE7V8QTXUyJ2k/UVAbhJ+/v4wCe5fUByUo1B51Rc3Aw7uv123rW77o089AAnzy0oUidxOeX
wVPLYLlNLP2YxBbxJ9Mumy3/+I0aTabfEKcdcdhwzMBGcKzjBUuHEiCsQ6U4FS3QDDzaePqGBY3L
VZWs8rk/Lybkw/awlGYAd33YDc/ToDPySGv9VkHIq1lRpytXhI2OhK0sPtM1g3OXErb+IJmCugYZ
qcJjB4MeOz8e9B4FdmgZNuvi5ifjSKzmcSRx2ro9hh4s21fmR/S4M+c0m8zXgzA+b1mXeOfqWWRN
Yk4I7FKcWrSs6cesA2g0MPi/k03DEG1gkd9xLTwjk/MSI+iv4Qhs9ytUpRe7J59HFTyo6oOrMwGL
JBYbL678VxzA5r4n6ouOGsACBrkFfCpyBYi3Pp8bmjNvI7xLXPD7SDM09Whb1OorDb+RqCZLvsdr
HJM3qlLPt1pjC57yA1xpB+ZAK7+15QPny350GJhZotT0nytXDbT01K6d5fcqwVE0wg1ExgJITmXj
1OZFoE+8YjVZwwhixhIrkCH7a4tzNuVKM2pYdZXlZv39WUa297M5HZVZJV4NANbIacUTt6U43nLP
w3VRDX7h/ciirKSYJXuVehm9KhDSisa6ltIFl7FVzFPeti76tBTG48fM3Nx14EFtMzWmIW2nczgS
jyRA9WWjGr3CFv//AgnYjqgxlBYRcqM7zRPI7AUoqe8ZH2q7loaegNQ/DNUOFRSozMEP0pEYPY4v
FsfY28vuaGKw5kCeU31UPOlk8OIHlfkuFDX5p1dnJjkYajTrcUpvCPmrMHeCTd2nvjoigaS/pbt9
LSI18u5asKPBg9usP1pe4Zpv+tfy2nOmU/vmQx5X6wMT655JQVdRFQYPnakasbMwBjQJIq3rg6XZ
5aQs5fpqs4NrLE9k/jpgwULSyurp90tF88PO2saRxGmzja9FGoDpLh+HsZx41VQSqQ2eFlB0rwWz
TNLMQ7/CndznwfzeCrdvjHW/jdqKnH9Qxpak4PnXHlxItXsUdhbiN6jI0YuLaso8227nr3aZCB0Z
SrI4kCnX5zvNtRL7DUaFnyxXIiXLMXL4Yfx1w1G4DPQTt1KAFOv6Bm/gta436dPB8FH6JTzGJsiU
sr3y/oHIuKKlLVxBswGa5vKnMtNPCBt5D+fvAVPLZFxNBxqJAKgz1+EyNawPxhKa9YccZIpOuSyC
0obSPbA70WTWFJ+meUwdriGdFgRO1UUDQsmtGgDziJFyXaaKJ5ZIz2kyOWZugfs2L9dJR1Av577Q
/4JtKyb4UdOfWgBTY0rJQZ8efiSXEF/XuGyNHVlnIxICoubx0OXfQixJ8QXJZ1CNT0t1gpmKzswB
F93cFLT/PTI5qAn8MShaExOZi+m8xU1KnI9dy4oLSJgi7XLsQqR+EmPte5wZ1agpGIkDZ7yvTFzK
9wx3/2x50EZ1AzeRbX15A82Jm2AYQ4xAgahEh4aAh3YdAlEoPx6ngrObP2JXOiMA1o9r8BBHOpmL
tG8mgi62RNgbrPq04oYzTg7HPIu8PA565NMYw+MOHxhp/7Ho/N3YJLbL/YD92/6nVQJEr5Xjka4g
cKgFyK+8GTN8y8kgPNL4xNf8ZzInGj21OThZhvu2FE+EjXF9uIX+P3kGAo8IaMPRA6UExf9yLMLw
NWOCRWrUfNx2s9YtQC5wBK65yL+rwOgp+CZ8QsRgVQOwTP/4caD5LsvkH9S/7yBJ2MX5pEeJym+o
BFfieYxWv7FxiekYytdibSb2GHtqBuPcatv1NlZ3u5IrQMcbaxTXOnPAUCHVqy/9DFSJKVhMoepA
B2QpHMpouNBuwmELiUvd18HuNUwlcZqmdTgx1kfEVARla5qCpzzxKirGIUFAq9klFKnd8vJEHicu
dFnmAwEz/ZtDO30YHqN407w7LwosFaSYcuuj2LuePk4d7Cygce3hDbeecILHFj/z5EzpICQCLi5S
OX5/IvNw+bV5R7xC39lqY9TOCKrOCI7axjof39M2hKE/kx7tdq15kvaBbU2zNH/ShaK5XZTr3Ath
p0Yx9Q6apQBZPCEEiIra6EPgVrGT23w5Eidz0iP5X+8cNtYj+tWk3/uH/DQdo0DL5w+EKKxcVZ6v
yrnGDLp9pL9HyUsBMfDu6CnU+ApI1rSGPXUYHffoqqsKp5NnDVqHhtyimSHIwUQPsCrx2xVHmW4M
qZbjSLVn8yEfPkSCPzI1AS26/dvZGecQ++3qMLn9byEPuTocaKeb3BTNsmo1LhbwkLoe1F1j4NNG
rGEMsyGfWn9UwrpOB57p/HiXUcPypwLvWgoDe5mk9A4DVff7PF0Iuv2iResTKbin/LgMtrXT7qSN
bpHh4GN0+ESE0RjJzmPhxLWdOO2MbNpWmwRD0emyQJ895WwXwE6IjdyFYq2YrvgtiRX4aonKY8ID
5C9tt5/y0ZH8LU+IrXg3geM2ZT5P9OgKEDpfd3OWZegItXOnUQVn+Pf2u2u8vShkQZIEUZPtqWrQ
wvyJQCJMHs/lHmH73Zin1ScriRAuiLOL6KKn1snp1d1nF3k1D8glIYyxZKSDdYqG/UqGfNUVyx5J
TrLOjpTD6h0s6MmIbokjinGa9EKFyYopGlEeTm8NduiXGLIcw7zUwuLRwwbatueQ771JSTBpXa6r
I6d1qqn6zzrbDbr+TumRPS/Mi9aaITUUZuLXxBCcZDm1Lh45z4SVpaKqZ1LI3IlHcggo6nVShfLP
SIA/8nWbM6p6mMvpQc5yCuI5yyjs72e0PwBoZCbculVYBu+8v7QZwm0mjgZGQ1/V8QwO4zy3n4Q8
PLBQ3WRPW8znP6q0c0IcQO4TUdMjf0Xs/5/+AmSFSdkzD/N7tO7PlJxgZYqb9qLGtu6gTAiKOBCN
RlTjWWB4HizsRo6Y0eczcpwoPCuA9PKRw6fo7CYNsH7pKq1iHZ2moR8q6njOuWK7qOdUhJEbqXjH
fhY/EYprDQOt01jld7mXnzRMYaOEaxhoD/NEhXBQhNh9KnCXm2lBp2EvA7mc+lmJNIXn0NCguPgM
U25HZXQVzHMpcZft4W4gjku8YeVrpCVi8t1mUJGJs3EAPTdX48oo0UGYYg2DTZFKbrAf7lm6iTf9
gOCBBRmZb7i5iadW1/w7YUQ0vfvpkk6OoMBBWSca6uDvuz9XllOkemHi+l8MwoOYmbE2BZwtDMqM
tTE4xqCs00692dmtz3go+MJXRQOPWEmKjv2Hbpud6OppRzv9FrmAe6/iOE1lthkeBwfoQNi5bytP
6vG6DqimNeuGdKV/1TcQXkyMVDRzKHtpufOj6doZvnBWfktsccHNInPcDhpzWabhy/EgpP1gCnMJ
7NibfvBPlsEuv/K7SH3BxRERsPmrnZ+tODHI43mmidlef3Iq/jacp/BTlXo4pzyJRoc/PpnPbn6v
qWLmW4QjKz07x/XR1Rh6+HeZSQevJI7/aami/Kzqmhmg0OD0JtU4QMH60MCPfykR4qiJxoSSb/2T
tam/H/p/NV3rJOpbVAnwPAWp+XGqefaDlqG5YvUKGwEjyynEPhSOzFaly0j5WDfdcY9BXKYFmS5x
+mgXys3Ilm1jOVw/biEQm4hm9C7J9u7fZh2TlmbAl5sXXnOXPACbrMRlLSIG/J5rLDDYpT2pvkoQ
pjObK3mmb3lpR6RRgH3YRdT+vU84NZ3khA4cDYhnsHl0VoCEf9CTfA8nDh2F8q5Rl/uUc8wmMYRG
+bQfhpSFO04O8DAeeGPLBoS+wHpxDKqbcMeFjh6eQm52BI+9a4Jj53ZeAl79KbXfmPvQ4/0LOJSM
ntE6gXc5tG13krVSO7fA2Yf9nUMXPW8+5C6rkFfR/eRm8WFYuYnIK7HRfpKu+63yr1H8WjkbnWe/
5cZ3+cAMJt2gV7jkXV6Mqk20RoQdWj0oicM9jWRvBPB9fgbhf50ix2jVchvlsczBm8IYmVahMvgf
ZxF3aOZA+A9pNv3iMhW89AjN/5X5lZBMQAOdopxXDoHipwssHK1GvxQupeBKUIP/tOz02nLJZLCZ
pv93o2HEk6K5RrtnCOqliFeY4urwRwJ0Ba9QdfrWMOQeFbhNqukePbPCCD/6pt4vDKYrEQoldeBy
fdQS2NknGBce9n8nSCpORBWWFuvfO+UfmSvpm+fypRzufTpB4dBuwHwCqWBNpDEWzL8DytUO4r5R
qx8i+P6qQWCYu3ioF0j3PgE3XivhxOYDas9wbrR4uwAsB5bv+K7zvEWs08n8XkDuM9Tzgf8+3ihL
IAyieqZy2XDdvv7Z6EKgqNjEFhsXygqptp+wZ3+kjV5B919OZ51Kvs2zuThudDBjRx3pITOGJ4uh
ggfXD3fA6T71MkivDW3M44ZhmR+PjhrjNWZd3cqbBVKAjdv+KiBTj3loM/NyhitVo5LCeXN82g3c
+iOTRFNbT1i14gNnHuycDnUHpjdY3g+KGaiFNRxTr2+R85WGYLnc9xulAFHFp7/K5DcV2TcaXCI9
CbzXMWzhdSq9DqwuOKYf2IpZEjsPKSAI9cyY85IFqsiLdMiJAAs3zRtqMobnS0PUfBHYyl8GBXGk
njy8irJTmHYMwv1mEElRsZiiwrx6wCjgYkIpk+ttdLRH/SHETwXbafpsx0WfQapJU5JWe7DK/EEl
BxUGipLFpUCOcX/9wU5FWxPInnHr51DumxM7d4IC7Hz8snMwF0krYb0lFJ20XTavQ5QeGdz8jahp
mPXhPw5JkdZMEemfbGMDBye6fV78kOH2yMYTCqoNwx8rj2JR/bCLoGdzNXGKVwKv7bSR7ljDLc5M
I6mpDjpDPdDh/mEJnTvtGyaKc+DQJnkFCY90Qq5vCtC1sIOV3jW0DEC1GdY/et1Dth7AvuadE7QU
kvdpDJgp8nwId7JKJxgXGgrrUKQ2pUL+b2ctr06eC1q1fZLLaOhELkUI+/xZSWLonDxWtR+V3D9G
pGFvd6S+AyCxWhshaf8pdYfcdwKn4sxHzYWmSFKDPDu8WFFIsM92O+9kHGtiGBJFCVkryVfxrgTE
ZrHMThHE1fZSoisDr5Ypfbs/YJqa8fo/D1R3jpYUj0FRdzLZOk/oXprxhnYhzQkGrc3EGCdnSTsy
Tlzpf5tmcJ4cBdcO5chVUGDXEtffddONiPq0tyh8sXWamMrZwejJZkQFgLTOBi1FfX/+y0po8JUf
aPrgXTaX9ObO3xlsZYSiMr9L9e5qi18/HLG5YF5Ti5TCQGUUXAP+hWAUF/B4rdDQ6hvMN8hz7n2j
DP4WqPykGiB4ke2ajhi5TvOwYYaskAZKknFP1wE6L+FASUH8obppGVgcvt6QUQUoOgH87IH95hmV
0WuZ2shERFlS17U2HZLgY69E91OHWPiWbvP6O54VU/j6WmJJFlpAyNSOcqVR1nH0gTfGjBZkkLvz
8LG7PkdLwTr6SVz4fbdZ5pEUEJWN2yOpJtaFeLPdRjNTPC3mgyvJgkhE1MYAKxOjNbgUwiwAYWmv
ep8oWk+882LAVsvE9gW9wrf6sMQCY5O0I1VV7S5cgxIFRI8xkrPTEE/4SNSmq9x59QtZ74Yao8h7
SDKNTJtzBJnFQ2xYM1WhzZmdHgv7r98r79UcihNXsZf+gaLZj2cQ+RkQn4xZS20fLz1oMjj7kOwS
Hia7oNoTDFvWmg2RjJOS3busF5+1w/wHGqOnOwHIt7OgrpchDj0va9FvCJre/PJuzQqW4kUKcgGH
npOsGHb2W61YwBUn1+oPOazdrLMfedX0ldG38yYP3/AGDa63RJ9npbNQvYHQyUD347a8t48ejUtb
SOzi4xPOUNLZNkE3gQS2L+2B3qlqhf5tMrzP4cfvSh/MadQGmzNxG4AS8pZ+CgwNAcd/sBTzopUI
PWr/GI0Ybsj0lC7QLK4d6QaSzk0JR/Kc0z7kasAltwiV9r0R2A+MsQwOjY4fIdERo0cptHScUukO
HLn5pb2a8simV88DjjZ9g/SarRyDFIu958MCEHB3k+Xxcg4XQBDsjoMRaMyiIQEjNgQDfBmd1U/w
3OB6ZVnSYkxWSF56kkteAPwsulO+uWMqlPrjyZprQL+3/trgityvQu9gvnAd5+KaTfFLFZa4uil0
IlE1NX1st3DP6S9qM4iTt2KaMEj7NTv5T1f3WjYhvjwPo0J/WnpmM6OeC1jMLydohRfn2MJOqqVj
HuxFLPc8T1WufpznyzqxxnA7XkdsMYeUr/jSZnWD8IEAAWEg4dICQumsxvyf8z69w3pxDx6m0jcu
Mx8P3b0+9T80/Rcpvty0RqWSW1q2lbaWEMf0tpsU3CMfqTAG9uUUXt0MZCTS1aIGxAdRLVfX3tJM
S/f+ZEciP9+AZRY+uWYGzxHzyTrs/huBiRleLWdT8zUxoAvDYO9Xk+Hque6bMPWcCjDI1TVH5k8T
62/NkC33ptq1XfjHeqfRRCuAvx3E7ildSyj+D0YantSPU3NtFhcslchm50DUL+gnqzKPa0BJDCTJ
X2LyY/sHJQQfK6fr5KFibRE4T+4l53IaBDpEz9MC9mj7+TtrjljtGrVCGUAK8Z4tqLAYEl7J896q
Jba1cxoJZpk3PFX1/34mt5XJ+BOMtLVHP4wGbcKyDEe1z9v9howTGUr+SwPhPdSMCkNpBe+wiQmG
7845jqh6WOs+kqBKHH2DwkR+BbYVBw0I1uHE6uDmaaSUDyTlgvOtm5nft/5/xoJkPuKNWREqg1B+
l7Jz6/VI0gKGQB/mwB1obcPJDf4ZgZa1DFpX08ZKFiuH1Z7foIldEQzamf6ws+vQWMfet6F9WWFS
ny+1qqZwuiLwTYq1afL4kfV6DsY5dOo+U80obi0BTsMSpy4hvJWLXAaHkk7o5JZZFhnYJhtZe1ri
BXCxhOqL/LebIlyWmc1Qy1dOmnBx5XeWYOpkAGPWV903qmNnt6VcB5lyMJp6ap5UElvptBVxm02e
swtEgoeNxUjtwmd1LXeaUyTb2/jdNDnb1oD1+rc3PAzw5RMg9EMo6hKcD3ihI7R0gOj4R5uhpOYt
xk9eDSYtHShfbEAXNCJ3l5a7aeat5RdDOXNp8FsQye3Br6fmxzoXyCmUXRppUExiVDz05c2//rbU
KfJMDJnjpz9mCfqhWa5c51We8UXkc1yF6OshxxrqP5jczElzjmvqxfoT1W7QGUM2Y7MPm2ilx2a8
05YwKGfc1O14lGIfKWlwFnq3GLuAnqZludMdFaDoTGShFWECor8QnRYZY7WOfZEQ+qiCVg9y57Lc
IZyRShWyi/9jKGjI2whrFkwpQwz3ekKsQpJAIPlZkwxGvtWsn1ARhqIpFabyf5PUCP+ZyHok/MKa
6E9suVGDJ/Vf65HlAeA/3eJx78B1Zls47fObjiz6gEgGIqrN8ej6vKkS8wUHW+Ry6bRP5i/Y5Ran
5L6ScRfdYH8RYlviwgGqPK6oArLYczuN+u/XXbuzdwJkbGCGBblfwJm9cc+mIF4AtWyJL5gz/HLo
b+ic2LX9hnovvPtBw95mFyA7BqV7g8wzCvP/Klfqr6far2wsZn2bGeNwx9PgkEzlw5KG6CuHf2wL
DJNmX30+ZwfMeEoTwixSJ5xU1UPuaR4HrVcxN9ZRAXk91Kxc1m6V/iON7F1QUd82DeYe6q6jXCRT
dDHiRYzijBqsMxL9rj6T8Eq3o707KTjEe9yC2jVkDKiQ/VeXIAao7JTAlCAbC3gQW6pCa9jTvGpO
Lu+W6nzCTxnei1w31TGS6qZUMJhb2otGdpionV9W0Y2XPM22eEIDBbu8heydkAb87fIM2g67UvKG
Y4cS8cBCJ65CLg9JDvIgvqYMKJamfX3jis5cIoxznTUstUkbVlokLQcwBCaJU7M6vntVan4Vvz/J
Ezbfk2Y12j+woy7ZUSZZn8/n/Ldq96IFVSzBlqehAcV0qhO/mwhe2iat8O0PcGtIy4DdpPcbNuN2
rfk3EY+4neaatzQ5qxlsykiRIRRmpJY92J4Kdo9vdU/Vd6P4jMPfATb2QpchfAMGOELW+z7oWkAq
aHujdMC7WBsu/ytajo3efLtXSbcgVKbJm+/69u4bYBnSyCxY+leEXxyeTSZjrDdPl4tTcO9aT0aO
vq/TgNd/Wc16lGH86tJ2f6m3m2o9e4UsXZLdC6Tp19zgpZju7/JE4mzoureeCq/5yQ6FbymPznR0
cgc7UpDmXiwSZo0tmUXgHqb6tVyfoAYbHh9J5ouB+mDuBtBbbgGxYeMKm1/TXuAjSSvBPqB+M9AS
9wsVkPZYpDfphEEiwcAx+Bv1R+xGZyx0NVdl5wX5mqm0qly5qVYWZ2MkNm8l1Uyfmz78Ke6PkqNB
d9MUa7+dnXGpCyk+ujGROq1/G58jBs33bjndCjPhSyBDl9nrgFo9CkCT9VWqjIozVsfPLSo7oCTl
OV2v4VM+WD5iVn2e8p6jJ8QB5CWlCWFZ8N9LBy5tfy+SJEOgMpaAtAbXr1Gc/5s3IhTBgSeO2ka0
xYXivlnE3DC4aK/4YDA8iEZAC+PbQDFt1GUdCKaJ0uXz/GRIMvtRtuOv/nV0oFGq++LcAC/AmHh3
g9ANMt6yVeDlLUc0laVEJigesF3otZma9qxCttasLWvQ0qlkjxf+3ElCm3Mg/2ri3/hFKWlfBipb
Jk0CpNAc30mVCrzMB4ezzmDZ4G1EY1RPThdeqltT+oZuBrhJKXiFVpYB9YcLXTvpo0y1p/rF3P5e
EeqTe21TCnlpw9VgL8aLryN3rHs+b8ZOYXHWtQ8Mp8/8JhJA/3z2lX/1R+0fcy/LNYkxFpEOJ4e7
TmlYsQk36iJaZAPhJMCMvQXzT3m4p1zGBK8IXIngDsrRmWJdu/bTKy5A2jDZ0H0Nj+Sr0VZP0nBJ
8qlv0ViPRBdwqJEkBI4fiq2B6/6HgVMpBYEa0W+hyNu9CWFPM2QOyVhfr5r5YJ+P02KmZHQSATIS
NrvWEqO6/EWVU+nvnpueXHds1nKFaWa5YcXHs5VwJEkT6nN99iyhXyJ7bCHn+eBEcn5BZMaCLapM
o1xkghuvoAuS9HDO5eLtzM2AYu3xPhr+L+u5YbR082RMGJTRjNAMwuNQwzONCQVbiJ5qjCowo8Qg
XWEYlQpmuxpcY7Et5jMIInt2IFQfMwzUSkvs+UvsMrKR9lcm4LhyP1reey0FIDP0juMdVn6SfASX
Kh3Is0cdoEtlHK86BQrPWlXgaAb/V8cHz+2/DnCZEDtTs2/SeJCM31ez7AbJO9emEXtUP1FlXQMU
v3s03kjn0/kSaN627Qf+Ms4qXyG1ZVCb6l/utgedyaeBZOi5u/yJW8fIjbTH4HzM3fZaF5F/ta1q
GhyLMTKkOkCIJGDyAVPv90150pghYiwkGu2sYffuAyEztMW/R4u+GuKgN7rbVa7oxPfYCS9b/bhS
Sgq7l/zMFDNa+unr71A7+BvGIrfayMPzUakjNoJpNnEpugq6IUT8w8qgVNSK0aTO8aTsMcohuEer
y5KaaZm/ETZ2zQn9k2rXJMxra06EGJgOopVRPvJi6sEFOW534Hs+DNXkZAllXtA4y6HJ3jiR6/JX
fxtnoW/M5392+AtgFS1Sgn7f7Ey0eE1S/VwBSnGp4WJvfGn9LFiNAnsfg3M36DSmWuoc8KRUfMvY
6LuJ+PGp5YUuf5uep0ekXLc0+RbV3CgcvVs9+9/4DashMcuBovuLm5B4EPNMWF4zQfNm69Vayz8j
hm20P0EGlcB+qkhXrJa7TUOk84vc701uxn/gf/ABHv1KpC3NJcjSAsnf6b5FxZmmaGGp9YdEcGfz
QCwPStqk7FGqz3q9inctn4SNINN6LnfZlHSIWF1dS0EY44iLMQHBCCbjWzRzBhchEYgVjxJNLXzV
nfzOASNJpsJ5KdNb4gQzzyH4GFuBm3ShoqOorzVUlfgzgK6jejhSHimdnCHjzUsmDnULNaPtb5Lx
kESwT/QTByHQrMT0aS3Sw81qn35xympL2Tj78bEDRQi+SY530VXFxn1agvHFgeAm19PWZwESssHx
+y2nPbnc5Ov/kLWET1hG9icxxAd+wFtv/LdOb9L6QxLntRq5aIS0YEfdJVObnQ+1SXBEMDFVV/Os
4L/b5Nal4f50HJHQ/0IdswokjH5OHOgYwNfY41rqy6QmDS8T3wTkv9M6MOhKFuupyE7DSbjEeEsw
OCqOhQVzdwCxoE73DeEHvtIiUp6PTZssBVqJ1U0SMcNxRaY5OZH3KZlNU4zV6CVLpjtbovIWtQk+
Ugm69w6pjL5q/BznBiRGSRV266xEYiUO42TBlUpBWnWg5cM7s29gVN5DQ/8Sd+WgM722NFh8M0L9
+yTGHzwcF7qpRdaxppFdLyo9Bm0hm074CmEpRV3hKB4m9Fa0iLWSG0DSuSclEnd41Dci3YdUlW/9
VQPY2oYLy8PraXVdsrTlNSJqWkctMpjyAoxog6Xq3CfvWvEP0G9rtcWz3X7QOcYt9sMSIhJnezU1
0glU7xISMihPCgi4hWZUQV+H10+zBDUSdv37dSyQgb4BYHfehKjoTUzMBb40F4fcugBH5Y4NptTA
Eq8nO6keI6LVWVHA6AQuG7eiDSQk69snwp8BGwAAI9pwdwhmJMrW2x/41Z9p4PZQi4h/w8wm9BPv
ov2skRNkY1Cw0Um2IDqOuqBiWfBi/7IFxQJYhSIahJQ/mMam4ijbUafYQTcUFl4gZAI0uCPuWptt
FtYKlmtEzY4o2JYjamyBQBhvyCiArr/gpgOMCNcN/eApyk7xyOWYsVmwps26jgfegXpAjUbMbIfB
QXRGpOzk3pyU0LZG1fYR1waz1i4Vol38xdgK1SKwsOsw47F8jzZYiJkXIDq1rltdKSnA82ttmGhH
FYrO31gCDDMoRWxLOJ5n08OtOh9wSany5zBSkjZWE0wp2ZRoxNkotqD5i48nl90L+sbrYTy63oDW
3iDSZSt2ly9DVPw1qRSo2ySjpH+0hwbEqOk77yIzJN/Yif8r7HhXXF1j8+hzq0SDoA9Q3mYDGuHl
L/2eqytyh1QuXuAmSa2d8jt23bEW7EGE/d7HM6X2V0MAa3itgI696H/660q4fTL6YMQUUdAGSnLz
JZF/pbeEywkAepP/AxkJ6CTl48xV29wZ9vbeNF7GZBK01PzvKgmnUgQY9BB3jlob08rx2BNNS5WK
I8Om1TJoARm3SFtglsCuPNmWzgSTfo7bLRYJjwYixPMADonG/TmJxHhiQHp8gkeJjin8Ld8t7a4x
t0V9U+DdnZjgbJalzD70O/YU+k2Hu7OFobWgdfcg7ZQQnrsCOGAAX+R6JbWYYg8JeaqbtB1ELGGt
qHZlnr/dw/VIvmV2Fzx6YV5SqHf5jvxHKJAHaOSC0JGS3am4IJkld3PL7QP5LD0sEAyPhGjKIMCT
MKAt8EQjrYC4Mlnoup1NBbCB0NrF6nsSN0vdbi0B+Fuq3a94Mqrzc5styxBRAKb5D6S1xxno05Ln
bJ26Jj9RDFJ1ZqAwosEH1Wh+zrDVQ9wmEzEjQcwd1s0ys0BpZG1c7WHGh948yvwuXmWORzoRsoEW
Tk9T5+srW8IQnTMQBNqGWjU+D8hhlgDdzsPQ4Uz4sJprIg+d0dXwmKOgPEi77ZKbQr6YIINd64Sy
SG5Is9gpDzJddijso01ILgd6JttA+TqiNXxuYn4NgcMlycVdLG+JMdHnlkc+HS+QUYCsdqiCjH+L
sDQaZgRw5kmPTljPkK7+dJOvBDG8OxEpqJh7toSF6npRIxAg0hl3ZulvNE6v3s3DIHBvC9XnTTuE
m0j1ee1BPrPrL9IImnAJ6LOs8aVRXyu7tZ3lr2MQ/OBDcBfeN4CwitnIG3KxgR4B8E4X1EK/nlpZ
lUB31FJJ4HCGj0VSJkaFLu8LY3AoDpoHzuMx8+lBkBkHSZsDqENrJa10OqlfMH7k36gaNqa1sJ0b
1v9hAV89XZXSA2874TOs5wAC3e4SEziwfHYFsCZgyMyz1mR1+UsrUVC+Xmh705xWwYg8DrTv2pYM
NJ/xI/oTuTDbimw1vfi2iQ0ahWd06e0tdAjYlL/kJVme29E8FgKHKASXyFzwHWYJdBXfNEz+Ugn0
TFllfKySXWO0KopPdmmnWYhtwTymaiQ6qemv9C6M6ppvKGyiUm/Rj3Zmx3lzz6SsA8fDsJy+tWx7
hAeipf1dkZknd37ecHW3D2kP/aPZqRNwSRZSaFhUtqb+wwZYtoa5Zb8AzwEkmQtFmfsAX1DiaIoQ
DzMfprxlZUh8V+OyoioQ9FK+92SmvqNZoxiLqmadAeqSsHfmif4rGyw4nkAdbeh9SD7AriE8yOF5
ejFG309PYbapUEGC1uP1KKqxwRLfWinYlGJU95kKdxfRyvYnVdIUW4vWt2mR4bEnS2RqCVQ4jDAE
CK6YrGNu5dFkLcx09j135JrfXd0oyVOqzMlk0PLb6t7QdHvRzPFhA0Kyn/8iaWr/i6+H0JPRWOhd
q1mQQBkjhMs2O5NVsSDE5lyW0jYUQHlTmsZWwJfz8JLrlQhKbvVqYbCBE9CwtMMZGlbn25a+T2T3
tqvFVgaCif90Dy5Qd6zzpAqqK/dNY9ykg6RIatwTZ8iaqQhzqCNnr8NmSNRqEDo7rS4nBQZxkpaK
3dITC77uos1XnnbPmsMu3NHOBC+k3oOnx5IxyRw+acrj0uaxNi2YMPYsdq4meNJP81AE2FvRKmbV
nP0rA2jzQ/J939N3mrimykaHZrDq7VAGD98LJg2LE7/FOw38M6j5mXb67LQw0mEFr9bFvoa8bn2R
692qlfZFSVR9tvUGqIMVrvkq/GUPvawcGY5DP552VTk7S9mbAKndIKGOJTTJSlAXya0gyAFgIj3L
jaUi/9RHBq5koaHtVJ0pGykOayut37StK1FDBG8FtpxRtJdeOyB4Q3i4t2ZFSyeIwV/qLjwHCuxp
H4GZs2ONPj0zX/91IPs/mJZFJdMhbmG2Md0Ve57tXHd3x9vcGWt+Xw3WdXasSvoEzZtC6StIk/RA
iSaFCxrAZnAQngienyitQiYUPkjWgcs5801FQYzCmFrx2CtVOEmxuu1hcZWmWwQvFhh/HqJd3duF
BDFJ1HAZA2wq5DyFC6t7lEfSuomLkIvifB2ccchf8DhzLkId3ByfI7EPF33No8hYFOkiL2+IiM6D
rcBd2qSRPwmzCXWrMPJKqaFB6STYtI3tfnwG9Vr0xf+uuzDP4qAGsDAgmPy5zOIrfZhxXQr2g93H
cEfNoIe2xKYwCIT3WtTGkCh0iq6Bpzy+PqI/62CJnNqdfbSXrtzuzY3YpeTgr4ndc11+T/99Lexf
qJzRtB7qp1UqHRTnDE5+DRRoA2QYNtf66R0wIU1OLry8m1pOWFHHRUms9P8BzHQsde7ERkzZg/BQ
qzYoPDIetAdkh5emMjX8tHi5a265vQdE3Q5ys/EAKw0cSAhpbk1sNqPfim1tOGUk/dF/6TaaLuXn
v2UuASBvUX9MJttQQjH9I6y7c6SA+1aQfuhUDHHKw8JvgHbBRn6KRqYO/Se3riq2SsrJ0y+W/zP2
kbiGO1dKwQ2gp28WKPcuwx0NsbJj/3x1XsivvzBjbovCvhxT6bbDUshSq2tTZxRzsZ4lCOUF15Sg
B47FmmKE9F1GmnjYW0wkhY+j7zCndSVSTQCmx9xUHe2W8or9lA2wrV64FC2LWPSP23ZDutCjWSW7
TjhyZ2RapP08dE+lrqbLQAoyJhF3gZ9/7wn68YBIG9vvoXW821uskpyUoiXsDjHR67L95EwgX4OK
gUGRRWN12Qy3hoHQ/yoAlMgmQ1RRswaEOpJ8JB4wihjeOxwXoN/TpWi5LLJknbQ9xEB7Rnc6UJfm
JSHzNGhQLPb9OhdPOm2EGxMMYNtvkOfsaqtfdowOaUsvQXKnsT1GRb5ISCKLLgAsGL999dSSWG5E
Sv2p5HPlX1N5f7lOJPUK0SWHbstwGtWlMIJw8iIwnZoUQxgPVVfAGNOePp9+5RscFszCYGgJI32r
yZGxzYZQwN6EFRiIEXw2vWofStuKQoQcA1ykxU0qQAGWU68g4DeE6ktl/DRGTGig21dp0xgwgyVG
pCDVV9YD+NbZDRawmIL1QQq9BVeTraCmBEdS+aO7DLfnmVN1c4k5o6/CntoAIta36SLmsqtywC9i
g3zthqTjIlMHXiP2uh5NReIwWmeZ/sM/HahwM17AP9QrZnFpOe5REBC+r+3DlQ3iWXY+9QTGJNPZ
c1v358+FO49mknz0VxPAG3ZsZsD5UXgpcIzDg5D68euR4j7gQ/WikIVIPSqkZv1VisrZsaAQGpBn
P0Vx2ZdklKywHtdtchoL1pJhorHBy5MYO5Pk6J/CFFwhTUFVoGu00xqYkf/fJVlC7sAqL8bvAakK
sR0wHYO17UdvfGzeG+SOUSJ/ULeeXi6MO2y4v2E5vnZwCem1VO4smOgtPVLo1V8RuCdve1s6ubaj
noS21Rf1TwBEzWzMmGz61T3Xm37g/yZH2QESCtknHScfsd/wlqzDvB9eZhATIMJYorQKCIkdnO/d
oa3P4y1DE8r2yiCIiZDR4yJnrMm/OL0LF8LZ26fVRSYo3efBMCOxkq/Lmz8JdAk1aeVsSxTh2plL
m+cDn63Z6I7WSM7yKFwni1yjPCXTHRjSZp4q8IUG6CxckpI/dBhWooemOBsnwrKPxSn/hJ7e0xjI
y4EMZsi4PaluMjVP4zPOS536hQCnVex371usJ/AhLDbK1NgUpYxU0NVcYVm62zRykRqA0x3srhgY
eBcwMdXu+DXdl5DzrGcQHSjf3LF5vrFxmEAg4vDGEg1qXgPlTwxFrgjrSxnZuEdewj9bHQjkel6k
FqXtayT16xDpC/T/66Z3mvvptnjlmmq+4dhEdYLLfjG+WmQyFc9e6k6CQAjQiPXZ0PV1D9qBhAcn
N4E1d3SBhABmmJ5GjuvCsAr3TecirM4r1W65omXqIbfMiCes+Yan7e/2i1nN5zF67sOMzu+0b5A2
U+CKPKaZlR28SX9TT7Pf6+aa4vLjWeip9CLV64Q3TEzuIzQRPFWcsuZ/Ostbq5WZslzESoSNLF0e
HIqG+dBbHU6C6IIdgj4fWyw1nQvLYceEDzaVAtkaQJ5vjVK3geDtBF4gU+Vvu+qW/0Ww+7P4DSWn
Ir0L8b7FGF+oLvsV9wrSmKKjyJtbLACfJ/Dfu/wqyUasou9w6T0OHLRYWIWdlKWVS/FzE3JeyG5X
W7pmg8fM3xE8AmZ04tZWbz4DVslZ8MFioLj+dwIrmbr0PaTjDfnjTm64DgpNulg1lGR3RsrcP+fb
06DKVpHsPeRU/xmljH9/LOHLI8iCm1Lm89uurDO/utxywYPXWVrBWCK0kZNyD+oo2njwer1dTBBw
Sr7YXWVSGAQH+w/QFvDx3wr98a+LqTwRhFQyKH2jHf8sxP42CNzbaPyANfjkakKk5oBSNwfI+9Bt
ujKyDQFNQ19EQIyyykA4/A3AC6caqlAxVqCr91a7yjuEZYwvRzhzhHN9pCMnr5T0pJM7Tiv1cXcv
rNV7FQ7MPg440FFL1I8vpmeXzuirWvP+EG/HjCrfuimKVjzyaOHBjKWCb0bpmxmpgLbuyYjv+fWz
v8CPg9mQTXLfh8izPNLCGvaf8e2OPHrfce3aUk/Xu4d7+Yy2NG0X4lkMQe/MDVqzBOzzbW+MrWqs
A63jeI1Z0+vLo7EGImf8k0j1VmDGpyu7827ulax9wxSW8UYGW6e9c62hcrQohYWoKvAURjygbfa3
IxJW28Uhe/OGkAIAvGAf92t87dD/9UQuPAkfDQFT1EuXoGp29zZ6fI9DA/+XQzwfiufvSLBi52kX
lLcwq+3Pq9hnzHNk1ZdihEnU4PnPBLYOcTux+7BH6KajzLyUjU8CoBJloCCsmJFU2rHr1htELzS8
y1IKpZ361fOX+jcOadqQtzweYlxlsjarZk77JZBHLdY+xS1oMQAR4XUOOYoh0ZzrN3ZctMzTagME
skYyiel8JYcPTQFlQ49GToL6oU8lfLmHGF78J7uQCPz9haIk16qT1hQUB4u1Tn9qUQOSey6BMMlD
L4yBmammTe6kHdVA4rL9OJO6BvncSdW1FFZQ94DCAmtx0WHnTrwCM9x9+eYzrrtXx5cZoyvgbmQJ
o+eJzqyHuaFpwzMKBDpyDm0t8wXm7M+ZFOfODDpRxTxMQCcnaRu3uqb0/ayjgStldNVDHQqAIEQ+
7UlyLNBRjgjAABMvVR6IJ2xXHbm3L23LIu9d08eGIBSNsBzJ/tK5bwB2qqAMvh0/Pmc7my31q5zE
tRV7hl9Hml2P2VqcYNr0Cp6+QPLGhxoLwVDMeSAazuiDfDxceTaPnpMbl2CqUY2/ubKb+BGYIIhI
2NLzERTlUpGqAqyNXwySTTwztYbnSUXPEfJyB3KJOPQTW1niUWdUjcgGWq9is2M12Zymq+igV/l7
sv6ad3JASnS+3cvA0euKzB2fkv5JE1Js1OOPvH4dHWXDp3nsyOZe8cHU4OcAE0DJ6l+sdrswYqeY
nYPoQUgIu8wJNselRfHsnCzbF+ZSEjHOsRsQlPo4RCQd3DC+AumRNCMCRixFlY7ha/UtzuoJ5uHs
pl3FhyRBD3S3A7b2fY4n8Tizr1MXWLcOL1sGDEQsxLq9Lfo0NT6o9HX/1+66B9MPdvTZ+OUyXe3u
ZqhMF1B23ONDfp8zx15fmuuviti+Ocfq25dy2CgJkmSTFKjhInkUF8GlvzClzBgyckkB1STrzcXj
BngywWAaiTLxRNYVd8urZHqwhn5CODIgIk+as1V3SEAtDUOmxph3esrdha/tyUQZZIr/Q1Lv60yL
x+lvSU1+I2OWpg8zfDBwnGRRH/K3mQzhF5wCLtJudXeMzkTWVrAbEUNtVD8HvzsSEdBSbIjmEDnm
5wpwJhdk3SDp3v/dgTZPAQM6WBTe9dw+JAD2sVLoflhgYrJdsfL/wivGawU4kTZfhx/1x6xa9YSK
hQk1I1DE00yNwITWrrfJxgWalJdQV2P4nsExAP6RkTka/ly9mrN9Xqq9TV9TZSWBBHn3RmkljuEi
Vq5emKmNGp/v0Kn/jqxmsOOEuLVbG4DAILBCJbZxnStCuFfBOBWKfx9Ea6lxUVMtfz6juvQZA+Ox
U1deVj4lc+gND+j+evPmvR8j7HicDwobyUdypBtMK00udy3VWrwN+y1ksOBCiwD3BT7gjgxZXlfR
dgxc/qXkYrapqR1n/GsGLywvbNtGuR6pycMuPsWgxayh0qfRvaHQVVQfyurxLvTewNfQgLIUsIYQ
eUK7e1OiEfSk86yNwxPojeCNMookYivT9aMQcefdM4pYxmTqrI+uJ09thL9+CM/O7XU/2pZ893oF
O5RO9o1DF285S+FosUmDGj4djUNd33gPZUahzPT/hPqfHEIzenfFBxaUdxrz01+xDCyuP5wiJiqR
ZqD9BTKSgxPyh93JfpVLG3g4Kz/aa9Lgv+1+p2DjzRoMI3ShL3WSkubNRkuFIAl4pFu8ZOP9UU5X
lvzTD6jSQr50qWJKrX308hQVitEEGDO48D/GLcMIa6UHGUTOjCMasiPni8qewL7ApTlIVG+9aV/D
yrpUYqRQzrfLlUxxu7EEgTa3n6kpg49kTeHmHkFFctBWwkhj3nn1MDgXGQYd2e2l/tUmgi/+LgQa
Di0E1QAhj9OiA81+HLOR9MrrS+t5LAAV84ruhYPjW4FDtBPe4wCXf3B61jhJkvoUsEy83lIZWciu
k2GHo+PJogSOeBa/CIyrRd5cY4Bb+vCkI8RR2Yz90hQhRUeYFs7fGrEzg9eAZ17ECrLndWIw+KLY
clLGUyEH2KZWweyKnqAo2+sdWZdXZgw6jKul/lJBaSbHx8P5htpNgOHaNNQio5OclZtewap9pjn2
V1eG8VMj3Ch4H4Ce5TtFZpORai1sOorEPe2iK8RBEbMezPu6+4cvYsqKBfLK/na8g0kk8D6LUiNr
tWZGOWyhODBmOCS6cTiwMdmW7Z8orbU01OsQ07OB0i+en9PoRLBlcc/NAPZWgUy52MvIS/L0pNXR
i5iNr7tf9wXK4Bz1RDtmFUyGp8EVhvDuheNdqXHuhRrai2sz1hNHtqrnqfZ7ipYqGZzPtb7hoFIJ
LQb/GRgS/P5TuXablSvAKOZz87P7gTopGLRc9d2f/fuKfxGK7KRYxyhWnXG1+nF0CmUMHbYw2LmM
nU9ggtooIGFG49Ai521tPL4pwNdPmV/vqeGPenmUK8vNQD/4peTu9/aS9Z3nhvM0ih7DNWW6lsVo
iARbNqk2Xu2iWWHPwWn7D2s2VaHXf0NAmHS4KxjRz/ElPQBJcGHhKPzy707m9A+3RuliXVBwQ0Dp
HOEjh5uJ02xbcKn9ps4WDIrv6ZB5tkc0Hl7lfXCRxw2hcJ0/bmfIgBEqQLrRW2JD9o2JugwmhwE3
NU6RSc4tVvQf+vuu/8JsQbJv8IHglQR1xy1bfoRvaRXeikhC3lkMBCVHwjmRYJTYLAp77lfS1PIT
LqRUYGKB7GJMxSELx2KEtAcftCnQFtrmUJN1M17247y96XcKLTlWZg9eYXfhWcX65hdC1VHrCH6j
xnLcAvvI2lwxuL+3Lr5v67Ov3HqlBVAk66fa4ydg/3+MCNEnUeOwlsVm6ZujsToDEhmas2ms9jjh
pypZnni2kJKkvuu4nKzTlRJ4I6QLk2RZIT1yqdwdawuYfHslPQ/xarSUWk3LSXyYkgfXzG9Thxfh
nXK9t8AoHcYEQvQVHjPHCdvEauo6uIAooLqD1Pbsb/Pzrz7WqQvOoUEdGq16TQ9v29jFeyTrqr6l
JipEBES6auBNVeqJaX+Q56twzlC9gE4LIaAM1HNG4NVT3f7oYLtyo+YLKwwEu3oGkEOqCEk1oZ2J
V7jk60qrBRInCjk9OJ63uwUoBGjt1ri1R7xA2QmQpPzJo0XSggM/hI3+DWcx2wX7juIeCsNwkaOf
+qLMuHCJCa5kNZG+hWkT/1i4kHU4C4RCVzJH5BPSl5kJy1hxhMWEZmGRRf+3chBN4JoPGX1X++ER
RByGO0ITmCzIwSSYIP3QNJ8vie5uzyxM7cZH5tkRc+/RmRfuvh/gjHhL3LgQAgM0vGMAlvfE1Ykw
vNE6huDG0hEnyIHGc0oSIukiHE4J1Wi0GmPO/49Ln0hZAdQ7f4XQCTZ53jeKTbbfUAwfwq983v9l
7o6E3eAJ9xQLIyXcoMF+V7bxM3Sl2YfzdTNSBwFBvOqXY+UhClLQ2BEyDqeyv4g3uM/U4uBZ9Atu
rLfPbvn6PB1ezLCVvmBjv1jLrBU66xwP9l0qLBNiHuAAK566FZ39jDIGYG75oRjU+1P/nXOcEfyA
/DWIhy9/e7mUrX9cobTapc/wVJwRRe6CS3SvAsc4brOri/x3n8mzB/pz+/2JexObWWD43JwcPBhQ
qc0wM5TeI6NSxVrzRatCEFuncp8+f/9E5jsWjTQv1FR7IY1AQZZ328IZAO62e00YIzfqocDgfiNC
4TP9jaSeL2ivUcdbHCEXf5oNONCy/IUpouNoTWe+Z+mjyO+342KMk0rxwkEN61E9lrgz19/uTdiP
PmQTw1Qt3x/l8XwObn7eKcvHhFuWLEq2YzRf5soR/u3ggbaHxUnHYiwiHD89k3bqAvhviniolM+J
DZV2UUFqkJnBlnfxqOMD0LGpSZZEfdjvBmglpL8jfdQQg2LLUOgg4955gg96duowFyuHTlQXi09H
6mXNCBxr12xAelNepxMepoic9GudWwAlKmq5DVSqug9VqqnawbtsHEScVaMxC4CuD5c2h+Yrso3I
+dq2J9I2y8Hk6SL4eHzUn32OU7/paO4UQykwCoiaEUaSyFT4IEp59GaYw7awbB0uAhn54qNbrXA9
ntCWboeM3cPualjtOyXGpo6iRYr62CGi4nqfaIB0PfNKu1fAS172w5UVNDNVnBzNlbqk8BjodkHr
n1fA1RoRrjLV7tQ5Bd04e3EEAdd2deWQBiERAfzFcHlVt2oV4RgGdKZb4Qm43k8cwNDQU6IhGsP6
D+CRMvKr2LyWWWC1xswmbHDsPKZEb3uN8ym6ElmnK10f2z3tQyA2ol0cy7JiM+41olThQiyKUc2y
+Rih6rNZOrDZYgDQrXWvSTyME037af1xytaS6bQiJIu8JhqbJfu8lUvyLfWDq0JFvVvp16Y3qsFh
BROmg8f7Ez17k7DI2y2jZ/u3mXtrjKk8jC+jntOaj9aHnTggcQ4vt1mpkZQzKYVEFDD+Xk2T9kFF
6RWvkHZLL/0TBd6GQLjJzUvPg47CpjF4xAPvTPeT1+oKamnpKhtmebx0XLdkBW7DFy8VOJznKmEk
KvUy+eINqdOLsZ6RgDIVY5iZJB0XAwBqaX03kfYbveUhGrpxRcPlUUn8eRX8S+ZPYW71ddZF2/Az
Vpdm+HrGFbQ+3915kdlDS4aOyNMubOpjc69pMNbNUfAcxoavbdHRK+MlnYoFo4eF7UBFnj5INaS1
CTgEQHTg439/NmoPLyQL/1vjHbExGWqE7IBV9uJxn+7rBqy+5hSjrFG/nwhVUnRBBCtbUEodcoX8
8jN0Nx3Vmbpq3tT2rNr7vnAK8/jC0FgJE/E5Zzz1jLP7H+ygkiEKSG+ae/hmyNpJ+QZCAZFzTFo1
LluGJVMhp/dQ7Qncsp27ixG8te2H8Y/m1YE9jb9YmQHwW7G6uAIBFwpuAoxuWK5Co7uaKsgYgF54
jnDjqseh68kGLcTB5EY/htl+DSR8jCGj/k2mDc9gR6zxnSaVKo6RcJXbmz+r4zTDSs1SoZaSxJl5
FNIxpuPh/+HW8qHYV1135lTXl/xVxoEo10pPrVcqMYssV+R0W0EDboDIYOO7YHNf8rc/BJWF6m45
HYcshsZkFzMepdqxLY7VhI1LELWbfZnTJqPyIj3NmvGy5FUFPklzGG2vODUqIBFyxqTqs6T+hhc/
PAvR8nVZRR5iP4dDDCWdJslsFJ0uc7sztjzN1AgaWXolg2HjHdCgNEwqs9jHMwxTe9GBjTRXg/BM
Dp4CJUfFzYc+4eyHoFXD5k+SgMAJim56Ko509AuGQ2tf4R9994MFUQLeh1IRPA/667BKUelqNKS3
9NePZKgG3imCuqzWosIfnoh/fvoLRJDXUklEYCbxs9jow7VyCa9ykf0LliTA0IO1E3H2ajq7oGN1
nbaL/e+ehQVCaR8wsviqXX1wbuMKyzRSOAQMt1NxqKPXgF8ZT8N8jWAhVdXMQyUzURX/hFo2CJjH
TT4IVt1oVnMngfusRzFklvV23ZNVI6SOz4mD/qssomRAQZCfL+OwHn9A9lgOg/nqjB9HnoBqgAJX
Hd674NgKEmVA/C6QMEe+Iru0X+X/IvJ5RPN4kC0g7jFT4HpwhLX5XmbzMcU2BhX5GPYRjibiLtx4
NRwXNJKN1Hy+rcj6emXUmYyHR+S5uhYZoU9jB1HIgtiRmqT5TZXxOmLCYs4G8CnUyWfixis3jkF6
ksWd6bt4Y9sARbMfPziZ9sJ7YgcZoGo9er2IYze/Ac+LU9dRCJF5dk0O682q5uwyxPBthbpDcl5y
SXJL6ZeVNyULC6TW2zPDfbk5MyUoXoce4oJrQaVgbVVtsietSfM0xenwSJOxIioUUm28Gr2UOJM7
iM2MjY8rtnjLOSkqo8T1okzmrv5cE5G6NJ6r6Uxv6aOgEqISLIBC4v9KBihNpDoQm+sQcZnUu54J
3jISG/USUjjXzWT9WPms8nCNM/v+CIK5exeJrLxoMycd+/onTSfVNZna8eeYvBhHWjmNqQ7JayxH
KmsZFHsZPqL3UmjSSl6G3JdG0NnwFBPsTN3pcA5vJoWEJff1UaHeVXTpGgtSW7GsksUI8cj/DndV
UzvDFjnJBgzajhtYLS9iuRA+WX951GC+JxXi21hDYvvg2rxZWeE2LdE+Ld0pPHfvfF+B7oL9DNh2
veW3eF/r+Tw+iSrvDwI7aaZftXra4qbj1qTgm6JGEjwY9mUEKA7ohv2fxPo4PqcuyiXFBd4unaTu
nzKbVZBVm5PPwis1m34bxTQxmbxDxl5lNSdSaVKMq2uE81PqQ2an/xadPL/exrEgXeVNOM41MFqc
ili2YqTm4CmaKfkEOvCwQ/Ot658J8psbEsJZPd2cw9INYEmxQmkdQd6pUSIaaxMvWs4924L6X2Td
6TOjPUMekAeCSCZhBZrEmPSmb5CLVdg6OMV/a0bFtlm5TmH0KIcGFRX3ID0GarckL9F2Zp1QVHFq
Sx9agVCdHeOnwm/F5MsNL2+BkPaDk3PKtYV9hRWzHeZnRA5eckOxewn9lr4e9erArO9dzZt8M59I
c/8oM43uVYs3fTaeEEM0aar8wyjGwXrcxEKP15malRfb1T5kIgQvynK7NW5zQXzp1xfv5RD6AYD8
KjSDoucPQJvfpfAu1IHb4IVMw13ygjQkm0Mli+gbHUyT40Kfa4uWsVMqZRQ9XhLIZUQXwvEQbaVr
IfGrLiy9lD2XkZe+kQGXiZuheet8TmPOSG+/JoU+pnBCq+ukjZ3t6wIAW85E1yRCQOMWM96O39Al
P0k9w46iyAJ0sLn9KqsmwHhKwAMfmB6nlN2NTOgAEmBzRR8TAGELACefxYKLL4WTOs0Dw1N+jRBI
w+19k19mv6ZWN4AcbUidFjCTfviOl0DXEK/W+hZ0d3wwRPTeJSNfKx7gQLQoH98+fx8WQuzd/oUX
wQ/8jRVkbEUgI2Fmzh26U1bkxWOFu2LcmJ/6eUcCPNuOt+pv+xK+Ziuby8TrdTeVeJYJ824Rc5dI
U+8HqVXg550m0WGDZeOdrlbLi/zMEBKmtM4QrL4jHQDk9KQMZzigXM7HHX3L+vaoQYJqmuKIC61V
xV8Fz8NITI7BNwOx1xIxI+JXJvmS/dYRtdPjPPKD+Xz8Dy0UsVOjGIZnfhYaIq98xI6Q1yPqV4fX
Qq3tf11wuOzXPMXwLlnM4miglw9q12UnrUnNd0+CTHxGwRU+9cTGZXqe93YklYK0YgosZUqXpWgK
zDvkH4TLuny9UAqRfyrehrcTW1L7cBNIVBMB3OzObNfzcWgaFTAsmVoTQXz6VLY+ZPYzZR9gxebU
fafrPG8s+mnzIn8glBpggCmIGkI1ztZDMKLTPhny0h4RVbmtFtnR1+OAIEcj65XwzLpso1Rv1Gwq
2JTgJnZ8EQ3HEpIMAfwmBw4bAirLw8Uv6Zw0W5y7nj+LuWfs7K5JGjFmc9kGfUP8I6DZviTsAjxW
dD1H/qmlLdPGLM9nZpj4zKodDg6zH67+34GQKdedLMN5KJSNsigReOPSyQuFn/Wymnjmy+Z4NQls
WWHSVN/C6zL8HzuOEXBAxDxT5DraiVKWk89035OOYD3cWbqQiGBsCRq3jA8TlTeMROJ4hds1mKLP
k+fbUIXTPlTS6xPzbNlIygPEydcNuI9J/cavriwTwum4s7gXm8d4g7aoReqM2h4Wn/VQUKl4VSJv
2JgGZRN2m9JJh1ax7rqxJzEO1gIHoZpwwHh91XpXOYlRMu9vgxEKsGMY86BW/OrwLVvfLt9dNEB/
mUI2lFY8mt48n4bHtavKnrMKfHN4sh7ivZln5Onn1JjAyEshxFzUhWWBJL7b6lfFh9/MwYGXQsnd
oqJ2/YoIggkigak3Q2awUZWDZa/K4LrRmWMM/XbtSz+DmFZKMqzXkc6Kr3Vb4dTzDTflJHJyMtW+
LCTITz1EqCf61ETaeuzxohfs7P+Nu1AHYCksQ0CfFR92WZhiZGyio64Aogqs+0nk7of23vvVNL1d
MpMUOQyGwt/sJW5eRThyCb6C+B+Z0QgMLVIF5aB5HLwiGbji7aQCt+EGxVOcMEGWQKGafpXfy8jB
E9UY/P4JW46RZulMmPHbdtGHa0eNvL5bl+/cqe+zFBtGehhFpKE6RgtWrgitYElrHrC0tQaShm3c
2CM9IbeKI4adz1k2yXnuqcrdSYJiBD2na2STQI/9PdFsh7oE26g9yFcyPnmVjtL3LSQSK8wVuPXB
gxVy9zaIV5ii2f74FK846RM1BNsailksfaIwRvA+mSizPJE7i8tiS2tJEbkQEm9WlcL/bGAxeZ02
6pV/2aIwNl0CVclGS1DxysiGIwoF9QDoY6mdneA9TIQGpBQwp+0+MXxpLkHmvvI/bwaXfg9nclCg
YlF7lsrXR8q6xVjCCSyDlaiJQtCvJDaotFaQXuYpiAfN85Ju62Jrznb94Z7yGewEPc7N4X5Nzx+8
72x7s9MuzD4BiUgt6z5UfFdKjiHwknHYA8QT9OyNPMQtq17BqHIgilTzi5Zf+t3Mm6gaZWKJ5jhM
fAs2RVVC6UdyzcxNYjhTqbw+Mzh4imuVCVyoU7tyEEV+dPghmXqi+akdTMVZ76mVnnI+z4gc8Em6
Q3QJW09BfCzJ6xANF4LSW4pqoKKBYmtgMf4sgyglzPlu2Rd3H/Y/TBQDfZEx0LFemePmIOFgPTYk
KHoEKHA/+XyrkVnhIS2thWqCBvKWdz7yAYSIbplkK5VJeB74929kAkwaPiAe/7goI3T5XETm3JK7
I/s5kNWyQ+S7bDHolOCpbxxwOXitUQqAATevfuLwatACZKb8ZZw6PHHF3pYs9DJmAAksqVdNQqkK
m5WnFeU1T2PYxjXiyjF4BItC1gAaeQw2AOodofcTj4sxDwOSGMk8ISbLSTTEXyeGNWO9CUy18rS3
qWwJTt0Ip3ZucwPgWTpd0JMxCetNWHG3XKTpg2cW+nJlMdlzDzD97CUnl4LeoeD1NlI+bjfar638
h+WZZYPhtz2TlbkiegKI/zfO8Z3SVxjS36Go9CsucLgNxPP/y3sfeQcGZvbB3kgAVsjIx/nWMiPj
7qFQSsjTZlKd5m844LdXQV9eg5gLcdKbvkK5Ls/ZwM0ikAvkwaQ6/g2WeAWWwDniQkK6vDQlAPX7
haTvl5gdYEbhjykc8wds7xsZrMzy+lpG+zPeM/8TRe+R7rWojKDjd9iYmo6RH0Aqw5j3of9CEuQR
gceeYtXZROvm6/IyG6x27Qc2bVBIyyef303/Sn7Ya7TMrQg8UuTn7WmxRcE3roNi/I2Dtj+g/9cf
/UB7O02n6z1U0ohfD+kYqzu025QJo3BEfL9Ak0dMiMeJZbSBP/doV+LLWxMMJ2ASDg2TG58pDlYo
0oq+9ZHMBx/p33jesI2JETpFokwYWxQzDRcRCAoCOJie5MIrEc5tew1inonzN+MKHb9oymDKP+6R
05LW71OPtHhuMeHXACFE/Vp+CChtSH7pMYg/vlfSqJumoYMc3zf4Sk9DVePtXzSBuNrAzBLGZ0FS
jiPArvlfUQ1V6I2SXsVru3Awybj+WbjckDnuY30rgLDPwhHAcxGP2t/dQ/pUervglW3kqeGxvX8P
91wwlwrWY2XJB2Org2YcDcx96N13mPGT5GhKdhgCJB2kVuu3Es6g9LVzmLqSddMhuuMQQPllX5Kt
v9lMUjOtz+m/No0E1l22DupLKiu114Hp2j7PQvx7c4kH3met3zPiLTIvSCaj9n0wRDnnGlOPDeaa
MMznQMyx1cWl65pLQovKiQW/ujC6WtcK+jaCjr2Kdd77niQP2kVcdDOBhbJSJ7SbWp2puAefr1Q8
F0K+4gQ87wcE3KGJ4GKawvuJZKmFIcQSY5TCJjeqokDO0XJgKCILyTt+YpxhlEHSfJ2WdNsIbNaz
7i+Zowanc9WeKeEPrH2KJBtNm4baRUmHV0MNzaeztSMFmO2GZYm2bRQWhCfbNWEfYoBPkaRq2m5x
Ak5E/ZMovVZNfUTeVz4i7HVe82DyjxB1hRxcBFvEmnzHYanJdzBf1AOp+g1mM/sX6sY2eeLqprCf
pwLFTvcqZuAXyT3HZUm9NXZMXXSfEdl0s7rYVRLMrrq/5gmlMgIlVHwDhON0yH6lVo6Rbg/I0Rtr
19zW+Y7ZNTk7olpa3WgEuELCFCMZGnrOU6oDSyzNnyMNGO3h1XxyJ+j5MVV1qoBV7xxf/pyNQWsY
617geV/wwXDEho51A15I7W7gU15zhAOX/jZgiMqH8XDBSE3nO7+1wXpKTRzB/V641G77aKOh9e7T
rbS4RNji39gU/mI0hEI/04fdY2YjD/r3Ar7lYBsk3lqcRvsMvankzwlpmq0h+P+7Ncx9NqDNIlB4
mfpmM6H875IV0OLBy4v+2KjJkOD+nbJ5jHKHSGMwNKk9qq6gFcdgMVC7o4GQ7f3x8Ns7MzoJMlXd
YbqCROcqZWrdu8vS4JqqPzR9kWt1NjA9zjhnQQkLIlcAp4suQbYAJxtWm6n74GXDPOXI8xfZbWUt
cMXWW5fGXpYIgDd2ZbYRUsqZaV/eGEr29IFOzSLI2FVOlAiNhZOBcvMOxuZ9nSuJXUGAwRxgQkJA
RDdFmqvJvXiZF3Dwr6p1SlwRpMI8rJp6cetyO++qBEuqEfmsTX04c96kpCgWOFIfMsmtxmvUSGxA
4tVOkeXV0DF+PSEWx/1KWD2rZt4aIAWxcQYlmE0Qeq3sySUjnEeDXVPKuDUF7DVQZysaHPiRmmYD
q8rcK0hJxN4MwjOA2esiwv+rd1Neaic4Dr95JAQs1kyulMrTQZmC8KtThx5XUz0KiK+DLpVp12we
1YtC/apKv9jLopG0GIIBgwxfVj5FYnjZIZH2UdgIoJiMWSJoqLwWqhYHNms3k1t3Lc22txN31VVZ
7DNtNTJgFuYikjTlN7Z1xzHNymLI7iM8j7U+uyGQerKejLYxBRMDmVOnIMCr7cEwZAAQXbVhbyFH
ojdcynq6ziliv8w2W1yZMUtzcTWnvrCSTxfg5OJJAzhKQ0PrJyX6iLtMB7BL0mhFTb/6k/flXU+v
LX9+maBsDYLjcmAIWDBI8LdkKIJX+/p6DpLNAQcdFryRglDOLjb2yNp8EdXh5gWla4+BrAAxUbzv
SFfmUrBjV8V+bwyiTsjx7fqnxCTFnGzD0RZAXCyV/87VZYsNpnsezDpyJ9Yj9Y+/LIrjawDq5DiX
/XY+vAuOn73o83lQUy+OPg2untThbc+y0zeRFvjOvdJE+CUUIusfwpmUPLna62L1zDGITXKHzFnK
JyngmJsNI+75Xhih7JzaDb9sJPArQ/57H96FjJhxa33QY11M44ajSagGFnKvxw5XrluJOx8y1AIr
HwvvmZW73fmN5s1rjcoVG1M/l+d6mHedF8wi7T7Qzh3+uWoFA8CPQUQ2ArTOikoG0wOrfADZoq+t
F2kE1ttgWZ/rcEWG7lxtjIn66GlifKkhl+GNvI6Z1hcOyVLshq4GZ9L06f+7/7RlRhNlIUs/s+Xx
qaZoW049sxHxdaAihsuNeTmDSuOVvresRrhq7HQSoTXqgvF0mFDKGM2w79J9+AkptXK987dIQbyf
/Ik+rnKmgazQnVnCbPsDrVzyVk/9yslfhSigfVuoUGbBJg/REQKnASdUznZ9+5ifZZ56MyblFzc7
EQKBy2jcxmkF/rBfVv48V0BJfKqbvbn8j92ZfJyiyo20wXgg2c9lzuQwT9i6PA8VzJNnI9h7VJHK
/SOeRDNb+GrOa0AC/eklmwaUvs5oaC7IdY04wOv2aO7Z4cK8fyZXxzH/AiAUJrs2BCOzMSZvIi03
vpXj0dglvUAopTNxaa0Pbxx+XrrniHG9TC12UnMShSb4FYjRnSYTLB9QJcdimJs2VeEdYoBe/U0s
q9ReKRE98NAl/+QhMUVQLFPBGZmbkC4fhvLpgE9B3NrPAVWL0RW3/3FflA6QVd2oU5x5a0jt9TnH
8cMKumEoh/4+t+W/6LdKVHRK+zxnUG6wuH4Acx36z8e/wZhHw0TvHQLfHVOK7Cw1yxIy0nunsBId
7irAGN8vsaXRriJbF8zedOmXl1wX/f67MCxyoElHvxqdJjyXv3JGZDZ16wlxnWalMes45yTN593e
PzDekK6pAc8vMric1uSJ0QqWAynD5FkuIYKMVEAlpn5DernlzwEZYL3H6MaE/VPVsuh0LxsH0a48
CSJdqU8VEfNkrG2Hv1NzAomdEXpYWxyDIY4Bl5TRyD4tyiXqv6q6p2dxYgik4aXVEW7sZNbRJlId
hARSocXq31Gku2uo7vNifx98a2/xdcymai8cF7aID/1ss+r+TaYaXno1wCF0we9odI1FOpJGQjqv
NSB6E4BmwL0hLiuHbV/8iHbZWxStLoQrONPKB7Ft6wXvVb21i2BsctQbuKEfrlem7D1Ypki6Qh3P
2d0yaUdP+kbvCbMJ5NqzpOsPGsog6MHfD3uA7ETpqtM44dtklLxW7VlEtK5sSuMIucplpTEWUSuy
I0nehlzWj77Ec1YVrjk1MBdRUJ0LWGB1xg4GOK2q8WJ5DgvLOlrf4huUFOSvK2c6n8P/SSdb5fpI
LApS6Ygzqj9xKdBirSBNexAbNo1IDHk/ue0Bt2Gcl+Elv73EaofCZ3qmxCNvtZKXNQE/9TPUchSA
aOegqJt+vfmutOhXEl3SJcEc3MTdtKnCGPvq3Qk1EDjvQxnyEGmEdWW6b74QRE1MIjk1ICLK6nSB
6PSeC68yNec2s8+Zt1ZfPt5k3qbF3KZ4VcPw4PS7pp36/rucWmc4Xlb2QZzdfykX0HNzDS4nN+WE
JIjpiS1dS252O/HPplr2zCF2GNrciw1BCBZ4WA5c9pKcbXGR4u+YFLTl/aNhSMCLGEucjnht7L92
5zckZvlUXey31Cux9tsFtmeDAjc9QDjGzhgtsYb864R9yDGCBH/17Hcn1FufJKUdob0yXQvPbkkC
Tsculn3glVrgVJrlRmSMMUpzM+vsKQ3xcfX6+rqy4NwxGZKhKpKQk6cHGHMtctBacz2dzOKUg902
Cdg76TrQT+tpnwIrRtJp5gfe4vy0vaQAlTzSdipywnONaElKsIV+X8lxjD9ZyG8FfM2/TECuOBai
srBhOlzhcIcLfFyOp2Ihq0fs7zq/+SNrTVKl2YjrgDxRHLDtytDcfRAbFtFqzD02ek4ZnCeaFljy
53n1VUNueKLpi5Kuk4an/Kfm/aAPaWXumezYVdeSAQjk+Z+V431ep+piOeTfbBcrginE+GAfMxXl
+ViiCVQwx6fxrNFNmzcrLfyZzJg3VojdmGXanX7+EivKRmrDZIeOcXE2CvJkr7dqrcTCBus4OzEf
GuGcTL63fpIAYl3Cz9NV+3jYqMmtfk+CQchxrp5tUKte5QRZ1CyAimSR4IwegjLxOlQw6hD00CBe
ejua0tioKccQt+5ecUPBu2yfs6wMWbhpb6QZw5MU1WC4SXb/rLZJobNZGP2PL2AsVlavA+oRM+F/
kDknl8MSC/pzIFkZYP46WFv0tolcmS9h+VsxfdXT6lp8BxBiBbyMn/aJTEv+gY+GB5hbc9MpYKn0
n6TNc7+a1YlLiYouwNcAoZcc4j4hFBr6fq2ov5uZ+9dk5QQ56alYDc4P1SfCs0gk5jHxjrBBN3f4
6whs0xQ5YNZwhVQBKngp/6re/JHgPUjI7qUdZ/l/TJXmZmoyTO/Nb7AE7UeyUhrwAOSXQ2yM2xCn
s9h8g5ZsemnFE3F+9NYwMwJvdCpjLfntIS3JTc6GlZo+2q0LNnSSZy/Dhlnxr+r7oFzPa5sT64NK
33duyAonrkNUPkrSf/dv02DtqyOrtjMeqOHkfiqKFV9OQE9d3Aiwqv9TOSLM+iH9gPPpPkdwcIha
o65RTFg9+knhMddiPP55vVj0Q3Q1slDUD4KKfKd02pFg+KRe6J7WhudgBwVs74IwkAmkQM4+S78H
JD/K5wXcRxUAG0Pl7Mz7Yp6+buXLlTQulZjhtaT2XFsH0o0y++cppPwIIhJHKhmKVu6pKOTfSkxA
KJ+OLK3WEzmyEqF+2njgM+15zmmUUmVIzzPr91qamDSXQFae3Dh5X+9Io+WIVEykDVQLFLcishj9
25qrQEuNcuhbbG1if8TFCc2FO1NJBzWPMDo2kUi9+prLIbm2vgQkSimxeLM8VMo+zOpKvbC15glG
x/HWIqO8PoJ9ZIBWc1qIyPWISYCGevzd8Mpxnx2Mzmau19h+2ftDtikscqbPtjD908iZTrI4ZkyB
dh9LAd+dlSTA5ctWgaE+SxBHQbdWhza8eWEuZxDSkMVSGBwY46GXDsyQk3TEqmG3qQk8emeSllrA
OPNceN08ve2YOA1AloqYZ/z6x/ChCnw31a2YOhIvHxQtAyF7khoAKQbvFpxKkGXcqUzGj9e8P9WF
SpZB9I0v5Om4XhDLYR/mb27BrdTM7hRvN2pkmm6XGmwRseFcB65QqI2VOWx7hokHbUq1a4WK0Frh
Gj6wGAhNpilxA0afR260NQOkJjh8y2ApU9sY91eMOB4A69sjgeLgWodFNXhTxbykND9zkY9+4TIx
RvnrgKs7gHlaRP6EXmnYa1N7taaer6N1dRHBbX2UV7xXTfUlJhUYUaDiqCnlqc7LAsQTwfhpbhBu
+vkYw4lLQyfCzl9bGRYg2jihzONV5wUJuavRWyOx2kJqsFl/XVQiE1Uqzj/VeiDaMbt9G1KYH2q7
RfD75T0zs7lc9r7tJChGwa7x0htOWOSt7mw/xhK6fRgJ9286npw47FXQUoj0bKcK+aX/CcOqYxpd
KzFeDSs//1lFL56jy3u8Tk7dU0L0qzx8pM409w6FVn15o+YTAOzjb7UEaoVavzw7RYsGrqASKPg1
ZOLXBRgtcmY79xFqd4ScGSWNKGUHL0eoSQEctCkzbL9MC2j272YAYZFjsfBl6k9AWl9VlV7IyEOj
RkQRuI4KzxcIbE7LxMWa5DTw42OJ4ku4nyIxzZKWM8aMm3d6o3u0HIqB1GC1lCxym4Cs6ljAKFwK
+dXPw02vff2Edep/i7NDPFSvRAByMVRY0RIYy7RGW++KwFZ2+ZZj/xeGsTy25YEWf6QRGok+B4lW
LTebUT6SPIi97CT8/KXgkEBDat19G3+K/Ow4zzefz5bOV0umcs1Q2EExqs4OxPr11ov9ReLauGm3
O2/uBUs4o1WlIxGGDhLsxjfg5fAYkT6pLzVBWE1/cr+ominQfMJiwFaygioMtRdf6qbGFmR0ktwX
y355CNcuB56iLNstyXCDElUtFBVMRzhx91Wz/GeN3upIBahoN1QdQuaP+wAWItpz78uHc96IxiP6
7a2OhKdeTJpsKV1pphOp/MQB/rqmAZe+3MNx42ei+e5613iuGvlqG8YAvGug76bw5kaWBZN0wC96
mSGsa9ZY3yRapSYael9iGZb7+gH0RlDWZv56kOYIrELT8DPtOltizzXiD5rZJmWtET6IOgwSnF4G
SvvvT5VU+CFiwIx2038PnOp1WKN0x3/l0GM1XXlw/ZtXyhm+v2nVmIjrVR6I8hFFq5yfpFn6K2B8
OTZYQ5jDzZxClwd8dhQAz2QE2r2vTPtWGdS+cL2HOUc/ADdTtYPw8SvZ07RsRNjJzjKGj4MRT8Ui
ATt69Cu6oqTCsbcjBD4Tw9ZUprBm5ZirCLtdeBAl5CEHgs8EojJx5mUluR5v00IDb4Y/xvF9v0h6
ZExUQWuX6bj2qYMiWGw1PSDTj9QOCeULF81zxmiY+o7RN2asts3tpEqyob9fL1SP0dfs2Tzd1z2I
h4cKioVXIOM/sN1RL8XeH1QGxHvJoFGdwve640cizNeNxXmLsSYkUH+BrHlcTYOBqDWc65JG/O7z
6wG0XtXxINPytDlFJ8l74HGfeiQI3QH88ImwRQepvMtLwFqArt6GSxJ8KDrIvwVS+V+L8debAU9I
BPIhG5sw6FgwhfXdEKX6Et1etzvu8GQhkEwyFufo+0sWGjNSgUfBaJxUNAHQbnzLhLon4gHjkhFF
Nv1NQLb8lMHcM5rPRszXYaUepoWbaEXwnZmGTjn0ihVJXyYsK3ZyxcL0jGRPXRHIEiNGhTBXRVEf
eiv2Szv5Md0wIplC26cJx+Qfr/XCk9Vh3Oc4LK10kiQA+7amgpK5ZA2+TJZEMz/ctEsX+iuFpKD7
RSkD8uZKh8+WxTni7NhflMASd1q8Mx7lsLItaRraiUJzVwqf8QrSHb0wMIw3wrslDv9qkmWS7NXE
NPL9ZBQDLlFrAO2gWHh35f8Ho8N000x129996ifc7aKVao/Lz3Rx3/RS6+QqakChucTc+g0iGD2H
4/yGLMjlkeElb+WEqIX4u4u2Utn6mNYvOpf3LfmGq787Cgshb9uaWL3A5c8zGPNNr1rhPscQEl8Y
CnKAf+t8SKsSdl+75Hdl8rzUeu76ZSPscTmhCYaPXfmCPLtK6pySDTCS+OvLcHQusZo9R1n43fQd
kb2I7E43l5R5h7Ix9oNYp3O2ZiIlhh95TCNaudmrDyBffavUGlvn84DvKUv8lMa3oyWYbkwGefEb
jIFfZVjs44DLHKksJPZYey65g3VgqZZrmrOY0KCyRYL6P3/LqkjNFyq80cpv7RXEOrWrs+qBlJ9M
2leDaD9BMuTrd97l1NFkY3KNbdb3jhphxTW+6PNl4xq9gTrNoq3PkqAGEoJLjZTJ7NyiA6M42Q47
cGmzYvhPrq05CaFdtE0ry3Mc+vXNQdFZqmtYJ97K1DCURGFg+Ih3l5bXFpzXpnP/n2xdD7rBc8R0
dV6U/Qv0Lu1zEULTUagUXvL/O82upRSogoVHQNdMXytXopP3Jc4m9RuxrZ2Vu7Hma6iPx75ymMBc
QqnALuqCybepeMECywz+rI1PqEjK520N2dmVNKjkUWiDTc7/WafDD0uRWsj3B3qzHVjyLvI9QZPV
npJ4ohYJj9qvwWT4nDct6E/3v2HS6Em+ik2HjnhIhWdtcB/XOMH6BuAmn2PN0iy4ceqCwy1LMNpv
MHBgcTEWpPMg/a72Kwve5rurEzhswjd225Ui+3JtIqI5yi/OtEDLbQnvYFZqdzLLkgaV0bfDXFZh
mm44wXZ/ulbBKulV3VY9NatLk19VnEGBubeTOAxTCkRvDSIwVIneDkA0ywvXomPVVhC8snwDH9Sc
vsmnccd0S8cLByMAONspVWSI6nGSiU1hxLKCOF1555vvrtc47DZY4Az1aNRqiMRh+2l2en5gOd/1
t3RjxAoaOR2t0WWwvQRJnf6PRt80vhVeiG2l2I8e7PaAQ5QaUVDi28cW5y0llq2rd8JdxZRLT1R4
MMAxEM7xfmrwQi4A7JN5ozObXq/IZ1Ba/jCtsFs5m+Zj/aTHZlL8TQZejEjFKsVdouenbcTpoDFc
voTQ5y0/k9ch+Vu1pUCg7Mm6IGGb5tvNx0RBDtAcQe+2N0ujNVxBH8b7kKtsldChw0qUZNxHA5/+
zZvK7fa3RGb/GxaEtC6MXlTqfbch+UNAgDlHyHzx5A+Q8AAt5rwtnBwKbuKYPoJhYdy/k3uYluPx
gyRxqqM5wHwG6iqdzY0IpLO7TPuHAXvB5zCkCyBT6nbiHOH//PYVS7kmWgYYgX7KxEh9rmQ/dlMJ
6gzsZPd5ALrmgTGrCzsE8n/SIuDNC+w7x0PPiUy0XCRv33d+DLRDGH1EEvKoRi7ZIkYm/6EdwoOA
+i21n+zFpdZcaKCgZx0VYjK8Q4hfpXhRN1Ycy5ZK9nMlsTqYqY2k6Kg63mPNul9NqLq3IbSWx+on
+zWKxMbtCaD/KknvKJ9gxwMY/EnGJMEhCv+eVL4XhaLBiu0d4jyiwiWJhfbH3KhCudcUwcd9Wddx
GMmacTe86EYz/esbntc1ayQcKxLWwo0EvCHi6mqN0ASopg6xzN5RsN/0/ygl3kuCH3L+ghUFJP+Z
weCxS9ZEqe90pIWX2TPSZapWsjOz4q5VbSgFZmn7MC/bFLBCP8LEEhN8dWMeJnuXrX2s4EzIeDOB
emhOwzrOKpGsOmiDDE3RcYFFYUkng+LYO2rxNGGNt9QA5eHKTZP29Zjj9NvMkEE0gnSUh53Dviyl
zubDYClKZP6uzjkQ1VOvR1cfS3qcTYWg+i9LiY3cj7xUtr0nbbxiXrR8ReJCvqhK/gM0vNPm7PiO
VgT4MwEo4maiALhOB+dYFXjWWbqhWqWZvBvorovfyBrHcVIa8yLIRgRqvnpXgFP0UCGafcxYk2aB
FySno090fVPTsbCauuiPPV1o5BSwvpYCsQ6RY9vDOytYiVA9UqpgHY/QstpzjOCjMM0Kqfv5WcX4
PAZWUWjXKFeppr66xMdZd7kOhHjegRZ+iCbkZBfE2qkmBJ3TD8FhHp7ZJMA96ZnebbpgS4l7BCOB
k59oQYAE2JezbhXu7HztHH5VZSwkb4g1ECbsZL4bwF3NECtkokQYVHPeYR2lzIyXbN/PYez4GBPP
NEy9RPrHGXFN5vQAxjPqgaWR8OXxTO7kaNe0eluVqjcMpWZETbOmZpAnjTh4YCj3zW+4VejvBb51
5r44l0pTH4JLID6ux79rrHInGxL1pp59euXCTPPGy0OuuhTv4QtorIDyzuK+YGdasTE636mswaPX
CVxy+CJ8OrgbqeeCFAoH0wTDmuSSvMxmwisgeZpGZMwJEGgwIt7ZaLP8uVCeV66vJbvRtREDGFHg
7F94Gy/HbTJkZxn8hhjnKBxS6Dh3I1xryEZ0Kn+7+fce6tck8aFtf2XxoWxrxQmAZDKlCgg0pu/c
0K4wc/bWgXvWQD/m9UnyS2dHF17RTtK/gGYbmga/Xzn/2A/gQL/E+fmhkWSBnGhlBhx6pWIkGdWR
keHhg/p6xUH2ik9MeGd6jN08AvtZwO7ErC8MWUzaorEA08sZnCPxxuq4YwzPzSrJpuHoKGeHtoRl
vyDiuw03eJr4SgFQDTK6R/l+1Ya309e90VLDKLRQM1Dan3OKBevMCfs2Vrt2AD6yIC/Bj9PEeV/T
EK5Hp+GMuXKlqDHw2ofROdBYb4VkDuLeIpDvQaV+O3R2IytrWI3ENTapB1+k5dlnjZBGZFfcXE1P
o01LCSg1C+yzoFB/EBH65K/ZH2UWBfwK+Zoc0iDGpALU8nTnWa8TXr/7r3KraT1wNjMyN/zrP92h
fIM4IhlB6e/YFnzaBEHc23ltPrP15R4tipReK3Na/a/Poi+QQWCQR2pk0aQrtTyXZ4RT0mvh2G84
o2vABw1kyymnIvmn0JzcqMQV41KWWn6doLMkWGxmvgqfjV3KdHy6PQozIOAkt9uFDwpPZx0DA8z3
acfB7ZCiybvwYPz+L53hyekq4MnmalBqnA5IDbHEyUXHMJqINNorBnenqpp4aX1iD+izQ57Bq9FK
VT0/A2ggbW7XE8OiWnYAIXyPvyH7ZqnvXmOMpbkUJluQbE3wjQ5/chNi+0Epse1xjgiGpf/3I34U
fEEOG2PvF+igCaZp1IeJcC4kZwRmvGfXYKUXpl/vV9eKKXjzMRwbTTjveRENKur4TPaGJWEbj1sS
8uPYyCp9DIfXQXkVhopK483NsF6/feu8ne1Od/gcZzMvVkk1p+9ewKV2/pE0eOms23M14opdy6Nb
F3pPjMD2doz7Bl1pLsRMQeuqJLBdPw3wXgSzBlj9qbzBZOfVHB1lx2zl9St4DeaaAv+yGiJ7gsTT
6U/aovXP1bdkQR1YrIvU83c6xUeKFCgqHeVTE2RP3lMGVt0AvvwHiRkfwu02f4gwZygwydflKr1J
1KzDpvpp+0sUgWIYZx+qr1Q43j1CiSAW/cr2ocleuiDcj+2Wy8wVxrS97zj1UAIDj0EiL72CXep0
X3sQXZlIT2bbhr3vlGRYmrfF8/LcLAY7lnwzF2F5IykzblfYfJKAPsGshP/lJGp6fYlsGT8+ddJH
aA5Ah3J40q3KK1kxjmVbB4FudFQb2+vAJdXwbfQ1zT8MM4i+0as9zWLVstADet14MeHq/CxIKl7z
imExFea37+f7LV+9jpb0K3SM1/zct7Zu/r41eIW66C4vaBys6+Hx7phXQWqCBXRp1vxq+PgI9NhI
vF+cpvQpwUjwiuLOF0QnxIhHv0yeJyfbusb6P2Po5AprsGDNsiGNt2itY0lv556YpYowZenfVVcv
3Yo/ROAzlC/fQrk07kfRBjQ8KerNEOELaFH2Y0b143s8TqHLmSRS4Gm+hWBNhdJl/6UrDa5LfJoJ
U1OIMbHM6SObz9X+hRRgyMXP41wgNP4ycRmWSxyQfsVa0BRQQE2sQyFlsD6PRU90IxZaQloly+Qk
de5dzC/xIpLkj5lK58LzrUmytooX5PuJ9wUwriBNFJVGafWv6LB4S9A92HV81+yAmjsbmfpy4OKy
6Kub115ebhh9//+5v4YDu1MBflQV1+7mKXVn0mjYMyBkRBXH7wSpXM5v+hcYND65XNj6m6lye++h
a0niebDG2K0WzF0GTHKcZntERKIDu0Ff9OlP+rjBY5EyPw+eWcWp/xbmzT5OOUODErub+x9MLr1q
M9DZtRvxPLwCmi4ecOic6JM9rUk+0dMrJAjVkLFOOqBezmOwicDht79uq/nBl+Pg+Nfloj3bJVGb
BF01J0hd2usbnoBHXwG4a4/Fb7EB7r8ps4M2S8aaO1dCa3f2fZ+5KceSZF8xz+gj7EbyCxvYC+x3
Zibf+U3CU8LmFGvoLmmXv8qkdmOIA+8P1CFUSXATCI7bDwSlOzOWO5SMHF4XtzMQc+FYDOngIAeo
UUkkV1aIYPNtFAJBQz1v6t6q1l71f3DDGEi8bjOLMBA022w+AzoTvPGvvNZaA+t3dyFXQyGv+V3C
ptyzuNtyv9YaI6i4Jreuaomsm3uwqE7k9cS424jAwtF/tZ1k1yMxiJ1uTRyPMOeZs769kiHPhKnF
MMDdtSh9o1lQbcSNZbgyfVIABCKbXKWvBMGPnankqHGjTSjYcz7Hb4Ml7gKrDVMOsuMnDiXGgK89
kwA+Kjf17cZXoa18gveIqU69lqy7/aqq9hXuxAzdBFplFYMX2Y75kqdBmF/CPw2F785Z36vgFVx7
7x0OisLGZQ2HRAhDbMhDYnnHL2Nt9T2rUfBABBdOvSO42ULMebNTQ11o5LUPRH3UMV0JaVBoI0F0
NPwrX+CGBqLfLIoy0RmMHwjEW9sFwQqIE4PNkxswbbL94GvdCrs8JNjYJNht3brxCzI2inwUbS5P
3PlD7+2Jv4/DS+lCwW5agO5DnPSYh+ZE/mi5B5iVIHUInzk8nvAUFhDma9RWbwNJ50jc2ArhWZ2L
jzkNQg0RwIekFjVxyXteeLXPOGz1H5jFV5VtHHN5eGwVu8i+/ZR+LeHk3OIylUiMVsjIjXCgOt0r
otwRRhpt9jD64XMICu8gL+2tAeCanXc9MXxusTLQgKwlPP3uzhpL1lGpihDjoC01kTAm9rhzSPIJ
RYsnZkugo1NYSmbn8am6idF8MA4bn+3hTj8FO9n0WcHKQSYOVVDS0Ujqf8I7iUJXXSJZUxnQJrX0
0RcAtHHTqakfEYhZmUgf7Y/bDYLA0XPoVpdMWdA5R6TDI2i9J2ENeeaUXGNZNMA+EemZBDo1oFHn
ueYH/M6pcffZ22VwtqIRVuGGn28Q1q7mX/1mxJ/HmfhrFTAdxARCfpHswG13klXRG+wQDdM6kyT4
krc/rgpKnm2dh+QnussvxkpRR+4InMp19WRYvxmdfIC9X2p+0H9GYvPQv6C93J4wNacG4sd8EWYj
Gtynll0j+Z5ZZOzn2znjRu9HJ3IZ5HXg1ByIzka9S3uZlA2+So0pxQ791i1a9XQVjGB6+GetQvL9
HOjU+oiIxMVbhFwDwMv2r6FcquU3kR9LefejgigliO0wFPNLw+B8GdkHQfvTblfDfTASqgFGgBZA
Kftg3vF3k+pJgncsuz+HX19hjoY+cLRxUREBdOdgVD9ej06PyXCjBHpGo94SXEQGo40XbsR9+Hft
U4euaFJo9TVR+dw1nPN0F9EmTxGBlMDPj3jnAQYj0B71vVpM6lBQZ8vk7SQlMJbxqQHQaWSCIupm
+lV6dFcLH8UgiOkq3x66xYPa3Ne9cmwbEs4EvtrZOr7hSjB8jZcQ2ulfMQpwYcMuWUzELMBHDcZW
iOJZX+MlSR/aYCLr2+WcJY6pDK9Hi2bpEZfR9kSPxblcwCmry1LIvvYSPR2u3a1BhnT92Ia7F+Vt
jpXZhgAkhVAWHGBYpzIwfbAswvXvnlw1knqF6P13xu1SsrgqJRlwsZx4OxmtmzOrpEIG7ZlPKZ0F
Ml7ReDcJg5zZtDkMME41KKcPjcyI+4JGMzpxSrKRph3wm3qYQ66FUfX9cO5jHcwKeMr0uVqAyzvN
qSEKGPlxjPyvxH11hPcUBssTO0k+WtCyyHTnxyqkS0BYuOerwpObDg/v4WERfnC+2qo9oFBJviPp
FxOh68FAl5NzIz701KfAoy68Fk9bzuK/LpL54mptyxuDWv4FORlQWbTiWcYp/EJszdxfamLkR/Iq
4aKBuRPYBGiwfQqSOO4bdLksnc0U8CVs4nHlHOHwmFjonwWfH1tDVG6kI8ZmknagH7b/6/JfUXoY
HKFTwXockaCX/KDVrdm21cHAZ0EXx9auGyq0AYkcJ0ZggiEewYCCaVsNWgZMqidJsLztR6lGYp2s
qOaiKFGNLnNaeu/6u9apr8MUKSp67sVc+8KGBvcfraBhx2zh/YumOVXGvT1zNaqOdoUW/jRJB0I7
rWw7ALkrXkQomP4RNFYwMMgRYSwcfxfvE+lY2S05bw/SMGXZBY6HKIjQVSPFpcVeQP/PFYeJSg2b
kozK/1y5HrDai6wnPiXDV3wkDI+Y6KY0KIdNEsgjO85gC4PpKfcjW/JuUMZ3CmtpQaoija6nYrh/
m+M2I0CK+/lM9BXyoDmFgM1HwJabDkqrd+ZEy4i1Gdg30j+h29/YB2a85nsGiVEMjCo4SQt+nbli
6BuOohgq9vhf0RjZvBkC/BAGlkXfulJkjH3ES3nLdXYROK583S3SBQUyNePoCPJTdDfRFDhXxQvr
kiAJrndmpKQPnZO+DJk4hmsoT2fZbjGP1Q2LQQhI/0YnhcxmF9RhfqdAZzGDUGaGyCdIf5DQW0qG
2vErH6ED+/ICNtYStgLmGkosVdTuvHyRhvqKeJoVIHItUYVH2hourwCQeLcXtyjaEtvdXwmvMVOP
+nfflwVCWuIPrShCEdR4aoPPuHVF1KYoK/bewLZpLFtJ7+X4VYhK0ihgg6gp7GB4OtynzTeeRepn
Qs3jOfzOpwRH+TZpvDB3NQNaBtX7uZ/RI7K8UGNQxTlJUzB35f9PlXtANcQKZFLh6CCgdCydhAWI
1Ppyh9WvBCZqXQKRx6r6XwQXY9KKDVtZT9S8Rtvi+Nztb+mGnp++oppkZ2xWfdsoZ83f+PKJWPLp
GJcX++XujjVXwgaIA1SttvIzohnFrpUhL9L19WnAbbDFht4LODAqpFc7A1CLfVhh9+RNpCSt3K2V
XoJ2MRiR9EBazWlBTiz9Fij+xM63EdJ6E47/2rcuQrnsODEWRcwn8HeLNfJmQD0gNPP5rGSoBUIO
YqqLt+ulgZ5qiQ9iz24PobskX6mPQexjH+8ZcaAESsEGs5pxNIywPIVLFwTJd0MRjSJKNYmKdzS+
Lypnw/sVSaifTLmox5A2vLyGGWQXb9KM0Pz9/LTrFON/A8rjnD3BLn6l1WevW0LaFDUw/ROeyA9u
BasTevbRV1tkTVHY1HiyrHccFJ0l5uS6ep2HkjXpUwBOIhD0bRY6JTwXhkNg7KxssNtdc3Oncq4o
kcnBL0Yacf8Fw0ldhawoTQGfZSWRcbhqtcQnoLnsUNZu+77OtzVcv+6G26h9jegdpT6ix3YXTFEc
2ta9hLxm2G7oNP7yzrvT9Mn0a43xvW82hjVGzsRtxfHvdFYegaPnwe9eBpPokFTVuyImm85ZzmqS
kn2/ZMLYc1+FFt5FOhSqHc+KkeYVD2vhLqzba3vZpNv8mIlQ6lxLNnfn55XiQhlPMt5W+MByEa1+
3vgiXuAb14eg4pU7qF/3bR1ho+vD8cqSsV1qqGO9zscQX0te7vZXH4rqopI2mjhNtysgxReo0X2w
0ZJCw0z3+ovOuu6GOpDesGWe2zc7RR6d1OmBb2GVklNd+zPa+IALpD9WJmAQpQqlrwwMHnDBE/A5
LqiQGB1UxC8BYKvOltpOi6VbLBUjoKZW7jqi5tqotIzMdkRbv2VviCSNpmcZ1GnzmAXfEhgw//Cb
uwE8xJNOcGmoLqdQVfTtR99FUAJ+GxyohciOo5xbh0iBGiliN+I5qV3/3qvQMEajc0frXrh6Bz3d
Mtaty1GEb3M2pxoOJFBSmpRwZZEDfEBrKvMXYtPOYGjmDvdrlUhUXp6u4Pj0zY3N4Lrwh12qycUN
edI+GLwxgOKqJrath9LLN+FLj0lQZOIPRqOs5qNmM9Er6NYgcW1s7EaxKkp8M+xHxeNKQ7ok42uu
hkNMjuj8F4kKAESciVLHIxhZfvXte1uD8U0FaUU40QYj1vjrXZCgUxym0n572M83CXZdoXZVhUA5
/IWFseTUJSxw6qt5gxdtnLGmC4Wq1YScmMxfIPXOA+aq5TksJRsYCxBNu3PRcYW3DWlixg2FeALe
eZGA27HoGUY4Je8UmZTf5SKrnotJCXH7bxxFKXaJuqC0UhxRFG8BTrCreUPq/RgIax0LDDG2YoZI
MaN9pqxsyANtIZQEtVPinUbSzrQ73/lP9y0+Nn0294kyJzOZDT7nLWFykRQaZ8y2iJ81eBOuzrKT
q6LEuBkmoU9Z9hZuUUPD4rkd2ADGxjiEcusTNmArf/rJQuV9jStd2M9OrJ6rYHC+Vfgn6HlTfgCC
1b3jLfprgKicKj5XyhD4Yy8Q8yb44uIsNcLsmpFRsfK61So08snVFyc/TXRaexmAT3AzsstK9BRg
+z4NmhbO4zGrg/hh5qEQ/Lye8lFxRNbgbK2r3xuxYGPRBYKBR0EzuQVm1/GgY0zbGVaDHQ6aVtWE
aZMR5JcUEtVF3gyuej1fv0wTlvXrRVG7uEmu7EaXOrEjzkgiBa9akIFfH0DoQ98kcDerclTNADj3
3FDA0dxPSlbVORHurcaicRnG/PUZrvnOu69zsOpHEalbaODUz4YKixszRDC7S45etETVp2T25l5v
+zx/+WwZEPrV1/XeK1ynbGZeo80m+PVuV08cNtRrENRTOTBvxkMrGdKohPR+7x3aUaXgsFSxFLQ8
a+KTcn9OF4VunqLOtpyO2+gye9iya7PCDo1H97D8OaRW7+IE8+JNzleHZp7A8Cu3pWX0nc+BKv6g
P9aGNy/2sfw30we1OwNipsoYuf3P+F66oigzzmitaCapC+6QbzR7lf8zfb1CZYPLpZINLQEBwiiN
Dcf8qq2TCG6lR8UPbXJqzu0dc7ZxA28411DVpjTbP6d45h0dRWBIS+kSOo3TC1Wi6yXRIzJNpbeW
fMB1ESWS/YQ5qdS72C1DCYvtV7VBZ+IWhL/bB63LhMXCMyaC00aL4CJdgvdIuYH0zefpZYJdyb21
6JjfpxNf8gb74JvBwNRFwLCtPnwxxrV/eer9uvd++MD5RV6PemX4pUTrPg3G/D8vFnGwV4IzSPBb
9OJ9shtjG+0y18KrEabU52WCWwzZYfMUwRYkm75UAbfeYiUUOwARaspq/A7jebkl4/HnlH/qFBR7
rdlpDzkj0GQenhNw9bOsOryurDmgN+9+GTvwcvMy/iVOG4LVXGTcfuvz4gtVGoN1WRW/czGXWCKd
+bfQr1C7XbDc12jFfiTxhd29tyRGu1XEBKRglg5UPXhgcJ+ESonOoL9KN/aPpgMjzf6qUGRxkMqT
3y/GZg2omDouPToKu7HYbL3pdVeWxtVSPL8GPsxOUn8pBhs4pSUEJijXiq1QeHgu+LYTvtFMRBrO
Vp9Ac1Uk72n3x3B7HUtdDYF0Rw/yFQ+yWlfdLfholK9vye4EZfYr29MUqRywBRhvsfIs2gaKJ0uw
CN5872tuOVk0MvYzLWC18xljAME4z5myrcd/L24oTGoBtSt3IUViyVHgArd4YaWulc4bcDsiCmz9
3xQtU1mRhgMPavnBZWEw2Jsah+WaxlI6lE7ZKLbAL5kjGqY5CNXOF1wqxogit6U1kO09gQQvWOH/
VBeCLzXOOxkRuh/rEZOBGqeTZzWAmS0EUVQulGSeTQMG2NQ60OWbFjzoDMwGdGRMN1AL823NCOOD
COICDsrhojL9DDGddXQs76Q1lHhADUmF9QYEt+oSmbmauMVo9MszP55lGEMaevWpk4FhYOUJsQyG
EHLLPduWCZk1XLP3875UwiCQL/6JJwnWgw5IP4HjOTrIuCpY6kgF58E+3jP9B01zRRxEjaTLWq/E
ihAsHR/TydbEmJv18i27YKqg34zHCEgFVkdPtBrYD2fhCRuvQxZAHoZflPc+fHKDXovx/64qKolr
WixYRRs0LP2Ph0Zu6oiJSteFS5iXM4CeZOxhCsXmNRbyAjzbqU1CcPR+jj3bMwVLi6cIGcpr0/F0
271Tn/Q2aiX4JN+W+NFkbya/zWkrw8sx0TD0k6Gm8neaNVt7swKzC7wh7vG6UXyhFGD6fLhocRZe
osfVcCPiLFkkPVKtFz6uWWf1q8LAAVM5eCAHQrsFghpRKNDXq7qZFddPZHno1IAtBeuEPYs1gVnC
80uohAT8WwNkR4BCQpDr8DTzRNiabiL9Zx/PWfg0DPd3NaU913ILG+8l8y36TqyQXA+NysN8zJWF
9foL4LBmRbrwnwf3oSk10vnkD4pgRJn89mEsEs6/rZyy5UNl/NTGOkXiwDzH7fzLw19ViSipV0y8
Z33hNMnrzuEGm4Vgq3a/GLNqH58hvsaulLd8x3wYY9TArQex6Fq8RpNMUbOyg8TVLOVOG9jojU2y
vTxT/64XzGfzNQ1TpvqiUwnp+9F8sp9FtcuhIyuK7V8fzPkKZZrYH6zIe7I/Tdgfxk3+26lVP3tS
T6CUuG7AmuMinN3IyyIr12JBsRWRoOAEjU5BCSabFVWxtO7yHEaIcr7bUBhlYFUZrqiV4z9WA8vx
Zc/enWlkAbeInd0tAQyxPYrvcm+qowkB6A7vZluQUokfNFsYiuvT5bkH/1g1Vkyyg+2ZODmx/h3P
iwMilIU0K4Si/IWoQbjgadH3hGmMSDf0EdfZQD3d1viXZio2V5oCv0V4uGLdV4Yqxo5BMjXwhiyd
lWw+k5Zqp8yxHRmzWufv9AZg6h27aj/RRn4uu5xcpTDvMsLWrNZSzhQVM9Y58J/XHoX21F6uo3TP
/GQGeMIcyDG7eF5XgYnWMawXSWxp9U61G5CZuRMdJjreYCUldcAfDQGY/RdxtCPPeDnWOBKVftSA
BLTjH9dlaDg9Au7Mkby1h+E3aNy+gtFNRCbTYTrqMnhWa9g7mm3q5BdZ51qtTi1QvinVj5775ddS
Jvi/7HR7UQC5Z4rvt7hDXPNUT45EtNRaK3ngNV5FEXuP8jiiJrQwecXB1bxTz0OXS8dGitfP97IP
z/sxWfek+KhLkK2sFZPnmfOTihHn0VtNeReQzqCLSwCC9RRqr/0NZBokFVoFqF09kittuGwJSb3+
5ZS1/99gBYu5ccC+IuQaFRBBgTiOBsWTBpFCSEEAWQ2O2A0SnSkJkwz7uEVF6amLVYvj5sQqImV8
QHcYD7UApPhAO7NTxnNTZSB6KBPWaoxs2VqmpEmwzcgIdeO3EGGQwKasWZvUK/HsCoL7iE3lXFhT
1CJWwB8Vc3rACdYIx1CXxqDz0sW9w0JWHg6X/qzRlfaaXcSlSkPL0tdQ6Jv7UV6OkOK7j7Dqul91
JuBAcw8OoqR8UF5OZem5HmmtYy2c7+iQCgstiDyNyCbFmk0BLP+mbRgyFw2G4a/U2kbxEbQ3pNGc
F5cItAtC7NuddT7Vfx+ZH6nyMbnqLfpSQp5oqM2AUNyWZgbmhkM41hZMXb+lZlI1Ncv0WqqvLlyN
vr+awZ5xGiwbHrfmQvVILThSYBcR4yhVMLjg4OiZe2OkxM9Y69i9/L6j5HN2BrpobZGdHwjflJ1q
CC8KaNb0OkUK5XQ6gLpkJ69+IDndErdtOSGsOkqwtUH14opsdPgX/6bn12OI1Kd9OgaR690qqLod
jRQFjkzn9g8iDyhjmhQoQJTQ8kvFIoHFAJ96zZQop2Xpe3BuIq30LvaCBXvYZHUNdNo4p3EW6nJN
5tJU4hxuuCJH4/OJuVr+tAy1rnKE2oeaPGXuxakJAaCWKO08d3oRrO13BkcIUuQicAbM9qXrNsX6
ICVSlgwlFCvN6lypUD7o1OcfMllGjfxfQfjNXBeNjEiBfKExV0hli52hclzJvJSXlGhcYt6yEDEd
NLfCgy7LkZ9HPO2ijfh9eykKJ/H6OXln64WL45BFz3VCEd0o6NnMhEJZCGRRKR7R2y4hv2u2Mkf7
AhgTSiDae4jxtMlhEcvEDgGuOCVv4sUg4gW0nrKiiB0227vI/hnvlQCxDGt1dJk22KHzmtsSrRrH
QdbQDo6+g01Wd2W2SRo3qTIOXgAbRCAnX1n9xkBljBNvMEe1U4QhEAGd4b/1sLVPRFy4vai0haiL
GHR1ESR93m4Fd039Vh6JB2eE+YbW+2HRfdaq2/0/K+vtNvv2Yu14HIWUy1aIcrM4LgSNQH8wreDD
SD2TaCpXNfMAhv2XQtIHa+IbxH5Qyj93WMLIl5hqIhW31c+n1jKydtApx87edQpR0cMuzJlfdZlC
jScXzEZpLBdt8OcMZK/K2Et7+YvK/qlQ0zYqPvo3FQxgq9/7Iab5+mE6ZXcE9+1/2Fsgabub0G2J
KHB1/7uhKphkYhYKNLS5gfYQvWm0wh9ZWeVy7RgNDCfwsrBZ/oc1awH2JAeq+bYCcCVdD76mBfCD
hjKLHiocP1eoUyB/wmUrpm1A++/NJ29KmZ1wCMTz8UvvIJQeYjdrT2C4meq5pdTVeZEYWCKlvlG6
cQdkthPmzqpbx6kNDnK2OYWkPEM278wvy6K8PjTt70DKX5MvWI3o7Y/0OWWRM5TaLx7ZcH3dVLDD
DhvRc64PjUlNuSusXtH6LCiZzTK8WMSaJmBrpnSHm5YR1KXMNFEeDNJqwt9CLn+3qa4g5adB47LF
SBYk1HbGTqO04mHqRaBgt83DL/adBpoMel9acxGImjC/T3DmNjIieieUuYDLgDbefGQcJE86dCkT
NwNK5Trpxu/Sf50n3Ffzhi2YkHNYC9dsdA0uwHI/5Y1hnw9Rcbh+6+nJfFHfepyQKMIil0r/nhP2
KN4Af1HaSZhMs/xpA9XlbbKUHKGbKU+Sp0edE0lZd0sklmh9ywk5vu8FBOBvKTxuDk8vYdKf+s38
cwGrWLLV0HC5pzoqdt7oZjjhNMAOwLaP2mMWNhTt9DQUc8uLl06BtZptis5rXY939fZBGO5FhbZc
75Usp8g51CLT6OAyRLZGVUjZUcAyxoY2eH/48LkmsOEkN67vuSkHTq5KRrsOCZY+yrvKoOn8ENlr
GNusy0F1h3sj931FA0eD9kDu3beALdrtDPTHpxehI98ZXuZCpEC6loxiKzzOL+ZYuUtK4o9c+lqr
p3Ijm6qy8IdMw9Yz68Id32R2LI3/JFLm0m7kluwqE6MDAFtT7wZ+MbZi8RB4mfRROcTIz/0Jxul0
mSvx8Xalt3ZM67dUoUDen8SdWcH3HaPaL47KIBiDcIavQtLfNXzoA9Z5/7Ju+TN9ouJxT/oYZBlm
KBCkDUtFbyP1UGD8WYyN+GNUrk0OmSUxdPP/DnwllOvrqaWl0cZwyPHBTTycru3CvrDXyxw1fcRD
Jh0pSx915VBU4Yy4DneMEmBn0uBvi5bmtZA8gw41PtqcZw6x8uz43xZdNazamHIN75GNucHYD7iy
D096ZJu0VUB0xk8T/c9GwH2cBw1FsU6wufF1+Tt8w1yyR8jqci30bbdgHdscJH3Qr4web6OaLGj/
c6KJKBkz9M+VLN0IUBpsYbV0Xy1NYKsmhvGcGSndRbFPVb4Rrj8nLHxfqUpevmLTa/o8FBRDFy5q
fTnr2ZIuyJ/nVaBoJc9G/eqi8oiRsip7hFi/YLzcl3G+HUJRZFmjAt81riyD0pUkO96ZkWLkKpQv
Xd+92vlfH+vssVaYomh3ExX4c10LEoDJDFKe3vWdZuf35h5tZSDNs/txK1KGDAGgTEHgyijUTsDe
FZkbE/hdNlQ7Q7IUH6sTsrNLg43rDTLckoAHI1oJY2uU6WkrAWnb8b4Te9Khq9cQp4YBWQfQeUOz
YhM/J8BybEqD0MDmt3tpo7BL7ZG17ywYDDVKFgvNyAifrBxIU4sNUHlQ7IW7Yk2I2jrXM1yZ0ZpR
Sj8N1epddLiqc7zU0Jjlt6+QTqet0UatBjxvHYVdvXxBRGsaLn/aWS6B2LEXpZK0ZKrwDtvARfXv
u29zjvGCXCPT8+Xw/0SrZRFF2fxFMOgPHE6fYC9W3/330xXwY6DbcqgRv9/84hbTbN/6xhni5H0D
JHZvZ0QZwAwo1LxVFAPUShkvAOUb47/vvZnJHVUXmsSGeiA++7SXyM9H8ExZAhx0eYVdTNmms8g7
bwhVWZhs6bxRP0nph/gjdrjFYPrjRoRzRNy+SJwEpKoBBGQ0k8t+KRMiy2IbDS6ktNlVqBt6Qx+N
hIrBHQAcMoo0+gEzfRpWzuncvt6vw/4zyfrgp2fujeRSwHb3qR2MNiuCRV8AOwzfAqBAXBDWk9oI
//52uBU/S3LRC909EIx7scTsA1QNNnzwG+/wpKJBq3Se1CFXNdWtaFLDDN4p0Ai3BPrlAbvS908X
enyuX+rYkyEzL4tZez4IgIaztY9pQlv9KFLcc9G4BX3dIkLt8iniofzsZzeHPipVXkEGdtwAqoHG
owYtbCELv9GsjbOYuNwQ7hbm8nALLpA1arcmr/k0Klkzu2j0l6WO+uQKWMZpw3ZE4JOtdEiVdRxg
TU+m7Uoo57181r9stiyf8IKDjqA0fZlThaAXAy6HilJ3OpNYeiSx8diROA2xByPXo/puXaN9fFiL
EsBxSKjxCqj2a1xZ4gjXCuWqnU9vjf0MCFMn/bgtV9NrjorlBIJQtZ5dXPAPS51HlC11FaJet+ol
OtTnG7HvawP+Px8TL+7oYBO5mE8yg3wPc+7E1/LAQCryi7vrANps1iJw3uaMuHt94XqT+ukJjWM+
K+zC0jq/UXNkUw3NTQrkayOhJKDFgNAel45VL/R7vdLkS2aCNx0iODxDv2XNAkBUWxulYev6Cpd8
IgPsJms1mdJi/FTyZfB3ySvlx/RGa4gLcgZ38/4fZDadzUIxfwFQsJEhB2uuJSib9f8I0cTzHbgH
qla9O5cGVfMkj305gvQ/FeiymHKRTRe9yEr/vySCOIPsgou4YwSt0dJfdmxLpet0SOMgYexysGPn
uqzV6FvdQw8RC3KKlyZIYD7XZMA+FEkc1R643FGNxDFcOxESreDVNJWTFE8w0mhc2yfpEBKVmKNi
MRYhBAuK23d9+86Dwcxdc+FD5VyiN4wZq9vec2n6sO85Nxtn177NhRQ6yW9k/Ve8Hj1Y0tixfql0
TOVoQnwtaq9R6uBUtWtxyd73J/ugBgCMQd64aYwfEA8tMUAbZc3Aob3jIMSkgAXCVehiaJZpt/eZ
aUm8yyZxVOqepDRR028s1sy2AkVO/SA+2vnz+lrd85h4dmzkh/M8wTVdyRMvGCJCgx12B3rF/RHL
L2hpuBcMkmG8jUL5H3W8CvIM2aw5IXaZ1OpP90E6F+ErxSKl0a96sHmqU8FNOz//47T+1PVlzZLw
SO1aqES6RrnCkSJ/M/IEYXW1dNlVhV+dAcnDivq15yNip1R8WdcmXmx3/hfklFzePv/kuhxBz03X
IC45LcN2Xu5nIdnMr5GZ6vMrKnfZbN84Zl4HYsLl+avbV8pPoMogWvyNrGqSk3r6cDHRjZZhGpHa
SLu2j6VihL5er1zTeS6FxsMXTlwJQ5IxyZbJhJragQzBOdfcPOfHlG4nzyHVmes9rS2s74+64Nq7
YfLlx4RnZhz8a9ukHmtEgHRN6kjzF0haWzEoNKDZXtLB+9FdL0Uh3BurKf3AP47YXZk+CpFZcpLV
LRz2pegDN1MD1J/Dx+zw3COejj63hUUE+8U+pHZ4Qx5v3x+4icii5Asd2sOGXWIxcGaIBIDQkVgo
Wbe9nnxnA34+/ck2JZn6S5viiMZwBbcUWDYZS1mJuMb5WmUTLIJChFJMLTqnkgxbzofT+JvnjB1q
9sdeKdMZAZJAAQdwYz9E6gf+u3PFpJsI1ivbfh2RswKp7v/cLMZFnBurOzVmVRO9xJ59XfTi0+uy
PyOmWoSeVqxsKvcBj1MA+McVs+P27hOZwtyC2EbzKwIUWn/5VPnjVfhiMEq2RFBzAsZDAPpaEnF1
ls/mJF8lpiteJevOPc+HPAo88GZ+RD75fOuHeeqtRy19OsXR/7YF9PbRA9WHaOTEYT/UDAoMD7Cm
RnU0UuqU2ZMfLdWF5kw0PkOzIEPiJ+ewZSRyU23SnnOZS/Byr4NRXJCzaAHCCTykXkYHzzgQK6kP
grc2L0xTCSDZCcxxBGvXzN/j3TWEnF2jKXvANmqWFC6lZotwLx7MsB/KyN0iNUAH1J7KntSMFYi+
Bq/cz9GoNU/q5ajngfgJy8/BPDgj5NEejruYnFLDSEhlC4FYU4+KniQPFGe3wYG68xdLcAtGDpgW
hFqQJEv/GZpFObzJywM8eLGceU+miscoW1PZc4+x+Drq4X3tQ0SE6TR996qaL4cmRTs3a29EN8ZK
tY7vq4CaSYmMXK94I9pjh5eXIKkpPuLpeY2tp22Ei8sLlnvqEUUtF8ya8MPMsMTu0YT6keCJC1P1
dCoPfpXn718cEEldMJ/0/PwIa2SDfQpO8bCtvRO56W2en5NuxkuCevAer7FPfVKqreNb+2LUdjwW
01HsA0rqYoCAvPNIjUoz8J0ydzK8NGlEzKTWgmGd3xR0d7oX+l+Q0JkJlQqOjIEoSZeQq0ERmyoR
mZwyEt3uZ3N/FiyRtr0bvN+J1R+ecI77dbmfCp97+DW1oO6qhBCP5td5PlES9IxD8hPHBC11s/oz
4ytGEpezsUooCRGUKdo3eLzD13Fyf/vczvH6zuGFzNU0rH0TIFQmzTIoyI7zh0mwrB016VGLhupC
N74F6hlE0PMucwie85scO+krh3nwRidNU2buB/39ON/BZvMd81M5Ko96I+jMV7HbJwjp7h5uowlK
+lvaP7Es//O+WDO0O0uznbAAQdYybun0e3Syr5v/zwqgNRdj5Y89z8blqzbzqQOBrswnJY+VdhhZ
+Mtj0AtatEzV9Rx7mwPxVVTme4ArUOxx1i+H/o5J9GTI2auSsyezIOqGRm/LVb9PQUCEv2d6Rtzn
EbgAOgkBKJ09E+A1ckBoEzDXLnwz3g/ZVnTmlL4HNHy5a+CKpipdt2s68UWBYePuu1dRr5+E7QwW
ZdI5E7T0EVW1gQBIp0Wu2+LoNx1g++7t85wXC0nS550BC0/LEe2OAj4mr7Tat9g/SL6zW843XHAZ
1lUedK4eGFE2vZflpZrB4HqGLMTLvxoLWrtVZaw6PnST5u+XjTH4RWprS+xwEC1bjChgDkdawL81
sEuX2ew8UIiMQyCtMfH50l2PP2GAyzbvJP+SlWEAFpkvvWJvMdb10TZZuci4lEB4qt5gnpUIbj/z
laHcvvkfJdLBiQbAKWrkvEz4/I9lpkO1leY8ShPxqHLgaVzuW2zjZUefFu+wallSW4JBDVmSCDaF
olPvDyY22zx9E2+QwW9FCAkcpSnXihA0O/UiX6kB42GLEM6dqyP0rBxDpAsb2Drc+4aDphpEKX0f
yY/BAr/C5ElnxH1V9KVykpISSJZ9LeYNhNyoLZirbQdeukJg11S3L9aiKbKkyZttBV/EaVb6Y487
HaD7sRE05NPZkfCJUp/aLLSBXfIMYFBUmbxAiCVVZa09LfHYXkFXqurbPaHc3uHyBCrQ8GwqYeBi
dLHckbVLd50lCiaU/rLtVNyLXpFOOJd+IshYtsnRH19MEYdkWk8kQTxWiAin2vJI3429cS9OB5FL
U2Ck0V2qr2VTKV4/BDEsvqvWRUkogARldU5iXI/SD8BMITWXAh2NFKUFYW6TdSFGhks1ksFeW7sE
nWqBGRsnMP82VJj3uh0NC3NLnpPjzait+RomF7dQYZ7KLdMS7Y3eEdSLDb4Ayo2VErGE+I+nqK+h
8HUFlQ8ftRdVlosMtkLzzBPmqNqsDflTo6SK3zj8X+Ks0KBuBlPyrQ/64b22Um1NYx1wx8/Usjwi
PzcHtmiPQRYxAIpNJN9jIOAeojuUtB5PD01YjtDctSEyypvsHOkaVnmOz57GLuFR004EkpX54yoF
HULhXVh36Z5KjNEhmYaoeSlmoFc5OdksYq8VWnvKZMlcekvSYGDppXEjYFLYa7r16ZI57ZKjcAM5
MKGkYkQ/qemlWRhA7iMMhpTkz92t/GyXGUn1YyrTZWrJqYi+JYL8eZCrWqbJP/aIgIxFgLqAId6p
leFWMIYzNa+e25CKEMSW2sNQ+w3z0dAik31NoCZOSFsSF04TKvnizaZXW+vrasXGI97PrmUL8uY6
M0GvIoU904oeqDRA+rdDiCSFP8rWQz8Xp+sBiTn0U2CqJ4gjdaWwHJS3yYfvy6WfUXMGP8Ebktdx
jvm2hcU+Hlag0gF/0tskNNWOdkyzft1zU+68VvO3FHR+zihPnszpbBIKVRF8ZM18u1yQNkJThb0u
LSSDi8wkB5lICwLpTgap7/ky5s1Jhy4FiwzO1hJ3jXeJAmwVnOpfM3SfjOK6g4wvtmsN8K+vALwO
Wov3SEt4W1fgxG7WQ5P9wGaxiJfKyMPa8iMdRFE+ypfUSk33orka6mZU/czzr7txb3lNOSz9GC0x
Kv4Lbwcmz+tOAprQ82IL+LpUAHbxcApqMmrn0tbDTiUI3YTECJ1HTjfnQvR07smDutMb0jJ3LJHR
hZ7wdWGbx4RtSizr26R1BoWH8UPSrrol7GdZy3aSP+m3FABJuN8L2sdtMdhHchpYSenM42DGcLYh
W2VeJsn35QYrcv8UD0OGdoI1RnKqS+5U67ypa/d6Nn/PYwjxWB4PKwPrETr56X+esH7j85Z1CsEx
xsH4dOh2R2Mk4XHbtQ5i/XktbChqKafZ00gA1QKxPiWG6DDHlGMreiWB79GYU6Zs4kILzlXpGn6b
UIL+Zvl3YNUlC2xOmKhNCMFuSaW/qGEuQIk0ZAk0u+ggyZNVo4n20yQarbeSAf00CbyDwwQOu5vP
TttWKykaMa9oYRY/mtNY15l2GRKjArG6NLVIWq3BLvlZOWdxdz/nvkOQAd46KpGfSKticvUlTZOw
XVakvN3lVxu5ygbTnsav3g4XJ3BlWD5REtoeF6COrHlD6N+th6LKsX/Ojo/8a//wPuZBv37lc0E2
zoDIe0P6d2d0APSkwo7bJsd75q4lfrQUCbAVzTvI6V/QL+i/zzkmQd2iOPongB+cOZCL95IGwMww
FbWx07mW1gNkGbhIxwzNWz5IM/xy2YcYDGPTXnKPHnxBcxe9V2V6/3+i7HhlQgFblzgBZX1nf+4O
Xm5vRX00xEUsX+/Pw4P10NP6TK2thr6/AIiXGtKLffIAnaOifwyWs98ffKao5l4/sFkxZL9qSmtK
hlx6owU7/ya25sjfO1/r2cSMX3nuwcsbZXgPShGhGb38nehYxCNYyWpON/QyEcHjMlLQ9s+hFaNQ
DBYTgis7FfZztaY8MUqDItXRpti8c1TKeULeze8hGpptrJrvVJgHKbYdKO7rnKgvhu8scGvLx7bE
PSJOEj32eKShrgyqcZfMkM4eqCUmBqZFLippfhRQaYHZk/7DqzOxc/EzpV8Ll0l3FFCEQJF99+b6
xIdAYtQpW34zPqb45fLHumrxIjEzXuJQwNI0ZMdujFnGr2SELeYNZUuckPeCHXLzJv8QseufsGhX
oAy78RYiOWFn7cfidPrFYNdxnnligaQYgYLHdz6EsMtSaCdZUaLIimkKkaJjnlWp7lykP2lkLKnu
qaHeNpElvdQ67yRmm7oL0o/SXb9CUCKo5NJNYFyYAy69XcLay1zGYh40ZYPBW1I8azPfSVqbQqP6
tOc2cUYPc8tPWrs35GoO4uk/OVlE9h6VgDZ+n2LbvhuE0nRM7o4HtEnP0wccPEWluQFxF5kE7H1A
sK5Kui4+TCMmrPMI5V1suczBOvc4bcDefNOPZuUnV2KoWhDPius7cOJdGwIXTd4EX2eZaoiTjDxQ
BW8umFYBXUKnq/nRzG2BA0+NGZSqEza+m/Sk699i8CoRPZxNT3ZN+s1EBqHUKrZ3rgQK1N4all8K
yCQzZ5mtyMysl+kAtoKuzYqEICqBS37JtSs6dLL+3vjormeFEgHo+cMG62WQkN8s1aiyBNuPHEr7
E21jDlqPrlq0Md7EQfiISgy5zXqqyRBjDUaKa1On5MVf07P8MSfNKhoHt/G/n+uy+Vh0v2l4IBmH
WQPLh8hDIea1+qexIMQtCy2K+3d0EDfBujN9h4mrNehdkeVjFOlS1eiWtjBEgLXYuwYoKDGR7ifQ
f35CGWi6l/xP/cy9VG2B/L0Ldzo7K6zbvsifwFqxudx8UAnjGBZQG/udYbkR+RzSM3jXvDQSGHCp
tCnESsOwqjWo35FhzqWTBSPbVN3hAOHp615k/p4BPCvXMxoSeskT1hrtijlcZ0wTXxKh3luksxVF
SLJtV2kDzyXv/eZDZypK7Ctmn5TP8bRcBUJXq5xPc4STFHRxVh/q8cfd/dBSbwuti7Y3MExKNMTV
dxivogtxR5AQDyf4HCzaWKXSDo9JKJr0RI/n4zxCSrmHbfaqvrczoq766EXDrF7fuHx8kv3u52Et
AE+FutZK5y6yqy2tKscvqdtCzzLLd/RnSejpowkUuHjNelt9R6RRJn5oqg4VqHDoL2vT68iLwSPo
WqmfoXc3dSKUXHUJO25H2PxBsespVGe4SOncDCdXAznpLkRPcI8fdWuw0jTLPIGPxmYbG4MDlicK
BmhAn443je7FACDm/7PcJdp3Dw27QQYl084R6p2JIIAmnEyBDJyVC8dPO/cYsE0si9lBVb1dPFWu
ML1Saqgso7UttJzM2YIoAHNOjplLZ6HV0W4GS+yBfZoz4OHHojUxKrohcYEgwyJtuHIdaPOmVmjr
AKJ8+v7DsRxD3/JBn9+B0AJO9LpECOl+YBT1SBzb+cRQ7yMETqZjJNX0W/72ltOdhlEqPqCICC70
qOY2byAa+dp08Mokmsh1iYxWIasfJcXjMMkmp1h0UoDpbXr5SXbSTEYAg9x2424oOOONkyrS4j3o
JGy7WcHE/GUcR2kLxDdyzrY7h2S9c1sz3+55zLbI1n23Vb7UyrKBfQDLH3lU6toZs+PUSJo0mBVP
mUe7sfTpRgwtrK9ZP+thvkbpqjgJ7mHdy/Ix7FEgNrzPmFKzeHGN9wM+NTNAc5eEiKBZ0WoxHcyU
hi3dBfQvHMWSXbP8/LcLnGbwMiZs/SMrAsBtf7+vW/6/JtK+ZJtZHd3GcsjOhoX02ibOUfr+tkGg
AG8n8p4XrIBpzOa/KMGN7Tdar8r2Tv+T5cBG1/aNOxctVJDbbvbeHezJoY+nSLyKzvme9CM3zlHm
KSI7RnqO3nGpFwNDhNOiXhFfS61Cpt6SteOvDftt6TNPiiItA4qIPmcXge6I6P4S8QcQSREL7kEI
eHJ6LFXuKCpepyZE3Jn8Ut7RvZBYaAtSpiukkTyI7HBjGgEU/IGDoRo3aTyN0L+Qd2I85m1Tp+Gz
rGLlVm5oxjy0tjnaeqJ71CKVe/vdemSePBBsGRZ4LmfhgPErzDST5SRNO/Uvur0g6d+5CgbVgxZu
kOidqzPhdXa4noD8mBZuxygBH/V5R+gpxvoZdUv8ubMfXk/0L6kubLvp6ZReNjWo07eloXiMpnwV
TbDjL25KcfKLPf3e9Q7y6DG5rggMf/nhVCz1brLz3FtdPV1OiRhSzaRSaQJ5eDc7NFGbAgC0winA
LP7Zqdt0qd3w5VTCelh+sDaG6YuuUMZ369UoWHJV7p4pu1uGN7m8UVR5g+bVt4/SvOAZhohZzEjP
bR3iFC5BYDrNyL36OLbL2juqwew3U0keo/DsIrI7RSLSovzrD5vuiiBEJh7JctE0xwVyXJWXd1fu
muiJ4wnTGPgnwkpRqmsmOMNCy61uEGk2gjmgUrOvcezXcMJXpbIWh5qQcA3yr0LM2xX/46FhDARC
yApQxXVFxa80pFRSkuh+DIDZnkqRsjmPvBVGLkMQe/+z7m2XcnIWlSgyeqYF3KLnOUJM8Mq0iWyr
0VA56ooHs7I7FrU++Ey5JYpGkcGNn/NXovvEBLg86E5h3zkfQYS6pgmuctXALgGfuSI5LwMD4Coy
bmqPeq0nwkGu/Wb5gOtg23IrCp2C/0ksiFsPyMC7GnnwNj/8xMo0fOPZdWZdFmMnXL57/YEvFxPg
avSfa4YHwcfKq0Ppbabm6qkV36wrAIsQ4nWqSzbGP6NWLbSywmgGakFtUfeDfNcGsin8M3JDwj8z
yRwajLnv37XwTXWoFm//kMgVa1/e4/TkhTjtWw6oUHnCtCYUhVnFP6EzrtxEgNIWovab4CPSvp1h
dJHKMLincDMSn/Bw1SCfJnVOq2U8Oimu7ngJtR4qVvjnDNKrao8lnvudFlOQ1+ERmLbTU1mxr0IM
0pbi1vAnxekl17P1PJSIptbpFGEYY5Z2gjDsJvkS5di3lQOa+KD1lyl/w3qPbw05h6SEULV/XMdf
8rSo6qKrlqE/c7TwVTj7NWjxYw196/rbrSYnBjeFdBf95rdeaEieO5ca1tDQkF+Uc53/l8oa8mNh
jr8T0GvfMmi2bJEsdgXSdF9hScPkpXB7Hp4nTJOh0YUu2WDdSb9kespUb3ARj+ajGiSI0wlcUWQC
n24aKb62Ig0UT9J4TM+5mp95Tf8w7s24WU1MEea3Kvay8ynZ0rxkc25cN662Pt5h+iePxy9FLr8m
FMjmR1jWSBdxRv1xq08pxUL+Qp89hccpaZj+071XCW77YWsMW5mKBI0JYM3MZebN0JWuxxxm4NoO
zig/fvw2eR8b4I7IOasFfdUecAbnFKpv/3afSVvSkYIsRAK3qPAPH1uLJ23Gm1tJ8eYIzKJ4lNb9
nXCqAhVxp+Y4IQUQ9X9BXbuIPLbMoKRl8rKOx4sJ9UUJBKO9sTJimZMXlrkj1ltwbj0cokBHkgKx
qzfbY28ckfSd7WIK4zuzD+USNv1YM2VR3SLt0OBTYXQhBVLXBa6RgwAZCPQHwILoUmDJz6SuZ/RQ
zT1AKWudoB8B6zC3NdNVQs50tD1Y1bCERh2BVWGrpbFNmbQVDTgRUpvNPfkaQF2tdYMrIekF0dwA
bqaLTeAftd24Rke7O5ZME5TMLuJUJ8yOXHUn5w5CTcufIy8Crks0lbMs7jPVRH0Ft+vOvmdVs1xI
WUzb900GJm4F5hQ3GRNBAa7Xft5z9f16pRoYLFRCx5EHLqP7dSRCoORBObYoifeTtNxyXp+3P9hQ
tk0yw1MouZgmhdFT+FT1NRYFU3gvw5qi8rwFmdZTBvrFD0PT6IFKKyH6TuIx3SA7N+6FVWIgO6jl
z4zT2gC6tGIH2rWio7NWNn4lqAUxqla7ShjMsWw3t9sAcuKZP5BWXSWk596SMrnKqpyItnNBy63r
ve29MPm8Od9y0OWYolzjXpmztUnXD8tujyWJc9+2WWHJ64A9lU0rgMhtBf1g4XUvG+Zamcn1rtvw
G2EytzSHMYRGiLgU7Ed4N/cW+jWneGo/kF5Ly3/e4NR5i9Yvkvpwp1qbP/FB/qSDICA/9wWvXNVL
JuHZJUZ82WYTVgxrh4s63Uq9iURR+v49wzAbrV4Dlq4y4rFpE6D5ZradgGqPRYDxRmmvikpekT6J
6tf2DNLnJnO/O3CFK/exCAwANAkgJ/KEGPQvWcP0UlvO/ZeuaMTxhxlP9A4YbRlG47VnVApNgAsZ
rhnBq7X3Z0C5DDzuunnAw0y0HAaC5bGCz+xhEB3+nWfpKHnTx33GzkKnJQOrB3+TZF3R9uNF1U1g
RzL8zWvHlK7SHi4jCZbuYWiIdB57xu8+tl376T+sh8rP9QArpB1m0Pk1TKZ1IUjlYR0erISjSp3B
MMR6YgBRFHjI6oaCxSc3ydmIrL12wHWi/6RqKKcZ5h0LFpfT5oSFO4/8tzbzbpXiqdrw6EUKBlAX
HeEBTLlly3OFVvH/9/mj3FWZAn3kphBhgx5yS56sKoxTy0K3r+7dzp0NbFjKXep6OhnysHnbMefl
Tdu6RMCCRyv7s9j1g2t1cHlWC1CoCSAIUNQ7yPeFmtnoUtrhBIZU5aTClGU8O3+lYQb0zfoOnq5v
5vjHOVOXD45hj47Dwd69abRPAqdibOOZbqfDHClbS0ACV526jaWTzxlLudBozzw2TM4+4pWErPWs
AgpwTsk3y63IUc41crXZoRDiCW/UWmCsfZEzigTuertduCrcRUkniqw4ka2sIjCLtmSEdsToOwzl
TX0nxbOTc0YCkKf2+Bc9humoUQ2fiQ9mi3X52xyMQaKYE9s3fJnN2BpzVuocgVYjJBMuihSEFKaA
8kMDglmlSnFgF6/eLlnlbzlPADYdJTN4HvreVqbD1dYQjtU7JuJ3p2gfSfzNukNW/AfudpatgWMH
9+IFF9IO0ddLb4PrzKvgo7u0kbP94xN/FR2njmPS2pVThnWKoIATiCwA5G8/VQInBKoUxuxZ3jOW
so0s+7Mno3u2O7PEX/YIKJXooYiUaEeAj2ttpdPz4b5DMo3u68jbjJHgCA29w5PPcR9K1XPDY/M+
Yvmk2DgY4VmRd97Y7bnkmGYvsGYr9aHFiFoY9lCebaffPwSSzVFqNVcjNXO8yt8yudvTNw9WE8x2
B6KpUx3YrNwXETQQ/L7xLe4NuKi99fa9Nyaw+TY/V1u+iolrhfLvSuXqQOpiGUlk4ef+TAhguyMK
Cxq2JOv/XIUaDnT6gf7JNVHJYv++BqmEEpH2hy4cHVj51hd5zZhnTGeyn0QsA9lmaYpE+aJ0xF3v
pOrGCYEqgGAcdrWCUfGXmcE2sZEpfNE0FgkAKN5slf0r2i1xVVj4yI1HtfTAW/D9st3bw/Nd4Nzc
e0HjUBphe6rfpwN3vQ8uOl/6OZECnZsWeByFmIZb2hLH7PfWJEEJyVnGePJ+D6ZGbd7oEXGfvSGs
CXdxdIGT/vwtXjn9Bwc8ATZb2HaEV5fBpLvS3bFwmGcxSzd9fl6Zc+K5Tg8VQf1VJFpie6Cs2MXz
N/YpIKf9WpLSBFNalcO78Fb2pK5R5nlw65MDXNDaUJagBQCLCHgfsvQamQJh+DXlrXsjH/ws6lEF
kQp240rS5/OKxAG5QtB8R9A8JAc57CMOiZAdhCi735fJkxebQd8DAbSoCAGfdWNU2tCHAcI0AHYJ
pm3gJEdkay+EajrVOE+oMLTItYZrxJox6fYeeMaXEQacteh+c9anpunoHAekjqseXKDE58rZPA8L
TZckzXUZUXVdWaqyYweS5/et/t0GqVZ5mcwO+RcfyaD+vukmWWKNOAMTj/lKVgFzsZf/1GhDk0Bx
ABW9tzCxiguGN24ZoMLM3T6NRiwhqj9zL3BreadIOSQFn1bFa4k8y8PT+hXVO+gYrDwFm/u7Qb3r
0N8PVn/qKzrqeBzk+fde+jbSI/B4/Ju9vOrFYAs8pY9hkWQH2XWUdZRfwu63jEVgB+kSngmchv4a
5ZWJrOC6+9+GjBlbAV1XgY5bAS2sULHv4eija4vwFdxLBYaCG1r5zGbDQwXwM22YEe7b0FVN5tiB
z4H6KoCl7O2ckT9LhOEznwdcsb+YUT11o66FwPHjL1191u0x+7DCmXHeTbWuLGlkgVS4vO4zwF9r
yYl6STwQFkUf+C05YCA8c02qi9dX+mpDOfy5MWKcmlRgqSRFVAlqPZm/NQhuaxEcpL0qkQT31vol
s0sg7lyp16i51GRwPlbP5pWK0s90+lhIqYFh3o7f6722o+MabjgBfSqpsqIDt/7XoBVANlxlPUtR
2OGEdw4Om03zT0uTywu5YOLlbSnQopbGgYPEXVa83x6M2GoVaZaa0/crTy4uYLeoheYF/hCkmcSI
dRkqFAxEctugfqLkGgu90Im0TqaOlvIoWP/2cyb7BoKElG1J81kkZ0339MZ3zPBNqE+eW2vNdJto
hZPi4rzrKRK9c05+6moZxnb+bqtjJot6yrYhgGSI/qjhr9dG/5nP0lJ84N2LfdD1lLttjznLKhcd
UnXfnfM1a11FT32aZWcme/n9hrtrI5oY24qDrhBb8LzknfyaDuRflherAwdSZK9uOBURbnkXYVYr
v3c2cPxBBZeTEi0xBrywfZsUKhyx9gb9EHCtgFNi0xXOwN52/0eit7wk/+JX+xigIlY976Jh153F
PpYI+wzuXd+jbxrVBtbLExqHyXmS/VhtDmYuUKl4iLMNJY4N+2H99z+Scq5MoQKSTLQoltAoChux
89eNwiQf3xflNU5y/6ayW+hHOVDkqMPcgU2esgUMci/PVh5o+nE6PWG5Qo5IZxNuPa7p70OlSNlr
I31wx8K3Fcekgt9TUqpljgqVF9tpx0ftDRHHLfBJDqe2gZkPXOCGbOSfvfmYrxd3RsQR4TTErTK3
oBl4oEKSrmb9EYtm96hkJZLJNkb8rKbH9REgnvHZxlXPHD4zJm34VdxUbayr8KtdBtpj48TH1kbE
s1SNYD6YJ6kVeH92f1p+w8VOGUBnAV7nu2CtdSVibE0gEowcCjR9JET+I2oaHKpzaMDAIRXgmGX+
cM/3BfXEWTJK5msTf04U2o3Hd6vRAb39V77P/9U+XJwlGx4gyFEbqzXxDo2SbfMtA1Bq2egtIPib
6gRu97AW756+lYeFlvmc8uR5Y56oC7wvbmft0MFwPMsoBJnUGQtewdvnlt7eocjGmDu8Hjh2/qOB
tWqYUECGv+21MlUOqNgR5+rIHJYVJrhSDaJ1cjl0ihI41PeVvaW4R+NZ8tYC5sFapLkW//eTye6n
nWGCoEr2WFuMBOUyOGXKhFwkDeTRTP0mjfHdLCZuQbFhaJLYRbh81OhA4gh5O0MlYyPKRVaAsxsr
72Xp4UFC+FYmZlWT807XUbQ49trSULR/Q2VrPTRfViN2gd517N+rm+uspcbYhyV9tYEVOFcXnJ9F
XBaMV3yiejENqeyKL5F/4Qz+A+CzUxILgRuQI4CAfX/dQzdk7bChE6OE4BwzQRdtHuLlaKKmOfNR
YZTIiwnw9AjCjgBN1DGSVK9sosmpfsjZ3xedKYNaLMlbCOfxJF5cN8mGIRQbeF9+/bmaHQZp4aP1
h/vnYnqO4nMmYMCFlgIwSD/ekQM4/cwj24Wa9RsScdNoX5N51k1YPbQgKuP/ezAK9lekYogt8rDr
imd48c/QIGnctmI1jLnWVTsknjbNWNgpMabwp2a7y7qT6zjCIPeFcEMkr5QyDZhzQAapUJsXdBT/
c4bQXQ4Y2bPfE2pzmCe039IZFjx5lF4FWefA49G2SBsnN6eFn2HxxRnOxXWPISsx2tXGS05KAPQo
blTQ42YhiJaMUYWwBOXhBHNRSZ1CnrBspPhsGNJyHuF3RbsMCvDD2XIX/gwguwaAsk9pt55p7ltq
wAOLeBUlq47+WAGykNUsYPUxFo7Pcy1NGLpsZOJAnBEOevtH7pFo050vkxGci7HDtHm/D1xopXKq
d0EhdCWYMXiEAhME1UAHl/Ua2b7oGsAmr7H0Pwr7p19Z3WYuq4NiHrhe5Z4bsnHWfl2A9qrnxvOS
5w6Ce+FCBdT6YXOyVgDHDAo7CQ/BIXRxBAu2SGFZ4OsVRD/76L1VCN7iB9NumocXnWXC8sOwg77c
NQbZNKvoEBZud72dpEBpHSXjIqMopxtFbeXwZjg57U0pBVeapQQnwnlDZUr8eokv4OcSBT4QQ3vW
miqWPN0Y1kfRSdoC6LZn2p4QfsLVrIoIy+FYeZppGW6VwIjB+RuOvc9hNOCrea9Nq2Qo7kMWR5xF
uBZFVTlseInF06s0YBW9lvyiFEs0p8hWFhowkj+C8ruKNvX3+HwQDTYVvB9yZI92B8ILEFOHpcWC
vZrk1HWU+xekziQjzQkWw0NjGZqqq/LI8M5ot+JPBQl1OZBw4ugPeUwExrD7ujNuLYlWPkqpXhSp
MtbimR3cyloOFrLb64Y+XiAVerWIcGv5XyJkUvG3tVImBHp6Kg8L9H6THL2v1nnE37OXalaFkzi5
QKzFUlxCg6QYjvdDwcpSQI3jXqk6iy7UHFjPX0vuBR0CK7UBgyj1cnZOsbkVIQkw1g7TtIVJrmAz
56mP8Wi7DLjeBPiZn0GNq6NiLzB5GlDM9KdrXoTUW+TVSFUmGzSV/eUFoiSPTsGASDFzCUcZ+joQ
FZ+3Yr83RKqcVCrR9kgQYDHp4MIitkiSHwhsDT45xHPddvibRzlFLj1qw2J2jJvfqUTxkr6eeEJ5
Xd5O6w/0Z/Yj7s2KjIkDlhKZqr5ZzcmrSYErFTWSclktBIWWJUXRB8ZRVmc/tS6/rPxVE8iPIDiK
3kOzecZOVPVd3jexA4L6ORtehDU3uI/Sx8ANmFR6lbmDtpwdVpTGoj1MYhzgGdQ9EJ1GbfiMgHJ5
lojp0MVihLWFOZ9t3+mCG8NamoJG+ZvhDNr4eVUMaVGG1GPUNjLRYoBsMxQwz+23eyrWTpCemSIc
O4vMd7pghOb7+P0qeqB2RKGq8dMdmH2no1cFfZDxuA7Ch+wVv4VLNNWfuhrPWw/kK1DVKBb3XtU6
q+RwckUUHHgGB1n/vImwfE3q89eNFD61RChTabXYbw9QD9eOvb96gK1kWYTQtbeAMdTj6TFcwvdP
2ApYTSCB5tsJ1x4yFp3VB6s6+Dw8ay5MAKVc/Xdm2Iqm/EELzkNUIkLQvK2DXAam4pspwO6kF6ca
RZnJYIKZ84DTmjHvn9Nkm0EhDF/yB0EaxN5Nv1JRXbmUlsuHYqyOGH/JCEHhykU/urStYMYUT8Mw
8C351lR55J5vlu3F//Mbq+EeoyfvyZDgprkttCifJAH7aN+MK6U6srguA1NTgD5pgM5jtmA630zj
MMLCCxjNrBiMOC/Kig4hHcIEAWcC+Ayo6HDvcpKurqiwQZixH7ETQW8c7hUsvoolQqSiQvqNQR/L
/aGlqxaTSX36w5ibnLriFy1uOifYGQO8L614LQoGJ69LnVeenwYbWQfU+xPQE+bSkSWcv0WVgRzl
R4JB70pEzYC2NYULhKckTicmr0M/dpvMMLZSeAnGPynQNvHKW9Vxerqkz+CVUOXOg3EP+IQCPYf8
A/iMQF9GsZa4hTMtWXE5lJPUbPqlMVF2Ri1/DTHN8WfUx3Uutn+K7YtAtBToYL7wJX30nUONigBb
XMWsS4x+pY3imS8Afh7umiiop47JVijYQwoPnCCMNlKip0BJywKUs74zPz2PeKkjwAygNDCfqvRs
uvNEkfNLLfERgp8s3J7MCOqd590ke/x1WFtEzSPFGgHHfJpQeE9VWPAqU8Zgr5aZLIa2Ajomafua
jvcNFu10MMJsKXF+staBK0ZlqoIFLAR6IEFI/cAfD4s3audCYfG3RQTLaEIr0PDXD44HwWK3qamU
SstFk6eKUzpayLg6LIissg99LKWjGdlOvvs/BwCICMcreGlDzNbA+nUVp4U8Q0f6ZFEwoViQgr/W
PHtx1/LH/JMgucFsCFsQQP2yczImFEMwCimQk9ST+lyrg4qhNjx4ijcxOqfE4TOwpjv9/S5BIjT6
DQOpUncIrPehmk++TeCAyuD84RclvLJiWSj3YyA4cp2hIY6n3LlZa4mxrTuVUzP6VgaicCoGPLLJ
bCD77gMoIMuzy3Fme5fhMdUpZxS6WGlfzPU46ZKauMRbuUwg8FADir18JoBqB6CGnsAFDiS41VSq
P86ciwZ/buEId3L1POZ4oj5z89Zi9zBqEEIn03nifOCifPdmlaNlgYiVXUo/grFeblMdJYN3ieHd
UqcBOaDhQhOiOj17GbI5nfZx9J2wFZ2fqDVJOr3ntb9c+Ogp/rJ3nJn6vr2IgikZSitjMGNsIhN+
7GwNcrGZ++JCAPjgVLnXcv1Q68CztpLP/nMJ0YlydszpU+S7kou6sqwfOs9tFzoTyfA1MfZ3hkN+
ewtHDbueUk4pV1xeNkDm1LfTKknc74nsGXy/c7jsrSTe1yjrz2Z6UHrpCESeJcKxyf2wesLxKc8X
xyd5hf5onNDL9E3+mfWFDnuzycgigy7blxfPtP0pF9oE37yW9BOR65xHsFQC7KZxZPZYyGjqGceS
TUYobr8z5Sfw66PytR4FFSjeeH5X3rDqSjIVazjKx8ZWfxMBc77QzYTaEOPGVGknk47b6rHd3DXY
sokqCg3pGTdixRoOOYkoGS/Ylg73IIvRgxjXfyIPRyklYo9TlbL7wge99fDj5pV3fHkSAI5dXYYW
B1E3ytxFquMNBC1ip7pMOAxZiFfPNTL0xvsU40Wh/6AZ9TLDWbgfdZSfGAIdXxtNfv9sjcBvgIn1
28gDw0Q1HV22Fwc6dLxBL6+NeoeBlSrfXsB4i7SKATYxoffVIo9j3j8rG3iLbWX2eRr/pyvypRPR
jpiNMoGIeoxS+K7KrV3BtlS+cHtrLQ7BST9pwnXpAbxg7djXDppylnvdM73zQ/7TpB7+4frDrJnO
Gjy71cQx7RWMaoU5Cla8VNdsPuaSAKOEScMN4pvYOwXq6/KzAMxkLyb8SNi48F8CnEKgELGBRUKZ
PB8mZrP+HojLs5HF0ouGY5OqsCEJuDWPTYAlYHzIzGgOsnzFMTjOCDJapV80cBlVlR+7l52bMEy9
mxHvzz6u4OcV0jhrwTiZKde0Xi2Hs0Y9XEmPEbqAOaOWI+GJR58cXPIRKEaL9P32wVwwkUQ3g4Tw
1OEBiWt2ZX+MlJ5i4GwcXIFZLyPUctLXUpxmoiyfmdG2RKdaGrTm/NK2Gx0mRc7gTIvHB0jRv6Ua
lSIB6PsEIg4W+Fw2pMNNYBzAt46dTH0ECISiZ/aBacs2Wvxn1T3N9Rt5rafvijiXcMb+97xOm822
kaKMynuRikvbchVbk9DZFSt7HEUt19AUxlJy6TZPlYDZzxcULqYEiq9BvQt5XRghhWOMvAYKlQoK
25R8shK2wumAolG0qiSasePd4zFMgTQUbDUqGDxBOc2lO44c7Fsl6e9vXvpds9HkdJYdkwSIPLzx
UErkdRjKlYR8IVJ0a4Jli2e6s4q93nJ4VCpoZTmhJGzNpVHv5smQtiV/LxviAhspg1370Ey5uO+W
uEH5rNcu2OX//hx+rjRN0KXkYuoz+XZZ4w8hpXpcLY8imLmkyJ43c/j2+OGiUriGzb64YqVu/4es
RN/XpWQ00vsy0aNrarQ0XgGKbYNLw3pWsbNiH0ZWgP9zRMliq/ouNU7pcsaiA5hVl9riPQA4uTLF
RyZeRgy+CQSzO3SixHG7ezVFNi1urgxF2BfEJnRxhPEL3NcsPTdPpgU6SkiJee5iDh97OXfj6xfl
2ZwTWx/gA8HKKmRiqCjKVXsgRNvOcDEI1gc2eZrpvcCcilAZpHBVR07980tTxwu65GIoI+D05cdg
S/j5AEwHs0WkIZ1bP530sN0jns4GcPzkCLnYkDEAEzN0hf93u7pKPiZI8OA4BtLfAH1HUh0jhNN/
gaLP9Mf49jCEGByPOBysdYl+K0EEPu9ukaJl9b8Z7pyPv7y0P9hlQwWWrU7FY6Bq2d8CuzoZHATR
n50Xj+UZzV8i14wCAuf/se4l+cKjhampiiFky8OjmtZdRhQ8iNp3JVJ+ZyRqhxWiBNUmpO7fSSsm
ndLshGAI2D5cnGoU4n8PdMwhub1NimkNLpvA69+8NYzKCNYGorMpX9KrMvqZgq80c7defL4+mmFr
WrVgOPmUYu3DBO109YA0rnmRqKXpdHc8bZte+OrlSAyu2SgL0wnbxfHOu0y7dIyBmHi6qNF8PInV
aW+oP0DVmsdpBy6jmBwhUFv/3rCRYaK8MBOaHLy1H2/z/KO5Ef/KrUW48nmqWrY6Cq+DiuswiVkC
uugzV2k7BvhlmBhYS7dz4FPO81imNRjlnsy7k7rryBGPPtuVDQa2F2I5cvpoaWue+y9HHfWSr/Em
JS+stzP6isp4MiFgZCFCIuJjNrxAHiXqZFhTt1adbvIZdfslHJKOja3yVJDU4xZnM7DdQuDwT3kN
dVlvmz04umdLt7gCxNq4ekitlevrxGFzg2Un4FkwPAJN3VP/WN0kqAFgurdb+hBwJ6Wk86S42d80
AHYpQGUAyfmsK3+N0b9kd7azrdzdV795iMx7uJeBweLqR2n2qocG10pbu1XkFQMv8/GAXAf05hg1
hk+fFayntxxnhrQ79Oki89XpyXhLEACK8FNZ6AGT9utZqjn2aO9lLOfLHCTaP6X11toeqsb7q4Sc
iNugonosAceW6FLpXNHtY+okgDgTpCUgMtf92f5vspTqwYcMCPXhgdr/PkyMQCSdVmKX2K5EDMlK
niVcPo4l8pUq7U4P86a0wLqpYpfYmwhQ5S9b6D8dWv3lI0EkjWG4cBnyfT2iqP8H3JZ38hGcHjrt
QmYhcm9IuKSYVb8R0WA7jxakCfT9RQ7xR+SSffyEtPDNrvj7JDD4RG91cExX2AuBVnBSu7qcZnZq
ilr27WUDfROi2mAcDBQgLJjoV8PfVa1grNqny3Nf0yhnfVWdOIb6Ezh6JGA7AKZ5DBK+T2bNjssd
klPk1ZKRiULgNH/fQ1F2zhS1I/O20hUEs99kmaa+Bs5ruVVLLp6S0h8Kgs5cAvgZHzIUclbl3giB
q8P/27Zyee/ywSNZr/TuVj33C8WvNkHayqd1dd2RuJH1Xzhvq0ppQTYHBzXkePfym5lmoZfnU1pc
hZOJZy+zVBofkQtGC0R4v+RBIcLLB+1LbY8jOAAiJ6YGibsA2hhzTHjkreBh/HlTdM8cuoqnyDgw
Kt99Zs6IHNAjXELkYwLh0hepdAGHFaToAg6Z+d5o6CV+9caYtX5lfbhFREvIZPebK6r6x3EuFtvq
UufK076eWu1VrUXlSiBJO5hx4tHLqY60r1NkJIgqiJdI5LzBfKlmArJJQJ0DjwlUyILM11qu4HiL
9jG1RSe/4lEhVSCyJ4JmkxweKldJN+zrflXOMsibZmTeRSbDImZwkvU2U5IBgQ8oY4lxU/Hc8JkV
gShi0wMNlI/CWqzCCEacdGNFpTaEAMwSWd/nzB3ydQl+F2mBK9KPNSaXdAbzAvUTDfecNWqsCMaP
LwfuH2uhwbrN3prOGVSBuLmjnwaqguClxO+HXRUrnzNXkD/Z18hiUBdCc58RgVH1H+5DPL+d6lWv
KVp7dRUPMc9xG3Bn7BUonniY2FI94quSIbgChX0sk3eAhcpZu2oc0RtJJOXIjNLOGIikooiOl+n+
lY2ea3S/BdUuxfhcwyKIE0p46OyMniB0OxSggLAXoYYyjFth0wf7a0e2zP57kTJ/iqGSrxxHHddn
nAt3pw2JBwq9qDeINed2c8fHHB85A5RrWXXfJinWuV6S7igaDHnG/4qD3cO/Zj6yyRqFvsIOp1QE
IzFw33hp4pb4i8M0W717QaOOWdU4d5iiYJWp86SbALW4A3R8wSdkQ6XGiz669jnF+aMkU8OBPHM6
Nxs53PAcLNSWd/aeRh5aAjLksT/WC238tvkVz32xJlvHFFV1H8Yn/Ewq73RRaAoV9SZjddOi8AYB
6YNQFZEYtcbqmOX0uERnNijhBBiNrxjEWbxEy3xawBcN8DVsa/q2z1qiEMuMPf/cLp7Pkjye/CQ2
O6daFRdmY6RFqOrLFVxrQplI5lFE2Um0FVinN4FByRICYn2P94hq5lro9rWdSC4NJ6lsjp5Qa0qh
ADRW/hYgPdGDT+AD0qDk+x8oIakz1l1DVQRzQFN2Y4hy/1lhjhK6Sz4shGYOzY+T2l620pf0xzlZ
DVnFfDYp79E/57uXMg5SDGUemJhHaT2iJOp5CckZORv5ge8Hh+AqBFYQToukztivnaLeak4AXoqw
RIOoGurqKo+GxaBOetkqEXKA0Xnl5n2ZGaZygBg4I1U3EkCWvh7xM3fH3Q77XNkyDEFBv8YW1BhM
QC4t/vIOp+Q5EAepyXZAarqZOf+Tngc/dx7iT+YGE2ekHGePgJzIet1qBmADr+sruNDpaBcDf1YV
mz1vbDguLV+kHspAl0p/wbv4Y9inD9IgLc74y+43DcLKJquBMXD5HzN8fpeyFvY9cItEWg88Qqxq
wX3uBB5nbIRq9b5VCFsLEzrcex6e3dsAt4YROpxS9NTcMTm8smTFgDd7z6vuapSlFd4jdKtmA+95
urKhyiqAIpK8j4wRRMH9L8u27OczS6jN6WQEW1FVU/3eY5gzT9x0hFhW728GyREo+B2MErhpAEJr
N7DMQ3zXTNLDEFsdfnGyAlK7R9mpzTjCcHcHSXLaMJqbPOAhc+/IozR7+5QUmCRHNsGv6ZAhrka9
cXgLPNNHfQsciYOUshBtnVirXGZ2ynppvPkPmB7lRbws1mOFTfioZsDQovciM4PHSeFIBVORz7Rv
vn4Mc9+pIfD+8FdKJUbKi8tne7sMlIu/w6fFdvCcp2bKYHE+1XlCafRMt0aCwoA7r8m4guVjWbLf
n2NK4lRLhhM6JdOFXTZLSXXVD/IfrxXbBLq1gSbZ9AVZGDrRRPouyzSgSCZgEmJe47ouSxEmcQzi
e/VPDbppC3WVlVkY4uUP/1/NoPf0y6CthLoCaTztpkr+JvWKps8EghKbrkkmk/nKZndwdnYASMnR
415Lj8hBC0NVfJpeSk/91VBA192Av/sj6LCaZFE3n3vv1K7xSPzGNum5R+44yrUugLYDrUj8zivs
nVS3I8Lzkyozpwo0c4IOJATSfD3htO1318/0bTHwW5ofnZegKQ/6M8OJCjS+T0tZZfkfcegIV9f6
z/u/biL0CQMwW5OSV9tYzxAoPqcxSwoCIafm4ZwI1hRWHMhpAjafxx6Vm6/OTGdM9HuvqMYOBQhs
/QPFIMC9pDy93xRf4A7iwEcEHUVYghmpNOp2guscBsFpz02j+hOl2LY/tgB69F5fK1Y7tVxexX8v
pyjuSWYzkHZtoN76k1c10jBc0cNkSifMYgA2dEkXDMd3lAqVneLqrfioc+X/dkCHWFvbnKFK9bM+
QRnnEuI01sDr1xgHlSCllz+Cm8gv2oI3Jx+95K91AErDHLXUYGtBAQCXaBVhG5FbGrmVigQPnbgC
L6RqLU+3DDgD7UJDCsxlpH0ycMNbDT65ZcHM9dX+p8tGjDJIbISbmzeBkjVeKGPDepSMiq08aUAp
lLrBVol1sRXRSZhcxAouE0WJDiFk4OJK9VM4iaJk1f0V2baGnlJJ3fN6KqF8lM934cHQ3ClzkeYj
2HxDO/rTa3TIh98fJicrpjr1nxRkZMhRyK8Xkb42wo7WkO7tQ3QIaYhOWbXSeZKTY5Bxt462WDh5
xWtDOoSt+vHRJWIM8Lobg9CXbx1j8a+OX9Qheur45PjcLruiCxFr3vs/IP7UWh+UXn7sbuviXD4p
LV4ohoQlr7ng1Z4uMS5/kevURC/8QDu9R89VilhjJ6LbT4ZSMxP1Y6nF0tsarhJ7/0lVy/tKp1ic
JPxXHjMK4zpMgXSBYa8PsVIPpeQ6KYHfXoJggLjw94yOvX2Ob3PAH3KeLiWarFOo0uwNiknr0gRC
5QeyGf5bIjVDSggin2+N+O6lBE62V25BCE9TQskssT7+TR3qcaVvpOGOJzULK6OZykcp8y4RmAfj
YJIeUetmV8h6OsZFAmogQKws4lBtxJiJ2fnN9cgxhKiNRQQtsUcBlXOAVXN/xfInAnWZl/0F80Ue
+3xMOaOugoYpqvRcuxKOu5p11V8AJyAhjWihXWobEGmfwZ2XMZYGkXAbepqvKwOr+VsaCvPHbpjW
4490q47f8RkON1oFqFP1UhORuzBk53XO6iC6eLEvQjo5c3SCKMEEIZraHN37lo4o0yaFaabQHikY
qYcPb6eykrcEqb/YplbISoDrdcgnQmjKuht7aKg2aRDQ9oVIFTGmO2hDFK4pjrY5j8KZZL2uqRxs
sXxh9loIjE2gFLoaSHWaKENbgiOTjE0YBYP/edf2PgRjYKeJD2I7cGjLB591vXA+qhvJFD0aVAVi
Jly5U6IgkkwI0E7zNIRGpL6AcQUyKDALFA0ng1e5YJPuSxJtgPtzkzYJcnkkl1ffk1TrD/cnawFL
b5mLtTat2zKGD5ILnuR0aLdy7VMbCoocnjBTJJpU7ESjMwxHpYtQW9wG7YIiBtz9XRDu9KpW/q6Z
BivEQVJaUz/gVOcTHX7DP4VbZBOfI18wt28YCbFTKDUA0R2z7H2MaYcU4PFvmWlGJjgbi5i4Zszj
BUW8qoh6OHbkunTHKoArQNJiVqh7HKaUpaGZg7ha4NrFkXHXIEGphp+EWoc0As9uf3iv5lnW01Qb
o2B0ZNOGfNhnbwW6hNhcUds7zlXGi+1/CTn6EYqrTuDkgvA8ytBAErr73cKITHpMCdkBNeZGhz4e
UrdUaQQptrzJbNuEP6mYQLPhiVIP26ka169qM2XO/RkUlV0Q8AKYZCxY+Wn7FNPCnv9xt+5o+1Fy
tI8uQnjMvkIoBGLPyEafLWeMK5ppnMi7mN5iftzfWm1pT5inrwpHwGUpIQ5e0GXw7hxi2Ofg0htM
lQ7jONDtWi1TnRloqZ0tt/76tMdd4h1ylBbaLsnvaYnW3nQunyhXM0/Ri1589t/D+AWALhY8k8Gn
kGG4V5F8hSGaerRq765k1A7++k2h9elT7wcK3L3UpNG9iKCDpGyEJBeeCpOMdy5wnzi8aDEJ5k6d
1IR96vZRDAjMcUneNkRZpgk0iMQhYPhbI0ho12UuPAsp8TxIzl/9lHJN8rpmT46lqNNP9uJg4C4Z
HDfnklyuaLYL69aTN8rIwfOmdnI52vXg5u3pMXYrpzwpGM/m4VkGdvb3dWZoWPgBJ+IIvkIV+U4J
uFArINWi3krhuS3IQjEd70i7/uPuz5l3hL1K35mJL6845RiPW/ExLKCkqz1GBALmVSmCv4mbtXFk
N1qCjBjIbUU4tTElGuCxJ5xmFix/TunEfOnHSWQ4H8Ip3BAnzPeUCPpDBE9t1jm1Er0Xw/6bYhgL
3ceb+SQ5tjG1ejNtyAAtpvKfqDbhQVqC/CvmxaGVnxZBbrb3EVPPUzxUolSNfUwdqV8T/cS1gYl6
YHnSyaWdgunVvBn2YHH+EM/Z/lEZW8ukoqR9Ukx2xTS+4OX6Nu69t3mLOnTjXzDpt/dOJmXf3EIW
ubwrDXEm7teFYrc9fWoHTTUMpHPuHrq1wEkYLgUV/IlMDsr3Ff7cR79ywK/6ysdrI7fbi3hq57vc
bqvYYhQsRbpOLyt55yJcye97uaDtVxtQ/X+xq6ul8IxPvJmOvlnXmQXBCWgtOQ8/en3D2bCyFOUA
Z7QNTeDrbyH+mpziMU3yDy3YGpSgeIwHEF2L31OSAJW//qp6SytJVWjGu2FK3JDfDUv2LNOmU0zK
IizYmtGuBp0ALcyxqhnDg3g8reHaulJ4FpvPrZTPgIxRBuW9GITyhSYXfZucyXiQUn+tTbmhKSex
kpnLtc1y6PKRUhfCjcR13B/gPt6kvQLaXxsR0dJJg4B78GghlwnmAwqSKB0dT7ern0JFEEVht9f4
11tjjP4svQv5kr+81PAoXgUJ0Sy1obZ2E7YwOoNO1OMDyLROLjs0ZqXuzNcD1dxTnh+n6+tYIEuK
zvgeGOjVmBBT6T6l9NBu5iheZljds8+Wc7Wz1G6ROUDJT2y4VJ87Y/6mVnJX3FKWQK4mmDU5pq5Y
dSlPK+Lwy5Cu/netydStqH5qv94oKCRic1ScMBLlB1aJEHDmy8UBbpIWl8zuE/4FSayeXFRFXTC0
u9hxJOTWiaqBJjGKOKhtdB18t7w9UsifoPFQBoXCAjkVy/eEXAK4k5B9wg7pot81lBGN3xkBE+v1
ySRzW+1W1DJYApRjAMi//CpaCyD6FQs62AXKXLOu6KDGli8nnWxxRwqsSWBUfau1LCb/VN0k3CRK
MSMF+6eavQ2QqucIpF3uz+W912sRdZ55tgRDhdXYm/EjySvNtOe7MDvKJ9C9+U0kkbpgxsQZ9ReB
HZdeXGVzliNbBP9qBNB9gNIZbV+AdONppW8t3vO7/l+hU/U0idQF9L129Eqqmy+CldFt/3V+DcZa
K1rG0xqWHEI9oUpjamkyYcPN/GiAABKSUpULV3tVDFE9sp2CIBCv1pkbdY2owUj3FpKq+bIRGP/f
iLalvueZrh8EahmEPUhfaw+uJ/TwXHElT+MmAU/76iWgDstP8uJu2WVMURZ2ok/Tleyldn2PHBsB
XhxNL8HbZcFPwnES9JH/8QdlQaf2upLa6uw/DK5E/x112qgEsjPGjpM5dHZ+N0QsmbEITID81KOH
WSKJEed/+674W1Cg+GxgMxSgyPR3xzcP+kQ85/G8QYlOT2P7aXb2wlqNNITX3Q7baLijYqNq+U2N
s3DqkrANwkUh4dwyyY94R+VUtYkWc2HOPMWy/94MjFXNFNByPlYa1bbOo4gWzTjNRZ/YO5/jN5gt
0cuwU5VHQO0/o/HPQ4yO8LZAEOQhYfoxbLxpfDqnjR9zAqqQoZrDyWHKLuGc4JzfWmBwYM3SS+i2
nGCiILSET/ewMcxtNwEnRp6lbD8so3MVv6AHNiTpm5Tm4jBZlNhR+sJdYQb8v0PkgmwLkSnrngt+
7134UN38fHpUvx2yBN4I7l9oblHXWjkNjwanaIoZ+8etmJzd/QUviMdcDlM1G0zL2pvp+ZGDDdH6
vr0TqKXjmneQs4fD8ogoeTjPrldFoUhBUzg5uLmNxEeESUJALm5dsWUwl2+LBZv6Om+wgBW2U+6b
Fc47htiRxlurmmApfHbbaqyy80n2rsQVaXGa0HVOd5UpdJo6me55oMkWn8vo57qwMh0mRvA2k39S
4X0pK+Rf6drGDIdak5TP17QQvFs+R/+pNQDa1UKR3LHqzN0gfJeclaDfIcDn6cNDnvQw8pBgCMoR
6EohT3Yf6zKcxKCzhI/PYQtbzpIf07fvP4qiI8XeoHo8bzG2El+PSA9/bWtI7RtbGlAeeJuyEwN2
DTMWRx6L2yF0uU4b5pxKgtFvGrC8ReSYSNytABC+zgdk2p43kveojv/oPxroMyMkOxB2NyQKF1EG
TBEMA2nYDjenglUUjLgjSJi3+H9Lgnz3B3gnRNy38w37f0qyx7EpRxWlBOPOov9V9+6mKuvf3Izb
qU8MAK27ddgeRx0FEyFNuU8fvj1BLnuafSyBg2P/Newc5YTy3CqtuZQPFjrLDcykZA32N3dKyDc/
R/Ruv6b7iaiK/qeAOTMu5PJMJXpWriEWcCzPzyy5sh1Qi7W8oILfRHuzi5cJm6D9hQUu8JokR27k
p3mpoTO2QIUs1JUzxObHik65WWKquafXx8FJ75wJBTm6PARjnOh8F5rNTAzqw2cWE/2eDp7E+gix
G7BoxWA0K0G/5X9QmkTmEa6ssKAM81NlTgFzgTE0d9tFCAqUp9vtIRGOfK8MCgAkcJIQIj+TqWOQ
XGUEids1S03g7+ha2Qf4ptsB71M/+7qxX2f3ToWVQm0b/0wrkOXBwQZmuiWfzN7Yleo/Vj+gF31Z
FXztUj0Wa09Y/m7nH8plImLvJALZoPfnEXe+gJbLhViKhZWqtNICnZJGr9Em8J1ls52mce4uQjgv
ZhbuHpEB+wbGlZLXuMBs0xGqxaxALKbj2eAOB2Z9mKH9NCkR4ke4x7+74MTsNQt6zQoW4v++Uywn
wwh6P0Wfbx0BDsM2JMxQUhaf+6i0YHiKymYCZ1ksPzGhKLWlrxe8FQ1LFd35uZaxliPtGkveL/zs
5gCGuL9V4Y+01rz1pXVspUdSYz1GZpO+H+CESRxN6OzfKjHYHK1xgHZaBycEUryKRLpBxDWgsguU
sL8PiGVHG1O/v7S3Bx5F/G8bt8Qy2ck5qhHJqoP9uGS4ujcpOiKtdkHQpKCOswUPpIJKZ8DUjwyW
m8RD9H6c6a2hQQ/kban3WcuUK+5Wn4JKyIHDzqQQF0bxmVE4LhsefOAsbyFXYs4vSdEMPxTmv8QO
VRwK9F7hk75PPa8ByJrNddS19nNz5aa1d4DHdywaLLxnBMX0bQYSrgg8hcqeRNzfKWVhCg7IoZeR
aOWEn0XFt9LLmtibq/ZzV0wGi7VppA94iRXbS6yUGvBZ3AuketMZkTFdnBPWGQdV4X/kyz63sdSt
6hAHnS4jOyOxtOf1Mo+n/I/pqWj2HWbO8MjbTh0qE712JlUZqyiynPoM7N9JDrrr/7pVMXnaOVGK
9ZkpT5BlQ3xmvDVpEg+kL52dLYvlYyin0So6mcI8ZdDW250qqAgvZOBYOzuY1MKQTfcMBs2ZPJAN
LWx2PO7fHsId2wkHXm7g7geTHPufbbHCXtpe/+QA7Ab5hxCI+u2vkQla/P/2ML3917tsXLuEGq8U
0nQ6Z9UDI8HTcll+bemBJA0jjX3mDTiEWfT55yN72qHcrYmuNi7vMDyIRAx4NegrMvvJV/8EuhSK
dYZOe0lUH8kbg7sxoyQFA5aJHjqgr3ykb+/LfpMedGbyTTFwSUOPAbRENF5IOppVnPuG6GGIsPEs
s4uA8srBAZ5U4Dy+QjGY0xeFDlXth+4cdoGgJ+oU9Hb/lBPjpHV1j7idgyVr3+7+ID63r82Bq/9l
KdkaGLk6nEyhvJ+y3sP0onOT72yuRMigiE5AmxLEYynw5kQgFzALj5KN5UJXHdz2MCkND0sHwwbH
zPcURPRcuDmRbP5B8FCIYJ/Dv9a2IR3gXRk80M1jxLehlRe2OqNui4yOLNhfa5xAqdOoyF5w402c
TJYXffaQKiaCOQp6+sXCSq6Qi/O/BxFLp9Ba4BbmgX4Antd1JNCAoj9T1Z48jjL34f2q1qTjCUy1
9zx9X+0AEMWcQoCsTP3LGzLrUf/07R74H7Vonk8dxvCMv6+6o1cQ8th1g1Yd16tk4qHiMN4T9Ujs
YeUsnZuK9otnsIWXyOdMyOCD+1jtvIhAjshHMuOVYEPD0Kf5vx/Fne4R0zCqmkpOWfN0lvaI+O+A
JmyiRiEfR5K06cYzUR5Hv2EdBn9Q6NrMbTAQqShed7d4cX9q5H6g55wP9yEKeaznkPhRb9ZDIQdW
2mF/lHnTjKz/iDY1I00r5ZPQohNKZwN7ilLf3dm1sAP9QecxQ/RJXkn5XDr1XJiL9rWsn1mMvWBH
t990/y8zZf1nzh/lUFzjv5vWJ5FzDvRU7B5Jz5V4myZvhOju+clTmiVi9ZDJEkBfF5qfmhcOrn/f
op84mrWQAepm5XIj+2sdc+u9UbW0U7ncOLwerU0ckssVNGuk2nm5vNZvViDBPwvkicV5BC+7w5ng
OPdJUV+ZkDZnV5/vWl6gu9NCddz6l9GepyhZAsemOcNhbulAkk7L5gcu1QINQJWPSutvR7ovzJry
xPv17/cl2hlL77m3MxC5Bs9D1r4zjzV+nB43LvIee2Cn+YIr4AdCzGGfbKh5zjxh6L2MhabLepEt
JGMi72veduCge5T+tL/mPWs0LoW5bWLhyE/oufclvFbQM90+KCa76qd6nl5SYGp3BLEyzRne1tGN
Do/dAx999ohOszHumty0yR/5ZJ9aZcKWqCKx6pj9VSDcRss/WKg4GW0iy8y10rg6EYfoi+mNxAz8
eG/HkUuBZ7uaCgTspOe2Bb6eJpxO2twrIH93dbhI/qwG/+ehwxY6TOoys8eanfXF6RD2lXPGcWiG
ie3mKa2JP3zoDzmz4HfoDVr65N+XkEvwdOfVolIkJbegKBcRx6sA59uOzHApEq9un5zrq7g66CRH
g+RCqUX0iqjxIWGkRiTC5VdwvHMWr60lo1aZ7v1uKbZvWv+nUrkH5V6moC3dtQLSyoJ+X9JIQ/79
eC7VZF9nfsbEselznSr7oRF8IoM7WzMl0DbUrJxbEM99dzMpZfSYoj856h38EPXtwe0CIJwaEkKg
aEQsghppFfjUuj3m6gcfIj+jt2iooaG3oPBCRz3NXlE/ZPT/FIYkwNTN3kmCmXKOhvAXX+uuOx+d
SeDr42MWnCal35zvsI8aYvvPkky5wRlXOTAmsFdBs3dKjNQKv2EKc2WHFnvtNUWRr7t5ZABiJomW
SmsIWxYRTP+ILv6aMPmfMIz9aoXdLzF9QS8fDH27MkJZb3BA9tYNp3zT3g1mBClI3Jj48xLAU7Nz
9DVJrvcdAHcSI/nKLO35j4GsmaBBeYNaZcNqgigQbEuSYu/JcRJmDWeFnIIICOW+Q9l1ayPtK0ZA
+4sz2x/v9mW8JcL9Nq17m3Ru7JTc6NOd3+oaOPkQwk+Cagvs8svu2lUF7bmJBDNpzdlqyt+D0k/q
lGp9aZ8wL3yfcRAGvOys8SscquRsQh0WC+dqe7SeUpVB1sjiW17howfqN84Hje3pY3ubD+ewUi+4
CvA/z9xuSdPrkL4PsI8cU55akOWxQ7Y8OLKCaCi29tPhf14F4YA9eeLtwhyBEbxkS0G/O2zN0BM3
eb6C/qdkN4LBs+XgWPIolIQ9u22/69IjaIcVF1eQTVe/VLZUNF9mBpLEMKkN2IJykTttrLjU4h8a
EVhiM480fB7O4p/+eVTva4g+AASOT6/eXoeMrrdR00pNkDWmlH7lthzte41i8Di4oMsrCyWHfrEr
qI8fqm9rfnaFUBOC/IdziTCo0LgA+hd4ZuGcQx1OX8JWp8ATz4089Lc7/gVx5lPm5Vh6Nb5p6wXh
8xqmuOiUJOWD0CxAwkrSQ960o0MJE8ZmPBm8Bgh6ndT85nKrvBChSvbl/fyWXrSuZx+g+ZX5RH9Z
5bkc8VjNm3kOUiVdLcg/6kzaeWBHxdvR6ePiK6D0dquQhSWiI+TuCrGlbzAgJ5xb0caz+CUsoE72
jvd4BabjOG4G1JGjIc+ExN6M9THusWzLr90lC1JyEoqz0V5BwhsMqEdc5TaR7sLdB+120J+Hr4IZ
Hv8RYiqMe4GWQDhwtT0qWGArS59OQRTSRhNRy9UTFkzeoVfpymm6MdaO1MW7P1hPV4FszxWF2oBd
LkES1WdDnEU2hhp8yHZ3fxf5btQFxPOrtybvf9YnFD3FX3/ADasHZhgmURxLdu65CSHPL6lWFUMp
q+o9oKUrwULZI2urgao65HaLMoxLP3qnUzBZLteCUIWl5Yy8iIvaei3Q2b8+veu9B7mrY/1rLyp2
BdofOnN0T+QqSoi/Vz57zH5HQUSlGAnPAYgdtXGz7gmdFJ+BAy/7R1PUbrtgVra8d/CPZEMg4cas
wBWTVBZsvutZfGaP5WG+dFiOP8pJv+ID1XDP4E3zCyPCuMQ45ee0MV9AZYQsAN68nVZY4iwc1jJE
rBBugpVIwAQQvOqnfs63sYnOca5yB2WdaXBEVpfXpPuHW6EgKR13XNIfFIhRbd2lw1Nmho/6brbp
lggrsAuTnkhwHadv3ETLaYIN6NLOcAFlcvChOvuufLZHDuGX2F+a3DnOrTA6xRKBDajD652zisCz
2OI8rSkedy/lU0qsxBNtORwvp/isMB913o9wVzSj+erC3uxsV1jFZ9X08wUky9ki7SH8+usEMjJ3
yq70DF03GQmBYRUxJ0nVeBC3s7D5USFPHC+d9xabsjYWZEuMbAe+8Npe2XQfxQAkkNPcAV0DuOWF
P6rINsAZvVDZPqyhyDmDilVJXMrwUZg+MDmQxKbx2jxehnfHrO3RkLm7y80p3WPllRjKjx6vwu2U
NIYqb6qIzZoV0niZV5aap4WB6QS4nx8LyoID23tSiRDqzyZ0qK8ztG3d4oIldNoEH2nlWrLKFUBa
Ll0IECPxrBhvE7tISiBs7nRWd+CFN/23errcsvegsOTJmxUgydevZambVL+kuxOCc30Ri5KYPhva
ZT18XcvQUHGmB+4sUXR8vEZ0Bib+AO/D/oYc/4XdFGBPe+pxO9/7PTj69gxqBs+yd8LQf/PCCIAR
ykGrs5lRlm1JyhtkQ4m8U12bqGOX+az2uSGxqo5jnS7O54B+lT3cKispypZtBIZFAchtIJfGRQD1
Fi9SFZaFfZLnhmlsoHNpb76GNWsxW54a8zS3BoCLpDAkua4ZXo+IIhkuPJ9r4KocLWKxoJxL+Xpc
YInPuskn1DwFvMEuTuS2uEwN9ueIjLBV1oYyf73YMM6NxV4QyAmZiWt1eGtKiuBw13mgRZUEJLYM
sHgSwnVzrdyU5NbU7oBEv6CLzEMzoTr9CXLypvE9eK8bn/bnLUhkyL5kBSnOnE8fZpIFi6lE+Y4X
OAAQk3XzHvkga0PD1Kw7NL2G26GZB4sUpcfKQV43HMDD4xSQTjvnhFBNJUsP4dc3Cm7hgxcFntiI
Obi+p4Q2MTG38uxfE9coSo4KkCg9z7gMANDS8P9zCHwD0HkNsqnVGaMdOB0yV2qO0Cz8lfJPmwXo
+U8MmDZR/Iq7wPapNxUhx5CQ/P0/KOcOAqUH9CpwHniJgVUw6VZAcGwd6tcRXdz9R0MkcFm6U95V
KALacxqICZcVAlKFSKo3HsBT3f7luLCKQafnAP66ulg+1PZmBfx0p1nGMEjZslvKnWTjYK9raXDN
tMl0JGZAF8QifKT40/sNkEGjFx3krCJvnAz4KVOLTpKF+k5QbfmufSo+tKKssZ5ElnlC7FoeUgp2
7zwXiw/8dP5lTa2idkaOTAPQgvKuc8AWSh5JmgzCAcWKR8BQlJidHm4x2jXdlvdNQx3xnetpFu/5
mST/lGu5gdZ2tNM4UHGUam6piLGNvrUqB6cMBK4wr/p2jt2HhoZH/dozNDgrTnp20EAogdyaiEZN
8AjXxlEDci1BBYi1pqS82XnxNSk5nSvRY4Io10864GYzJkmiEa2pTFjIewJZ783203We4a9UiGs8
xxj96l3IxnNI7t3O6iDg+myQMjSwJk5uj0V45/kPIKRPX6o1SrJdW0ZZn8eNjyuwq4ewFakOufxW
iZVgv5qi+SySVvWDb7NZNGSqMRgWNBLhC5MyLcQFgLce4yHPl31Yim0wPJxvK/U2UnMaF4ZOlAT2
OltKpZrXIZM/M+hHd/3D8pZKnv644XDWvLo93YVYc5B9rJIArcWFhyNlBGwFQB0j1d2ty78gll4e
kR+oo1U0OEDCj/NjXOyBKGzcLxscsy1M8cyP5kzhjAQt5pEDidNqx69gi+NzRbemT0MdkVSitSu9
VV62g64Z3o+CPDX6ZTMO16IlEZXemZhyc9OYcB8gaaHHEKkXJgRa6ADftBn6YhBJ02VIgAy2O23M
rnXfp2t96psHYIiWh2EIlZx0uYSrS1C+qJLrOzCpBPgQpTxqKgsbPBlWpsH0/yepp0+6niZ8v4hW
em3pV79CK5doeq+4/esQPzItn1xm3j3ZzwouieO8RMeVuUqqDE9ABthriQ8Qd5pf1v9oP0Pg+s6A
P4uaM0gpp8mNcfZTozpDkourhZXvVw6fEMxBkQ4AcaZKoV8dz/fxugwtIJUc2j+OUClzVDmzNGos
Lw0ccxgMnApcsqGZx2QnNrLmk3PptntxwVRyQtf0ErLwwUZuAprz99YCAwhUxegTXNCHAa3YuTmr
UUmYQ5Stg8qbkUMBsGahBHmVEdhabISYZfZmclVp6MgVB0miexrF37Y2QDMFefkqm5tRdk0TfHCM
KTlOsaehYjxzIcca5esxGcLEFvSTGb3o4e+y5H0Wg6ldo/+IT1zWxLMdYJEmg7eiClvRMxXy9fKJ
Z8ZrElIbBrwAT3HPcNPPuVq43UVsoWZzcvqeibdSHSmqnGUYB2MQ4smzTQq0NUJ9BK/XISSptFdK
Ob/3O8uyUjRklNdhJXsEjhVO7B1qvJ5qPvkT7ACGe9fvw/nSYnPlm2PbfYyDhYUT1QECMl+yKEMv
09GxEbZQVVt4UYwOkWJVSGUbCBq8d4IBS2qc0+cYhy1E37K1pm1+CrAMD+uotQGCYZ7VTfwFdbPE
c6tAHV1AOBDFFd9lFD7MkbIOPXQTeg79ILXT4wOYcYMJSwLmpzD6TwSHTmiAllzAfPc8tuOI3w8S
48IkzNakw6ArqtTDnM31K5GAhizzrRSeaIF1ZwUwA90HZay+K9HQpKIXSIUHULqFoZT90KTyL8D6
QXG44FnDrV9FDFwmvgEIcr3SB9aWdwVZD1iZC9TNBOMeFIHH7MvGkIplJiPUc1b6q+exTqJq16eR
Za7AlZE1bph4c9BQS26en7nhGP4wlusAUWjvQzg/DNK1FjmN1BX4A4ECw5JwS8l2nTWVLRX/kD98
J9up/ZHULgaxnHh0jdu9PuSdTd/8groF6kCCZffZ4/Dfq4KO8my2v2zjYt1EwF5XO0Am0Q5AAcDY
MBesufsTKxm2vE4+SAyXXu5BQwmcO1nN1FKMI9WxgvjpTDUZF8YiNmRz9r+uiRM51qKlLeTC6vJ4
ivWXJNbBMO+4EXtty12HhL3dyZrKjgzzv6kxV0a+gpv7VWThL0Z3UzuuxTrBhzPkgbCV5hsBvsmY
YcFEWXxS5I9g7bEsL2FNBZr0tXdyKVZPdpCckggUlCCvv4ROzG3lkNdaTmj1yjtM9jIXIk1HWIfm
P88AvQ49UQ+heeWl4+G8nlq4Cv75CzIyyxdZILkgCZfaMifZ3gJv17RvGwzlEHYO/ZDtd3m2Chp+
RFDhVX3gEQxAu00A4OY6pduamK5VXDdpuXgvafgg0Wj+clfm2wwCDaAtDddt1RR1ktmCSjvRyl0h
z/KDp5n81m1OhZGVVguizTvZBcPu4gmH4BDLwqV1iwtQK/ziGQOLiXbgvklU7SRRequHZF5igMIO
m/0yQHjusnJEEmuFF33O6bANbAbBK/JVEiN7ujFquAZaFhVHxpGxppQozrEHZOLxL1YiiySAoQ/V
JzYpZv9qwArv7QcokjrsQHCD/nkLmm8ATfMSd1VwtsoJRqJjI6ue7emoF1VMA60XxE6fU15ckD0x
+HSX31qB6LO4y4joag+nALwOElZqryDheN6FDrlnQkuK1i5va7678IVTeEvYhAeY9RuFhf9geiKV
TUsR5lhtIOn3R5B0cuOMF8z3Ak5G70WiE1XkhFop0sUVqQ0zTSvBXDd9DaSZO4Of7YWrK2WhqXqc
yDyMmutpWLX8TrHA/xTHzC+ZFWls6RX3W2YPyXK3KlabXl5WbR6cu71DAPQmAWkNTeYhDmmXE25c
QsgY3dwsLSggLc3+dLtAWF+oMv6ktJCZvjdhqtB1Vmkd03N6ew7I3H/ol+YCQVyGAWk4oVh/v30/
KTowv2cdWnt15p8MrxfAYcmjdNviLSwHCPVzaw4CenEzrcDHVpT8jvpn1e0SELtnOtQQmuXS6s0R
Z6mjz4eNZGRP7u5vaO/WPqMHAzwUyLEhsRSbg3nIPrF7ZMumCyLgGcKm9m2pYG6B2/5RrmwHtwpH
fqYT00oIV2dm5zGjxP5AK0YI8MBItFc1upPw179/O9pmnU/VrqxS96STK6QtlywbzLPvnuiwg5FV
l2/NvwZspCk01KFEEJsxeSAtaBDQKa35M0VtWe6zqy/f29r0IHjQSTf4UA4e5FTe2Ul25+37KrND
GL/BcoDt8ulBMSeWmhFWoTbKmIPv2yaUUZQStjCpte9+dXciKmQQsEqOC6f7x4AKMBWHK6TTsoEu
maeiM26aki1Dz5BVf2LTnIp6LkOm36pd28jZyXeL/8jfxvtY9CNQOQw0z5jQlOplmyogCsPgnuIh
9vpnAj7kt1umweg2QdhltMMnn6uqZ/KSgsTYKK2sUaTbCUlkS1+VDapNhoZ0BGpdearExBn7Xvzs
i4aobZggZQ4V5jED8N8mTWAXNZulRKnSv3ZMhbYLtuYzhXAt41voN1myQmTGpJg310od2bRafcqz
atJj1gYayPDDyV9sLUfruHK/VGA7rA/y5oXKoyG7sAqLI0JHUQuKOgCaoGRzNrbWOB36WKL/M2OQ
8EU3ZQBOyNt8CBSTlVD8L1OmTfbPJ4+GTeXKk7Iz9p2qy1mg/OfFjDYkNzMc4PvP5n4rZsxkrYdn
foJoSbnmxgyaEKG7O8Pjq17vMTWptaGEg9R/H8/IWv0DX/PXvmLjPh44oSCCqLPNLgHu+ZfPjzd0
mMrZUwwQO4MZDEJXfZEGODK2QOt0ciQsGB+ZoLduHRGvsxyuc1QtNUbfnz/hIKLuMHv+c6/pA1fa
sTAeQCB+wR1k73ErF3+t2rAy2bZgFPvoR16+UnGO8bTCTAQbFvwEjSeK1hq00e35VOvTG7HEpY02
g9TRVE1qHzUbhZ2Vs5BFT9hzXmZl+mMMmaqjx29ejvTLzEw5I55jmVyTIW+NJUyicbHIGH0cO9Bs
sVkR4AJa0BLFiZjlR1W/vZP2gvNQhDYWvpWFVMx/zWerS2xOym13CIZAApn5IflDVpl6YRMgijJJ
vXfKb91CcjnddRKmTAJFBDs2nIjdjfaZTEppwdBzkLC1STFGwTHmybjl/50sJQ7ZT0hYLm4atB8a
C/9qwdHdbhQ5AQrsthfZFvkkOcfPEeC2XQngug9jeIX+P3R+irr1zjfpjVcqPqGU079/arE5En/5
oMkZqS3rYo6X+eN++oPnqnew/tKDVN1vlcZBPhTvmEpbewAChO7DHdTamZhbWmjnPMq9W9dSjQCH
Ww9IXBqGVE3shq2NMy/xjBSm/N6dqpD0RdPOBqZvfOacEeOFREZ5wxGOQEjA5ecXd0e5MNt26PjW
PeeUqM6n1UmK3ITCD+ETZGaL5K3VsKYVPf5ONxWgfQYIlhW6av1HksrRqjNpvBM1ZU18J8OwNdyE
iWgW3XrQUANEQqcvWdeBc0sycdLdtt9OnVC5TVRyjjKpjhDinRKwRXu0ma6U7N89FRCxv4b1ceYL
RiEc8vC8UbgVifyMfBIlJXyI1gv0/jTza/r8cTve3B07MH5sx2IZKMB+fay3zvqyLCoIB/C6guTI
dfv+6aKwU8J+mFjscGZgoP8bvlU05se8f4giUq9Zjohpqrhc2Tc9NPmYLgNGi83HV2mG7sk+jmS5
7zeU8o5xCsbsZD+/fNciAkzNt3h/5W1ISDHIwcJkHRMUVSilJ8E27DeUrWsJFQ9oOsa1JcNu8yrw
315iIVGhn8kWHJAqGfpAFxusixG0sKRLzWrDyZSGRmEoWpmX1q6dZDKoEQE33xpMD0aP+2BijNJb
IZLXTsS0VrgydYB4XAVnjj75jDuIVfJsHX+4H1Bcppnq+CGbnMjbxNU31HbLok18lqQ7e/fGUMKF
UNaqLXHNLLykVX4Nfbpc+beRCTP3eoHXAWkNu4hmu//FX1K3lGE6P0xxcAYipSKf6K7n425Ost8d
CI6QiqKYyeb5ePDkvQKJkY4+lvRoviJHZ+9finhEvzcDQAgaPonLV5EgjR50TVkRbD1YK8ebzlzx
5LNAhHBGb7edHojmkYgTVFzp96LCApkX2foNibCnKVhBt+fJ3mOnTl3AGvd3DG+HksEfDtK4WBO/
jkyUYJR4aMt9blOm3VVanSoogBZKPsqA9C43mWAUbJHf8x0jTHlaitVAuXLq8b3v0h9PMG3nzUi4
ntsT+1ZUWc0R8P8hUHUllKvxUK8kKiscfZa0/XtA4yR8i7DRRZ+CpxTAwNk9Rf0UGZ4vH6nkmA5M
7vo0+xxYEpeXy4v4KgSmIaOkJQWmLlp+GoF8Od8IS3hpqSoxh/Yvh9DPhJfHrpaz3HnEDyOG5MN0
ZhjFWZVlYvPUW+XLXy/0CXoT3mRZvBwwjTH1KRn8Tb7WYriBZ+VaQZGppKs4r/PyLhWPxQqAlgmv
iuQMEGcnBwPMSd2MazJovvyqMlxl37uJ4lBF5/nIh9gikIq0wztlkQjZGiorxTqUt7leD6SbqfMJ
jYPSgAB7+WgfuVfkEM1tamrKLDbbCHS+4DXMiRaJ7dtGjrriwT7rumwJJ203pITbNqbgHjJs6+TB
rPL3TkCAYJTlL9c6I2E2ELSb/7QMZrUgo7fuwuy8jKge5xElt6eyCpMN0WnNamwA2p3JEkPP5HXa
mYs0b35J3ieyySfiqxJmCWf/K2GnGmPUrMbMilfo62LqMTlGhuANDUu/iksLhWRuEAnu2JP7XnVE
cG0l+aKvZhYFbAeZ+C9V1IQ4vIVr2RyA4vxIVDVxeTLg1CtMZdOAhPSQgatHMFsZu7nfK38LR0eX
nUuYe0AjyWjiSR96K0VIImLCnxYjK+HpjEzBEfFjHHTk4nfctO2B27BFWrSNERyMPmXaErT/kOX/
7UKtrNnvOUQ2mXtEpII+OzuuGrggDCAsotmXC7wSChsz60BRmSq902u2yxNE7c+JR3I6qgUDNu9n
bcOqSyTyzVaV2e0pdZJVBB4U0NOeSbX0SYHAVmyy7cZGNX1AwqUbFIAH7nJ9cVfDkGB4ZapxRIBt
tkSgIGC5t90Bjahtdzek6jSR8yfSBFiN9xiP0Y7PVuptp30wldixSZYT7GXfuy1xmg484mVPi6yi
f0Sg7oyUyK91G7okor6Z8Onqa8MIPbsjKZx9au5L0oC+5b3/HOdjm857gy61TZHpTslzY8tmSpFb
VCBDKfAtoe97vOwP97pQ/Db9DSCGlnLar+xFNCXsoa7EEfo5QGkCzRacW9QsvmVt2XkouK7mGwC0
hzp06l/byQqv9SKcoD46oPyZeRo5v/cR8Ih120dE2AZ7wTU/sOWp2f0qDCKuT61KQW1wWQ1s8qQs
JY27QfThBU9ukeby2TC5Sj+y3u+jlz7oYOZgh90oYEV7I/NkNY3CRscc/P7fIIWBiA/8nueBIU92
Y1h/W615HVW3s0Vh8qVl5Yyqa3DMbp4VzBC4/E/eCbDu/5FgfvRclGWlaONh6S7hF9gwIjgR5qbQ
M3VqhipwPiuQzGGFuzBvast7upTlyp2BTl3ykJm8L2ioLMXay6inB/EMSo5QRpu6NuLWk4EaG3Wo
DOmRqxvg/hmFYYGjJGzzLpG8DCitFk8POHL6xpPla8YugJQDDXup0sXSwnyKqpnMdbskG/UmZqJ7
sSVe0yoy/6cz6TT9aSFFR9S3LBNCGlniHK+st6ihaLrNzzN0WSWP9coOM3M2GzK1JsN6cWkrI3Aj
NrNGiNFKzgkIYwEQDz91wyIuKyrPs883P+ojc3Hd8nYldN2w+4Z7hE2VavUyy0SVGwVnwf/nbShX
lMcHhiJnrT3kV4gNTVr3n3YgBA9BT5+pv/JVA/6ttfIFA/oIEh+VOFGvQN7evK90vJAV8L72cXA5
qyBcZp5SL9wxoMWbp2lwjnOp+4fzCfDOAqZ5KJwv95psF2rqVkbkzKGydf0H3YfRiPdG4iyT0S84
YpF0bqAtVwbHEiF1EOr/ZXnJ9amBmM0SjBYsDk96hWxqDc+heSeq5XkOb/ZI2lTe/pCOD3Au1qdg
kl3L1AcypEH/QNR9H1/jSPO2lC4pc31izX4p4lg43fkSw02vyglOtwVLRW/nRJpaXE9O1mV8aQJk
7+1PrDZMx1/ys5C9TMlzk58Yz4vnxSi8ye0VuOdh8AJsc/2ZcUXSKJWOlxVuoAc0ErWadkbip+VW
y8I25qg/2cWrLwEj9p3IHHfVUDFpyZyZ7abE2KTsxR/MCrV2nSyDtW30T+bfYSCr6qfWahGGsFjk
evMXaQt7tWLRGzFTIypjQClYxfn6lZbJx1ybJoH02zCaugfo5GFCu3hI5QD6+BP70YTv64TCUC5y
S5b+cuE5mmVwzfNMBArgOxE7jj3Jz5saJ4wbosi5ZEwYaiB3wtKC+UB+Oz29pKf1vAilFHm7X9aA
/S8E1chsF0R4MI553aNc4I0aDtk3JhvUxcVTzC+b8nZoONJV9WTUE58hKRjcfqsjcZMHN7L55Nm4
qGUP4ZQZVSnwafqzCIts8sD1Q+0UiXRBE23UcN2XX1f900KllF2UHcDY1vpyDLTRGtD2WccrlhIs
5JMasnBgbj+J1gZlIt0BTbwMt/5DtemlkwIzHDxuAp3v+NGSm8d5V/d+h7aacvuSgf8Lp/tm3ang
PtVRtmGXqldV6U4l1VVfaSoRwgQgiWRyBY3KfnMcgAexbaLaYdNaKACKleoMtxiZs8/alTtOC+n1
QT1DhdNAnOFGVyiQ2NOWnVolU5ZAQV6S+CQfzvpq0Yl4H0cODnX8danbAdkqXiYJxD/tPlRRwCaz
5IfVaiLmKNICN+S4oEsgjeG6loIm39a2dh+M4uFTKbGxJiqWDRe/49lqzfemn3QqDt/mHMfMtMTk
yZC6IFO1m1qOYhCEsYwVzAVpJTLbYva2YLTQnU7Em6n7igpZODfIT0H4HdnKlzh3NdDwwvCfHxce
8bbagM+RlkXnMecsV6EqQ6pdHnnRqtNBnDZPis2IR/Xv4/iTijwvQ2/zBF5c+7HoZxG7wevohL+n
yHDIViaJ6dYBZGYNSOjsI2/AESifj1tQtBDVB3TN+yjfwx9J00Xk+PvkUkY1WifgpBeg1gkGIdIg
jeqiunzmvk3KRIlU6Nh7qgs0MFGbdPwEzCK3/ZT+f5ypb2IbX4jas5JyWvE6mxcdXwj3pyGvM+ei
7/PKkAf3ORCzEbNVqJJ+2GNebhs8mlR63EIKApYak7MAG0Rh06JY/LOVWBytFPWgTzsWANzcWHWZ
ZkDNQfdkZ033qBcwyS14dIp9WQV3BmetGo9nAKemYvLi+UB3p35iLUXEWSolygid6gZsJZGRAj9M
NYXhCOg3Ad4i6Cf/D1PrNNaC31y2m1XyDVwNF4pyAV4ycScQdQGBf46rgKXI92SQdrQJDxcQ8448
S/O3mwT1ZMbZ/jD9ApJMHR8xRUaMx3odyNu9pvrVaM013XoJIOL56HpeN1f/+tFwreqDEAB3FK0o
NJIZgOzl60vVyL30UctIl1jaGQVt5aQMCR5f5Gsh1g2ST+DrASL2D07m0Z1AKFtA7S5XCQYv0FnF
nOWH7M5TeDD0KxcFjQ3E/n13n8tYx9V534xvD9lzLOBID1qZ0dRa6xVGAXJ6zbSrEn1yGbPCx1Nw
mZbpI8XIdcmLY4Yd4PpgaqqQgao43WZnQNd1rQGheQQEzDx+p+BUBSqkCcCFBZuVyjhYttPiVWzo
sjpGnZxmd1k3yjBWePcHVC2XDbKdAubAFdgrkC/LX1BKRAFpWY461ijAFe+ZtxGi3eiwMXDPwiFI
IeszDjASJv+YVI1VfdkS3VvmkfkzTPKGTGzFpteYbpkw4uU7usuA+lz7kbGerqbDkJQ3k+OGCsbF
zVue6bbYa/3SLxGOeT++CSTikXTr1wOZNxvyk3xtU3qONfUjlHTIrz2G/C+QDg048VMVCpRuaGqa
na7PI/KiEr6leRwXyCSmGYszMwC35KWxnhcBqPzgl+vBu/LDer7S/LHbQGL4CS7p7nsLfXq2NYyB
RMGp/rF1Uvl+lPh1A0Lq22O4boThC0xFdwGEw4YTBJatbg/dBEfpcLGtclB+Fftg3he9N4piysZf
NsFocvVeKvl5pX9WpJlYQi8qhtTQFw2OzqwS7sQzyucLE/uXli1D2Lr5AXo7FHBjZ5+0rvs1VQkw
Sk1rI3z105nW5oBjLubXnN7m8Vvw341VG3Kkr8UIR9kpiuQTS8udy+ptJSLz85JgE4LVeyVWwcUn
rTrSKhcBLm9uVQ/ehbocMqLjPaF1jffSS2RUeboL1czIKNQFq/6tFm5NZSe/tbqgEtatRUXz9utg
hGhd/uEULTJNdOYj/wP01TSWwsJeh6bQ7FPMYOhiKvya82FKjWgf1mbsDRlcUpjDD7YIvd6u/iPM
AATQ7fLRMPCBMLsH8V4uKegrLoNWgiHPtyJcjI3xnLPJtG1FhP09aG5GW6BQ2Yu1UFam8vwpo9Zm
qXrtNFPZWMxd+LnRuEpMNRRNCBrI2dMRDUnrNNrBvbApMnVA/KCvdJjqlyQxF2hjQSigALS0IklF
O73HEAbmKEtzc27aKMRIPyEnFX0KBANoNuZjeDDgb6Gv04D9HTgQG1rKW4oNrRxlRkFSjmwzTYab
Nr/VQJ3i48ykc9kU//p7TjJUXe/mXImIIifq8Rjibdc53QPMg08SAgRKJnxJ5L6vHQcSlycJtxZi
bupg3bjMb4B25FwzPzQ/orpgUEzG/r8f0J/79Jon84HlYA/yl0PfDRXOOqfIWJvQFxu6DHKrewbl
VZjCJ6c9pQjWzAXC8MGfSTyaecssaO3wIYcASag1ORQL8Cdy822G2VfvOZtYER9ZHey5NbMm5zC3
pluNVPRNo1c6rZdhCSV1rCLKojJUPvy+Jt+NgwgqfHZDMhNbBfyPttNeF2yizPephZFZ8I3Ld5qW
j1z9QuA4uusVkEtZxEk4aZgOg3zknfVSNInNoPLE+qdSAeY6qXv0uYlaKALoe0160+dbj09W9lde
tlukhrz22ANx7KQWswshu6giyzXEGPUrHGm1uGV2m8QYkhEYoSzPFJuBYPFhRZvwhmIGQsj6L866
f3jUJmuqWE+ZxUXC8b5RQn54++CArDAT1FWvz8WsSdYp9p7aTdKagbCEKmnETfY6okXSbS/0AvLj
i2dDWCCRaoC3CoRGTbdrwzmuYakNSxwp60wmezQKQ41HCtK0hzALMN0qDiWgNmvMbL5JHycRtn5g
TJZuH5/rOe8SHE2Ij8npTd98DmDaM2N4d3D43uppb+vsBbcPQ2E3EnmEl/BibiEl7dAL+XPZxXLl
JktRGL8uth6KdUZ0QRMU5O2X1rELasQB77OFmf5ZLT6DT1ypOytku1XaSYZXOgpCOjv0jsk7FF74
edCXltLZV8pDg4nqKNOQpHEzUAaNBXCBUciOkRF9txpupuhFvGBJLQSpR3sojRB+Yz/LnN/qdsg1
G4Rw+vrdR2GHasdH0lt4iNrpQ0OQpk8dPShMsrIZunbw2etYFvWSau2yhGnOhH7cMhdgCkE1iOWT
t+HlWCvJx90MXjqwsIDAsvkeb0dLeFmCm6NfXz1tSmcK+cv6ZclreMyb5K4FyWpYGoYGiVmQbtoj
pHWXjUNG9tQTgqmQJC2RD70hcGQ0gQSBIJQhh81WtT67IaizjrhI0VGKWIBiLZvG2XVKfZABtua9
dVol3ghx+VIcRTYAOGOlq7RLyUj+gkMxnfjG8ckOC5ypqAu2nQU+/LEh/h0PbNwvviJObPPkHR6+
M1MHTivI4D9EklRjoOSSr8wucXgpiMiCx9VIX1X8ljHgDeBLwKQ6bWeVI513i6nGW6EI6BZm/3dZ
AcIrGSaSvFCknvHWUbMn1Fr/iXVxmIkBBW1t4yyzmIW75iNWBrN7diGNZCQWTPDineHxXhgMh6kX
mVFsUmsBz+fsBqv9bQUk7JccWiZRHKrT/5acYbVPwEL7Y22FMzXUmHt2mQ9MVIKpAP0P00HI32p0
JZOUC6AQk9He1X40B1FoyctdqkRn3rYn9D5RyMkYqvsCdnj70u2SwS54lRuvG10l56Wr41xvmUma
eVHTH4pmeKZdeUkiZmYyhKKD1EnEQMYh0WxlKcueLGUlgmKNQhypYuGV3Lj2rsw4J5miP6btGEaz
7ED91XUWAxessbS7DjMQqItlWBITX3KZC5zolLg+KMCKvJ3YKFrL5MTF1QJWhPRKa35SibLj66ZY
3QCqqUkUqfYljE5udK36jbkY+JDAGl33qaiPnb8VhLQJhAuNImH26u1e0XU7Jwk08Chf4axz0Vfl
lp5tUqGEQjvkwhqHtXpOGLFU3+tOxVbYdMqLXjudle8zyjfxgljdvmkuPVqMjSMxSpMvh4vKH5rZ
Gt+5xrShXmkHjgc2WTeUBdH1zBvTQAReXFSUyctztefsy3SVJBZR5SWWxZhNL7ZzqqVYyZTNVlsJ
Q8KmaUNh63N81Ce7sYKDdGmQrXwcPY/+ZW6bDZuVe4CoSSFcbcRWTh/zwzf3FJ5TneHEshYqc7gT
sFvilY1RJ70G0FhIdx/344u/IQRe+3jI+w1OAMlZK2Gch8pxnHAjDqmgAqPFZWVGTqoarL5/1f+W
wiX6hv6U/XXWxhSejGazGal0Lvr0cEElD3DierHyECPf++Q8ZOAE2t6b83VWTuyimbmtFkf5X+Da
Y0wZSHuyA986akmEXDVluFb8/VbdxIIXSANMkWI+JK3iWDuk/D1XF7KbD/BiSKM0Ae+jMZWDXeeo
Z9/kzCqqakedh+3NNk/x1WsMqPnq4XYNLP6KSqlFPhM35DXpBOpAHIGlYCIm2TldWNXCD7UsvrA+
vo9Y5UVAdik3g84TsniZt46fhrtbSMUZOQSL4mNMpzRIYJwM7FUcwFOjKfDUYpFnHHTWA+RB9czN
m3lFvPxAXzW3BDk6LjcDSAsT9chBhAt+8oT6TlY01yKVkKrQvTFVSAI16Muaoy1FdbZOmn3+bffR
/BamwgO+LzBetat4uV30YKicDhONn4cDV95a7RfjO0EmQhlXwwBsRvrkz3171l+TV3Z74iu+7tMx
G301EQCKBfMHlO9d+V8N3uZA2bB29ol3KgbDI/xz6M1MxFPBD6rgHWS6HrkXtuvbChKKJfEtF/QP
7vMU7muyxXxrZJiV/Ag5ObwoGszdPlurmEABfu81Fz8l+p7SOslriU/RnQXo5AOx0rNam9GoKSQY
UHjZ5Kq1SQKpOnp4MC0Fng7pqofINO9NHnYKYNJbVRLJl7ZRhH7yZ4JJ1BWPIvHOudx3N55Gdvt2
QwMymYmdhWwP+jXoYMzAzmED6pkMcyi2XmiAMqkuWaLTNZ6+xl4BCeBj/P3IuCqn2sdvun7mOgPK
Ds/ZplrRY/SGSSpCGqPDJUWLqHmwP2mSNUuAnAA7fC4cLZ1BsCq81cMtOVjN+x/3w9x76D1+ZtQf
Wwybx3iZHBoDf8gbDgoPyfnf5szgs6FIZDBaLPn5Uwp/TGG/lQtSC6rontUqsrsKNA+Iv95rRqe1
fBWrDsIlzS7W6nHW8QMcNGBsNoJ5dUF/4K78ia+XX0XwrJZyZzNOsvhu9fNTA6Phb12A4hArDCA1
I2lFpkL32IlHY3zCBS0JtX1BMm2uuYj0DvURr9B3qSrlb+e4UKCQB3qDiYxpPpOvg+zeJup5Fs6X
3LRBemNHT4dlPlCiyuGR+LCkQppzVk+F/iKpOLm2fg58Rh9rQdSb2ed6y9Qzf9M6pxDzwzUlHPFf
nBV4xgswHtW3KtSsRbWgCD2TbUd6ScDGO4fPifBwLwZzGsH4KWgelzB6VZoEjEbUN6kfCm1ZXa1O
AtgnFie507msdd3w7L2+RhcgNJfsmvwoQhwpAqpCt/XL+dMoKTTt/PQR3/A0H6X0iW2KIU/wW27M
Y7jEmT7Nem/g4zXD5d0/fmK3GJccKX6yjNJ+rTycgjChSSLjen3VwtvayzB8HOYb+IdWqvfd+cAu
YzEt3vfLMUQNipIv8rTeI7ut5iJfgrPcgrXlyXhCbSx5GWlfSuQYdksgdZVB4S9x/gElj/KTDX3F
tuhubYvkDvmvsOp0HqBTPUkCHXy/pOoCT3q2csCstpHiey4FR9CropBR9aCZwrYCSy9U4PvqIGtP
OR284XjWw4TPoy2YChavS0DisYkN2OUaYXQmkyuUESbdUs64tR9bZ60C1B/KuSuYja2/WqQcHmHP
6FqJKOPEI2Q5aBhPNpX2UXYvuG37md9PFcYOjQAMK+JPbb9o6vpoIk2ZDm4IL00KgQRgONWAz9Fj
Vsxl+j9RLSVBaNMLnuN95XT5PfFHMbTDbNVirIMVLtTdos+u+2yCTPWp/mKUMFDi16GKDFImaFOS
P4fdyxpudcuTQ3z1oXmmS8XIn0CUJ0GsTkCJFviXxKHasSgTbbRsGcbfEbT+HtYut0qrAxwU0vPV
/JfpT5JvydUYExBvIKgZudwTpIWAiglRlKNBGHjiGacHaFcyjjR6Jqo8lEGBkeqFUwaGNhmPo7/6
/NiMBA5FUhU/M1YhqOcTogZ1k1KD9C98mhXKJ+pEUAGKL3srsY5VMZAxFuxL0DeiRey2MttUCZKc
UNN4WhIAe7dKvvwxy313LuzBhWlFjrMcdDgGv/ueD3vEJcy87efInmSdt4v/sjBdbwioy9VOZucf
AsmywuVp60JTEHf0aWF72AV0Wl5DK/H9aP2RoGmJBdwN/7UrW3xctBdV0M/38hFQOotICCkhYV7/
K+2sCjzAr4SAyDWhgOJj1BDBuwVg4ulM+kdMChycuiv5O4zscjGiTPFQhnMn5p0tNxzsHEH9jx8f
bkKRioqiyC/FlMTD00pCE5TACGXZFjb60GF29H/Ys0UsRDCXIjKKOHQsVVqK2p6q5RThAfXCltY8
yQ0Ve8CfqaooPJwud0U9YBWQLCoIitveZUHbIga8qEjNtm+QwoaWwxjlo3lPaga+g2B7RmrXG/Rz
nysyY5sXuZKvNa+QAwaSlh9Yp1Zg6fhnpyuTRqOzYncG4xFApF59/UBHinTu5fXuTBTwBZ5R1w5R
c8em/PJDWTjRMz/JeS88+idGXnYUOQzlYU2xwyFTQuVJdpbSk/I/5l2x/n0uGjnBpmqkYRdRjwjO
sA9DS876RoZrIRQfAsFGZiK7PVFslO3daVkn1XzJSCLTCp8YAH1O78Cqy8h9bHPVFuZEMHkYIkmg
W6LvIoOnV2gEQDR9IeCz/jqThcu6qN+8pEYBp1owTvgtJlFk1BKVoICW7ZHc0FgLit1NUrEG2yUf
l84ELK0uLnxsiKe5wJ+zVEyI2f1m0xNe3OZzycD0khxi2LtL1pcbIds7CjQQagwI45SVtg7O2MVV
QdrSmqewOty6HWqrzVU6/2CDRHrcErP1+ArScDI2fUtIzs1P98FfBWfCyBLF6mAQzpVhmZbKcVM3
v9AeW+d3utriRlHU+vj2XdYpYdgdwB9fPwEMU7FF3NltkWWNbFmhLsaWDg1WqMFNxuxDOpE9TJkR
/b4pQbA0TXkaXaFHPPdB6gw3TVfRzDf3W/8mMozST1Wa7w9TPE3WTdFJ2GTMSDoLvozAJjU4X1hc
DKIDE3XpQ3zuU+2UQxDJVKRKcSZJAoEmHw4ErInyKRDru515PHTew4/rP3Y2otfhU5aVlu1aFpjX
g4p9cJXGx5jypIpR1uhkLkiTacBwsW3RbFnPOUrR+iWE09MNiohZWy/oQG6TmSqK2x1jxacbk2zB
9qjibkeEdMybIb6BuZAeu0/1STQ+P8lY4Z9U8u6MvEkS9+xwHPX0B7o7Qyd0meEBHRslxUbEkPpF
bs+XvY2U+P9xWI/P3jKPVcR5N4VE93SjNqEA9UicPCIxxxC/UBMER1jHhiUYHLUBXuuYg8XhEgZC
eGWw6nooyaI8k/W1ZBl/UyL1fX0r3+qeI5IvKSfWDtVHFcEjMA/pqiG6NBq+RI2+iTDVOU0DqmXc
z9g4al8pTgrpTbOJBuVoh4cGNHYdgMVtWq/L9gRtTbKDtlapHlPRjU0InJNuWzVO2EkncT7w30wV
7OhosSeqZPh6tVSKEiDUf27x8b28yozUBkDmfzN47kVG03servMELhlRLBjw+ixVN01QVxuboiGy
4g9pc7x1jpgePMdRIH1JuVOB/Bc7GZmVNh91Psn1lU3qbAwD/AhqeeuOa6ht0jZIUx9N2ZdJuwck
TWvotG9MhyoIjw6RG4oOM3tGt3TmlwekCq1ZsaBfOVKzfB37pYvu/22nT7ZTCY9BrH5MC9sS5qgR
rF0gDkP4DKb547e1Hh9aqzW6GqR7uPMN1QIZ1pAATN/IJM/9lw/Mpw84GPyLc2lmm/DlzqFKkl7r
dtpwKIuFVOLk9rh7IPQILKkp1nptbo/J+g8HdxH/fokiqUw65IEFmOC45VxFn9BK3ZUtYRUtB4iO
v6d0VwZkn6KMOsCRndZidOfH/szwclMT0yv12V0csVpuhbtNIIrAoShOz6ozlFgTIH1xZBA3KzSo
zpE6ket+9XPl4tQvwIlwyKVLv6IWuSVqovdMqcpwmCbMzvpuJkONKkYXItr52xlLSEqQA+RdAL2F
mpRmxICy56JYOAVdGIAa04cOjDDisM5jVBW+mmM5lIoul0UHwvzgy1hQQQwCongL80x++9+1nofD
pSCBPTv/ie+Vd/XAA4J2/F27iPYkA42R7SY3yB3SQ1FXhrWwZem8GsJEIvnqKjsdDHzs74NCdgnG
3MXk+TJh+eqa6Sf5SnmFezdu9amBXB248vhhfeY028cYjHPqOFw3Tei/0tYAuotSKT2kXRX0KnTn
kMCPw/hoYcxBslIMHq2ZM9i34df2P4eddXp2nllNjOqZBzw96AMmgi3GfI4IFtHRYbPhRWQcVNxl
rBQNuvV0wdghK2vF7Ol5H5HsW9JvJLHR0TroWt4xyoGnGq29UBJe4ix9jcJy/WuOTeD343VVeKik
y9RrthZvLskGZJmXBGwVgfNR99VAAR7HNVmA6/fPVHZNMM/i9EVHyxC7SRKTRegQZV+W2NQxe/vT
iol0dw5AkGHLRl2tI6DINo9B6MAyfLswTnTr7k0dIGsXq8It+WGtED8gpNikVZhYXsWoHoxZ3jCp
lASzbBBezxYlKFnjTA5GGpYY/PwndZezKBdq9MCeSHBNix3E9RdPYyKUee9A78SVB2eTcWi++qHQ
B0J5+yneaXLIfiYho5HeW4+/VCDrvYyRAd5xJpdCS+vH6b29Cet0Z889+2A1c0Kb6mc9273nneED
04u1NFdPnk8Jy2uwIcGdstdu4EofcXfR7tX/fOXtkg/fp7cGrkiDC097gk4YGVPAk2veaRJRJKGi
/pCQ+WAEYXZ8pq0wDCjMJSlw3pSJx0fJG6/U5HTctOBklMChRXL3R8JDdMh5IkOG9GmCpTocdUuX
A8m+OalWXwtltMDXg4Y+MlwOnKdzzz+JnZ+lIP2EeugMSg6hMe24SVTzThWQhlOXWc3Z4TNGS//n
1wIEZmuMIeKtoDu73m+hf2QREAygEAG5YZX2LWKwo4n6/TUeRn0kLY6Uzctuy2pX8bRQlHk4t9mk
nOUK1CiTDqFe5p9OfipBW+2pi5g/6oFwbAaxqKd3zslm1587oloPzppnaTiccDg4kZNPRsTqL1N4
XGV2qZnzzrncjcJBx7l3dOUHWY0rHJU+KGkdYYeNWKO0OBseXnkASitbjq4bw5yZIsSTL6vHpG/I
97xV7M0xDvR1R43A/LC76avIIl5DBzPr4Qg4JAqRnPn2NT7+tUdaV07G/tYX4RwyoLjcbAN4LNHt
THs3JHNiqeIAjZJqu0wr6lDz7VTJImFyCjANqCuBk6idsg/rCqvzGEEDDGQbiafjIYOWI5OdTWGt
O6HM0iNqUds44gL5RSwEIda7kVpOPYUH1ovG+t8yWpFlZWn/mV1+znwIeW55eJXW0Qs36Ah028Zp
srfNErM7q8YxrDS3VZk9glRECPANhqLrm/7CYoQwaeLY0Z1mZHJLVSnz2a3f/laYPHMe7tDuU2Yg
sNhHsbO3xJJC+3Nxai3faJY1WtXnpRmoPOMuF1L6r5SI2XydCkJmKkPUTKsrXKXLSajLMMuv8YSy
xhZoyPJZZ52pBtq40BYtWWAmDiB4S0pmg2YI6cPE0ZbGFAQnQu2Qiza2x7GLU4ou6FFifaUk5jvO
rD0X1kqzmhSDPtfScngkZYGwSNF7LM077Yz4bDozw0esXH+IZdZVbzQQaKRtLvluBBSCxy8znw3W
rFDG7dVCITjy01L8Z90Ge082TtrDH10by4+O7iElk8jIARsyZhCGTJLDqTsFFqx0PZ90lJZri9fy
sKeWzBLooJ4oNxOZK9fVBA0ng5boBUR3UJFAOxgSp2luD7pdDovg8707a/4wWjyyT8lGGPZuj3H6
jRsjX0tlTFB+Zla0TQkpFlYRWhP0bZNrb9y2FnPPalOm90dbx5dYThdcWE+HVwM/Ej9OwsVOnZde
0PlwNp9LClkWwfvpOeJBgAA4MaF2KHJ95NB5BhgbZzhe7fgs/WW9AFOY+ZVQObsa5I4jz0BTFqIW
UqRY7P/uJIQRJbapH1sjoSlvfydUrlTHs07o1W+V68XLea1PN8I2FG0bdZauYiIjv4q9EWEALsxA
iBpAF5R8njLBxOC8NQ3/j0srcatNHEWFKdvjZMDelfYVzk1j8yihvrW0zlnZFdo5a8zO6uPmL+B5
j4q4YFpq+UNOyMHSOI0yUErBQzpTvaWD7NZlJh8h02EaLtqB0rT0vXlivEhf9KrZ3bd9JkBhbqvK
XnIkWPRAPopIebE67AOL7Wwfaabuo+L5mYBrgldqLQ4ceVjuMRjwxZs0dOCquW+hLmnUfa6oVNZK
XKzerb6sBMk5YF7NI425TKWKqqoQcprbpuz328/lnlTlBOfGz03qbp0ECZd3j8OP4BFOb/OLkL/A
MYJy7Umqzt5TC0OX65Ds9OMu0O8WDQ0WOf3bRhUuNy9huOnkP/3c7OisMZX4h3wI4WWpU9xEJikG
RMizhSdl83Wr400FL+6db+5SieMPMs747U1HHUKbbGx4iQCNr/TU73yJWJ2thSduzYUwOvw6iKT7
2aRBwzB7H0Tfb1TJ0lObmv9GkAj0KYMoSCgdY9pXV8HAX4MlpD+Wj1lBeJ20ccWVuya5r0mchB/l
7XRYATUD57o2ALy+TrnjvHqXHq/J0LxiogaT1hyZc4qdvVPGOugFfmRTymb8wbBP4bqv+n3DPhSF
/QFwarbhc2Uf6aOMNdNE5+HBkIEhv6YeDTWKjNJf6eV3dYQ/COpSQ8C92QsKi0HnK47jQwMcLyJY
r6D/am4T1NLYR3e/MavOxJOheSY9JYH2lMYS8ROwt6gBAJt2KGsvjGvAwnxQzCeQmcYEK/eUJC1a
9eMA09CzkN/rumeJ9KB8W5Z8QbBXvzZFRe5gheDPaugZKwp1lOG107BBr9Mdhwo7b3h7IIecEqqP
ho0oJOzV94/TRjdKFspeI4UGJPkzNT4KUwzJAWUm8kmp4ggq8aERXmB8Nw/xSZ8Cpka16nx0Te/F
BCcl2mD0M1zdKcKPMwz9uN7KRacxxLaoYeT07uO1r6PanBWPvA5GnFEZ+6Xt2AIpKd/0KeW8UD4D
HYweE1Eh9lanbPCoa+d8xeWprMlO1a7nJpS3/ZSzupkovcPJISs5Pqxx+hZHiKZLVW9vcomhextI
9+ln8GBX4W7NJcKuYHbHgowcTvZecmFVDUM9nzw23Od+ykWobhZM0f6n68Ran2l+8ZVnMRp/kBcz
OXbyidHvt/73bDtcV6b/2dc59ngSCyM7j4Q5jc4KFzwi6oc+jWz3RMivTN3hPFf450UKP3HLJQLX
R7VXbYDbk0IIaVUJ4FxKAZd5kBsY2lNxnvgMr53F9AcwaEYAz42ycevW6ZyMJAf+GIhio6kK/ngt
TplhEwrZP6SWSjcMjUHXquzjYI8mlpeFgsVWr4uD6PFwa0ultD8Zb/Q/8O3rz2PGgAQtZP0SkxEP
t2TAX2HnsQu7HYv1QWfHEmkcG+gLSqyy6p24OzsnEWKEI05spzxOG6w+eKC+EwzjxVZaEtFMbYWO
l1YKU6tXSqjRQ/dDGPV5Aem0Uf5GnjTfZmgYIOQsOOyzujr2dRfDPJmkllR+/SUeVon012Z2pVFs
N+Xv4AgBq8VQrIjQ2Mt3bjoqcK+XiK/zJQdVq/54EKlUBgOyuAahc4NMOjp5uu9yVEytOq3BZNwS
4dYwOAeO8xuUc0lVBb2SpsbugpMWP0nTFmhnNSCroYO9NAhaP2igPS0chsoUat9RJSdC9llZJpAd
Atf99wksrSq82McanCNp3L5LHQC9NY0ViTY8GIEhVtxnrYjAycz2KzU3gUcvuvZcXVdTTOB2wNiA
zBwZYGmGSw+GihydEFiz4vy+gwijLtiRN/xLRK16LF66BOKTqqyCyGqzcq7nasawYBxDuwlpA8qm
8PG337sTj1ndfZdQOosyfrOkP7ollKw40DrCLUwm4+z0kyAxfXTX0yZLxMVa3cbX0t9wCwWNeWkh
X7vJpQn1Y2nUWGX/gwNtWqnDg8sOc5uWm5dEf6pHuiVDcUyDsCVByGdt4QsQZLC+JN/5jv5/O/KS
Mn9Rrh1mK9109tRp94gZ+GF4CBGu7GKkTpBVnkYhmlXjCY28QpsFyUGrJKAjQLk42DeqRpRvIumZ
Pp+xeEMyc9VEMC2GaMQZ7VPPxYNMqJnZYG5QISU9xWnVZmnzVaoMVSUaf+dzTMg1rjK5ePihFH0t
n5FqOucA4HrAG0Ewtm9Yk8M/SqucXGDZA2C+349tK/AVc8Y5CPLRx/NgAMGqBzGt6iMgqoNTpWyn
Yyx3oBMXf0tvCKz4qtXcQF4CHYyRV9ntnBQlVG7mDJL46JjYQXPoCPvuTo0tqDNeeLmiS+rvgAj/
+pO8UZMcCMIHMSBJH3MpicmdOfzdYQ87K9qA+JjgLhJyW9JS2UY5J3d0lRR/zSL/XIyr9sJSuvtu
/gad3yQLGtn/0XfcX5LBBO9cG1uZ2ok5qe9aqrxqzMn/3/k7NRVxWGer+1o9XXpted2nsiKeaEwH
Ok4r33aKwkHp5CkS+6DZKlv6ErRW2lOGej1DaBoATCWoYLRL/hhaidaVrpgRMDkE1UsiXSGFU2YA
iA29DmX2SE6W0g3KAvbqp05fLik3JZYsbBeMFNsYbcnfIUGsEYAhUpeUbDN4r5wWqkjMr7MUpiK/
UV7reBLC5VN9YAD9zxHyIb6tTSpUTRmLvLNUDTTpXFzUQChb36kNalq+RwEI4xE7BzOaxX/8UZ0z
KTvotZrj4h0/+K5yjH0NE/U8o+0w+J7Wgl4DHaQorOWeyxG93ezjKIIV1ingHasKvPP3TA/yDf4c
MKapSQPgWpJoq0yN5q6eFaknvBFQ5AEm6avIS9HWQcgIEMNPm4EqhmkiIhF0Ftfll2cNG9TQmmy+
GdX1ZEAjMfjRhLWk69RhxxM4dLB78mehc2SsnlXUfwFCrfzPpuC77FmxUmgOY1RMRHst2Fd+Vd7w
uUQpO2h1dHp/WafP4x5DdOVGZhfx1bpOe5gPT9Fu0Px92RufIdG1qY4XA/tGTDQV9Paho8nc6q2R
GyIAke2HHrjtxI4Qd4LvQUesEkX1o6kBTx0u8t1ksJtrDrF/kR7FmoVKZTy1zaPNpeuobWfVw49p
Q4PEE9eS6dRiuefeknTyhFrb8DtFIZB+Br+OKApfh+VI09zYSiwc5gI8v9ZLOfjfwVzG71btLQaV
LqnHjCMukt7uc1mG7gmdtpTzTD9nyCjmlZCbL8Z+iTN8m7wDme+CqpwZjtqipGDiJFF7KZs1HU73
vqe0edjLgeTLbOolk6cdakLQH8PN+VWWy+ZlkhlFnE/Ustmpfs98BhqcdWFYvBbRjvsGWAAK4MCh
nAMz1Cxc4rXG1tLhBX8wg8Hv99l+pxSQq+Fg8tiageEl18T712+o+pE4da+PkbzzoDD3vaZpvRC/
BsL4rAlaCj0Sm856abSBHZN6F4AxV5Q9YHAnr+FmoUgTDdwP63Q2lBDvxoDGwD+K84lifgOrn76q
6C5G3XrBejagsGLsG1bfQO9NJr3FEOwvcL43XXnNnUFpWgRqE1kdcfoIhOq/lfWDhzSE9RRN6psK
S2TjHmf3BmAqTAOp9Zgp/nGcds2Hi/lCuSIFzxwQhAnjj0uoTrHlZVEZvUSj9Jk6XqeHw4xpQ+66
mvDDeTybPZAaIJaqbEr9vEMysN5hq5THzW2gKJxE2hGNSvTDuYvtLGENpb5vwqbFDp5TfjM+5pHj
eCuT52BjZT0bx8iv0PKCCO06xYcMwVzdbTqkR6Z2brQvqg1gbOUipJ6F2SQayw1oeE0t54usRzdA
KqqOfwGqyny6FWtYXzNsOJO7DNBhkNGBgupdEIEiZVeYSAUKNgQG5zDk0NdGc2VGGyZc3Cs/ShSe
LBXe2wik/vhvkenyddY7Fb9La00prrtmYKwmShcvJO92+El4wsUUKTScEYEiyIBg36zLNRAZa+XF
NmZFs1gbMaJ1jmMfyhO1v82FU+Xq+NS3HHRgX4JSGZdSNH9W+T4iQP9kxPdTWdRIeTsplUUxjLAN
dN7g45D/TaEp237CiXW7kD2R5bLN92u6t2Wi2Z9Bkr71xZR2Ve8tSqnvjNey4lXmxSfXgo2aCQlg
prO30xgDP3fi4RxuvuJdj8Xy9a6wZgpi4gjWbnXsDz+ZkFdZpHgTVeulIJzr+0/jlcQTKKu2AS82
uQhUUWMfCEiJAqR0aSW1OhJFqTbjI0jqluOqey2b2ZtdQQKmP2Ua56BwsuGSoifULwiytczQfXIk
9HISp5o3rPJeSZq1y+jT1R11zVThLf/Opmy06Btb9Dn2B5l5Cu+rvDPiuwK6ENj9Cw9f9ZEzW8gL
w7pdXyH+ptDyY0IXXueSNnO9aq4qD7zuG2x60v/Ay/L0A1DODkV9eAX52Ohc4hdZTYH7uur40OHT
06QJn5TWGnU0oN7CGn/rveugnHtQSf3u6Qby+mTgbGwRu8Z3UXXFDRIFEu1bpNf82WTmJtqGFLjU
VhCd2ZEIM/02cdvApHBKnHyGgsbUV6/3uTMYxujyLzSB1Dp3o6H/uyX22gjqu+vEAuKrwj1bu1bj
VCOgkyq7OOvnmLdAgpsu86p713K8Web3rrjrGja+oK5r9rb0RZhUXg9ZfyXEWFmVgBXejP65tenS
3qOB1ZRwCOurUXYHc2VN/SZn65zioiGmOo7kHrFY8MZf+2bvZpUsMf2bMFgLC3vY04uleQsesMHz
4ItYX+Tj7p88Q3Y4CQRuWZG8aZkG0j996fN8xUR+clmlXXKTFh1Aps8Mh9zkJatt+28c8EPSms16
Ic+crvARW1mnaaoBknYmMHrR5jkJbnoqfxw/sDneAb3SkmrvMqqq9Z+7i8OjW4vH5WDVFcVa/t1+
fINIw2b3uZXaV0k1qISMicaZ6t9LenIzxm8T9aTlg/lUQ8amvB8Q0qPpkjWniqjGioN9giE3CPXf
X12ZFlSwxqi4B/H73YJER2ptdbcl8gYPid1CSBLhuIZTN9fAiivZakrr9sLGNi8rAn2LcMiKEcAp
QgyIX4YZdbQ8rZlyCl9CoDEw8AlqLk6D/otKCRpZu8A5cWxLtutb+fyg9YZOOtrCy8woMjUV6NIB
zm47BLrZ/bkHHOQaSAW/u90cc6gp5VAnSdbNQ2KS9hCJCZuPIEv2xSq6NFlFyRx65oxSioagekQh
IqHqLOFQK9geTWpiNHyLzBnXZLGfnPXHsU7HrOm6jlW+IGnsfZV1OMrrGyt99efXMMguqO02G+R7
Y0kbY2Qwhn1SVWQNRg/+H0IHjzIBtSIi/Op/EmUpl0DSU8jkVtChTiz75tgdMRU3Nf2uF2fvm1EQ
15/saTQiObIYMg15IUPyHLgKcbsDWIVKg9800ckPjz7NwEhO4CwZeorbEdzQgNQPeR7a8zeh3Yon
L0PaJNKAd586C2hhr1jrK5e3Rd0BdU21kSpHhL3qGfh3+/UbVg62o1GsSGcbhhbJozSKxYB6fBan
m1hzSFdmofKkGubV7yLkgYw3jy3L3ugA/6mNsYPStJUL3p9sPZdhoAMMTXAO3SjBVG8psm4HgsTR
2o9ysFmDD6cH5YZ4R8XZ39fjJI5ngY7C/adP8pdkbEoXjXsjh6jADL8GnZaYo1cp8B9FKnJE4J0/
0PXIDP3Vj3Rn7gJ2vaex6azLpJ33c6JRyAvosbvIzEbhUlDNsaRYPdX4MukznmAKJeiMUBqm5CG8
+1T4XEMTHpYkqwLYF31JxJ2RJvcUo2CdAVbLd6B193c5xHnukF+PgaQjAX9kO0UBlTnAAmbmeSsa
+XxrH8a5ZvqbNduC/nS422QQrIk6dbJtv6CmyfvPSPBaOHTPK/ZzBUtT0Ij5LD3TL+1SKLitfMAJ
edregs01lyBqu2l1KjLrNQbjGaCRjxzERhn24ceYLugpgoPrIR06gQ04IAV64+/sOg4lqD2qW7wo
iMzi0USPNpA8ZwrSSSphLFASG+Zi7NuaQAM9/J+F9yNRCzpkUzTRNfB3DGrtoJkOjyLG/3WEVZJt
KRwMP8SCjZm8KyvxOffz8EnZOUqeWMZXiUMKBkSoiaijNktUMokPgBs6AZfByC6J6YsO/1iYf+OX
xYwihL9onDDTr5OyYfToFdGycn7U6Gq3QDoOy9PtGB2H3y6PrrFoKfCtqQKAmxfFJzHsT4HCFhl4
fwOqxl+Bt5lAf/YNafT0tCMT47jiqP3nrttbzDk8Zs6d053zEzDkT6cLOrcLQs/65oMsp7FQlSNk
YssLXNJ9Z0rT+IcI8O5muGNk12DfWjmLbtdLiLx37mc5pQi4Cvdxo3QSPRFx/0IoUeZv+4KPQSue
Tlkhf3m+rSi3h27KzJyfrknQPkxN3aMimY/QzfiBTeTm9/2IlkqC1PzXCaR4mXqbd3hY5miOoyIk
P7NeFJtE0IFSLBiTpfOJ3WmMKQScfA+8qlbDikeR8eHZosBDRHLXO/sH04tqUaN/kfyoe6zejdew
s0vE787m4s8mt+YXX8YnUPCWZpWHuwVB4UHqvBoOT5LItdXA0wE1m8y+c8GtaEA7zrfIsizV0gaq
ccHxvUJaRNxQB/CqT8LM5z1jkE1rp3R1USd3jYdW+ZteLdP6ZWSxh72n+5xdd+uO+iMvjjRis5vx
Bk262tVS7HXa8Jn9uZZpOnUkCKZGlEx8958ig/ai84fCTX7+4Oq/GcbmPpOGVDW8xPY93ZTSBMhp
BMzm0XkrOhgl+jD/Lb0jcS7j2MIkrAMQBIjyOlmSVQXLX6uoBBXr/hWXlU7XE5j4+v1mYLQroQSu
2W11TBk8G6GkUcMgPhcsmmSzAnItfUuwbC9Z7Qdozvi+eZhtbC+fqOrzD8byQIMPDMGs9BicD9ud
o8KCng0BGZ9rp4tFNt2AuXC+8Ln37rMCgu/wy+bucxPm/th7KFkz1PEtwQJ/iuRt7RNkXIJaeXhT
odJFiWC8mYDXpiYB8UGP1Xgn53wo7JsvA4MY0AmynJ5MsUgJgc5TUwNT6TE/Vgtc9gh13hlj6oty
Q+iOA1R411hmHK1o/Uq8Jy21DCdidJj4qHt9cXrS+FzFWhYtjgfHIoctYqXUkZOCquPSv0adE3Pr
kJqD/Fkg6a0WtDYSKYuMZc4JGiOTmfseaIj5MMH8kiQxxP1tyarlcGrxzVUrZkERaOyds3GXYMNq
hujrq3E0ituhqBnD8EMsyUbfufg34gQWEqAgB+asJyWa9bg96PHYVkNKHQ6dS6FwKLbMSUqHbpdF
sbAEIQ1oriAAbx34QCr2u3C0+lPXOwfv2yAPcpJq7pUBijvmZzXhRxodU4KLO5lvQ3ZqAJH1oz9f
kIlCsRAx5BoUMQlH6XVFWS2/NfpVkFEOE7+CoekWNv2srgENdVti7R+zt13lvE2bKMrVbnvWs633
Zao7BwxFU7q8159f0yvPiQlLUAFrB/o7PQo0RSlEoyONMAggZ+AcFGF4vq62cMTHYxdBgbj2F8x2
tXRokrKgZWpTpm/i3i87Sq8HxWn+Hq/nsl0M0SXHRAGcUor/lGgtnqByjrz8FJRjQ7+M+osA01z0
2tq7gyku1cada+vZVhwWpuRXTlhrqR73RmsZDFT+uGt6exuUqPg9XRWCNyJS9lK4PeFkh4QY+8Ob
IJbRcAqdNTwyy7Oa8JCBIGuA3Xr+NkqDIn9K0BpaVWhBcN223iyirMOs9DZTMIpbN2rjiTxJN4rb
q95KnLuy0CUGxHQs/1k1CaX6zIMmT/w0xdvEgFq1zwDshKhSHJT7wnj4MJTNYkzEkIx+6vaXVXZt
NzACj/AxuKLSwB+45qlvQCvhOUsk6tGxC0EvVRQTR1iDN0MarA81a761i4JDEoCLXRhG9ngxq1Ny
6xPfSX5cb2iWXsL7ZhOkaNRDknUFOK8M/5SxjAWJWhTWpAGAW19SU19QcGVpAJMSgFeabfOgl2UM
CTN+ThXAQnmfwcM9DjhIpzqS2VeLRP4Bg3L97hhqcXIlgho53HKoadUR6r9Fn/0YR6kDZUOwAGX7
vrCyVgy0aefNZm0B9/ohX2Wfktgdmd+CEX85J9MMLDSE7fnRlVBBc5/cR+NoCkYUwVGE8SDmLiIb
8cMcir7KTaDHi9nWyGt0Cctc8/Lv7XRde9HVPHzM/9lDQQwoAT79vpR2WjNHoP9EAFiOM1bVIUSw
oqb/9CYkhtaxO1dQd9iKAeHIXpHgpvQTpqjwKi/PSNnknAcAUrul2FHaw94UAQMrwxzdTyElMNuz
dbLX0X8YMv03AbfhftnCEmPAQ1ps88g2HxJK6ql8fRm/inzzhuyV/bv3W1XqzPzb79urm2jk3NUT
aH7NZpKl8K0pC12oQm82KAGyrPRqYlZeV8WsbA7ev5L1osFW2xQU+8ap1l0rJycZ1zlUGJJ+y42e
ts6qSqoOtdtBlw1rcBDnyTxdvh9JtZMB5do900o+CofwNuhstqosq42Zuv5Gl2H/N1xiVvet7VXv
P/N/2HRh1OOamud3u/1L/5JoB9RQj+irqXjF7WMeImp/FqlArSfRu0+G33jChDW416H36+FqMdMd
rljYJ14wPw71arvlcNn2t1CCEHM6XG158t5fyXTIXKeCEcfEOjYIJIQ6/lh4Ps7lgKKl6Fj/W6ue
/AVaOp8idMPWVKTzcpQz/RJPuJ7uGVIJL+14AHtMvgbcUvznLP6NxvpUZDBoOT/u1kj8IR73Lwmg
1PTSlABlrt819JvLI3KZZrqJfO/FUt8IIUoVhubKrW2wMFo+F8efjHTfoMCuqkSNTZ+qVl511OmL
kAaQSiU+51+UFVfCVFAOVm+4MeTnIDu5km/e64QCxaRvgstyI2qcPYxP434ShN6D/9tb6Fq6rrK4
Ews+bbzAiMPWFJihpj6F89fTsISa0fiJfEhXfW5FWd5FsbVAYJghtv4A6X+tPTASwo1AigzMUHhf
UD5OsQNZLqePTJkoGfbUyLfd2fMApFC8FvdyCFkLaZru+fGpI5EVHMTFFeeCRAWxD+wrXLs5MJee
TGwDcEUWYnF7KEjCUmTFs4q5s0ni0bjcKP+LtmBD6ES3QyI49fG+0nq4oudtKwoNJ10c1/tKW8Ie
TsNP89afPCKJeZFvndzwthljlN2wu4Vg1vypURtDWoeuFbwyx6EPqsPrOZasXEDRk9yB3s8tTR+c
T5vgxra1v/sf2NJtv5D/IoDZNk/UuDnOesfsT5y61ay8l1hy8IuSMeiixMK/+ozc4tu2PONIcMid
9FAgHUfc+xZbqusnxjdptsp0GbRs8uip3RGDkG9+gMeNOHBEtb3nJtzfJGfu5o79M4LR5N7ZAvO0
QaH2QR13O3M55Ym9OtRV0E3SWrmr28n4ic8LL3Rv1E3mbaIDXfxq3jP8cILs45cfkCy9BZbU50EN
90ixk/wUsL4pstx49lortdcTCtn3Y3kHLOVlqxNwTsdHCDD1ngPbvw555XiUx4xen3OcdHHWESQU
Bw59w0kdJxgJCKYtilxy032WiqyVSrCbpnPEuwq+/nSLZymE6VD8Z51s3MQHxxWHxHLYw9hqDuQA
WoRZin8/6I0bBBpGqMeHYmP+2wWyih7eeDSv7YZxN7Tqe8YVKsFh53oT5RtkNttntcjIej6joabE
TqhO3NKk8rjQImX2XkxC4ssA25ME8HssLAte3pntbrXSrWwzckbDIncZU6sCD2zAsOKmQJhrnbeW
rZ6F00HcNPZXstp6MyvTpIv+oEL5JfbBhoJrLqWHX56oHX0K/OYNg9QRwxaE2k3KM99j21V99t1Z
rVGAcPbXEPZpJ8LXVvsUZMvKrwEP8Af78B6o57AHJjJDP5zGwrMCWmzdXTTgPdeWEEQ7D6o2Cwn4
Gpr7MH5YszcWV123tDdCOIfqluS3lnfrcJHGMg/febkV8RpDtvVVjghoi0HKswK2y9KX7ACqpPKu
5+quIkowxU3e4RgjXZrn+YHL2HhNKfjQp2xfQzFEK/9ZlAK8dizabCCAfRCvHEvCh2YBB0aHx1B5
Tz1p8+c1jFW4g7BXesDctEpvUbendSteLfZifZimCMqgDHpr39rnORuZW/FmJ25PZRXmZBGNOvW9
ENsoh4gvBId0zR6C2EmMr9S9URq2q8KSai02e+szNNoXwmnR+pt7LifvyADRtse0cZr9O2kc+0sn
8z5jOV1V+d9nNDRA2G9odTggvzvex4aVg1pN2R2wPdyZNZ5Tn/UA/8DYXcCqkA09ILP/ePGkUqJc
7nFA459vG/aBRmsCHDBLy+d8vh23qPLZ0nFTrprcnMXUW+Tmrg1D0J9W5RGgw3C44RDjiYMuTfD3
zpyWKDTYVzAUxmLn1MUu/hWbe9eSipQBpy2m3uUAlEnd01ELb214ulGbDmRrSjT44Lbz+zUcW3Me
g2mP5SMXHlf4pEG6TuwFFkFcox7nVPKK/uxK5l+tuFi7x4U5fqKrh/rtKuIQBc9FoyWs6MTttgQn
U33T8IybB7AOLJpf/24IC9J6T+KlxKvueC4FOuAUJIRr79gQ4mAp74ikfArVMcb3v19H72CHOoLx
02ijFQa1XFL9Etg5FiA+nIBAgiTer1h3WFbI0brpgG7V4mGX8sbXaMdEQ1VZeKNIWW1fCxiG5YLe
sdAGnvf4UkU9kYP69THY0YowXFAhwQN9rtLlmT7z4bQgeg723bJSTalvKNgDOaqk6Ocow1z8Ghw8
nILbLGC0LrMqejc/nBTm0Ws6eKyFc9R2DSuu1TmJj6/+RGoMA+K7WnkVkdxzTLCkQLOGvJk37MRE
nNMnHlJvh6+sDF9tHc2sxkq9s77mjUSmzxuAFY6dtr/9vcugFlLSu31Cb9Xj/wiBi1osbfCkmNe8
HaCRpMqrdXgUkRTOEYXsRYpErIhYWEwzpUKcW08J305kctDSdysLe7pBKS0EGr/BL6FZ1qMzS3d2
ReiQ70gcHm0Iv8t085CQIq9CNDk2GEC7qHXjuCRdHHG8EXQ8ZBdAHOoCZthuV4S5637eBwNlPwzA
FemZGlKe3aYcutUA+kDRLN0wmvE8A1W9YhtI1Q1IdRSBj6Q2184yLAs1PsEl/nu7HhTwEpt2FGOO
qv+dvkYNw3T7ckzEg1mdUFXUZ4E8gk6RFq4cOrzITM5SORH4zfjYGiQ0FQKYhWbUrX1hOmgT9ebP
Hok/g0BM9fOgnOMOBjtozY7uQzpABKY+jW/vB5h7Rk+q0Skky3/TVwfn+vbKsZbnYF5oL1qpe28r
H3Ov8zas8CE0+krBvVLfq5L6XLXGL8+YthkJxAj/bZU7oqdHUZ0e2YLzJCZYHR6YH4Fy8RLNiqLM
0KeooZVvoh/m24o1obB/VkSQsoJpbRKBezXM/HJCJwhWSSYJJncgWH+w1v750d9bQJQWBYbW9Mq1
KWAM+4vaPZ4F3WXvhj73F4JUoiP8xBWoT7pVx4yvQMMOI8tPmVWsgdpefkcsLZmXrcr5M4OM26xC
8RZqUdoXdtOzkKGnj6ba4Xi6PK+eHUfoXDESvWAUcmi7D70PB4f0Mm774be8EtAlS5XmCj7Mryp1
jKjKWehvwMzApscSSeqFndYKJ47nxdDYTlG2pX/LNbWiWy1CIzF1Uy0svmReQHiEGt7fA3sdsBfX
MeNhpwe0y1qliscAr8eCUZ9BiPcTFW0qyYDOn6Us/qeNnmoq1qYtJxANRu/VH4/BxYLRAC84TCVi
lYLaDBjbRU3fCy/wQ45d55MLJHFHkcV4ZlGICfi/IA16NZEqa5Yim8e0kT86U/aUAV0oKdRmamXj
lUgB4t3H3tevDzeWbN4hYs+iv07zjuvj3UdB72UHsdUt8chUQP+jPBG2zSlJY6gJaMWzDrNRV1QM
qC/2PEv2O+js4Xs74YR9sQ/GqBSAt4i9cRqIBnG7qKQorIxYcImFH6r93GXWqpbX2/fPoogaaGzF
mqBW8qtA7zvJt5c+HxKPYjAHwlwqg8maV1ktCJJDaSz6IkhZn4hsQIiu9HpZ+gbyAd9/Ymm1zmN8
1o3G+lN6H/YmxawmTn2JDozY1GdA1tbgiKpaLd4vlD8EI/EZRtO83Xs0qkMYApYHEBqp65d/vFNV
0i4HX35Ib0WIj88FNI4gZ18/DgsVUf4BkrBFoslhN/b0XHlviSGUmPpIsXWK4ddST3u2kcBsF84V
pmXxL022r3scGNO5RVzZLbUD5ZYDFWvmzffUDqr/jE3YkdwxQ1VCyg3YXBcIbzJz4PJX1bKfWjyb
Xf6P7GRxE8aj/JgKPXyGQBpIoN1J5EFVR48FfBc6QlXTQj26Ms6rBzMF4lVrGkHljDUXUrAf4jsq
e8hib8vACYnSySg6ifmR+RcpIELkrVmoIbHBn8+Ul1soNrNSbfeRR8MV0y6vubtW8usNZ4ikhkLa
wroKgT3TpJXrBpinXO1FLiAAgFT/HOlUAAvigAwqulXZnDvtS5d69MN6lzgD3ApUznzcMzHOHMl8
tRW6Ud+2Tk2lj6mcwW1kXbpndMe/bTdFquzqaRx9wmsjTas+dG9w+KJT4+fyFdA2seLSv9xDgJ+B
s9s8GN4LTboY1xZOHfHTs+39/p6p8vxoPdQiYqFRMhIZi/NHjJO0PBuDujGUCB+lyrvbFHhbH+cA
9pKaRfg9eKOJ7CqS6WG/Pmv/cGT9I4s1hn9dbtqhJlVP97GJX6DTZhqFhUu5C8XIgMcj8jDPNx1+
1rzXADVtCn0hvaH06knfhN75sWrc/0UxwSxm4lOhHtQblA2efemKyt+qUxhnfpa2wkvStx8T3Yvw
H1YS4B1NhSHuG1j8erXnAWJDVWohjybafrzd9G1u1frb24RY3geMcPNlEW1eFROZKTp+HhCZ7v2F
2TchMjYa06Tlxb0vOQnZG/gF8mZrB+euF0SiEQAD8G8wKO703wQBxiJeGCBCzPB1GRx/37USBcm/
ACr96h6dYExPgAxTkrg4V58GvX4IZi5dgvsrmuvZvnEW2r+7hMLHUhrqzZ/SUiWA7Uf40Tn1w9Bs
HIQR7FSVYPWxVrCFRhr5z6ITA8zFC7hU0Eg2kU1zCgzo/0vtwRKX7bnn+a6KF/GIJAsVQABd+ePG
CUcLmL9hEKngUaRnnYKgLyLGurxzZqzTcb8js+n6UP2ZbmMtBSXZieHb4ygIUbXegjs0sox5ym7x
6o3xvLapCHWaB8SKaE1X1MQkjg+PfDtImseG0xOTpCVAxpxyNUU8JEtj1kXXzabWxNeFozz93mVI
rN0zuem2Hb6Zm+CLmmRYGzPPEF+V0CugrEGtC51JDjvVhqL05nQLoECoUdEZfm+T2HErel02vxbE
Hb6LZQfHjOP4Fs0HQy6gU/9k9FYuOziiyJ59Cad4ow8pglwz7rr6/oFuz0JWv8oL9fY+i/WAaG96
g52WsRbkmG6jwC0eulslUUJ3S6iyuL8GtVkHxL3ndZ+IcRS5n3GYLPtu6ptPeQ/Nx+4ZGdq68GTt
rXEYcSFU5/9ZFKuTjRwJFlJcgYLegG0WojUbQMsY3Prze0eB06uFelIT2JrLcywIEZB49Il2TN6Z
nXwq4+xwMfMTwfQver/f9M0dSRNPKGVta0IsbaPKiBFjyqy9KMW0tHLQqs2CdSmj+rTj5BvlT6Ta
KojBrJ7ZyvRsG9ZM3ZCqsuOvait+PpW1egxLAcSZC634KnQaAXrz2FWEh7xegB+WePj/i6tq5ni0
KnyvCJxML6/2Tvg3i0Gtjih7oyzH1uFqxpytXBw+S1kP+F6IYOsmBsxXVJ7JZHVyzDn9kLBi6wHf
ZXQF3ERG5dAITHVRB3KIdZTe3kXE2bsUn5crc6oGqV7QBLterngLpw+zKvwYenVlcXSYauOhittl
q5VAy5Nd8RtCpjJBNemvzdHBCd+7St6uL8pkhia2THIpL6t1ziSsPWOs+R0upmdNGntQN55GYnes
iYJ8XJfRAl9hSH73ZZJXmxbkCR6wDKxp6l7tg5PLRECFysIeVIUj8ufm+8fFg89KHEym/x3xDSAT
pc4TUB3kh/Sxd/DWDtL423ZujU0bS7rJiUi7maR5KZZ2zsBo18KGI9YhYiwSqjslFE+CUFGZO4pQ
i4z72zCKJ+ZJKmZyTwzDjthQjV/mPR15qMWfmmezBhqBpBHN9hZTIzv3zt7Ln+7K1Ut5bVcckHrM
0tPhooWx1xyZ31UoI1zPJ5Mzj606IHcU4bQbXUDMSGz8kwyS0iC1EZkDSBKOmvfd62t8M9lU5xDF
eiBAqMfkamHSkem7I2r5av4XYr0cyPl7TpWThxBGQRQC7Ri+5zk1J2WNhE3DJdy7Y6uNjL1A7lKz
IKlJyos4Cucmm1SnNzvAJMg+aNETZMND8uwE3SrjiE6j4/kiSK7BU9KjfBV9tZOuzBTVjs7E8uu+
AlM4VEw8mJqmRq3brWMv5G06loqAJCZeOYsAqeIrGYDj7TSJP7nkR0T5p8OoHLwPP1nfryJvD+25
NOlHwfR0XhuCY6xPSYQ8fYgtGmj+DCcf5Gyj4hfslBcgJUoX5dLyui2n1bKaT2LsusiH9Eyytz3K
SwLYEDR9LM2yKFdgUUGdvoThkfUQn57FaISkl/dwypX/NYyZ4Gl+NwQ27ADuWbQIYk5M0JWj/33O
+jpGcy3jCiG8rKUUUg/0o2qDYueoAjUZi4evEZn6ryc3fxzqS1Y3GdiO0DI9MpB9gfDx4Ek/r1DL
CTyDpyessL+ijAuG+IlXq3lHdP+IJlCaWOev9sV+2tqpitu4J3P1rFJKtlWMwtaftpqDWBj3KZq9
MYHOtff9qhNDw0wwNGCZPIwnqtf5te9KuZICqNOD3inv9iuj52zhvPRb9f5/MufKAL6pKqRyDmvt
t8CAnuygEVnklsdSsap76ynJ5BYVwy4RTx8XKINpuDGbXcQGvYv6wjnfYgl9l3reFjzPo0AlKllV
TAifas03PF50ZYhqtIAo2g5/ytDuQwSJ6r33aJbBvfyp0scXFCYl6LmZYbJ94siR3C0pONJGCKv5
byYozHOdyXuBXh7RjzGUjgfMLZ6MFwHw2gFr8H48qtSPIztxZpLTodONaj4wLPil7bw01zfz54Zu
kD8wf6R6W4rU2C+k9s8OcAwik8ot2DE5lILOFaAC27qOuqMWX69hdy6c57rCbEOhWR4ZUTPh7tmh
Or6Jg/cBi+S1+UeDwR1cjWVtUaSiaTrzc9uTW/s6hxupBn0tLrRgQEElg0o+6jHYF5OSMHfFKxZP
aByEnttQXuLQOIfMsMdD6H/V6NrkQxbJvKywsNYlYcr8taFTM3Z0sLhjHOPjMNhM9b23c6gE1cdP
cEowuoBVz34hamjWwdguvMNcAvDm4tXPbOH0PiNWeoEuvYSz6/T46+xRh4CqtxseZfMBA2MiduB9
lUlWs9MCkzm28rgQ4r78jIrX/NUO/nM+fhd+LedNE6mbFGo5/h7rtP75ABDXe5OHXTkB6+zjHOtw
Q0ZmS2wrcZwdCPq6tpD9AemZeFQroDGa15dEGqI7MxcUD98jaNLEYsfLrlZAcWiJxm6pChfgJHW5
BVWd4bF1AF4zIoOgDojTox9wvutv3Euc01InZgydtJmVx9pidCJ8cwUG8vbwYSxYv7HNXeR3jPcg
zxHzMk5ld4Wd09HGVyAjUl4ydKTaewmbpUEBVqdKh8VsLZrqUMjWrrLPTg7wwpvpQRCpaYrunUSr
kFbVLlgz+L7m+gXjCxZ7pkkPFKGsUh0dPtoWC3fHAhUG1oj5l5yZ11dY0nPC2IWiHPOOp8tz2OIn
3kzcZp4HFZgZt4M4elz4LBwsvIlBYAdAUtLfYkV4Uf3k1CxO1Xo3sRlmyZCaKrosigZ9D29FHhEp
gJRXlFDMGsamS6cHbyqe3epdMOkWjFdUKR71VY7xdzTjug/fLyaiqMfbAl6QQvN/SN1CzQUGTmqo
xzZu8BmH6pje9QS7Ldpv5yj4vCo35YxqfI7c9hWda0n3GSMVAGKJV+EoqT3H9/yzuRQ2lDudnnDu
8DZ2CcwLwGZBCw1H+mxmrf+m9JMdQ3iyqTszrv5I2trKI49vWfICyiUKfDWY8qSP4wR7j/ohbm3c
Q170RzCf8SS8hTbPADTwbs8pxjsfskwRSXp1isKx4AOcIqteWq1k1rHoC8OM5IilneVFtxo/IYsO
tCnknmWdj6dJj09mQoKZ2Z1T7/AFL7bt7uW/VHqAowmlmcSCw5Cm2aSKYskwjDoA9NqoPz5+dFAw
lTVYA/7Rl9WMk1JgU8dChyvk/WE1wfU4y8NQPtmieth7nTTYuyMABINa6mT/ZiCDTVgGLZGlYSP2
MktFy23a+jomA2gUNK4OoUx7kfx2jTUzlQ0dgk5yk6Ud9ytXoVG9VEGK2XCxjB8Sq61UiC7dMDmT
ltrRiRoat0PhSoBwtovfEB15y2SIHPwosaB6yI9A1tK6Vy82nAbL/ewtR1FZ83LKSoRZp3qpx7mi
i+nVt4x32LmKLPqrhNzwB2VX+aHmkBtlOyaphYBs8vLTqko2LFLPM9vyHWAsby8rViGA1PmhA4Bf
9NMF+nZ11+ja0spDICT6sGpnd2IqmtsHar+gKZ8QGSPwnm4ShQUYEG9QMJz5lmPVMUHAhbsc4LOF
PUhTyY71oecw0lF62MFVPqb7sEPBaIlB0qYF1pqpVFLw5TqR2EBtJVQi2jcU+9Ddrvh652Gs0+HX
Tt9S0VWQC6nd560iSmr820V06HS9TvAJqo2Wu2x4jiJ1KxWRQvW+GMWb4LokXZK6hdm/ohh7ykIZ
s7NmAyiPIJOd+5HE0HN0FjbhwTk3hx5G+1Nflzt7ejXY4M0buBayPhNmLeq3eghc2zVzt3fFJ1gs
IcRHzz76XWTby3J307WZSEddfBFVn8/QqaFDT2wH0PZcN91OaA3T27ABenwnaXSB0bfzAQ0Rvm3+
bl6C6zdtjO/FhOJt886TuTHMt8W0avd4aMILFUddKLFSb6lWFuYU6JGAsY4/QCm4/xZUbLrmCK+6
vi2C5H1jhTTgs603Oa51R3TYTHwxt77/ihzFa/l9nKTHCOBVauyQb/p3Fq62Ut1CqKrjUwERmto+
PWvJCGs9avVGa0lZjmzfXXhRTcZQktNQVKHtpsX2wFBGGTUKTjp46UWGBSytOvs5e8cZWkGWLg5G
b1kX6OSJP5nHboED9s0J8sMpMkyzkTTtbPMVCpj+BcQmUu8nwt/KevOlsAhusF7EaRZ6rNEK4Udc
p4vcfwREEg/1ktCGBcr0ePBzAkcHd+5vIiT1tMCYC5MYYSidAeO7ODwGircrj+6uF8S5VsBBMKpU
AwjcS1OrCYG5Xp5Q4bVGTWd8XNC2IfAf+j3njFAHUcngxbQ7NB7GjbKTP0ckAwLrnn+uiP6szvJW
aIaCSKBMRiq1kc7bm059WThlA5gk1pb3g68mFPrHt/GUJe+vL+u6RYh0ETdzfQNpgK0FcafK1s6x
U9fakobOwpVs59vsBhw6j2Ac92cIQK5xCekVYYJx0n1BcnP5YYsbFTsYh0UjfnWF5P5U2SP1K5qT
V0KSytIoE7A5CwQvH2Y4Go6IWNOCPcPjf4CBpcSDdiw49L89+ZaZ+BOpVCHrQO+HOgZmfIhPszBs
wo/A9pshYWRpd5p1fSPKV3C4q9Pter8XkMaLRgAvuSSspX3/Ywmt3vdlDUHicnLMhgmCOzry9YHj
f3f17C7jIj6CDwSq+FckDyHgMMDBv18I+eLp4nAEU+FnPkL6ZSTxDlu1asNZ/5Zj13/aeSXz3+r2
dG3q21N1gK+fw8U/v1IjecaTZjujfZ3oZJrxHmf+vk9sIA2UoZZisf5xDJccMdGb0jLjjI78rBEc
Jqnj0lzi96EhHNjdTpLhZkBc5G2uirvDkr53NzkTScVZwgiOzOMVqVY67/essF9FqZo+4vkilbzq
9S8URjjMfWRp00jlUkebXVOHSCYlK4aPIup+b/G7trRn0S/Gf9QQYx12uxM/C2OcLBIMVnb1oNiA
kzsBlJmDkYW1pdIDNdPF40wgGzl7QMEo8lbqGJ93jYAs4iTaipYIUBfWYQCwC3HZy2zIsyKUMHSQ
5im7gebWIurXwNzKo9zuMp1e/AgZbXdvsph7PyzgNIFKKED/wAMMz8qGZTyso1YqjVVO838ng4xZ
nZ1bHm3IgTO9K/Ge88BO27gpAo7WoAflShNGbR8USSus0Sd9uNh7bYjQnwxR+a+jobyfGczOQuBU
0RgBIJXL8JdW8Z4L8r/mUjFNV9tazM2tPU1fX1EzMm1rDxwyFouXLvgjRJIbakNOGj31bKpTf6ud
pp9/vs1VsxpgPqBI30uR34gQG9S5y4byGC0Xlo61nR4GWwhQjg46m/pmv1PXVtYchqMCz+Hw3ZFG
m+O7dXaWqZiyFEJ6KYF/kfl7xI7vUllATDZzeQyDYJgBzuPUDRL+im1rz5uVq2k+EXuyEI/7S1Xx
9SSPFs6Gv66jyVgKlxzNZ8rVFFg64S37GsCtLTyYX5iOgd9nw0iqa9NoPms+d2+H53cwV7bwVkNx
K8ML/b8Wl6cbmphbmcoNHakiLurym49d2macCE4/R3hBk9xJA6tPHT2cWtPi/BgNm4glv6ze/ZzC
Jsa4b4E3njJ1tCxgmt/0j7xw4BF9C/DQgYR/hoVH0SM2ndX7ku57oBB8O0qV++eQ3N39xi6Z5SHv
Ll07myamG/gNiv2Qwgs48u0/3eCuoouluIJro1UZoeua12s3Yi8LF4Cvji9VjzWVXaUHtXgFb1Ak
pzBJZh3TEF4AP6VIl0jkSwcGEtHSSEovXVSl6pGYwjQHLvVu1EsutAak+/7Iwxt+MSqIR2CIBl/d
1/+d75rVe35TTBcpbdusmGCZ/WWm4ghJKpt8WOYWHMSIDClgcbN1ubaCYQM56of6YrOzk0hklKRh
K7hC3xtVUPkE59gimAXYqlJaxaEhKvWCkggH5d0RclJoAmWlL5y96A9vRF2xa4+/qX98+436/Q0u
kio633xM32b7HV3lYEEuWU1vijXJ163AVIFZVWrVh0ttdKdKsKKOqg82rsHzrigeT20vz47v4qCv
bWgg7MRfLb0Yqh0sHOJFN1/mFjm4wuaTz4G+3pi5S5T8Rr6iC+X7VPArnbHHlpADpC1AqIxYfuXm
K7Ipan2AQKAIWklTNeU8FsNZOn2229IAo/3INfkGZuaIsTD3+UvcqniRhYhcs+gRsxr1eKPZJRa5
hAsdafpoDB3UF3rLmUqRs81IxpA00vosOxlMFkw2Pe49rlm5TmtkD0xaJ7jdpmOO6aP2WEBh1aiE
kAw6SVzDBEHdP6qEqAot8GPsluaeaz7hWcgIHXCSpF2cbhwiD5XWVAhviBGok0DybZ1QE3X0ECx+
U2IhIPxw7utp0h3AlC/0NDqPgzrGiJB/sNvn8hRDVsxfy6XOZSaxr1yb9Hii8i7pXOaqKh7jdPBB
jzWbj6v1X5Vyq4RrYK8L40dGiK/O2d5xES7yPYDaOJImxYvJbwTtyjjMl065LKTP81dtGyl+yi99
RWyO/xnwBQnlszEQLzlFu6I91GYb3mrZ23f4x8HaQCDj4kXzp+Bt3EvUh/dsHh+NHSx83dyTbflq
ejtqx/vtZgjhjtdGi06eWT1AaDUjscx2ErBxBHejdJsBl3ieIw3UgKq3FtMw7Q8zRcIzrnGISNCK
aGbYkMKHVBlUQ7u27MWtMPSMj6PKthu3Fp8/FYBBfXjemq2XiIlx0RV56B+m3tbSdP9ipLruq9x2
H+/EYOK35RBZ7ktbY5ZhiC7wT4VBnzeZWSkyE5yx2dGiXHawn4fMgcr1owllqb8CxsxV3lq8bNMh
qtbTVwZTkBMA9ccV6f32PlIYOINM286aZupnGOOkLO5Vj6L2JsWptvmm/ZLQgxguJK6P6unu97q/
/lywo7G7hnDLfnfLOSTKZ+zHVCFU+zTP8G4IkHzJudiUvIQEJDaZmxxvxXw1dpCBo29sCKYe/0m0
BMYDPQ0AmEPjxPQqCerF9QXj4Ktar8/YTUOPY1Xuu4rVwcof01GCD9yGDBluc/eGDVnNDYKYAQ9u
9McuYB2XruzIuLAHM8eYnXpwYofGBimhryBYXAP5szYoSm08y6LQHwxiG1CGOEYP0NciO12sKNV5
RfaEIGvH511IcXA6OhM4tHs01/qPdLqcIsTgwyifpsNYbgHBJpZ6XnLk0QFTrZRGNjXn4Np1Zjav
cCpHkD5dkr8/JmO7U0baBol4BZmoTGwLOSAJnb0ed23eC1oGu+CgUXoFFN8LQ8i7yNQSFOpC9I7X
wO89elXASyDPa2D5YutS+FYFGoJOUogk9XVPffJOT44ciGmWFikIZwwL9W+3canZX4DimYoLjiy5
4/AUCl9BkGeUsxpRliI1roG+9vUzT/rjVnVvj4bzglVGFJ53+Ol1W5NK3jpdAY6RVdD0u6MFT/hX
lKWoLRCYSADpONSGjvJ/DdmUt2Qby7GaeiuSApvyd7g6nT7VvHpcaXsPbhT+LznFChTrcdsvWk0I
1B4KVAnK2oZOgvZUkJuKgocHjpyW8etPwJ0cWj9ltXvrboSwHLwqrRh1uR1F/lEdiyhau5z1fdYL
fiAItZsOpyodfX2eNTlXN7LcpxDWZ0EGtgEKJkdxN8JtoUTgiKsD9xsPwnl1CIf+mSfQYG/14E/b
OzjCC2sdgJPRa5fkEMFwtODzApmeeU8dUx0MaiPO5JG4nnP99Sl0mUemX4/3hagKrjN8wtKlahiy
m5FEuvl+pEHs6WGvYtGx+wl6gIxelFpQxdEn+M01Np31GYrRzNZm6jDmzlPIojIhO8PCS2ueIMTX
53/wSuIgAyu8mKyZTxR2hqydeHY7aWvi+7AdEqpO9es1oj4j40uhl+CI2wYij8kY92kCTDLw28t/
fk9u8IXXNFi4w4ref8lgjHYSC4q83rcPLaSie8Ii2xk5P1Yq+LruTR63kgW5VklZcx71nvlDlU8X
Hu6Zf/V6Mmp29oAmfCHeAqSeKplnTyom5CuuGHeiPQ++tldFldPzIrrPoiqyhWYLLwba1g6Wumt7
tvUogacW7T/5WlHvyT/iYgnmoGSEpTy1GHGM4PFAYcUGwXbmb4OZL7XcfKdgYamtji7EwkuhepAz
E79hhDWOFZkyOU/UZbDXzklPcoyPPX553fQrL/WCJ3rQMxg/9p1uAxVVGGCYVV8uraKIxG0NHWAx
R2if8gRRz0mmqUidvIWXrJQ+k7yPczvVQVQYWhHwxFRK0SqDYcD3rOgejPctacMzCIao3Va4hhZc
qspAxhK1DKHRaAi36wirtNwcObtZ6lqXlWe/+k8Cn2qPjYvLy8LIymnRnyrqXmJcJuhS8CR97yHy
uY6+XTFf7DFhO1YHqGsUC/x3Jx56N0PUqsyfuYFBlA9G7yD9uWZNFBD4VVo3cHlq5q29jhTOTu2+
b/MxaQQdVak8d2l03fDipAjntP+wx5P8+Vs+s8Nl3iqicf/k9dlCM/lAUiEcW/08a5L4f2N0S96X
DPmS5JigV1WE3HWxKw9/RvjTr73xx5fN+G8S/7CCbFdPNgUJD2xmYxUGHqbqgat+NXzmnaKSSuhx
wXlkYeV4nrNDixnm/7YO1DzmXI4QIWPByYsZOKbuthII8d/QvSrHDgSV8m7OeSgaCpygjIOomAP+
pjMq0RUIz/QlJzRiIkd2P+rdBseVkYuq55R76KpE316JE91NuZDSkaj8jQUFU1rO79HhNJmY8HJl
UzT42yKu2S9b/QpiFcxi78cKC6JnQZI9F5KMeOThbT+sN6z7FI2du5m9RJZG0rmyLlET0OmZAL5G
DcB++G6klQORiJFPAdb+I5/I4Jziri2DB7ibI6CdSvYJvWLN4AuxPwVzzVZMYYoFeSK9ih+Ndm6v
sttfJh8pNjSKMpklcdLp9+BF8FV0Ye+EsXVb0YJ0yguX4ymyYAI0wuiBn49T8l2f0v/M/iiTtNBU
T5F6zIrwvKdR2ZJr3oCN4ntN9tWd2KIT1SCdNYRNKLsQjb/26htfAc8xRRBgFpd0ViqQaVMlErh5
Ry1u/1BxeUyyD31oIHYousgIBoLgcsHFvGK1fWTR2wIdgbaOxHV3ZBGwdKDqUVr/LYQo2xJ7rmEi
nRbMXYWQK2PLyqnlDK9JU+fIFw9WhZN212lUmKjCg+ROVvroc4bpPSLzQaG9EhmBVKup3iCs/AP9
d/TPh9FTtesT0RiDdHi7Voj96zwS89JgKa43NbltiO6b+E7o4NqsUDIVl2ojPjRXPh8QmClcohO3
Znf/Jdh7ZpOhUWIw/ZLTC/8L/5GQti87IeF7ntVhDC61p8Bkz2rbTKn6lD92BH+jDdnfloRkWVyb
9VPsUJC4yObAcDvPOvW/ZoUxS6K0JYAj5S/ntj9DmKViIidko9kj+OaHPE9LDQ3PIUBy1w/KCXVo
zwTtxl5BQM4NP7e/z3Nt/Ce+6gsgFwM5rmcU+H3qYzauJg5QX9CY1yGdAjD19nmPBV9eWaGrN5xw
vnl0oat+kBkUrE5O72tl+Td+yDEDOty/ajweKkW7YcGp+m4XL3uZRgi2pFMtXdUjVxli5PyfXp4d
xm0L7QGWg5FbD07iOvwhCVIi6DPuYg+KEljCeVVPcZFAlkT4Ujz94m0gcXlvzVF7+ATVdNt5KOJ+
It5uaN66qo59ltwY21dIRMCq7UdgQGryLQrVyjF8Z/LHiyv0X9OzhWhjlgngWSQgQ95XLeBJ7/ep
nRp+sPKjpd5muXtQLuJJAqGRD1yOZdqArpK9a0tsW3Fv7eZLDP7IlD6smFP85u0fW7PdaxnRY8Qs
QPnk/IOeH6n0ZUAtHX9DbgXhqGi26ReGB9fy/P+GjyPhFUx70kofa/B2oJY/Ru1P4b11Vangzd0o
sPKC7OdpbXz5CsG+LnZKkKBVDw/jyZcNtoLOjUkR8wky31l2Z5J4x1YJkAXeXxUI8/xAf5MHU+Kb
oHJS4A3aXchQo+Oq5xEaE3qp+Kj/ELExjkKfm2LTerxz7xnw7uKU+/vVItjbl8Njtn7T8chQqHxV
VxgxFqrlOEMXZaSMok3JXYMWi6otgmbJD67+bNgoeL9qmcczItuGlBDBnUEfKD3XgL9NFyPIY+QF
svT3HTU0NST5oj7W9hghmORbrMeVSCLY+0rLSYmX3UZvBlvrCe0BRon3uMIQ3B71abeOiJUkOddF
fxu9bWc8rKUyr1UC3QAtX1BoI2cwKy48PQ7oQPE6EDyrbdaOrr2VqvOXNGaYk5eS7s2mBb2KUhno
hZrBOTsvQj6BZqqnox2ZSyRYFpkKbIs3vOxZvQLn6NYxx3m96ujNQXXykSmJ5N052GbXjc9DBgMl
gMmAHhyT/bmzjRnEvWKHDyeCFwF8CzaKdDPHzBE2Ltv6PMJgV7T7vbPNVYaGG9Nd4U9RGD3ABrQN
vGyUcLh9w+BMmH2qr384oM+bRBwNIvHPzw012FXivmN5P30ot2HG8rYMFSfPehyz20SR5MXKiKG8
ZgDgE0uz7k39Q1J3QK1tgBA5JUsICNqJISK6ywjbHPqiqtysf734YDKL9pFy5kaxG6fhlt8OBqEy
DjpJJHMLidXdUaRSEIuc39get2F9NjpzaiBjg1UFE9TNL2shBvE89plGWxSOj18/iADZOViC2WdI
r01+lykJSuAygxvrRaZHt3moI1AUZEHnYlW/nXe2toYnDFvevsJKVCzhaWuW5PHQBq4DHRPKoxjp
MCEmGpJ6SeaNePOFS8VWpuz74ZUUFhYkwqfAVedfZBqigtMJ+tEsuBolxhTPr3HL+c+TXp7C7fLE
7fkilMMH1ZPiOcwOSfSKs7DWHOxn4y8HAdYwrNXznN3lvSLsbYk8+lTeSbwHMZhoK0Lo7oHGNrRO
t/A/G9Z0s+wtwwchRFd/N7m4OQGB+9cpj3Dr9f42BTy5RmMqbWE6GFJNkC8GZ9cOixeWYMD4oIed
FX3yTuh+UtL8B9RD9Q682VG/0hpfs0yQ/I8Hy5yy5h1CrLFrhh/4/4TUIqw9zdpEV/J39xT6J+8S
r5Gd06T8VTxtwR0e57jLf4XqhJ1rS4SI5yrz2hPAEXYNsNM0Ovc/s7JvJSfrR4/lKTJvDjFskelY
8G6Omn5uwl/esDJiQXZbgPC2CFBa3OYpIlTPC0zvBn1OzqAjHjxd2HlCyQBFHr4qHncZYiAcRcnW
rZz785xrFgiDZMVIhAOvtbCWteoRf2ev/HRYt3TPQiAycATFLz5A9Y5tDZQ31NoFej/y9p3WIrcx
DSrc4hUkNYhw55jaOcaRAvi0FPCW7T/KXF9J4Hn0XgcSXj5d6DcG7bhZRqNUYnBp1vjIwMR02gwa
icbopJlTPrtR3LggaCV2F1XT42j8vApeAyoIVhzoAPuT2N0scDNgLv4KJmrQ83z85KPgum5GVM31
iS4BrDWsgvaYzNoxGzh1uCJMBHS4HY/0Hwzar3ti386BJDSG1wtiUH4NADtyKPVksdEBIS7HIgxg
EFbi5qUoUWG6VCz9iFHXqQ/LnVzWPIzyRoWYSxXeghm1z3C/MUXfc/986aiyTTe7pvzAjEy4v4Mp
KKD6/OWUXpJR1a72vO7s9qVC0zc66BNPoLO2R/VVP2Wgf3pFxe30iD7vSQ9Tlx5vI3ubSdNmXVkw
sXBDOEfryYbJlmFRbOHhT+yMZEYJVlWZ6EskplvCbF3M0oamcq4ULAPqrNu3yAVDTh6STfp7pWT6
vK5+nYSfJ3eMUn12foQMY+J9Tek+9rpaJ57+Oaki8dRXg9vf6TJF2YCyVR5wDkejj+8BR+9XLeTO
oG3feH7QP1fMx4/+Gfc7ix7AA4eMN2cpGmhC77TuvUQoXa4pcBRi7DAZtAnexnTPra2RPW7tyBlR
3jAfXOp77eL/YrAObCKMj1FAkeFrI/qimh5y8jcYPCaaKyTztg1o6LD5a1oA4P3RySehptJVsPN5
rUb4j+Nx2K6LT0Cj8GppwS0/LVAXViyhthiDJBlfh46xGBv1M3+y1HWXtYDhc/tOe0hBuT2I7AMQ
tVElPM5/m8OfQ5uyGYPTS0tqMZloLi9isLzFCKLML83A5AAIHxpKyv884z7C4bT9Axn0gtd52RA8
VrG7IMgescIHYEaTf199N4nr7MfX3DxTk57S5jmFsSmvo1YtviEkoX4Nkf7WvMmBb3qjFk9qAKlF
tMTgXGeJaqq+7/jlvTDkw7teeDmZYoZKUOZKoEBZRXfz9AISVG4vNzDRgWOVaQS0RvZ/Dz9EqRXb
1/bdNzCNZDWKGyyFr5oULCcNA3AXmghhmp8HlQ8CvxFeqWfrx/urPyU9pka/6OMyU1IB2VzBthle
Jl2KI8a4yDv8K/UH1JRkpWRwhwp0/0Lef200wcDXP/sNMGW3Cy357n6JP60oCPz5+UOxCMSkhVCD
bS7Yraa3I+iqOlrBurdR4etc++yk4LhgGkkmW0JkkVXbMrGO36/rpBPnne8Pm+X+zM8bRUJ9Rh3K
fmg7cYHCHsZBfEgmLdB48nAmWTb8/SL/5ytWNOpIGxdh4uQDKMaBtc2lxNr9XmNYANcgMljOrENs
4IFfq7Y7ItdPP4ouQdS5fUBHwUaJDqF9Bde623XILbcJx0DL7GDM/jp+ow4Em504i6RN8vOrVyB9
+rZ+Z3DQs78Yf5PBWcpV6ogaNI9PKWiQ4wa1252eWsUpnYPhJ9R1hWZ0orUjTAmkhIlcMMbLzXPT
O3fVWTuViYwZnPHhCYrBELLyW/vXjbLp3e8n3v1nTjetT0bYAelCiGkb0FQZZilgOrogse1Y3vOH
dLK8s8OfqRJh+71b53dLc7oPGAP+xoZ1gRBxQJr5LstuPtirehJws3Lhb0T5Ngfq6UiYcTZJa1wp
JKN+7WL6GyOCoZvSXifaiQQZHEpyW28b3q25gBbSNdzlZz8zk0WEaZ7bhlljWjYD2tME0meJKMiJ
xJ7Yge49Uqt4FY2nnYANkVwGW5A7x50PX0OUUjs65pCXU2Q7KMdeYec0ranj2f33ROAJX1h39nxG
lBnT3imSI5JGnxUroze3BFkHyy4aQ8JtVKfyNJJFZyqTM14BvorwMeoLN+9MvohEg/9EVU5I6Je5
EbHuYgys0tAEvNG7dZW+LL8+OMJucOLmHcfLfqVw2cMRFFR+oMgdD9wrPKeccqywhnyEOfqpviQU
Jb0uS4s5e3kvaYJfhGtAnLe8pSsO1kojA1I++CydFPhdc0abUlvEx8cTs61Z46BZzhBgFNTjAC7Y
mFSm5SAL1caijdj+VeT+MFRV6PlvO5JdbhqtaAsoMmy6bCh8J5WEnd6Uu4iSB2Hf/Mm9iT1qy1Xh
8BTeOzcJjMc9oNddqXvNQvVhgvRaOTROvP7ECHVEWtLfg0STZ0f7zxQvxfabZAVbjq9jRuhNfgOQ
x8rcLl/FtTYTHYSEnu24eGsFk2ECNuCW0AGQcw2J4HxCWqZEbOm/NcG2ZDWrCsnj5IlWLxWnhZmu
gMDt59bXIVJLvY4r3gPY1iLkjXKqN5pVobj6053CxXf4KFFR8l5hnVQ/qck0NLblxq7elUTVZRpK
lzvySzGIDpxfIhMaDISC7ILqDopiAuvistUJ+fdCv/zrsCdEbhmQ7ybbHG4pfr7F3t8xbaoA2raH
wmDAqU49bCcoFUKA1IKaykILYljNFBDMJaZDj7rorUcQivp+g0Ooa3txrHqmgtgACCbKodIgVKRy
C32+0BrW541pVGvmHRIx4+6H7C4xaa87LdUBcVHXrSzfCAibrXBMA5KT4CInl0h6x5I8Lz/yrfWs
ZHxmRN8llJkezzkamqJfN+f8CzeKC0NnMGng2bfTOQeokQQcufDaxVznTw/xSFxUy5B0Y3Wn6paL
Wup8Y1L0fY8VjMIOCjIRXxSQDVJH1tM3RmesRBYU9Jb8h/4EA8WpgPN6IuLS8eEEzgxAvgnzC1bB
VDUqVZEORzhvoGMGAD4wRZ+vw9ZWmcN2emvjEUl2InbOOIAphIgLFTBoiYc5UlaE7JhWSa5xspYN
CyD7PT7NzM7bpW+3Po8evlolgHwxQLjM5OlX9mdTbOtahgCNYUtkpY1ULG+X5+80N7zMj/yqFtSE
JZetsavPPFOlbjlJfUjw/bOL9zBIJ+rEx1luHWDva3Wl07JjKDjISeDFkD8aaBeNsm9A7V2DCp4L
PI5LtnDn0Hd8mVF4w/xMjj6nM3/J6NACpW4wn1vthfoBFRht7hUkyyXHJtKsTQnqibe1Bf+qLNmw
13r9PtO8ofXc+Y1iTojKuLU6oGaCSHaGaot8bJCFySXHGyktq6SvnpPItTGbS2Cb2KSQFq++3NvW
7IB5hD2V3e6AZbzWuIOxnm5Lm67TLL6kZh/gjAz+kKfcEJt7QQCGd7AKSFHcBGTQ6ATCMPj8F4r4
4pamv+xW+qwyCDiLeeRrCgZFNDLUGnO2kZFhKpXFAb65YPpTJVoAFqQW0KWfsI536jnhdJVuM/Yf
5Dul7ZrJ7KO37FKxkOsiY1h2GjT/zxssNCujtNKsnWKKwtcG/VTBXG9aPPQcXZUZa4F+VRYGL0/G
WDxYsDXAn/dhHUCze1Iz68hRtkrpfgLP+BtVsCJWZK4FKh7P6xooLGLdJEnQ25Qo2cMRLNmjax5e
GcYzRr9wxN6vbkW89OZtALx5ErIs5o2izuSPYPIgg5aIMRVjUx/xcvXsfXC21t/Lz3hxRttqykb8
qjTcyB/KAJ2aZrd+x//QuTEbyy4pVOhyeT5XFlnV1s5Bk0h1CyfRrPMuIlGahwGYrH2sshsu5iij
0BfQ1zkIHocrbniHfUfBPFx8FsLcyqfnV3gv7NOtXjmEqwBdbh6/KZAazURwfrRfvunMd0Oq1o3g
PsZA5YFa4+hjXRc0yGuXcu37UFAc1lwnDaOjrZrATiEb+loecUQHO+ndE0qggu9VhGB13oVRSaD8
gzPLU8d2Qd19qZTTsI+47eqyUvbIn8j5h21JOYZV6jSu8SRMNZxyERCBYRzikzqpS0EM1XNeVhUj
VyeNVvzVg4ZDYEqFa6kyiE3BfgCAnxRoa+em5hebyZGI0w8qUM21L0qJyncO3qawqRV49AyM5OBq
lJJ8sBhiDTXPLWgxKt4okNjTU7/kXKiZbeSl1CcqWY9Lqk5QMwpMYNC9Gg+otLcUgklo7B6xDzgk
X660JLVWEGAJN+AHYPg9ATX+VXr0mqhBZSa8RZKcKIGwYxt+f44Mhi88PgpLPXj4nh5UsPJ0jiTd
tY6OuWiv9BISWFuiRGDepTktRifrjUTzJlZnvQoC4lZ8q44oJAjE0r6Xzn+i8MPKgDVtwruunDwg
HSM+zzXmcLXDrb+fHzjeGMlDw9XBOsqPXhFet9tbTIOSVz9/fttxDOwDfwPIUtAc37yXoBUt3e5a
TSlct+Bwjuuwp1ByU3GQUavsQgGX0W9mCRWytgRcG2p6Gn7e8A8X9pevCr/37p/aXyeSHOK2Dm7B
JIB6Bqo+8dVhWFSNBS8XBaZymW80d7x4gbhtH1twwOgB5QsUt3TNyK6gUbCNSM+oZBInvgUSJeYi
aCGXVU9UE/rktUevR50L4pgww7IKEpF5XsnsWZIoHZ2GcEGskA4dTsm4r7Sk9yT9NAP4THqHp43c
WDTom5okChoV1QBLpPCzMC0rTXQOUf1lOIMYkD+mWx8ujmK08KerbpcQavhzMNgZHhA7rd0aNqJb
w6DFPjSxm7A19OxX8JG/z4Mv7fa//XtwSKGYsTllkEysMjoffI0I7EAyFvaVqr4Vr3p8S3kDoNOA
XlKXpYqjMouyvK8TsvSzSSXkwSIx4GO9rNSCFLl9VvRpChPJOJJz+v3PzApaNba494iY3XwwaNdp
Nkz+gQGW/UH/H3MlNPE1zCu372XrFkboWjf9qaHhxZXX3Fbh+hptBDpaIAOyx+px/yIyqOfUuGzu
NpNq6JYf2QNPe570zauc6P9xPbMYP9cRHw2IHW2Qu+9hL3Q7IUO2RN9ErS7fH0amxprDqbOblLzb
9uPeZ6Xweu+25GLlduJbXtZlZRmiYEabg3ozzmevIMHrNwwnwvn9HopHIq4BJs9lzrSd28BgdDke
PMvBz1oLPK0N68XjwAblaBVBiZ7mdG768Pq2BHt+IMXnrWSKRjVQMQVKLYvG7GbThJryxrDevrr4
glTPYPJ6QMv/JeScJmbee9o/2NS6PRcHZgtIzpVMBfFmERtyhMpklmIPAQLC0HihafuFTDKWmzhn
es6ZbSaJKZUytTUsIjvsVbC3X0BjJBFPvqaJvktkuHE1xgAQQ0KRfVlKYWijmX2UPCgYWPzvzTrQ
QxZaMnSg1+b/rIrWjPQku3kwi2qIVx/CZYLI29Nve7QuAGWYG9UE9lIR/jXGaY3viKk/5VHR7Jld
BE8azTfXvT6EJ7LdjbhyNQiuSlN1+efcsEaQXzK5wFxbEGvvByq2wRq3BReHDTKM+/zg7Z0OOF53
s+hTcAOa4M+bqD0ii+k8lU6tbwjd8ff475+gJFIq36xVlI2zmM+C+iYsTv8XchRSJ1p7bkzGgn9V
axF1pSRws2/MGm+N3JLNaz8b1mq/0dd2wsurOnFWJaWtd4aTONBGEx9iOGxzHpoOTtXxu3mFU3j2
QgiTgWMxG/n54IdhWV5zHFhj+nyhhKmNkVBpb5VbLL5iMbqIrLAcZUg99Ir043NUDfYGBYp/bOgg
GW5qeIxEXunXGwIomxuqIICgjjDbjvIDWPYJwVg0E9vU+/z9DBbjoVMjpMAf7L48OciKwDqXNIeF
3AcApOdxTxoKwwl0lV39e43iDj4lYg5v00lQ5nI++DYJHfgGC17YEr4wR4Sjd0NMcU9HS/L9Bqo1
ycd9UdR/knuTQm7K+0p2KcW5Md1DTSVgkOa4qhyUFoMZOnSynwq7I1g9Q1S/Uc8Wud+HAhQxD1OH
Wua/jKoaS4xZ8SfZxE5v28eoRZ97IEszKQW0zbqPUiHRvOajaOPFuNMXpsx9c+SxttBwtJfvBj9l
8feZvrRj9pfem0Ivd46cutwhqzvheHG7Kj8ZgxYZNXRuuo8kV32esLTMIcM/ZU1/3lpjVkWL8+lX
8l/nfH2ur5T7ZzdsSa8HNj7oU22/lTAgp1x2nBsPktadLCyrNaY9CYtsFIAmteL/OaL53G3x0f8S
ZiU+WIXXkqBaKmRBmxbs63aAQheT90Y/fsaHiVwN0H5kGuR5lav2t8VruJ3Oa2KMNoWihfTkQqUf
SSNZqWOwodtID133jToA6GprP7MfzvLGk81JwQaHTP47YPbNFiXLvdOxRJiXyEvd5Qxy5BMCx9S1
He4309r9tJZ+ardlZJAe84HfIhkfyHip39m6NeZXLAUHo8sOtDJ0bxUf0fGNF8/ABzNtn0czIC1K
wHA+vPF4zavXwWORCVFHGiiwy/DdpZ4KQIH4Xo2jO882EglZSsgRSy1yw0dvvYb+bDfLoQfmQP3H
zGRMnT4z9PhR10ZqsKQVgO/wK9VG/snzciiAFGI8h2BHnLlawll8OeSbIexDq8x73fqOS9dxsAkX
743zRLh80QFmd28+LyZJq6BVHEDT/sidoklgH7WVQfaFYPROC1WQWgaukzs8OD+lLj6n3WvONEpq
ZwctiamhLw80/f6QVk0Je8U6jFYJESoQIKyVdtaGSTDSAoASbeVXlCVw5hQjX9hVu/1+lBwM08rr
3bFoGBizo8IXHHtGORS3oHkT2reu3Pwbpq+hraZufiM5ELiQ7TVZ6cJbviWnm97bHEkG/XK5iGsp
jtNkMLkqgsQ+j6fMK118ep7wAT47t58gamGtRgEfY3X63i3iWFX76Rffsl63tihYES0jNVHwZmK1
5s+ag6/HEOfxU4oBAilBwEwWP7Bye2UqB6b5FI9jiHbX8spyn5R/+BIgdMAdRTRw7Q9ClDIhMBry
rlUw2+PccQ6c0aokkw5C6TncJsv2J5ElN+XjdrAzMz+1+/PSnR75zYpI8N8Jp03OBI7GMTvBTa4e
dov2B1OmZDqu5rWJpGTDtHYX93KwMThU64AUPnj5Qyizkv+hlwBQ18fjpHIopPiGa5E2lYyhNBQR
ZBL470X3OZEncTwv4+mLoPbTYeKYEnznk2F0XYX430yF2d82n7y2M7mKZ4OJMN9HkO+CpsXBn4n4
pLeaMtsQd06G7RaWO9mxJSzgxG/e6CAR70i79h59uOK0iW3xdCxi+zOZ9/7sMd7qZMkqEY0qjMKL
haRgE7UHdjkEK0kAtWOyommZ2I+DCJtkJtpOj7zypPzb3xfW3FKZfSmSUzbkYBmp6RfmSNjyX1O+
t5nko2y3/3MUdLNX6sfPZ8ooQ3E1anFz5l3tyf472w3P1d3tqJXjI+cLImY8QDF78YqVyNEOBaSZ
nzTUqEESI8vg2IUfOpMuhW6rvxTzH0h+40I5Sbk64L8fC0KXIxJMfVqdQU6Xop+uxDncHUF438Mf
25z4CAoJrqRx5SifyvTszIJwxaNbJKflEpsLWddU4cR3W9WKwbqEb0w/XKPlAidmsPIC3SbvEoL4
4YojLklieDTnfQpPPR4+BGW/z1y/BE5umQSu83kBT0zpQEYVoVfL+AQVav/RB7U7+Y9XNpnJ705y
IiCROkczRqY1PHzr+n9YNmRcCdNTrkfet0EVVDcQdO51LfIzCeuJ4nRM3fZfaiiBTDatt7GNJclT
eJl6BJPyNhIJJC3YdyHhNnxgKwvY1MD9xXlDH8BVYj9QwEP4M0JtV0Z+/X1lgCxPyn88r2BRcyuh
j7kkXiu06SLd72HoM0z/MRbbmvwL9ADnMKOwuyyb4byf+3/iIeMf2GXhV3pjXKZsDyr/jviNPK0q
BaIfAkyFUCxb3rrThmRQL0PC/oLUETReujRRWXTkp1e1kIiuJ96ChRxh6hVCjn4+av1jOdr9LUOu
jbAUzYFBNwO1tACV5H9a8yhFXQWOW8PsC1m2FkW2lzxDW2Ix5PpOV96BfqwunxFcTOb+s49Y/VzV
ufgKU4hgOfJ3p9FqcFgVNIpSktMyFiaHxeXaJ6o05hk0cBhjmHOiLe2cYYlKSwjNkkQxobzf+UUR
Fv+bRzm4u9b+1q6D2XDIjwgeDV/YPLbuqJ/lnqcz/V1pBE1yjgIpsrRXm8V2QKuhxxSE54fouBMM
sz9LGfYz56u8WzXxYGt3RxEKV1yLxwtULyST0M0dIgrG+XBdffXJYv5mZGQjdMGm1WnECzMZj2Es
NcVEIOobs7gJsiSuLPxHHBZZSAeSCc6YXIbnnMaIkoHaAxjVdRjee/+ocvlrslBuE5GkjngSxGjK
gzfWXScXZQ4eIvo+nXpTb0PqrUfaG+puN2tLVe9xNIe84xkcOKtMODwcbH8AUiaEgFJI2p7Bw+YF
hxhiBlY+6tbQsZjDrl6yER/TNytnVuvUyWyYDaM/lGqEoJVYnBVe5eKsvtNEQ3EBRwo2fQo6hsus
F21MSS/NCyvUHdcyVb8uhOJoiRgOsIYcgjO2UnJnoi6lkiUejnHpq9Nq8s3uHU9ij7+7fuoVlgHK
wwIkfPiXmE65uFE7RvTA8MNBrxLmakd17vr7pzFZA4IwvsxrJOzgLRs12qlqjeJqPNyPa19/TLos
FEedJ0AfQt5EXziZ3Ph2ygku/QzxW0xpUvY8fftMkf27T1r51HwcN6oXCDBVOuiRsVrAWFD6Ydyt
D/2XOjthN2+jwCQacf/O0r8tg9+BVIJjjzJ0o27eCsJ6ygArdb9ku9fV3islJYo0E8Y4W2VTNmum
7S40dGYtc+9918k/qiiJgiXTolK0nHLQYVskWl6X4EkgZHCuVqD6VE2l0oJyUe9muPNXE9t1QPeR
Zs1cwtjYGONTKRNcmrwDYuii0HTj2okx/Sw5468wVOuB9rj5vVuGvjgpwk2SVq8x+blBG24G54p0
M7jB9QlB82wzXAvGDvaQN2s1z0z1LqoOOea/HR4ImKI3I/HS6/lyn1bjsUpGFrIm8HP4HIKZGxUJ
+ruOmcT8VJK8PJZ05wwsrgxD2mPsk34HY18psk+RAawLc/FMt0np3slp1d7TEbXhmKoxBQRlh01l
tVmOmuKBT8rJYQBVRl8CIitSYgXFQ9phjI75KNgvGd8PpB/NdS/xjP36kGNJ3ksm5ATTOADClZDO
BGSmrjiv2Hcs8Nyb3m1sT9sTciA3i5ztUWSXYIHbRFVD1bvUPhp/diECwn2YDVqmKlZpcfpAx7Qj
iell1H4t971NMPanEMlEdlDnYH7uDSDY0MQiaWO0QCfWFE1AudFL0LTOneynZpklC8pqYxnnEMty
oYoqpnB1coP130oJcBaosLN7lT714IPfuARwZn/7JtTn1Ts08sLw/bBEyOMbHX9Aw6Su3+5kuN72
YaoGE/FkaSQcjNkOgL8odoM1phIb6r+pdzJZy8TQjT9EMaxkgSYp2Qh1CeBQgTms91Z4vJcFZqES
Vkuk3zAg35pG+04FWqL1YFao36NvCegl4MZ3BX6OXZb/DoYhdIrQAbw5pr7fe+8rRsHErduMV013
pKdgvx9aIldUVQbRRyFqVLy74J0WVVSstwsPNPPC7zXeRkZpjkLRYAEEgyAHA6p9z2jsBO6jZ4Bi
8gvoNndUe+07UjzXCCNYlRJlZ2qB/lt4CLbAuynqDwsbs1xtLgZMmbeROWwE+t0R5n5CDVpTv/YK
c9CyslAy8gL4Xq4YkYJWtbUj2lU79zEtcQpdD99ZuiTktjsIBzjz1O+vVNYq7z6MeVOpZ8fdhrkf
68oMlyF0NFHKauSihT9V2DbvvLjPYCH+LfcNPxp0RptSYIPvWhFl9mc4TnAWmbmKTCM5QwhIc5yl
Jv0S4ppVAVeshYU3sF37ROi0/O3uP5toU9Ac++bMj7L4S8PoYXGSLuuYEuzL8mlxpz1eU6dTnY4R
ex167sCQHtEV9BQC0ujLoQOJiNY+cFSq94t9Uk/1aljKK9UQKMbg4KAMZTx9IbQPVp8KlM78dVbH
naYy3dRpHOFYQJMESngvlXYZcH8duP6FedfHKwFtde+FmcuPj7uyQXOswT+rLfX2XivM4arvUfFK
Jw9l/292q0fBmn6JjN/4JZmCyIB3bAp4pVa3niyd8eYVONLkHd7COPBNlhpEzei4dFggpGAmZMuP
9z+DhrOzTUDAGfr07EBuwxkD8JDKKvJBS9l12cvYmau5eBWQJKMheXEtWpva0o+3B1aKeEv6g3ab
v8Ld9N6rggfVOS+yxARr3AXpi5hTGAmqd+blXDdyCGg2/oA87xjq/NHN0CpmX1rQgJn2OR9wAU3B
0QuhulEgywW7d9H+b7wW/24ntIRjxFKZJeME3H0j/ycoDY4oNVP6A/J7hvx2KLkGekP02FDtmORs
vAs81AHFz7HOuNFl8RA8DrTZxj4LqdlkE0AcfRr6WiyfE20clnP6ShyzH2YvJKd/eCke9Am8QWU1
/E8AZs9YI9Zti9wgkMyPr03z5XrOcmvoOSmQZhv+Ies8ZjP3ipnkgzrATPBfTS5hluOn0Oc+OLfD
cOGI75IapcXSadC7RmUboHXnQIpCHlDDBUpQAUtC8vow+KexOPt4i+H1y+74crKb2x6/st/OgRCY
vFvwKTed6jYnmhd37aI7bBqlopgk448QCgrSc9ErodjTNCMCAyHoBUOiWiQu1AFcf8NfSoiappmn
/qqXcBAeOiB8cz5ygXSoX6/GuNNNv9uSt6WY3L6mgfvYgvdkvLR5KY0JVS5c2wkq+k68UB3UjFXf
7AEIER36thIe6FofeTBrCl7tYofHn5cQofIPF9or0ygYY03DowLQT4TB92oHuGcO4cN+WTeheuTx
lLPXPyv9iQZm1rY8FYUOn7ud/KkFcHmc6KaR7i7ujXeLyqRttQcBax5YZMgJjKHrjPVveFX9tDcw
48VIdTuf/ycNAt51bX4E0h1RSFuJ4IVK0CkImO2MaW/g13mgeC1wZn09Tx/ICPYWmd4QcT3pXwmj
PO311qnBKw0XS4vvsYn8eNYWO3RkAIyPvwiG+TwUQLky2VFWG2DHTxzLdqgD/LCbQgnpysk/wwDj
RxkKyebscTvW0K+lhvtnm9H4x5uITuKrjg1c4aEXsBZolzZiwBO4TntadJajZyxIRSSxuhPGphUe
D/aBNPMBs5AbS5xoJbotqxTiGqXtp1yHRiN9a+Xu2ZqVTdsbqpWfGmw1FeE3DPOoHCQ4Ym/tnbm9
ycy4m7Bk9sDYebBGOnvKV7nNkIpKfPgMex9Ur4Xf5FOFUkRnozVQ8oT17XXZd79/Do5I0M7b8il+
707afVmgv9uZZCFIGE88JYT7b1KjdIpVJRk/uaqPycY2c/ErHCxsj4+4mJZdKgUzXv7p6AZBAfNC
5/RfJ+3jnLiUJnZI0hf9Vqt6FQdglutGhKEavgtKA2Z8WdToRAlyspqImUNuhTvVEnCyhBdUqRc2
xfqllztVfhd+rQOb1N5Q3qrYSkf7+IO1sgFQ4bJiotoWTcIhJXhP5IM+1wzUzNnwSl/W0qPF23ni
yBFmxUAtAs0kNhPsiftn6YSrLNfw0Cd1mZfGpGsTgXbkob5NhlHPRvF7eXPPiEiF2Wjx87i1KtEa
ZkmW4IQoj5T7aKd3lkubBGY537FQp/Zh4YLnkiupJUrMT1zeWD1TSmO8LNRDT1k4nmLGey0kgMBY
MRCwnghUaCG+5uC4RKx86fgY0u39io+IrvP7X8pxmKNudu6aW9qX3/t7hOi9D7M++vin2xLkqYP6
MQ3hFd5Kb2OHuC0PVPGLtdqLVCAmcBKT+oka/yh53969W+upk/OOCPmtCY8HAmaAsru7cbqTjOIg
0vAsBaBjpNc/xZkIzulQoqeleYFT5MlhOZoZUtfit6HRLtB88qaIdBm5Wzrnk+Muw2MHpJu8Revq
Lj6o6MhRGek5000ZUBVLpe7UiRnYZJTQjkxJUq9yY/zRIz1XztKP+tfGGojjip6ECaWrhSqpid42
PRQATCizhP6qVg62jH35xzF4R+nbGvd1iJe5vEggklEsMUfZ4Ssp6AcIT8+jDsGI5dmx5ztTXoL6
AfalgzJLq342UXmNXMXiQgCtYQB4vwutvn8ws9x0kX0bo+71SqICvK4WptCvQBpdZUQa95YznJHq
dLQwL0oht+uLR6K45X9LesJ2Cv+dUN9gmtD7Ob4XQKMND5nuKJsZyG8ijQKZNodfGED+/gFoHdwL
QeRGHX4cFsa2zzuET4cxF/nebVqPZ7QOh8NOQr9ILaccJA0sBt+marVmaQPSpwSIIP9CcGXk58yq
qOxDdTjccFz8cXo44FjLWx6ueDUVSUzLlNewDCEjp1jiauLRhc5GD0zc3yGR+C0iWj5tLW0F4LD4
fJMHt39e5pABdEIA6SypPKkUkV/5Onx6qz1QiVWnx8eUFPAtTEVPMYktl8NYbw/+woNi8jBGap9w
PWxmJEQq11bVREBQbr4mKY3nHunCnx/dr+61Q4NZZ2rcK4+vyKyQJrvZh/rfgpGgqWcez8I0Q6wu
sdPGL2837weq2wcdxGf8FnbYZIItKMpGBAMEYVCv+xCP2GY0zfThnKUTONGQll+nLGOQ0DlWWW6d
0gNe1KiMRBLQyg28zaIqvqUpgC3QA/4LoLsDm2HrRGKqiSa6LAXBV+Al9+kijHgkpMQIwfqvCic5
n0gVN9FE/mfZ47T2wlvcb5Rn6zbe5gnv/iW2zoomzH8cS4xS+JYhe0HoKzdAgzEtdDeuFR2/kJMd
YXtJsf8Z9Nlnu/cseJveRg3IO3bbcKw5J4TVXTJGXoA2WWU8XdoivVJQdnN/HAIolkubFR6hPiLK
MtQmj21f0zxasSJEClRIcSJeo2RN26aHHc/phnZwKNu695ikMG2lx6bsHCqz9ZTbfIbYNg2JFHEg
E7VqhPhNKLkDZd9pMInksg9eikqgjMebf6ecT9b2WTwsMrQ2N5RFqH7Dj39riRhI1KryVgftq4f8
ByLjWHekTRrXjxyTOdmj9zVDbWjFENO3FvmyVX+Hq2vPcsrudtHq/RK7fpv94FsoIB0Ep/iA8M6B
+C0nHHcg+JCQOs8TXTr0nCTT+2nAfccgaYndLyMzsd9v4Hz3n9LO0zjxCjTqYVSOJZuPktSpl1+W
Ndbhzz7TbcW7to9jyDagX+yuFAGJIowzG8dcy85lLVr+Z2jMA8Bch/blPk+Rr1HFQwG20KmanyvH
8qWbpllFqhS73vSoUgRwxC7egzQKdmYV8yeUirMCMafPwAELVQtZtWX985AmOo6G611wzqkzmR2p
cjBX1v8KB01ewsuQxueinhLB4ppcDhs2o7UrrrniKhfC08vdf7Q6AdKtF/3+SUruAnCEXOBJ2GxV
S84UR0v8NwzdR8Svi1+68Zb2BV5NrFPFF0m05w5pzN8y+/l4i7HY38UPILydztP+bvtXy2xTEs58
fWkWl+9oWz29ClH2YK1bZq6SYqcn6g5LRmYVKlD5rxQ7FbrLqwevWDY0KX1O9DFUKmO2muanv8Zr
kCy+KfsO+tf5bwKyW2wpMYpChWfPrks8oy66FXdA28OZfex3qnZT1cFkgiZy1M3g7t4IoOknJsoi
OUmToLtyreGVBZkmM2RbAsbhKUe90rLRT5EBX7idfjcSiQOGxDrbwNTL+IZ7YcR2dQivWVV6NE/n
omX+3lI+nGp8MvUzBsfWyk4bzLabIoR4JoegoxSZfoc6J0aj7/G3zcySweVvyduzdFDGg6mfQb++
kYmQ1XAiAiCJ5SVxgpoppjeIxoRitjxz/dXmXUYkACOiedQu4OSzQETVkOT/fnF7Iz7mN89wwZ6u
XgzFYmiKsafw6Ojac8yQWKREmsVb21T0oNANOdPEVIyqsQD090afhcSwD4kGDonrQjkFru0G22jY
nKdJXpNL8p/hLk3fwJ4Qb/cQxNKrLKQQHm8z3E0dKCRiEsUR1ILafQEglx1/0TNv8ebCh+Pzg3dG
dI1lYuQRwLXtOM8J4Qjpvzj7i8tLEBLDMBcKKf6Xrnx4+nd8mSah2py6Uivdyn2VV0OGIwJ49H6M
O+T4YYWOVU5NK39qUp58pilmYluxUiJkPiwS/oiy3jrsli38JjPqkybQGaOGYBxavG6BRxjY18FF
NcAH3YbGDFe7Dx25/qjpfiLfl0b8QzwL38wXEn6gY604IY6KdAkEOF44ecj2Q9ZSXxcqFkUM2ttF
WCisOw8JTyrY/N/fhEBubXDxIEjAw7xqgEYeVn1qoHiMq78X8BtZu1zQYvhpw1imMUdYLuSJQzTg
EGpgGzdr6fV2Sr/XgFza1M0Qq7J+Ke02cG0+sp8lUuQ/cM5Juq+N1cNmP7MfODX4uFKGGiJ8FeRC
Hw1MuKdePpmbnZv9ysluLPlLitS8PRn/6eOjZjrknGN6OfzY8ngmNUayd+LUFAg6hKk6upkBFpKP
okXtIpiQf/n4KtqWpAqL3RcbB+BGNB0g2wdWeSS799y+2ZqTk3gPMkEYi2XcSyVjTmLIVHW3mG9L
TdI1czZkgf9IPWyKpZk5L6hFNY6KFxoRH5USpZU3TBgGnTdzI5Djx1sXGPgSw45jNMtkIwlCegXe
qs/RkBG6bBLkGCjOVgOSIkJkMYmjTv/iEkWeWEz+n3YsMc4shyZSXDTSwEGtfhgMhNMKviQlP/ef
lAV0Utgrj84s/kuRwsPxBuq3SzDQemqHAphKvxaYCugOrj+XB4GHCIZhSLN2z5SDBHyxSFdz+f3C
PgPbb55APuTZn+jmFJ3rwOVgOBgsDjs+1zhpgPLd6q/MdyXbf8bOyLHWJyxgZi2Y8VRzXyT6W+cT
i77xd+KJW0zLc95/mRHWZQEWR/V5CJcwMNtbAyAjYdnqMSJUcawH8drm9WbTWm5zjyiq7hPfEEEv
LCmKY2N/VYc8I6GA1RyQjQWAiMag9KSlKrt5pmEwj144KnT1wH/5RDX8zkwhoJMFIlaD5UBbmwUt
PX2tiIPxgGAD1TaB/SrHbcO08CtTIZPTUnLRqX3ftiN9dHT5ZphnSN6y9nMgLFMV2dSf6DWy6MW6
WNTIk5kXSv77v3PDmm/BMTGHXV2ZQ6yKhJWzMF5CgTrmuuMY1EdDTwlu2B1JjjiT1M/kCtdwgVKJ
XkiCDW9MLK6bYbQ7mCCZQjhVAYZlqbFKdpBkv9RImxw6649N50Ak3o1WOdptof6+wYIDiyCF2waX
qEjoHzv7+GtOrmSwW3xXUW3jW4mmP6eRqul/JYWPr1sgAJV84vKAEFpeQ/neaMJPAlqn0+Nwig2I
/gxUBdwgWhYNZhiFLnSmYfKLpeuAFgO8l4WgkG4V8/tT5m8unpzQi24Ezepg8gVVIRJVVQGaM/N+
OUCpaOzPUpVY3nt/Im6X6K62QmsA9izBQklXurEt70W3wqhNeUUd6WSteyeTHH5mG5sCKwZZDzFV
h1opG1uyLY98UAOAkI0hz5JH5f/BRmQikvCFRugTCPT+lj3QtGuvx7aK9CcIfrBpHeklqcAeala4
/SQDooIWFhDw43DkWGUkYSo6ZwAqtGgxrBDHcfwgr8VDfXgDdjfqD2M3V9kgEWrnaKAZXFpyvJ48
dKwd0pCsfntrCP5/ay/IN54UQU4YDyp1NK3VG87aICvfpX0Ds4HCaO/hy0yA5Ad0mqFqpPlue5/c
ej4lPbqX4hvWCeUCH5YgNfrBCYa1PkvrHhl2i58qztZo2caqoOqbXe9YiSQkoglcSYXPM3/aR2zG
PFiCrsQ+HXqFuRfrpUVn2L7/02FB66QDyt7A87VzW9ikUz2xJa7ZfegqfWKIwkLnPpSqA9yHzAfH
ImfU77T4xpFkbuVPRqV0CzjLWW+wg9wLFPNVRJnGjdNoqEOSkoLWYrl1/jOuOzA5JO60x8cyARiI
aC0MpYLSoSY/qCaofx0aoJGp9zsI5rrbxrARpAu9z006gdQ4RGwL6kT6jEEhniD68fmw8y5MRDWt
upuX1n/6wNrSKHMIlgcPqTy523JOD9hdTFxO8JwiIfVA5sUnEuBtE51tf8+C7yG7EN6sgSCk+JKk
6GA1RsayrljirjOAYYay+NuatLSLFqfyIOnEjB4uAi1MmB1NnaVAbbo7c/m6rCTOkjO4vLs7RTrs
U10exb+OYOs37KdLe1EcfIktGLXacGRy73VojU1yEf71tT212jGTTrhleGFMezmCM55iitSrBX8A
X4PQ77LLIF3imGMf3ztXwvCwCyl/yUBiUmiNDxJjqfibAZRGr4XgTfumxdzAWUWs7XsngW0qjOoy
0se1p1/7qYeERuyZrY9JycYZb1RULrT9GG5hRdRow4OzvmWf/zCloEAg6CAorDEMu28M2yZgfFBV
El64elmgLc6w+nzk4eDXstwG16KDmrBg0+QcP+xvFYMV845gO49OnyeJRBkW365jb72DKGFVhckB
kE9z6FuyFQsv8gs9ZiX37JbvNQTQyvRSZz3RLq2E3IM7s3Xm3354dKk2lqcMUqcd73G5L84FG+Tg
gJ/FBYH7keBneJbFiWqYX2TTOKZZvrYluVrgBGWS1BH2iWxQXwPvp1JzwlCNIA6/AsfxULa5uQf6
Ig67xzdDRDv+metkVw4OfnIYPNqOvZ9qIpwR4vlUzInWPxK+gDc5/Ukno2Qt1i1WX83NEygS2LRg
NTLeYavzTUIr8avIdZIfvFsPAc1GI6OuUAYGdgrKwxN0fzFw3VUPUH3Wom40aGkGPyslXohJDm5F
A/X91GfGRS/ceiiT5Us+idvgnpZ6syylEya4Hq64duDOopWTgmk7q8ykuVD/GOdR6Zu8phn1PXEH
ncSgvTfe44a9jM5ba+xWKTF7tnGgpaWMhEQD+Y8iHM8TR5Syd2PLXFZl0ZrglVos/DBNiOjEHjfx
mcdugJLzEmlf/cysAW0B6HtsNywTRDCEIdPP4enhRUUrIES7Ccp1j4CnaCmXxUE3jGNFM4RyIuiD
4FJYO/NHRwoWcZwRnN/5+QRx4dc5q3Hh7vRq+ipBELDS9aDxh7yEOuDUPP8RvNiKzihml8CQl0ux
ARDDn8v+YvnX4I6WAcJlWETBtY9b4yMljoHHh67iJebmTD1EPyMSfCa+DNWFv6JyCekaeXO9jZuo
sccs9QjAeySn0C1K4Ue62wSsGBL9WCpdn4G/EmGUcajr3Dfuu+NMslCF6FGDanCfIP68i3q/lhLy
VjNGDxJWKyqERFO3Psbp/d9rh/dVvKk3ZNaZbWcvvJJgZ4arWflyyyiMmXHFAulhQwIexKMIYYm8
SEd3kFCtc2gP8P55LUYp8ogjXcCPzV1z/cG1vF2//9XaVIMvW6UwBFOzZacDogM9I16y5CprDZaK
ulgua/18hZ2p1nUXn61L8l0QsleJDDhlSRf9Lzb7inuDJgUuoC/04DhudL9gShs4fO6ExgaUOR25
XzCmp2kwwLrQVR6lr1dLj3H/cogYXKX2VbDOuRV0voh6LgKihnlSwHJCzFSXsGWtX9pWQ/TPhvI6
PsyEQ0ZtpTvWxywQhOoMlCO5GheWZFZIgXx0D1MlZYWtXqq50tt6Ojg4lohTayRFYIrg0Y9c2Cuo
sgsPJhDOJuRV3yKxUHkb+f/7UrrI/mpfSO6MfOVIIDBp1WsVrX94sThlCyN2vHcIc1DsWpaxRVms
4WL5lti3LRXzFZJ1ZaHCLZM4GtA0Fc/ryYB33mfaLHTAPVt+Z19Xr82qKCHsaFMRom+hCSFg/DS4
ZgJoRvFwJ4dvGT8uH538MgqFByAmRGbB9uaJuM1itZGr/sCl8YcyVYIyW7V0V6ZZOHyxwqkHrmvd
jfnGswnxaIAM3cSukSzv6aCQtEsLEza3SzGh04oh47IF9gQnwkHOWSGNlr6FLFRck2UNK7kCiY1G
n/HkuzJCNwnEV4vrFj6vxXMoQDeTdCzDUpPwnLvg6lTioFerJz4dqo3EIgfc6T2BviQSVz1bbDh0
PuUjXmJktYfJ5AYKlyDGnmN33N/L2vUmJI71JSr8dQ4oZBqJDb4MoUY/r5Pw38IdUJofasnXF0YM
Qq+MDLru2HA2AXJIG1pBNZtEGBZlqhShpwWL0FFDEGlK+cN71rik2kmJtkdZrHWRbJ1KCsYhmAWB
xwHtaL4cHsQHBD3jNG32Kw9yl0n9URRiL9DUxWh8OkRm04xU9miBbThq5YzHZ0b8/mxICVfNbXwW
uOuZiWK2caiz/A20SdB77rndYQ7J9BN44J14qOMdFriWLLtIbFVWMY26HjORQt4+Aw+FfGjKIg7p
ZYKqi8Xb8DikiUU9gGfG6n/iiGakVnOCb43YpmCfZRER7XblkLCGLOO/2Pxtg7rhewTKs4bY/2QX
P7FQpxIlVINVmKzivy5rOv3DSQLKLlt20ZmAEAYpY+mR09vEThtnJT6ZuCpPW77jVV2IBXg5O6b+
eBZzTTgbjxQigy6WTC2kwR6H4oNL2OKo+hv2Z1YX+8J8xSxFROCzCwjl2aYe5odKA/qfeq29BIvR
WojrG+pSRpoc2Bmt9VVP0Pceks8d9sx9sjzWwWBOawSLqbvW2tMqj1JB0RgfoG1zDZ9S5WoTtfN6
8Go54RET7dGQo+9XjML73/zZRjfQzDXcnn7L9ZEjZ4FJdYReKlqok/PHbeXKj3UHsJwuQLnrntDU
r3Qlj43vxJ1RHX1K7cTMBf1Xh7mvsRjqsdXNekC/kzKsKlufnbLTNNOQNIVU/N/yAgEiZFGGFbtA
Z+3L94fWdTNNVVKtB7cBBrTS9kc4RFRLnwqmd9Zf2uRhtakuR2P8tOdbXbH9DnebzyC4xxmU6vtp
AFamwMfFcIVCe74eIoNsq2IwhYLzfIAyt3/h0JRaUOTkcU67CDXgsK0MuoxbirXRBido33Syt4ZH
WgVcnyxcMSiYZZ8oZFhUdX90Aaj7USiWpm7pc9Ck/dFRojSu5puTDg6ILoOQSI2fVmzp3kFlyO3O
XyAw0nt2d/ADhopONJsNtclTxo6bozn/8liDLjAAhmpNpTHilEmDXwll8zT1Uv1BBRelLlZUnQm6
mLU3IJiJQZK9J2skChWO+4ltGsnaeve50CE3Ogf4s8LaM0tcyKdBTXOMKcwzPv9W8Ux6TndHID2L
sJoPVkrrEU/xrp6v2akpeQk1Bh45t2tGdqUdMJpuJQ+6xIJMVz0vC/iOQiB8poxk7L29gcE20Ors
cPGktALHJaOtxOorU54fwJaReo5ngnj/PXTI2tdmci4jbfmTRtegNXfBi3Yqx5ZSIMQqvhR8Wu5W
/czkblF2/8rHX+DOKH4PPkH0U8S+lVTEaxNjn3V/GpPd70hOq7VtJN27hQLRoua9j0NsSY+pumZ3
s+dbiUvuMW2xzXM452xnbYVR7NZy5gn1G8lQ6hnXtoV7DUOQ+NbfPgq4p6RKpN8UHiRM1F6gvPD7
EBSitdOebb620pnw9mJGBtSapnunVC5oMbMenIzvl/NLjJeSm1y5Fgf7VPSZdS9U/qjQSrQayQiP
IKUwxZgV0l/jWYVWgyzAOP+dx0P+qPywISUX4OYlZOSysZCK1+RjcnTMUL9ZN71Vg6h7cJGGraLt
QQnTrW5baDKNTGX/pGyVpkmAPgfswixTBn6L7xj+/rw1amrWz1jxq/ar3U4B44wEYvNIJFkislna
bc3pkXqGRBG3FpoIDh7CyujKKpSrEuoW90kLZJuR8I+eR4K4fhWmahsoD1MVE5pLZxohaAHlkKtH
oaE0MhLpJ+pSdsh3VoDi8/opD33RhPNP4yjqNXq2h/O17PAGpo3Mr0YKDEwZ3tIfrp2H4kmyu86n
Mevbre5kzywtkVy/73S/DusC9FxfbyRyVdrgPZkPz8qWR5JQ4xyBR+eYnrQiONDf8DDSXhRIRCIR
Iwj/+ywYylr9m5w9gJUaoL8JcqfolumLumJnmVHwJhEKJ6dnF/zIgPrStUHX3vaSaprjoCtzudTD
iIXvJQfG4764Fru86Z/ywAJ+0XFTDMwfKEs+KFb3sQLhZJHUNFukig1AZDGL5WQal+eC6o/Iofax
etEFOyQOnxiPGY7cVLI5xINSqPlHcJa3Li0VVuwP3aMOf8PpCF/2uWOaPkUxENbrIZQZInfczTZW
Y5sVy9vG4pXyW0BDo1Gj67+BapH3PnoxUBL+VCV0AgRRj8A7De1KQwDU3CYXUDTuc+VjLA5VrVS/
Z4LzhMi7E2WrbIIHJfTLFsFWzADbEeBFkSEmWmdgzBejFkb+VREPj5KVks9LtbaiLThYuVFzNRhS
DpiQWKZlZbGIUPy2WwdJs1TdpUb7aO2AsWmr2WL6aK30vfS3itXe8pZIbJd43z/TZtqTBL+6Epbg
hAaXbQO4fnYbGdTovIes9E1ggXlQNckZAX/+piXnIXKUiOhMoVNCrbFDNA3vGv6XXAqY79c4fi0U
4pDtlkwpHJbctemqOBRhp/1G1SdvuVTxRD3eqp4QVM9Pz/FtRnwIH6Bca9/unRtppdw8ZjbIF+nx
VjN1GiCoLaaXIjqeeZzofeyj02sKJAeGRCLNUrGuCYp0FDNfdD+eXhOyH/pwquagzvsqcW9ZD/33
tDcigc32Q3sMg5IHX2u6LuqbYMdhj7BleSg2vTBipUZP3mL5BUh5dS9HCJBQpnLAysf4oHX5b4Wp
CN5iB1u4i5RWXqHNOkL0ulyyoT2RDyrVTioT94oS1TWO3ilEiPU55KKyRe/Q/wOXepBf11phxW96
4K+L1bZHk7E21bVFKZieC6LiEMXje7gtFPeiMnA8y/onjQ+W6iQOq+ovd6/seWjb+lGIE+1cu7di
6p3R+NnxbQzOV/HP8ebVE5AOFRclyeQua8D4uk/EaSHwtKvakXus3NXQZWMecxfbcKU+LsqGtWVc
0PuEjkNLjTGGSyqc5dzZY0gqwJMkh3ylaCyrtGPxIBIA6TvFyzom89bCvZ/Glnwfy7k/TRcZZCI6
W/JlyrEl/Z77Mh8HAG5Fo2PL2dfPQMjsjomSLdV8+BVPY2ucwAm0SK4V4YLDwzUoCLMDIsfox9n+
zbgMzlcpyQhh+Cmpf58bf5zd4Kndfhwk/jmhnYfe4q2okKsURF8IoW6ijTJyjGR3rsgriPEqHDGD
rKXc649IfB14VXtlqpCS88y9e54v5gG8C0vnv+21I+s3G9zcniwEYM7lVY/3QGW6KlBjQd9Nce/i
0qVWkS+P2QE2NDu1ClGrIkst/uWRYEjtqnG7AA1SBsatncIHS+z8sl0lGNPXXzdhaK+LPG+F8nnw
PBEEOiTiGlmgib4FRjuZQGGzw3U4Rm9ekiRlXDwrk4HsnmSY2B7g8j/xK7NxEzb6/aOyliw28y/9
NE7HnIYPTvLuqPeFQpcGAajU6Vqxd7F7DzrOyOPYwYVRndlbAT5jrNp5bX531NeKeDpQktcioSf4
QaWIAc90HdMKYti8l0zDONC+v7SwE6NiI1X+JzovYMedDQsoA9TqDICK0XqCUbZHW3XzRa3COvc7
gaRdas7g3ktlGgFPvGAGLNad69YrwjZHk/jaWKOEOQ4xQTO6Ae+jjH3ANEuCiyywbQsZMlx4ZCre
ZSk2nn60g6sGYMt1KfI2gd1meFMqj0cyYsEZUpdfm1ykn6gLFFbT5e/8W992RqoMw4JR94wmfBID
Wxd2tJsu8GWN0pQJ2rI75tirp0eMQPnhkiBswDOLjDrbMtUXvCJ6Xeu9QzltWbHCbFpVh2UgZz8J
vXXxzpRma1rDn1fUglfzlT6tA+Q37KIing/wml/pxWTd642pBPXPLBt7rz0aL7TErRoIYtTfMub9
ONtAMOMwnjQ57bo/M8jWSRlrCWGfxv2GzSWPEJn+/ttLHzvGMa7meqkXmeFG3SgnBWvRJNzCRRpZ
AsHzULdN27MOB5HkRWWT+QBgf+ftvbp+9OSFxwUTzYTvqS+DfoR2I9XpHXl2IYTt6OckK5gxwF03
Ks+uQ9Vd4vD8E3h87/YsIryupoHyInm0TfkVN2i7850MzzIPfn6xCgYfUJIycJOv2xIWbFxF0kxP
CFudJOkRmV+aSpK2IdpnzkRwWBcWHq2kZS/ySSCzD7xAmMwRiyYEeGJLoANuTAZxI8qU0bGYBFwv
ByBiGMw+FSckvguGUOUBp5QzNk2+7OIR/vNRojguzW/0TZpCNmx2gkOREneUXyoAXdQfcs2wlyoU
gxaJ9NhbKb5+4wrTHGeSc2w1Q8zphMTkre6djKxUiBV16dm4YnDtFw6N4A/D/xgWip81IVcJxANe
76gxN4wcy+GOLehn8BsclwghOZhW2KDmboX4Tu6ogtjz7ZpYi9mBQimnkNmhNch36LZbbvY6mcZ+
F4eljnaDfaX39uMRjMVC+hvwJ0Pm39twIeGfqvCWaTbpv91G6ztnxLUpHdQE5G66iuOt4aRusnPp
5g60RHk3KN8wtSHy+RxTmYR3sis3qHsdd9ti4r0xt9S43wTOYTGA747zlOZoZ6+pcLdrKmcid/e+
JN4xd+0WUgIvTiqUL+YdMqibNTLifEW1an+D5Ai5BwSQ4lf72mg+fYlWvxNg46xE1QUtEr1ItDcf
UmKJ9rcdYaArBo6niCjkR+MfhpEiSYzgfDgwj2CgmmKZYKaSmmIZMR5fRyXlSM7EISBEljb1j5kM
fLVF51dFjNbkIgPj27nrIWMlBFfJwWHFPykDxXwcI+SVLYRSQ5vT4+x2aEpQeyRpcIrwe6J29+hY
bQ8L07tEH06IoYyt752vyewch1Qw2j4iqANNLPlcYiEgj1rbxUot0AB4NdpPwBz157jZJYObesuL
yUuUKG5COMacDck1Etx30ngzLhpb0tVqc1cYzhOK13zJQBXhDyYf9o1RHhJCwqdP8p0o5w3vCfYD
HvJd3nOdbUaHCrFWPnLBYiWARIj5zoLEylpe/AAi3UCqmR3Ghxv86zQOJgtDnmZJ2sqxjebTH3i3
EHbivlVV2yneu70ujPq+CV0z8iRWMAhZxYwcqNqeSNG6wRwq+jeORZYZC0rAl0XUUZ2EZhNycWHT
OgsO4cn/lKBmAjWGxdz8rzcQejVpYiyD8rnFa0LyPhHRutUqKsZ6POqmL1LdAobVupgQCxtAeYc7
y1+6yJsF1Q8Bl7PaQ4iQmV3fQRrx17WWYtS2jMHoE11RREy+9Ek/gKrxpFO3z2ZzXaq9d0GyUaK8
KpBCJkcWIu3peo3lIurBYdEWy8SyqMm2CyspGoa33NcWcSWNtfg0sbUy3uHUctluGzaAElsaiFzm
tlfK2f7QLqb7+Ua04cev0Am09G/VW+/KUbqSJCsLhPObABInyIAnEvYH5Xr63MkKqsn0UXZRbh4/
gspkwtsn7Faucz1i63ABVC7ypfV2xRtX4/WZ3LGAY9inykIBT29zAsFDlp6T2OTZkJBgODn0j2d9
11LsjiPLIicUHuK0oBXCigt4FKyWWvJ72HBIa28/uDSULljO7tW2gVLDu8f3/7UgkLXWEu8X9hr6
NlLXYNbp1iOPCNpGu9X76lXqFXWNCVBSKss3mh+txqI6bjWuVWDnK07LL1QzD/xvgwjhFvX5jz2D
F8wj8ayX9Ne2qsCuFLwWBAX7DU0Mv/J7bnqvkXQyyI/i9Gx9XWuot6tKJC4JcY8O8PhTeYDG2O+E
6RqIor0KAeZSm1756buttfpQB2vGgdx62/5kRQcA8juXKUL+l/VzibRKhOCkpR2T/4p53Uy/KH9n
sLhXL65mys3ExNHh2h4N+fhHlJg6FFrhW+HtSbN3jWcrFwDD6jKTzxRtwxIzdSzTAO+MgPiNWklY
R+LM25gTrbTo8Zue2fcNnzJKYLKsf6GIeJGjgM95wva2amXHXalk0OzIZBxbuFahPHNUzejlXhJQ
8imqLnLk3sLkmIUGfQRXUxejpqBx739XQa1vjR3eoeUk7ypfq8uI7gGEa0Nmw4B+dz9DSj1StTz8
olfbaex1Ry2dWOPm6ZQqQFT/tOpMCLKaHeOV4rtdm/7XfHmcJ1MjaUs2+onOvowIK/LCfF2RziBN
GEWNB9TYGSgslKOBiTfzAjlwqa/TyTALFzUORKCMbxmGAGL9d8gpnJ23nNtvzHybWSEXzBI1hUaa
pDdUGtYnOjN+vlErZa74ersBrTJUtzBRxKBJvdWGNs2Zo4IRXnEsknhCDSV35+4w74yNM8oNvF79
wJWq1wiNsWLji1vS6obBrE6jyigSkqS9FtILIBg5H8P36bRnRfaGyFrsnfYhAiJy/GxzxcuZOTak
ytUt/uX+CPiYOTWSfAGDYDUvrlZxTchL7s0whCo0ErYHbd6N1idbv7cKkZU7dD0o/I9o9UH+u6S8
5FCJQC0nQWkFDpt8zI+TMT1koqJ89P7GPsyRuMmSXh6l+31yCQYPirWpuTV7hQu3JthIkwD+YI/Z
B6M+9AucTMPqh6Zh0flru3hij820EiVBC0+iuTz5M2mW3kD7uhHDvHkaGoh6cpt4XNlHhjjxAwLj
tkOLihcs3hSRuKJg7v/aEn0rQiZDRFqUmMT76Gz08dbgRo+5qbn4/rgjHYwdzfMNbRKpGVI/XLOe
EAtg1etHlcYmK7D548CRrXcpE015O/dh7zSiV2cLQN67abFY/dk11OwYosUheLDYGW3tcaVyF9ER
V2H2nKJL6gac2N++qaVBxe8/RuZbohgMILNN6tguN21U6XykSuuS1dCAwP8SEuYRkDv5Vya6T8FV
2lAReUH6V54utTcDHOHC6wA0nW2KRf6ZAzfLgMK0sthDaXj4Bwqi9xox4S93IjOpCMTh4kECF9Yl
uYHJW7KkXEsufm6cjJmTzhGve9kobQkyTmjPPkyya8lh0NgzvbDOqJAR9e+VujFb06hewZdJ/K4a
ez9c2kQztJ6kC9XvbbcFWMpI13hjbmRhU6nGXUu3gsUz0WGcKWpO46l9LwGGeEgiUcyDMRE0tWRR
Mv/Nq0bU42g9u9PsDeayhU//1mxTXQfV2u9hIi/4TO084wF++uFHtrICHiszSdWhrW/1AVNoE/g5
EPOkVEMfS4tYIwEynuYV8nrZFwQGa8hAgX5l7I/smg68ZuzGSpD3rm47T4kQY30wuhgpqM0vzGO1
bzQ31ukP0kTJkPVLzfFn1246WlBA9kaRplawP+fHLv+r7gI7oJWzvCamRnGdgzcD1EozBLHJp+10
1f/o2RQqDHBrEKirWg6ufuF/PGCmn4J9L+wWdUPNKsetGFN+7o3HGWIea5bg2FITUXCRg9Y7aX/C
ruLDbKRcan3uaqqPE3ja6JGKgOcflH3fshL3YdhRd+9n0c3UxQlf1Hjiepgacuq/iMpKah0etZTB
qAS31ckauayB4NUTGD4mNiGpLil9GQsg8EpaSiB6yU0xAuuERHE1sJElL2gKLHSvKGslZtDyMYlT
Fs4ZLI7+iKAMxXvmrl2w6ZEzTdhxkMWUtAGRLZbzNOltWzU+iFV3WJ/lK0d+OoDVnydSUBreAJSQ
+4aacwsjJNa6kEJUwhlJrEBBKLyidjBjlS8/r4P+dJbOA5FFaZvH/2FEZIjSWPFFiQPyMRaFxfio
qKX7eHNOmzCyBjxHgGeD9PSLez49xD5PtAH2nhr7vl6VcltVy+0NK5AUQ2pKNcSJ9c7LE5L5Vr8o
dqpyaMl1M9nkjcYCEVhYzVbDakiRe25osHYa2uzHYTB++ly0NVF5idm6rDe1fmO2MwR/LyLLlzcf
+5AtDCpxllXPcdHJTNds22/cTZrL0SX2lOLKf1E4+YWlLXvE2QRcFlwspRtV4dfsCNTV1N9fXMDt
gNkb+OO+YvNeacMsOJLo8tmyNrflLEz4S8jrZ/6QdVt/ZHrF14UzRv2L0FgJPLyKpAvl7sedtA3X
OUAfWgl0y32+SSaP4CURSHxXcuASzanBBcsC/ADEUCzNlP4EFBIhoEnT7lb9eDbCwenR2wqhZ1Ec
IP1qfhmpBXDGWJbFGCK3r99NJks/nutoWWvZRDrK/LIZokIsIPfoTVAkMxh6Q2S61S7FHPiKUL3h
JLF+m+GNuU7EJiVo5T974NDgrY1d5XMILJWfPZHSEhXd+uXXNDOKUOkOPcr7iLRHKnxJFALAvIW4
tvxjb+riKMRRcskffPReDQKpFBqZJqFoxi7J+XyjCMrpBAYJAK6WMSbcc820Bd7nYIreWZEnywl2
qN1fkNC1eIBnz46yMWGsDiaGiEwWijHgyX2WzFEvDtnVYloHxorEO4ffgUkF2B1I7V5mzhWUuNFp
aeaDnVD11l2AttMAqGgj2Zo8Hp8WUngmLEOvWjpWVRi8hRUf/Me3Ns2IFzsgB418V7W1LhjPOZYg
/BtqH66JOisqTTs8mxGg50gVqSV9NE/6GKDp6sNXRrd0e8xWA/QE2TCxTjSH9RFBLiOd5S+pbMhW
uQ+n57ne7gElxofh2skT7XaxKLYOQUmxMHAIO9TzyY4duxYLFr4/9MOa8B3y81dg/9vA6GXM93uZ
hRcOJYUGDKcKhTtyrl8GIrbJts2QU1jvbdTCWzvLko1jUyQkZtuBsYvywr93eJsKHgID5p1YsDso
VUGrE8zhWiPm5ZrQcjqjlcaMYxDXNPyFrpDXzIQpxj9EWvAmtNHWNugGTc/IpzHcM45i39Og0jSp
j5GkMTQi7Cjwy88HRPWET2Adm7+Yx7uGKIbjlUbmPtfS6oR9th5lCJ62EKY54Ovyc5++6JywWafh
RqSTQZyxqIB2UwsN96Lj6FzV/c3qPOffjvS6em8rXqf29O01DorMEpNeG5EqV9CeALN1CSotErZY
4e/W+1Urpk3LwpSglf+xs1o4PXZG0uD6ayBLlZW4c+YiJkIkQug120cwVHYd+aoClRLpiwN9VXtF
RFyCPdSO4FhQ4+SXmGGJ/+w3mlpj0QVyNyv0eVbeHhWBlaSqkWv4ICBbxImta+truVtG7EAsazuN
/Y732zlWSGPhIvdtsgUG6VEClHJ28Qfoe42CD6/tGeh6QkbkCk+jp1sH5yCom3Reauhn7oSIVRK/
cBvVrpr4VbaL8x2lxPjgUIgZC5pHheI7zUuFOgpnSUPoJSrtwjVNxeeVMesKQKtdcEgqXCCmloog
1JQlzE0WEyfgv6+Duh0yFth0kPkGQV1qOpCy7MELzQugO/DymLevIZaJgY5KIaf0At8a8Teubxxf
FEc0pL6cIJweW69N7WCtqe7Dw+ikpeLW7RnrMvT/Q9+SIoMCoDJtxr+zquVnmNe+5oGElim680QV
6PWYipBg/gcqPKeMSJeGypwWkVDMgm6pzH+mIh1dlqStmCuTraMXv3KYXW2DmPZdI2TsPDGDN7Nm
CVcnS+pZEeyGeil5yS3MwlPoXRxwiZrwvP/ybnN9LfdOyWC4VTKJkGhrHolW4iSFWUy0vEQt0rYO
BMm3FFu8j9yUzmQIqhndtiMCsVRVs81mHFdK/lSayZFbN92ODYlUb66BF+JJazRhnI6a8UKnQENK
U7XquxKL/LH8pWumh63PdCTK4bN9rwh0x5Nqj0UD6rNvIpyvImxyU9Sqqg/UpNClEUbdCaTTUjzO
pnIxFqcGqRqYvVcgMkGLJQL5vyD25L+i/B07LpUz1K/cR+pGRm0WIscGed0GcfVCL8kn8mKrB4GK
fnIS5aFg5ILHnBDUVOkrT5Z/Fq5aBUzUJzc8tgfbfWH6eEHByPmfoTDnuLxGlaJ8JCeM3SMzOxpf
loB5fY4rmsj9TTkuMAcqhaH1DisdmSvo1tQgCx2o6K3ekB3PsnMKPfBYZiEO0qiM1/KaeUDvETC7
BNiCOoqgAjGRb0XTIlsEPEw5GwIahqdF1iDvVdFBxObemlTWblNF5C7GIE/IZTFTlJMyh5DgTGG/
XPsPYeU51gZrjsi8zZhf7qURsoq/GqU3ZWVI5oHbipTl+9YbIwyTHWJGnWSu3ROZb4LM4Vwp/9NK
K4/hTNuP/AMvyc0dBpVHDKZWGAhQgae26mHOfAgwBJAWdcxnizz5YXCrracNjaU3nVRhBr1HTnqy
7jy5ZNC1j05B2+Do42/pd+tqIUHrZ7pCVimH6bctLBXYGocjvjijDuNyGAKHi+ZJvgwIQZpr+u12
B1qsRvKdrleIlx6Gcv/hI1+l6r9qoi/v5R9ScrXIxzQWS4vfX/EpW7hpvqZv4uqd+zFQGL2nIC+r
uIDenYY0R1hCV47MZecRKxTY/9TRsyi3kzByHvKUKtFwGJfBPQtx/zcaqYCAIAKf8ufhoKm4OtXo
oiSI6T9Ligxt/u8Hhaxt1dJ7vUt/sdOwOBkWEvMbxUKJkwApV5neDQ/VvH5jnXeXkDsNEQ48O+7W
dv2k6yEfIRJm06XOsdk9z82yqTRLAvY9t9WOariRTFtDsbuarrG6ei+UTcN0FkWsue9kkb7s9Mwr
l+crUf49UwuT+sbj4CL0VM+alUmW3dpgYLt59NWg/L6nkJWlPYmIiwqDILRcdHEKXSkLccck1o7c
uLnuJ7elmb/4Ccl93XN/RNn8ITGzxMwLztK8hmXGpSpCWpx+/i1qPqo8Nj39oQrdirjJB1WfZUBD
0532IszvWnOKR7F49a+2aOtkR2FuvQ6Webbf8Bpk02peNKdGk7vXGmcXv+m8oCY21vj7VGlyJ75b
sZwdTSu6UY0+Fvz9FtvVKZKW0FyCx+EDOBzbTIMLIxd5gmnu2+IdbDt4zU3swAw/FxKFpJ24Mi+T
mjFB0RRbQ5eldVr3d0otY3OhAP6unDkjNXQBx9dUg0zRpFWsuMFjMdNrps5PCzrFKlQUlkI3eWdl
dkrnPWGlJ46TsFLGDQXZyUXKFbZp6ZZGcRKeAvjaj+S6qkQC38tIATIrdn0Wtewaz5Akmwq5Go0l
PjmAVaoC5gPZK4VCWt4JFO/lQ9VO4gd4XJfja1uHmN85QuIS2E2u9JimSL92c/MZUpuNUvqeqkr4
F4SJtrSJg9oX2wtYTV1zFVpV2w5oUogzNzsyfUCe8AXzn3PX5C6zYrsaROk8HvuzZkcPiP0SESPQ
/uBIBgXdC6LeIIC+xXp+lrdOm8qod2dSYmAKDgn2ZV34gKpud62wNXmrVH3Niypr91sdDtaZB1z+
YYS+R92I2MZLKNE+QGpFyJWOgmhBruNMV7S3D08CvFW2TOyiMAysuRkeciBs7dFnkZ+RB7OoPV+0
NWcfvMAeToZlJOQfKgMF9aZUUU/FBA6KX30uVSVSlROnsofweNWoxPjbnA5dXYSkkQamlDyY8+Fn
tEK4yfI2VsjQZC9XoDZFAyc7k134+agsjeFDMnL+EJWMnJ5EGCds661kGO12Gu/B8GA8Vn9/ziZZ
veKQfUOYje+ZNYym1i5N/HLI10XszDs9Rwbh4TABffLhlIR76mSavqwlJLkWCTkj7p7SrBqlSFKH
uqMvCdCUikHCqtOwopyXFUFJPJBogQmB4qx5+t7TLe/Vb6WTfCFnYzKkcAKOC2jY6CYZH/eoQaCx
kAcCyvaW+dWAVhmYlxgEPazejn8L/3u9HbGAfivuE0ki1HpQg5R9fjNGtmhd7I1oEx0ccpmcmlVs
Uu7vSaRXZDao0VGKZ79A95CT2LV/9OW6xauW1GJTjEOJfjRgy0BrKqpU4TjLPB7e+dYaaGnZKIB9
b3tGzKkb9yv1IlaJuOY72XtERodQMGu88YcYeaWwD+fnbkNmruhCzj+rngP4Ey3a6IzlUz4EncRw
BsZ9SPDo3LZ1M/rBnqhmU3u82TNRxRiOOEyI1R0Z2rZrP2pnFJ36EzebF8AJBupl85tXDF/p9wRG
hYuMH/tx1GNPpPDrNf8qTUZp8XysU2wajwKVqCXP4hiqBHZRnxKhS7rnpyXB28vNCv5TrteaK07a
rE1HdjkWoVJGwgyOiEenWwQH1E/xRw9jgGYfa2m17wJ2FRHeracuTIx+D5x7k8xQ7gAsHnEXQnKi
8ZN7MPgVnQmIS5a2PFd6VjkwWdFizqrplDAbcQ1vOzb3pqED5hKtXssKZoktN2IuMfwQvn/n2R5s
48DcHKTepRmORuCf1lhvAVwp7h4MkUACjYAoTjjoBNvXoVbabM63rhR4c4wNVk/9aU3Z4LXsJexp
3gcGsj1NwD4ZM5v8CHoFOL4NcwAWftIg2e/qmEfOhpWNY2YGTULDMhB3WMqLA8A2eoxcu0zqtRuO
2/xJVCMj9/V38iwnGdJYXR3PIDUF4/U189impJuVON0mNtEwuz6d+LlxsrEiL5blt5smiQ56cwVk
85YjQcckLd1Yuf8yNCe+khUF/SSZvqQ1y0ZU9Hh6heAz0nKhBuWg1E4xjVUD8FTEumZwHzIokWVU
IqecfrKvRPQA/IyCW0IKRIkFOjFfTVQaTFFGyOB7jW+dAnLwuirw958tyMe+j/y1OTctRRW29a8w
jVm11Sugto5J2ztq2r/5E8lEC9b97rctqH5lJmuDQE2gRA/B0ntcUbngSVenNqW1waf10u1lhDBz
a9+v47F1X53wHgwPeMl3gZSxQt1guy9MWrmS+Alvk2MCW48Au7be0NhM2+jMPCE/Hn1u4SALpzjw
/JmxlwoWGmdStMiI8pdh3H+dr7b/QUchKGOAXfghne3CDhb5u0/kaZIgxpQPWtZdj6fVaZkrtef8
c/oS8IGzGGSuzrYVBsw+//15bb6/LDs0elnHCCaDQIBJibxMFpxL/94ghT6JZ0VMuOzSdGn5fQ2q
Tnv+gkTMqQ3U8qKfgsnVaSJSaQJ6IDYbSt1MKSt+7iCoRVfNot3Ft147SJFqzLJnEfW4VZEY/eHx
YEyGC9nOxh/sWhpoa81dP2htSB1uceYMwx2Na+GydTaEiOEbLrcG++uxE1rdH7H1gY8IczdyqOke
vqNEJfGRnpBlu5wfWjn88q/cQDYyE/iaPoa1u2GwvFvFpqLj4pW22N6S5HpZWEeFwZSRyjIFFaM+
Vw2RGXjjOIOGMa8cDoBUz2NId5XMQ80IjO6gmRbLJO6yujVPqnWQXxLKCtvynS7s2sc148wEpU99
K7AKyAWLF0JCzYE4vr0yJ1GH+5V8v454m0kYcw/2yk2c0HvjWBOelIxZws5r5c3DpFYagNnwRQws
w5FVedUn77wQltQrN3tbABwl9mLcjIAXRXMJ87VOulfD24mLyBMfhKz999447kcsahKa4RxCvnfI
R6qR+5w5NMWl6EtHrTDdCyN/xwGiSOLaeCxYFr+WT4Adn+fIXm7YrXtZsrsIdPEV2/FNoqju9Aqa
oGomB1jwrrg9IW6LYYG5249bHYERHFK2jJkQYx2D5UWtSSnGU89FkLflwDZUN63Bb1apn52PA7d9
SsYOeY1gtV+N924hiq+EQj+57LpofDBmLYGwCG5wVWuHhT6YHh3jUb1QqZoebtGDEUFkbDbgusTQ
3nEdOIauatAyFbgcS3fImy1r/gVHfYPr7Eiq3G8NzLIpfMCUAIrFAfwX+vann+AyChOJARLUWHAl
ib7EX1584W4e5w7Y6R4H3oHYao3UGZEPwjYHEhoNuZ4k2NBO+Y8EEJ6K9WRHXgzkEU0AWPyE3pvh
lCGc09OxdCZuDnyP4KCVqhTb4jaR8jjS/bK0z0kmf4+fjLwNAyBRhPT4c6mO6xZ+h5dr8tA2xSLO
uiBcHh53OxV0I2LvQF8eTQIwgvjRA5jI2T5RcBD6n5IaFyDVFBJO7Jj9xFKBhc6qwMDo7Q4cKbed
PfwEfoTwt8310NASvb2smQgDpnNvpsR3Be2HCc/uhKdIXdIesBLBuLT0nW7j6/KC8z79Kl9PJqk9
Cmo6bCJx3g2czXfgkS9zlmS2rThrYG+UADm8xFijC4AHYGAz51r5rFCtu49b9Se8sI+Legg8LaVg
R7yxoa1/gGHN7CyLmCGwalhJzT8X2VSwvgXHpQcoVkr4cJBp7WeHoVqbqZzmqC2pL1HYfd5RvFDn
GiZu802gdoMMW6dYFS3l8lt3xyl4Tgj9Y3Rh7NeVfWZZcTrsNB1bsZbGVZYd91Jd+23GPdZUO4ih
0UagMrY2V9XtoHB9Lb7Bf26HXv/DKeaJhuKNDvk8BzZNqsGxFT3J6XgYz0vwgu0c4Cs8OJ4uQBjn
9FHByZdeFRuqqNMQtO0s1vxtirqTQSfWr+/QIxn/Eua+PGWrVbiUC9ItMBhJeNaS/AIHavAU+0JV
uzYFbEiynhWJNZLcoHGp9ddnAOkmCO7LV3ma7h8JAEJVh3qIENH4+I4icMH7hvoO+HRLnM491o5g
uk9LXk33dFqlYpWkDuunCu4EtA0E0npPilSCWfv2wwpUJKP7Go9/GIQkWELUKAC7warT8s2367K1
25XwNZ12ALMcade7rTSpCfxMNXf2I6BKWUgQwwrE+9bpxC2ALRlDdnbkt2sSo5FiCbHOvFSwz7IP
maAPVuVNwgys1BSdtRcfVDG81mkTIqZfaGzUOxXmcGXy3rSdfgd8ltejKTCM436O0KojSQ9Y34Rr
JRIjTRZ5eMsZPrlPFs5KhBI+gNsJXM1SRFWT1Onb5DxmPOWO37rovIDOTUjDubhzYEXnk+dMa3ko
WFmh4nEkdvs6vYs/NmtwDrzxlVTwGfrFZhAlBgwSWjMD8itpFEdUraDUjoO8iYlRUO3UPO4DNTUh
gvbFUOv57fMAipN7O8L2dW8DFokRbLnCqE7a95Pw6GzKXZdHnbhQ363XYoxgLiSkaYOfDVgxkd0k
1V2BZV2B1IzQqnsvyFMU4MqoF3uUZB5kWEMKrC+mJLsT0PhvlcF2n5RwvU0r/HDt6+cMsLEOmYR+
in39aTRX49E5rPZz7+DsScL8Fe2W2NtVQ/ZbifTpr2aoDL8/gVpArXd52g+Z7x5b9jhJBhF4AjWu
g1mFRvEvaBtfvf20h2YC4Yq2hFBqEMX3nq/7iLueia70a2mnOr+kcU+ILVh/PdZBZ1WwN0e/Mw1P
7Jfk2Hz+Fop+jEV7d4pvBSK3Eh/SCwiI1nTPzX0TlCmKiXAcp3kVMR5fCy9hMGROHK9xejbYb+zM
glQYDLx8aQ/pN3xwPEwg1jpgG8RjKZn+YglgR4Hn78TaYS2OFmmR5nhS+GWfJkjjMktolChe5VAW
oNsxSR0qbAgvIzbotoUbJ/ozRc++nCVJXL5BY1F8qdU++j+XLumqXdn7LxRgtLbdxdpa7S+BXlpe
JQqglmlamasYZjFsOr3u+ymDvdPjQJSKSJo1uPAQpyIe4COHym7f5m5eHyWN7YQANpoYcLp/YrzS
VmxOwOfa6kb5n5wITQxTr2SdYMyOHYJ786cW0/zVpFpPEzAxBEzdodH1J/Z8qDCM4WYRUgEzGoE0
Gex4RC7/ktnjBgRl3KUV/FcCknH589LI9MQNXmf61BfAGyaRF2hfb4ut2JI8NI0oi6U6baJWruE9
bHGvJ+6kALPZYTgQnp780HUfsss/5dbt79hqh5IylJiufDc0suiSxfRTx3z7Kwevco8JR5+T71dV
L0Np3CTmrGDs/W0QYYV+uPyRGzuLd0YhwllHSSOPZdOPfX5X16iFdS8h6Z9+YzJpaFDXnyMn1kPG
GbGwfeRY5G7X36jw5PUIJSK0uxwE1hAUB708qenxPdib4Uy2wJCMt/t52ZdaqGm84W9G7YA3+ZKN
rYiJFZk1xBbhL2a8rE/EettYbkC1kMfFRYZb5xN7HOILOMvahrvpNIM3nclSd9FfGLNc0qako/kG
lsNg070Bj+880tq93u9OjTM3FXXhO6xmqgtrK9wvPodsBVK0+17Dix8wwBj6RfcUerlS7JYZyep9
EWqd6hVRf7Jk9SGWgEGLLZ62eMS2penNeJrViSs1s5rOZJVzJ3O92x7nJidY6cs2ZsTsLSpYtgYJ
Ts70voHrDXLd1IW+bpd7PApSp2GuC3hSEXtNpj2UWX8hEKchAEyl3OWcZYC/OicLFH2FpNmSe5TI
PtCHdtJIuozQRjlfcD8M9Ygj9NEPJWNtc/tqaNNeXO8CdAqPOrn40SdLz4qUaceD42dVN5v8dUY0
q03eWTk4sbSOtUl4ZgsfyFlpiDExOEL45Wgh13BbpHqAhbvs2kiDZWtBLcGROdndrl22D+wiv+QD
jlvhsScIRlVzux497mILnAJYLs/circlIkTteG7F0/XtQ+eUQUFTs7wBP69EujsG5V7b/3odL4H3
cxZ2o1BRoyJin15lQfas0cMh7qkgiHNJGblLlNqLdnvhzH8cmdMQIzvdiGK/2L9+N+VI5nbfIs2a
KCalmhZueL3ntoAKWz8zV/tgoTHbdlJgHjyi5N1Kxb7V+9JYKa4FeMvmMoz/RJcV9Xc7nlu+DjBu
zlAq5pPA2LP+ej30ELigEg5FyRBbS5V42904y+ZnDs/yf8VO99yJMU4oPooaitOeDn2INT+4RfYV
DEyzeZjNW3jzaJ0H+in45G4qMU9bknEpp6POCQooFtjT6A1ggT9hUhZ5J0y8Fpsg2djWipIwCiL9
1Fvt8zoAc0mQ4S8mU7HXH6NfksEfqyBiM0xIU3XAb4ex0vAsfN5sqnWqzLMgsz6+7JpdgzOeqbsH
+fjDwI383haZYMIvqxfRGydpGTW+ZtyqQewTnCXZADC9NZMQSSKx5AjHl/dRmlT+1iEGeBB8+vR3
pe3u6/uR7+b6n92Tgypeehc8i0kTR9BreadYZwU5mjMJfKhFm7shDf5UA5zTXOEYPBDfRDwLO9CJ
FSafhLVzYw69fT6RlXUZOHS5M8Jz4zIIEkFBAp4X0+Ds9bU6WUBgU5CiGI0aW3F1YkQHfc74Oroi
ul5EE3jX3JRMJqUPENxp6Zh2gDhBbMhTAyfGGqwi0Y3ibJcxZd3INWgaX0A3k5RAQ0Vx+IB3bRVx
Kgg4mxEp+lIU8Dlqez5+ic7RIj1c6V5GQTyavWxEeYW90N8pRxVewRViHS9ARS90lk/3ub3zXoev
lZ4IhdRZa4OWDG9LE79XG6zoVkWxMElu8scbz7OC+l5gYiRSPachum6DZGbZlxjgOcJZ4d0OokWG
9r+hWo+8OwM4umB3v8WJVnt1kUs96DoN2tnRmSiMYv8m851BTdUV6v7aCtKi77iW1umvjoJUrmV9
8T68sUvJu9xhr7h1YTcO6gJL/IX80zmSmMK+6JzOC/UC0QzOSSAqJ5/rqg9J7e15hAbCmGhvF+mY
wBcy3UHHvT4s61k1BMG8LFhNqLH8xqDH93MQ7xME3fCwqUmFe21iZ1H15f3iKn+/kEY5eHlBamix
1TKe/FfX+s6KonHUBw6/jewVO4vz4m02fGpQDjD/eORqiubTyBuuMH6VFe+Uq0gKI3S0u0PFir8A
VXCzHN9LvCDZgfOQM7/Uw2YufNiOdI75eq4W+XP99/S8raACdMZq+rL/XTw6OhV1DWLSKa4kOPrq
746TkaMA9x8zv+OgZJtmKGu/tvVp8ef6Dy0mGcfC0/RBNo/1WIETP/pzm3oGMgcHcdSTgFEhqIAG
U8+04gQXj4lJOtXZOl1MWfh1xzaJvXHyqODQvMjn9/0HTfCeNznFrveD4Y9x2vhVHchxqX5rtsqh
qVO76Ftx+pb15G6I3JQLQH3ODGsxp8sZCnFUqRHhbFzc7wUDddYv0prq9r7/q2bh/QrW4bG7qUgV
guzLgpBTtZvHUpPxE6ERM6vOvdxKiNwk8wDyOnTDxXdrad5wDykj4weoezilMn5LBM795Ic7DUzZ
7jOAXWR3kT0OFNdHGZd8l6XbwJylUtMp7VaJwgHNIW+GGxVTHLtsZpjJ+fxst1JjeDAW4Hz1WkWz
9CKM8vGqBt45F6Gd73xTHPRXsRvalzxDMRttiQ0y36uP5kJ0g1stKp4KEX1/duDvdp+khdx55GxL
mHCJH6PK3/RQmT0V7BB2tBryOWdPzeqjv1h4pANzTpmWeQTD0q/JlTGXV65TvoePHY77tf7pVi+k
UAg0ofJN6IoXDMTFAvQHxviIJvcuyeOIHsXc3uJ57x8KW9zZE0/0rTgZ3h/dQ6YBXNBCNQkmQ2L2
ztugg5w3hzyctungou5v/Qwb86W+rQGs3+lAoVpq6GAFodgFMRytG8oAnH0CT5TvCWh4bGlQlUqS
cpWG+vbAn88qm2cP1TfaPTc9rFfPCzvaZcrygIiuO++OxxIOUydv3c1WqxVKt/0WTz1IYmHZpLT8
l5sfFvUBg0clXkoiR+G/jBdsmlTr9DySG2z5cfjzjnuq+uquimMXmo5Z0+euRwMroDk2q5LMPupz
2RMh2aw9QFQgJSI6GLrz6iuB51f/4kZv315kzh4zahVTbFIrc+yg56CcUkF+2267NbAueYuW89AF
WHoqsjMumCsviZ4TNae6dvLsWccKlLK4w101fMC1btf3crfiLwpfwObwjPiNV/rC6j3Xf4Xkgmye
vczN/LN8yMC02a1NVpyfIertvnVBz6ZzNwf94Rg/PxLPC7834VyGNBRR6bUbIgwwFm/tqCEtct1W
drr6mEi0P6CfrEDW1dmjXQWaAMHP2DceBFp/Z7KwlrBqDmKbCESMoTGCxRafZbH+3hwmLvb+5c1E
dgRGk1Is2WjY1ECxozwisdAk9QKmidhBe73O89ehP6QBuGXL97yVS6e1HuFfPgzZOeRlJcSPD1jg
+oLJlkNcDF4hBe0L1gQ7DvQDnPoLliT/yA2zR/wE0e5oRfsgo51VN0Kgp5E5yYCPBf1WboeDJ+oa
C6yazFL01EAhQa8stqnXcPso2WbfvY/BqLoHiBUvU0ZEKZOQuwELdQllyD3AtsgvZ0EYfqxPq3WN
VyH98h0uxf4xEtu08rJDswHnhoAvYgYiR5rMeS1RylGdvdjmt7fHgJMphS9kU/VuO4gcBg1Zk2g0
xGcDx57XC3iICgVb+tMJkS0P4cjT303e3gdTFJbIcF7We5eUbyASeLjnrzbtd+vpHT/dFP6afQDD
wv3cP/yENOOH+iun80yCVSltaSfwL7k/ANyl9Huzbz0xFldJBpICZjsX708vqqb0mWDLAhQhoHmr
A9uMLZQ9PKIYjOv4UiLt3fpusTcvTsany0qqp66SazINhf271tujTRNWMrw4z/JDtYYqmqbnCZJV
9ei8yIye3pkOfbqRqnqbopKWXBuwhS/97CsnjM2T34gJVuMuEFBe9Xyk5U0B3eGeCdd/CzFm3Ueh
hC2JCN8YufApSi1uyrZQ1jf2swspMbwbebMzNcEfvG//3+rjCFFeKRlfXTKF5DPP3MT8SUWRV/Ao
vzFM8IJ25QWIXVXVmBtgVmXIXGAxW18yxB6CjN6gujZ2N0qh2VBk47Xsmbx67/vV1/zo56ff2Avs
CuYqSqdGjtYfJKE5uvVMvUeusDLj3sxvYCScgoQoYxZlVCdBzI4a5wWLJJctNowyML3IQxxgt+um
bUaTexRVF0f7ICApDSRDcWMf0057sx5gK+j7nQc0gf779L8XL1WfDvXb6QLq83gOkG2BjevGyhmW
6TE3zARgFavqllJ+BEix5cuz0en2t6wuIC4Zq2Zv8fbDBZbiGu/MkSlN3cGtpb+xFlD6P2ghwc9N
jGNDZqLx0JO0lXE3RzOpgtskid1c/B0cwsteXpOGNJO17lVX7y9a6qdIA3TX3mfnjup2Bm+L0MdK
75jWHAKPlWOgsFgolyOE9to75Dii5bl+ekpLtjTcZ12qG6w2TaAvvCvrMuALK+Lv85BWVFUAJuGU
E2JK1HrNw5aDoS+kM/VZQbRRZHVyOW51ugyAPiWQ7sKWh9G5LBEqqtaKGSjtDVp7dpnXxpcALYee
HLiArf7rSeonRYKnklYNEvimmzZGD0BpYB5aMa13YdIiIDIdvsj21jZw4FmLWSnYDdBwMofaCE4b
DcYf2/f4pDd9VnPNKr/ya+qps7qpxmYCLAHkTVfJoof3LaRc1+9LCSc8Cmbki+v6HkxBfIomGi/1
f0rk1kjz1cJHFOppoQ9clDaVfqfzJOAH9JZ9YsKkt1kgZbRgiXjzdwS19XG73hW0MfGFnmTgA54C
nyomH+xbO89NLJH8rYF2A7QDto/GAmxq+CIZQX7yga04irPyOd7ihD+14KrAfGDGhWKlug9TrM+V
LsIjZJUrOWSqvk1OVIAD3ug4IszT2uIV40Rwx2EEL1783PSgMyqrJZGF+q7zCCjB2K34NDyRXKMk
dTl+joHvOzT0olvDFCCYgoTA3rWOWQ+dzCd5SR5joCEIfLtPm5KjmIlfV1KlNR/HXEgbRu2eucyG
06mAsro+oUdOo2ClhTqKVok11gBUIGUGaoPQ9J9RmalTr6GVZ7IqBfWPumqFe5xeZ291PeQqZOhv
ivXoZXg8tCJRuYSUbVb0orWdLNHD3Cy3oxDCN8j5ecVFYYQd4T9xF6VndBGBisRmh+/Gd7npadDf
R9frAIQGcRb/7Wy9Ia/iE6nWlpEoas0/4o04N1j5JelfnKnKH8YSKLzqAkyNd5FlghPUYVghPM8U
okf/NO19nnpRo2ZKbjm7UD/93nJUkqsXEOwS9F+o+9BQrNrBLn0/qmdyN7DkLZhBnlCa4CdVVoUy
NIc7cAF715e+YibnOO3eurVQvhuahGS87REM2L/xTXzyadCXY2hG16ZSs3OosYu08f1+BRODI4hJ
ZIHX74M2VtyjXTuT+uVWWgYrd5kRifI/neNoFBtNMHbqvnzs7JREDXFwKvOn1rP2uanhxxj1peVd
01KF3mtvr4/4XIiODxEZeLU6oCHGCN8898GKzVaE6BV2Qfx14W4505RUuXqP12CprMslAsj50nvP
Qe5CExggJwf1+TBiIqwD4XWXGwbo7x2U52EWLkMZHYX0mS7+wFhzWEfILXInS4rYItR597yyfhKq
5jh3sADBMsEnwvgBNMgB9Y2jaNqdQe5ObFnmGqhUGl5zeT/bm3QLYGvSh92TS5cE9UsARxFvhuL+
i6q3Rh5728y6XbSrvkM5Cw5o32tN3doxhNNPN7a5FtRIMAsJvEmP4Rn9WVNfHxkRjqVrbOq1AOCr
y1SEaeVCC//WBOi+JYeu6VPzx+n5AE2k/RkDU6XNClcIi/Xvn8nqWkJIiqivQyt5lEMsza2e4DM2
89Oa+gacZYnj2QMHDj/1XvbCDO6/IfNBTsLjinIzQiS7kTYS+ze+GMYQRFqMrslMDKdHbTn2RKzl
+u4kAqFZRZv0Ha4c06rRPiU5gJEQGqhCwH29H7DKa3ZrJHg7RePgvr7GzL45ii85+GPtCKKQjySS
wxAKbzGNxcphy3s6rHqsFaMpbMuOrNJVC92pH7aa3CHO4N3NwjwTWi7uPUYQmUbidPZhjdbWmXgb
Uc241SIL9Bd9DiwEgSvogbwQ3X111peQz2FaiuGPWZBFQywMU/bpZFgMg2N5LekyoIqXTn7piG+x
ykK/dLfa1CrBxJvijYz39GPF0HrkkVbOHTMnhDhreRR3Lw2Ijyn4Ij6rEhpkJYg8OTKV7ZZ+//Qr
C7hE50bQXVp7a2t5cQuLHaLE6QAz1XzH2uZqub/cNzkEFi3Cqx+I0uca+xNsjGc+WqOG0hQQoEDd
wP7SIM81N3/I8WmSQ/afzQMReBN6XemqHDTGBp4c/RsCfHpLsEa9l0eEzxDXlFknCHhRHxdS4qYi
feTn1IGJ1iPmn/RMnaOBkKRKzqCKkD1aIc88cyVLPz3bf6Dv+TKD1CXZu61T9+qhGqX497Zk28oG
ZfUbe55nYXI0IgdGHOi7jjhj3AB3OLepdvVifZDx+3jNGSTCyGdgPado/FqhpVOF631+Uj2SrH/f
qNPt4QuBR3ypkOfgyBScGcogRtFH9EdzvxvE3Zg4HxnthfOZ4IidlmUVa54NbH391EYtqOfs9pI3
FTwAEdMml6jd66miHCt2IdCxkoNmO0Q7raNEZEbANz+Ji1g/NL9BcgOkg06oZVYuynwB1csrTIfa
H8ClUlvCpD+fyIt17rGXKQW1JRA9iD2TTBM1MbtMfogH4HUQkeRIDPXW9Zr8DmKdKmN9IMweOJrc
mMhG5kCu9fD0ckK0tZhx8SV+d1UpSBSun8XM1BrN1cpMTVeV7Aa7JSkykWRdtrUbJu/AIL97N6Tq
CVo9+s/aWEKjS9gMazxm31RM3022AhPkHJL4uGmKAckqrrPEQMyaGsP5wYd+i3CcqJZRrjSBQBqS
EYxMO+ogqiR13zLKEJu1b27ncs6r6WgOM6MlHLI7sOB926li/gN1F0dKcNAqPS7YbZmaRS2eqA0e
jAiCNPVVw+mZmghJSBQvM/lSxMSh+aRvlDkLlA4QFE//26ZFWgJ3e/qjrvOElcVtSoXVTajDlXUW
m2aEBOqUcK5f4VpvUu/Dj8sFRumnjFLBAHCFoTIiNjKRuty81t9MjQFZt398uy6tjulhpLyVGXDP
cNg5sLkVS7qRXEshoiOCAQfJyHtKjK/C1p2t5M3cNQbGH5xcZW+e7JZkkR67yqYkvvJ8l5qLlhLw
WkhJdb90GcvuKnvZp40XCoX1K4chbaVkpgto7e3Ba6C4vXnOmF/REFG2yf+zeCV5kcX1gYz2Pw4h
MzMJL8QVGhIULsg04Qw8g77uxPWs7hKfXXRTXIWeSlkktsVmLAUrV7nJXOTBZ1B8lpRVnYu3Ipt3
FM8UpT9bmbON07g7a7a+uF8GtQ60SSCxaadm0wQUE9YXjyyWsqJVK65w4mugXMjqcvmrzRLkpKv0
253arNg8ErxC/BtDThcZrkq9t1+o64Nspqb7WW4RLCUjeVnBaPxsGkVE9qX3tOeIjZ7LyIhlVTnJ
YwCoZ8eIcoT/oMCKFhAOy0X6eO4u5ljy5EpiBCmHExKlZ3JGYEeKxuUBu6HS9YKG5zz7hPPWtrr0
QZ7tTxfnC/X7VC814d909F/WmIbEJDfgGik2vp0WrHQFo+m22AhZYz3lE2YMIGOEiXtOZPMEqU1K
k4Ajo5GCkfa3CbUvNBzwXbjzRiHSnFmhkUMjnw3nRsa+NpO5P+3++8+6ZURC+3dFlaq/kyXRo/Jf
CxkbSHehrehBHQLbn+pztBO79/IAbAM6BBuV8TuSS4UOkdoh/BvNjlr/KamEI+EsXxXb1P24ZcoZ
683YcbqyzR2ZeMtpel/9SRwhHzzaIUXkt3JKrOrzm20gDpNjJC4QaGs9IOq4ra3pTMTXl87uj0MD
EcpmmGAOjGi5qY89FBXgUWCk5vsz93yalRcB5Y4VuwUyFn5Rlh9mWZKb0pSZ5PIf0TV25vy6aMA1
VDAUtmLVqv82UKx7omGed4euBUwokY53uj3VhEXbgEiY+EZUAp37xZOg80tpBtO6mgk7qCYafHip
sTazfdIJ/MArOYYrkk0Dq6Q0dOZMu/ZzNAdH9Amg7nHXKxRelJvb+mT/tLfCb8faIda0vfql7c9M
vTO1cpjwDfRk2sAL4PTvLKPQaC53CkSBE1vlolG2HbT7CEdTLSGukrWu/IxkPwirCzxQ85aspPOH
dkqQIbS12nJsmM3dRbj3lRQRC0qeb8Ufq2kX44T1+a7oRlTnDB2aWuIISc6a1Fx9ihb9B6np7fK7
ClwCNNCEp1nGXV/apvX98SYdj1PM/G+cVa9VMY8TX3jVvRydGFEZ95k//pSAcr+iVjftkcFmMksM
oYcEPAV5K6mGi5KR4vydb4CayV4wiYv9YkzpqTAllW6EJsymtkhuAtH5KzaEgQJcy4+olVUh3vte
WjSLbUCS1xXBEcvIXCBm9hip/FyXtFnzM7O29hdGEKHQz1T88kcTVEhcdHzRJdZ0l3fF5kukasNg
R3daDc0zxt6EAX2T0h80px1XsEwhaxDlbzb4Aj1BSnIAWwSITtQnxd0OudLo574/T03RBC07lHEE
pkzYrR20Yy+6INoFAsCTGPeXMXpnsF8zqETtfUppSVB03qtr+AfqqF5dT7yMx9V6W/xp/a3hyU+8
+NiR8yJBQcwLlIX8z07Kmu+yK1h9QQM5B9VagRrFhAQMBrwB8JQtaeAYE7vqEDw+RPlotxLzwxc/
NKOrsVA5ASulSE5+fZ//AdkLoGpKL6zlpTAGk+7v9XCk9ZPqUDGdZagny5VB5ukbsdTu1kQ1o/Vg
u8PCbQIsMtPEPXIPqHDkwHoWoTit5cO/zB/JuI1hLmiCshcIyDPJbVkUsw7qFVWIlJVFevra7Mut
Qt2JLFGJlAlvKCuMQ9Ay48y38WcHIVEUbA4Fv29DSW1614n8SZ7MIPwzUVpGxfVCJzFPT2VeY+Tt
qhtSXTFTuj4MKq2dRlkk23PyT14LTMjUVgfS74luvbumfAMoMRYpws+y5L+I1OoSSP9iO9yiHOlq
XAA/Y9zlIQHP6bU055oOhxcfo8oFp1HZ0F/lFUHHxVI0vMlOL5D+lHDte1O/W41WNwkicwhpuQgV
ST95NubBub4enLebFxRNo6V5/jEepW2ljGY+bKc5VOrtc2QKZbo/Ye2BVTBxlJRsqiYdLBw+Lou6
+tXgce7FHpMM7a6OD2fv6PXXvL++1g0qlB227jDEb/EqKS13jNDQ1X89HL3vgbCdEPeixVepwLu9
w9wEjLykf2Cjs3b6j7PJ3TiZHBcX1zpqi611MBu+qWZdi3C7HIHUL9gZNPjywJE1NV4kBrhbfGy8
iwTS1n1/7Z/REsBSLfK44CPaF7tzreZRjyKBhPJvuoD/7mbsi2qOgaO/ebBnNE15Z01lOXwm5DBn
/FvmYPvQfLoproA7n4uTD4iiywkDUCpgN9s2l+hAPOdN2+tHakRq6C0el1dvtLeZ9niM7893dafe
eckeCvmGkpB4erLaspb+/yACc/l+3HuVt1sqbXO3ndLVypU0eXapDpUi3NISwdIqDYKuI98T8Egs
3kYuURLMUEPMssOUz3/wqY/8rsnEldwcXGP0Oq+9gNi8MadtczjvbuQ0Ku28qpSJGRPgpPKTf4Yc
EIbguN4Jcw6NXeIqSQL1s81RLDl93HyACUnZ7EON+5qH9QiCyogBN4lsuPhTqNv0sTOm+/nOnoiw
TWAKHHMgT96OJkI6YTn/X8CAYYqNatHuqm/Zsjsl021lKxqvg60xD+c7IIQlUS3q4fP8ul9fGYOo
uex7BoSHOKJik/8g0ElxcMXT0hGUn3cvz87bVKY9awLw8s+nZxCUf8C0hDkKuoyVyewlFplvNjEu
ijkoepEPkHgLXadwXuC0mVvtG4ncciDzMEAhM3MXjeRT3UGlSgSRHWf7izb6RrYJHhB5/zuLk7nl
zxOk70jd9cVowoZpAvm0P6gUF3yNsL2M7WWo6+qk3XwG0vupblFFMwdwMUCRF8PmnudeugPIqsEa
HrGX10LG9cagC0UPZkc8HyJysc5cGXV4V8VXclHwtcXGgyODMb4hHHrCLpBLufIbyosgQHW/JUQX
aXv3+VcCZD+PS8MPHtruoAKG8086fs5KToryYMBRM7haMTZfQQLXHII4MuSJisw/sQSCVRvOrrGf
lJOlKwVUaoC22TAvKcrMk2zK4N4siBBfFQlyThu441YJN1Hi8qa+aODxAZjdEpEbckWUAXXHZ9aR
jzfupaesKm0zjtX2C7j0kQqCAIQU00gw0M14NzOeTCbPhiOqvceBlnvZ3XryuIEsAxaAfshtbT40
bmDtjOsgZjyG6M5gyJSVgGh2b0XYmTFMZIg4Zy9I6zTcdwB7FTWmbI0vIj3dRbsPOUq6xwC1NFcU
RbgV1/mF8KSuCT1NJNGum6lMvj3gSCougyN34TXuWgPTRXbuM+YdhYpOlNfyDtuHNJoH+rINCXKt
Bas1GDcurvgMVNlGFdRoeMC6beyGDflbeedTfUkQmGFZ22T8HP97AQ9CIQxCVxapy8wxwVXhDkW/
QUyV8T/44q99s23sNb3YBwrAGKcGAcIUacj8KxxVOI5xxhCk8827kyn1UNFC6y9AlZEw0g8Byt1i
jM3t4ulgDDeFlPU6n6CDDZGSh9HmgTwtKVq0HgvakGm3tCRq/2e5iIfVD/swVdK7j9Lt+m4r5IHo
YMohFMutrIC25WBDoaEV1haMMmTh0o04iK4kiDwzIm2OAXAIh7QuOsTuADpGvbgtWv0N3OmIDeM/
0xahEKyfRRD7S8qe+Vi/VxKgUD5tQfR6LS1uj/oaiPMi5CmSoyKo8zMSNWPdwyVKaG1cQWPDTJPV
ZnXThhN6sauKLw1B2eUuDkCgSLa9MsL28odk3FGzswaDKa1trrGOlYblWgk+fB01fGcQHdDIrOA0
sgxb4rGJXM9SGZPw2nMw6dHjiU/XVD0W2OxQmDV4TwZalja/JaKGNOL3B6h43VlIS7NPQt39x5Za
WGt4+BxdW3LFTG9yyKfQuJnBy//IP30I61Ic2dSWT6uNGPI3BJWMmzhjgw2jsddqs+rl9D4j1rRS
AH6MpmvBCoCwV2jJOaZc3aTiR5A5nmgkc1hyAHihheFR8e9dl23qHedhujGkbap1Jlxgjvkunf8S
+GtUDRht/FLOMc18AEMS34vxRtWyKjduje7tyM1ZFqnX5iiVJFgRFjoxyaMrfHZ2oeXt4G4vB3nx
L4Y8dfhmhkpFn2dluhM7VfuVTyyqIZLaubRv7euUQcTjcX1jPU2UV0fANLcaGLnNLQgcvMWfpmzw
1Op/XF2r4FbwCBEEJz4Jwbc7E9i/eQfTEcr5Ee25ocCpKdJjpYC0WD2IbQ+n7+HGN+5ZfMKCzLoh
9CeeNmKYYRzS011yTwC9uWCfA51TK5GW8AewTws01kd9viPD7Yhv5Qvp0RGZZmH62a+hxu4crvjl
nHedmhNHPUHUwICVQszeEkUxl3JXar7+2OdmNrlDijNaZaRb2i85PAWlZTuwu8I+jtidzsi1nBNb
vw3HQjMUS2In3b0RdkXJnWymZqe3pR2rT1AX6FHPHnLaeXA3+b7+w7WAp++HfkSaG6nmIiZ5pXsl
lSzZa2ZBC2/54oy2xrKuR+nWrJN9jO6niXeKEtZjdXwfj2vVpkSWAeaFiYpoXmcgix+FlV27NlGK
5UtBS9IggCBezC605dTdIBNC0ZEWQqOOCVhoiTwYYNRSGuatyE1OAjnpf4lqbsLC5twnojQWDXpZ
DOvqUbfi16HZGc5f9DtkjF/SNP1E42qPfWTZtkjn9UakxHgMX1ZZm+AFDuyoRPVpsE2bvI4+U6Vg
hGrIBQb404pHpuz9PVwF0dcCFUZ7VYJ4tWES7ntGYO3aTHcvVEJa6uglMdMiWCOHOntJm0mHHiYO
9mFMezK36xYYihb15ZSpQhijFfkLOY2+mYlclfZowuo1U8SejicoXwKtd3oGWs/Ed6MkeOI2FkAU
4qyfnIvktgXMbuuTIuoPmml2QbMkKejNRmEyQOXfD4EEyYfAsbgc5kLjdbPLgkA85qTnhC/C5/e7
kgPQw5B4uui00t6YI04QMUTCMrlfwvhBSQbZzQcDLyyZb1SjVwXHoRCooKAlzYqlD3Gp50UnIWbh
iZ29cOxKHyvIwhW8gZUdiAF+SnigNOiCdDSfIdQeXQeSqNXQR6BVqlciIsGLKFbU60N74FNry6sq
CQeq90b+iSu/3J0DIAjog9I+aMngdekVS982a+7oFre3HndsIdqGBGWMqsQx2SG/zhNO5iXXgnES
mifdHSkOYXQ3fEp0eLPyi7boIlJX58UWajWKEl/yXbRqXBcjWirfWkHV1MeGoekEYczuPBadKZbi
fgWEmvtVdRgGbeVPPBNMjY0NwPOMPRDG1IRLH7rcAiTxcSTyN2aaumZD9KPHRRomB5+QLYgbij+S
0fAk1udvf7jaMwP6nTo9QC6X9L4JDMS2kd2CUSKxUaGgRdAXJ1Lv7OwnHooac1/TncWkWJW+MKqG
Cu25WYwAe9/Jq9pnp542fGtVemWbhoBrfvLk93wTDO+LnOaZm/MT2ELzQjM8E9FHbiWuZfThhRZH
VB9cFPNxqXVZP01e03Y1rAh1oKe6EFjwqo1rlK60HA2AdVjCzRqx4IIpN01ARLnaHm0QVY89qxY1
X9pr6BgWyVWWqPC4fYc1l+5YNCoV2kMagAnK8lyWFxWuMWRxtYt6+lBSiYdMXz9/GSPB9yGo9rua
5w6hPojiXFO/KhLNDW5/7Svp2Kd9JHOItQE/zfqRKS8nyuqBzlbN+78NLp9NzK3K5HuR++QDgcVI
Y+/UMIdSgu/o11WmEBy18lQLNT4xaBscJ+zJhGytsCxu3Z8EawK93aNpSlCS+loMAbnYjpZDsNG5
vIMFJWngAD/Rq6VnJEJCb+YA7YoEkum3UnyNDwxDuPmHuDbBzyxziUtP29ykfAhHKulYBCs6Lt9O
cxrwFVEBkZMOuHf27dqSyBLWXKHYPKT2H64kpMbCzjUwCd6JeCG0GdJi3kxa2g6KhW8rAjV1sQfY
jgF141xMhTA5l2TjTpsMfviHxNjCCXgANAa2S95mH02W832qU3y26aMySzeO9w2fA2r1b6xqpV6k
543FWs2BbjepunM1sE3fxZXneqVLay3ELurLKywIS709J5S5exQwp6x7W9O/6eWlXtOSlgffAm0D
42hxy/U6KJmtSRrxCLBdF2G9ZPIVGDMPPEw33aWQK14C3D5evcBZbHMjT3bIwepIZlXmlJZx8YME
wyRzgg204o6Tb6hiTVQ+7Lq8U/brZvGj6yMa5WAWJPy91EePaBcBaRYtdNoFeGUnE+usEwNBwUeP
OT/uVeHAHxqJnCsUGdU/6PzGF4dXDQWAU1uvfYqOcP4fuqnUvCpnrpVOjuyZEF3QMH/6umw7wyfz
gPynJKkPtpvzpkym+WtpNFANnznOI44zHSn25Stch3X9GKjw7rZuhO0XQDcFSMwSte2AfsgeRFHd
fM/0DUfn96kAb9/hglE5LV+rmp+KW2OdkQoptARYid6Cfam6JMLn9wxXj06wCyZwklbf7RdqtC7s
3ysHeRszQRsVByFrpMdmNfmFW5ltP9guMx4fuRxK87Hc7NCgK54VWENOCsOMEbeUFCXEjFPbWHOy
5gt3+ah9S3s/I1W2IlREIkhzLMxYyWIXSFP0Ux/9CrkPbwFffoIEK8tr/qiDpg8byZiIYZbu6eZI
DJBuo5QRsnVhDiK7eJZ9C2ogQ1fzp3KbedudMWweFoIBJaVLR9XUjqjOToVz2vi9JvND1i2RAamK
EM9pmtO+zddDDBjV4FpVKL1Wtoqve7TKnGx5ON+LVJjudrq038SAH6z+OaVZQqO4E6bFnh5yQ7t1
BzuZelsC4I/5dY2WsIermnZOGUMNyyOkeaeRAE0omFOZqkihWrcEyXa41E8ni/jJpYecznNiqWZj
8RyaifztpwaWKmfpYG02ZNug/YLEeYGZ7l6uaD4LK2Fpl2k/B3O4a4/2VvA2fjHc/MBznDhbdpkC
HZahgwlSsBQOAWH1CmYuHqEtggjhn+kt/+PI57/dXb0dR5ndFZvmtntDPAOit7FfKr7iSA/vhIgh
BYKSa++/cmWnrfIr5kNzvtKMLF7VBNgjJ9MmmOiu4utepaFwUvGoOS1DY7nSqUCEE+4ud/RRtFqB
YELMNxtZ04TDMb6VYedwWVTIygZALn6AUIVdLTkWfZO8ywjvsxN5ENhADPHbU+inr4OqlM8mIsEw
rs7Wnh+mM1RWUvgqeSbq0WpR9z/TUqasv2ADiab5kevFVuDaMocdUikTYjpa9nPinrQnAxNxTgrt
RjG6K6LQSsFpdSy7f3pyrN63BxLuTxaCbHMVikIGs35W6pIV1SgIungiYCzCq++z4RtZWMzheA0z
cw4Mv7fnHQaTsqiCcsqzkz4o8Rfk2KnRZBkyuhXS9N4/Gzk4lhjVriuVyqLNCoYtKEqDX4XlWoW5
dBZlRIk1fViHMs5WtfbLzk5lEY8/nky//dlh9TbnbLg8QtieDRNTSK5ycztKjkmbYRarBFX/73mI
34UNiH3q31eAsPyMp3Hcm8H+cFGhkdWsssBWvKfJ/RMa0HZjkaFH8mXyT2dE+lOclG+tEYd9IwLp
Os+W88C3jawqp/URsNjOQaiESWpLFnOJ1yvkjsCJa75E1KXS7Jswwzqzx8UEnTPPf9j0VJ8lgSiV
ORKdG6qxD5pHDMI7AekDehvW25mHtOnd8UVu0Zzze537UeJWSbyY0LOvjzQCjrDB7g81hYwKvDBi
uyClfOicMs3G6JBsgRWEj4x/ELnE0VpzlLIXZvz1TxnA5lobfRtIbjJ5FUhiahoSk+fj75f8+kKn
wJn9XcOA06GnRT/OpOoR5Zy/DMcQJ04X08kS30LI5XSDfoOV34Xa+ZqlrzKlhstIrlNLihdnh2Sz
7POcPYC2SIPaC1XAGDonOEcANLu/CXoCdH/H5B0Y8VgNiDdO1pQPrYS+plBFHT6NMXTFhse25Qhj
0tLBqyzUvjiceu9AhXXB1a6QNSCK2FiDx/iC+BQOcW4mBn+aQAjnHY+8mBP3kJym4QRsDtJ+Q4X0
jrM/ehUvg5F0rThzshxQAk1bDXltYUaaD64OKlLSVJUYlmyaVMbOadhSsbtYFbDH0+8eG21TeENl
BvW0x88ynt1JVNR2Pi5bO3/FwiepEZcvD5kokkqP+Ms3Oudi07C/ZlOAAytEmdy8T826yL/vYFCl
fU5qUh+WpWAXQ9hkOSukdCGSZgGu95F8roBcpYZ+6JNzQ3Iq996AcXyEPGp/uOmfDgwQZHRg1wQm
jbxIIGYw61W08owg5Dv/MSOA6UGzDqbBNGZeT0H1XHjLdrG5a2D2AOQmh7mH7NkXfg/9u9ioFXPx
FU86/QC91bdXb8b4SFIGnEbsZC5EXavkskdcb3jXc5swQNCzLK2BAbc4Nt7ZiLhcGsWk7/YvwA8G
lgGgjbsfd8G9xXidQMIerrXCtYgr3K06RhtfZ3Ep6b1iMrIuzhvwih1jRgAqlJlxHaQS4yc2UOo6
yufqp04gS0pGjuWlOcNXoQhI2PESzdZeP+jIY/y1/z+lMpfCLbME//Yq8i/LzdBAA0ozqAHgZIFD
vLU3rp//2+cVhVQromTZQutJmIQmBhfW/8eu7pUkXUtoiB3mVHEjVKmXxUP1MLCKURahpgDBssd3
+vRNT9EE+xYUMWArUqmRCFP5JyvhG6oB0qxxIC9U3xYc/m3PJC8eeXVfmY7sd2oq3a5R4cQF9B8c
AUW6qbCQG7TEuUyU7kTHJIThRG6Zm+no1GGDeTI+CvrXWoRIAx7heCaSTTjnS8Y1YoYtnfvnoIXv
IPlPMxKBE5deHJ8WJAHWhW4A83vjXOu8HBasXwXwaPSv/eJ6+bXRPnOomO2b4MdfVpQN5bY7ZWMG
8U3wA6klrZe/NhkyqyHKNP7r/jOnSqpPtVywZIyuFwXh+ObZsp5w//MltGu7BVkOf7oLmhv2IFOy
vvc53qshX+bHGad3DdGAchaW3K1qQxfvhD+fEwgsAkBeNn1kS5F0WN/uLDTzwInc9YdkH22wPm/s
VjtnmTmIzTxHE8DHitrtJxcrcR+RQwSf99O4ob2plPO0fSXrKxmiWjvghIQQ+7OM0BcZTo2/cWHP
pFpD43uLG8u7FnaqnsTKcSnbaOWhxHNv8VXvPNF4HQmzlNh9da0qZBQLSgNX8pwsmmsyvjDfKWDc
qmt+WQ0OvFETssYBR4weyx+YP8LvCSZI77Fe/311fg12XH4cSFtKD2V3bjHHbAlWRlGcPcOi6aLp
z6SOj7/4B3HS3wsIyzWPtNipQI2Rb3NA2tRqwB3UI5s0CtpFcxlyi1Coj+1MHcruC/3krjyJD8+N
0vsRbvsLXlCDRyu2EsN5hvWnAF9uNFpgg8W3FVph6m3SdjVQGgKCWgraaGUJ0M3KASGzyyHOv5i3
8GE3kXULTFeG7PuRDzkPHdj3JIwn0J8fECNZqFyjJNq7qdj2rNg/s+G2r0aL/vxrR0+962eOwVVI
eG12XdwpclRmhc+N/NpUlEeCswK4sRGa8HCLm6kMDfNFIr3n0kT5EVVnTcV5Sa+3Eba1GELGPyRt
aLWD+Acp5yz0TqRHJ3TYkb/+FwYU1gEsqtk1BEV6/EX7B3QLPH7Bss+GvlzZ5L2yZq3wXtdSk6RY
DxyR9VgHx8+Wu2VanYSj3KxDdl4fvX5euI3aW7BrQ87jWjjE2CFoQw5MaIwDaKncxxZx6XPWT6Qq
L28NETeT6Z0jLa6VhMKRkI0pIrUZVlRmmqjeZr3HRiKK2Ca5kMWQxx+UuyZVoKvdPWN3kScr23CI
fvKqwitcviKJ9ofbEJRauktWysXu3ciNUxjV6uSXeZ0JPqeOz+QD+XVUJtFoXTuoJ3jpX23xrcvV
uc9mRMDOD2VJCQZK04gkQSMO2PKO3ytfYkm2TtT1lPfYqbHgICbmeNM4BwNGwAxwYhwXEul4fy56
N+o7F/pj2vDvW+0wI2dmYq3iw+lfIkqqbE4LCpg52xloxbAFu6ZICS9EHR1JlCstJXuDPeQbUrSF
euS++jrGf0H7Npe6hDvrofqxGl0/q8EGP5JL5VJYDs00ATQKpowyGdbdv+7f8etuj7+NAni62v8x
w4ny2q9Xw23+aCjCs0E+QOYASxW3c4zzmxxmdeyvUR0xSOTkAx8aCBcaA/QuveBgR1quD6owenMO
C5n5vhMIsusFzDv2SI63e9Fqw/oMvlAzy+AEadM0hfDtK7F6moyBm9C/kKjp0bLOLqmMt+HR3SXo
U7NngcAgW9h544les+XrqU8sB5e5cko81TxgRY712o/qvnoelhOGWdRDRCrNnSkyld20WICtEBs8
3OhmhcpBeDKUwT5bGak8Q9I8ZEXzXEWLz8FiARqF4hdf1dlg6LHObiPrX5Uod6tx20twhc9oltZ4
xZXb8fv+QgNHEanAANqJ4poBhYFHuvtbu/ev2xaw4VnqMKGlFS2aXygx6xtLWNlrF0FljpCLcBqQ
Nqn1T6UFutrk4dLG+pHK3OSJw2UUJ0ED9v11+e6ig1Oh57+N3SHnv1RCEo2y1hZZHgwhmFdCaJZ4
nLLEb2m0WbMdqbpyFdhMsGrr0SHGVmq6sW1yQ/cAdsmmkUeWED85g6pC/U/xcI1WnCRVu3ZUkkE/
g+zvNOhVkAVMXk9INY5Pv1VVikFO4DjAn6Yq6PfdJkPTn0pgWLvUmTroASt5Mt30DtpHFk/hoKxD
tPsiUnaGMikoOBFt3LkPNSxye28Fm+NS+d5F2MBqe9ZTwWq0ggax6GOz6+DGf/6bi5VsX8HfsP93
mJXCULVH84wg9+P5TyD2fGMHcQBusxcSsai76gCS8Vhg4KkcQkgPh+LNu+QyvDgXnLTI20Gt2N4W
wfKY5q6V6QZNcuIdNLJlEoz9kmwkcAI0RsxZagJjpSDuov0DFSHSJTpeV2n7jXh3oXrHWw8Xcp9t
DZ3u9f5qmjQTMacYcBH6gt3029goxjeJOt57U9byVeaGgw16RokxP66OOkeOeYylThgsubTUWgSY
Vee69l6kUm6SaZTvq4FwAiS+Dj1BZWVmcyNayzyXkJB3UVNfGp4MjCtWFWt6cBqQ6TdpZizCgy4/
3KAPltkPP6RSTmyCZhCdlIYKlD2K31Grswg+/BnM4O9dOIl4sY1uOorPCHeKHbv2KqwIkEpWgFDA
2CW080xuQJyc/IRGtx6lwypZT4W91t9W3W1F/wASVgJBQnWAjIKC1pkD52ahpqExuy1TDqq8oYPW
FNfE4nSjC3EdG0FKLy1MpclUwdl7cXFjhQU37wz2h+dbR8pO3WEAIMYUIKQAY1Y/gm/3UV3V6Ho1
SYDTpFWwYNF9hDUEsMnpCkrovhxIgzwhtRjrsYZkEgWVBn1Mu56ICg323RQv0lquk+PtMCWpuPy6
wQ7+EYOCqWptzYJPLF4rYr5KmMnKUHXXbL7MWnwmerzkMCeDMU3g+PpBPoPpI8HK4DylzBnEm6ma
oy2BVlA4WAfAjJdrNmSLmXVi7G2guRS0h5g7Bn0SJFM+Z73d7wF+uyWOrWrX5OuyddL2fhVQaHXT
lz0qsfG8if0qtOtxh25COpQdeKuVl6hJNBzMPhtUxnsoGPD2S9wfRJEGbbH6i00UP27DhFXJxBrY
DoQkjDOen+MEym8i0/XJX2MNopj7l9hhiQHWKLXNCmQ4rdfXGIanZM6diZ30zaqJwGqsJPnyMjEj
lbqqqQTo1IzWHjkI+OhZrTl1btKkgL74tKrqyBwE5u8HfdvQRjYVA5PWqVED0y26YQUYhHxkQe4o
EmPADk4GYC8jqd4skKKqsNrA00NlOGnONwSJI48eY3g+HUf69tmUq5kGW8iXWuM+siWWuXTGWDWu
rZRIxnaL3gOUYTHA06/XvOuDsonqSmPVe4PYGz+Z2xG6JsbJGTJtS7D8sGl7cEY8czTGB2VftyR0
9KOI32GAADMVCtA7DqdcKasS10Hbh0p0lEkfUwvYgeLWI+MfhYYcDCqXFpNCrx6zxZB1Qsj8moDV
mgacw/aPDHgpkgaOGybKhvau8RtKomdRcHtrRVBACr5soK5ce0tO816srVJkqALm56d60necPs7b
8wpb/x8HRYrYUZw3kBdFTngSMwvG86ZsvBJXG+Al6su7XhboRIt0VxjmDmK8MPPPMeeci4Vld9+A
pC2keHwN5DkrhXYDYM2GH+Ni8BbihaaXIVJoPsyd7qUjBqRHwd8jXFRu8lN1Mgk7umMDXJL0HlDP
yPdshoQrYo2acrn1kHWnXjmrF55VZ9AVJwDaInnjdEzhmVCy7urWBysMD1bstI/OiMShkD6yCEs6
sJO6e4X7v+jIygAOtDaLqi+TBfGSHB62eribVGWfdgdLL7dWNL6v5d/POfxn4S/n6u/VVhsB5Cge
p/fmCQeRGtCUVH05/M1cG7DstMbz5MhMSuqCX4OPZAD/OBMBAoSbECjHlZAgWX2ssPlZ71fhYzFl
ouP4FzxdjWLpyH3XPgP2J8VvCU3REOTBp/ZgzIy2FO8pzGCpqivSCy/DOMN2R+R03PjIzTMsyDFM
MH8YqK5yqnAcoLTJt4S90TgomPMzn6RwjSSM0/qGfMYcf3z5WcTIuIqNvYoeT/MnD440hFN1pB9V
UkGF/Xw08e9N7Oa47UKbB1s98xXyOiNo2oSWopoLX659Ued/wWSnZXYP9kQxfj9o6aDo5Cew6VoX
ghgSD0RTeVxt4v6liCF49RfKwb/CJlFbQWBNRprQyV659L+mAD4K1349uk9/wg4TpYgKYKyQhQo5
0v5s3QsC6FlqzmWv94HdA+1MKagLzmULbQMujkXOgpVKqESXjiE+zwHhQ5Fi973rMahjbVG3vTFQ
aMptdy5L2GSACU7p4lbUvXy1Tttdc1eEmc0AteFhJjFkqQgzPwzr39PkFC/Ek89f7YtewNt4/ZuW
Mas21dNNfVKK9BAHBR7F+FkdgfTPCzsnv+9KdmPLDaaX5qLS36BkWZegrzfzWKGJsT6UR4zcbYpI
r29mVBVcjpKFCFj9eWc55TxH22GDyYsARbqwfFfKsXKX+tVCK6gkya8gPwPs8IuRXE9AhjHibLVl
u6lbXXNgTMb5kDZkak2FC48HyBp4yJqKkaoeDc8/PYKfu+ZK7P2nPshqm9kxA0Sl45j8hc851zN/
gEFoQfV6ef7VuDc88RE0ADFTNU/DsFjYJ/okVKJMBKv2mRyADmdesAyDflJbfKseESqYH3KkXKf2
gsX0U1F65L06GFWpGkhWAWnMT2YvB20X2Ba48QKCUKF5iAZ+RfhrFfhpzMsMjGxd0l0aBnYWiLEu
f40G4kMtHlwkEGu9CkKH14mn7UUtEKYkAeNB/rL78hky7a79d745RUkaAaiyZjaLQA0LRy+BKKMQ
Ivaym6XHqax7beS1ft2sIvy+MsvmTMd895AUntYkRtj4XCRALqOQ9U/Dqdtt8a5YQ5ODQotgBytD
65ZjOzZhp7AJqe5UNhbPz5GcgSJfdHPda56sCSZx2KamUXD7D0Xt0K/Rad9N2ZYvcx5KV7idHT6V
7tLzH9jE1muvX8fSK9v8GozAjQ1urk9AZiBD+ItyN5oiaDrfh6oPkT18RygdQQMtn/baqG2GxwHa
Ovqx09NwB5y6J7f/EnfCevTEtJEHvMquALhZtnO4qDycgmdqM9R6lH78Rh+geJJd0WMKN/TME44E
FIcgMz88bYgZpyX4HPONgg17hAWh+SBMtKKfUvaqb9EXv512zvqilqTOx3HP9JS62VSog5/ObWQa
tUPSbkncfxDfaOiCA8CsrGSICGIap18TsWfr8P3o9iEdEM88j1CQ5RLHpGxDn2ffYfPZzG4kGss3
ZiW1FH2IDnrjFtwH/omle2HkQNNdlQW4Lf/G1Aehrc7ZklD20YLWAEN6xtgpqh7MXcPp9LIdXAcd
fH+H6uq3DKXtBSeTAFaUFElDFgUlK55crt7YnCAPLco92WywoTSNSAimvi2tHD3Gd0rZCI9JvhWb
4wR8gQscYPb/hmNvKwBZOrOY4FYEd9qPvEQ46aTLLVMBKb1kmDqDNU1BtBD+4BdEAQZ5H/t/IdUy
Iisp9Q8lYdG/FjWKyA4I/HtdT48zcTkO2dgnAq+XGvvQSyFRN4slABnbsJJuU84O7/IKuybGfW3Y
5VpZDkWZxr1l1uWrJkh+KyQbbdm0sINCmj7waYzboMUC3IE7QKcRokddRhBsOh+rfJ4KSfSyZoXM
CuEjyzdDKbe+5lEx+ujfsd+RfcsSJ33+5VTo2FqnzpIoMV3fxMBiuL7OcP1lQmL029yn18oY6O0o
fsbm4vlADATBFkYZIwBrCWaHCn/NsVttdnvhERnjdlMLH/BxPfUqp3ACESmmJgSUxVS3DF0OnRYV
8DaWPRb5C7QQDEIWF873VBHDpqi5mVTENLmU+2zjqVkwYEsUoupmBU7QeWQ1yp3GRiXRxHbhhnb5
t05XIFlj5L8g8xBf8w5dY4XmnU3kAsxfgRjZjRlukRhJ9nBjsnjN73/CQ8UCYsSrJpZKnBedsTrw
Fkwp0n2Pgpf+ye+ROA9S9RlvG4Yg4/v3Lxb7eO6OXz0wb9OSIeo98HG+Y+W65X7UnlmND9MQz27y
yInG6Q1dIOmTl1QtHjd60ush96zhDjLEzp/6/8pjwU3tv+u66r3boshKdNOY28TszLFUxQJrOEVH
p1Qx8psZ4TAiZ9wnpdLNKYCR6D6pmyTIPkzqKuKLnh3SmF9+C7wrD2e2fd3UXUAFwxtMMbquqztV
axpm4VokpjtVgJqylXzgUw0TLexyG3DS/NRQormRw2Y8yjDG+xuVMTxiw+LMhWZ/hDVZaYdeGkQB
3a4LtLEHzJUxXxD/W22y/AR33v4+K+0XUY5UkBX6iD1LIymz16FuffoxdGQ8SXMmlT74unxNjsAk
iduS8eja/cnaH2rCTh1yu2+1Olo3nt3oEDSIpwBwK/xBCTxteY1XsDctpUTEvhLa1x5opbtcEMKV
V4zeQXSEGe0PByciXgDS7ZKIR5zpnEl2lHnS9tl2IMm2Yq5FhjR6rYexymoc+m9CW6tnMrN3OWcD
uYJ0266RWfIYyP9KATEhtI/uQMHZ8nayBpk9Az2pRWCzmQqUZzIhLaZJWpryS2uqB+gqi4RWtd5W
cY6oOUx+c1EjDi2rcBklW1bJubyYNhGsnQGl9DGppEnqBoPlIHjHCAVj8pz9jF/T/Lv6o6k88+c8
vQNpDmXDYDNjibSPHNNmUsqzaU1utdAqMnVWoct86ZZrmK8GGPjvXMeHjHPfgUR3G7dUdPUtHtVg
cYwxbl0ZRL0y/f+AnMqBl20wgf8vtDWVu36h01dZk6aybtpJ/3h0SGY4k779OndNxgwwfUcwE1f2
fKkbu5TnkjpjDi4mXoV3z8zyvxuL6AGUMg2zLoSUIdOy6sw1lIfn8yil8LSKflD3qa4KTUTmOEcQ
FeG0tkje2aKeaWQf3k/m3P+RKgS0/e1BgQoTQQJhcXeF9OKESVV38AOL+a/ji0ET2+6Oel/2aknB
Ul+mPEyBlg1SXKiw6o8EYX3orSOIdlAzuw7cUB/T9ya9FLk5OdN/qodYXHDAwsb1ovutxqlRkDSM
4rLMAIgvyi5+SJg74rsIHM8vhHn/sknwgiHTXwwgpO4N2A/6tv/Co7cclwtvbrhjgUGAioSpjPi+
hXJzeYVtbKD6uPP3xo0mHINexdyRGiLNgaKsaMunvd9xyYkOkf3Ce3/SQsGLeD1wakb2rBVy4reh
HAHd4Gq9/EVrcZcdRRBhDiVGJxFkZHY9gPSJzThqj86blKf4YL2UyF3Xyp8h31SojQK85zrI1Kpm
pgukUQYUjV1n/9eh99irWdpcho+H37XJTbHrGIURdr9JVZVibdcyfhCDsdDljKRMrIe1ReGXkN/t
U3l8EllmWvk1y2dUqeyEyPsKW0+NxswGBG4x1n/+Xs9WWIPVbg8wdt9vhwr3Sk3BAjy8F/g5Upc1
3E0XPlT5lP6pllFGdxFBkolY+hDqi+FNCVppQ7MlGljE9QpiHiXSRPzmu6NWdr7CSfbHQx76hh/5
Eo/o6JvtQ5/CEzkMzL/TUFIjD8EQudsSzESV/Go1bPrlrlMzqVlCUfVNbojOM3cl0jLmD/GW5ifr
bz7VEPCjWwoOb5Uq90dSMjiklziCWo2xzeKy2OPOSxXqJ8pSe7FDyBkzpTjuMp50THJ5OgvbiXz8
5Zrnkpx1nnC/ys8gidf/Hx3RXQRDbUzbD1BSfC0b/YiVWxWg14HzPhl1B0mX8HZkoqZXk7YQ6i/h
NikkbfL6lyE8tixygufV6LstFeAuIxBBwAanuSeMZ+CmyMoYwcDG4QntZCrYO9F50qFKo+cv1PRl
pBHH4TH7ohsqSfX/D9+DzBcOrBf5oiIt2uHCS48jlPNUgiB50mlzTiiXSAKGAkG8ctbiWmFWOP0k
jp9cko0apWARshBiffknGvaProxU/EzAPRez3RZx7UbAxHw1944VRZRkqvJ372NBGqLUCzqaVGAa
klHzXuzWuKNyI6zKDqWlEuHmiN6t+EbjnbiKOjVEbRd0bO+Sfp8QLc7887eGH9QMkGLUUwgjPgMP
EmAj0+8Gb0qIXGhz3mQbbwRGEo4Y08qiNOl5Z8cEehIfepE976zD8yg0eqFUZ65O8shBZ3+FX1OY
56XZm3xyJqqY0QaDAxnCrYm+sFDULBuJ0hcxRanee1wtSaDUpqoqRep0zvQzTQ3F67lyYGglNoPL
SqdhbfgztIjZPygSb1dpwi5pftFhs4f6yYy+WKUhvwK86j8MeuBgU+h+Vf/xP+Fta/fO/eUaBRUu
xM39C0gF09GAd3utv/s+EaTwACM2D+WMLR6iGUWyDQwYgNsHvel86GSnE27+P39BujG/RDgEc6fy
808ji6jAWGeyxClI36KxW2XhJNmt6msrhL8zLMGeuDsgMhPzb6mjSzzucy4flOPbC6nz+n6tFsN4
5XuIlBXf8glg9mXHhie4K/8yuV/4plrwRM89OXRgwGyexLZWbputaRtn75L9ZRTK8FJx7zJ5PwLl
R2oqHwpCjq7JkamJvYnQqdWS9T9f5Nfq47HbiVzKtF5Gz4sYEmNwTDNDH3geJTruczYCD8fuA5Sd
DzGldNH+shFqfKpg1dGzXeXJ8jEjbH2Y/FmpVVpX7H+n3iWbUhWG76NsCbhYvVgZuJjbJSgWV61R
PqR25PI+8h1V3DJKMoq3fytqd08Q7rcgtclm0x9JwP9K5xkRMMd2J21/oZCi21qERdXHFs05qDK1
Y/9KoYZLQFuicf/MQkXZ5UMD3BOxyep9R6niWm1aalqBV6zUX0e6kqJDEdjcVPBDal088QEF2ati
Fu2vDY4fy35xlH5Db/5Rcl48PHXZl97BkyIGBCpNeLjjFeK5RnqB/eiMnJ9Nw6oNLw0siXtt0FFA
z0pOE/lWIcAhrL72jtCQXa7NUiYnHZ4S1feMbfeBI0zPdCvrQHFm3r+iwdkqV/rL7QioY39FTXkR
H6lQixChji3OlL3begunZzeveH5p+M1jcwGaqGpw/TN+R/NNhwBBRAktZ/yydyqjV788RMyOsQBm
Il1kJRo5rZ5fVYEOjuhd18xCmjT2o2bMOVi3Wm0Q8V6CeDtWR0ECDokqVmSpnGxW4QX09Qy1aUjm
vqwajFoAo5QCHJftElURzZLX2SxOLOZIkAr41CfXQGIxumQ1xfu0UpB/mQ78b0ncekiVAprdD+Mk
fW464Q9/W7CHoSzdO5hQZfbWsbBu9jclE7v13ET1xlEP5eWAme1PTj2Qyw3W0PQb9w94N/ATU/nM
h2GFnMXqo9pWCMj89+JnxtmuN4BFGrCY5EDV6eC4n831dY/+GrzzvM9sgegsjc8NUo4NfmL6ElEo
suJyqkfu7qcvdZrnzXBp+SjCjSJ7q5xsyAXF8hhGA0HrYuZt78adpERNzmAOdZVJlfVDrE+buuSf
8lenEliugJ7tyHNgncMude9gFa1wVWBbifmHFR/u/LUSv/Mdly/Y0pexFhKE2/tQ+EsJUYUeNp+P
mRgEq4X6OpyqM7mZVhYUCelF5K57toeRSQqP/gvSCcrpgt9G+l+UtoJ6LzzrBSsBVAnk/n+uqZRm
MhciUNuM9va6uzR/rgmnM9CnsMqAPxvgmnOXPxO3i7/C16zjDDn3CRmce0DVmuv8KftUERA2f+55
kCt80zEQZhmHW0Gl/RMXfzE/kIH3eOHWRsXgilUNrwLuCXfqAA6NvKEzWa7fuNa/lWaBoqlhvIqf
abmWKFX5RWcP1IApksB8QHMewj7h7h1ELMW/3Id9qNssgzHPYpsA2ORZ8bA55aUSxQLGi4ilONaH
el0IjzsGrcsq9eX8RLJVZXZYKrbe6AFdOLAo/95GFPBfYvNqmd1oHspiaA5a2/fkg/mWVlP1qkaw
ooh/pAIAZ4OKT0a9hSVBdx1TgWVHu392+XzpF0aQyzN9n+1Buddt0agwsKjpsqQokSr/5eI+OUBG
NlN7SI/aAla6MP22dDM+Gd6VuFJlWw79dHSpvEKgp/lH5Rc8W9t0dpjmgFAbSx26VDIptYiJmZij
9ITayjASm3tp3jIv3T+ofKy4Upx5QFC7oEYDT/tLXHDBcJd2e5GwbvdJwrL5wedvcd3lRepBf+16
SELygMkL0LnR9lAqgpl7LKEQFp8sStbgL3/szwBh4t3uf3yny54n6WASAikTVZNQnzjflSIzEWhK
IGrLV//oLMAIhYgTjSQtste3bfAOvW2ujJyxA+BFt9lmryZx06idqkGHKEbaN33az9Tv60RujAlO
9xXC9TYNz6Wkqr7drcaL/Gi1z1/sX0cIppW8sEEwNRz/W0wca+iX1VdJVPMvNDErXy33SC3u0l8J
JvtIWAr0ZJJpi50SuNoPGh0ODrBwqB98dGDbXdRDVCvauQwPmpJ0eygTnFick8Yt3xjGDe1ynGyX
SvxifTtTDnPqJYeBxEgKNoqHOmrvo91xtbiIs1Tbn2iWBWfxeZwcviz2uCXm4IPFyS8ro57zthkq
IYy0Qt3UtIYBCVLnw6W1IwlY8t5R7MVIa1tHJPbBPc9zVWGWn4aHu4sHG9/jDLJ5NWc8/t00eftk
RPIry6wNr7E7VH+9iaehOalxaoSHMsKyPLgC7GFXTiPg5DBWVcRgDmhe+LWCPYKsWb5DO2zocdpw
h9FWYIq6GVSgCsUD+67vLKPTR23ljFSgyZjS27nYnPoHA4Sn4kL1FIJOPzGd1g5dynmIsttqtFo+
/vACBo0B21SkhOK7VyqODhbU1FskwZPOidNUVaB1Gk76Rry1fA+/wM3s/dOIIZIubvVy89u65Gk3
cuoaBOZD/cluasOq+qJNTugwkSk9vE3u8AKWMQ2JhbGpUQVReLYjIe3dSouOtfo6eCK1mfasxm6K
cAu6Qv7hCIOZ51nvBqkQGltkRBO28oXC6ERr+xGFqPBcV0mZvoNvfmRD31coLY4Y0uf7QhZE45AD
uHJLXxdOtEf0mWP71weXnMVC7Bn7rY+eBRyAYqp//8Bi9Ms7Xa08DTRs+8ZRolXe6kSLzx71iRGi
/geTAltvEhqP22b0BAtPdrSCn/rNF2IgIlEbuYNdYuTPceCQf7TkZpIcw8KHgd9822gvGwmEbU38
0HOU39TxoRHLkeGDII2PZRKIlw96mWF2ugyUxju/sP80xWydi12zDcNtDPk/CVrPnBylWpDPtKJx
6JOz2UmQIAa59XseN8neo7irIcoxDRJTgQNsvIyZl1S+FRkgxbjXBJWPy8kop7FCAnihIFfU3wBq
fDLimaJ6u/zQDYow56U4ME43scloSxbns9wRXOx3FI/r/zYCBAsjCJX/E/hhzdhMNC6H309g3/nE
TWTAJO39nuXJYd8P/8oc0TgRwqRJ/ajVrgMPvlAoS6xKgddt7hZLU5WS0hgWaOkfg6T+GAXHlYtp
DdZiMOHVHaR5cXA78mZIjwWLfybuLWUItsz5E/XD6JyvfJATHgEl+VTSflgmtOWzfFeGC3Vgt8wZ
ZoTqwyEUtC80yO0hn6ccsTjkGagVon+gbAW9785U5orrNANa9OTBRNtaqPVObbLHpTg+FCahuK/7
T456nXcsRHC7Pkd9mZGGg0mafx29XXf5r6dskPF1trSB1soLeYlLZ+4gMAbrs5XevfLF/Sv60sVj
z7B1LOGC07ppXrobJi78h1WRlOy2qQ3ygD0j5ABx9/7rDLMQ64WoQHL34zUrNFB7lauYoYqNa/TZ
1+iFKxDQp4FFQxtp+pKGJ6uoI+vRiSfxRW7VdzRhe4QyEmiFy3FinXBHcSzAN3SZMj/4goQU5fEZ
z8T17kHyQ8/KGgIUrGzMBvfy3KUTDVf3wk4rDcjujQPyHFidW8A4R+/LZ2MxBq/W0XHV0e6hTYDo
KO/HunJOJHadC/e7VLCcmv4A2Kz3JWzdfWCoQlGnSMfV57RQPMDeta4OoRu8NqcjyiaF46TeXr0h
yqUqzpCVzp7evcpdbag/SaokzYmRHa+Bs/jdoEae3hPC6KD+7WI3yFtFbPpcdDEYRCSDz1f1Gq08
5AwmARXtoXD1ybtPRnzT4ETuGNL+vxHCzpcXIVVeuxbGJJEY9PC1Vdk8gYnApQBsJgFwjzCH+0zz
1B9BeqnZ/TpXXnxdzNXVlHhVGbYsxitWEY4tvYrC7BWP1PwPOwvQBgaZRYXFJzxjLlWUT12V0mM6
GqnGRSCjo9RfiHA+OjG0rcMe92SCSIi92/nKahfHT1vfCpiAkemomqHq0pFHGsi1MdPZluBRDrE9
PhXlFSsiRqbPrphbiTPTWulHCiLTbfLv6xKtSr7AZmftZvEAh6KXVG5+bLDIcLrxPK4tP1nP+kWG
Jr6g+6tLQACoGxLYLcy1GYQadeLw8WvttKIC8wXjpCmCNV8dEqBw+Ieb8sm9OOVdMAbWmYqx0W5C
Q/VMO49AF+Jv82bzL0N8Yj8bD/w/8trXZ4saKge8Pr6ZD6Iv3WYgqHVeUWnw1hetymPe0+xTNQpW
BpWJtOQgWu8a6+uZuieUheNYG/G6a+s5gBMKB580SuV5qHosJotdHINS9OHgB18lZ21BAYH6DSer
rRHpCC2uBCdISMgmHRi5u94ECK/X8x2K675DJyOwjQzroBjE5cTI2p619zrPMUPgLoMJ9D8axeyR
PQuzpIxjYBdcc3xU0xCR85vOTQwzRlBZaA3mouJbxtYfkDg2+VsI8OYp3xxgTh2lsikHu/acEod6
P5V3YYLrAU4QT/Qj1zyjfOPwFNZyzlrkdHVobXj3PsC81MpsP+SyDhJtoNnD4knUvaAmV2rXrqGc
gdcssjlwbRQ03JeVOa7QbzoAFXdAE+5EtAkxzSnixyzBuSo1BskF5WnAEB9eQE3QVPp59U5vEmTA
+mx+ECAYjHUQT2mS2aHS8ZaTN94pNsYWTA2M4D7ATI49H+pp935QV8o09ClN/EfIwkIZuwFu1k27
CCnfZvUSN8bFJ2k8Wt+Ojo7zWaLBPhCbRIN7AGvFwg/mxKntJ9ljEHWBshsiC5+jUqoyNOCMnJ1z
m80bnwK45TW93X+0PoGIhIk6Mi06fxXn8l8Q9HeujukTdW246995KBUvbmTIAs9pydQ2GYCg/uok
PAT2Wasz6FORVXcRPTg+S6zTPlezx5UpsgzghJbkEU4YPgmZNy6zTgP8bhN3OFsjYOR7TmMeIKcU
UUczScn8wPUdWJmvyCEl0fATluGJOEkgR9ha+AMsOH/l9WVDvcKl0RvnPSdhl7/lg31dS2u3LfDU
zP+u+HhvnB9cLqMXCzPEwNJKHfdesTa8RaN+Q4EfYTtG9613EpSFLdF/qTUwIv5By3syWE+FGsIh
5BsaYuy5Qe77sPAKShkkR4ZiVQJNMcL1sNg8M+JnzoF5y61gZWRMscuuKE+rRbsUmHhl1WxIxYyh
2nccrzsJjLgYKjnA7obKUbyfcr1d49fWf5xdUrO7tA6a+TuNiazs2JoQwJwzqgNOp0zo+1OSHlBP
HjFaugOehjG3nZQNeFx9iYUBMNhTP/PvaNTD4NPcdaIPCo3IwUVOIcMhg5Y7QHA6NgMyiV9kFjRR
MxHuw2mi9VKQotyO8OC4FWF4sjuqK5wr1hNVVB7havXHE9g5U06lO/l3cSM5OOkr/B+b2JwTy97p
tkt1aKWJwvk3yxitqMsmL6sxCFMxpQBRfn5EhldryMseYwxnVN6NaHNbwdp7jsjn8MviodCcL0rZ
aki+tZpQcW4Tl2qlpFMJpnTcVbQWYXdGyr4ONDBzadgI0jqFPUmdSunICF0mGkLX+VfsFuCP7eNq
NumfuqH5HmKn6BZHLW/iY8UixV/egIS6225s48m1TdN0SIuE4JL7pfFcbVNBrxc+MEVVbZ/NV7kh
YRsGnt6bivxCJfDbDB1GzUM6JPrrjatue0JH4PNWC10v4fnB6yyt3/lZO1uYuLBzAEEaeae2FL00
49M2NG1KJRgTmt+/amZcBQLpvgKXCudILbLpaskufOLRa18cWpQwWTeMqsUq0i11gPPH++EkUlwz
pPJgTuW05WZS3P5iEleggr3ZVPBoB2LyGrUcTY3lx0BK/DRc6IYHp5qJfuthuCo/+2/n/ClAZ0mu
bKWJpKvPfbD78HCvQiicyDclcjqqQKh8k4nTqU6osp+OssDzEt5tWpiz5ilITFYuoPKt3tpiep6g
9gcBIH9oo4BFO+rnlF5ohxkSc3xgGS02S4E3R1RuJm0Qss9UdscFx5JlPvWOSv04KAfM8efWZJyp
aYbV1IFF7/XJaownGMU70bqJ9ENYYla4EZKUHeT/MPUdJhIN2tJb5JEppnoFEbvVc144LkVMuSYM
wPW9IMnIyBwDxfRcU9DrMUr5yQWlkp59GouZ0fmLISkatKON+N+csOebAfZTGC1jtrzc3+hrAOMb
Fc1FXljVSvkLqKY+D8pqcFfyKfgQq8+93ykOEsU1xPin6OUC0FIvXFpC4U2IrosLNDsqvQ63MJs5
bO/2eiO2WAHkSwf7Is2EfmKOSCRCzQT900H+gAF8x2krZMmmVAcXUzF6LPbp9pbQu4OYzzV4z6Bl
rs+0MNlf2+Fra+dA3cXS+wt79prv5YJTcbaXGasEb+gsM2o0kDA2iZMuiif2HMS32w9HYyFqX4Eq
mQ520usTfcTzdIsz1lHUO8hC2NlcvMwPPa/lZvVbduEDEWH2rezpFumekiHv7p9P7+fODyKld7LF
TZLDaNH94r7niwbO8mOKmeNQUED3cxTlb7GzxIsIhExz3fVJUNnW7jUn2WlxuLFyFPDkw1jitOyE
i+XKL5I7J3hT/MgrPlx1NF6HHMOCTvKrRoXUWtTRVo87/Zq7QOQcuiDPQ1cVf/6LLo3mbIgLq7F7
9Wp55/cYCvYA75i1cqTp/zmMAfDyXYZXOxekXwavP0+1C+J9YlHEmr9xQ8ZXWh2io2l7SqQctFmx
qo/PRO4aKP7gJL3l7PS0BCy/UL6JjRRcydswlD/tT9wVDm8XaQbCLlVXnm6+Clet+vyOEdYiOc0p
rwJBACTW15I3A3nQ+XmINKZs6yidpF80elxW8BdfdI3+25BJ9zQzf6A2hYgFcl1U0Q8EUUxv4DHJ
lzMzjP2fBqc+DM4SWUfpwwUTleQBUwYwk6XcLh+O3+Xbnw2/yMpdah+msbSjjW1WVnpWGVn3LZdE
QjRM11eBcZOEeCN6/RYZix1WuyqVjCQVQkfXVYyeamGrUq5sNzZdPV4i3gg/+Mf+oe9sQWicgITG
3lCJmJtPZO77DlfgcefH57yRC6IriZ9h6Pnv3LGtSKxKBMKpDUBGIdi88bKmWISVWDmdj46OXpa1
fZMBCL6Y7AN/MHh2xKuJRqTxbjQsDtj0HDIX2FyfmXtN2xs5OOE6tLVy9NZYRced2geUAx9mac3K
xCX2aDT/mEGvKoPtaVpXUyUuUzs+QZGHsQqmVN1zm5tlXT70Z7AKCBrhkc9V/d0azpBRSnOrJ84W
9+o6myxt5vH77rWlitsvte8H6M1HwrPGwLyU+5TgkLW09gcid0RGWqYaRg8OA0DOJ4JQluAw57wK
kTz+D2El1ULcE3P+e8icVFbM83hCpq2hD0fdW17i/4wqMAM5uX11/Hk9OyoZSRCW4FxNhGrvQh7p
+HbRAvLJATy99oGPosRdnOOvexkhkinBTvFq3jufj5V1MrWnySDnnCW8Nu2KAavyKksFG0fxCxbI
igZguVx4eJMrglzfRLsW700o6QYY2h/6c5oXM0AkQZqwZdrdFTIMXnV5d/J3/mF+HxQUsZ2HkbLK
TPoyttH2QiPjIeI7qSCWPjffFIT6Wrd0Q7Aid4CBGNDML2uwLe5Tra/qArzZGxbGplKLQ+sq81gP
Pqof83qkovemO56TBo6fxF/CZlGoNRRGMu33I1lnydnr06tL3OazTQoXAjIKRTCaVvbm+FKMRDqc
OFRCgNaqxozK1DrbqSdvuzjmIOKBWItuq4V39t5jY1We8RsmUQDhJ6Yb7JpKNpgo7RUym/QyJU68
seyfFQKmARsubY2AWQBKa86YeXkTcAIC6JV4talX3GYwkKkooCtZBrfrMVTv5ukp43hZWEx3TRql
E58QUZ7mJyTM8SFLZNV7cPGHjM22/o1833kESe2XdY+9pkpkokih5rr+HWV7Hn3ARZjLAIquXRfx
fL9mYuQFrri5cGxQt9iJlTiucV5hQvB5DvqlfdpbduBFIB77u/cdh03MXKD+SG/cPugjAOqtMOfz
P3jLwVIcJxmeQsdJUSNjNHML1YZ55uix09VAnunO8gnx+J4Db5T9AzN8Gl6yAxxg0ZV4ontMHtbv
2z5oOHUDnpJnQ7/yPoj4qpJMmnCP/b3BrHd4WbPrpjfN7bOyAjykhOHGb6qY2OCgQf7RtugmWjP+
nbbdfE3S+AVfAN0Qz9mEDXmfJyFOS3sj836OdxcuTCTdjii8vVK29eWJEWiDEQBrRiyLmOuXkkQ7
pXCHbaHZKQp5EaA1Lt2UoVQjnGnoCUMDYVchJcoYh7EHXSf/oiafCnoKqJdqXUQ6xA9by0ydKbHi
umTvObUIL/LGEgqJ3ADSLcW+iJab8hdX1dfoE76zy2IzCRNqKZ5sh+Y6P3OvylbLYn4YjZ7H5v2e
Qgm/Sd3R+Bw9srmumQGI9dHQp6fUJzQBA/OF4GzGZ2zJu6zcEzTW/NUgFSHb1ojuIU3CbG4Ha1Bk
sAwAbrxb//EERcE0+eehZnxslD/k+U66HZnUXWrqVSpfsB9qHtxUhO9bSu/vJUTKrZrnLOowRIhC
9WBkcWhArQ9Du+eNUREj786p9B1F1xp1viviopGVeupNo5zCLW6dceBx8+DygOuba1sP+nGVz0bH
7YsfuT1mBHM5QGV45nx9x2kwG71sx/MdeWXPw7LOOQenAzGb0m9fwDIFtkr1NZ5BvObQbxIdDp9V
JeTrPhOkZWq1uWRUBA/JMX0lSSYRzfR5gKrZ5D69D5U4PjEBGB/dEuPTxY9Gu87R1+hPqB7d/PnU
qAhTxd6kgK7xf26p1NxapPkSjEKIpznEJ9Q1+kx9nDtkFYD2J2Ppv0HVc+ui6xworgveatq1Hnf4
nbJOQfxPzW4ePhm3ppNF1jjFeCLyQgBFxCEw/KeHzMeZpVsUloV2dM48eUQoSv9Tp+7ERTjhMKjx
aZfF7cnB69podGEzDQZTWoO6JAfYF/Yje+o7QUj1Vn9XxjOCS4oJslFw9l2Ns+T3Cw2OFiqb1YqO
ydtgS0SfW69BviGKp/lFxbrG7KWrJkOFMN5MUy4EyNusuclJnzk6d2gtXO6xE+a717WfuycvGzm1
IbVYlBZK2KSbObBvrrFpj1BfKvTHgaA2Gin2L5OYVZYnjzlAQJI68jQS9EfTgu4/1ViLbjJKdAxM
pmApGaHcb+dhAcQAHH5T/Nbjw/SibvuqI1TG8WhQAdWcperScGjzoRvhUqHrBzUvxeqCqVsnhBx9
FNdS2yClX28domtmDLG330ujVNJ7Cgh/DK7Bma3s+MEr4NkLO0CHKvG4b+FWuVfzg9FtplmPMR7I
Y+E1tDAW02QDhrCR2V7ke1KaNwFm0mHNsO8MUQ8FelPjS6KM1o0mj4j1pTbVYfwBXRMiv3o4Wjgt
RDEEwP7zOC0DZ7NChhz6ofXKyiF8UrZo+arjDAoWJ1+M+Njc6ocq7HOLGq3bcn7NemCL45AItDyC
O0jkR8wy1dsgWyLaoMhtOmnF48FC7DA+cJPGeuoyG+inv2BLGfCpsZs519DEaSfDBDL8juqBeTFG
4i2ioJNpAmrBKPxCcFxo5n4IyKdR1ruou9tZXoB+Q2lmjS7WMPeE4VHCG3S5XfnylrckIKRPAwhN
YiNPnJ7+zcglLNyk45C9w14qNAJCwUMZUDlo6OJjQrgrYjAglblaV0vU3QLcxXZmZc3/Fr5pS4SO
2zv/N462VX+E2Kd/vtgZbtKKHHuTl5RnOs5AxA6Y3LP8Gk+bUrLEhHVyZ6DbHRVuc6X/HSnQWiih
/XYa4QvU0tRMhkZIeHNWqrgWoKRN9y3BwK3yefPghWURvSBNIEHc00CezeQHPgKThtIJSrEzxiym
n56w/o64NlrsEaJr1wSs3tcQaQ9EHWDKj+sMoHhe9khksBdN55c7tLZDdYoZniNheJdvP+mMfhVR
X1SanUw4NF2Y5hxp/Hrx4F3yW3z6TBc8e7GRbxY0JO0bPWs8LBi293Q/oWYbh7nneFJojPt5Oc2m
oZnWvtYmaC3VNI+kI9T400FyZy+niMJ29/mONj4vyarVozPiZBevxxSLGvpwlDm6RlHfQN3gvRBU
piUYUxiAlnQtUuSbtnU+ihph8pt1bCeQiYYWZvvd4H4Wq0x1zsAn51wvgbxVAMIdB8JANl4DaGo/
pcfgu17sgPBvfIqPMYF8P0ZChmPnU33VnZeJnLOfZQl7qUQLWPc6VoFfLBJuwsa2XbOf7oac/a+O
Es7TLlrdku+RvcgIp4Q1m8aSE7Kho/pf9Y4hA2H2j0U6UwXsfyuqJiIVnMTXnFWfyScilK10FJDo
5HN6u6XYXLVkc7Rbv4gQk3W3szfoIPW4I1Z+LMjtaU7gj/7EqkaIcVM4wVgKzGoaMGgO7khWlrbm
BVx++ObgPXmtN0Yw+gciEK2r78Zdcsvyyl5Nv0qBBltuWjJIddAamnkbXJY3x9/Sc/RzgPg0F/ix
jnP0X6/8mATDNrKAt4eunVV1nnwp508N4UkXbtYiU++Ve2jPIv4l/QrOv35c3b6V22DVCKxUjrUo
70EyJW2GcstqjR21ZzaAFt6XB73kHtpZ3H6HkPnDiZseCLTPiyA8A+p5h41FZtYKDkYSi5P1+sVX
LVJt7+4CZ54BxfTK98GnOfPuLDGF/ocI9dYkq6qh2w8keFGWj9IrhmQcDSaJ/A6jAQLKPStPimaR
ZmEzAzooq2kR4RpMAfeypJ2NZpKNwNodVSqhbLLNRhi/aKR7iMKwxjpYanslPxrs46mINO8HzfHt
zY/7PIjFWvym+uJ7MVWAWVA3qk+EEcQrGPJgmGP11KOPqXLP6rxqzfKgO9aQkcb6sxuEapds52UV
CFWUfTlu9nAqT7Tb/FHh+IxXYUuWRgaGuKptTp9LHb0BfMTVMLkEpdJD8NkhFlm5xE5VWG25xa1G
2tbL6Cc6oUjbFK6zo98LMNJ0oMKUCmVi9d+zlymaaHQi3sGhOXKgHmSL3niAqBhMN3JEI6NcjbmZ
niMD3qa50zyGcJwba9ikkwGfUDObry7wgZpsLDI6VHX1oQbwxevJ3LlQyrEGctwue5o05ziEZGK0
k7tGCtV8QxTFJvQCD8K1iQtDAUgKkwh1nonMgxdsZ70ahYydEoeNiL8qtWO97S2oxU0XBCqK6E7H
moAAVQIucP0W3xH0CxipKK/IqI3AJ8qhssUpfX8L8E5jVa8iDW/nTC6yR8P1+0VzEltekQYx07Bk
xFjfW0jTUSh5U3YmKMn2DI96g+lq88q+lOUpX6oeP4KePAG4VsC0gzd+OLgq3pCQCNWis1GmzUEQ
qKeQdWJLrxUKsqrqUkT8/TvaK1awnKUx0RhTWENKbTVes4QDufeNTQsI3DFv41ag2Yv22HYsPhgZ
uhj9//EP9XK9BGNcAW2c6iluOnR13huOE4+gDEX8uBE8WJIaidvgNS1HWi0rQ6/dP+JSonHhWfK+
6H3VPJddRxR/UtsNPDF/3H7w30eAQdIRh8Arb8PAdHmvizWwG/CzdHOImbPQat+KyrUeqpZc0YN3
57FDuICN2pJTq936fyXGWIszfNfmRj5mKgKTm/SGVeEuOEDv9ubROaoD+fS3OzZOIU1hP0afn4Xf
hPbeHyIu+zEyNSjyR5qlgiFFeBVy0r/kZZLyIXdCVbus8Ykl+gE6TLres3otWysOZTDxvSyo7dwh
raNJ8H4DgYpPyvj62KAlhcZAhF//pngvemsTTglKscomeOrlWgNHsd3JLSaZ6IRWG0e0Cb+B9Oc0
nlQWWI/CmBlv7zOVomGQyWRmast671p9oi1ZOHsnJ/aFW/M3PmPyfkHMkTHkQ79+Wz+gtQJMgfE1
9LsppgyoDqbvsh+sBL8dN4vTUDrMlRtvHf5fo5kiPZ5FGCn9YowK//w1fjLa0YtPxnJ8MsPek9lA
jsV6a8rRSrIy7SqcfPUUNl2uiownaQrcYyg8Wy2fjjfZPThOtwQ1tL/QDFVDaVXvoWzHwoXkbDUg
CVvj1Sj5BAAuV7kkHsxuu4SLyYpMq0ZvycIArAgWEHwJRVU1Kv7Q+P+zQrIq7gjYSzMtVm7tITie
pQdKEXwa8+2wFyU+HJfLqvlshM8BwruXSjLknYRrOtW2YmtvAq8+oS+6qpnwbcNVV1xu5kiCsPSm
QrM56Xb7MiL3HHyPVxvcEiGuUmqzXZBQ07HK5FuevL1r3FN5RwUnVt6zzp08HIRaxGq7l/9ZFxNy
Rqo0akLHjIcr7C7fskFYlfStCmSiuGo5tR5f981Dlpd24w6Uwarw8YXJa1W7GyMMPRJVUuBGt7+5
DMZto/2angTptx7bkymTywt7IWv5ztYoEDPdpA8EzTLkL9y9vEcd8l8x0n+vDWb2O3WDLG15H4bn
EIk2z8dnePkplfr+IfM+uGIVwBviT7nppoZUv37IghwWXg7lMadS7l1EFYKk2yvQVvC4SDv5AjXw
AxBElfE5lK0DIVTwW2jIKAggqWPIDgzKb9WRGJvkXlLHMgfvHSWvLEm9AlZg1Q8Q4w+aAS+4pnVa
bV6OgIav3XsWPM5JBAz01pGUGdj0n/922WhB2r66Smp8r+JBmjJxC6X89y+VMQ1RZACzjzvbdgf1
s/OmRbo3ga4uzfTikKWXLbcHwxhsQmwfVfKvEdtD1fej+6jgdex8QswkxfBEjVXwwGG5bwPQSEpG
MCV1TRtulYAnYhkDRqsueLOHYisWbsgET1YMsY0GOtubq5B6ZLnFV0tO+sgrAPtpv0XxmX9s5Uab
n3wBK2virZ7B64nuINGz1Cqgr/WZXBiTSnr1zvScW4TtrjDoPjnd6LR6Pl8lIAhzSri32ZSdZc5v
IpUYgr5W7/wKzMfO7kVe0NhE89Eno7jLn5I0uXqHvmjPhM9Joxjnl1zYLuKBqWZrSNyZkPIkrESz
GSZ/3+lorLx+1+VWCrG1gRFvcqm24s0SPX9c53LxhuCCXbNUPlwDpoR5ZWAiwsm0kVMPzUViPAqm
KBJsGbhSreV00nuiM1cxGDKCbIljxqWR0MC98x0GJo7Ciy+YFjaev5IMoN/n4N+FVE54wGufIjPR
UiIgsao7WipehsSB0VV5iHQzwn8AcZFaKDQAh09SE8wTlVwf665p3ANPRj4XaEbifMIKuUZ8TzGI
3wLMvHcBz2UuPALTTq7vWOmfVUHPBR/wMBgh5X0K3zYw9cQIZUbPI3RuX7Tcz9cxtf/7VBJiqYx1
WZjP6/Xxuru9j+zHC5rQAYrjH7aB3+FliXn9gy35A5ZQL10Y/P+nchzar7f2N+qGdBnyyQexRlko
vpR6xP4/aymEMksCjXBSsBhk+NLq/Dwu8dSOux4jhip5xukgp4M4JLJUNUeyfgoLLBEACz+vk+61
KHSOGLvN0USun3Wm9lJAmWKqEws+PU4T3csG/eyoJA3d79WYKM4OjXK8sE3ZXTjiIO6lCH3nD4w/
7NZrFHHpQQOZ9XT/nET6YTrshP/1ie5j3AfE+kHcvFyZDMPU57KaoeH7ulDFGjsy81d9JfZHduFj
GfaCP7vNs90DwYn+P6FBxUELDl0MmY9KAjbNMfVG6Dwk/Cghe2Iy1PGMSiPGpG7fTf36BgP5ZjQM
SK94WiQDdb8nNEW7DEL560EvvE2z2D6aEv2LT9rcGxKXJ/cQCDaqugIyCGANmCJ7ei/USm3WG+vk
5O5ggKHOaE+CVcyZQ7fkKQ1O82Gxh6Hz+ERNlDgY6+gsF2kCg2b0SjW24Kw5pkLo/ulRO+j0C+AN
VFi6tWjOF9pT46R6igqDrMB28W9b39VmX9REJ19pwqPvQSFQLFbFVD5pI/gV2qGNW51SHaEz+VdV
dWlvxU1YghexAr465P3GKuMtY7aDCLyZDqFybktSLyfq7sPaxL0VoQPuT8pdxgahYrTGbFzaq+ps
GCcTzkpOiMPybfOmuRu6KLegNUjeeZ9GDAEJYLjleH4cnuirbh+GUs2h9gn82DdiV5gwGiGh1lZI
yyN17QtVKDSxju2oWNlbinsUVpIz1PioeSGO3e/kdRwxFnZidpcKfeaHvBac5/1ZDYZf/4J4aHFQ
LKNd1HAVsrVDzOR2YETt4uJ9AIAAkOyfA5c1rdwpZYDQNPHuBsoNkWVWOlklXK1qap2PgVQoPE0a
FSYg/Pl5EjQq7oF1VtsKGSDehBSkMdAbIw+2ifNVOnxpLQXwtOHU89wRtzc5TzVkcKdMb4tdbn06
U4FmBurtjBGu0BPjMIuK+CN8SR2OgCiqv2d6HMKG9yCC2UC7JumMI19JSCey6ppstPJU0IQNCElJ
SpZ57nW0k7DPtoiQICx8QF7QfoZTPZnNs4fCqur0pM/rkbmxRyjX9RGqEd5vsDZYKVyxdy0jdI8g
U5mrBEwe2VT+/oQ4+Lgp3cHKoNYOlUQ+lJ5F15gzwj8QhMszu1ZRcXslYK31s/WJ8FVL+3xkJrct
YBNKTtR3euMxAks2Y5mAxKXq+x+1FyILaMj+Yv50eD+9nPIdJRE6yEoLj/LNYZpc27XbsAaVkjhm
CByCi9JZCVPckEx3/vi0JyxqSbM5sw0mNi8gBzs2eP01iDIRZPYRodEKpwiCT1X0kk3K21KeiQAR
KSsfx/eL/AraWcVcHz9G+xqe7+IHfA5uwNzl0xxdRbzU6VcVG5dR/lzkJRkEBDJqWdJkueikvDIP
X5o7XglhzOnz+VN3bg+MlnV/Bsg5YAzA1Flz/0h6QHf1jif1zIwanMhXhm28Z3obEGK4Qdvjp0gs
vZevQIOtYgpl7keqjY1eT+WWC4CMbN0A7xUD2TZTyhngRrNydZKvGsx5BhMa9au95s84QrY1/+7n
tvH8mP7+bBskVVjVklMPvY2F/Wwiv73ie3HIvKFD3scWuypzgJegYNS6nWrHsJIulWzj9yZd5u6r
PinjqV94ulxQOUj3fJHLh0KQ9vhtcNncCxbdF3zIesIVCB8uoOBodXVPGB+A25v2NseHDTgrX6dC
ZdmaM/2Fqp9SULDzARncYUFwaLjDrSHkVfyPeaP6Up+MM1OkIFi3eKUPsTNZxUMx72O0AUW9tdSx
Jac6CTHgNeSX1fEUrzTzVJxi68d4zZvY8U6Xalr0JVqV1L2Vwvv81yvW7adG59JaVdjZqZRmoHaQ
56l/+Bx7WX2d4V+q7MnN8/1AaMqWl1lvHNZscxDOhWx+Z5wz4Yp/RPKkB+et4vuXR8umGmPU+RoG
vbPlNYvMVv4CPDmJSUQct/yZbuhee9Q6iPVHr+Y1N4Boc8xCii00X/dpslXKZ628zLBHy7PFOKwZ
48dNHoOZ4vnAsX4pDZ1QPPygB06/GJGzR3AUTF0MVD01eyrMZ8rw3TJ4wTDYa1jMINUGDCh7obRN
5RYJHkPw+dgZcBAxCBzf6CkwL4Ij1Xz+SReTktjKzlvaf+0XUUi5Gz/ZaezeK/S2G1y+WI8c7UOg
zhLII8x/n6sfvGwC3d+Ce3D2Q9LUcx0tRZEo5WhL106a6a11saKhHotVRfBsSaQXV/LGw1oUeL2W
gknHog6E5pL6q/R4touu89MW+HEd90QH9nEnQ0MFQS9r6fCxJ1RqAAzjnxdtePlZ+IYaq+iPck4B
sL1yrVveoRYzH+NigvzCCD7vb3HXF8DOCDvKs/ioLRlBfMW0C4Ko4PwcexRVPmQ62sq8vzvGycvP
zaLH43+Tp6qnGOAHe743wA1vHYnQBYUVcAtkWAzqvaiQOk+CohNWqfqvRMyvv5fRTvFK4zY2Q8WA
bcDM17/4X+MIqk5+ik3yduYrJ5oAf9ZzAI7zSwG8emFdZjXXtJaTK/iHSv5RI9BWcuuKEeCC5Gx4
YkjO2sBpU8ARYrRjeYWx7V+Mx6FL2njSg38Lm132ciVgJcfl+E+t5lZfP+5mS36lRXRznRJ6og6q
dlIWZMi01c/ub7pdQ5AmsP5I1AxPiEItUgRovLKZFqu3Heej6UV87MQrsuVxaezyHMZlWjvNsiJq
RsPh0YH1WmbuZvoYIe8cbWDMaTWBBFFzPUQwLx4MkqmZzeOIOpVR03BN/9XdYf+C0R5gtfIf1w2e
OmJhM9D1+yn0lyrQWGEMcNKoBJ9UD16sN5Jcf2dPovs4dFGBjPnaq209L3/OE3C6Nge9NwCbMxl4
B+dklTvDFMek6kQLlLwlvdb9ofbeBz4bZQFA9rpEVUPk3tplh8ikoWpj7wI9+KqoMiAwmfaJJAan
qSWVRg0OWKZoymqSJ0CyvFuHeMD/Z7uo4h5DHT5LjJZIA/IU7UH3DOQKqSIoOd7AI2/NjyyUJHcu
i50U47wkNbjdzrD61xvFUx9jW5j7bRM5+L3f23nUC3VYIkwSOhGdio1w9Y6+TPcMOu8MGtFzi1Hs
GzEQWmqzTzEhQAD1dHOLmhMxAF0ipmElBv1fU61Oj55FlIce60qC1kZzAj+wU+Fa+R4ySFtJL9yi
uRAL/31q2vCsBpXG+D4YxORL/RGwuqf7HMemlFnP5euwGFTuvnmtcKAFANl0V3t2aUBipoWRpgSa
QooIxeKqOXvJzezefPxFkzyeyCz/l23QDktluGkbxiYuT+drpr3uYHnaWHk8nSNXYlnTy6ZXZqg+
g8bdY7u4f9qKwL1fNStpPofsnlA4/FhDX06uE8tu4Fgu7OsIZyBaPahKMpCCVUDcN+DFN9AltP2H
31nBC+7PDpnuY+cHtqXtVI4GysvLWI8otBXDuV6FJsxijatphe0j5YHKv9Wp9Jcw93c8108+ByVy
89li1kaeed52HdRE0U/qB9RNM9MnKvsRwxxFfPW6nzvqC/sh8QIBN/eshIM3FmJxtd6/8++Cp0Zi
cMFsgolJr8HM5wZ5TH+jsrUjCrc0MqoUiwWr2jmZgVeBlS9Vswj8F7tmoShnH1C7Z2OE6zJGbE4S
oTIY8H2+9pnNDZLEH6JLZ9wevqhNlotDEQhF1+I+zRyCV35LcMrJtPn1iXBxh9hCZ/ruciY0mscF
cw3Ye75e4cyJp9niIWBkJvoqGh3+CSgeIZnYCi9daODeBvzVJkfPsiYNW6nAUCz5AzExEqkGekVo
Pc/3HIimgIbPJ3JZHe5DYUmr0OAxN6ulqOr6uL+0BckRw5jv00wK8ONuIeHQWw/ejuiaKBnuiLM8
EncNw/Ibij71R1oXdCmVpUJ4KnrC5LFIgML0+f2fTJRSEOfOXVOcq2Rt1DJK83fG6cOzw/q6ZAI2
s9j/sm8mdSMaV/Dg7/wfs+m4jYmmnHkbDhkijI1wTtZk7zlD0L4hID3JurGxdKbkLwKYZ7sgCs8j
3C8y5TRXH7WsIstU5Jk+JhhKUrwJtRVF+XEumtitbP2cb+zJ4veA5pLS2/duEPDjTzA/Z1dF3NPI
NwMpe7kBBkM0Z2sWRxJssXreMtKiN4PC+fyaP9oL/d3VbXejgD/ioxYQig8Znjk/z+037IfMcoT5
ygk6t4avuDksSp3JWVRnCXQQ7hwQrWqOMhGJkztqbyIdxD84Vha570JklrfJ2dYm5iv4nHoAkm+3
ronsP3Rf6gEXI+JodHO0mFO802HsLUtsTHcZeuGJhnXEI9hPQxp5IJCYAhtlnyS24UbdWwy2ADoh
q3yYKLE0BXxBAlYVHSFNJGnJ2sz9tczj+MFVSul+Y/TFtcXTfbB4kYdDj7HZLvAfXkU1HmktGXbq
XPu7j9HZGZg9/0S8amf6aPGoKkRL/Ihs2uqvzWHvbI2ONUaG8/jw8h/q63CFjGIGANW6BGDRLWpy
u+dTKmYQdaXJIGpTp9v2cy3YgGyURocST5Ms951wf9JX+PZtO+mq7ERNDwLQB8ZvzyUh4PByKjjV
mHMGBMfdoEFxMrPBcSbnDh0DnEPp/xSwjfHhiUYZmkkRmSIMSoFK41yUEGVcNVmSLKEnDVM9Sl0U
X45WMu/Q0UFkj7dh0k/4FOzFJQQ6UdiD+htVk75AfLNCfV1pl0XfOUTKo8l5ONi4nO2bifz8ahoA
W9twlVOsEmtxzjuWzrKBwkhuYgT3U5Xr/OGJolm5M5I9aVjSIwSlcB0GkIl4Fs7aJr0ljRZSdsYy
rtKEtDbv743zcd47YtNRys6fpCbG7oqU2vFoTSaKczYbx7AttmEjh4BUT/cK2YKAwWrUzA0jt7e5
uXuu7k6TFpggNzFivY28qdLmFMmAG8BHo3JZ8D40pnNKF0wl/ByYKg1uLqmpKW8z3LTEuxbxXwTW
xX8g0ti6g7d46kYBYuGX3xSiNpX/NSFjFoWSh1S2HrYY4F6fDGhvSyVeEawvg1vEHB6UXkXZij1u
JPHkF95HJoNfNGWvtOpK0ag9EG2+WquCe3wSR89ITa2V9nESGgPcZSGloeABoLyrxcIoAJVj7ZUo
/TM22+TX1//uUGRItbgAwCAKd7CcIxVqst9Nqcd31P1fVhwts4J46DpRCR+8RPze5rUJ6BNT6vyj
C54jbWh/7P9I9mIpg0MROcB7+D8JyuWxHJWxsu161MpM0rohWwD2CZBshnjDddvaSpO84kN5BxOz
Zd6efO1X6554HFnfm2O+M8h5OR4O+V+Xn0iSNcabuVcFIR74qRcKwvvQ9LnCR6ffKH5MW0VVODuO
DwC8cmc/Cceal/vE37rW/ukEifSJqIygI4hrTauzghUIceR1ETWKmxzQo2Rw/vneHzpQh7fdHqsm
s4e05zwCnTv8Wc76CIOWPis0f2hV+XAqqCQIQ17TcDLIJN7NskfxkX/05Zqtu7SN7MV9CU20Ug2M
UB8T6X3SB8ovhNeFDFLo8JmCkHLTq39x6MhLcs3g5Mie7iCYcheTd/3iVnC8x6L6we9Yyef4ZcXs
0K/ElEm1x9yCk2wvMVuBjz2pqEMInIBK607oUb/axqKJcsTRdqBau3hu1vG0CdUrZd3ZWFVuUacx
s/8l9e2yNk449m5LbW9Yy1J45I9iuhvPF4BXxQUd7sVYEsYcVttH3/+qnIYX8Iu66tpZPEvs5Gbu
9buuXR4DOO9QGUJk0NMi+qHsxPZFWiXUy/pIuFk4XlUQgBxR8j/z9HxIrHdgrDQ8x4EHZc8O11DD
rjIgoDnsSvfXtbXdtGa32sJwAsaXqwr/PKQBRfDDKcxSmjieOVua3COtDHTs1WI0/pkw27GYW4GI
AkP/72BhEhHHRADg3eq7sgpM4aP1cbIl8Kug4buBpPP8iQVO6GypNkLgCjoTg8trgKDN8ylDrxEt
liQRwAH7VaQabvbdRR4/aFRDOCjJKX3w5EB8yNDL0INfREEF4ogINvaeN7UFi28hL0QQPUjvtUbK
XmUpHpP1UhLVjFhK241zbq5UAh9vEPtNXMCnjLo4zCDYmGCcdgeApsZP/vrg5xZlBgZ+pJyHc2s1
KMCmKY9ilTPwba1dUR4sFKsvZTXgAS7ThIUUSS49Yq95m6UJy+1QvA1ukqzRLV2kQstTT5mcXklt
Y8v/nMzT/pCCl59ItMtOwGhqPXUwvX/F1WxJxEWN+f9BnpB52PS0//IysyEN4S9/LSTIpzGy+D/E
Yb9q+sAwcQg6pu5Hok3h0uXjAvZH/SbUSmG1iwzdytQikdpwH05YpKE+bj8UQV5rxCwGqrkXCDd9
2Dsf59dRzrH7jYgvmsRYkZZxrs5CskzrRV1gtGXykYTV8dDuAPkRLl/CQS5XjPf7POuEDJs5YXU2
0nA6mTwPD17JqEJnxSnOoYnnG51dqsfvZ9m7cyI6LPEctLwhtKH3sojB7bOmAHlWjKUq7pLDoeCT
yAAXRagrF0ubHghsJczqoR+lggPkDlP9YVR6Vu6zxl7lzLqer1ACYdZJltUgnXLwEHYlgCXrwpWy
/e4/LWP68LNMMVuj3FXMjVakvcXfW59jGVEG5Sdu0dxTMj3NG8A8DOaAgRrzukb4drvbMt1Zh9oh
Lt8l472jvF79H+QUjvmH/zQIYg9Y17ehXJR7sdw6QdxljgV1fN1BTtpDzS/8y08EYHH1rNm7v4mc
PetM+Ka4Wg80/FrdZ6XFIj0lIVmfVG5mwhQ9COOwNpu8CZCmLhh8qZp0kiL7vs2IHtntlFsFEF0B
52P009WO7EiR93vAH5cOHcqeD5yYAw1HVulea4uA8tmKGrSL2NkYp/qeO5bL4sIptItna6mkbDhR
4cX3Lb8wt8otWq3EXjgoLKlwCBl9iA63Du9Gj4xlQu0Ls+ifOTRdnnXDyFI6agLO8Fv/+bPBhNhv
DkIrOLJMs0qJzDJDweJEAXdz4RgehXQzb1bF5VW19zLpUkqINRIOwkpkcVTQQhkqpN20Fwehmgrm
WV+0A5HWPJn6srmXIRWbfKbChK1uJjlMKZ05XRga9N/OAVsHSMPqjLuWKe/DOz7lC8R5GwThu7xs
bCaVtCjQ/VC2D9dCkRMIjjZchm56SnRg+9cqE2NF9qTFXBLZqnPZTKDgLc2MxSxerqb8Hr4KkSRV
XV4EspyIby8PIT+sKseUj41cUkrq7ojCI+mZsh/fJ8gwuLA2eXkmyhZNEFWegcHx1th+KNu8fSid
1gf9QVGnKTNCKipqYlkZV+TBU/xTlGRuPmcYBOPP3mpbzXhiEyM92Uft5nN8BZHQ2NKzNWftJmY/
fpiI/XxcVMgqndIKB14CrUyl7ic4zwAwJ508fjsYMnABSf1HEhJscoh+3QrVbE4faRRQHJyDWJKU
SyAEJeHNFEHQPndA5aR0Mf5Vgg0w0U7S03pBqOPC5G9T7p7/TZKia1F+vOh7YDX31nVKIYMZ3qGR
VkFF5K0ICuUGA2kwBhF7LH4l0YmIvXsKjWhRIyCnZNGxA6jHpqXFb6DUBOU98atMUFALecCGdKTN
XVRJlIHkUi6wZSdJJfwSU9VmWhKGgfl3fOXZCH8BujzneicqDraUeWPz+ZfraY+Jy5EKnNlCPS8j
gND+JD9kXxinIRLNhDMXJ66Oux/cTAAPHO1RkQ9BqfThz8wfCBgbC813Fj4up3S5A0U4tV6qdSbJ
ZmVdySymhjiW3qtPHChCQvSJBokl5BgDafZDe3G0+bG+M9divX1rC1WflGbvXMvHWNmh/k9HXgph
jIOAB1A6vyxeLJrrwzBvUsKEpKYUjgzDF2mdKGFm6AX1d/xJM81OoWUySVp+mRBOGg5C7wvx9bHb
FW5C8BPRuoQ0e6TVBKsfvgcll5jqopByuIJqfiDv2RhwwfJhJQdt/cro8QhrNTB7OUdwFV6bo/50
sBwcuV+S1YNiEf9jMA+aj+3nlHyITG2yPibE8mYPH2vjgtXb97FWfRngycKVH5oDW2X299smn4aT
FTXE4cdf8Qtic0ttd/H+1dAb/FzGleZgu6wwvJfhXck8e282gV4L6VxKCqmix7isDehOEEveuLVG
vyN7qmGZeMHTfgy1a1A7hwlk/G4HHECrn+AglhGQpSdsJUrmhj7u3wIi+00Dtw5hT2Geq41BaoGi
/LwnGWtEUjCdsaUF+kKDd2pcTGG64WoRcXfWbuI5xNijnP5UQ63VxjqXo1minkVYo+NfnnBzeW20
DiwMK7Ouzyyz7CzVIJ8FIaAb7QLFATPEdqQBsYP3fo4AMc9yS9jrl3vhbXaG689+znLqSF4RPC34
3T/T98vKwCogoVx1IrTOMODvS8RXYTsZPn4jcGb3LVaxrG2Q4PXA3d5U2qJ7v6OBfNEBWETb/h2+
cDfkHf/Is2ounhOCW5Dyl34H6PeIuhmKDrM1Bl6YRCu1mJTeC4XhOwXpiKUgxbJ4qbii684veegz
f1E8MuWAfoXzo/+I0ksg8KSEkq3RR6teC8/+3cewn2qKwq+mHzvAgoiKPNvGlrsZWNEMj9wkeWBK
ZYjcxyzdh92tv7exTsS+RS2HDclXKYiAw+07xwr6qYRHkodQw2M2BOsW54NDdE7VMH8XKBSVxV2z
iWEFTIFlT3eBPyFn1XGwXcWEUdEwgM/CD9jN78XYqP63kzdcpwFAZAcvQ4RW4XqQreaJioCQyP7/
Bw4/saVjkndPxhNzg5cdeTPnRsduJtxaTz4/riYP/R79voPqNLL+WQF+ZnYewX7gg6a1MFbLnVXG
25jaq7H6ucaEK/SNRAxO2HXJzZ1VdkRxRGMxQoWjneIhRmIsfaXKrpbEAPKNBm11QblNyOKXj0PE
hpjA2+3aNCandoCQHfjwf0l5+svxt+doLO+US4bCp53PCo3qybawvQXhzhMs6rnvLVeC4Wg1/RYD
/Qpl3zQg+iehCim0/2PLAeeVn1PqrywElLY+ZPgYjhITD5CupHieOGSpJtsRtauOtB+fDb7vMzru
EDkL9Ie+IW5k7vNJCpIx73KgFfNHLe8oanRAGZ0FlVAtFN+CRWRtK3YH0q0vG9Ukr6kEzxYJIAAq
Z0we26PV45RVb9x8o7R/raR9Iex2X3RPhS3cXwbBcgUAUvI29y/CO2S6Teynyds1dQTR+btfr1hx
45ooztw+0n8H22h9dqujh0KfnnsINgtcwWfH3agApdMtJZC2LNTto3rqP3Qi662sB009hYddat5M
jxTqo1CxjKau0uQ3tkRp5L9rPl7czVBXjE/vLc9egddTLSt6FZMYv0PtEFhaC7q/nPdjAqdiu7Fl
rlH3e711KkMI7BcKFnNVkP4YOWaGNH4pRDjal4ohiretnYgyKChfCDb06jHY6YCJBrXinZGJkrBj
TL5Wj4EkNo5674miRjk5+Vn6TcLtFMXw5qYeb3UwZsTXnN/TnUUrPGP0lemmK7IwONdg0edOIq46
vmKPoQlI4bH4GSjGJgeaxT4OztM0vI+ajOJy9saPgkr6tDjK+I5cHx0MOt2ISdKrTrtJ1vaiJwuw
qxwXPTwTutAK8uH80W+96Ate0tCCvoGLIrPvwJ2Ir3oafUzj1ms0vA7BUb9vCEI3DVPZHMmLX/9C
mVkpFF9glZFa6l50yPCT+utwHilhZViD37vEXFQH5F0PoqDJcTWUgqC6Irs4AV2okRrVnpdQic7J
lOCZySRdKbCG7itP0TzEYafJZYBC3sB4CC0+E4MrhGfaNNeFGdKB6HSC25mkV9jVP5cx0Z9mczN+
WQkm914WAFxBT/X7CBTtr2p/9+TzcOee1moBciNu5GSyAHsw9jsf0mDQ2djew73/EGj3FjBPDLmJ
ENr5JFyNqq8+7Nm5qrWz37eS60Fi9CRDHzYPTlnJu6w8lPN6+RkB0TL6XqU7gVCy5OMxlFJK/bg0
M3bmM2FwWbZ9Kfe1ReAS5ZjvbElu+trED4IqvoHlzi/u6uDL7arD0zpHyPewpCzyhdWVGc4dFfyl
qgRy7CPGx3HpCGx4iUMp53bauNvfPkU9E57f8gQnFHMxu0lyNASiQeKb+R/iwkFlkvSXeyZTY9b0
AVjNPljZftbQLWuzpr3WBsa9+FRT0gVbowQOxc52To04mOp6P60ZLJMxjOSKx+G4iNHmsRbhyThY
ikOpfmC1j4GB1rX54ayoFk78pW3wnJS7iKyPf8ANGTQqFvFPfagXm0yx+55qLIdkNxuKnNmCWnRB
D0mZUP2IhfbiNJqhNFRRr2FwbG3oHZ2r+mZBUGzfQBv3jCyLX6SZgfAIlkQDDwIt9vfRzkSDJd4/
fDAIOoBYm53DTvQ2+gcf7GdT1vbBlq5pdrKbp+L0biWS8VBeSwtygi4RuoTZ03Q21LR+o4E0bjXm
Zcv+fgEmMaxb4j+3LAst5movAsjqs1u6+aGMypPDd9ryLf7aQpXK8JOPP+Xi2ZAVPfQxrPPqBb2K
QhUoRVzgLJWn9J+oh9eYBD9M1ihuf1YevDbe4FaxikerJXe+CUbekgOpXQkOXClHopEEVq+d/UGi
pjNsVF8DwcS0W81SHdhXD4dADrHkBbJJvf83mMnVX91+6N95TOwkfQ6amsQ05XWdFSqtCbZlw+rz
a0AJLLVZeY8RVj0ndovvsj6dZOeV2CzOH/y0nRc9GJWDmSNMPYI0qj0SDJGKp+u8ua4jFnOFf4yd
Q02Ljl4RlIDFrU8VZrYGJFXdkV20yVw8lw7h+r24TtP35ICH+E3ls5v/sUXFzao799MLyPSKfo9r
k8OIb1m3IQPJ0sR7AFGJeAMf+tlLCKogPMt9mPd9qCV2io7pdETazc6e873A6pEI386MzrD5HK+t
RQktfmaSeqeMxnE89OMMJKq9WwC29Iy4hkqDmqyMAcAPgf9R0JsT9R35JhGAJpjH/PYhLP7tYufZ
YCWt2Br2wYcYY8k7uXSb0K6zI5Ojx0IUG79NoPxeV5fliT8/SHLau2Kg44hmAq/lIWDjyKK+Em9y
sjigxcAO0mWtqDirAfkO4OnlSb+BLRbfaSxTzuyk9usg5rqHllJaQR0ykTTRsPWDAcBYgKwyUY/+
U4neD15eqIQlPVFKih2rQDJdksCkVnWAq9usyuQ9jzfswU3OPNU4ZG2XWe2BohqN3k1qXLaqczKp
dXTYuBlkgjr8JL06/8tXZT4IhrygLogR9LSpWbDhrQlYGoFW27QWh5DSmOLJotNmlFHPFKT37H6r
3ghGWs1n/CAqAMUX+EBcSMm5p+KJBpwIo/0USo2ytYVSEiJ55XTnCsygy2/UNgTX8ndMVxh19JLG
6iwCiAYdx4Wc/M6pNrGDVI4x2/b7ktNaDoBUIxmc76Q3ucJE2hr8Qy1EFF8AsuamoqWWZ+gqeK92
YJ4j1J+0eSfaqnfNwi78HkXsni9Engz2XutM7RKxkx3nhJpZafGTP/0nd1P248u0Ik/D16tzGuom
40IanzzEUmhNoaIw+RHITZT1OVOZX6P7eTPNGe7eV7wTfCgGRArc6jAeQ/5g3zwEKBCpaLcnPD1n
ImidQ34enTbV/ltt4YobtB0sKXn4YN/uXjaUAyj8/UXcsf/p3CaqaQKq/Q5DM8jWRuMcu7n6X2b1
dF9M1+1S2K+CTEuUsLTzBXZAwme0EhsNt04SA3EY9TKYk3C2mNFDJrH2IJ6BEPpDtfEl2wfriN6a
wpvF5ih5ijxUvOSm0mvCQ4fVilA325OcQPFFBEausMelgnSOPhxuMQGm5awSaItu5kCj0jX8G1xx
ccovXo6oE/QpsJWvwkbNUuPS5oqmK6gMoSF0prDUXdrAjefxMyEASxlnLNFWnOUJS81SnxWQ6DMo
ecHIMVurFpFXXQWc5H5/zRdbNxp0xpNQFTEvZRRquLE+1yoxi6CNoqQG+hRCPoP8PRt7Jfhp7q9R
eAXq4jX/vloj0h9J2gVo5hKnua0AnZBJT+cL511zB/kqnbPHuWrWKPVM0DgXJgb6c4QH17KfgyXm
yerEQ9uBS/hBmGGZQz4yKP+q+t79JmpUlfhgg/9bntT+UHea9uyDRlJ25VaZbggTEjSaapethJaE
zFwtLHogzVMzJ+tHNxfdWR14X2WuIkWWUYpnIUFa0YS9TCgUPP7pAPQC5cNiZsPrZciQC0L0DJ/P
tVaK4i+LqBBxAT7q19wLTbYVCE5GTmPQGAmb3aCDSHGOnrGLL5Ya3+teJs0FNfTJGEIuZOCwsO5o
fQ5Yne3uOibmeWLyTk/9/8XT4HlN3a5WqeHYw5JhbCnje1k31nXlNKCsLXhGyNHOaAUDJ+AqBVno
9/imJw9gqGSMvHgbr7cvMB2diYKbIfWIC1SPDdK1Tf7EKpXEU8Kdxr0HcT5wOr8nB2iOlaJXuEUr
LGh3VJ/R+wDxTDAu9MOCObP2bNByNF6blLGaHrlbCU8Ykw5kMCQjipt07Vq0khD/2bYlKZWx8GAR
PqMiJMPUbbQdTXoCzw7ORRWmTKJtM8NiqvY39guQJq8IAj3a8k20R5AZKqm/9/OixsK3i6y0KhDz
tG66qIcGWCBYhFZxgfBpOqYkffyGjm+Urr5HaQvDjRkF3G0LiIPE+YE838OES70BQvBDbYYkPVvy
q/13o3Vn5Tjp4tI8OgFm7Az79yPYXcqomq7vlldO/gMYcu9s6aygaXSdEWCODSYSX0ZQWPyk4kOv
VfoNTZLlgcGVb+DTKclQ26MRGqBDvzvL/q0nkhB5KW07K8i6N3XlPLNX6U7lKnYnuPNBPg2ggBBZ
8cqz0SCvdXHQOtEHTtQEyWpqDhNkmjlAJ1YqSNXSIZEr+P0hqzbOvgc6sHFC64RlFKt+ORRfMp79
7q/kXyE8t09YkUvpat9CnemVhLzM0eQdQ5CfrySNe5O3vILwehEVhEW7ue89dWUbzZKSujmjs2pM
78MqIm4Rb/Cw6lWSpYusjDz9c4jfyoIqk/fks08pyilRMxqQEo6XpePDyWGPQzvOAGa3p2GrBSP9
+6BlBxOO48YSpg89gGAHmnuXZtJ/zBqHPtXY4w6W9pjZsWrojJyvZ2P04tmXfz7hvDlTOZPW+yWq
hSUl4tq70KdbQxSg8i8FJHSEmLOEvWArOO6v6ur9D3F18R4DppfXrbKbncOGJXdPWfnOqYX5ZjVu
lUoJiQReNrVzI5i5jku6Bq+fo3tyg3eb9DS/XuxcmaYKSo+PK8EtdITsX4RgW4kajT7Ec1/gaeup
MihIJIYmQBYVpuzh0It65DVtao8HRCjYTOGyN0gOIYzgQddUYEEodJ60Gs3k72tZfTskjc4Eg78G
MbULhKRLqEJMdCRnCj5lG/24szR+zgV+CB05Zju4ANs9L3Qtt3quJr7u0a/0GXNZQKP+Nc0ynq1u
K87TFUEHhkqXECIGqUyQrNFxuZeudQpMYuQSXYx+QB4gYTZKhlL8FY2eL+oFRh+xkLuY5brk5Mmx
SwgXQRC9o2HlIu2T+uE1rhuhETZ+AT3VgJdK7+guMtbH8VQoLteQyX0UVYzZxfen072TTLrbOqvI
31Y/HPo/v2lRpVQxzmw+hdvXg1RS/VqwyCWN2aiG5DkMsaEgW7l+TZVEcVKo02oA1lv5MIJri1Vd
aMS02yrcj0ckKpffEVg2Sv/f/5BHizzgLlMLbf1a4X6E7piaO/edCQuBZpKh+48JQdc9mTapoMZi
CSlvaTnGkDGh4qDPY89yhYbQiwqz+W6SfwXfJ9R6ui6oBTeOH9WMR2XRIHHG5xiCoHY1gusT2WqW
Y6lC0K7m4VR5D4u0aYgvrCbpePgqXpVZNUqhCME2XYzIHzc1ggzwfuZyBHOUjd2vcNN1V9F6N7XU
1H87DJxkdEOwTf0qI5EEINERYY0Q5kv2kDvH3YgtM4fUrU06jVlH/QGTFS6cmY41YY3eK/poij0h
cPOCBcZq4qbXgv+vwGsulI357OvoTIe30FdBbDBO80Xvr6nrhdRqJFFnifX8ROXzfUMmIz4Zq/FU
pRS2/phwYYjWkCOo9FbmltwvOVkW0+62rblLUttXbmsmeiLi6cu4AIHqD8/3Xao0AYa3/VrFdnG/
titJRIDiyln620c7ZML8LvaXb/n5RA2Yg28uycodFIywZhHv0Vy2fCyHud1jmQ7EBwaMFq25q4E4
KcUY66oj7w/4paC4IAPnIF1swCTYttcIVR+lDA3o9Nx3JaYsy+D2cNds94rd0dcaPF/QCDqUc/OL
+jJgqk8lRTkuE2DFq3U5ZXvxss8z42i3yyoo7b7WMjv7y7S1Zw+DfXkq1vQFS2H/rzFRy3EMBVVX
gvuvOqsccWHKs7gzORFgcI7DL7LvyTRYufZ/YTgXruGaBInZF/9ghoJrXTCY2DKCODXt62sIhvxk
X1TPdDgoiOmzIJlsAaEzXJbknZyh3A2ee/HWmaHkXoDhacJuprM6EeIAH0mlgipHgk+qoNV1qslH
l1N4wN9A6GwevgXiC3hmH2aob2iPgyfs7JCRrv5dYCfllCbqUaWnpNa3tKZCE1igawNET5aMIl+u
0suloBWdRc8zwrS2bXz8xCiiSnBwO8TelTxl3M57fJdy+yvnUfwKeOjhLonTI49p4jS4JpCCWXnV
sFSfzw+B6VtfvpGfgo3NUFbqjPci9z5mO8E4SEUyIVbnMugcXJBk6e9qC3xMxYetaSthbcd3oHX6
YxFnhjG/7pAHS/VhGPHlUZOL15A+kYRi6ut+pS4e4O11fW0nBBsKoJsNzSsTmVtanmEjXaqMMlxT
i9n/ZH3vqIkdGOBqGP9s54yKluwKeeiqAOuqy7H3VzZ6fOnFykyR4fu4fEC7g6NIRIVgmkQ9/lZU
dqcmkWQimGcL1Z8/RklaigII1UV+jLn9SBbtoUcWfyYryqoQzEn6mU/J0ZHaYPQ1MId+cS0qFSX8
xvwlLRkmgmb4lV53vqodBy7A/9PM9CTYP41NlQnWwiNBZpXbdjNRkaLPI6ZKN5iVlQmhg88WgCfy
x192Dzo5UYZGfo+rH0QAbG7agI3EYuKfNBEJ2xgFVtWI7lLXcCXNkjO05BhRKAc4C7gpbGlDBHKy
g2hcL2FJrtOTd6x88kSSYe25Np1LmmGws98qY94qryt+vp50sq0J8So1v3RAUgJVclxIsYe0NmRD
v7V3FJEDllc3oggfrso8zucPPEv5HznqNPgcK+ZrE7OVpNYNhtkLjFqwax33lo4jnA4Ga2SgSRwF
NO9HmPebdIt5GhVpNbrqIrFSJspwwxjVtP45AeiJmHkzjAZp+p0B/nCfV7hL5hvv5uv3JssHeu8g
UgYz+FDpKTzEwOpH57BNSW/WtDpTjY8cQgOTOxhWg94EyD3clmoEKaDeusB2Kn7I98K5xOTOMV3t
j9eZYMlgD1ldtM+11Lfr5Fe25sNZVEs2DP943cIWgy66DyhPR/jjccCk1Ovml+zHkzfDjHu7S2nk
cManArRUbHudydMc0UaDtek5uO8MW8eR3G1jw9XFGpV3HZtChEmVOasthRUxXH3vWMyoWkk5a2rZ
YSOqgiIm1KydhBhtZ0NPh7YPaNGCi7l6huqjcvltXzN5ejbRGk8rkNGncaALoSXGlAty92oQ9bNA
+OwhwB+6ao0YQYVy8teB29RtbfvOYLPri4Gs61/88xp6SUouhxzgg8wGqyecaUu9eZiHD1Ypn3vD
8q3p2laG1e7IlU0K4JMnzDUyAOwjsk7rPJh8nJZfA2aP5hTdbDorf4BV4z8Mt9veCZaXzBB2ulUS
Hut0LvEdq8zMGPKWxRmNNM9IY79voMTOiVnAtmRws75wIXmQbMsR3G6Q3DtpL2+Yxg8zD9azpxpt
MOEVXllhTYWSpKX+/qaolQ2UwWDWdgB8p1vTEbTvS3qzfKPf64SRh7NL2uUIpolSATxmWiLWhwXc
Ni+TVxknQbM9OaxCuAFUOvsVudfvC/ocPbS573WTCi8/+r7uBwA04AdYT6YSygvkyWuFg4ADqDl1
LjX1hXP9fGgMkwa7w/OnI4KhzbEpn7/1UsUP6EZAVHz+50Sq3etMKxznPUeV4o+Stn8ik2pLMLBm
JFSJrHLYdskr/N/BiyycKEf+T89M18SefWwBSd+9BdNVkdZf+FWLfKomeMTsUfUfztAhtQoc2IOH
uFF0z9ZRxwjyMtlnwFyq5qq8LJYx4vw3C4TPx89PWtAmmUSnpeyVYr3P53Mz9r4FP0BR4ThvlT0v
/d5ve91YcRFLWw4CpF3YKpJCxoGyVT40GowK2+A6uMPEIDCupYXywWq0D5l7iYaN79tZSxueU5Af
nbHKvXO5ZrLc8EEtoQsxkm035DVT7V2SPvqLsCnp53nocfXWsOiR55u+8e9Oho5waMljT4ZqQH4X
JhqadJJk8GX2vQLffx8H/Rw7AjhNlzxpyOlstiVye/mqGHdGJqONydpMLd3CtTw5bgiLSKOBVhjL
Zlc8i4X35HIy8ZeMWxKH2HdReJnBONAfI3uTc1EhEGhRmAKnrTChTflrlAQK/vcDHS8ze/s5czX1
Zy+nahJtYkX3f0wE5q6xXN9Pmrl52BDHQ81IZSdlsQ7Z9sQewVifl8O2g6zvsLP06Myed08mnaaf
hZ/3HB+5+HWuFWEVBLADZwcF+dRp6PeabDMy4UEJVtySw955hmNEGKar4kfCfUJG/C4OFQcbZ4mi
L/7i5P0aEVyUJncI8QFSLRA4QZ1ENqoJXlN4p1mdOJl7RtAMbXs6xIvwNHXUUUJcWLkhan4fmxiZ
/8TvORhnh2QNAg73178A4fo75eHKPEr5BFS8VyH8qGl742qYwxkgx1hQzhQUJ2sVlBEs7FMQDFxm
JOuDsQLMqotCuD6cMUIUlOZe+tNDW6SkuEZFr3fFwCMfTZe7ofhg+kDRKUVcJP7y5GTmsY5p1ev9
T7w0HGfabRRxzmWUMEYdQQHbxavoGgaFlaztlKM7v5XxPIGGNUAGWfk4ctI+OASbfYVmV1qNqL8q
TbQqyAQ9LgsePrpnIl3Q4JxrEQnAvzORear9kxR9pGih7J9Y5J1xkN+QWEfDqmX1hL/Ptq212cqd
XmMgg5gnrA/fQXvBFwpwhk2Omf6D9Aa46YXiO1D6r13/yJeLKfQs0IAYwJs3XdDG2N9nS032gLnF
h0DIWR4z5PpgC+RWw/+Fj7xHXGFeJRyvh1YdrKVKANro9wYt5V8/oM/cxh6i0PzEphDaEOUcqKCx
lOa6zQ5JtgX/xjI78d2Rk6gegfqwT7e79pMKXw9NFOhZS0h8lrrPN2D4HjTn+c2Mhoi3tnoYaVPX
UiIc97vKRBk2l48rg+40ydtB+bWpGOfnn5Ic2tEviMUHpHIsw9vYaINWvCucTs7GJhbMFtXNotCg
YMX51u8brMBlDeVq8DOVRK95vBeTnTTHyuduCtu2xTpwBySL6nXAg2eYh/rQPwpXNDeb3lXPrDt8
3nmU+TICRYkrDnTEFLzlJR1aOKxdTELWsH5R4294kj0uTfdGSv6c15+pF6LmdvIukU+W9PWVjdn/
HjtVkbiWvHDDXuRcgkZRLuKOCVtXKBSvysDFOygAZZEk87B7eEy+hif8UFB3jVfTsGbKM/ASEMqy
ORIpuUgIf6ymRG3qKQa8ypM7SuHqsh2S9u581Ntq5mlew+RVoo6GLysLJ6HrwEKJ6Oyk7rhBFR8Z
ptriTyADFTNAis9iQ8vHNzV9otXSl2KwYfGgP1R/gfc9+zqJjGrI/L+hbTRgsIISdy4juOsnNwdQ
RtmAu/wrIB8KMRI0SeDaTYXfL1QoyXSPVtsVl60SEXKV8td0gJxnyzEi+WvtOfMfiRijI1jhuT5M
y/NHjoyY5lGmKOU3vy01M+hu+C02L8QoQ8fBoVSfE1/XeJg4ZRdSY9CaIiQsufIsRHn4pjEXSecx
cQ41svtjwgTBXjsJp+zqdhb5NaTF0fVZQkhaPqq1VNc6s6zJS/kmbmitgzXplr9RsVtKTDECwgXM
pnxZCAki7ACCJlQbWF2tKTzVlgdF3wwgKKFHp21hJql3dJJ1X2/uOmUINsGX9k57A/gWZ/G/V1Q9
k1b1ohY2PgAzSIdzG5kwankwYWNxdqsLpny6Nq9I3Rqk+ytzMPOoMn7893zNsghC6K7ehjacJ0w9
hp1C8Q+DP7EBLGj4iWrnZ+SL59enae/AcI3HeCTp/hGr7XOFPxUr5Bfe+JAcKbo9vMOIkEcQnCl1
qUT8EEpt2TPfRgyKmkKLs9fgmvK+nBoeZqUFrelzfqfA7Bj2qX4w20AYGk941oxHVuFU87x1Sgcv
0gvZail/cSyG8dmFoP7MdOZooHyfkGS/kqE8wHdFC9iJ9hElmhlOWg+97K/xo0WCci2AaFRDS39Z
ZwbJmb5vv16AM7aF9n9HjXqyI7DZ+U4g5lzyLW0FIG9VB7JHDpOh/puT2Ycl1uMPuFz13t/Ut0qx
VP3xVDdqCwpSVuY5W2kIUd8mNyFz8PQKDyJ6yGhCwzDVAzRysjoIGF9K/zLh5OAJU7VF3MCtRC1N
2nOPvPeixeIkYA5CcKrzt+oyDqYl7UHhDMwCaUCe+SriTu0c7TsUhoSapG/FUj/GOljzpp34OSWp
r0G2NZpIYjmfTBTnWExXwY5F8W9VO49F8QWEOFOVryrPqq84ohF3Eyo53OwdD6kwFBqjt9erO6lr
qqgbjNbcn6FH3zCSlW7tm9X5+oZqzMuFuQyhWmKgyihxVHaC6mteQWAfXD2BOH4ZRKuNQolNDMB9
JnZTmntq+k8N0f3SgN5L4ILpD+BHLpGwG3Q/Wl/N8y5F/1fqoKNfLZw+0NRdFD7yPED1ff047skD
sBh4EyyRQXjSpEjkrB81N8TGpLWoRV/nD8LwnwfmWSIVrxXKbNz5l1JInS2NQCBddgIrkHocSczy
BSFEyNWndIAYUjnFdPRU93vUpx3m8hrOtfFcDqv70q1rRzz9ek0nE2yAyqzJnrMZPVDyJVF469Pp
i+p9jH+fBm1mxLrYenHZ0YjxCFLYwGGyJHWejQCLPuCytPncZ862l+7JHYPahxK56ClGmaKMr1gp
AxXJthKmGCU4IqwtUbtw1aGtdeCCfgDMJyGa0PSonXwerEjYybx28DPTUeBMz1hXyGden7N9mwKp
Lu4DzzhnQ2dckOFPoc778wWnbV5pgdXLKPFfBrH9uNvqf7hkBLJtWGV/PGegqwpon7qpMG6WsIio
HB0mTTsxb+qRy9N9fb/pj1RPIAop5nyR/SLxB9MiVKkPNpvox+K5nDoExmwuj5i8ASKUgC9C6OMF
wEROEqxm2IgOyk983rSnnlf5hB+C6gO6B5ENyUrxVB3HdCMwG9NA0CDipIvu/2+2ciE2ClW0cr6c
2YE/tRE1P/NgxjIRfHgouM0a2trMrGFr4X+2R4ghOYJhaDMbm2bQ7/ytFJdrZhqt3wqCLTrxv+dh
4TUgW7i7kfZ1rS36pepbbWFMNsMk4pNy7CLCI2wCK+FEcwtvPW/LTbMaXZFeO8E8urRxG3PXZl/E
NzGOocsINZhaj1D+BrmgeBYOkSwU6zWZoEWqUarVRErqrjFTKDxyr6ph/19EvS3ekhffHgNR+FwG
FQW72p0kV/APfLEVP+G/KUXOSUhFSV6t0HFv+AfLZJ1av3AysXlTOE/ivSUlNs76GLJBQfzfCByt
WSF50Rrj0pgrXTlcYR9LdeLKGxCp7vKgL+F2pyYCtx9MvWB8GiZbj4T/WWOBBJ/4i/9mf4yz6gvg
RfGatwWGHOfEFO3qTD0l2h6warQA/aE9r+zDJ6MAHqUhujYsrreJ+9G+elkHI4/s4dsRwED1xLYd
OPcwInIba8DyFBxdF4tkfE3bTIgoru6FrbTVa27YGESYPY6sERhAY9+vRGGAuDhnbF7mgizv9P6O
2hVzB/W3HFuueV0B0UwFhTfaMbPCWPlECguYmIZFvFQ0DuLAnCqsMVe5G8JHp0hZGKZ2lQRj2CIy
QlvwmPutZo0ZZwEn7QceL09Vb2+hgfyamNohlcArKuNxfjIzjSbbHyrb2bomBM9wNwGchxfhm3KP
W6Zp5XF3CtBzzJ4RAtNB9JwibJOkJsOKZfwY3pyWE/LIdZkQXgEwUv9zAp/5BdNITfVEh1otBGbm
pU0RcKzgBm3GQAzDF75bkOEL6L42B6+0J3ui1uTjRpKbHdRKHzkmW5wVU6ITNZwJqkfdtbccWDtC
isVC6jHaf5DcEIqmjAbEAYXPGDLSSQaxeA6BlbZsaQCspjKcAxziI228EJARL0msDgcXBRNqj/lx
YvaDdrine1Fe4+ijriOQu9++3kG4Q83+xJV+i+9Z/HeVusHOOROS/kqJBtpaB0u/1JKm+iq85AO9
bWS/rUTNpxe49Sm4iva35rJsMQOolHMQsTebyfUuP59qSrleCP2k8H1pHJ0IQXGWOiVLmWnpnDNb
KZ5GsEb/T2fplOfg8BGuREGkkecdxu/eivBkmr+LlM2CMFVpF97HV+R9o5R6IIJ8Yu2B1fqww3NJ
xufFmvN695U5SkoISjGCz3JFBAy9373HoVbx2w9V3YTNiajdZj3/rh9LTOqHDVw8Ve6TlsYGv8UB
WoDxf+Xu12N6rjDY/7U58y2uS2dfk9vBXFRt+jc8j/4peswwo/0dtfgm0zTh7ty8oZEL/bnKmxEA
13QK6CW9zKCYIL1qLAfO04Z5+B7Ig/BW+Q02AHDFxRnN3vjs48NThwYpNaP8SKJYjEJr3sUKJTc6
GQzspsMG9Ue/a1qc0Ba6+BtJ5y6b7lAASAtgFvBIfTey3VDhNPU14CnfbGeAC+2+izPWeSV9DCSa
c3I8iFZxUyu1xzfaSNC60b4H3/anmppuR5eXnA/MrhaDFqHUCyv9+EPLc5I1/KmuDWQ1jFl8/KGn
/L3kST2v8GVxWBNx8owpADoS1dn6okIrdt8QbA5l4nlD1iEmX/HI4OPdssano9j5joMIeeJSYDFK
SaxUOnZ12/6HzgjDV/UR927AoqxdcbI7IPuT0HuYEHrsWg8yeSgNx5Q28JaPpnQFhdPzm07T6ZE0
Nbs0oOdRwekNrbkIYCftli2L5uaNjnOAZv1+MJ/FMffqMX6ohLF9AEh5iHBNuPzMcXKMmfimmgo6
LolpeHwPDm5uCnXQ2ohC6Dzph6DE+7It/V0JhBn/FXiKaHDbUXhnucCnDXOTjNbkM+gM0lmQJxoj
J9advw6uNVTap/lTK0U3Ll4eyQh+4rAsztlocxSuyw+RLhV1Fu63CsGXI6cWBKkyrjyMWKDtNvLH
9cYM7M43fsOaX6Ls5Qd8uFFMuPevx2Eu8aLy4jIgrorv18sSNItz4lCeU9BeZT4qAseKHhtjc22V
txE/6NehGVEAPf+x7gV1/rPIExvsI1WSQJCL+WEb/GGbbvxl7AMOLSHheUiFn5u8K1r7CYca7j4B
/oSXCdZPq8wLTt7dt7TNXNFthJDSkl9RyCWQlHcRiDhOJ2bXuzS2a+0WuoKhiZklrFnOYU0eNRLP
J962C21YvuZlI7JnDK4cVFee7VcIG8hjYN/AO0Wnm2qWhHjLqypZUjZx1/ia+OsMD76dDJHnnOub
Luh/MVmMo4XBowtq626gWZdVuxgfnakP/BDA0El7o8v11sGxJWK3h6GzJzHjCc9XQ9BQsKcib9Gm
UWZhWltlpFRjj6GjZr8KJEr/WJHAkzIAkDGn3QiezrbkQXvctB4K1rBwEIChYLuvj103sjHGuQZ+
y+TESZY/Z2FOqkUu1DWf7onwTD5JuFJeIvq4LRxnaAAwC4iAw3e/jeJZ/U2dl9gu/Qptew8x9Nyc
POXzu20tH/WFQ+0+MTbU+VqlrTpLAoST+3N+0SKyBFRxql5LXPGL8rH0nS33UbI7RXz/AnKrJj7s
X3fj74OxY17529gJkX/lbveYg7u/e+ztkzVP6nIP5KCmjaLdNEMgcqWaBPUp2FbTH2EP4o+V2i7+
z/OqcPhHyABnea2Pu7NOrbb55iQ67SZ1IU3WOx+EsD2qwKTo563c35snYnOO8Nc/M5TMZ6nu4Kx4
PXJLLg/DWgP5Z23OzucMQiNXW0JGhBAQu/25GHUDLJQA7Rp/rS1JeQuQK/mYm4nTbg2TeUT4B/4P
F9JIKAKx4x/0XzfhHciGHlc2GGV+UFnM3oHG+HOGJDsUvvj62K2WIniGk/51fjiRw9x+w4I/qe3y
0WD0S0kbfGrzRatZYkXBLIuzJr4LnPiu38MlI1urRxKHlmabmoZF8G+8jZMxn88xVrdQmzc1m5sI
wVNzhQNfK7/TGFfB7lXpqUJVwftD46cIOqy1hfG+5DyTmJmHNWyJ9L3sq0GWJZCttlxhYzYqB5Tf
Yzdhm2L9k+ggwcY2OIrS/ETm+BeRp30ZcybcHlMtKZsUzlfOLNLdsvjLHlhl2kRjaq07R6FNbWNP
lcK5X4LXG0y8WyNVksHkxg1setjfXxJm5J78IYfdMCpTMMf60vdxnQF3epA0rCVI/DCvspPJ+hWF
VdnF7Jv91rl22mY6anlDwo2T3cA/UTUtJLp+8azGZC525fytSz5OojBwNJ4/NLkM5Kc69LO+5vlq
0Eqj1PNyXXNW//6UwZVlFy+iQ6i0ye9XyJ6D5QMWlqLJSgY2C8SXYL6GHbQz5UVoqo8R9Z/VBQla
yGTZvfvDUnRPwzpWNzBMJ8RVl1cIt/CQjGuW5P76MJapc2HqgDjE1j81J+kM23YBrcqrJ8sJwf56
kz+y9MOaXy3DnF5gzJYot/26QoLPwSw2i75kZEJa1GVywdTC+48dN1l2fHeYnA+yENpdlOiVh5h8
yfd0xP0L/dAmWV4Iut10+7XyV30W1duy0lzaMbpqmQc+6AUzTDC8sVPnvuxe1C6Lx7cVl/p5n/jQ
+yoUJ5OpKNAbYtekYb+eoIGAakoAYBRgdy3pYgRKttyFn2/oJogbg2m8YB8jmazl0x7JRnNmYMsH
c8IfLrsiubuCQtySMlP/DhqPdm4XSPGCf4x358WlCODj9AK+WerDw8K4cJB1RwzBz7C7f1elKsY3
OWQRer8Xj4RLba1J28cQxmuOWPqRwCkzwdRZ5Mfb0B4y/CF+1wiUJHEoSwAkum5w1hth/5TNdYIE
QazW1Z4O9SVreHThHb2R7dqDJw3fRfMddQctj1pbp7ymGpglVwMF28fMkQVAni8fqXrjey8lb30I
dGXGMb61x/MEOmVhc0n95nSCXVVP4+BRbPeWaJfJffEeFpeYK/vyf/y/sRJjKsbByQZ1yX965Elc
SaI1cVC+QAU4P72oOKwLv7FTevSbIPiMLu80V0xNZsUOEX4ArLXAZ13S32/IbwoO6Hjennrgpybz
mbm/rnYdVkIvpoavw7JNLRGdbHqnateGY5toe6p3De9iFovBa+MFuRQZ6k7Ks87B4Xuf6883xaqU
/74xjkP4bnu5J3oj6yF9lmmiHGQ7nmDoYxeQiHV8iegWz9E00P+9x16DpQQ7TVjpJWN6ogAaXNzW
tirfTO/KtQimypx9hoUeLAYB0NvuHlWCLv/ACJheyWvQx+yQZHbZhgPEr/MP4kIAlBYyVG7FWjLc
L+raTiPb8peupTYUVRpQbcQa2Z6MqzfoJj80yvF0LZhRYF2MJperV8z94xU11V/AqBjUhPAIOuRA
jMNmIJTHvMJQgU1tcypZTIvh28PPjbMyIyTSicYkZvEApA3kL3SmahuS/dM/fksREPxOjgIef3xb
aEUTx1z2tYv6YJwnr8CUSDK9yN2Z6m4LBQnC8arg6Dk8h5NZrxO3F+H1gXcIgFyyXSB3OOfFaTee
olP6NmPuGKfy6BA8oDd1lk0YhbCEZA5VVfuY6hYtvIXUX4ZlxWVeIBf3byi5+xwm7QukdWSNn5ef
8C+MPjtULxpyh6oEICMFYzDWP74wojR2Fl10BmIj3ILqEEFGrwS/Zc0btfbGUJmDjRguBKmQ9GAJ
2Epr96F9IUxkgf7//Uz/XaVHzMWA6Viz6i1n5knlsORUVDRiZr6oQ7WVoV6J6v3jxq7sunvAgJB+
sZ4mZ+Cykb0MO117rht0TN5lx6NB/2wCoo9/2B4DizlzLKhz20l2oxaUVQuFjeXHe8a/Wtpp6Sn0
xqGVV/TiKDvnPHWNMZ9HehEo6RCMDKdQ2RoGW3oHtp4NX+akKul9SMnRv7NHU0puny4N4WL59fME
fJdNjHCa1MMfXAjVNBtK+Akf4JAfuPSa7gYvw+BRpk04JG4D+2KC5mwRE5p1BZKSP4h1Ses1aaxI
d+dUWVrby1E36dL6kYOcpSTTanysxKb2hXX4as0Y2NcmHgWyGnwsdO23svCz8fDYbmibIE+kc7VN
90kmviZtq+Eyqd2Q25p/15UKEdcBah7kqZL3meWWJ9pC8oWcNybvsbReP9/zP9yULspi7FbxxxfI
4t8s89k1+6DnB7u24IKc/7mrpm89jk/w7q0QyrReXAnRpzLNz3sc26ol6XcQ4yTKXiwqQ0dJYQoX
OnO1CYT8HEq0lrVAIi/fzeYD+ZWHRl4FcgmGir51UkdjBwLqLFJ8jDhiopKhg1ApkUCgrYBR582t
psf1FiOBgD3vo7QScs9KtuUpPe6hzjSFYCqDHMHgbqzVy9S7aEYiUqi9Y0e3WW4OLGuwmm+qyvQE
nbONtOjFbcswIvr02MR6+grtXcxMs2YR+M+M2SmlyMu6j/3NSmvMGcF0YJJ50HCHfhOW+mpL0Ach
wUE67NoQty3a3EiAMdPNevoX0+DV0SLllJ9LYjs445l4DLBk6AScsT/NquQpUj7uILbpfPml8+QP
xPIiqOjLJyobuP7z9aVtUTFyZxhAgOch43+ZysHM4FJqOsOfoOtAWynsU9X+giqpw3fL0xqRsZkP
IaIvqAFFi/GGXyq1wz1rfWssxfnjYIRzG+D2girXkCzn5fMNLoEGNp8A12xxJcVkLFsMGS5n23CV
1DsRy7TrXARzTt+4PoOufa+ePu29eOosJJObJpErk9I1NuYFCasC/4WBeWJVaNxn9SnaJhLPF9I8
/F+C+0qIG+Yb29PPWRklJb6/KCycxkjM8Ujz7QTUYmGxbfTPXYHHB5ICKVnuyhbQvK2UkdOlxcv/
P/MsN1gnDBK5SE2uzNALX4bZXwNVUEUfie2ASnkYAqSbb0I1FksyBcSTaIG0sUC3CpQzlRaXILcE
4fq9Ud2yIeFnqgWo/1t7QMXAj6XtXTdg3tngVHe8MQtM6E/qQIr8T5JY9dHCwfBhXxKNJpGOx5rl
QhWj8Pj6TRdvXQfbsiMTYxpUZgKjkjiMnjzlYhPT8JJsQzdlJSy64PIiFYa9y+biAchXXGQ+/Osb
pGajGzPUaTO+dILArQiGxtGiygOrGYv0P4VAvHV2Z88Fh04JdoVIaCG39HS3V70/OJTwM7LS3ai7
tPy3QNFVYUhCHvSm4dHfBUjmmzNASmwJpQoiZoyS4HOuHWiY084YpMb3IH1DrUfbLM1Un8UVHlEv
y80AYiVMwyk+HdGET5IvTeR+LPjMHabYqoQIMihVoeaXDU8FaH6somyWEUhnzCbRnsb6TSC0O/CT
vb07PvJnQdttmMoiYMe7ZFpJfFwtKBkTvl6yxNhEaP9dvKvnadkIe5DxLd8qwjHD+xjQTEgqXETg
vgPgXnyucoTtyzM8CfxOZ4/mBRiA+8GxZIo4ceVCdWiEBKS6BEYVxlnTHGi2+qatTBeknAvbwJTv
dRoWPB9qICOrMY1dnzHFRo0ck4M3nL1jfsBYLh8Yi2Pg3tsBVIdX7u7HN7+ojf+lt94GMJ+0ZIuM
78LVlSqTevV3+S7N3wUZCaERXqKL3/Flo1V0jgejCkWJzlEgdEmtI0f3fysoY5sjivmxpbJZLL7K
Y8giDrjlvSaSKfNclvk+/ptM5GOhMyRkhyHQD1H2OkSfwo37gSsYpR5kIKJ/EQ5YurdimjY=
`protect end_protected
