`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11888)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMKSJF4ybxqqynmhS2QDZyMomYG
NwEXErRX79D31/2sINfq+xzV/Btggw+TOlaeyE+Qm1kgJzRCIeDqbrQotdZyz3Kzm08DHRPhrWf8
hGCGTzdgAAXIbXRpafnrxPi+kMoGwxrPBCDI51eMq2zeHHZbyFlq4qD8zo3u4h2pZWzhv6JAY3Em
bM9jkB+watnG8r0lFhof7uaHY7Oy4bRCgpUzyjbS4tl8MrdrYY4S5hgq+2NvZlcHnMTm1Ve7T8LL
KcLoTbglm5pK7WBBsLqmqI7Pxx893+lCw+mtG7vTNIlgydprZLWyuJ53XI98Un8IIhVAvS8PWhdk
hrnOMh3hNbpijDUgMPCddnPKjVML8OBg/Al7niDQ7mY4MZFZZxsok1jDPtDv0UEXyMLcrHs7oJ6Z
9hYlqMlUab8irCbEcJ6oMuBBEftnWJdUurBLamwaWUMnw42eynwYcLaJm+MRr8MJ8HFnUjc773Qs
vtHq3+nyidQFGenADw1SLcl4ht5tzxLRmxW5ENd3eNr/Y3qFjjEQiwSXYat/xLEYyKQNZrtNu9QJ
GI/qw5aE0u0sbWSP0qWvzR6KdNriZ65kT7ygDd4haxKMGw4hZ+19j/9jClZsyqmZuUvEikdB/EGt
DRduZM3O8feC8VY2Amdg2HgufzN5knoaRKhlU6zeV+R+0LHgeycfYtns28o0km9BpJFW03Ww2yPJ
s1sNCtHVxAXRjSUFWVZug1NT2Qe6P6wpCHtobWb57TLR3v3TMUZ8grRKYse9eSdvSCdEQsnaoQNU
vy/t4co2lPPqKwP0oj1pmFn8FkcV7t8BmPzuQzeGcn5L/VrmF4XOLMuHt7smOMZQUiVD513m/y4M
FJIoSZKNY3/xhqvbUxdDKRbsxvBMVF1pTzmYHClvz58IsYkhHZXhSH9pzHEIzzSJii5h+1YTmLy3
Ldlmtqz3bwo1dTrux2BSlp9LOpD7iol47zaKdnbkxsSnYMUEB9AmKPjOdRj6vNgsepali2hsbviQ
Nb03YNTU9jbcmRmLdO19bh+HZvq3iTotf6Lw1tykzstIJGgF3rGhbiMyIpC5xy6Jqxo8AfuhS6FX
gvzqwUxmFXnXm5hl8AhOT9ZkUrTezGcVrJai4EBwEmdkeVNQ3d15y50bIhxMZcbQcZkMq/khncLH
2uEMghMJfCIJRd8l1cQJprarC+KTysl2Tgxz46sJRLJoU5Y6t/Ka7mbe51kmMj5ydZ+HxAz1EnaH
i9iFkjqC0tMWIkprnZKUlr3awFW41X8PL6Yzhh70CAhZKy19XyDrOSHI2QagWtzoPgHEUXuwqUNj
OypLecxZLqQBwlewsdReLsaGB7NvF+bt+bonp8kt/XytaJNOu6JobEQ40Ud3OP9HSpyGB3EYixBo
rGyrgKQ48o1kAFsh9ys5YFskNLKds5eE9OfSrhqlCu91ijKRv8ay2gvdfnOeyYWWEb53KdrWzL8X
Kqkq2Sh66yhPV7CTBcYT62PQS1vQC2+hzKafXTIAtqRHInd0xONutMHFRRP7A9WV3aZ095vZ3yni
S8Nv4PfGlr6xAx++3nKYDcsTk2RRQEkCC73NXAKDNn3O7EX/Lh6gqBMR+uwqYWsLHTQysY6rO11b
PM/9s5WFzYif5TJtCoIEhtiuk5+f434sfpEct824ExTW+IZ7o3M4EZctV5WoLCg6Nemt3HpGLsgw
CqEhiSiGap1OEW6BOAPmmXN3Myg/xvFsS2eeWVARK6h4rr6f0JwjHa+to0G8T4OKlatMgYJOtX+l
qNXgfrUnOkG8j4Wc0TKzGM1nDYnrBpaSPTtn7CTA29IjqEus3N1z0oNsS8uWnn7tOJJDM5fEGSeY
quF8VbzLj/saqSJzG2VpwoZTONz9LCz7yqufSGXEdop+9BEqEe5SpK4ClTXK6il+a20bldsaESlk
xorU3ISftAIsnZuAp1Sm4TiJ83YZ2yz+knmMtb+EiRWAUfXN1KZA//u+MI60so5PMyrPXrYq7wwc
g/IG7wr4ZgAY7mOuKRUxLchXWOupQ13JgTg7A+h4WYomNNw2fRJnhFeyNi20Jm8386vugR+iny4j
g6wX53ZspRNmiByHV5luffk3GYzSdjxboZhiA8QNDnZFWIpX+B7cduVZaJmtJah1J46KGQGhB5iY
399b3dbuVjsnD4uyp7bRiZGGQPvTWM79eUOym1iyMOlMkYmLLohDtnoOXClIsEZkHkib4hcHqhrT
wiimkhoeodTI8OtPf1f19b9d8H+WVF6Ctzw6WcipMH7sTaP7SE+CJVx9JVoc66BEmKYcsLWyzKtJ
eM2Joxv1Nke30SdfsRDdPlG1O7ov0yimN94Y86U+vvI3N90oJ6q4wgzt8sCBQ2C+GaelxJGqR4ud
Fy8LZbpRgWOiS3fjJ72DVMxVVwSzCVliOYiBbheDVr/5UEqMfJIN6r2E7x2QYO4EPsjaC/M3v1+r
cBbmUq5UFEDx08zCaK+7cz6YIvPxnNPkvWiKXYgP7AFffZx48IPHgPY0J27NpffUSupy5T2pvI8R
10qu+EoQ6MFZL3x3vZlWd8VIoqbrzj/KmWY+uZOYTPjUJ62U6Dmvh8AvozB6l+7b1Z1QuWT2b7eJ
PiZxxW861aIJR2xwGshxFeLzCzvQkxkNyJkBcwnMySJb5Sh5R+UcRDwAwfF9F1uXzPnad4PLR+jS
bDHXXt2sa5AybU0gXx1DzRMPUSAMEtcJPtb6oYzWIyBvH/iphXnoSK29ZAh0gwY9ug2SQdDlR2M2
kT2bBdsiOcLUQhuR1jdOKOIi5+h1ey2aOqzfguUXDeThOCQg971CH1V40P7KQetHIkyJ66y1NAjJ
XBbFitDpfJW/VK97fBfAi2X8kjXxUthJRKdf6gDtNCIKv1EHk0q9eUyERc4BAN3pWNdpyuaCF5wB
LNwBF/8353/rF528ZKrYC8cFXUiV74ul6njybIrhsJ9MZVSiBOuslViVkrKYB2+7eTGDYsW1lht4
uHDSUKVhhnhtLlN7YRUTcOWLAwKziCJ/QuN5ERQol69GVFdW7oMHByXb5SqrUGPVXmi3kbZeC6oE
/Py5RbguqS4znhjGbN99N/o9e1SagvtIhBWcXNO5hj7yMObM665DD+u+3Q929Ljb2oQWTOFKQMM7
etGH2+kvyJYPvlZ7UddeNqWYRTBH3gOX7e6FwLDajJExzSFoTaoQquZaY6UWlOb3x2F9oH23XBGK
f7s+y7R5LTFw8kN+0zN6zAqIffPUve+v2t8v96NgSIvJcX16Dwo8hNArT3oVEWCdEix/DACPbfuU
AZ19kLaIpBwfqzSNtoAn5YOR9jqgQM15sncKGumgrqJb2Bv1LAXnG5kKdgxBtkBI4ILU9K4udP+k
H+1eY5CxD7GWPffWgVQyLHrcUCjutFURycCBP0SeAtCJVbUfy/RFS46Ehx3x6UaoxORr7TX4dWKM
/05VxJVUx1zdgMyjuf2BZTwApQBFDoP1a9bPdezvUjy0l9XCMnFvYWaF/G4/0197BbpR0XYBLH9S
UVbB9vV0ITcXrLEVbk3DzRXcN4hAvewIpOXA7TQuHF50HHHbxSsGxAmNehbe2q12oCadVW3KFZ2N
gqIumMMoCm9vC5+4ICGwzuZ9k5aQuEqDSPxTrCGXtvnrpjbnuQF8Hxe94juw3dLeZjTBFqS388PL
yv2DIfaA+Xmu4dDBIBYS4a9xx6zBnVMz0w/pSVJVpXEseJRRh3LH1LXRXxoejMd05fUeEfOulZy1
kyykWNaGsPljkziZjT8CTGQL8WlB5EPEB8Ncvvo5B2rTbmluhCZM8bPzd5QkJphUbcT+j+kHZ3vY
F9uQnkRRDV7xrZY1MiDWPfPPLXJxpY4OfWGDdDfUAeU0w2u9/PcNuWN1O1vqY3XsvmWxzQA/IGo7
DpIPOs2LDmcf2Rd/dgNMLG7kgiKhNU0Uko2BJ0zbRz9pzLoK0oZcIFuqQ+tywK6UA7tpB45AvI8X
mg8ht75+Yfrjdxx4t5Q+k2VCaozJ30L/GCUMbH9zpkKjM/pYkPS1BHDek8/IGfpXyEq/LowJ7FLp
jT2IUbMKY2LJ1+5eOqqH46CKsGQgaaMjB28IiKOVTZt0b4th4uWD3azIcnmex/Lxn33+mFRro1Gk
OsIkEWtUKxj22dr+EnG1pVtv7w78gIIM2EX08YciMpUKAQtoQ/+hcR9KAHMLGr8HN4a4bDwQgNZM
Rqhth36fiF0DtQn/+33/0IFjy+58URecZJieKSt+yTx1zhhfO7dye/a53SazOryX5/7O5FiQV5Kx
U5/n7bD+OdiZ1yko3wgZ6nROaKNqygIxicY86KIENW432u+EKJ2RjSPSqtP7pJa3x6SNyJkn5UeE
uALC+mYc4pNecp2wChdGOQDVDKTIsRxLpjaWLEdU/EUkNxZaQ28VoqjiFPq221sqNeUnTFbpKwc0
ggxighK2sQjyL1kqx5SawnArJN4VfPvOnxDO8BRFbc7VmxY/ZJVOX9JnOD5doneyxgbtVKe+eAOw
AjKJoCKQf2qfKHyHq8E10ctBD63AQ2esYNbcAjSimfr8tIQRvpmuR+U2fAKs18kdLY8HlTNaNCVm
Tttvv4jp6tNn9NR5tn2cyvrQPunjpe51CVHpH8GtmJf3APJNaVeQrONgoKS1ruUm4FgZgBlIHIJs
TNPEzUDfzVlqA2IOYYN0PBM66z7cGFuYlqHh/BBPHPy2O8zI27jyq4lmzwV6RRmbzBcHg9Hyvesq
HQ8FRFqv70LDAWk0T0Ah8tfKpNSAGfgMD4ivTN6FfjLzO5DI3rAsVeuRxmgOfZfICHZBLCJ1ZYG9
dHIHpx8fN67hCBCB+37Dw09GR/mWt+cg/HebUGFN7r7pN9eExm8y2fG+55ahj7+NBHIvApPLnNzR
v8reZkwu2sxxm2wnnsnXeFRc81Fu7OCj8++ZMdNfYakgUd3r3SY+ED3gJ/BQfpDqF8bQbhAnhtgJ
BkHCJVnn8pznBfYsuGeBfj3P92EyrR4i5SAFFzjhZEOyJe9SRxFGuBD2avYcRJZ3qyWyoCU1Jskr
kTiTfn8CNRQtEjk0A5ALHTtGIhAUs6Ms/qKBZnsiew54N1X5BniTc/WGewGPiZCfGxKweO2DKpCz
GmDERA+aOcFFm8f0kW/cTsChaLFPJ8av8M2fgiNNQJ1gXxuTSmA1lIdAzKDycaSdIPwaQoPIJ6sd
9M522v8JEFJxd8ASQejnhQIBJYACBsAyCuGbGfQlR4zXOnlw4JAXCkHqNHZrI82tDag3CRvj0yz1
imfg9mtLESEUa/ZEUuMqyWmy7uehoNZZQ7E0lQirjtQuMkLbA9fly0bnm4+b03P+hQkVdaOP/BzI
kzFX7CJPOwnuvcso1HF2LWCjsD0pV2ZT8BobNx0kJf8/oIimCbNk9rdr2fuxrHQHXfSHIfGMJMBs
YjcQmDrdJOWNEqjL0/XviET9QMb+G0YBqVpNilyy8tBO0jbkLFAt1YDMntaMIhX90vacGyGpXkJv
KuwLlsSie1o980jfRyPhuDwieYVqIaJRP6fgUOfRu5bWR0gXwf8lLY4dw4X55FJjE/NxnjddllG2
uSllPhp6YH5Anqb3AFZuRjWCY2lL3cRZFqNUWlR9rFklDa0gkDULrBTCgDCJEN2OQFW/Ux+apYlh
ajKO1WQ/TWbr/ZNkNevgmA8opprzj35ZHpihZSzAScEorFrKxvIHeMqrb5LzLXGIyoE7XJpGhxaN
4artljc+yQwHStLNsCq8KlWfuB8VEqgwrChWVdu0tE9AJjuppTiRj9F2g9ujhdCExi2OpZ5j4Df7
/v8PLfOG5qHxzPUcB6errQ7udYSuE16leqvEs3WQJz6VPLNKFOctqZajuXQJo3LNGSf2f5jb3Gwb
VIkZyvT7GHxp1OSFLPljtha9kuclvnuMV7sXPfNIWfnaXWvp4yOy9kcsjYY7jXvRzYNOpokEZ1eD
G2zr8FjH3ivni6m65JQqtzMBYqOJ/tM08xw8XKi4QggbrfL7eCPAeqn1cnf9XXCbnRS1JTupAe73
0QN/sao9zFWMCg1/wsePbbeItx0LscbfeIXSIGNbjZR6t5TiMvDeCwcYN1DZGZpgFaCURcmNjONF
UK5Lr+CJoIopGoSczAVL1oZ9Bu8kW1IRGbkeldx/xprlNzTGtGcMTwSeTSBW3pNFOuYXF8A3WloF
IsvkUN5zpzv0ePKExrGqZFMm8/0LnW0dYzv7KYLu9P5hDX+uUOxA8je2e7XvMXVrV9LQtMPjfODW
0ervcKyxo79l37tmLoH8yuRT4rVTMENt10xRolQRHwHcCfJwqCNEK9aOvEMYkU4Fy+1I7rRLe6+J
gzGvls3gH47gW/SkpyNnT9jI5/TMiI6vGJ9vUgSjjYsePKuBAo61YytXZLoyvV5PX2Tim70Tak1Y
64W33J4EX8hjCGHV31O6aalCxaKtjJbPsvLTFEZhDSUDyWDgmwgu+EbqJ92u5aGAKQKBUKQr4om4
cHZQFZUvWZSglOwh2SMduXefXei16UGxYaxGABREwSLYUIKBxu2vvLl1effBnapFBQYyLki6PhLX
wN6zLRUBuCePCMQiPtQjYVbvRgTNLa9mfRIZ6k4W4UVeqPbFoqYoWM5r8esdeNoHowORb+jay22K
qpXpNfvursVmAurnFxsL0sLl1rpIzVlEMV3xHeYxIoIeH3kpG6HDUe7d3XSJnOqhyNq7K2PRhgPv
lJvOVem0lt9ofKjx3ZYOTjzA3R4bZ3QCg9pGZ7wk+OjWK5Nd1xTYh+3CwPC6XozLUJj1VfVi6qoV
u2nWHSn1nc1eJbC11ZTHv88NQvsNx5kDVUdeDjDt0IVnGElz0s9z6PpOgQ/tj5sVMogziGBDVWAa
EO91WcCcwM4Yud5Q4ONr5sx9v3NQn0QhRGZbdIZyRRKQQ0lOBpjNar6b/E3xQ14d7zEHTFXCVzAT
zKP6eg1MYR55pCSMlGJxMbIqfIeo5bu8JA0pCiv0E/WdANm4+qdU1NYy5wV/4+6kaYs/z5KkYRsc
y480hSusvEiHfXjPnsvghaVM/ruJzEu2NBpagKStGBiBB0XfSKk77uekHGZC2QgzpR1U1WakkMpd
pBm3LFdnA/kKNYQSHlZCfnwAcxBMoediQ14R20ZstXzP6iHv3w6mYZsutqgeus4LotofuhWmQWqs
elsWnnCX7VccH7NYSNUY07xcRkUK2nuLoTN4M4oQaobe7y72rJprv3Ie4zHUnrTVyYXCEh7kiauV
bpgIZrqykTkzaJJUVCvRtp0v1iRi1rUoUEJvQYUDfHTenIzqrv4hRFi6Bqj2Dm1oIyQD9ToU/0Jh
MjEmIfYfOkMT6yaBJHESB0NUsbWTCRgsEYiJQaQQYUO18ALS7dSlSA7csm7ZaY9hVzAXiQVyAQRC
Q+qtdQB4H/cqfTo88Vf8LHs+OHEvQBBqS36CsS4u1ZeWlycoABAXvA5CTkCFVhI5z1q4GZGHfqMa
fAeTj93gb6iUefEppwucF8HdBcHyNKguCzkOIbkYp0LZ3ewwRhKqe2+yZiFjQcgvK4P469AlfuYZ
w4Pj9fHVYYfUa8rcG1INM2H2zm3I0o0nZPC5IxUEy/9v1Ka/mwVN9itdoGBh8924EcJjoH1m499A
OsLPU02b7K9L5ONlcuNQ1K41hw110N11QhhZsRqZpp3DiMaJuJH3/fAi1aXRIYomLZoWyotBZ1sn
FH4ILyTK+YhnUXjBK3uxdeNnMB8JpQHxXMs9Gh5Kh5jH5V0mM1RiqK6A7wNGJkIyA/VuWCXCR2cl
zcQrlKi1N6/igUjupY5qXEq9zYALZkxsu8mHohhQSTBN5LG29Zzqb0udSybqK976zmzYcinGepwz
oiG/PsWdtbj6KnaRvRt1XQeKW6YpaSTIpp+yIUGiaPDvJRVWZH25GBkC0yPbgc+VOEt0SpUrGnuD
Un7wFEjFg0cw9C4MpQOmQ1Rl6gFozIDMsMsgqDqA7O6uvQNmRSKdlHm2My/7V+25eulo6vQ4DKLI
4XMm0n1oKJRh/unDFBpvyJOfTqNtJou7b0OV4iUiye8h432gfYIt8HEk18ygksXTGrRNQFX9/h/E
z6HOPBAH709b8Hl3WtVVIZ67vFpoTyxh0uqN5uIi9o0+mu+WwKJQh83b1HIqEDw6Iwyg5hAUmgJH
sQgxVd95dVyQwuUOoTJrBvWvXyW8Yg5bPrcVCwpR49ziPZht3tG4q4HVpsJTWSzY92FVlKWlpnHG
HezBBBRwB0CrOKug0A05EpbTh2m0iWN3lA8s+fFltsY5ukIWc3URsyz9YFK5LN/kCdYvJnFchfOQ
BeV8YJiWn1s6YBPiRVfGGqwjZp1FLPeIkZ5Hf3Gh4B/8PbrW6E1lKVxYRepsypBPkuP3RtEfmY8S
PSLX9aruo8Ta8yocmY0oZ7Ff373jDQVnj/afSPUzsjKDbtuy0pTixS8J8bdgc46oR3WyEs9oXozY
bZMlApBxEhuhAlV6O+5Ic39C8byp9jyjTyS8KH9hdA7d55dfeilzvT4GAJYZRX1EtwI1Sry283BQ
5u+7SK4LhU56q/UcZjR4uTVxn2YGLOPZD8LJnKz1TD9px4RPaV9WNRtGDx0AAqomNroRL8tvh46l
O8uLxFIvc9uQLnCU1Ln9rjXhwVTRi50G3GL16S3D5S1UNAkPWcVDOVmBncOpZkqsCKvw8qwt9jN1
h9T5sew4IK8L9Rmv2QyC4u3NAM7hZR1htzf6xSMx/slUrI7bwIfRmIptmk1IbB8Ibyx5Ej6IbC1q
rwvJhNgYNQGNJi0UETUi7HknRSBZa+uwuwekmeTMyfdaELJtD8M75TqWe1kyjYzrc1xHdut+ywBA
xo17DA1PhS0SDlbypk+e4dE93e0R8qCdGlF1bZMjm/cDwtWtwYQSQVKuPBPMaT4GJTs/LAlq9ZSW
DBpVR8rYtYIdoN/DV691urGRpQaATh3AvDLO9Hp2mCVAzvH10JuVT863WE3e3ukb9BS4IcCLGqOd
U9irTQ0U835Wwr78WccguduWSt0dcEXR8F11agPlR3otRdFCWdYZRdZ0j9G2uAqf2DC6NeI/Kz4c
+LOSB4FV08nbibHhNadHpEQvdty5irOIgbemh14+HYn4wuDJsFNfV6JIqiiKJ7s+rVKaF+RjqEqT
DcolhCUq6mLlnXus8d5V8Ae/rqbmWMsfMz233uOtrWfd2vjqvioHuCy3a5ZhfaF7Z2mQnX07yB/N
7MBrk9fZIcI3kEwG7XTkQkkQRcmkYjW2m2rD+O6LIyBDgLzq625OXhMq8eQNf/Zilp3kzYiWGH2P
prY2abKdI2/VsegJRCdz746tOjjLBzQ/8qqRN+B2gPwYi5hZ1yi1z1fC/94lsdBVieUNyGA7s+vd
vvJgD7GiyYh6q4rLSOvN46cCs+8gtBXb/uC8CEWy0dQCpMGkmpzyvY66i/WB2P1jR/C1i3G4Pcz7
/oaMsSDnet8wJF6v3a2ihYzD6yF1qPOU8Ohfn0xm71ONmkVIIA/WP8aiApg3Kn/TiQZCuIygbml9
7arb25qjg+okxLXLj+DjryTlTuHbIJZ1B9TCC6gESRMRdCOgTJhoNbDpHjxx9JzqH24Q9S1zsaRw
QcX+WErxPsen2XogVU+9mMXhRQDZzaFwgUJK6Z+CRIO5Oogaj7ejbBo0kHVzR2Fx4Q3XhhxFYvJT
y7ztDUeNSh5IQpOnBzDw7pU+Y6F/nstRbi5Pjb+vuwfrU4iTJYjcCGT7g6ceVIguzshLoxqBhCFX
GFPtdezzLjsAeGVj1bqsa8/fpDx0bnTINPmAVMDJE1ELmNG7f6zb5XanKazM5hW58CaDtCOsB/4E
HJwsgyMPjroLNhIrxGLQ7FdZtUT3zPC+YuYZLUSChkztigD1cXEs8nwiGV0GS+EgBFQqzc/1mPAZ
sXquYjfPqTQSJtFwUB8s0Mra1jebvdvO//ZD2ugdm89N48C9CWVK9K/DFdiCdfikGHlZHWcDZpXK
yb9Ep76HZGmm3KxmG7OC42o3uCvN95vOg9gSmsYxj3EzJ7odIyO1iQLxMMmMoJDvpbbT0GmKuqNL
gyhajOp+LP4dYlp6xyFdC+dlBNU9slFCH6xTssbOodHC7sVNPwHJaBPesY3RVtw8jtvNOgejyBcc
CJsDC/IA1sO4w0sle0DpKlHmU8erw3to4W4v/DawP7OwT4HfroBxxgPZYT2dFA1WILP7nvuhKQ3G
LwEGywwVEc+xHWIAmn/3Xfsd7KY5fyape2y9gHjy+FLA5qsDeX4jwHg374CSlslCMFz2m34DYpo3
dHkfhxpLm2qUNE4oOI4aIKcom0r8rdwWsRWOaWbAoIkBqNPCVIS8DM9tTtYbxwiTJCzG5OEN1TGd
oN1us+LKjsMX4ZGUelWbSiXy4w6gU+GNi/WHRIiErfqCEGUieZedpgxbAkr25BOQP1wRvLzfToOO
jTsxEgugtFIv44zDqlKrb2MZLZUbS6dkDsLg1IgDvuTvJzgEk2R2VM9Jv1AMHfbYCF73GaPQvhrX
8N0bsp0S+fZ43QodsGSUkTtkN+rdf9oJ4/vq8GQG9kHGMWJR5eaYCMQZbc/4HMik285MIzA+Nw/p
OXjT+FfliUKLdSoxxar1c+TZ0Q1CQ/FeQFzcmpPd797ZRjM85eBerrrB2Xt3SCRywyDnZbgNJS0V
yeCUKuh3nhq3BYjKkAHnmRVpMnUpLSej7xRE1NhdzUkYE2x8MbhR99Uso+FZ8JaRs1nr3WnPssAf
BafbRH8xYy6X8RX6CvxiywHTe2cPeYs5WT1vdmq6xEaCVfceibFAkptJ7HOu0jUZMUBS/SK2Ozvb
D3FUuPfG1zrqWnWzXSef3/djtqKNwvOItQt4M9R8JpgCClKORn8R8rgHqcaIj9dbSwcjlsTmhjaj
oHuSEpKV9IHWR68LZ8/WRmVoirGncITJaMWshnAZI7WD0ZjsM6rAevDRpoNRIspspDkG6k873DDR
UUvXt1qWazB8JMQGC922jxoxICSR2D44WXMkmCotpm7dCo8G58fd3uIDv/I2vNm8A6ppoZ/TVwSN
uQcggFB7va93NtYw2H2naVPsOri8MVZKMdtuenTcm/hcmKxu6fUE0pbmfFRmT7vmBZhY/SkmWKo2
DDnRMRcjBgZeJZroOOtD+Z263E54sJtPvx3YxLSpO8GkGlHeTW7dK4DPTh/AvXZpjBaXhYD4vVfR
vrSdiuG4hSNKSZUaux6tHF/rwXqpdrVRh2JnRa/rNbwl7vnVtBLd52k1Gea2lQgdfJ5mziVGEnkN
WbSu1Evh24AmCJT+U0qj5+Gkr9VgHdSzuCdS8DpyF7feO1QK1Ig40I8d1j7MVKAjJi72RKkfUcc+
13q8MOZJYfA9rTFlpHKsCauWTqdoO1rFIBnFGfiLP1gboCB7J7ffj8BceTaDcuC3IA574/OrJlIa
jXS+haWiWZoNlwvrUciK3Fkzm786q5ebGz+oct9nMn68hXGW10bgaHjQRCmRnl0lopMuoN+d6yuQ
Ky/CMR5BYkXco3Cx2D94Q3jY4uanwR+z3MT1Wsnq3y4GX67N0uDRAaao/nS5ILpE1I4DFf2PcYII
15FLh8BlnqWKZr5q8mPWv+Ek/dEqwtVIjeQsBzXqzd8t0ARtNo6CIErAGr8V2bR3jiIoFKhJw/kj
5D2VJA4P8lceHEudO0Iq+QS+5aIyVsvbInj/blZp78rqoyGmitaWA41giJzIW04uCd2YEw6DuFAX
WfiDzKzEL1lsv88bJ9VQuTzDNrt3bgZ+AgfraI0OFIwVUKKsmBZGihG0CNI/RcY3o7DACTs6vzsa
h5ShRLoJImGlnis9Ekxnlk37tUkE6in4cLy1RrzOxwn6orfSyDeNxnuhcbS2KvrgkamQXbBQXs0m
b2oOvMxWyiAi4YfJ7JJW1rFkaijSArUzPUFGwhxjNiaLpK+NirSt/J+BqxL7hKarVe3aEGAviPQ+
e1HEF3bW7py9UMThA5Ct/DceCE7ceQNqNoGw3Llcbc+nS8SZjidteWgn238Db6xU+qNwoUfeDbWe
Wv910TWLwtMrv7ruSA7bb9NCGFvE5ARf0BFOeX5gslaTNM9praiXaWVP/xjDqUlOrupC5nXd2Szf
FIoMJ77hDXXCGLexrEqT/mEv6XH1AileKpvT6wOsB06cxgN4t45y01PJyQIcQ4iZ7JowDzotXg9c
eEQu/yzF75eydwiM/pwD3p82IZLHQgiAJnq58wPrMd3w7NfSim6p+nYOc3nJu612CwMKJ/359Eb6
UVgZCGbVEGfBOFNty5ZLHZRG7cn73qUwacb5f02ogBpOAUKH1Cw2tUOxbtY/+zjDTD1nwxhqJGFe
AIyIKzZJEhXvpBjvr53lbcrDD1ccJgHhrz4t4aJAdqqbboKDW5HXYpGqM3411mmmZ0wMCXw+r4u+
nwbpqzbif5GPxl84D7b30anChLUxV9BDwDgL2I3AzEv0Arf6VDBH2RX8sRSmExPj9ABv3j3wpsKo
W2kBuTXRf919ikJrgDe74vUxXbO6wxAUIkLUaeKG77b6Gb6+MVsVdi7BALUQVw2sm79n6pUb7K/a
zRoDGi7XNE13uKloCl3WbpqntV8mtfiJ8WH3Zx7DXWRbWgRywkvaNSf71bRh48DCe+4/IwPPmGB3
MYa2HmCXeuZ3E5Hl4mnmHQyHnoo6UdXpXchRdZUYuwvwPKOsvdsXUha+zljXMLPRlneNhQNVVdxp
s97pj3SfsbO/I4uB2A/y0fwbcFy8K6DFawdpiO3a/IuJSzaB76kG6LqJyduBLYHa5DQVTuO62VMM
lecfrUL6ze+xle6NgEf1NavExQ8xoLK/XVp8ogqble+ZpxzTwfzGQFxV6BU9JoaZ4vZkjdQxrQVQ
ZPw0Zl/6UcTHplmk72wFxf71BAE4LIEP6iaqdN5tTX6nxSbcUTraSLMINeEB+TjkwgC6mazSyx+k
7VCpcSrNzboIspFarsOjsRWRv0nEj63yH28tEHLLySakkHNy/vdGRyt3ssdgFfWxCp0NBaxVnYDF
PLhUuHE738pac61dAA3bTqM06/Avwbm+5Z5owEZUWoL3rjlhDPOjzMGBrkARQwzoCUocZdtEdq3i
9ks9enyJhXK2tLopxiAbw3Lf+XWTuXdx1cMWayNFiPeu277lNOGYBTvTNLgWtftZNBS8dO3KK3JZ
PnbrC4O73Ba6pafvmlFv5NLkcgD4nlax2c/Sgwmqn691rsqPiHCT01bY1kljEl+vBqY2Ur5CTaVA
JwifGwOqfKFZQ31uUx5XxRbMH8to2IwoyeqcjFytvjUdWUa5I07LTW7117tUzfIznikHswu7DtUH
t6AJcstl+8bAuW6dRidDmLBX5IssArNl1mzTFKtm+J6Gtut/zlw+wYNTE3jonNZAaSyMz8etdoCR
XrWppFf0bvFoMzOYvya1zOkGHsaMXygsAGszrNkP3bwXMjVv/rNtundtNedUqjWNSGcdBL1per50
MFjguvkAMU2oACt80B6pWWsDwRLb6Q4RQ4ibteJSoCaiKyj6/AE7hvD6QbNWw0ttHWPyB73B0kVO
ZHjtImQFevwffxjKCtn2Vt6cLB46VapiwjuGnFfGU2sgI4TSo/JdKEb1G3FP/KMMvrtThHn6fyby
PSIovYakybxHRg4iW50im9HOZZgaK8LXgMB4a2HGHNO7fZ5cmmQKCgIVSllezx1n8SSY+XpAZKrg
8+/5acTrLPH7Z/IoySENLXEY5+VizeM7fr0IQZEQdbQjyOkuTyAObbzGpor8eZwvRRDhT1zNPb48
vCMXsAdUYEriX55O6DbGWHeOowrjqTZAhF6cAzuOu+ZHC9kk4dwsqFVswJsKj3bo+X0GWbx782xJ
zV8tCL9n3D6c6GEMkJQOWRxAdY3r9QPlz7ZHiyG6aPrE624M0bFa6Bi7lmiPw2rQADZucHHfInyS
m5759yiyUpv51yC5N4GqnT9kjJtezxdbD+bVVayP+d+jrnxoqB73JVBW7CVptkWuOeb7wPLxOdqL
l+ktGESXk3YZLv2MmfdmCDN6IQXXsY4UqXWz5Z1QPnH8OyhovWxuYMPUu8hDGeruNRf1rBW2Cr0W
WP4IxU70ErHp06h5eQM8QNS8ydKXIdlIftSOSWk4oH3mUpnoW6lSoEoj94ITJq3QZdZQNX1W7GBP
/7zBGSYmn3g7WVUXGL7VpMU4T/mbgK1ejk3Ptcel6Koa7ksNPDcuFheo45/SHov9R/p7Ph5kKVgM
GBp0Au/vGuxiezkpb8TgMwP1JDbTorAil9psJ8KhkiKc7gw6Ha/Nn12vZT3ihx4E8FLkfqONES7G
1EEI41kEPOs3lidzecKT3FYa5miaR5LbWETHRpYB7703a5LY4UwUTeU3LDC6LDiBSUGQ81iCdczf
LoUA8LsZAdGG1wCj3RswFtwINKdSawDgEx5Ir5dqGn/2pHCOvoUBRV7aJ/m4sgsrX1gk/C34WQME
xTGqrB/Yg6S5GWbKheUMPfLdMWMyTIl/Uqj3dKcBZktfGPmQlU29yCzr/deWR9PLQwyBo91EWYt3
GszZhb1rc9q5lWHEMWsGeicGqUI5Hfn4jqNWeA9AlWDnViznZ/iAT6AXKQt9KlkvyJ3cQWYjdYhe
xRpeIyOyLXNsgrtYBFeZHfOJxiuiggvEkLix4BHxMBfDLGDj4JGIn9plIPzjT32yed472T0mSRoV
JJ8ZVZLRhHNN08VVdt76ccPhTqIan8sKlqfLgVYoj5GNTbrcC3wc2ojW2J6LzmLxM5WedkgKClVU
/JR8npsQJhmI5JXzWJcH/Y2nBTihXBKaKZe/s6at7BY0f1UcjLkxCjaY6bysytT856m/B685dE5k
gWWTVODIUcJ8i0szY2/KBT29JvMS+D3s5qqnLuFdvEtnr2vBwv1lJi7YrW/QaimSnTC5iJWhAl5H
PqzzgjD8Og81Gp7GaqIeF5DQia6ckxSLmo1Im5A2XpVQjKQM6O2DG22BNsk3G9JL26akXxtdZ5Rm
jYfXcfBFRa7s0Zea0zBc+GqPtUhWE4VWEO0lUZfdRu2iO+bSm15cIC7u5P7q+etDybyGSwjtqGkO
MEzVw52FxE/kuC85o2IC18AjHnZVbBH5SFGMcvexrckMiNEAJlI4gEchLNktVXQNhER2ImB5FTfN
y5BzSvRv+2PaL7iFku4EDVmbXfLTfDx/kjL0JdtfPa9WPuiXdk4PWpMDpsSdcAQTl+Ve2QyNincZ
C3XAbiPlqyK0sAdXrAjaIE2oKoNZAj/D+eEF6xXdVS3qFcyX9OhN02uP0MsGbS39K9sct9FO/VDW
oLQG28/DIMEs6htEe9jdiroKRjUQ/z6wYVAhC8bQTFvXqeRbB3tzWRzo09XMqxPOURuzuozY3tob
VSZbmJLCBF/uPQiWj7fDYXhR/MDAVi/Yul9U8QRdOWE+xKP/vDSinMWkhZU+VP5qLd3tiW9A0A32
0ppzPKpdqzMa0w9QkikUzfcu+OT72zu2vH5BOBudMGsPTGwwg6Oo1nuDxgGEfkmTV4EdKa0hUbyX
liwLhnowGBMbpOVgAozaWGNRfsY/GPMZWw9AI+OuvWiHtWUOCQA3WIGzFM8/PA/90jfI5PCgtLa1
rOcePfRiPgenrzwbbO51djM9KzYoi3wfNedz9DPgeYm5Y1IGJG+0dAw8zb9t+7my65pth9S+4FVT
06DoAnhobJo2qTH+17BUqJgIN5rdwp+pFQC7lHOZ3x0=
`protect end_protected
