`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 158432)
`protect data_block
wrovcHZ5qwQL2M/nAAAAADeCTRrTnvnNgJT+JPGsdI7teFmN/P4zEkbuE0WrQ72kXRZXgtlCVcrg
pgPNkRH8JyJ64eFxyZFG+Gvrg+AwpIT4i/JTNGatESHbhPFgrp65ISH8Ldm7bRH0OOsqoWlos4H5
N+vZqBOPEQevZ4BJ0EenOFJrHj5iC1IxDYhMUFaADWI//D9ZBITbj5XuXXtwZtPTXHXY8sBBcVBF
phcxbEMmzdLpd0fTdq6nOj+5o1HIvj/yemZeDdCf1+t6UHh4LYl1HgpyQ7htHNVk2V1AYB4o+e1r
cIYSzRgW8w5SN1Fvim6xqnS/0s2SUzCY31tDFg84CsKgd1UDShKUbstD+L5fiw93zWkiXnB+yPc6
7ctpU52oT6MckvjDGod5b5vwu30Gs+yjRJXQulL9JmP4+9nfjLIvRAYL5GdoEYbPMMjheLSSF50O
5LOjqvh5tMJbPgM/+APIUAVzQsi+rq5J+TxYZSvxx3uXBH4HoriKJEbppNXXx2NxNNhMoXX892o/
v+gRir3bHUlLnvXGlAS81i5RKeKb86JL83VTb04UyeIs3tGw3SMpVjoDCuHYjwNrFk5a4EvJZxfL
PxedMn8qNOWsIU1VddOL+zgLaPF+1FfWOXtJWRV5G827tKstQCCbn/SKHQbVKbtk6MGgIlzFwoj8
jd9OQgjd+ISAMnfQfHe2gHHSTsPCXnnihua9gvKKiwm49kGJmnDI1uFdpWLfNyxwccSG4BbbuUr3
wRLCGW9/n9ZMn9FdurdrAZqwzHmL/6b1Q8pBTnT4Rq1BJbyWIlr+2fsksuMKPXIP6GIiyv+RJRYD
ksmNOSk9Jd+r4FCUJayAd0LlnJRoxaxFSAkDCDZGRixk263LKussJ41D/nTG3VRDBANOrrlzNQhx
z/KKZqUd0dPnEVrMjx86MYTn7uT5YY+x47ajxVksdVblL1MZEE4X9WmjzfoaMUL8ZdNi7OuvFK2I
4ISvARYTQLVbcMmbmVLSwd4oJniwgbx5itCrnevSGihWiiz/fpdpGkppW3Q3h38tiY+QtrizMfYL
JFAOJj15S/UpM0qJaPEc4lrCXYUZgMfx9VnheTNRL2XLyrYyhVvBlWXhuFVFWAAEkJfn9RyZ01pA
JQEy1LgftHgr9B8PJuRMochdf6EZmG0vM04AloMub5SOB4LZjdQtAJezuQ3HNXo04V1hRI5jX44Y
fEb2mi8Mux9VZKRxQLm1qSF8OdfjE29dhvJhXyBaztaLmLTFKTcD7KayJv7Lcyy44zMVSl/UDg2s
RV18tUuNBvrg8PuAgwERE1qnypz7fXmYs7yUAAuAWqGEKg6M2NaEX9bhoTAO7Yd+kPTwNfDJPZC/
asmXd3PFSxtxrV2rT8rVDyY7/hXZwCZf66638yVIdJihCB3klH0w6fB6ixYma/lI6/OaOr+wiCQq
2VOgQuF5hZHKUnVy7eWrKOFK8+Ug+NtzIdADozwRGw43LoZZO9wJEGKJQm2Vt/T6t+hdLk/YclS2
pP/T0YDgXYGkslG64s9uGPB+uQqLE8L5KGxCViNBNWDVdAOy2yo+Rnxu2K48Hm6MJxcDzOgCbV4K
3ZNfmFNwBrYokNaINgMRCsUv/Ju29ldJxS3Gmy/K9AT3OCJwKPvqvLEzT/mecYzsvexE7bEZXyvo
yaHcYwsQsY1lhaURxSnzpyeNa33NkLPVcaUTO0M/fu/4qDczPEyxesIURK0bP5WKsqo8EfXCPEIw
NWjpmT9Sn/INiMxcGEAe8aTbOyepdq4nI4HLMj0w8JM4georyA93RpPVzzcaRScm+FofS0eWyV1J
WfA17BBtPhX3aflty87CkEo8U+RikT8G33iKIDf41S+cah/xRd5Uo5Hzjgfb/4bv0zTaKioSrrpM
ZuPZ2b9GPv7lwDjuRbAy5/KRnpYkICLM5oCMWTC95W60q/dNG+X/VQMdW4NDIRmKpm3GNBmKFxKp
lequMEPE/ikW1x5lRa8GEttP1qaUnVWSJlw0J3lUwzvy9QswFkbs0PP+0hZnb+3gehh7epNpQdf1
vYUBHnz47+OjhdQQufHyJ3ZIW5nM9HKdjpnwcHjcZL0KXfqujkeZPpZBCSkrfKt8MAyiC1RFRQck
gtjZc7cUZnLrUPcNo7PTWu3+4w+eR5nmHjssU7qvg+P5juxBrc2Be/Lr7qF8k8lgYP2flgablVIh
SCB87Fnk5H7EKNu59AW4lJxKCps9EsXoWTtgA8WwPPcvWLC8XHbS4xFLDMYqZXH1m0E1OGntsy/T
IrsD9H3YwpANaGWQxzTJGgxgnC5R32/mXNfmJ2DWOSfpcFKQOtWok1IuBF9vlS63DYcpZyhgkNps
7xxGrQ6GMvqFmJRABP7b0b6pmF92SBu8psxrX7L5ghcAl094zNgVTpbDaBV468oqeG1mnDSSplum
Uq6VQ3EoYSPFhrHocDIEsFqq6RNWzDOHvjVKjyejngmoXyUfT31jkprjs+6oIHkbG55OmWYKv0se
SmdVzDmNLu3aLGlj0w6+/M66aTZ5cq2hYfsWUtBiXFJ/Qwp7E/5G+cvIPulz0AFbzonYaRyIoz5F
8E63UQQTCxJYSmNZqNb35Ep+EA3a4+/gKgswZNnYnCq5UpnGnGRavnpgWxMXKHMZwyZGZV0LX8C1
/QJB8zUIkmpfNCsgXkV8U4F30Ua4dEVtYR+d16DtwzZ0vE+zRZRt5+8Gg1xI7PQOpnuSX0DpqeN6
C7T6cqKnQDG16y9wgQrDulAUVVTWglt6JHcqtiV0Ccran8PD1rXPCtKBU86DpC11uFZwTk7q/zVb
germ0eGhjqOOSA6IKshjdY/zb3d9BeJAM4tgqc5SlHWaQDguxaxZ7Hek513Oq5MKhIQoOkrlVFWV
kaDgf4mSBWnCdb71iSXwFTK/iUFAncajX4d9PqddK8HUKym3ybwJXHU5CDxAaczv/40huPLQZhLI
AquydRUF9bKvdignDNDyA7Lfgm7q7jRPcoSq3IPFF44OxbbSjBvtOzHUYOIEvwtOxjYZFLScARX4
j2sowR0a1dx06+zJY05z2I/7zleS+T8dZ6c3Ii8F1MzTIBanNlB4q0YySPsUOP9/6vteYMrrOT+n
tEJnKzvL075aXtC4tZ5Q8ovqpb+iu8wYgKuigdzBs9u+CQ6n/JdOPOo3TZDON9wARbjAtFnzWHWj
8AQWWFAOvPkko7ReHaf1xi3/YAnwSHeJLdnQaAJjWiMDWpB9c3hMC99US2kYP2B2AdahjoJpfYTl
yThZBbnj8aGq0/BOmigld6FTU/667T5l7s35yru+HM2eaMPzejzkqjdPPRbW+7IgFs3yGFooY1pJ
nNGMkUYWR9c+jslPUw/0hEuvyT7tuLVstxxy05zFeMqtgMF+xkFPabl4bvO9qMSZ8UxJQlGtZubW
Ig4yOI//8LWX5Y9a8ALShHEmgQQmHZ9eGgZLkAawEKHyRj5sUkB8AAbv2xLL0GjwaJBH2mtmWobM
AbKGbjkjWYuSHqCoadxaulguEsmXOSZ7itVaTDNTJa4iuEF3K6MFjtrVrix50FQ/bWkw17EUTwZ2
3O/lgaf+3ZIO/iwpnMqhbkO4CpjCRUW9djPIH9gRNIefFoapxbVaRem6THNTkKiNwn2KZ2nOr5Zz
0spYx4tjP9QUsYvmCY3rYmSR9xL0qg/GGmLfa7mGlyC+WRGRSIOfWzfyErryWKgWjVgwiUhV3GJT
jaRwEVnpCsK9OSci+bhgyAqzgIOQ24V1z70ZG3GbVQ07LDxlLzDtNfMd0MrArfUWcGr80RS57FAf
gI1b8ulsNjEbtMzFmiUI1gRmGcHlQTrC7vFbtfSv4kd2LE5GN6wMUO9W+1U//ThMGkbHnYfHbnyd
hAM2dc9NCIb2sts2djvREwL3gZq96phcYsc7a0oTK+RhD0vgAF88pAHBTHkPIP2maRiYrLfLfXsK
qYXOs356IbkA/f5Ia/mVSaYdUiDuG5m0rZIHYnQ5eWyMfsVKO/4TfPgY/FoWIAgiYTSnIApfPzKA
sGWZ4DkLUw/z14lsiyZlxz5T2hF/DFzcVyZUJZ8+mnC9Wy/Jk1ZISkYc170Yyvb04F8DJwsMpstV
2F3J83Pw/eXlD5M0YUZfuVtid87K3FLTr2YZ9AiCebOmfzazRAcaWvFbqRxMF/WbsjqU0Bkn/FXB
xFwjWhGsRRF9c+GVK7rqK6RLETZUqfm/UIXsZbJs2iV2Ad8mJqtzT4atctxSsaqN/W0Jd1p6Aghq
4gC5fEg7BLeAcxeMQ/dWVmbYdIMCHexQbtgy2SAyIh3ZrwOKJc7bDJZon0yIejynYn2c+ZamOs8E
/Ht1lzLY4VizCB53oIXl+DUR87JWK8mH9rhculOl7p2Numt9FSTauUOtD8Ueft2lrY5f0/2xNCqP
BVFwLEOlabmyKItTYVm2i8KvTDc9AzNSb1Uz2ZWzbhrUKqCJKv0cZOrYLSbFt/c1UifqWaWgE3PP
Gc3DkLaDsDgWJIeBnQxxR7e0dF9Ual2E+kuX5eoHglV4HzBPVoVc3VQxFNkNaRw6AEQiK20rN+c7
LJUbRrW6UZC+CTOtWpaJH3s2G32xJNI+YRmw6AHSGooHBDX4wDLeIej2oaOJrUebidnhY92HWHud
rNrnX//F4nbr8Zdc0Wc6pWxNalQxg950jCi3mSV2Pg7thoEIvZvsx6jRyMlFQQWkZxEQZKU5bsVR
+gH1GOkOfcl9cmoOYxunbbMeY69a9wpcBD9iPHl3Hu+1I6gDf/hwp1y1xehCuXz+AIfHndNy6eil
7RVI9LLVluFDjTA0+b1VYOCiT9DHH8E643fBhSEDS26+M6oPO9r36JKocl0ipy4PktScC5S33QbD
DvuKx429iP/SjKYhk8puEihftaWn76UrJY04Oqb2xQdBe6Bb+wiU8GB53qpT6Dy//ONWjjohObJH
N01NTs2WkiC0nMYvj0vyrF67LUuGy4n69QMTbYkdLOYRdti9em1YpwAs367fmkgcKXYiHwQBwBuO
NoQl6D3pT6gNwTyA3BU2UhuQKi4AZxlW72cWgF+Uh846MRiSlTgC8OIgr1+cHO1qsm2AjQqkHF0i
zhxKw7CHuFmsrGcmQ3xO++24MldjhOjEzUxLLaf6mYnnuV9X/bCPN99GgXtmVYPdeHWcKhbEp+K3
+i95ri2HH9gsiA+4UET4MOzFSKJt1+CUbxkJacfw6Td6VGW1WtpoKmMwWzWAfgbc9n7CiCbNACpQ
rSwa+Bt1Xd2gX/Ob8iQ15fKqDlbRnX/75dg6bZpuoqvsqPAfK2C5yA4vrdzoeEAGvgrUjHSzSOWd
LB9JMHc10NVZOqES0wBK+BbAIhMHMtE8qj3kESNnkbf7L7TVRLvoN2ifCJv9AtTl0rot2f83n0Gv
jfRJSGtfLN/lB6v0TS64dlnfW7anyrYNtFAe3gUXxsK9r1uOwZLwetZ8QmrNzNT3YbMzYa2V1gfq
fXH26V0pW584092Oe8roMuKVuHL3YNVKsbc+Pd3Twqx+ehaOAoTQNXT5P97CoXDidTXpUyyjvfZq
Emglws8oByzz7jEBPCVSgJ2DzrAw4xGt0O01Rw99z+8jZDLLngYXQJlqQf6trlQ/UptT5e8CzPw5
2i9fKsMY8KdT/55gIJtClxYBrdS6nhiE3mWUINsGxzZ9SFN6Wkm27AhGwJO8an7mNE3HxmKsF7rj
MSVsKyeaCVS3gEx6qR262il8WtN0uCtVgQU6djxdVqNMaQnodzrneHG3y1Ykk7I9eLbbRxwKhJhB
Etho3Ygipu8/qBDR+uhh9ucPcZzyBTUc+MCz69jxIqRQCv7jvGj77YvHbvg/WoTY8mhVQB0UYHv5
DdkB+Igj5W4mphcoSp2rW3IR9NQZETUC6XXRbre7AHWM8TbqPmtRmW4FdGUHD5x516VaFuM53uXT
EBTxp9eN3Sx2n28izhU9qORUJZlNRgPiuzswx3PJO5Sj9mb7VvGJU6rfGWlrMN6XDnzAfQ80GJJT
lbha3FkChYbxYPNHHWnS5z6AQNfImvh8Dmr2HO3ZxJP9zMOP6kgpagx3VtucawA6jDCa+M99MAiS
5sOC5PXLhc0hYiErN00kV5RwEA43ab5GMXOcAhUbKbVuYunTNRDQT2XjoP6SUpIkMYhtKbzFGuZQ
7AkJI+y/x2GOtFAbXLnaZYxYMECFKBilyVm7H1EkaFF331reGagKklCPmYP/z5nV+k698S7DbPmp
+0bqRIFShgwzMleQ1f3xA7Bf6ZGbr2quRQOyK/SDSEAQv2pgFUGdvql0k7PmtJ54BAp6GXZST5Hw
rho60jqu3g6eKSvaZqBuMXtN7U507KOvUhgOardEMGafTvZFQC4TEhDwsgoMxdZG6aFdJA5Enev9
YcRY2Bw5G7HYCSYdh7wbYekA7Reoa07qgPgEIeuDJlztjBld4WHbbZwSS/WzL7c2A/tRHylYBHh/
dxfhNaYB+JQCibkaSirfxlOXgLdmQxl+06AyiM5W39o52xf+V/9y8EMt8pqyKMrQ85J6W0KtueNG
ebjqtC4jC2JO89MeeY0cggFG/mpTPSYIfx9gggICaoYEA/XpDcOQTUyqywqvMdHlT/uT+UycvALw
/0X6WmQTyCP5L640/p6hRDbr/WpYsZUjzYVDEOow39P01bkZMYlVKItItB4fgZIWtLKAG8ftJEka
FI84lwKL4LKdQ7zqrr+DATYa/Yl9ABu/hcvoBU3PyaOJXmAkm5LGn+i5LOwmZLe8RB0+OfgGl1Xs
+x5LJSLlwtUtS4X4LxVRuP87PU3CIpdEyrLH7ZBVMF2vDE5S8/O+ELv3g/7Ed1GQQQQ+6OJFyJPT
CJ+wyru8rpsfKdMhX/K3fCpD/RqGeCquOeyZkOheky3n7/4hxMF4CDI5hyvkfyf72Tq0jOAQ+iLQ
tinzmcCSap/wU1wCDtVxWukKc48XZUEsA20xnMAmwVmpb/fRcE8XVq24LESCBultReg9fKYe1P8V
Y1ms+ZkUGKardNxDex8tEOcVeWJeiRcP6VqHHPu+QXgI7W00Ci2hoOoFP7vbEJqeldv6SWTvdMm9
iCDoqOf4B3G3GNDRtj72ZLHHwIKJIBJWaWTEx6qubuwKj+HO3Wdi4vEg1k8HdhNGSQ6tgkDeX85n
t7V3j/AsMYrSAzX12niAnMhSMTY5ZDKtiWpt04P0eACw6BOkYVZnj5+bMR2czJqM5noUcpdSmZOE
Y1Vn/sp41e6q5GXE0qrDJl+9ootKzfDD8/8FE9rN98Tclxd8BsWtaOHgrXTYhoLPPgYdxJCyD0C2
mMsA5RZ6TjRmVaYmPAAJfPVCUSZvJMBs/Mbi/2PMYQZZM1zM19IeluuoEKjQYWmdoUndK+3AubfW
py/LHG5Ecz+6tuRK+ORybaCY+UIfyUvzoaUc6h1CzSjA28fL9sfn8pUCTsTPWzDsdK8FlZQWH11G
/K4KSZ7rZ8EZ3g+EB5m91oHPBM+atg4Zw3T37vSSPv2v20FkmBckgTs+8UdgzUIx9QRRbr8GiiXe
V7EQ8lNqWltppjxa1BIEBTUark6qp9y/JoK1ZrgRAW/WWr/35Tct1jPWoz6mfywrBIr0wlkFGrKd
7vEZFEnE+2UWOSTuPzo9BdTzR8vYPbWhmWoq2xW/ME7DCMDMA+Wu9/3Nyc3k0WfeWRQmuxad034Z
RnwJ5Mil9LefdXhASLmF9QyCgOdIIeT1uqfqdy8b/liVmvJMKpduxQI9uCzUCBIrlQbdv/vlWxXe
20bPjnBmEK96SiF21A1P+ev9WEzW0QGcVLFHM0dmkcRkqfJaY780Nd+gbGrFX1s6nwkP6bDb16Cy
sI+cSKPFU3jaAN+7iWsj5r1wYry07nNvdOXq0vFhdksEOJli3c4+dtBRpp/1ZdQMM0v0hXQe4JRW
BHjieNzPftE+CCvX3Sw1AArW+87CSS3yBUf6G8Io7DlGE8YlH0h5B/8wTGjyw2EHqA7//RceCL8J
KJjvRKK6afmeJTLPXjPheQ8M3A693qNxFQaUmcMcvLBzmg+WSX2usmawAJuG92ZKb92QL2jK5ZB6
WVik8IlzdFxEnUAJIJ49/slViIHTRchszchj446gSgNwIk3Y2JYZJ00Fl3iN6NGBskqYp2GQxruW
+kMe3McPpskgHX52M9d4Vlc20LPhopKcNLPBH7+4Y1kG8U6sYP6zZrKd273NOgdosSb9uZyE6D9q
dv+rCSQCQFKCQQeV9KfGDe2iPktZF3i4UGHcqYCXpun71oEQeVdNXGK0vtYt9N9KVWtHP3KYD/ni
/BXev1ig3Ng/GdGz/KJt6cqy0NTnAzHR2gbw2Ha7LqBQfQ+8q/Nb8oVzqK00VEOT1VbVbET8aoRa
TH/kibMymxz5HccbzP7p8EeLjzw86NW7RcLaSXcQCvoeQP2mE6EZ32nDTWq7Z0soa/DyRstgXEVQ
E8o97wdVEg05WtWS213bom3x9fjQ8h3fLhEMNUTmJGz9i27Gq73pRkEOe5CWQThj/oaZk/4ilAzW
bb2qBEWV8cTjG9k++Q9aFi6h5lIZJuXZ9eaTvVYD2Cswr+R3r/76K5Dhaw2nc/OyGZ3xbkvfhV6m
sHeUmIXguJTlUchAjlJSP8U9fe5kvmVY6BLAdspBUtBzy+cpf8tzZvE7teXa6/VwU38rZQRhN2Wa
gjymRPTk2f1uK2NLW1hSpam+ekstjvsa2th8mASkxJJuKqXIxYUkflVcm9S/z5afxH3BhftUIG7D
fnc8gn4Nue4CpE1xbPGu2PVygsy6dP24Km6IWTlf5dYkHhhEoYiMxjIaaKJupK2796KT3ffQI+4v
Idl1WkLxGPPrLyJt9h3uGrjj5UzOQOfxC9XqusTT4v50lMuWkf/EkkfjUMWnGQqIRiBMa5D0KmaL
nr92Sm0dX4TYaAM+J2Ab+IqUWmzr0l27/33nzHqSnVK/XJKJihWpDUmJ4fHqCjlXCCxZ2ogB1ojc
f/p7LemhvOM3MByX+41kYrUm30w3ZFKZwZ9u2ftDoBs0Cs/tyV61GU8U4A78SiWAyvPuxtkOGwmA
ndO7VVsyy7fMrhJ4qHIaylRaAIBfIuwGXiw1WFyYsYhKHNYzBtjjM7xnh1OLnX+xTUWTnA/70s2p
TKYhf/6Igmdl5Jxum7ETUW+0ulzUsh8Vz+lCms2MpnVveOH+shW83zhXYUJqFHFPoiq1xx8eayA+
sLeY8ni754MnxhPrFC58iO9yUbnQhFDvS9bHmGRYmemxHe5zoptujYVwCK5YoAxBa/huhuF8c/2p
CkRnciErfT/gSwOjemw8iTg9VPzjMfVC8HM+EqRzha4kKK9K62LSUvkyQMXMjbI0DM2MA/Nq7r6T
4NGn306ZbD3jo2PoFXmoc+aGyWWApUgd4f5zz62bJj1J+uRWT9syABSM2+pinWuU+JonLgFlBcJw
5UI/+eoZLYJqvhTAJWJI2oxrDpHXJZP8ZsrNVjz1luaw0WVAm5M4H4pitE3MgE358y2CxsbuhQP+
FIhNUln6VgmmDW85+mQCkinR51xftAVvkCXbj7kS0KuLdtGI2Kw7r53NVzWs6TuKk1UMr73XK39T
B0MMZ2jSCNyQI1NakiX/2jPYVSpUOcZXcU7jA50TtfWbLDfYs1Ituj3LXj8edEYYy6IvfVjsd51+
sTNpX/ZXwvEl8zAKMslytfjbXebV08y1mMGpCmO8AG5won3PnXluTeXDhTB8GWDQoSWUFhleMBiX
Q1Yj3yi/e2kqHUsh2dLzAyTT6GH6LipiCWXX2jbzAVcuzxMPs0qftxsgCSYI16kxZN3VOhofkKvI
0Qo6V++Dgo2ZLR244MCGsqKkz2NP/KlVP2NwjAcU5trOU/1KVhVO6upGsjrYRAF7ELsa/BA/Hs4/
RYs2mybSubzQap9ZXdy0hl/nEwNchuVSXBMlFhMNcXLWpqsXrzooVBGGWoLjhHrN0MES81egVt/i
yktLuLh97a5/ohxjoThiskhe6LxTKx8CwUn+klh/2a40A4duOu6zlZTX/Day4dolD0b7HkZotmCo
ic+FljeUTzVChtE05AC70YCJH+EyqQnjbBuLNkbve+9lRQx+CZ+FBYv91SbLoW9wviJhSfKuLM4Z
Ua2FnknQT8yoffCAVRRhsfs4NVbQqywkYUmN3NyoCFLsDPuvNgyMMVL5V1eatXXGA/24rxBi2tra
umtg5pV1DuZ0o/2s1+kETjK6kF/HLWsJhI7Bt1WKrwRWvL20SQUCU8BaNQa4okjrGzrobkMFy5f5
+xB+8CSrsS/EwsafpPLBWEWU2ym+XJ+caCDyGB+E47tgSKrCAdRz6iNufxSxjTsB62XJgb9354kU
JYJ++7YHDMqXX5XdMqOckcmKMSsfYosfYDhBQ2dyvjKagF52Rwbht05B07C7JtXiEW17dLBkdGeb
mUNvaQ9zZN1X0RuabWCOfSC8rkuli+Cb04N+wfy5H5e2NXtHDPYpLvYyXJ7CLiYZdzdmOolwl817
ilb55bh3XhouNOpZIZXeEyBxKJrvtUi0eyBLQsdOTKXXkeNYgXzz4vZgvmmIRNdpAlEhWVCdV8VY
nX6+Nb+/cH1jeQynlAz4KvjNrIfhAqQ5VRTqkfy+nx+TGRDK7GJxsedTO7eD3xu8fszU+4Z2M3qk
lCiqngeIiAlju7sShmEJ1ok07UxFqwGkQRX775wcCfzqUe0IRzOwMNNH6reCm9BS5mnmivk66Q2+
0O4JPblWESBLglmdX9OrUkmalNf8m1EsMFTPjgn4mOhSoseU1G4Nl4GvafsPRNnFEA1ZEAuc9GXe
xgD0Chpi3GLOZNVwk+VXRzoNRkVXl8E1ssZ475eGcvRipNJ2IWf2hOSayAcg5TiOrz+uDCJVqKQ4
gkcKUKqVsm8HuPch2BV9O83JDsIp9oerbCFHSOtdaGDtzGELKtZNJlKopR3S7NhDNvfzhK4qk0SG
RN1k6nIZLOJkO+7XClrMVLIWhmh2syPdiBDFBTTwnJASqg86iolTbB2TeKdNvHfarT7uIuS1JVS0
FnPmxDDOLvNjoAV6gBfKpahVOmUPNK29yzGrNWkEWtzUbq40r0JUAqV2yErMWFqPqdIHel1YJYOQ
nCsInAC4ReRBZ+LpS+HeVE7eQN5Uc7glWMIC0tDHh+gE5xpnThnxPlLhMMjsu12DC1GO+uWe+isx
ejMq4rr2Vley5yqHdRXXKVF8oypkP/IOYThQPWEdLMPcw1SsAd75nUHa96+IAVgPKol3+tFo0RLX
SV8LgmUf6QHqxaIkSQ3c7DfPcyMqKhh0qS1ZFGxCxzaHlgqLVitaphfUlsSKTI6+QRi/nBa3Bl/8
PkLHSrO77pUR/yctp6N2SAEpTJLDkVZlaZYlSxdwuMC4fKfYAgY0E4qKoAQMgzWRQbI74bGdNIkB
INm0WXWA9+PkOVjEAljIp3sTnhPWtBSpdlit//goLUERpwBqJtQrb3yw1xAadze6toiC8ewdLfC/
mQ/HHPJHxwOMP8k0Rp5+LWMCjCEk2aRBqLVayEZIfVd3L9KQgnsws2DG2HDUjIUh3Bf7J87su37x
qLwhuEZJLekX+yp0Mw13UU/IGdFR7GeqHEfAXfcXhk3Q8KWgSah1QWPcWILZwTDgow4W9bccCxVa
ffomSZUwiyGjeQN+vSoj7yJO0dJh9nrCAo37XBCPe5AA/SLFFPwmuvvLVojvNCv4AN14twi0eMCB
MsvPOdlyci+AktwDUayht1br+NKg5eoIi2lIjl476NWBk/+hNffbITjw8u/2Bi6ob8xSyP2lrtr9
prWmHYZExSDA14gRhaZAy5EhfPsHTaJ5Otw//qWbAP0Wu2SBL3jO30HyV+LnVmlm45+OHJy2iP4g
IO9Zaq8CHlM034gz/qbMUxnfbUHQEiNNxGcql48VV66rNCJMlG3Ftfa2PFziXswiS2QYLbdB12yp
IqWMifZYNzkkd5i2t4IUZNVi1opPaqU582bGhuf0xEfEkXITv74KNXDKmO9ZyQhoRotDKzQiWZkK
2NHRxxbwVibBPBXabCG2rjuFSW2RvT/7yxwD3MGe8Fkf7jgKRIb3dpi7eklpkqhUkrdih+6nWkne
PD5NswTbA3Wiqg3jiQJ6iMFS8ypiCmM5bGXBHQLSi2hx6O/AvcPFP/EOxQozSNvWiO1prjD+6ND2
r6eJh7YcrTYM9aqpDlcMJPf3oIrxwQHT9H/eAjaJnMF+9dkK7EoN/mPPqMl6oJXTit3CqDXVotcU
Ux/OrEYORe5rRuYDkgnYBDNpAADKspSx06DqzQqBSFJKYTSkcCO1JF88+kxNsH/tXIflvYSB/xG/
6zR2Abj+xZ7t0cn2GuDhR68pfz0wl6gh5qI8bt9LBCin+j6CgScYLaHKSVSQ6ijDKE0HVaR7PYqp
jzu+9uX7raqYEML2Yfqd/ID7uLtOzTJqaLLO7S/qDk7JNWAFA4v/L2rGJAn1MVHWOFRj+F+0eV9k
Mwytik0IAiDQ2DtYsTrgNMvw9nJQ3EPSTyWP+0VgFuUwq16RxIgJMahZVmtLaU8r2HM7imc3IeEV
/cjikRuo44TwsLp41UnQYSpkzxo2EuK1ctFpaHuGXkn0kpTcAAVnOEgxT15ZjuTMQPb2QOGXYgy3
fQGYUJOWd6ACM6l1oL6m34qfSxAMPzrjIDfX8K9bauEPrNDlLj3P525/oJLzddpAkW2Qc1mDXr6m
AaRtNR3U364IgCmlvMqkzIrEv/HWa+6Y1G9wpDSeI49W5uRs/2c9k25Y+YMQEygdTpgA0rnALn3w
yMEvAMbKtIH727U1WIFKVHuLTHjFI48hD+r84L7Zz7Wf5/8hly7ATdYXHv3JKmIzwVixZoPzxXl5
Jwvks2GX+hl7BgXPb39cbadVUIzv/s9EF9UShS/lPEmP2nc+kzZ/irNg/rvEN1uz8qGhr3ad59VF
eulBcJByXV/sOYPN+/RzEnx3UxOgQG9JZzqyjHGpNPSuVBPZ/u2LFsjisUr4kNd9YxOSDVUtHOIt
0Wca9/xGqdf3Q5IPASUbKoBZvtSUI2ZOzY7vNeouzol7DQ1zqabn4li6Q+2nCKKZne2IO7VSHfgK
sDYfSByGYtcyGw5f2WLEZpGhgqSG8x9I2Qvx15UZQ3fS/BAcnnZpYHu8tH0RX9Yzwd24SnYYl9fv
mvTyyJgm9nq9q4BEG7ljXcaP/2ib/TUEWMe2jC2gPUVkbKnNfiUxbAXnV8/UH+1rxxJJ3cFViF/H
rq1kjEOOHOwOIIdbsZTVVfZtFBOYbdB6R/Z6FwyOOy+5Gsm9LObYbS2r17iD4zvli8pyEv/Iu7U/
IxH6Scb9YVstK1j8PQiRIucTlVcz9/z8U6RMqvaggdbgZEOqXIPQKFLZHXTknDRhTEB4FWaVl3vR
oC8RRgrh1WVhSg0HGCjqNaoKBkhTTiZOEhnLCOy00aULC22T6O/XzsTbCE5v1oL02Q8AtNwXSv4T
h2sVk8UVyxqKXtX6Xgeh/a5DjKf0KBP3pyfeRJuu//32ME90sPfgaqkN65ulQ7o1iU3Bdn0gNUDu
KUZT63LfOUTtvVQA9/8f6NLZ5/mHPR221XZJ5myb/mKur3m1S0pcJ6xSqt8QLVrxyFVjGwISmeFf
AcfgJ4y11R3wfKNyCrtiNWf+NL2HWh3/ykUE3E/ZYvdwd1w7YJU/u/lCvCxwjru8FsnHcKMGI7hw
hGqjIjGCcD7TXIaQvCc1EEOSZl2ly1OLkKc0nLJrT9QgY975On+G87pzLRbxF60vQ5OcZ8rpZYVo
ntUIILxvl1b3o6OMEQN2F2Bbfn317eMS1p/kKxcaCltgKyt9Ac4GosJEIlWKcfI9f+PWHVDc8gK+
LgNUR4tvqZOGIrFpUlBlrbvHV0F2ZQJnXEZ4rjlpqIFJMHVsberMvvpfSK8CrdD/wof9W5DVa3qv
EEvbdNoaLNORzPGadmG19HSn6KXV7MbMnBPhz4TNu1RPTt7Jkurf6TlMyUSOAY1fmKngNlb0PkNC
s05fGSDjPJbGITYYd7/c4auyWgE9CLdLSe7clpStXO7cohBb/HVDtqQ/RfSEqDLFDOaL53tMddu8
NvvTG9ZsGo1ELvD1KGSMXmiCyIBD5e315peT1QvIOekx+7hB8APcoFYYKfG1NHQMls78v1QjgyaZ
qbxY9JABT9xe99OpOBD3vnzW6BrUVmUqXQBIq8xHa9BvCIV0NIgyRX0We6aTN/X/doqQPPLfV4Af
mbdmHKQrMvgYigXQvtB/fPXyG/YCXxUfDstjvjxmbmldtSCBduTM0UF56DPqqybHcuABfz1NHfC1
H5dnEXj8S+8giCo5dbWixuoK+w4wl/buPz5VnDdY3KS25GGp3o2WfE6g1G3CdhuAt734slTbZB9U
Aw6dcAnwGZGGxwzPZSQg1YNPf6RWNKGRFOX5zJ12oeuKeIlRkoht/uBPbq6HjpzyE4O0EhUJB++3
8BbAt+g65Uni8lqI5JBIV9s4o/CqNyr8ESAh1aYL/Srjy6iuGN0O0xb1YFXtLu2YFTYLfWvOANQr
oFu9nVGXYrNUVuydymPMxLpu9qZYSV4RvARuWFXF/O0sT0cAI/H2eiCaZD62Nq6dRqvBK/4ACPWc
G2uXYl0U7O8CQ6EMUVeWPidPrPYG9DYvfTFh5Kdv3GUTvKKX3ejoYWhru1JFA09CNFkFiE4JAhuR
F/y66SMDi6ifFEvBsY7RVJamoUomciitbY1/xbsk5YhsrvBdNc3bqAWJNGznK+cR94F8Yr8Rorcj
N7rWyO8fMZPkjvB2flQglyhZLP5nxRw7ZSZSfLF1WGEvjYwm4HNZRd5tF+cX+6sTuuQn3FRiI1Bu
rxkJYAXAsjASKKioINr3pCixZkRNKaQd6PCaRfEBMf7ohirU1HNz2FenB4BTak8KGXbGHmRAyp2i
PA9wsc0H3YLTtMzBAPLY6r7bf93NEAFI/IFiqpNbqFbypWZAmhYc52epZk4ZLrmHFMzaLh8PfOiA
+dpJCPGma4nnrdMiihyyse/uTQYn3m/8nWl7IKbI8ypROoq9uaRr6ltI+Nuw3jckr196+Wz6PvmG
5ARsSpBaoy08qgMy4ZMUEIkjqNhFQm9d3NKg2sk1bN1gp93VjxWU//UHRoXkTqZS3+kOIubv8qSP
bp2x0vrvfEryPJBHyzJSADKiTgGRupmmylwgJNatOgFMlwVx14D1qjP5LtZAHc2j5F6Hvw4UUReZ
kPSN6j4xfWYAK+9Q6QF5mfI3RKpPU/zST0gxjWBb9JRFpG1k2CRbRsW787715lQUykTTktP3P9s0
gz6e0poXhl4FF1iLlu+b+EZhNeAIPp/N3Z2rSHgoGpKVLErOGrD5FdEriGasb89mEoECPZ57zFbQ
QdDW3v8RuC8PXYUIy7xgmzy9Bx4DZW4PF9N2wOQ/5QAEnAWhFwjHQR+MeLl5xjRIgpOqWugHqXlD
Vsuk7DpcDQlznk9e90FAcfguqHh1u2HyFE2Gsawy7oU1lhY7FRqLwwYQz0ju2VmDZo58hmGZRkUA
ghruIi11loYDuP7+U3f35SZ56hw5+Q7ih2yzYtvNg7IjP+ktmd5xCieCHgWUAivdUgQmINl1WVyw
oPO+IKoPqf+O8uy1xhfU9mHEIh9ZbzUI+2HDl8lcv8AM6tOVDh2jl6SiFn/WMh6W+XXm6LO4Fsr5
lF8GlOgIZTBwGEk7bRMmEj39/6G9El31LRJGwOMNKlJ+1cYEV7U42ttla9uF6BjFneemnprwR1Ec
xlq8hNL6X11DAGurMPyYCXpQ3nCMGHlv9K56Absncjg4+VJJrSwmhWNx9v9lgNIEnlYimAIcRxP5
+OxhTotsoPvNRKJjz3Gb6EW90zcu3DFaDZAdGtjsmE2jv0Y3emSWsXrvkdheMcD4mBUvYPZubVea
HOUcHx2gT3JXkglybgyB75qwCgzHjMR2eUCQkssnTfaAyDC2LJzQWUIdZhXYw+F5cF8mU1ZYlHIC
l10qrt2vmtlsBoRkX4aso8TZ+h630IqdKtJo/K56AM1+WnDifuzLdQ0InImmLwEDvwLdcP2mY2zH
+j1vMHfX2aLiHhzp1RPPukWlZfDOw+pL0i0e7mxT37qNga6ivkSXH3XRoAzj9HJqi2SSO2HRH4yX
3veKhmB41YXSDfnINn7c00amIkb1+4ThC9XqA0wYRYgBL8T9Zd10Zh9fpKooN+S9Pk1CbdlXae00
YpCgeko0eNnLenxD3LfS/XPDkqsTJGqyUxc03ISwzs+dBcv2zSvcF3GMMTDRh4kgUpvRAe/+nFGF
JxKTlhD5dFiunbu++JHYEijyBikwaXIlgKyT1TWEqFx15aWYqQcLftraG+92HlsSYyQbfvYuuqau
ym6dRMuRzd32sdt6Kpld2QRH31OcuICK+Nr20rP//LSSmoi840gJJEaPK3zy1GrU+a0DdsBcfJid
fzxlSEZDM5amBgnTYYcI5yvnSnN7X3KEJamj4jgew5Ay5gxprzJiVo/kTNqA9MSbZ+pf8k982CWS
2RR6B6PdZ7IV+5JKvAF2jbPk+/pz7R5lj4bZgCuJKXiO/gdZqGF1G41vaX5zd8Md48oonOjyIucH
MEOHnUxa8rk9CNv4Zo7ITryIgMBRmZQ91k9dHkYFHfmCeTsTAIUO8yJjJmINAEcfWLjgAvmseTUR
c/cg3EbFxDJ0nIanQMx94AcYg5whMgnY5Ofb5AVCuPIskrLHvkeFGVPWK9WYR7A7KTzxvrmeYqXy
ptR/gF7G9vXz6axO5SQVkK3MMeluLFxr2PDFThKMqr33h3B41sl+FWlAmbkDgnKEYiXVmdF8dyg7
bcAdxxCOV9mIxI+R1HVTRbiUhygGYKWPhcKazgQ6e943FewTlD6K+JyiDrhpBpd52/ppFZ3MyRtb
PMVZ+nKmGYWNqL0jBCA2wM+jMCJPVB4WmDLNVTyeyAhkOp5Dv9WRdxKQrSY36WZuv+8V2PokO0wB
HWy0RaYa3MkPSzqWETU8tyL1FIIfy6bJp95se+1zZ+oJPTolDWhGwoYaZ/b4WyDA3bf2unsv5Krl
MsArbrxvU5J4A9N1jSgj4v5Mllwo3qMe1QJNvAOtOh1lrvEPUBz6xE1tiFMg7W0/rMWDNK0R/81Z
sm1YAAEeNVy0cEu/5GvRAwtVwZo9z//clZYExHSY3fE7q8u4KruMUBtgTbGG5VHLx9oc6oXfUlk+
LmkZySIzI3RdY/QWNfbt268RjqYwi4P2S8vm9Pls3LcB4o23/EvjNZTNFhVRqORHWrqxSriMfRQx
Fok4ErDnu+zMHtW6mDCt0Gg2wiMQtBxj22JYwYTX0653mlus3GJELWvJmfkqc74IKTKd62RAH1eY
ajbzSkUeOfRNfbTyfm0RbhxWV0eKtTMnR2/Avmk+rksU4lWClqNT1NUVdkTAmGuXmh4Kb6aN2iy2
dFqyEOn2tMSMhoC4L/oCgCS+79KPgyIWJTHgcmdjx2Y289LuCQqWKQFqgGEvIJ1h7tR3PuKKR28l
22XxCnVWsOisFBr+w+5M9Sh7PbMNq3TJ0/u2nopSnR+nc2tA50VWmkQw33w1XMW27oZu38L7gy89
9x1g0XE+3eVt8HfIJk9I5M1nKIAFKEPykciQ/qiWasnfc5SZ6Z5EG6hTojzdDju7iN6+TEYGM4Nm
LhLSPdiyS7k9mqVDmVI5wpf28ynx7UFf1+RLNR591R7uWndYn0fsNuvbvinUcv3GGRoawHWmNrwJ
SquHrFQ+6Ne5h4lOqAyZtRU+9X9GsfipgRHyeildm5gJFSxaYsIHDAMcFh1BkiwOozEcWhgwPaAj
1STyLGdzdeymSSAP8LyTT6jRShuPRHSboWA+bNyqCEzklYeg/iuuUDG7Crp2RVmoVYyeajHSyY9s
iUWpXrlxOve297mbtUzlfjoL293tI2MNL0HWa+CajykA1VSEm9tLGvaljsOXCXXGV2Igm4tCifmf
S4dz/L+GXQdco6k/uEZljoDo0qIetfhVlLrKYj3+akuvjIz11U2DuTLaR7Ei7lbFnTaHyvx9Sj2Z
kPw2IPi9nX4BJj+i1WPmvFJHEEcNijqwSM9FoEscfrctYYkXs++54DN3iCtYv1sDx1ZjGgyDcBja
ffiIro5g6slCeL6nMajGIBVaVIuF+7Sq95KTNLfG7a31hfUtVpIcZfPbNXuB8DCfYg35dloZZOZo
g06IR3XO+KwpYZ0YldNysTeZ1ZVXGG9TIyfIoqr+DDMTwLqK+Z3raTbpZU+NjnLKBBy6n9nFApE+
0cd03ZcprD0Ej9kCCP/c6ppDxHb8XM60dUG0YQm8bYLjPBRaxJ5uB81JijyfUQMJ15J5pNFpaGSG
MQo6exykBdKVnYb44THwrYOs2w9zC+t5Hg22xS13sacR3AXc5gerznnrcp6z7CqfQUz45g5U6ms5
tRs/VpXlDUDYVc/vIqMcrgqCs939jdK800K+deP7g3tWyv+ccEVgbQc4YPdmL++cgGGdEVLczimf
FfVKpbkPg8onG2Jhz62MtdSjuhAxApiyEtycD3je0FaAyBcOsDQ0/TfS8X9kejwmGb70omlJpytx
LfYrlib1aLt94vnqxwcWb8Q2TvsJikUdClNdbTN5J7jMPDGCt27WiKzLpQlkSZFQovLVrSXpV74Q
KZCo1acwRHAEWvg+HoKxjFNXKMklZmWHVAJ/2hP9GtFK7YIBbjH4CZ1lPnI/1b7TADpwwtEG6EIH
Lf9nRZTQS2QYI6uTQ7hPkGa29u3v33fbsMy1ljdayCA44fDbY26LE8+XsuC0ngKFFipteo2TEjwn
7wOymrwwhSpgWpWTJjN4CSQCeSs/WR35o62f9XytHkgPZz4KKGAzV30+pLYh2f9zy48YW2K/jWcI
M6FZjPZdPZal55VAzCcaE3Jl+zrIcGtZ7w/S2oup3WJK8mnzycvXhiRBPtsGB2wb5bZaXoOkSqnw
8v/0p9YchN3t/h4x71PycoN3b3DduKeoRH9jr6fqLH3IESWso9Z5pmE6z6keYdK4hWZLKBzGcIjx
NHfdk8XA9Ua50V9V2X5Ropk12FOVxK0SNxwKZTWByKJDIiyV1agIOGaKkNDvaR+6m2uJzg8ulLbL
aBCbqYIFGh3ktJJI8AFjaCQMMg+NSmUnp6M/s3I6r2RZjsIRGCGFUWkGFaEjSy6DtejZmLK4jIQX
/m4DA0cBF94CDC/Ph7J7nC8DV1gHzj5IwTdoUsvPL6G758XjAan5Dc68F373cKgWwuEMN7X/vVA8
be5K9RISHq2B1Xu9pXz5pKtQcXp1E0hJ+uyoArumxGVdqmoQrRBEWeDbLHlj9Mw30X05HHOzs43S
okvp8+RghZk+k11ua15HoY1IPjYZ3jzbFNBkfZNZkfAsPKXP4vAcoof393jamvz+5Cd72aB032tQ
kcQJ1Md4vyT45O88eaDtSCaxCw5H874YucYe41IuUAtZQJLGGihkgC9cMaS084EpwYXqNqkMv2jT
HaVBwmIczTVjvfbZnHWD5nMbbK20esNd1ClcO6yhyhowrtW8crYa462xIRof8/xYd3lVYc0Y53e9
tCyKI09F0wp7DwFai46SNDOzZ60Izy+Z715/jZ2Zws0NcZrjVyFSmOs/wtozyltdzfGFZpvXfeMf
KDi3ed8shzI5Ec8jEJsF/+POTLEkliJ2yQp+yk6l/f65w/J7zjvcRiX1GYHkenSMFAmgDkECLkp6
3feTYwyQhQjslF10pk56apD56Df0wXOhLqQKqd/TMWUT0iUmWlneXuNwXJ/8cVGhIIfVpsYLLMcj
XGaLI5nfPX/WHPovaD4t82CbORvDFfD+/VDA4tKt2xcSXUrKxKkdf6PdfisHbHhiydthi1q9IjMz
nXYSzUmU8TgbLmN3bQEc2imZLXtokkP1T5kh8Hc8QP/PDPxvOeHy5ZhoTIKG6Bvek+tz6GuZpXx5
QyWWgdoXUV70hyY6fbsstRjrSfMHCYcvP3jgMe2tQKl1JiFC3axoX0JtmRn84D/BZjmaRhzW7lFY
kzCODfxPl0pDb+sDDlkY4ysWF3TAbhtwXwyARYn5Bncy2m0NY5zY52wqmB9MmcD58h0b+t3SmC0G
W79crzzREK16V3Jehj5gmtB26ko0Vk/LRBsJZCKuob3ADppGvUkRbFWkS34KEUQ1/QdIlD/sMg5C
zTJzVUeq4W3agx4YTprOi6XQlCz08lnqH/3/EIwqMgDow7azUWQgtBayoW4zlZ1S57Twj3lzcSh5
tpzmCyHHiiZPmASUmwAP9otVCso4x7TG7w/IMIZmVwopZipAGC93CVQK9Upe3iPfSASjxhzRra55
oux0R3KNP6JGW1+3zsUG5zgyKfDY/RY1+gE5dV6Cg3greQIw1BsH9Z/bcW63ufwtebgxwYLVz/4j
E43NXseM41qJmRzWXv27xh3BulUUZIqiR87/sLEBZ+BWAltis71J9bdTPPxibebz/ky3m7uBURSh
LfmrJM2ueXb3kKjPKYRREIPnzCl7ZQVuMXRBkcXtpK7sJ91Takjsj2dZs2Si9YZaXaqtSyGlaGyd
Qnmhrw9uIaVWN0LcY0NUI51Ky67QkW1aGIaPJ4A2R14sGANYxbtKF7RRMVmp+3w5o5q+EU1pcR29
AoEmU+yJjYA5E2BB5fgrXI+beGB6Cxsnq5j6wlFmmFpvslt40fT4/pPSmwZAAmkGXQ280z2GZg3m
53m5ocXNnrMyRm5/jmOeqPAO7CEb6iFMIn4b0VDZ4gDi/xjOjVbrefiGdNcv+LQalRil4R2cKxFi
8iaktRcpTwTLEgtIa2nfUzjVdrF4f9aBun7hImEoWNQcXjReAVTq37Wg1onjR1/F6TmtOGApCGni
8FD/LDluA2dKoaA+9BjJkJ4Iu4yVpr++XSr9c4RU+jxzSNjDph8P7pCoNgD1d/MmqHc9CsnrMneh
jYpCNCxLacVh8/m+nQO9kP6ubh5F/k30awXfspmoOPjUD92lMbxnqu9Hq2S7lJNdoGMNc+6pzuCK
938H1aHYBvlWGREg3GDz+3w1x2Yc9Yh2inGbXVpU+wteDy5yIiOpOL432B5+8HZR6w/H10MLKbtP
gnjuXAi45VvFNcXr5mh1tXRqB7rXbOph+0cliTXbLovT0dHVF4evPWNLmrruU7s4i/J7SQhSN9SC
tBYY5tQndYKX+t3A2dpM5GSN7SkRnUjdg/i+El36IUQE3EM7s4PccwtF+0qZS08Pt/FaYwj/UJvc
3HN7j4QZpL8nC7AwOorsaXIbdHThLzwZBbqBrgIzaPo2O7EISDQpV8t6S3dMUyjDvwK+EQZpDoEV
FJWxSmc+/ZlIyEjS+Z6tbMc4yYwAU+qCbLVHYezNTTSEYLTPIXHNExwsCpPArlOH6j5oM8sstOeK
//2gm82qvecP7Ltq7pMk7tOzq64wlgrAH0cKZ3F4Io5fmpXGYuypl2NCYLYiN9DbF0W3Oar47YgI
MgvaraX2ewO6+vpcnkbm1CeLteBmKea8eNq6WmAORm1avacR8hc4hwaGxG3VCtb+gH/d/6XfvYn+
GoJ21BHyeX1NnllE+VCtGQ57GUy0oKY61NSegJfRZz54fmWctIX8eCk0kd28KbzPTYvtyMh/J2Tz
r9A6D769GW+Ru/JSabsF5YA38GVvoY/ZN43oOYmf9t5aGUXRL3Ue12Kem0fmIJk3sP1dO4z2Y2Ab
lFyZZSJfNkf6l5ayDgOeIpMB9hNiD9DfWGIlllXwBUjCXy/IBemc3NiTzUULSmR4CFElcXlL0Ljd
evfw7Ge4vI5UOd3jmWa4bz17I/raPDfyo4TlJi/MV77Bd0NJTLuN8ihF/4Brxh4gUAvOyeYo+/7q
laKlVKzEodj0ndboyFBiN7p49bNK1+6Vh8dz9cmsshzyA5bRw2qY892eFzPpkQG2X/0fZ6JACz8y
euZEbsi/OzDYYeqZ5Xb71rTwHstBtoE+CgkbwxkNnPgBpKPLN0hES9ELHw7sMAsRqd5GpzqL76t2
pPIKWdV1qKRp2oG9W21UIkrwfbjEm/n4yXmsnnTXsC1zF1L7zqmhukI/1imSfTOKIyx2QeJQA9Qa
UzAoueiSyy2Y8JDsiQnXd/l1G99ETUYb5JkJwf2cxgWFX9kIHA6NW7OSg2gGFQ1MsqMqrnSgaqt6
3BxhdnGuS+2oGJ8hMXOFldx9ipU2pmyDQ0YnMnVsMphwwVXXkL0MqZsaPmWfEa12xn3Lr+vG9n8d
L/YD3drL23TBZaWosGAxPuPYzXjN1tnKpxQGL7u0xJAHNOPacMPgBWxbo/osnFVfAxhBUEj7PdRG
30CLqBRn10UcDPrFFZVsqLOUzxZHdANjWd9ktpBeB8EmYcdKIdA4usHkZlt9TBQICqzTMYWd+Qlr
uiRR0gqDJ4j/E4KdfxwTDpnI13HBT9ywzPZ+taoSH0KFT5hhurMzEtwNYfBBLRk2Gv//CABhaRc1
9G4kBcz0lOUDjfi+qVbBBtkYSwkVVGpEqYc02FEORFKCrJ0dCBkmwMxdB8hnonbdwHTTtQ9pbQvd
8RmetNIkca+2x8sN3ceIavJC5SRRE2nnAbRY8uRS+22GSv0eKc1/83cdZinwHmVDMj29Ts+Z4OJ8
4Ju45UXH7b85pFjCO8+hCI8duNu6tLD1Xz/anZ6KFZRJaoGPlFnIH0LYqiU1APEVFP3cp6icfv9W
qeuPd410R1a9vDEJDIInTDQd2wU1rbeGSGgXYmVkD/hM9ZQAf3VNnMdf/kzupRVmM4cw7XSkHpuW
5yBVwWF6aZ9lnjgUnPwouW6YUQmOtvQr4cnNNWyvRaCDBW6mzeHmqglr830bieh2vQbWCBNeMsc9
PET2djbT1pCa5m79SudpmUCw72NKOSznXxUVqcFf3W8veJ65OaiJ6QGB43cIaoiiYk7M3wo6le+R
skqcj/BEIyhfQf7Nz4y078zsq/4s+oG6U+jRH7ryPlT9rd0Fy+XNt2d+XOfKGGLZY5H8bwXQTDT8
ZD4JzRpbn13LeXALLLUjApRsZ/SEwQvcg0R7KlP4f1yec9uG0Ay1a/VOadC5BkIFbA3TL6aCXNYl
aiVAWpiDpJsDXfJVypbtBj7ajlZy6rx6HCQ9uI6ai1yv4aIvMPPfmMRFvdXz3e2Iip/wAL6Tpaq1
HHb4L0/9RvLsHy/8p83/TfV05fQD+kVYkc2SL8SCvtb1yujp0j5gXDNOF/R72je8T7tubmUibPJr
6tDhXqplyPPvqO8uZylnuXw8jcqmdEuDqGWDL4nzXUSktJHF6n1iTV7vKOnCR8xKYZLZGcqcCi4j
lLVem+CRhS9d9LdHPdLhgxx8J4P2oaqGtfA2iS7pDB/dPucEhkcYPUaXUSLWzqUh9by2XvCpsQvq
3kV7prcx9/SgfZahhc3gkt5PAxqEF92mbsrP4f2V1BK82LyPKfdNRilCwdNOWG7h2Je0G/tfFCB+
vPAQuQJDxs+CHeJ4veviA67z0AilwagtdpfNCOBwjTPY1RcU3fSawf3fZfR97Cv4EJcCRnfZNfoi
e115Og2mGtRYYGjDEZWulg1Pzeb9gbySaRzLzeeHvvDettDYRo/RL+kLRemLdypvPryVgYs/cPFd
5GDxUxpnseD0snpEfYFvv/+kkASlubXSqbJgs3vDu2Zcndqg/oV6JY8UJ/KklMQ8KBLQKxTEdPI9
+VWK9BgUaoFfn2FROMn+KeE02QJDqf1X+yDutXqoCPyRf2D4eLkopeYX4P1WmEiybtHceUUUNnQ6
HL2h7qYshfDJUoprHehnhfVve4hE+16wtbobiSJuK6tYsr4F+cGzcM5rJh8cHMsZ3zU+Tkx6SmfF
gOAqR2TsKknaz1ZDKjVUL7hBZnAa9UdyWfGKL2fap5G/NfzlBoA6XahRx2dbjT2iz5KrHhLZDzG6
KQNzNysAgkpuSidfGAns72+H5GqS7YWBCJYhpcm5v1uON330cF/ZC0p6iP2dYQBL1nR028LgJ60O
CD5+hyax5idn1THqSJrbUHr6eJl/hRe9gH1fWQ7xo2pGxUwSS/7rvB7vJ2bP+y8DDLV3RS7By2Ua
Wn4pSFONQ4LOylyaTLQo1usJjg3D2rlutw/g35QM/9zuSgzmW198MpUnGzf8A6KDy/fI0ljXKZeL
rrIOAbuR3RZE4qc/3exzhTs+vMAWTjfGF7pWGncDKxQ3RE/9H4on3UF+eLv3z4CUIOXpJqny+h0l
KLuc8Ocg/BY1U1TzXCbxhlL7L3mF3Cj2l9zyBu9jIv0A9VZ/VbAw3b4b8sQkS60wtI3tcIBauqt7
3d45J47HzluTmVX0dZi9PIQEC7dytXhdyRV8Xb2owpVrAIykKavgAFxdsGnP21yi6aCWAbPRLmVA
Mv5fFyQeFERNl+hV03W79/gIGjXVU1Ztds7BTVZsitx2pYMqgM/HAEWgZ5OiM3Uj5g95dHygRGCK
j8OWghUlzBf3szAhrFXimss4p5SM6tVQWNDGS9rUweiYhTnnY1S3+SdmYrLp9MX5jpikGtU9EG7K
OcxcRt5cr/RCYMHOtDl8wxZ/BMr9tFQmVPfZ6L1vVhKMB+6qDngUt3kPYiK/tGZD1ec0eD8WfI9b
PP/I7G1azjnNCgbFph9EgH/DjxrOB7rdcvj0Bjdap4Z2DGzwPv6IYx6vJfo17MRHamaffeViateI
T0pQIBkP6hLNLaL3IAId/jud+sf7s+LrLmzbfqFpbbprq1zfgploFseEl+OsXRMKUEW0j/C0+ycw
ZvHhUjqDXMgHSjfIhhtCa71EeYnu0vmzTYyREqK2baGCQlOYnkuk/4j0QqvrQNx/x85f9KokmrCD
4XMc31RyfHCKCcb9iuL7gpRZxmuPz7oL1XMNfNrc2e4wIxQSH0bpvyJBIo2GIX0YZ4HWM9kNUyTZ
84f1h0OZKODec7m9XXTNPiwI3lWvhDn61WVs1i6rC0tJv4wMf70oPFFqT6eSDNXGElf1zgiA+Xn0
FLLbrJNdQrnzMjl+0Hq4c2GjvCVUKwXxCW2Gt51T7im0OYade90zCQuynklQehf5+lRM9Bt1+i8p
sF88hIL/Mpp0Ul+emuBB6DqAWZpqfmsvJ1H5/u04PpVhEJ7Z8tgnbhg0pcby8qwOu0LSQ1Z0VvX2
9kl/EvSLJhgIkIUaMaHHILRXd6pP/ycKH6ONaLMfNsWmoCLCLXsS0LY23IOH98K6lDdn/vpm4JJh
tyj2cvbV/IFFUulQaaftA3Vd6dGl42np6mPHcnq7bYdTX/FNI5nYU+6NLZMXCJLRtNcdATnwmtQR
/oNRfrc009SO6IA8aTroQvAWq8Hh9VIuWf4n/MMV5KnApOrzsd7NdR13dVjS828zSRMYA00LVPIX
mzX0LL3qLcK0/eMESbG13WYX8c/ONtoh3BegPv545VQ08Oi4qyrDErO/8ocNfPgNJqfgwwwZstV4
mSLR/B8CkDzogHDHqk9VrTcpCFTDHPss5WHe7Pd1Pl0PkcOxGp4pqWakkRXWebDSgAkU9mRk0UkV
QvZXbEQ2DDldlDUvBksZfl/Vv8U9CDoqz6o/m3h7puT45hLu7D7nFiVM3lBOMcyHG9VU/aRjPXsL
J+lPrDrRmKi95Ln/uKvZZYdn7l/U9BCuRgl2NUlUrn/qqe4XyqZhXTeSb3EEdvbM0gQSusLmyQp6
3W/kQox/QVaNoOR7dF8ikvMhfaXHl4FEvNho3VR7R+Mihvg8Xy/+5T/ejydioyW4yI341gE11yAD
DWFGdALLTLKlv2XfyNFuMPB5ER1oFccI/FL50sS3hhYhJ1XqzBSSOVxWOlobClmLBW7zjd1bb1Hl
In/Sngg7kfpvKQ9DNWqe9b8FMRh+LPgjkyF0+D7DiwKfojcy/SgTkywWwBnrEJAp4kVHIu2i5pkV
hiGP3FfOXrVoBlOesMExNuJ/7ysiWi5xol7lnSFMttHjn1uYw8Clzc1ucswTuCMYw58fTasD1Sa7
YqaxxOXobCgpl/3rVzkhnkqm/tJGkZxdyiALxhwdqpjCBwxzHlI7Av8EFiTa1ZA184jJCGh2gc+x
pJuhaKwrV10GmRYyex2g1jjpUOom3RPB/K3nLk57Yg5g0ZEJGDM1f9qkLrnhEmmQQnEdlD2ilS8B
PPRs3k7OgS3rFrK0UeLjaeK2+l4doSXHTD3guwGlrPbpXaHpoQ1BWWPAlnCqjurEzfo45D9Uyhs1
EU4o+RzPU8kk2WE7EeDKkPMK2Yb/tabIw8MK+gYscQZGLxuyi6duJCx/EPKp5aRzyKJakfyVlDb0
+iIk4hEvqKXTu+2yycaEKFX+WpTQykv5pjs7iQWj6mqDgc/ufDG5WGrVBHHPyyz0olVfNH26oDTa
heVZJV1O0Om8ECoKjUhbPhpD176EfiFZ+7XLVuAvMCSza44rVa9ytYzcBYyaarg11sDalv+K0Ejd
r5Ho2SR4XVmnjoqFb7RbgnOq7EM1X+UURhBsFmlWR05h0vjpnxV6mhe70CtN+r/SCwckhKyHJS88
wC9YTLgWcyww5MvwFp7d4IgRTtWiuVKyzsOKebtheDha5vS8fk3cwfIZsXEERf0WmZIE4A6E6TRx
ffsIBL0z+iCNQa6ReJ4a0DNpH3vcQE2ivxmwpji7VFhVZBA7eVgc1eCPNPTKSCh8B4Y8R1ddyuOU
S3gfNb6T4HcC9jvSza9Mx4mNOH2Y+NsaGVqrr4BZUpV9XPU5KQrwZG+hLuZbjO0H/RbUUGZV0sLP
rBqOWriADixpeYevdHTA+9tMZnROK020ORq2oBmiCH0nlDQ18thWXE4LlAOfQEHE7VR2j38pblVW
txdVZcnWBLRMFm8/lJPNgxR7a7px8gdz1Xcg9NmuHPlNPyfa3Cby53d1tetNuwGyguML/lgljcap
TgEnbNJ/TD8siSkYDDA4euEHFj0DtSAvQdCx7ZbsOLO+n20akclQjF78lg3zHj2dGAhnIzki3qse
p4eIdrM3QwilJR9h0U2AtEgSFO6eK8dN9iOz2sL+sEQoWuIordV7qkW97o7bvqIBlJSqM1FettKG
ZlFR/F1gCbqvM25wkW+XS2bP6KJg/6fMAUUCqUs1bF/tgo3iXSBIAh1QJUZDGUe/GjFRggVx/NxQ
0eUUfIRG9m0HehTaLM7e60UZreEw3rxgmYwYRtAcb0CXa7llX7NmYYJ0GvBv9zj+91eAw5DIDjAL
QQE3sETP/Zk4C03UKbY6nvpLvVwsoDtmMp4wx3TeyJTF9t6CwUjUOt55lfV/3x9PHu+LPT4XXMnU
CHIn6fZ1CyVhVP58jUr0N79jteJARjH8b5K+PvgL2LgS8gSZGY7G9lmeJdusXDQ3AVhog3Oybfh0
NY7hJuulvLqdSV5QJmJnJPLcGwT9fadhIFZvD61r8Ami6W1Gry9VJHetp+o1EsLQNq4sqvE99VzX
hKxta+fczozIn28swkEGyz3RZc32jOR82pzXDJ8YowdYvtUJgUAc1tE+grusD+S5OAUdgH0psQ2S
r3Efu8YiHaXpOYNLOKuhThL7Zi/igkTRpyANAjInbZFheH04UQ0qT5jNwGzyllblFR7cQvYr5qcf
eGDBDVzL6F0LWPXY2DVRq0QDTmN1tJ3hiKhEuCBowqHKZBqISFoUIerg6PYR3aYIH5XzZmtM213B
/wZ28vVQmgv2zIRgtBWDrQbXPoU6eQgiGiuj/Igrl5B6Rm+9yUu99dwyv5yh7jG5D8jyXuSu5zI9
qxue48L0klclTEq/qh6Sldgj9FPIqxIBucWzG3c9haDb6TGTPdig2HDBFvk3JPXIY4dTK79Br5Fs
F/q7lVhTe0tTVrC33foWBxBESOKtIrNCkU+tTx1PomBaDqfjBZY5oyTHWhDcjBktBpugiYX4xsex
T5CMVbrD/rlBnqZhNSkp6O8f+fg1dwmdjCgUS6YDvkMm54GQMspl1E8ekOBsyFiw3xkUCsowr6XD
SjTYS1WD0Mtw0xDjXEP3h8AIuUML83TCFRZKBO+QpYMCu0pw1C9H1XqX87sv02rZxuddTnaFOLVa
ep0bDwCvrBXWCdpKrYL6llOpjIu/Dz8FLe28Dj0LmDI++NnNG84RbYUhJ1P2VIIODYDhegDKfaDM
2gPiCWk9j3VUD2lSr1I9APbThefMM6rZd0waaYflikQCU76Stw0yG1MdIpuZSTgtazXNJTkw1KSi
2BP1eBox1VOhQSNdqAthTdbv+gjxNcJ4xl+NliBhDJwyZNurfL7vm4htRjIvTNrlaxEmPwQ3PxDU
t7Un27mZhJCyAV7EbAd9IGeZXGT5RHRhp3h8Ve3WyZIfKV4z+VUQsixSrTzdoEhgsrgizcEbvioW
Rreo7HftKimP8sMXURkCB0szpKiJrAqxr/AmSaBfOWOeiR/EmXlMblPLWp0WYXBTkev93blFNgH1
SpNSV1Calm5J4tsiSNWJa9lBzbnfpJPP5x6bdVsJcGikwkz5KkEe5Fu3yWvX616e9jNeb7ssLnm9
5vRevTtrC1dK76cdZ5DSwwDS1Ct6syqLfAo4lVs8vVSAit7DyL5dKoYrAHh2N7RpaQOQdAu/bp3D
8jgx6Otf0CmDLTp/jgxLTJm9RVZ0i8UHhlx4+w0Z1DVdy8A8qrqWegJoYcbwE3dfa88yJsxJjDcY
c+VMKw9n/RNfLQL3R0kADypQmTZXvptoAMsNkaMgnrab8uEbKHtuWoBVL7ypESPeRrhTcx3JS6QE
FD91HSE75vI8uzh/e23tM9D7HHqwyfEro8h7KJvLH4/GItDLyzp55MiUTWxZSrfdA+YcILW3JFGh
wsWP3r/zKtEVhd7+C37iixp9UQ59kBMmRB3nbVEhqN+5YCG6TTAfFzJKxXv5cmN/uApejZyCT11q
TKQZbFW615P0Ig+91f/bDL/bnb/R/GUHncfwEBgHyiGGqFht7JLJp6GcqNIdjGW9Ylh/rVgMiuJr
IQhk6kuDSarqciK3ceiKK6Ra5Xg74UqcEo4IGaC4ohZbuV9JDExcpn7Ke05ZbAPLaEE28wok+hr+
ISZQBsqQ+jaeRX/Q3EPv5O0QSGYo1+OgCUIC3BjgT1NeT5tcuQUK4qWJjVOEtjmX7Ok2wVvJVQln
KajkdwwUl5jr3vNd++BY5tmNlmnJRT6FeLxgucuUigBJLFm2MeKkPcOtCKMhWw7JSG8w6RbJUmcn
MY4KXQZX8EY989DZXhVigw1lFQM/soGmM6sD5ShQ9CtJurneouzLKGHUYl1h7bTxAMID8IieNlUJ
/6t+8diXQQMCjxkZSbXAWqsS1iGvRS05tIFg74vsAvpL4vOZ8L6reBkWFUuDIMv2rYl23IwFbDxF
/C7pdzsqCGtLl/WDfBziIW67Vmf6ss91lkNpcDIFDa759UJsZza+6n+J2YaZjAfDEMFv9NnhVHgp
gLxG59KoFK0eM4mfx9/QZ8d9v/nT7O9542XGjmJWlbbkXZzWe00NbrrRLuONAVBN3MVpTvnspffH
Lc+wwePQmV7xM3e58DYInuEMLqfTJnl+f5zKPEYu54o5mu2s8C7FDrFMtMmOvJ1kdwshtLXQGGR9
LhcR/Z6KCDQZrcMh0icr7sKpdjlHmpQ71V19A9xUjq0d3HakTZngA4+tip8iI7ldX8Z1q6NAzOVo
AqdGETAg7cQfHHCdelhrrxjsgVg0ieLiFpMJ6unIiDn9kTHWk4/zGa/rvOnYdXQ5ULKDpAxEPOnf
D3RcV8eTiyWEvo8A/+OJLmlNJmL0AJ+8XIcQ1n+bEb/OIN31zSrWg06Il/QlRkOHB1ZSbzvg0QVa
dF2F972uh2s2JbYAIolWYfi8PRq/b61iyeLMFwBPPkwlIAduGTqwEvDCDZuuBXDLEeJYpBqUeqIu
eRhurdg284b7GVQ7TCT/7eeo1emFBC8DSacq/AQTw8UcZDt/wvC0qBcswNICXa05e/KMYpT5YcKD
k9gTbcbn6Z/jp5Bve2v8v6ixFh8m9J3m01SfLFosUqn0jD5txiMwuTMzGFoWF0U06oj+aXTsh+Qk
N5xIP+ndzK4GDmdPdrhL3ibpnWFRaef4Y2aLY74tgk0X65LVBcpx1RhwpuVXQIp7ufxCQGTNsmri
rjOEjEInAoBekJCeAX5QoYJTbRwA7s81tvBnCe2RB6d4z2M4N6NLdMNLQncI7x2OVt1bEBFJo9nj
sQo9J4AFkw+YmBwfKO6sC00je5viVN4Tbj+DxqHJBg7JRTtRAkYgB6nyBVbXsmAiA4JIVAirCHWq
QzMIVFy1gLGSRYkLVSTIi5VFaKmWQ1FAKoXa7H1qAORxUy6CSUw1ERHdtqOTEhWbeggaLdWqyaTc
frtxghufI9BP+BFdaS7SxkdTx67tmduRDG36TNMNjjcFyBVKowOaiY/B2v+hjSRO/ivyj5CD1+9X
+x5aFiz5VUExBQ/GuqpObvduSTFUczeLdfhkcOTdux+vj7KITIVq3dJo/QAwwEXX8lbXFwNn91Ev
n32BdNmKoJvsNMqQGH4zhQDiY36ymV3q6uQiCQObbEO1w049LkA9XXVCCd7zKIirmNNauKBIMUMB
+P5GTp8fh7s552lkLlHmg/yCe+TvZQZV+iAEPWnraweozd/bgCKsD/6E3st0YX/tWluHhWUgP0lL
KV44JjqfQiEP5i6xD5cN7cg7E8O88/R+tHwllHt8UMvph+jM/4/xgvrLDH7wn0E9ydzehDW3umuW
ND/UAuJeAil1JC9r+HD98TgFhi9AWusotGCUZwvZv62sY2NIFSIh6sjcyc4Imk8HOUXLqorUQU2P
IzQNZ1iDWWjUKV3Ft8xRImyfNf+luc0b2y/ugXzSYUHV1gTQWYU3x676bP9Su7HUCteBKaEWodM5
DA6qd8IcMj572tSL4ILsBgWPsuPAwutnwlcd72f9b215ylzsppQBkV96RkzUS1rPw8HYBXkyTJ9m
3dGk1S0+QHfhkYrNyHMOEx8mGSc0h1ERXlYZEfl+j6OHNbRAvc4PXkRLiXpkg02MCYDF50n/3cZc
vvr9WGMvSskr68AWtvog4896WE5NnMWBZgDyfWjK6jlBfJqHrOLheJp+oNDzobYJePVy7emc8sU7
uIcCkO9QqViLUf69jnRgBneQQJF4nwQ26CNi44hR6Eym+0om0X9gPH/UVUK220TeIqj0v4v5b+xF
+WAOeRLE5b3wCPLM+yBqh9C7hvTcR79oI3Fkdg240VzBS05Bo5uTCLJozJ7DkiqfAq2Zzic35XUn
za/l8Hhbwzyo//q2Vdh9NV4hweRu4qU8know0sIX7bN/8WXk2kpwcTwYzxz1M51AOwK956UHizG6
JOXYQlF3VWWhE5vaDDe8Em9b2wY6hez45jDB4AhSZikilE/RI1G2gLw8WZGoFSMscAx+1cqhfaCa
1Uwl7FPlAazLQvYTHug34N4TIOVsMZSwlTyDnWubMI2WNXXyNL4zXoUg/7RjCfrUNEBcx9Xxonwk
X/Tl5LyyCdqcLpT2kzDPbOfS4E5ainZTY4kMU9kb3QI4M8zoEHBwqkI26lV+W4fYcUuBnVR98rdd
0f14e+d/QiT0lYOQQ57y+IiO+xmu5TEZw/J3bQIuwsFqHH7iEM3ANp/qph8lFysoExh6N+xMrzCp
c1z1kPfysGKlEjPqy5H9dJK1kp2d2Jqouc80T4eJsatbSeEb8JHatQ5RcAS7NjxfvqEy9MFRdVVS
Sw0SK55fzI62leZm/hgaAVelLkfzWK+MyzBRuU7mZpbvvxd2kA1VTyIpNyeVRvpzREg3kAKniKpy
7T+KF3ABA1Ft6KDOuvh/RTVMwZWFyBXeY3k3JTeCuL3BTiXdf4znYRTY2yQPRdrQmSNAVlF8qrXU
TPsSA5BF1kiRkBcW4QJBMlg22H5vTFLgMQ8gER7JIAt/+UimbidzcrR7QBmoReUo4ohEkcijyOCr
B/e5P2YMV325iWLICREgPJOTDO7LGTNs+hDP7FeBEZ7sgfUL64B9pORfJ0crc+5MuddfLbekcJx/
fnyINNl3VyO03MeXr12D2/nlSX9nnPkdjxRkBgF5K7WHDHmIctH0BTW5JYqB2rbgFJLI2Bwl5EWc
LI5JVRBh/iAGSmxZe1Avrzf1vAoopV2sSMKQ712CMENoWGQRiu8RZWdSGIf0vzlyFclc4Fipx2E5
gvTJQQ05d0SMXwfqg+k+MbWh++dCoVhZwfHsFzOsHXBbebb4g9rsJBsrnxYGxuqaifnNXHxpQbS1
ysufaDCsgD/zZx4LSpWtlJK+vRQpTAJer1rgaticjbVUFJXyJp3O4JCBcacJAjJmpbZo970JuDtn
Z9M04BWAPeK57e1ZlhfODXirj/Q1c+aoQLPa+ShJYh7dPGfreDxBjvAq4kq+8jQRTHBNX7f2ACIK
mAF/5CQLOsMWXeiEcsgOMij05jcLtOCAaK2uG6Rf0SZ827/9gmXJM3yR1hT3yYVHFpO8DlzoKKT1
3F3MSn/5zEm2M2a2eHFcpsz/au18QgqQIrUPb0VlcenpR7jCyLooMpIIWGiT+YJzQQ18lWKPd9Oz
DAhGPFLwRcp6F+TZZZc7B3xlSc8w8O5jEYEsqUb51AoHKnokUYYe9JF7/jvNfvxG2c3mlJulSmZ0
gZ+0IE2G5GHF6G7EuMZemEUAIa9n/0fpWhzzI4vDQ0yFzbnW9yaKsC7S2ZPmD77yGWWMOIzplsMn
eUBXZbwOn8Wd/zsYI6sTCkB0v3drMmKWDksUEnuFQ4royFW332MO5m69kTri+jba7fKth/33QlGh
Cefiz7Y7W65a8yfomI3BJXALTW7lek4eb4MNGK0ctuuKvUQtsrHuog3l0D7F86ACgvjN1C8o95jp
9XDg6LtdnMWSJJS+bCaWAy2UL41K6VTvn2DFabBJL75aPzdfSpmDPB3es3t4owSzvo1au3B8Ngz1
WoRAhvs9frkTl7b63MThOlt77R5VUdRWqcLRyqYAB4vaU76zDTvD5oULPjIDtffgKEJkFIjwUX7m
afzRYWjTq+5YGhF/w5+qVvdFyjPGxsyOfggQ96PXhs3HRHwRqCCnwQxeCWqvPboEfvVAqfJDHT7j
Gr7QdBtcW6FrlDEWC4HUXX+DJBwOYAaJJiWXngP5DAs17J4wWBIAudkqjQPB9/Y0uE+CC/pKrEJ4
DfA1cp0lYWSI+yyFJzUCWQD44TehdnEt9GZZk6wrRgKr2wVa7sRmw8smCjqYdbRxjtQSXD2RS/W+
NYBJ4C1rusn3DzSoUSo55HZKoklkncBuHQtXXHtm/DuU1SvwXZRSabP062Rexe6cFex0il3d+COD
3OxAS+Loj5cWlqychIPSqZlEDn28xS0gi6U2+Wb8M7+X4XA2WK9V7Ecn0iWnJkEdX9rqC7oKs3+Y
exZ5nJC2UpUo+qt219Cw3lAlPQH4pfJPHQZhrR1cqMAr/bXUrINjw1+aXcer1wplhXHGxYMMr0eb
qSd7DtN8+LqtNbZaOxfT84I6be0SHfB+KiNpu8IL8pUhKS4RIlhqvhCOy/e6bFmhaOEWENiij8uD
9mNdZiq7QIMv4UC3e/bI9Y6OtWN0Z/Gbk1TxNqNpj8+S4FrIUJWPWcJ3TfQI0tl0IO1APOVcdr2T
eaT+WuwvYSc/NwAxQd4ibRciwPa7noS363Wb9TNv7kk0vjVaIC2Sg0704Ic3zdWFr+D2cML1maUN
C8lWBhabJnAFLzJOEr8IgQcQa/BpZi5PAHSGh94RujKJXhcd8Wm30v2v9Tfklt+Pp3BS/AChqhez
+l9mNTkpIaVuIdJFAB/gXnbeF2rbMIBYtvVjFJLzWl8U6pN7qZXI7SxUmfdo/+CTbthIAjbfPLZH
d4kZ2yNUG5ilrngw1E7BWzkfti8LgnYhSvfSgsTy4DRAE6khRMdIZnCD6lxBxoQ1n2PiiytPam5Y
ngk8L9O113j/fhGemAraHZhmv+mfqQXCYoROTmTDzNST4dsaBAIi5XeYUCOXTCDUTfK4xmYnIJh5
0qobPMbGekT03cJfD+sG0k5XygIDfHDG4ZLzJNkvLBjEVT8GlXNrvA0GwpiiaxvZkxnejL+nYMPV
/aaqs5Yreb97+7AHiaJXpfdneajFT0X/gHjhg2q7+PchE2Wm2WIwz1XHl/J1c/4fpwv3xOWcW4hz
AHxdn2nKgVkV59w8sLr33RkkE18yB2gvvmYibYCaczaMdJo5zJKZgy1RJRpg2lgSypQD1KetFIsJ
SC686i4qKMxFPaoApKScAfRQcnhV/ljWlSQzbsQZyUszVDWryZ28YOaK4xF/wGmoY1IwaTaH2vb7
GG6SFOE1O3i76SmcjrqJMyXjbwUxyhzLfZCzV3mxNysZ0eKvRB5MQ38SK0alM9cLwD6CmFBCpniE
Yc4ZkoNxM5ZMrDyPjtWc+9U7++KBKX0F2/CUKb7uUF2LuGhXvz+co+ossTh7kE1cjhmlqMJxRO64
R+pdb8z4mGeRT2EyJXjyFuqRMmOB9R3bxhPtzK/0eOQToc2MaRbBhAEm1Wv1xK6dnn/JkcVP1G+y
Tp0rnMOD0yup+eALed4IOjwR6w6btJ3DjO58pqk3VU276JZtvVlHAWWBUEsQ6xT6BLpbgO3SbMxr
6X1IaZSYn+ZViAvQlCNwK1A/sD+3fTgtCi1g0WZT+WEh24b/Mf2e9+IFa7AVYnCUJQumNY0wED3j
/jmd8L5f+GymWkewApj4ECF3JXXc/zOxLmiX8ADqUqmrrcFcnxK1YS0zG6xT9buchUNCboaeNKZd
6JVfqnRboT8I3QHljpTzlfsPiVArHXlIdwbWFUDSEDYCcnYqA71QqLJVACNDLG72ZK+STlReTYAi
36kIor1HQyynU6oWPbP6WfwMYXddxeg09XU/bHnOPZgdki4xtoAm478nIdsg5ien451NtdNBA1fd
8CpxdiE6PAlV7GOoXNtp8MaBLJSoxtUPgdQmx3MFa/AWqdF5arFMLJcqhbwlnhENRdvBQnVqaudG
CPGEpBYunD0mtg3CyxcCexFYCILsQgPIpY8fIJL6jxS0ukDklCXnm2u9Xm2oimYDCP2APLKiD/o+
de1hKjODoWiXL/wuaEVde50oAv8J+xMaRU+F4QrHs56VRrCdafZDNXcosYHEbQ9s69Hm1FFFXXsJ
0HDPYSkFbC4BT0FplzWKLdjIubAY2ch58IBVwUqdXC8zBDaG/Rm1UDpqh6o6oN4CZ8aSbcksQGY4
Ume19HcycDqRjYmcTt44mc2tJykTG66EA1eYh1F9KSg9HKfezkugHQoKcCnT/4kFIOoyQupWfpWG
SS3iG5elkAAWuyJ8PUNGGi0ooJNKRGq/GF/muQNWKKcVY+ApX0UnOSFGlNzc0Cm21p0vuB6oaGmT
fSFWOedkh+Rm/pZ5XefK2IRB9kV2wzttotJ261y5wNB51yJCJYzufeQRUsWEcRh59ISjj2ONnwJE
ehr9+UrTKpOE37Y6SpPxsiCGYLlPkP+OaSRuF0juFOLahUev/Ijwb8Gdx4HRxd6apgMdiZRrhI0M
7Ou9er9ge9RVpO43oTQPVFMP3bkklTby0lTFWH9sISqKtwFMvXWS1CkL00dShgxFaPwzUNiB4t+z
P9aoL7CQQuYPBvSPTQ2AuPOYPekioxgT+MRWrzg8nwPklPtlKtmX1GsreNd3SJgKWMu/f8hO8Geq
a6+9ZGxD+KqAwcwwWwleUWVVL11mq0TdKszS9a0AmSwJpHOQ2TQ0eO8XI9rD4K3VZIhCV6PsQFqs
4WiIOwPut1hryFJHNMVjQVLkYU0LbJsRkdwbTu7IpzYtu71AXmxgVdoW+zCkCEFexYtuBHP40/XF
VSVyMVkQxNrtcTFD2AEQCipZkqE8KxthJ533uwYqeQxAOE2xYK2nPg0PePoNBNKw/68iXs5E4pPd
ckTCthwpMYCzad9RZuZZajUvnPZo11ojLaiNO+t7h3TOMaFAAgAQYN+QhNkBz8pkBXVpZV2F20cH
apWI/CiCecADTZ3DrBrkpus0MYqCWgEWUQ/M55AKFaRyvTxfgkPhDtVZ/EBydQdjEIViQAb6Q3m3
HmGFvMRKx5PfzTM0rRnMHQgAFefxfrL4pUAh0g4RZG8k2BcRe8EsPjgCdtOtekAhReHoxZjgNkpg
KYh+F/G4ujKx97MOAJIJcpg2n/49hM3wvi4ndG9BM9CobzVhzsSt8z/ZZdrjei6fmnZCS0teZmPf
cC6KRGXttpZkiat5ww3A2saR5u0AokH5gWv4IXX2406SPp0lL9/cdf6xzFtiHSnLPKQefsFBludd
laWQmlJapU4ZlJ8LF3CphxclK0CLZgN8rjE6oBXpbHj6ohy7MyWrLWWj9gUaslDx9FSkH9DJAh1o
BeMEvOAu3JP/ZQ8TMZDp/EoSiotYiUJBNnWALjVfzrCY0hOHMlSpgGzZjlVPa0nhN+58IDPsz7Dg
5L7ce7Wp9OtffGtJ0c/f8l5hova6MkDavBtzkxHcuuLZmbKtyFpjfRNyRtBFPjtjaKrtl4rBl683
huxNv65tMXKeNXTlKVt4eZyiHQiuugzyobvDugbshXTmsDg0Dwlee5H8BpyGivkKijMo//LVHsts
/puMLq5FeFgmpYYiuVkt2F0MGgpMpMjERa0ZquToHHmb5Qt8YsbwLPO/hyM1Q2dE8E/HuG9cH+ER
KvVkiyFlerjAelYMBKeIz4RY0oUbYHKPqf3Dc6O/Bb0ep/a7Qae3S4LQTdHIfGWiSTqcnzX9Kzee
kMDtN9BVg6Ue2k/dokHMSxaTMv9Pd1hQvvx3kbQAq09NVk0YkJMzt8Yag2/gJymIghNuPwwaeS1u
eH2lXSiUv6GFBukV8c1ZBm6EFEt76P5m7Q5yY1/5pctz2yfKk1lhjpFGvJNbXqic7z1KgUd/8uVM
k09yImkR0Op5kNyVnO6lasxDzYe13+GTB+WxVrCkdZlasdmGKwoI1TtoEpYONAaxOBbUq0YzS+cn
B748ByPVG5LM0VJAbklXkmVRkAA9ZySjJWKsWes7kdvyY4JFLBmOsgCd+EGu3sSjChUNxNJxebnd
isLhIxyH+PHRtvkWBWR0CyGbwiE5AddIo8XXMCXCEeNbpLCTg37iR7b3CfXiPARhRhen5kSX/riU
D4hc2ekGBdaz6xjDZHFBu2RNpIYmi4zyUQxshs7DR8RYRbuMOtccLTj5LDQyJlFB5kIz5nh9NFu6
Sq0qzZlRqTUYNAFTzEC+QYDyQtYExRNYVA24vXFdbFsqOJd89wqOV/t8NY7ra8G3Jb2Z54n5Ks90
HuuxNthODBqX6hIdvsfuK4xgQgobSnxqllVH14lKNLMuZM+Ak9rj1FfBeScYZjtIoMXh67A+XH/t
exuQsfDDCg8l2RvOBVZPxDtwSZrDhH96F4aQqwS7hPp0yw0J+OGtjNiXSCWROFkXCQEFxM+9WCfS
14sGpHxRzc9wY8Wip1bP7WdvIBGE3sUDnMyOLeI2Q/EvWnyHN+kDl4oxVdaIBD+STF35ZHJCJpui
1/9ARe/sIsh7bBHD+OghYPH2K/hrnhcBwunjH4It8hn9h9d5YKa+H9WA4DgAYdq1MgrIP7qNF8F3
MozyflE+Yj7BfFbWlebnAWX3odaU827dnZfhztxSpoXWxcay9qaksaFNwdxzh7o3jWdPRhXjBCbR
OiAscOsnrIEnRkfzSJww0QR1Fsm123i/FrAzwqZgPR+dy/JFJSKZWlwDpykS7Ku34Psg6TOQwkMD
iPG2pJF58/xwnBWghrkPiEt9ssHm/j9XMnUSML4x/YKPsfBiOFYqTqu4xUQ5pS2US8dAdh0LSic1
TSlpYrD2R0F5rV8TmBjNv9arKQD7j/GusmzHTQGJlJM+abc6QbdBVPspnHZAcnOyTjzfUsu+1C9b
jJoAZqiY/haQ78AsZcfMY+RXzlXCsO41ztGvOrZRSLXi7T5VO7PMH2Ga3QWrO2tFowm/ZgtJespd
BY6UA9oUpwMF9PQ5veFz2KCqwuNZnC94ON1iwOm4blkRGFhyBnVyH4fkrqkJOGq650rgK2Q89Ppv
prixx+e+EEpq9mMzL51v+DvU3QcHVEelfmyoy5+grlJ9EzM/qsADEufMqD9e7/iTo0IjgQcjwEqm
Sv4OfoFopw0S2wNdQ2JuTDYOPOYTrc/Z1MI/JmfhB9R1enrkkmumvvcsi1k4Lb3PSclnq7JShFg3
IpJEkHWQr8YnO6Oloq2d9slfEti01v1OfdP3wxtyB+K1mvnjzQFpXxbr4lmDYmi/mPY1gpPUE/ec
s/YxMU8Fr6XJv6QEGzAvynNdY7Dw+qkKLmtrhErXf5+7mDzTj9TV7jdho66cPydMEbt7ki0a4+MB
7+2q3qL+/5qAgnmLjf6OYSvWHmdNALyvUGc/ft4rDxYXdZiptU4dZcKW5MeM26c8A48p3qVXI69J
Z4SQjOBtsO7g2lK+B76uTnEpZnaPowacVHSmWerjGIMTUPXzR5nJtDsuWHfQ+i/B0b1v4DZqzW/R
XUA3g7rnN85LkGi71VNQ9j7USv7h3FDsX8nEvpLp+rB7twSsoklE7wpnfjX3FUXPcl7MQ8lvZ3gK
qrr8CKsuhh4qvk4oY0J6/kf4kbUWUSDhHcxv4amhaE+dGkMd2xt6Woi03WVGMeVSUpZE1rglyMf2
s6DEbtom0Be55EK1qYpzJWRrw8JE++Ku3WvBs6PsnTWZoGsniEBND7tOsxEF1ZJnxf6Rm2U/9cLY
fDAe4pPdn35OGuxlzk+S8z2pYPFRY79MFGU8xeWvFK9IdgC3hSXtKlAQstme0CS6avZ+UdtmHqHI
tHsbHph2YuP7vR2Tq6RvNIukMd345fRZwVEbxeZ84pf0YVHrOEzalaKhVMjzXOfkZS1BZR3pnHor
/q769XNDw6rbYu4IIck0hGuHMqR4edIoE4//nHalkWXjFscrJG5o6cJ1ETbpTk5xrFaqgbgF6Sgq
baHzpjiW9iESqscDy73eKg0EbvbQoUwH0l4r9r+9V9apwF5tdXmzBQQSLmFaP0+9Ss7z509B2lmA
uEj1WtOPaRz/pMcsAvMhwrdkvQEJQy10KCmHjGaVrij+2PWCrucH/HFRVKbjtkt4rjeRjfO8ahpK
Uj3xRUKdaUrcsT4sTUDpAO3BUhlodnmctZHWfprX6lwZ+eDtnVHnRj3GkUTwcKwqJOBtiB1kWVCb
w9MfovWOP/wffxV/+b8XfzD1O0upfOxWCWMBrViTEfz7FHunxUURd7RSxzsWBB2t1A5pEwyslz2j
mqLbuWY4tp0RgHvqi5fghOntWef1vKZ/9gqrMAIx/arMz6nJ4Ndfaq+3N2THj5qBVI6TWOR1nxoT
EVYMtpMZoG+bHS/eQ+76s+XtH1jbN3UJEyqq+U8BxOI/NrKL3bSThLdOF+H0wVVxS1cf/ui8INpU
3SQt/kGQZ2sCHeujXl5Kva3cK9MJIJIGlJnIsk08fq4qbQ9m6qqPYBdUZVagbCqX2yKJ/yBMLt5A
A0duWu3dIYWAHQxexpi5MxL1usGkL9Ypmn9jN5amxNkJHq0Zw35mBHRv4qHfUyCgN0i3OVfs9kEz
gWIgGB8pRMuJqO8+5tJIvejhGzvefAzXv3VtrtoLg9MUfTKpzHzySmvxRe3rG0UYZHc+J0EdBUb4
X8AWZ3Lus1OgPO+L5Iz8x7LyEBIDMgA5NnZ9aBU0OMmd9ZPqUu7wlQhyjDVhLT7qOLjQ9nerT8fs
AjBgYja/1hRc+w//UrSXy85XQ/OGn+SPoRqfPpHNCeFqlw/gn/CV5PIo3QiBtMTtmakrpP+pist9
tMqiQT00hdCV6Lg1JMNQCnkbzh9uFnB5rbnHPJ/fUJ182I21k1Xk3A5mPn6pzF+PyGA+eH/mhQZl
qeS2xtR5nMxxTn9MoV/SjeSkMWJ0WWKfIZXX+5OO08JfVDW9/naA0s8AvAIxbibQy0Ux0O9zPQEd
tKj3nnV9/y0QoI01kZGB1E8S0lEi/VrkhOys4bfo7UDtGvxFniI0GlfwFMYIuoP2LAGe2y7huHPH
LJ2Vn8e28kHgU3IXeWg9ccJ7nAYimd9iCDhk15U9NWQ2APSSO7ittYt1r4NWmd6HsBRXPvbO0O0P
8K/IEHevz/dacivCP5hnGwmkUjQqYOiv2jK4Y/uCcUNBJPMVgzLNaTm8fGXGSLWLIQ5dZNp9HFnN
Ck0BgQ18k4w/jobP1AI9vJFv74zoc7beqJCPvM9mYSUalDOHwtGFqmGruFjpLVGocktF6lEY2xuL
LqZheoTIJj5w30+1zDf71Mw9CsdLFPlpkYcC+4H+Mmq6lh62MFyqC8Vs2v7bTgug3Hc2avTTMDO4
oaeb5xfNprbbTe/e3xRk9wU/KA8GRFD5T/NmYEWUwVS/DKgR4H7LdYh9cDKPtENz9yJ5EtUBT2AO
r0oWMzncjdxR8mUjcIcB5AJqfENBJlCloE4MzPjHbsahZcem2oNkJmewBVNlD805A4NizGEWLqNo
OWqjz2zuYHOqB3hqQmqbxOLiztsibfXOaLcGR2M3EAxAGcLdEE4SpY8kMj1tVuhTlo0xu2k4Qc0e
AVKseFC+sV+NFxr+1kfETW120IgX6T1h9wq5yq/pGU0ptU47a0yxBVcs8FA2Rj16cbXq2dzkehWl
9kSkrZLhmA1y6YqY6cHYEJYQKT7WF33NSsiBIUInR8epXjVqMKQsJVPinICLTxFejkijur+0zxyh
/dwH5Gmpu6xOsvfvfQV5t7vuFI6d6Od5RB1IkicNE2KxTJzZRW62uE3+ET6HGby/xoB8bvjEUrnh
PEV+SijUMgsCDR/koqjKO4UXnwVajhL5jXP2CaJosnvzihr+vcsnN2sR1gjg5+cs0BNBFq80/ctR
teUKLHEjw9HXPnAyULreiK4SZToa8NOh9pQdMh900EE3BvhCPYy+SI6YQHiGVZMuBdkXZndah9CK
mrVYY7A370WTcLsO4oYJhgjKe5PA70cIHQmDpcU1+NQwS349s9sa8KPtg6yegscLQKEgx964d9LI
U3B16iL0PudYRJ+q62ES7vGy5Xx1Eps2p9Gn1snHiIOu5uIO8Vai6HdY7y/vLJr64mrBQOfwGJIU
xc3fio3dmv64Agxdd6T06JnH4s+5JpsW8XZsumdi3+CP+UJ1ZbreELiqhrxNGlPS52XSAAfyO7cn
/jRgWB/vZSLMkR15NmBTPOKsezbqOsGx8VYhCc6HbMnV3Y9QSGtnIu+7XuJgtcxUNjPN8TuhAxNG
FblBK8rTpcwsTFm6yEasoyI9kBX+8j/MmSY6/o05bW+7DFB50BOtaDVSFBCCdSttcCIuEjaGxmRG
gSiphvzslQy0NrbB7BDAFsohKD5KKzP22rTdguQcHnnhBPmMqtZZb9ECotfZOp5I9orxBIdJEyqX
6FzlpYxp8KU2h2bnq4bfaN6lJV+qDLKbbv8NCD53xg/EZNpP7JC1VAzG81aIXtlvbNrSj2s7GuRZ
f5uPtVMtyqD3AjPwyArk5uymvuODl2yTbQwxA/ZuNdF5GNtxwCMByzaO7oDsc0pAEXJpJ8BxOlvi
ExYYBiOI2pnljRBKT5475XmfrmfvPm0BPwt/+x918TtTFjsAwHD1mW1VVIq84wovD4Ag2nOlSWs6
mzc0eUIZEr82mjYPr9HqZul497DnwxuRXT4AgbBvX2I1+mF9JzCT1//s7tjW4BkmteYhNGYg20K3
G7rhfIU9Tmj2ncLH018ygFJK86tJtSR3RXj+yni6lS2DHZ3RffbpUf/Isjs9VMwoEdUl1uyglQpO
SlyrVjNoc+YlwIQavaXHeHodOFWTl0MM8jZv+et2Zpis65HPsFlJ7FMtQFgdoFnobUNBJo8UBlLF
Dy6ovVA2bAlk9FAuCxdGdAFK+e0zQmHRf2TtaEOrqQttF0FVlSAssfkFJU8e09h/V7Fo3wB6xQXu
EkNi6LyMsrIzBtmi/IEAs5ciaG9ZSX99lwjzlqaDOJGVnYpHSN5XNxYSgH74bTgdOibyY9HD1Hd6
ClG55w7EmiuOnSy6HTMGPr68JaChwKBZuPIqGT7RmGZvq17JSySEKtgVhDoADhk5qba7OxazVlLl
GdmjiI1bWfAZ6rSNwCVEHr3IVu9+BFty61WHx+z8fpsuOE8fPOlXPKshaa340zTgqVkfrHZfnDWZ
8j/JkXJVgX4HrqjM5Wd77EWhbfXBNZGOkIJETKKWom5e6wX1CNh3EGFp7grY4UcifZBO5cJL0nVR
df1vKt+bl4o2ol+5eR6LmZGlqHVERLbayIffmxZBsxG0/0xCfVaInm0s2fYzIQ3PxkT21NXJjaWz
zAh5WjVky1T5zHFKHdTo5zXpCFsbgIhuc7/ZpkeC8SSLcoft2eSJ7EtRZTPsNWXXrc99nGTcU7Hi
L+2RFY78OFu4LRcsPLC7u0XLJ1a3Y6XhWI8GmFTWl9Shx9olCAmdfakLPmMXdVs1Dgr9uOk/hpN4
QOZvKXKrKTZaEmBTzIGjQ8SIGiMK8IcNtmCJ2x/zhnAUk7kvCEaExw9fun6zGoFX/eGzpHPiKN+N
ZLveEkYKljbq4ZsQeJB4IWUwtNKMEN1FSlitASWeVChcuyXX/pQt3Di1xuxq92Bh93umxgxI1mJq
XBQ2a0DCojSd8/AbcWBHNu7V+RhvqZi8bkCQmFABx63Uj8Yehocz23CKjnYnqsWNoKjlx8WvuK37
XSXvwGQQJb0KDzTLElgrEIvRIBUGUCTzgfR+n8S04m6tuo8LK7Dga1IsE2CSSA0V3aPHJOJQzoG1
OhDelJLBXchRZ0/RpIZK+BNhSFmZLZBN/R7GAZqx9Cg/qoHI9MkFj7DpsHaURYfmgQKugmW4AZCB
iwIpd1vTyhkacNRNLFuoa+HG7OWwl0ph9p9lgFu0tZbvUyXSohScYca18DA+DOqxktlMXk+mo6A1
iQ5x8ez3Y9409IgmXUoBBI2TuxOMj9hCfT073ymfMC9vZGMzum6+e7pLARF4VOWofxct7aWNHHCm
2kq/VyCCGof7Rh02FSX3Tfi9rRv+R+hFvxrIQr6juEXZG3DEmvOJG3kL3tZi431ZVTLouCBr76QK
NvKg9mK6vbSGx1WMMKUmSHOtPvTvjtdT82ODTkngXnmubqPn2VuYSOEWJrLb9JERb5C0AL1YOvAD
X3qELTV/zGsr/KjRRPg8zb6LUTTHmrUAZnGCbNlcQSRWms+aktE6M3x73+I83/AXMyVfN8Wrko3R
lVCM+Xb+wwM9CB8tkuGrsklTNUnGDFM0hv9lvpsMmkOH75gQV73Adnwia8iDbH9zAfOPaOzunm3L
G7bdq5RQVk68w162gg+YqvcT8JC29beiiztAxR/Wx121nGl3QtLvGb3FbU0FBVv3BSjF5fkAbG63
ObwpXaBnGiDsphwIxlkCL2QXGC7OzArSxJK2e/YacnlomouD5N4GIhaaBjQsINGtYNxx5HOJ41kR
sxJxzfFQl9IsK7aSTfHMB2QwkealQNDz3TjA6y3lgQGCRhYS9FfcJovFxaxH7wdflf0qrSpnkmb5
GZrixk5SSATxQJpZ3nPB98XjwQzDRao+ocCHzR39xlxldYLnmb8aZWiLBnlLTNKVUT4XirmSIptj
K686K1wLagQfhxMp2bKJT8zuBeTDNasTwuMYVoFZ0hmTJQnNEN7lye5Q9OhsTAOpvmerVzeDT0rg
pxPHGT/SHJsPh2aikuFmOBVT61DlA93QJ6fTdSn6JfmnnfJLoIVUXBWZTWv10LdPhzkDam+FMSWb
cR9Xunn3ZSdWs8RGZl0C8LX6aNg04pHirBfHPNKPOu+oKTiySPEuOgNENo9q8o3V3a4CS9tU5moB
gjc+UWTu5OLiYsnrYT3l4WxNYpRyI5zR/6Ve/2xC1VM2fXHyw0CbtSNjuCoaz9onxghJfl6bIDiB
VgdOB4YscW1kPPYC3ZKejA6A5aApD6c3j7iNxPxl2SyiP4ao7oVk39LHnDC8kouIsTTa51nHDf1Y
veTK6jvHPZG/M1gUclfjTt5Cq6YL3nz8MoaesSk4bnbE54+YdrqxS37NV547fNHdY1o1HFpY1pc2
lwW3eFVrrD3JyhIcWB2vz8qm5R5vOZQLNRvyzCHKvOyvdFofmDDBJjsJ1IyFgcimXBla7fSjGEmo
sA3XgGcB9IrGsOeQfDWbyJPn2AhCsh4yJcBJ9LffsAeLfjRL3JeNkldjhcXdztED5/18f7m29LUC
IMVTIocnUOAuiHgV7csIWuuE2HcK/lz//q0kGn4dTMF07gFUZrRD+VP+VAaBX4BHhRVIHXorx1p1
8KhShx7QkVItk8b51b6yssx4+Z4/6TxM/6r0HULKZmeVusZqgvNYMVKzZaUyWB/FkvT8qSAF0vKE
wDQy7juf+ygnO4glRYoVdOmd9KApth9SUV2xAnXxy4T8CddwesHRym1aek2QqZvOQMceKNAQEJzC
peggsuSwSDeMPTZZBjPAttogF3NDd79bwxH/04oPQ9sN93C/puIKg6N0S6pVbiNMdy3dwMJ72Evi
9nSN2fz6GGb7fT7CkA5C9xh9/1sszwMjSxWXJr5Vs+8P7DCh2hRYnW3Nk8FK5N661JhOrI1aGp9N
vuASxR6aeQHQvOWlAJ3FLSeRwkZTVQgHMyarngfZtTHEY0y0o8unazQXPxLMm5mFs4hFAz05Q+Zj
6ri3jr3tLUURU1Qa/feuRrnWXXqQnjPBqrsB04Y8NejwB9raHZgdFGUn04+XTeU+mI/7ozC71oBJ
edNjcZ0g4FWlrE0Yi3V7sL6GiHOpOGGgjNvSDRSJj0n7g8SSX+Ofnb56KTR7+VduUgC6gaC0TI4U
CAvqsfAylyn+QSTpWX0cBaDMr9m6GoOEhI6AKE3NIOopeHRqTUB3v3oPNmO/XHBC6dvDo7gYkR3f
F9VKcbrNguaxe2ALJmyPvPXsu+b84JH2hltm8qVbwUWqC2PvHpS9gh/J08QzyilMraUq1SKJ3WWj
S1woahTqJVusv9Rsuq+ZkQPp5f6FMpPIbVzb8QXGcZ4WabvP55bHlZGjACQzP4mOp6ho+6u7GAQH
ui4T1Y1vG6sJK9xg4oWR1gf3Skjoj+oCC6ybx1/hejNMovTG4c6eNjQ+LyrqhvA5m4CRUVRQY2z4
Euo1BI1+vYqsI42uk1bkmmLplUsJ8w8Ix7RNlUXUWRHpfSILQ/pD6eXq2YzR/CGkOKQgO+PGJm08
BlzMGkSJH7SIqIpTHc9PlFa5xZWj3UNMYVUjRdYd7n9g/eT5LevqJQnzO5lXsdiHj0+o2LftZcvA
pK3k4i0U5iY77LjYV+aAl22+6HFlR6Zz9O0tW7OXfmLvhLE7bPFeoWmYFKbMnmrJ/m92AfcHdmv3
bn6UKij9KjvOuMEF0t+LUOKx5ZTh30fsyKljbhx8mCwUi20AhZhha60DE1FLYR0/vxpXnPZTQvo0
tFsvIItvAXEizDVChnrQ1MvviYQcgva9T0oNa6GZQeknl2gxf4DmRBShMZAeSbgkK2GhScg5KXrN
PO1w4SBNb/rqlWeCG0oh8wTLH+4hz4PZ6pPBQYKPZqHrb2mONaqKMpgtfXLpYzF5RMlgcBe6Tizb
b3yiUryV4p0Q3c6ZR1oKbTJ2WLwilW841SeiCZ2/pN0hTd+MsO8VQUeZ0T/2BFXKGcbZXXCbl6PL
wl7/3vR1jYUWs9rk8RzxgQYDLb5zMaTPe5KkP4CRMK6vQkn8SzMRtlsT0DETjsKdIQfCh0XeT05M
3tF2iXOZoUw241F8x4+N/dnyPKPD33kOqjJ2t5WhvUtg5oNvyQ1sgNywk5DYOMTCuZEFvCwYFFoT
OYS7vmtqEjCfC1wa5p1E063vJTBcwZu+AQbksYYQOb9XZfy9RE8GlEXFG3h8pp9vWLvcor6T6P1G
Mks7bu3NcvrF2PhnCknmbB7pQzO055fWJ1wf8xr7K9mKQV9VQ1s6al6H1i9UQq4/faDAElhG9vz6
MWsz/S3Ev9t+Ro9QR5T9wDEaRMPPgJhl/i5/O0EvJFuHK/GDsiR8eumL1T4xJwlmDDsLhUnp8ggT
3Tiyfr5hXt+xHi91ajXQJcuth9R+6Nig0Atuqb7IlL/oMLPddba0EdRipbHX7LPpdvKS67RCH7bA
tsk/txqSWvFUcKFFIdcc37b0JEuntVCl5nyuPICI6JO1/tVqzC0/BVvicSIc/S22gG/qjcV7cN2s
VevAQbl0tR8+7HrWbvutKzEA/qWYSVAB0OaBT+aBuuEtKHnFyKPQ1P5X5WiS4KvW9krI87pXUK4a
lsTXLIHrrjMu+tATbGeFmtDFfoSufsK8kzD7THt38NAtCBf7QdGs0Oc2+pFB+zcxp1jE8lLJlog6
z+ocpwXnp2J6Yl8/YROhAuqTPnUWVFYyJsSls6MJPOqdlHsaLxzb8FD0b0dsHX5NHE+H+HQauPgx
e0Zp5SMih8leA4qRlmdjSS3wwcjH32GP11+qUhhkCwgNB487PSpQ66Sk6Hu9lEchaXPp45SIXw0M
D/kUOotYBJ2XypNYV9Jnof0OyH71DQN/o1Y+E8/sXVIKijc8VXXLu8BC6gD+/5RXI9m01a811t92
s6Bp1D99GPP5DEhgd05ijBbgajE4FHlZ7yoLoHC+hFveJJ43MLnxTuG9yVhRj9npsgH6Zo3zLL9S
62/cXGH5Q8of3MtmP+BAL6cI/FwZ1CejyzhYw8l+a6Ol9DmcaZCxZIFjUkeZeQKkWM8vaAUbz7gj
QDjNmCRc7bDvlxnrzfWCgOiVGBSis8c9Zi3n/CpIRy5Ho6nWqwMgMs52QGzcSSOhVV52KJnHfmzX
PZ5burPdUPyM8JHAbrp4GA1HIf/lINZiQV6JPOLaZUknGzBdxpXUFuB43Fu5pzFS3YYQjfMhiaAh
tO9VgYGyFh5IXZPKAPF4Szg16woPcWAoy3bGTGKeIUKcick5CV1QsEpyGYSke/MA6S+QYH2fuNsT
Mqw5YQGAw6aPh9fYKIhjX4PzM1qHK7pmtDQ7xRriAJAWC9YgT6C74sNprSzGTuieAxphItAyDDZN
BZsBvJz3CN6rGVMSw5H+/QeC8vjreKpV5UUdrTlSDLObNhUcsnhfJ2ecDqffdaELLGfHShHccan0
OQhbOcvdMkh8YygrmodvXhEZgu1yjMd7d+4T6Mw7YUsQ2eqXzDtslOpnbnspMc3MkyDXzX4Wt31G
Y4B0nbQo1OMnC3UIkjgiyI+82LEnqyX0x3Hg1Cv6Fb6qzAVIgK+LpU48O1K2JNPy1rn9PxyzsFlQ
s309sgCWX2s2iLdQkBiNCaj7LDXFbejDexyNOLJUFAG8mDjU/80r5KdDP7lKhpdhRhbth6Jnlb+J
ed7MTme2FsMpmjG5sKhGUHpUouIk2yLAnfIm3p1oJrPCPO4PkuKg60Eas/0fnurjx7/DUa0fdPPb
iOFfjP/KykUUaZB7DLU8BwUwcVujRiELRRSq8POMorNMV2O/wOlTErTSm9E6n9YzhHAPogKD+0Mj
+kbp8PoyPq0FCm7x3roKb6OwqQ//pExZuCZT17LCPBoewWrLKdr9ES64DF5c8vfFsghPUMf6+6w3
sv5YcOovbK2z9cf9jkL7pYMHWdT2RAx4o4Spsjw8pL3+yxq6CnshAHlJMy3TlWQIKK/4RNw9OtWy
OoLR42ztZJw0dtXcqXcWGySOiaIRjKdfFP9kp9WAAdp2FIntxwTzHxyBzklFkTyWTLY7YCTr8OW9
6rmH0VQG9ocx2IAflB2yvUKaAraOa9BlwNTmQhQZe2HOV7CptGgd91ALekg1GIMOLd+7rlxCSfCg
K3bqadp2pfiybe+rUb37ZW8W3V47HP4XHFfd3dPspSy+AMmaTul7kq9VZb5F42hCHYU0ZwFcn/Z9
qb/A20GFdXcOIvTm0WT3/3JzHm0h1+tVQgsha1X8VbPWX28vNt21nzUi+c9jz427IG43HXVW/5P2
oyQa+0aqRwRSscKuJkxQJD7ye5M2X2N4QT6ME4NOgeFda45KweI37ps0J/uasFXC+GEpMlOtmg1i
6NL9jY/c803BrQbKlKrVNCOJN8X/mleuGRUIst0olFpLsp1Y3q12eLesmnDU+COPc9vzEcmtZB+o
Nxc+kl8Y11j0+/p/c/7tMh46XKZALZUc6YkegMEFgQVUyoCPV1oSAiiddd52cmOVrtt5jWle5Im8
x8Rtm1q264Ss75AptZQH7WNJqWZl+II8qqaSYO/HC9r+uitFEG92iyVtht5VR2WL3SV/sGPu9+9a
6QRK1JHDZj9E3UeMFq0roAvcAyk+NV+tg23ew6LX6GmfPRfz0GO/dwF9bvDS32w3E3HBQNFTUmAb
0JDBIBOmrNo/NdkS4z7utw/e6o/xQmHeQvFNEvvaT6wZf3brTdBqOKSxNVSSgVPk0+M1UQfTampq
8+4skchCCdxA8WILgottC+F5TLEJf6oFsMp/Efopo1MNre+wi9fSO5icqNaoMwhajLnZZXXgOuJJ
fmJ+MGhnv+h970ILMaQ+EsJcQc+ej6n9ItLUgNABpfWiaEXaGG3wc2tnp3xJd41BkjIDKqiFiJi2
C3RVx0tjP1IOywl2omHk0J2DkS/ERvyZIM5QHpg9YJisDpAStirJmZazjG/7L0bIryig1NV9Rqs4
V1FL1LMaMi63rFEHLgNNLnhCsqzkyFe2ly8KA72LublK5ibyC/koWjFbOARy4YUnxXzieUiVaKMH
b1QsyahcU9wPp5/DpfmHko/BbuCNrVLBpFZHZTluEcowsL6DHjpSQrE519Nma02NNSedZY0vgR+Z
scOPIbdj6gs81GGFuY68X9SQUOu5Yn0uZPmInegBSuPD8iYDp6ZdhQVojmrAMuMqDgiYdrkKzFC/
nH0+HNPM+2uaCCESpuNkZl37jTTSd2M1lwtLrRkdT1618/AR8olTPYWLx+TEyZ9Ey6h/3Q6GQ4vF
DyUUKCWgBFPdYPrlQkDyaerhJI9u36xKCzh9anqoolOO2TdPchlP1/apVK9VaF6brHYtlf/gP+HB
9/jheO4ckk57SHjUyYwMCoUBIWSVAHOAxalHCJYOrymtM9OdGUujDzGVpafs2/0I5VMSjmeexFwJ
UtTbdjMdae6jjNMBW1JL5e0lFusax8IDJ9ZoBMqKqKlj3tnf7ozKqFe+DxwSoQ6LlOpNo+SG5fSD
ZiA4EFTEiG5U/biv9YJLuyC/BordVSCzhlUqQc13GkjF8pNGiwR9kJj/X6hovBUluPkAAP3wvCr6
nX5WBoq6ua7dj7uGcbLgmu3si6S+S9w9RcVqGjOSVZezRZpm5hiBds1WAM1LK7BdFLdHYOHyOiWC
xiv4EfX1UO5C+9hGXTJtAzXfq4toPcG8IiXRUiKpUwn4TebpwaLoYtWKiYoqgkIjYCwpub8lNDGe
EpxhwmBnj7PyNtYZcV7fYU6xgqgvOC2yDUAf+SkYjK5HAN+ASSfhoj+kGBDUWaDp1cczjRUGxTfH
M3IkYZ3AiG7ny5Dej43rGxGzTLbegdzJsVb4Q8vCBxhSOFL2kaHdn+U1IsVACNCF0LpjstFQz4L1
EAsybujdEp3aEmKL4c+S+VmSMhw0GKfputtj++xG2/7eOLsiaAjZyosMjfTuaOhIO0LvVOvlauv+
Q9PgKgQpA9PHwBI+fD8wUGKi4FpRYtWhod5Dln4wJ+80ngukU/V9NGh8rV+KT+X7nPKDWfNdztpG
z4S/BrbHEjWA8YVtH58uXusqprSsQUg3TMw/NW0bknn+AJT9vnsQ3PnYoj6Aar6hcmp4E60OM3X2
al4s5w8u2BydeIgNxsnVZ1ASA2yHrnh/KAQjtPLAUROVje6zKQdKMPoSurPw9sAxNOehSn1pRWrn
PePpbacyzo+UqcN8vCH3boFW0wJu1ZScEL5Zuzj8/ELrrtpDIT/KmCYHIPNDXSA4bSgdRjwuo5Di
TIO5FbgqnOUOTRq8AivoqCwZDppVcXJ9aWOQ9Ko07b3EFuY8PPZI8womdmskGjWobc3+9i6LRhyS
e857sdli8gS4ghKj/bXD29dzZ/O02+gNUNjohKkZBowZ1fEXY6I6xhlMa7Vf+9S2A6cFV6EuLO9L
IIPHmEnzjfW7sm/k9oiiIk5tmnxpwlxE26LJgp4K30fWQb8OzrD7Hnz0R0b+k9OC2wiN6nLL/LUv
iT4M8CxU7oen7o7Hm+aBBGmMI9tKKM9HX5QvIQXfu08GicqbPF5IaS6kQnSEg5SIsDl6IZYjB2Bl
0bIcicsAyZ10nH142IGmwkLnjd8a1asYzW4yeTDopKfg4l1wxwxBx03AzVcsU2nJhYrSj2youEqM
eo23kapfBW3TGah5vEKuWvTryl7SayYJpxkIi+nkV3OjyyMW031/PN/80mXVx+iYzWtdNKqVA6Mq
HHWRjFt7akoJEqQfFS7UXRYFG+4UsqgEWO+Fk9fWF0VW0mKA+e9G7J+mKLkNjjkZYkL4VHTl55C9
kGnL01qqyc7RlZIMEWHBd2nQaEB07DJgfc7V34Dt+1b6MP5EnFYzHp06kQErwWEB3W8JKeDZipsz
RAqIB/zK/7xeY0ieMYGNts0obZUlsGpsYLwv+rhUjTCxRJXT1s+Nrpc8r3et8ZhAb1k18zGknYon
EdKdBcN22dbWHcxYxrr4ycfN7SZ1/+G2/wL26/kfu0LquFv/Qj9oBlAHhtmttVjridAw/dn1aOpd
ERcEyI94Xx8+vli3PBmbXvyc9JzxPiwhGSUrJxqjR+Ptjdk+MRjoCSEWZs4/DPTgZ5vBK1Ha4gVJ
+hAAZjw+Tp3gTb1onCMMgdkrOe94pnERl++mx8x2RG0N43KDEdspF8PI9FByqEEFHvB0FQGGmFIA
oSgEdq3Tf1mimb3y079rjbYKEucLhbDePAKsyVY6ZAWejE1/aAtItTCbfzcVX0FB1LLHrAEM2Y7P
kfFby2LWLl7gxMdmu6vmXhHvpizd7VO9GFD3nCgJA3rFICNkG08DMsOtHmKM+P/RywrqtT/Hv6Rz
mxcUsrLyiRboYDYEgAz+6LhzgUPcL/1GSIhFSn+b0VxwuJtpnHGXhLOex51UNo/cXmCf1liuxKHD
OrB/dSv0R7ekbLV26KBTM2WVve58aQj0Drot3yDk03c+uKd3ifOj6XrCu4K+E+yatpMCBcLX6t/0
UhPqQB64kVecS2nktUxk7CBLps3+LS4F0JfDzF2TVqrR1x9eXxEqzqg28sSx0AThHa7zexzU6bU5
27rIAM4M/q1CRgG+/QUIY9YDHrcb4Wv2eLuTRLNH97ldfhJvlHkthncyyEQtLiVXCouI2sx/WoJA
TsxWcdMA9wB8Yn1j8bXqTQXsGYOcIZaYK+GTirRi9SK4uFj5roxFxaQCa9r0QkdKjRaDjrdfAnMl
yt31QcWOsm6Tmv8fSE8lVw0wcVyB2gFyYhDOyRQvT/C6DZUWChVymc++S/1elMwKc+HkOpFF/txk
ck6Ye3W5HcjKgx98ylmpb0tmdpGPtS5sPwR8f5wDbza7gpQu6ZmKYYBCorEjO61k7Oj+4HO5ohYN
QJjRG8otu5BCMZyxf4aJBBKKrEPxHOj337nq0cL98inxGxdenwbCkH49wDb7rrZyPyYJjobgaksa
NnTEvocCVKgIDiRRZBsiJWAlUbIszUvdsB5yNi+nk93R2Y9BNQoWU3Spwchhy3pDB6Js1CQqeWj9
p+APkyf9UUwoMxEFNQxRJO3Y5hmoOLMFhMrImuo6Q3tFGZvQmbPECkE/rtO+Z8nqZyv4HzkA0ybj
9DpT/CvHhoOFYb0k3f/2tjc5sllY7M0kXn+n7HV1i3q83zJBBoc22+KvsNnp8ieDPTRuDTm4hm4Z
a0NDt/Xa+Q+NL8+flQjykereP46uLxC6e0HbNH03XXB6eTCsnlDulHURG/BYbOTTvjWO4UnWPv6+
Rnt8f4gJ4LSVSx4PapnaqRKqt4410CkQXth0avTopwwXTwreZOFjF6i+Im2n3F562KqeMJHJTtqR
qHZe9WwWJDY14fiEjioeGPwqnk6rzT3+Yb1mdMMLNHq9JF960HYktjbr8LlUV7KwFQNz8QWfIPEp
Idt4CkBJNRwnhDL4IkhpUUbf7BgAJ1u2bLrYO/S7y+J4Q3O8gsr0I5iwOZFJ/sp78wapcQ/se2U7
V3skqxXpB91pDUn0+I+RpnOdt52NGSTSrlMUsNLB9y5R1Z8+/udtwzjoOF8wDjlfFCVAegnASSYN
hgindKM8B0l6zqbZs9HeS2fMWmP7QIi8swe8V1UtD5Hp9jM29js+stvj/6/ugl+E5GL9hVrh+Cj6
hI2J0W7LzLRRRdIoj0blqvhmhtPhMf+hINWbEP3YxyFpCIC4ze8vUto/QiVyWrmIS05Uhf5rVv7D
7Q6XIq3YZaYmCBZUu6YWZxBOHljzZj7qG6mWXrgy0/D4t/g2P2+nLQ6V1sJoGCzu4DLW4HNjQVpK
7VEN1CaeonsY8BYKa60DUnjY483G0WljewG4cg09BF+uYIAoyDzbOPCVWNqeDvtAd3Yd/0bF//UR
Y+G9u7eT2zE6Lq+e5ByfoMzJn18Fg0/hPRqAY4nt1kMjBK2uE5ojRQvOcQo/aqZAcX9UtCKFYLxD
4DYMXSpG9UioIQIEqKusDU4Ubxm7FSfy94T/mXlqq7NdQUgINYF6AtzZXO0CS5jGnRKhraa2m9V8
rPUXxkyO4SbJlqFQNebiaAiXhEhWgsCFXnV0vR7ePMfHJwHad7PLBnRCWHBWbEdHsKOUUZKXat0c
jzOLHIm8+lJeuHzvRGAB8kJP94Wyvh3neO4dKILdvq+uCjQEjkArmZ6nOnrJZ6rMH+E/AS0XCve3
4g9aEIXfg1sv1zcHiXAFDM2lCjpFKg+Xc/AAHWUehBuXosKdx01U4zXP60LW24FPuzbxvSqJTw63
wNn3H5OZEGPhhmaCUn7/vTLM0mC58WrAWy4YnJrX52a7sYqCe/P5EF/51PPk0Z4sRtYfqxWlBklT
rdmQXzDRiwVUyNmLm5zH2QDA6RWuscC2maDZW/DpDWEIpPkS5xYWMmgBSvfdUl+x7Nx4tRTj2kr0
j+kJx1VueggiDGXzdwNwfEG7OZlR2a0YtU5ghaqKM+6NS678rBi8zhorcQ5GP1tKQ2vnJ3FinIV1
2G2KtKiWt999DTUdakxq1i//0AWWDVLwzB1J2L7Tojl009GuqD72HXNpUqOcxMLb+qfLOQTe0CYa
H0E+G8Ft/nJsLYpTdOQIEvwSgspJqstKFU/2VKJ6fWcvw0sYn8LQTxccGClFHj4XSqjv4KKbR9rk
HgJiEtYQFdM75eQp4BtoVWIrdn0myywXM0WeQmj97suCshBhggqq3G0m9jZ67ahYTC47SUxkt4zM
vpu4m+Pg/N3q0odov+f1wCqskoam8/F3pvkd941n/ySEqn42TXwvjZ0HfP/NaY73gX6bxusJheMd
fsXkKzyX08PPbYXsgqk8jyD9dA+8TqCV3SvDFAIEXuyRqPVpjRmhxfs2n+2OgOdd4RKcrjlhlqM8
nzl9V4Bhs87rk8HynbT2+kZfgMGA6WGidvJMrrEJFLmmCq/SzNnFdRXyn9N1t6klNi0EoUH4k2fC
iRzT4NmfYH9S4VEIyT+cnVdTEtTNQhFOocGbwUegXRViDOLpAe1wBEi+GiEfOZb5HJ5EUWVpgrQj
meL/Db0dspLq3IswEkVBnmzhQziXPxvQcLK8PjqSfhLy/Zhx+yLtD4SG5tnYkngZRy9MfedBhlE4
H4LTpfS0tHZTuU10O1ZXfu4I4S777x+HRMwLOGkQeBT/sdMwuGwKgvb4uown9jUXAb2ZKn1y3rMp
3RuYzmq8zCjCxN/cTtkRUIR8VIVGT/z4uD/TCmGYa8AWyN6nt3/3iOi9m4qSBJBrguV7mwkIDaED
wrR3EW+uTS8/BzIGMI6FTkCdADmAyQlk/0iA3mfZulbrri0BiYX2b2Z4NAoR1t0xxl3tdSjzojIb
yXTZzbXPl79ia7IzaaZtdJqgUXv90rHhP5bZyP18FM23gNuZ5leuykVkbfFsZkHUf/uQwufABhXj
7yQIjSvAKQDDCHhyIsc2l061uy9QBSyWKnxJuQnoM9PxrOrf9HdkolE4s6PqIDXwMho8Wc8qiH0L
PPg/44U+/Gr1S2aP+761PB2RHx1UKrSEOfWQtJtrUA2FviXvhiiS6hdN3rorvaGEadlvzN0ISWEU
e+NpWe1hbLXWIDqUQbXFzhcZEkpqlkz56m04Ugb9iUVcf8iA0zRJnNj1XOD1pqvrgwoQ9ICU8ZHq
VDjvGzPsR8+AhClB2Oy+U8yORmsLcm3hhylBEuXDAm8D5ByKv1kbMgsY1nRhYKjwWS5z2yd7Ci9a
Ogft6BeYrp2xmia18SbqJP0jcT7V9Jv5ddJ5QaJvEwveLe7zAFZZbCVJiWVwAiKuLi+6dH+Wn+MU
CZoKf2vk1Oqjai6HECDQ49INYeZD5COKU9A7Gzlq8KbQecxZh2+U7wooP9J5hmw5e2dw3ZnR/Cqj
+iMJn9udG/sWEVWG+WNfZvSuiXqg8PNr/K7ONnzpejU4dMccOvT0bADskzZuO29feEoxJuX+ElqT
YZT71jf87hJHN9L4XEC0kqysRZ7QDsJpcLly/YqwlpVFfIhJxpGfAGWq4DYLxNDnPH9eGpEm7wmD
pF1SKWjNOGKJ+jfK1x1we0Txj0eIX5kgrgM8yvslvZFdO3qTZEfYskBwuVnAeiZJ0j249TI5/Nj1
eEOJ06DnIVpc0XMNicrom+NfIqUhKXCGJa287nBIE6Wbjve8lnESbakV5IglByZpkJ9OtxuKz+n+
ju3jtV9y7zEERs0t45Tx0orV3Y3nHmHH9gjamn5ol+6g6xxL5PtMJD2BURCVW1Bfcs6Fu11kUf0C
rVrF4kp1rcFJsZBGvs+J5VlDFrcjt3EXHNTema+hZPyQv71YV/kkh4LQxod8a8YMDgDwytjcdcEp
6aTZ/d0gKhceufs+W6UN1WaRfbITsujH4zpd74zdvG0lf88JI/V/HanVCLPOr0H0Mv2jsG+RSML1
UKBgd/bhGqU9NclxpccH+rBy5i6KSvMXSd8OGEGgQI5P9NwWnVxZ+6xQpdvzLGSPXiVx+z/SSbwh
kn7JPPTxJGII7VbH8RxSx+5awgPIMKf2ulTYy1wE3n90qPxkYPWkX+7N0DQXTywqgvOwNhvAm+VD
6hY3zTq6vN0/zfQCwbxiXphe439Net8amzrGqQVkCFGHCKTKSuKZj3ZQJAADcYm3aGPwuIoNaVsk
vbW8D3Duwt3LHwBKyOQBjMv6sFsKWb/KxVDEwgav5/XzjMauIYZyv3pnMZmkOWWE02/OxgX3CwYI
rHpdvQonM5zg/HTJXplfi160Bh+cBAQDvYNjx/SMahMGhaUHZPEK+Vvf2JO9P/uBcE6gnNEH8R3R
VACtj5M/VlVoJluIQt5RBO+3WJ2U3/fpR6YymJAX4Z+xXqfWwOkIPf2x6wOMK71Pm6g9RAPhjT/G
SuVsYah8vjNp5sVxbdnCbjQnUt9DyaNoU2n70ncWZeLLCHx3Ppk8TSzZF+1Zv49YduspVFmxGPDN
AcfE0JPK5cIivlgaaLIL7D3QgUZ7f8wxkUOLop+kHNwL0IcKeJbYlEflb4LYTF+o2KbzBA5J2rpX
Vwbp6NIbaKRLAO4/7Qv2cmXoxm+3PJcVriZKaFK4uqJ9Pg5mLO9jB3UkkN+nvaX4UeOvctS/S1hX
vF8xsuIlill1H8IGLGY12FVxnsgxW6BrsQIns6MdUO8pb8glwCk+Z2KbFtwnJCqqp7j699Ku0Dk0
c8kb7TA7YER+L6MYCoJESltc5uF4GZZXLTl3xEnsb+dogJQ6xG295oAXEuytqUy6vi93eHvJNuaP
MFt5GV0hBvfaTlDukfv/b7wANNk5+7Srz5tIH/gek/6rZEyn54rzLEQpaJZBUpBKXRvptVn8eQzD
tJzAO0EICFikvynJ8s0SzNwLoMcJ3cs7XnqGQbaPpZoiFm+OadpAS7VqvwjQvszm6HxDGxQBM9Ej
qymM6cyWdoyFjQ/IR+11HnBoKydbqfwIx9waZdOCOqEU5bByqYFmpYawMgRWmamsHCJNJtfek/9x
KsBeN1Bfkq4FVHztA18ha5+DqIzR7aLFRchAUOGFdZFlPtJmCpVPMvT7wmDkKbmnC5aJbZq52joC
kmbxk+MqWg5pHyVfYF5n5znj+19xIkqlDVcL85zakrWagd6IfxS0l3VsjMpT5xQB0LgCvvHgIOth
GKTCG5hBg69aaTqOtJvua2z90gUA/9vVcbvkBVbfnlef4UwaNRoEXgdTXW/6P+8UkQC6bKrYQSjd
Qrjb7R+Iymg2lVVkOWvfw+PPmxqte6setp9EroyFtAKXTUyDvGatUJdzPCj4EUtRcnQI4zpTTsLx
LMEoGUvtRbXpHssBmw6VLf5mUivXAGyHyU93KAzeZyGMWVkm+qmP1bvwzx2ym3yXDguftdOQFsfU
JWedkk9M7O1XnT4dn/QpXuoovdckVX3LpS5fqIPqDQuLZ0UvlrQDTr3GMjRJxjy6/eWyx2CSyHJX
DEP94PdeCj81VASPG0uH9wEv5+CtLaS7PnDKcO0uGc7E4j7sKoM8zBa38NFtgSdvz/xULaQ2FD6K
/hGZkoJ8ULh2Vd2jUOgcuMSFMevzGpldvHRL+RP0ntlW+GzIN+au6SjU1WJCOP0yIVeoC5cS+vzt
1ZmqNeAIXgtB5ahNVQoSb0132BK1yzX3wN1VSPjOVjEwlyKNYZT82xfcUM/17Rj474KhU76EWpNc
V9EGP6WF7VXNIXuBeugsc/xaVnEbpzVtiNbiwaHay8T0gjkT1n+LDdXA+ZM6NH9xjHNIqLytGXxm
Flgvvr3US/RO2aXslXl9sk0zIm7u8tMKOWwVeX06lc48j+/A+g8625b9L1JJ/RBRaheoTDG3sG/I
9xMf2a23fqALVpoFbFap+xFue4AZgOvGGUuEBSpLYyDqTIAPUCsO323CRnYP3iiwGsyzq2rMjOur
JBtGPhOIDckSURFdZX4wBtag+rhgzNvJG5L8JWhtR1xBQmCRmZ7QPX32wEEAD7I8ZQtZW3UripfJ
H58OW42uGJjd2eOF4J4QuPQf1RZxEt0umnLLo9FbDU7S/bAT1WZvzeNhAmn4E2LSohAo0D/rT9Yg
ZXlaFCcaDv4fHloxJqy/1dDwbgVFd1ipqPoRo9NI874TsLIUY3ISeDWLonBD1RTojqZvWyU2vuOX
Uoj8ozWv/P8UGHYwki8jWv5TlVqNYZIs/bp5WiC+Uc4npvF0c3HUQAt+PZmpjQpkpGTPEwGjuYvH
ejdAFmTbXWL4oUEzwyk/WiI+O7S8/3W7UajnXuzqpH8yB8zmCdnLib6OGqptMUadlw22ZSAeGblZ
hMdrb8HcvTh+LG7/VUWmAiLHdh+xu508uEh4H1ii2B6/wZIWJFODz/ix2O3UUvWK6FiDCE77U4Ow
Z87I/86jci9OtAxgv9L12OcZMsafexFEGgoWRD+CpnWsJrFZnzSkx0DyU/MsA+WhQzb6sriG6OJI
W5TkqT+QFPTKfYiMjUKy2GV2BEJFMPrNk8C/AAPThSIWyRbXTUskn9/YUsOC96wRWjn582lceEWB
lDyEdcVKoZc/K/q1wFlQs1J4sUtDeFvOiqakskadCkPKnW+5kaAxUJOyY9If9ndI8cUxB/7hJZ71
11zlAt5T891HcCJZbe5S/w0YLgBvxY6rXCyncsNvKgqY/Nm0y7YiiLn1sHnNZXpqDRZ6hp9xF2vI
rDa9q3lzu8EWU/x6RH100tFmZOp1TcAaNtzGQZ71CX89O/oOsr6CGrJrpA7nXkJn3h3VzWoyYn5z
q+8HAltAaNzggceGiOQg+oPLFJM+nhr0zMUuumgqfM8yxKVpWGGmdNAa+V4THB0Jc0BGOq5OjBZf
HKRHYnjke2aJYZPhtkWoAvNirqRdYBkE6xDRfPVXSSIa22arzZtF4SH+vNB+z6st2Sdnp6ZvG1BK
LxIgBvnUlEp7IQLdGWqXHUa41JbD7wPz1QAgC8np/IB+5ZomCYx4NT3j2jvDz6U3SGwGH7VrmoLM
GX/W1gS9ilAv4emAOukpYoUlXPa9SbNOWNK6KlVK+gfVgPRv9JjN3oJlTsY6oCuAJo8XjahyyUHy
GuBRimOpnjdEnolW0QopMDGBdWfsjJIQSikBF6V1dqR65ADYVI8w6zgXTzB0JWtFegex5mep/W1W
gu7zrxyBcMypt1IamsO6pJ3W/7stHgc82isagaK2jxy3n6h09m4c7hSQ6GzP2NvDJon0QtGRjGf1
G7qdwIFJv8vSp5Q8x8MKfaprVysFvw1wD/kKghFp3XopDJuHtFbEznJ/lq6cgdqqWSsI8rHDhyAa
lrAWyhOZKHRiYVHMQU7Psm3df/TtrBNipvvh5aXO9kuQqqlbUIOF4/v5S+QQiS7jSQfEF6gj+cjv
VEZqyBnq2fxKv83EXfFfbCDk7kMSlh64VH4zO+n/93vfShlM/n2bhuuuopzbV8Va3A9imUeUvN/w
tA5DxPhj0jyb3O/Javjxw5KgXoMB3vLyYkYLdAfMtBlxBG1/iKzB+iypQ1tK4yWtv0l1P6Tl4AfC
h9o0WHY+jMNLnYMDswGEEhnibCbThcCs8WbsjbWTXFqDPVzPbwPKibvVHO9/vCLQJyDJJqmQjJ9u
7O5Hk39sS8hogkSrYEp+UG2oQjO10ns6LzXnyGUlCglgabZCYJ2Yixbb7CO0aDTS394jn7ws+w/q
6L42y+hErIrBjog4gSUZU2ydsJQu58GVDn5XkI8/Zf553lkc1tz0hJi8z80gmTKCdZEQZ2abUFZL
Ft9nAL+RVImkxxOrpKmKJNwGBGSwZpgyZB2+7NtdMXtvZ+wHVivDGK+lIMPpAoCpRn9Sf/IxxGFA
B94WSyL3GxJSeKt3JOu8DaudDUErcJIolrf1QaqsUyvcaZyJxUVqd5dBnyRoyCAFufgKDew6vmaB
fRAP25CAfGQ3chKJ4R5HOK+vGu/IM6hWZk1Hq+LqfIJ2uP1vJFwTHwKeO66LVhjhUL991SgbfTmP
TXTEaUhC/cD74QtQ2OCCmbd2PORXYdMui/TVZzrE6EFf+RxunqDG+kLDz5I60TisK2VegD7Ye/rp
CNBXz/qoHLxTxfoq3UR84EqA9FRjpgKVrHzJKj+AV0A6to7s4tSYggDI+u5vUi9HqtAwq+0QvbUy
kcTjjTtvzP6AmLaL2FU/DIdCroKGUnwSspWHqH8V5Zt3teEbLs3ph9RNK+QL+jT5SY2Mvg5pFp/w
W23GTRzGuTTV6P8Wf+NAdYTDNDSnkVnpWhoMsxgNEElL8XYT3EzY2kXumboo6FI1eyAwfhLaCAWQ
QjB7kWWjj12WdKYzNew6gYI3vSYyCQa7AfKZutfBYnTouAL81M8qOP9gQgkND8y+zQYMteOFcYCe
gLTqv78hujqLQ5QLtKL21Aq/Z60bP3IvJtZj20/poGY2GV4CG0iNP5emy0kNoA/AVbdjUAwr0DWf
oU1d8adsewNjp+I2bka37fbiNUKUw20QXyCsauygeUmNKeZJUvk511KbYqTizlRNxm7MjSQ2Zwlb
ZFFac0lm1dfcHl3G5WWU7+zdEZf6PZkSztPzPqKUAMg86sjAVfHHHobHtc1664svei8yu+C7Jpqt
iKNvYx1x4g3wHd5mGI6UnauGQqb1nKysKlRqagYHB59jPsNgc5RBEreZY3JDQ5TMKu+EwognZaTa
Ga8NNqoIDcz2O5qj3M9lPyb24azj4+banub0jEn0476QoarHOSkMRx4DGsWPF1D5qFtrplnaFv1N
5QKJ//vuL2dPplp6HmlC9vlOYHqOjm2K+XISoor5mvYXs2nft7T3PXoX0JiTvqGraazTyJFAICfh
504S425zVTJUaHmFnzfRiOZczGoRqwO3HygcOfD5m3qWSG6pHUL2YpmeY+zRd19mhUz+7dBW6Ka5
cU15nkXqa5VbGMO8OfKum4/rGt6yXOkh8M99v+ZNiOWsb8LMnIM7b2k0ikA37LGFoacT81gBsGIv
suc+5HkHWomHLsJ+hKkewupkS0+ZYCuFPix95jDVeK9iFFH5mlhAnh1IDe21XRJJJseIAVG7feZm
1yJdgjvbTQb0Qy8Go92W8vU6b9uThkqJSPhESuWjZELc7x1QiAg5UYaSnX1Orl5lVO1VL26ECNJJ
N2J9RYdmjsCr/YGauhqtpklkI9UEY0BmrzQUU6TTOHu/9mkKLXFsegW52GFHM/BsijmGvul+cgr7
j0m/zn5z5c4GO7szAXgNwhEyJHDIpjrK8nDbv1YiZubzxb/WP/5CrTFwqITLGENHxXsj/s/7B21X
sg06dPmGM6rJR1+BAA79LpJ7dfi5TqEDXkkojS9v6iXt0zQ+NNRh3wifQa49zOM/1gsYSKH56Lpb
gaTjEITuK8UhWWzI9iUeXJ7RpkfmYIr8k7yyAdl9gtGHLgHs4L8irxETnMxoxoRkOLt6lFOZqXPO
+MSVRrxyOSCwx6ps+PiABOZYU5GEoBUzh30PavwbUvhPi8V3plunpZFUkNsbHYkWXXlCL6Q4hbaX
RJyAZm9ZfsEdj+N60Aohfd3+ZKk3A7/xzWA5rMY82E+wNHvEeNj7H9GV0GUKTie6tbjdTKBQNa7p
8hAI4fPONrag1hTP3lnUQS32EjzqJqchLqm2gZQqfHnszo+xbBaeiz4Lf3CtfUnja2BO/7VGkvuj
5GLSqi8BfleUxjDaKfyHO3aSjceCWbeuJe4uhp68gIUBDeq7mYifCdCEZ1ZD0fAdSjnfPKm17YtN
zdpelGGl/zPSx7qdPZKGqzDiwMefB09o4MsjqcMEaWFN9MqskTvoZ/N//8Qf3bEO03IoPkUFSQqC
01TuqyaEISSEhC/m8B8jQzIN8eOYZidcTTOfKAB34Y964vXLq5eQ0xKalwIFiURYKF4pyQE3n4lO
F2FDAoqyAzTba2MgCYjmi/kS2Qe6+RXPkVOP4ZlRlYdqBJEVD7ULJ4cOSP3VzEXK31Yc42Yhn/cG
bz+Y99FZF0cssRSM0qulQmjSoSAUr99p7Z/nY22NNwH5yKRbYiPYFVA6EfcvBR4c43kHi5rnzbjv
Blx+uIfpqTmh/8iF9lK3PXMfroX7Jvl+DpHGgaD8WMplhtstQNjpyVfs3JSur2LDwd3KI61Aip+z
uEfNGAFFmhM8p3aj4bFuwvlfES/sQSAocE5sDxeoeg0y8bRUEMHP492JNb4H+tbMdLPk0xkKRa0E
uTKc2STYe2/n9AQic7pIiFKio4mC53dyheKAmoQNlHhG5SX50x46Y0LQjdbNwnRZSsrPBK8qEFsg
q6qMhFU2iWSJxSDY29fEgCKoc1r4oMVHQXykgSyQj8JKv8RqMJhTqHCRBHCOm1w9tPSOpyfGTzD8
3vM72oWJyrVojj2eCl+LrtBgA8qman60U8gVXBgE7PpeXgHZiYtIxGXNJ1Z+h7ubsQazLiu9mNUA
sed0RVPbOY4M566H/FmLuphZ925JFXbCkEjDgF8Q+vmKhxVM9wNRI9XvtwMnLEeghUe//IDsJbx/
1Dy0GrM+vBMXJ4dbE8ihV2r1dW+KGBnnPugkU1Zy9fevW+u+J8nVRC0HJbPAylfn9UMgzfo1uFTE
lWaw6WkOcZUJ31j0Ho9eRjZSJdWmYJCCYmZQGaaNhfKYNkmQjEGtEFOJdQ2ACuXJBORADMYqhG+o
S7Q+D1OwmiJJh2Q8JoeCls0I8trjftCNMhJdHLfn90MyNxrkm1NG3HzHBNKoNqENRJxdqBuOfipR
d+AIVRr/CnxR7IGB/qIzJCj/bjXPoT+bxouKgQvNmp1Um2j0LFF8vdsvm7L+Yf6ZXC88gOoDXXRQ
3as/Ryo2nEb8li0dgiAU0oflqnPbqo9AJr7UgtoM17yc7TxYWF16zScw6iQQZLwsTcrh7eCGnC/G
PHM3cofgZqvG6y1ojg0p/NhBIIseUAl8x5Ckhihny5OEHpRsajwQeaqYHI3Le++vNUhizz7HkmkU
yRJaiUrQh6xNo3BSpdLW/JNUcuI5R7JOGejlYHcSvgRc1RHVSmCoTvUPqfR67Kng8NN7Y2j4gakk
7udjDPlMRqN6c/goZpTYro9IIKSJx1sUgTltJSLai30rcjuD0vqntCiKzCeKOnE3+G9xSlDpwSSY
WvyhTgMqNQLN8Mq7Y6wSBjQjWSsASpnGH3PuqqHSOBgb1K4RAJV4ws4DJOm3Qb4dDUj4ql+jFOCT
kf6poeQNHAhWIUeSF3WQdOVSnJ5l7vLnwYHk+FV6XbmokSTKNibjNrkVy8q4iQ9C194slRdnYfKW
BQkJKu7j472ZMqXdPQLU8a/ec+kDpQBe9CVCx8HmdGDkY/vr+gXzcBKig7U3lP0zPU4YUIYWY6OX
jkmy0xFRJSkylJrs7hVy0KS2r1lj9bkeZTzxVNTKMBATyzQt2qX+3Z+9S8GKIKhy+vlL/IFY1eNY
/1pRxXgqpiw1AlQD8MIw5Y+1C8HT2TR8gxlnwMDS0S16l2wnKqvmgArw81z6TZv43loyvOUmKAXU
ExrWGPvPWJxXiIktEjy3gBulx6x8XUyCL9rJgd9fFOO4R2gn4hog6g8+HkvSc5jHxgTuW0k7F2kS
AMY+kL1pQkZrZ90mGWRXykkWNesIXtdZ+IIDH5useTRvN5LmGVKHQHU3lv6UcWQMeHZjRaz/RVaE
MpQVB8f2cGUfuIoagKSTJNvE5VwuL9rEi25iRxwTjLtDLKWjHGA9yTj/nTc1IU9P9yq13aopIUDx
uPbIVBsG0wNyTI1zQvshm8+rcJQYzsxHUkC8Cy82RoUEJFdhU6lSymUTbR/u8OBC8GhC5pU/2ITZ
4I+L3MTeyhYvbfkc7Eor6wYZNLrYV0thu2colawb884CZSkbAvSNT0+TmcLfOOK1GYdtk3drSqdn
bybztxlB32mt2KWiRTLnAQRId+u+GlU3ESOsQLU0XWuAf06j1LNj+blS+wCuBNsv5jqYLIUUmmhX
DaQrEwqDYlxD0Ruwm9Ic8Es71vehNJLjyMvSE+IeNX1GlRiwt5RZ5SgQ61qgA3X092j66Z/u7PA5
eA3EC89JmiELgmutGSUA3ARIWMst/54wiEaMLx2hX0HgRsggsx0xEPWp90uTXlSRxDL9u9WyKsWr
fo2p7yVByQk97WZzmOtGCHJT2VfqCUgIfBEHtLtiFkszlDk6cb5IzeEmM2uXHL+V6DeDlx/2n9W6
KLOvV2R3MtbJcFWE7DegU1dYVbanHfyODye2u973k58QlQ5ErmHxw2DCp2WKR9EoU/7WgUHINTB1
J1scJcrbLKyCehgcEmjBlO1gISMmrf8h+/1PwuZKdULX6X9ANIlOjlaVYWz16kBb3HzLsevfPvO4
aK5O+DkjQoS7feJvcSIlqbe7nxSvdVtnPQaPECoP9l/YHSfOD7ENCuN7I/levlmQOfZTa8daOje8
DSNu+2+MgOZSAH9qcH7R3nm8f4F240a/AuZccHYI3la9K14O+k4DeKrNdBq3sI2DrKEKNwUwHIbH
vhYvR3PT0Hg4/c+Yl8iIHSFkkVHqRyjD3l5CjZYr93KYy3wPXObK5nZJ2WlNL6Ny4rf0gmJFSwCk
4UW4Pdauoko0maP8t52PFI5J1HO7Gt0Ab7kmDQKpCtf/oQWjt7horbvT+1MYPQtmcrAsrZKZ8v8j
NtK+2UtqWZAR4AaQkRV69AhcS0nTVpTWjAa9XxAxc2d4AqSTAyPxbNEY54tuSG/cpdh4410QDNiV
/20zsq+SoDrG7uhZWWPoVjikKOrKzl/e6GNz+Xfuq87ZGw2A5Ua2CrFNRtuDG5Sso1FeoFLqzocA
61WllmGAyDHyH7tXopXKREHNfteJoo/b8R8M1bL7cGKZpf+ZL3VFxGzn3QIsDXE8IFRAU9IdXSe+
rwEFkeTu3Oqm6u0LWNV6L9FvTh5TTL+NuI4fFhcU1d++3Uhgs+VZmqpQRoKsAQjYokea9uAgfykg
HYD6TO2ehF0la9ZC8KVomOKmBl4x3UPrhHLtGDl1L7Xm0CAXPyVJEvqZSrAWnIxmQPB+KyeamRto
h7DOC58BVuZn4fPk2OW7/NIXfXFcbod3zP43Q0RSgctpbr7K4d1E+MKGbYgl2J3xR8Aww/Rew8SN
CiJflWrks7da+v8ikCK+2GjilGSMTenuB3uEXR/BXnHIiTfLypEnlIhxyMrLkyq0OhmbVFOpkX67
3ZOCtB8n4e+vGxCN3TG5AklCuWRb/6TgdMRwKI0v5EwuTTN2Ckg735wk68A68i2c9d2xp16dUlOa
AMOoel1Y3SMFKoEAeEHZ1FOHexu7TgnUK3RNlTKOIXgmtayoMqNmaf3uP+EE9hl8HT31HQ5sUfOv
aV5oAU9e5zDzhF3fu1Z4CobjOA+OR50R/jhRMbakt33d5h3hRKRR+3xx7seB3yCyV5nc9k6KiPUs
YC0vo1mqRvEwPdOHglg0GauyNqG4YQlby/0RK6gzlnXpNnSpsv9xK2NwNylvWAtDGc2FaOjQPlzw
YCjnwuM/Hbl+WPQHLyuV/RMp7pEqoX8MSE6LQfHlX0mDJyKgG2Qd581q7v4h+/YkdOpwLTdihpx4
z0php8aL5pjk/s9akIRTdRYmlwLQq0NXGZ8+G//dQQM0Q5GUw+QZCgHLnVEbYBjqk8JtxjonMnpy
BiNOOiGlJ5bIPyIPM6Ri1Fr9vjMNQTLyOnE2bIqqzmfGWJjWar5y/54U8tqpOCsEEtYGL3id01WA
NQ3OlJn2nYOp0u+rz9RXleNiBVd2iqyS1Bqb2UrGBvh1Ij0Fnzzgn7xW2Sdmyc9fgkvlRI/bDl9H
bc36/MkZnaCe5ngoA6BjucggcLsHff5m0H54S0Wf09WnHQvafkEY5etkjCeYpJe6AZ0/pv4FyXdU
9wDmMYnGXxlPLSpAuKvK+yAdXD9JKyw+E6D4bF1eOU5gOXqag94z6F9PRaiJZnaH6Ej6NUcOciSZ
GexPAUeN91BBxKHwUeUuyHJtzAKOszQXXZMsLnjmPDWBygrMKGRkaXS+faL2YPSdvn4lU3l2CiyE
fVfv6kvZZt/lA14JCpZcMAamsB1WouCAqyC+zy/MVBN2SCS2uK50uGcQp51T/XX1sW8eJI5T1Frv
t9cb4hDpwTc976Nm1FZsLVGMHGsDScJ7a/hrv+vJmNmIaHta6LEAcP5IIfGFEt4yFw+WssyyDmJm
ZZG4rksgWPWiijaj3oGpsZ8Y0yxqIs6ljxT+tWgzSjmAi+xmiMyk9cTC/GkW0WJzXBU1KD6bdeIi
3H5ZA4RICEBCee8mhIgj/r/wX+ad7y0MOWOJWEYxZljdFFWCYBN76Qi+iNWELOXx04btBnZhKtZ0
wiF6qyJBIRNUHOFUXD4PdF0Xa1tIsJtFN86yejwr2MbXZx+a2dLfjyLZ370uhprseC3QNBsleSeJ
BaPHejc85/QnZlAoa3apqRPhHWerIn3wbQWxqzYS6BGX+qZEsEaH6F1SSHP5awBo2llRwy+YxhQk
a3Rnmodv9Lu47ej1E1YR1uVqgY/LY6N2IEzXABzxu9mRdrPZOCsMneSYW1Ct5CTu7n07M0b/TTnD
gYEelnhJo1NjB8ySdv6eN1tW9SYK5K7UQRhwiqsimA2JJt82givrpcNxBmuaTIEpO91F8Vl9aYzq
jt/uIkfvZ7O+iYtFui5i507ncmgA4G8f5B84n/aDvYbrU5v+pZjLzycT7FAuruS69CYdGix9HwQB
3Zq8l5Mlwqebr486YicSXkkOiD66HILdRfYKPocn3LcA54718qkdYSk+MTFdvWTYVsTTWnXJHOyK
w2xmej0OpVZkamf3mOKHVlBPChPMRgEjQTvUzbI7J4MhHlTdPUjySwmqBMfGkJwwxw3FHMj1c7pz
C12+6rbJrPa04kaBPZPII51yJzbdQ7EQUGpm6ug4oGjob7ounOihUj58WhczKFmCnQHI48ydM70d
xtzWkOR4vChUkDCnpYgiPtlNhc0TM+5dz0XjyqEae+4r4CJrhD+39rQjvsYiLC1ITsK4tKf0id0D
Culys1poM5/T6G1cVk5ahDXCDG6BKsUiE37Vp+mIcdpzSY3PoAFooqj37g6vDRJKsxA+nK6ORg2i
QZUioYxHcRimUpfaF2HOX00/crgw8VVx0Oo+3V3p4tybV0wFDKtdG/Fq0KcnllrLtaytGwRB1SwX
WMmeVVUgODhMwRV/GrHDeXC3wTsk5Bb3RbrO8KllLMdUbeYBrv7n029UcFsZsYBgLZUyUeD/2eHk
+Fm/SleUZ9hqNig3euGxJvPyBWl8xDc9TUrDom0wzMycBD7cCe0GRLzgfFNa66g1AMun57/7S73B
1tygOaCBkSTMw7Qv2VPN473cn80wXqfnx2Jk1kWIHctVpbJruT+I5hujyN02LkIhXrd0p2pXRs1v
Ym5lztbK4UiQP8F0Q+tnBmJD21JJLlmd6sCzfP+yQppn8Z+Wt4iwkNvJr+ycYNwU1xetbpge2p8m
xlNsSyhquCXED+6s9kSYAqIG+f3tG/kttNlbmJg+vuzOuC8q7a3imzRTE30n2nbAw7cTleqWXPCc
tn2HPxUHxhdEn4Fg21HjqvVMMPVXOVDD65Lj3L/bzJ8Aq2NI5NYgCkKNl/q8YufPdJXWbjzbKL+8
j34Tvjvit2Elz0OGbVj8KVk8yxAsjzDrMix3YV0SrWme1iksjDdFyb7UQDWHVUDNfn5nnGqk/hA/
cbW/lf5GfRII1EaMz+/XWC+VVgx7bSC2XcQKgrI/Ey0V4Sx3dNNQuqkA7Xm37wyUQxHnlT6gRqEh
TK8mW4El33koipDY3MIE89AHn2ZY4z+CicG05cm65+vp/Ae/A9IEX01wVpM0PEIPBMGJzsbCtJQi
C5EckgUd64HI8CvCJF18q4mj8Dif1uWsFC+w/qKp7VlVJ3bCoP0ajAGcOxEpAwgTZoyFDo+mb9/b
SeQkhQ4Ie2cjO9R0L/MmOMzwyHJq7odTLyLlkkbYlTjGqfcgjqsvMzr6jUgvB5kU5YYQgrre+J9E
AArSIFdZAkdI5WNVf9YIo0ok7Mp74efanHDsh8WJtwuYiXmDhtFQhhYglLjcr0n1vI8Tt1d/WQNf
COAkyTIkHTS0aJaJsOgVOPoSKL7AEN7hHGaJKFPhyfOHcuIjMSSQtqPLYYX30eOrQnWC0muymTe7
2EzkbH8GgDQVGSPtTxooVklnU7rtYPq3MGQSRy4z4dEb+fH1Aa2CO90dJJeKs7ZHsNi+BF6ZJi3k
Y3qGXfqMr8P11G3aWV62A5+6uO5yvBlAV9+xdilq/pmYhoU1HhCwC4X7A3LHF5xYt7bvc4B85nhN
/kBRv46fYaGrmGSCmdBzpkkwjzaxiBZNjtYV+V/pX1QWdXfr+psdZP9k+skGw0RQw00rjVZMomnQ
+kN3iAqWhialazNq336CrJD07OnfrlUIQkvWwQCjIyZWvAylvHso9NMW7KuwP1FGifxxi2FeceuD
VFHb3gRlhxg+g2sJ7/ehN20j9XXCOcDHVc7n5+Z76Rbo+8+ZVdeARAJdQOjEAxS2FaYkz/oaR6iG
2Y6EoFnZuJ84rWSopBynX9hFKGyoOtAsGc4sEzlB5VPyskgQTImja8R+9tqNZF+ncFkplQAArIme
h23+rvt6IW2coSxVCaw4IV8EMduMM9+XzTs5QqNIKMDbUM6r5l1j4S0FyHDaphGpT6A59iyAzmHv
l7N2uMmOS67AuZQa/12gyj4oxp3dSpLuFiD2dRuh9S5BsXd8awC6yerb7J0AW2g2TNKr67LZ8uGS
XxHyBLX+rumWhlLw4dsVtBwbRU6AMD5WRlnW3nJXASUVeMCfhq5vD90E5LlKtkWn7pioWSSrMLIB
9e1fjcbq/64kTO+OrdSNCQ5CPQprFgcRtU2opF+q7CmG7YC7dWxAIHTvE1BiMDTiiOK/Bjw1br1h
WrymZ+srIw/FE2W/twBo8lse+2JOPYojWYetTAMxn+9X8TFz1ZN7tBQEPpdj9LTpCh1XEEdOIBgy
4jMPUXrJfb8vdnjLUDk3FzUUKhXwOHdysbBOX5o784J4MmByZuxqLDm9nP+d4uSBBXU0vBcDEcQF
7CiRAMZ/I2x5OsVGyvf3syNRifksdCiKovP4xm62jGZME6E52x1FfJ8Z6YV5Zgq6QwtBV9g9i/ZL
uLi4fQHI86+1F2dOnPlCPoajgsp17yPeUiwAJ7NC2HFXj8uf6SDFervjWiNo2wIzPkDgq7oVvfLc
iDmoTDgA4loYGugo96IVPWWQOigekT52zGSDvOW0B3g6DpodciVs02lCtA10EVIEbvbgcqMKmnAM
K9sVfD/6ulfESZYmrc6+OvEeOvGWZltTY7Vc1ggLYrL5Ck4YbMVOGwfjUoA41orKAerERYKGZJFJ
EZ0bhrp3nM4gL5JVBkL4TTtc7qkojOmL1ZY0BtSa04wm1GFsilSo90Iws1AxgSQdXxNxR8zV835a
fHi3gjGOVWQwn3KFX8Fu8gUycFv8M3HmiQmrU4XGsMN6052f4pVC3JFrYTxCh/bvKH9vcy8MdiY+
waLiE56wHG+qi/VCpqcDDRA7RT4VfKskeR7cB+GQEN42Yirer9ZBOBK3K4azEdI4C2SGAmVfqVI/
nJczm5wCir94wHErgG6F+9nkOiq0QHeAjYM19wMl7OCpXeFy6ao36aaEQWYSZ9v+W22svA6w9S0w
pLwgIxgrs+drUXrto6bYyl+IVAyyXEHIfSrcqUjWbl4bKMvqGvGvOfbJLQuHByGEUvvNgFpUuXDG
uhbNxPirKFS6Wqe+kSNNHaS4cej9HbaRI3W1ACWmh1Tjrg3i6sfjeDSf7LRGYuPUUaJT4+4hurfh
wzAYEyQkgMTJrYqK12w4aXUfG7P1kAGLD2zd9RO2rvvYyb3/elAYDVk23XUr/OhhgQDY5FhTXQPp
Aix6UJPpVzA0vvAMXhUDhh2nFZr1DIA6n84NEKVgI+i5LsvGoT4i29MCLI76IisxlmqVUhMozvXI
LUhuUUmgx+DNBJFHK5uKytmIXLYO3sC0fxXGVqychMrlgHtJx3o0NpQBuh1HIX5ckysEOC9ymNv4
P6ELwaHP/3munpAUkSXVWJ9MTVACCQ4vky/t9bC4gVaR+Y+4xriMeywnJqoo4HauBcQeuVlhdQhw
Xi7djIxpmuxoEO3BZ4ipraIHFL+rHQLbXrsmApWvhTmA9YQhTWeOXIsijYC5gQGLIya7JL9K9Mme
mseRRvBw31+ceJOkLW34KMMxR+jAO64QPNsx+nefv19uvOP+rng7FbohkjttyC0lOdnDsI544zKF
q2gZoXmnpb19jZTSP8ejsodmjj1tS3VuU4z66nXjdRbu0qhGzWi3FDBPzP5MnpG/IvE8xG27cWIQ
Vpt4fCtTTXkJIi2ntbyANx5DhiKno8wVVyO5fJ9+/cRRv9CEyGFzrbkjJYTrreYueF52ENft0jlb
QXvIa28L/nTrbP3iFQZIyVxy1Gjo2wz4EAeK9x2eCdHAHTeK+FnyQNPSW/SxagmL4QHZsWTLxn4V
M04BLmnYZ+4VarKUE+Ox1Q8FhXaM7r8NrJ5yxwd7GjI0aokv6MUUUhLo6R/XCFBAoofhl2tX9fWv
O4e+cdBPNdFY+lT2QqUKpeNC5h5sOoSdgQXfTWMCpwiCZrbaZiK08XXKOBqXLyXajbMiVbxkDGWt
YwU9QXjDpLs3tZob/pQGda2/8+KdU1wOY7QWWW4w6sP2LE8xDX4biiBR9oZh56CmO8Uy2Y29oP7W
tn451xbQ80KWQnwKgGI2qsMh6qg171jnkR4dG5HDYiC+ym1qKKoS0P1bk7y9s9TORuw7Ahc9yZ5O
u4SqUTO3MFDwqBwiCK3xIWehqzUDW6ZXHmQdyoZyOi1mxrVQPtla51oy5mvhIMiBWPdwzio4aJAX
QS5EsvxW92Dy192KzJFXqlVIeDtff8B18juXUuzcVn9piJOIwHgZoj1BLMHOThqtCnGrO3CNnXsn
kLBMp9PH2qf5jvdbe/YVa2fBwBW6KleA4qEIk6Ib9BCNY+Nd0w0yE19497aRF/bZln2m3mQY1riI
/hEs4dLLtxBmU78uvXOLuCriHW4gD4E2T7FNU8zMLfkCDhmj/2sIfqauSrl9XPXuRLZ8VjM8VLnK
wIAJR4u3AfRv+AkJz0OCacAUGsvjnuAqJKEjO4hLYOfdARPuYw34U8+Y0xW2hPnbBuWubeX8XkLw
bjSqHA1cBX+KN6DwXQsp0fQREy4XT1CS+1FP+BNDxOdFVnQrbTb+OZUVPMP6YAjwOqP2av4gkrlL
CPl1hRq/VAQ4xbibaFqcSROfa3fQ3h0dOKbfalTWH1ltG3W64GTv03i8vqmZNDgaQZwTaYm8KTHD
BI8dWVKChpa3Y9HXDgyqXn0bT+CGXRZX90er7VNXIZphci/j+WnPF6NgUEp03/MrVxSBAgDvXahN
/uAjtaNZnxhnkNsyrJaV55D+NrdJI3Wwfa/5OhCiYu1w4bH8VRtfJJn203vmKjO17Do7kt+hiQdf
nGMTS0LhEbmLLTF483BWkYp08ZnXhzOXXpGfaiXG1aywdGw91k6T96jTsVZaaToqHrzv4605JJUl
eYJhsJOaPcG96cwgHa1u99QnXKj0TohDoUSaEY4wYsbgCfgbRRxNpF8sb40O33Cz78azLkFLIA+3
+qPK7TgIY9QpcAjNEZuqG7eJtHpNG7c1xmI9e3sW5CH5NOp4G9vBOTVmaqpf8OJKb22ygxXRkuAq
zBT3K7cDyUm7Bs977/3WLm+wEnFdJ9WOa2JAicOHCyMPwG8jU5+9st+nXmtqoHFcbW4rGxSFb00E
ZOt33iJrymb6DxFa53Uo4pQRW1p25JxCGNy9QGWE0WB2mTDBkQg4/eKrvZP9sVcHypQWYeM0qkMC
e4fDEfacFGwqwPlZ0iB78dXekUsd+WdkkNKMmVoEt2XKbWZc1MDCtxvJM6iKs22g77sL1S20mJf7
CnFzdF5N2WSwyUm4JiVcd4/UNN++KiH9dFdZlzT4ZA5rKS81WKe59XtiOUoCBOSv3/9jzMGIouzl
K8eP3gJ5+w3N/W3ir6f6n0lK3RWlhlxfRELtO34Jb0Jj9jQDoVGG1oxL71cBLZxl8f3rJXP6wdfp
oGo+Xw/uu99cnKAVLNILj5bYJQWBXf+x1px9Fg+aXxLlRJk+cStH3hVsoxIwv0SP9UWXbYOXoZV5
fmGrFEWuY7IyLeItUx/Im9RDaEyRfNBNpeX0xTxs7O3lyALBPGrjS/nYtSzbQB/guSVz0DTOD5eZ
xw0wcXKhcHIHKLNvpaHbetZ1XxCcPMX22aXS9FEP8eNDuZBQWfcYFI+DnNw3f39NsmdZkFSCuuWM
igl8RYYtnUbPXb3nPfbaUt0XbSq2DaXiQjze7cxMci+9FsRa2CKwYn0+hgokWyoSaVcC8cE5K6PJ
sIuFYO3AMmHN4GWSLbGco6njvPGUrOEh1lDp3+typP+UGiXUv4HG01UkfHfqVvpHtF5ZHISnXq2R
CMW39BB0beHMXm1kGhwvmQC/lKsccxHUCGnTAM0hYwBsgTyUGFRrVJljT1yF8gLCWiOniPL6DctM
3sUXJYQj3p+zONWsvVa7sGtSsBekyYldr3LGTgZCJHYOkAIAE9QATAbJUTFex/tjxH2a385lOj9/
o7j21x6+1qqfrlEMNiP0u1009daEcNE6eiSMIx4PKsHBcdE5JeregrH3uEfnRrl/PlqlgVeW26WR
9BBFyR73M+mwdmjhV6pCnLlrZaU6+lSWkL5ZpCVPoDN3jQvxKTPohAaP1psPSQDRXsdMqcUuCJVT
FSq1DPeV/QLe83oPM5UDAbTMcc6vVsd+i4a+M1hsE2YN2U2ANrsxnsOGxeihyqAO52x6ZjSRrTBl
GgRENjEZoS6MtfqHZHgh0e9e8tnsdZflQxLJsbmKXRoUVGHlZpeyRKCGbdk0nIlbV7TDbPp0fZ3G
qpnnyRKGJ1g/txcTEQ3dL7VJ63mfdX6NHhuiDpVeIFRb2bFqFQjDH3D8YhwDYxPEtg4TnF0Qr6rk
a/OyhLetVW+SnJQfrZqjq0K/KowATurnUF3BY6wki3NfD1KW4WKu0nZfEoxBX+aanR4Rya0+trlo
zH7qQ4OyH+ko07S1EYik1LGnDItW1UDxwRwiVx8wt8sis8fZ/oY05eGtShFFHx9r1KWwQsgCEd3w
UAJUOQfCyBMve+EhaiFsXpWasY+gdu9cAETSMyP5WmTCRz7eGtFOATop3LiDz9dRPOts4eD6xgCZ
/HcG2Cao0eSs9uZJLg+h1aVCcoE2MseUPnTydJuwun1N1X5gqIixaMmbEnvDcgFhvFT/CHYvLiTu
vcgNoZnt6gqeOW2bdVLtWqt/GngxLTjoKNZ++7PaVJGvEVFePDOra/j1GjJPbRWLw7J6R1411b6W
aqRQYs3tDnwcSSyJ1DtPiO1WXq7OTLhBbiRfDOB/7DH9SnTo4lSIqGcmJ3zh0TkDoRlX0LNDfy10
HTP/vczPehbjuzGsKAijQyQja6vjojhuZKJS0f2mSvgJYMSXGNX4u6kb5vGUTOimygsMkqW/c6Jn
HWuaiEsRKPGU0AjQ03R3GcgfiLV9hWnjAdL745ENawui5CbXJ5Z4zMKjWTpICtzWQBR3ZfF/P3UY
JiqydW6LEXOR9JKX+sdcB6eQrZeFgDCjIUUxYnX57iNabYn7Fl5cblB5imY4yl45WlLzDLE+tTVJ
B5om/CNQf38CLjOYeBzxfHkIoCaB+DxJpjjYksfFVwynGL3uPaJOaSoiDg9yPZf6tg+7Tk742/be
ThVBbDsWqcdz0xxc0SmjyohcE6IeSy3vIwwwM6SOzDZGyYeitD0MBB2S4K3XK3JWB4Lb4qJtCBU5
8TaR74qtEgQ+EGZEgzNOQPWPScivzEnAOM/8ZETJ79keqG7smYVFRluNoL//KsZvlrW5Csd4pRfi
4v7LX/Rnj+Bs9Faav6URS24/ms5FJhsmadVtAI9y3lBrcjTQthFlECeN4uk9k62gQHqMGPxnwv3y
HoS7fhQQLnJWlf8bQ8gpoCYW7bpdy3jHxq5ekLv/QgTUu+C4sgrJj/mUeAp1rXgvMVsmutV9/7Qr
h1diTbLE06ZZOnnukgNWh7XF97EGcLfG2l1BNaKl2rWAZwK7RCNdmksTMiiHbiD0Lge05ZNNX95g
IVsmcIJG9WC9EpoohANa/mOuJ3d8flQ7yrdyEqJ2/B80Xt//zD4j3Rq+0cjR749BGFDRwWnIPgiG
squSnPpRzC8K9B1ogcyypmuZpAIbKz4p6V8bJxLrI9xC0VCt6ZsSaIZVdKX6cBPj9sIMqziUQw90
XJ6Ai9IEXwHknaJVUG1Rt+OQWyoMQi2KohfNscwzZG+dSEHisZWVdt8lH7lNi9K3HdbKYmfizuYj
RVSSuhrXpkmXentAp/dan0kdthnVu61qr0LJ2425ep5WDK+xAsqkn6+28r2UT5td3K5SpCPzDmRL
+OT2KCr4z3X7F4qKRtLlB6Bl6xSTGm8XjeDkAj3z7rKTxfT74U1diOnfkEGwA6QMJWcRiIBzAhoD
x+7DebCFxx6y2kKhWqygIPVKe95go+Loqws9/7mlwtii3rcQtKHx3kj5QPIc6L/Q382OQ+gUfe4R
SRM4q+tuj02mBPBp/l/b9hhV+2eh9J0BGxY0A34GHp1ZDeSCNOV8uehCFvGO8Ps3p5L62A+YGl3N
N8vTXPA/7euCQPidVHUrc0OS9T+MC5fINMVdrLQRruGTpktJRxLY4l3aiTocmb76vbg/QGTZm8Jr
8s3z8M2hu6fRW73/U+2iYyAxiNXX65CTvUdOiCsWpvhzwpcHAvzysfR9RbfbiZKMM/kyveRKCaln
KGTliy4TQcZPDx694PdFkiAd0B08aS/8mSISj/EZKXIbHJiCiB7e5ak9B4BUMjoC2jDIQzrpurWl
pCNmOF5FyiT4XeuhWDkWoFKTzRnY2kJja1T70fkZmmyWvezdNLKm2VimOIcAmrsJhJAUyc3IvoZy
0+9kSplibKeVzyXsrUOj41tiV+D+r7g/TT3AXACWWMnrARkpKfzinFiy8kJdgk1QAYPuRvNCpp1e
PW96O9MtcI+haLxdfKens1wRlhBJF164PzF1QmCrorngZ8+5i6zo0TQUpELSLe4xI5eIBxSyJ2kw
8XceUKyP7Oe86hZj+DIE5AQzLFFO3DCqZ7xOg8r1zLNYO7M3aR9PbKGONj6PUW3SbFH3CAx6tTS3
gxxOnKU8U7dZSKk1c6nF+FKQYP75C2Fs56jJU7+G6g7lWFSlJ8XoW95lTxvLcbUmsHfNocj6XcWi
BHLMGgb9kXxawO4PK7Z8kYdWTHlzpuPclTqUkKX0cIsutkxsSPAJ6O2lnLhMgiWPccXdKdqhx6Ns
FYi3pzX+QWBA/cSxrgn5UIiQ0q2Riu57GSlJTXQ+sX5bMAwkNAEguhN09hlvGZJqSo7QU84jfIAS
Un+L+sn4ME2eu6ZSSmzCXZTLxjT3Q7QBqlTHeSWwYk8yFEhWIURi/Avj9HmObZbK9FGmmEhrdoxE
lmKgN2LRqB28/16yM7PhpTppIh/VSV+1tUEUWdGlD4OCwY3Br1EXDql6IhGHeGc+KQ2MHQuFftxM
JnQFfAlUsvdbluZk3GxHwoAEynh1ZagTfp7RwSTFZt37ASxR7EUUiNmaDfZMAh23b1aDscxK0wC7
ICGLYGhRi6wosc5U6wv6MB6zJOosxX7nvYM39gQUCfaJsFyNj6at+YTaSGtVa9+gZWV9uCQYa/Bq
XcG20fKSK7CoG63hVkF+alOLLxzDp9Y8SmuDlBoQz/pvnl+0QRc3F83dGYVNe8e20n0tA61bPoLb
9qUb3DVE2+aMdyS3RastjhvXb2S0cNk17YGQUDjNYecV3aOaAo32CdGOajTqWA3680GpWrWPqn4c
M82X4lwhNOXFfi3G1JHPmSw0EySvyNxmVk0aRcIT38Ty1dlkgzwQU3IBbFxfqf9rIEjwyVqDayo6
bRwPAsAHxS1McoV51Mn53OSFDjBzu4AYAeEPbGjwVZLfXo10YsmtFGi1jXywxWqw9kZN8mz+l0OL
Ro2AgGDtOclnCIjKRd4UlZkjZwJhakAgK3Yhs7RZ5If7mFI9c89xM9HokOwHZJKUTpTIEKCOFo3J
tky9UH0xFOt8SXICZkj6jwTjC2d34ep9bdc10xeAB6ZTS53i7KTJv1BAFJ9eyavQmkCGbae8FI/k
k59nm0FLJkTFkPnWKBbUPGjfait5afn3CPoEY3OHVQUEvwgsild93TB+bbozkRdLzTnwamZkrSai
zMegd60wc0gsxf+nG9XWajosswrYhN6D0cNb00sLYJlbyG0GcV2mT0/ymDa9g9Ux5dDPysN4jPNO
WBzPSGWvyDPAAlGWJ2Lj9/wNuM5cdsQbbijQ3LuyGYXYEjmjEBzKMiPGq++vDH9Mg5IcFLM7Mub/
O7TrGawDKM8jIbx4JsmbD7sx3JuTrwG+o7zHbOcmyAVS4uzOm23YQh7CYF+4g1g2tyINlo/FlgYI
ay+5JSDFbNe9DZG7xRBGw+GNVmcMCtEY1/XZqWkpR4Dq91TYFgjiGbTfxH394HaTkiPMNUNsZCEW
vQvq92Re5lN9BbeIocNYN21e+XH5XPc84iGr38UKTEatkRvJBTO6E/7cWZgupraCZ5+cf5bjRh3R
NTBq4bR59JuJb9uqxBJCipUMCke8cgOGdzB81md+zuyHnI0C9heSrXiNapespBFy4SvCj0Xo1pYp
DI+t3nYxVPXAraRTQAD6mu8UyrhPboND0L0zuEjpqqel3cTsWaXdyTqcxEFpNR9KwGTNFjPJQmW7
F3LoJrzZeiecfee4TXX6xktCg9aAKfyRQ7K0hw1xfcc/cl5oEDcXma3iln418i2okmrPOEL8qpR8
mLyzBAsjt/jIn6tmgMNWgta/9YpfRTQNSWM8IKeRqeEeYjRL65BAOzJpy+9HPcNH+TA6GdaeOkW3
7imDTo9vXZjgBToZ+kovvxeOCsZyBZbq+y7G8tmaN6RjQvJa+o8mzQw+1wELNKRcTj5yyd81CTo9
s30Yj6p//7eqY4zYN7t8YjKbsogo07NyGkE16eGOI7Xz7qfGzukTSughDzuU4dw17Eb/ex6vD17D
23lKTqzvID+akguSmD1Bzz9NfpNpzmIYjEMiLRXQThs2aMmYUjyLnTVwd6+kkssumaBGen73oYm4
VEbN08HQUgeCkN1S4K0A9b3gZfDS86hSfyssbiilTfD4/pGgoEwqNofU4hkq5Jxx/3kmX0ZO1uzX
JsFk28XEwZ6PckYMV1pYbY9O8yqZT/GJtEs4jArM/D8GtOlEwYOIOjaWvNcs/lyv0RAxbHJMm5za
GNhbmvZNkTjeh4v539ZpuKRnj6fIkJV2P5jOo0o26ePlu/hpsNCdwzpDggQjo0gVHmkuKdK/kaP/
x5fmmoksEm/WyWKfit5wJVKFs2/Nkyxit6fn+tnh5q+3CgPVMkR0uE/O/kI+G7fXSrmyWZq5IYoy
1Z6mvM0g1DAZJPbWG0fH47R6QDpDUd9K6BHQz2Qs4/zYVY4zpiIVJgv3Q95aEd7ryAG+4S/STxDf
6kEkDbQMRLBTSyS1EKIOgUsanKLOQiZcTs3KB5NzSZKVrznZ4fVi4AcFd8kOZAlQNnhrQBe3yJuj
6ZVBxLHmuqcAeM1mee/WebP4OCZhkTj0lTNgJw4MQUfaI8ZDGGQCJ5aV4dGmi9t2TPr4i5kxC4dM
w7nRIb5DhfoprA74nK8zbXggk1corwCvSj8YKMvcqw6HSbr408NCckuOnv/VqTf1coXUTSo0qBNM
k7FiHlQtkjJLNDkD7nLhWooFq4I4z51egj8s7nIfYRa1QfgkB3edNkxyWUGYybQih3+dwoaI/uav
FsExqXxBufK/XIbG/wdgdIB0PlqWOoqN4GGZ9pqzqP036DE78/19euwegAt1ugT9bmgQrId5q8a/
0mo7mFnAJyUBvanE/GinpNGwHl9ld9OBOBftDXkyn/JdXzIx9pkAjWNtvFNgOYz9nm4/dx2mt645
5Z2bwcTAN5IDG/AgjQyoyQorNUS3nfy/U+vztOxlRGsz7CQq4rRCWJJMLfdVJBOE/wDVt/cmb5mA
Pa/YHI66jNvSWPkpSJBOCYexS+DXA6gRAcaMHGJ12FBB2t86wf7VbU5PCGadHwjUIP9Y1lRTjO3I
c7ZfO4tH60R1htjkgZBQIQ7RArtTgb6fej0tdPGONNsBwMrNVC5CvkNPVdePsftuqG1KQt5+9H8H
IvfOjBazSQWNFc5Mtau4nTUoihI/y302Gh6DBTwjZH8T6krNGr2gLQQkD+MEVPiQ6L63mohEb3Ug
zs5yvvbkaLAWknwl8NENkCCb0Rbi6CQyoaL2HANsPsB00DV3qZmhgPg1HneB0bbCEp5VtRQBm53h
OiEkNtn4cMaEqYOOoUx2aMPsXEMyD6Yv8RXAk1DmddrowHd9oqcegO3ofusQptZMdHEa2Jpj3/jY
ag5MPtGxp4253T+CROrYSec8UObYQFwu4iuKoO0i+WGYxwyk7nZLak6MRUv4n7XuIJneGat6v5uy
QPx4ZE3CEdlFDTtzgJB4/+uj12QrvROtg8xGqfoyOvqKS+1cIEJKp9w6us+l9MsEmW1qCfdJqn6k
S8bXVPflDKbONxm1GcbP+3+4bBUDi9/Dyjbc+n1mw/d3OjK8yyTQy1Ly+G4ZZHwnauseg+unmVVg
ASeHZkFLDyYfWF1zHLgx4uNctgKHbkjqzZNj36YTsQXw+V9YR3LPbV4E4XzRPvDFB7wPC/9zGRtM
pmSj/hLbOGaxEWio8W0gbeeFfc23DHtG7ZPHDWS4TIfLXGd6M16tBDXSfPKpFwao0Lg7hvyidAAW
9VVp9Revmqq1m1DxO9+79TyQVRFL6EgWSxY7HyfR89KgUX08sbf80HwIjJY0F3kSQnLSOYK5psvx
5ud7J78eYH9+FEnCYa8PFnLfkMWtLGq3iUVWlEMX1d0nfP8L+kTstAc/1VfPHbqM9KMwDoe8puJ1
O0YsngLlVP0CmDQSUbFiGwn8tfwXweiID4OYSSea3fEU49/bY9PVB+HBhmzGCfneDcVbaT9v7LsV
axwV+L6AeEg1vgS3zyt7UDoDQFGLpsj644ZyKXQH9IFvpQqYJaxilpxbTxGzVK5oJ01xnGl6foKX
y8uvz4g9rSXlpd6zE1WMSZbf6qVGbn5SNaGCzMhbE9a26UYXeoEG8drXYV9/9+cu8s+WrxHTPnTl
tlezHL/vgKr9yIEz6dHw2t7/g7zZ35LTZCFhOuT0YHpQVeXybDuhQ/WOeoYmG/d7YXrhmgJ80xzu
BcMVS7JhBpmK0xMxCs4Zji+bI5X0QsezdeG7jgFPoGXC16lc4/IAuE1guQIM1M0oa8AZFDSaz2M9
cB/0OZr6XHhSc1yaFwqlN81YmJazWXKV8/kiDaxSPH+AKNYs83At7WEHvoSUhLTokVLhoWxInOKt
8Hsd40Y9TSktuOpA+5XZaH5ahATB592jwDgQ1gvO9TJh1+7wBg6Nzs7ykJ5CuGPkcM5JQSECZ/CM
kUtyd/dONvgWAreQR0j2wF9DWJrRUpP8cv1qTw1ArHz8X4ftN9JUF7qdyxYV88xT+Irn5JTFrCl1
grQIFyMgz7ZjJkEUgr5xb3LyYHoQOwrNHySsuNzKTgl2L65PWsNfmc/APlA94ACrLhCj3EtRUD1k
u6WR9tumrYqUYdGopasGDVtr5DZVkP5gIwK3iialAwHLgudyHpns2K7q/Rb3THkVVQALvhTZmM+P
OWZABhdEhK8w3Fg4Nd+5/+G7jyhZfTNz88oS0/bvds189l+kVGQAJt8FoN/bN6vnXY0R60hP+Z6S
sI/O46jLB0Uk05SYlBnhYE9xwinE6qG+4CytQajuLYCRu+QLcSocCE9c3bb5XhlHEUKpp3mIkLbN
e6xXPB4VIoE3BS+QP+SvnNkKdLf8PInL2+XrXV/FZuS5G1BURbYhwGGNyx5qkZiVqfjsSXKeSQMG
ozXw/PRdcYrvhUPLBhGLdYgXd4pouDPI/0OGoxkGJLqEztbDfDZa3tGscbtpjS0BfuJO/CcXn5Jl
RnIts805acP9ZbGMJTEyoRlp4N+VZk0bhzqKs/tEJt7SDg8qYx7RHr38os6LiUJAWRI9Jj8/THcP
eQC6mQt8CdQ4yHQ4Y0Ny2GwrLtb3MjiP7uMwPn7etr+3YmEUkqu6Gg7uwOSvzYNpqjmPHQ0Dywwq
SeiQ9dVnL9RvwvO+WPRy5DjHeHtgO/h+D+8+hoLk4uHa4E0u9FLcNTktlKFlg+g2bJiUlYboSXYc
8ObBKBiMGRUOXTuaJAXcoQCOy1VohPgTZJmfg3PljpriCWPHXOWHw7L09eMDrUUrN2nVwifZYtsd
iWqeDFQG3GH7jau0h1xwzAPyMla6wW6SU0x4o1dE7NORoOsVw0POp50/Kj88BirRAJTRgNUgNFA1
im2K8pn+qlyu4/DSEtld4CJQSxlm+L2BlDmPwutESabig2SFkltGHKSG6NFgdHGYUJT2zQSQ2fa5
iQTik1nqHdR+I0tNUr4RwFm05yR/MMEEeaikkzt4Od+kVt3+ro2Ty8kGksJlE6BtDwqKLCWq5gcn
shkrmfv3nKFmHRVRQfDfUZoyOAGvk/TNBLYm3ed3W3tCcaTSVcKyjkaPjmznLjILr9qSbwa7Ohx1
S47SRU1gPYiFgM8/2qerleC7RNy1wUPoo595cl4Jc7RD4c+hahodFfPuIKfCEO4dzTXCfIZOh+BM
p8rS2cuwVloiJCNVVvWiSIGXRWGaLNG0/D3ut/WHQgTdsULvhjjktsmALzGyn3Z5pHoI8Gt2kZ0L
hCBFx0qyP3Xf99BORfkFHSw2AFd2t4RYa1waSk2BaPQUsmirjbKgSLiNiT2xQghPe++W4pw5Lrdv
jfT/19NJJLbCcznr6tJT+xwU0qAVbGi0fNUkrvjjSDiOSTFa9+Aj5LqIGCwyz+yVvPOGj0kSFzIm
B+jCFPPb1hRAnxWKEOWgOFqL7/8HJJsThXr8ZH2BvqKCoc8CaKTQVL6xSwajefiV69JQ9xaaVKAQ
AsFFQsKmVQHCKjui03U82pjVZ4Oaa3khLwE3TaQ+4zH3hY0GFTQy+AA7+sMqRVRl2Xz99ecDGgHf
CK+3j3U1Css6EF8UQJvaC/n2heDDA8Kjz69/3ImqGFyxXHMFzZnAthJdqC0mgfKBGKfJ1HZFc/uA
rREjf5oktrRaeUemrQs/PsIeVpCyMB3duDa4AYh4Ypmog95JSuRANINPjg6XdS/qHbXwIL0UAJfO
3fOZyfXSzUttG3WPUa2m0TC57Vy8tIxmuUPmav3oOZ5XKuDDdPEOuzOxUas5arKsNFs4ENAbbi+d
0OTKykJ88MhhDnFCffzaiHtZtUDuMJz6btw+jY+e7FGy++hGGT3RMsXrhmAiUaEXpi6dgM6Umyg0
8HSopo/oFcyjPH9fyedRZmC0RcvMtqK9jqYneKkk5/tXdTa0zh1876CvGZtG7sRm4tOhQe/hNCBh
gwPmKo5gyNTpnGoSPJsjlGOmhViRyIFBYyNkbkFI4oDN5yF0dPGPMferMLKTeN7k3l0fFd+NzdQl
Ccng8xI8MbwNDPQgg7KWtglUyBuojAWzxfLqINnasn0qxM2VQrCgDcg3WPzzphwm4uLLQ9XGwBTQ
OT3bF+ubHPPbU+5r/0cJDfIQNPv8cRa6n/FDRy4DxV7jvolMGl3jQlsF1sXyjCDY+gVSsQx0aPKq
HR5nFottI2cRI7gT442ok+ctc2ZG/9xlcLV6HJyJ6/pOcXckBFc8EACZO2thiwu1CLwY78wTV1Rt
9HtOiy0Kg64pq9rNAfHUmPWTpgaoSVT9uUySqcPqMsNIPVgb8J03yjVG7K+V2NLGlW4LtreMCdEX
1TZEOfa6LuRXR2/QvrXitkcFC+IWd4Sc3ulN/BSVm34CyWDwTIsPZByCSDJLb8ezRMHlkY96TP+O
a+rmS4lAbyob9Wv/ln7xu9Bf0AnrtFi35BuESam2aWWtPVrmxeDqBvRV6mbfMdUTVVZx2ZMQZZJF
h7VEuEX6VSsP4wQK+fpzKZRTF1bu6fbH1ep9cTXndzRkBBmytbRJH53wWBnUY9jpwfoJt86wImG0
JELtyN1b5LHuLqPU1lqs9CAWw8No7A5MLj60eluN5Ubu+8Yb0uQxuZfdVk8qWXgvTT6TYb4WdbyH
gcdo8tTHSvmU53q2+Ro/ZVLK8jsVOoS7u4vzJgcgeVQuwKCO19ElB0Npahx9W+9XLvJY4HO9hDLh
7/eKD90uFCZtTP7jOms4c0cTBpmkiW7TdVWux19zgWL+q9OteY3z1n6T6CJ8dVG+I4dCK4ozQe15
OzVw6ySEc4uB8mkwLccIHhhY0h/qWb99u6WOWfx7odq8M2cxh7lBtMxi6Qxx7bSmZZoQhHbOJE7r
nIatOGEZxa99fS7YyjANaedIvuC2l/CdJI2wewqRe8rllZMgi/UyXGtyALYUNLEVoqoJogtSD2Dc
04PeU/Oe7olZcIEAE0Jty4KFQ73oGUoc7SXvWK8wvTW4/H9ZjWthSH0eJ0uC8yTBRnVA0CkMbP56
kZxfAsMFLZDmThH70sDDPvWjKnLLZrNqTFHaFucIR7XxWmfNYuZSIDajD3lQMygCG9WdTVYNomhr
oc5MFip17pUm3kNTwj5qzv0G1xN88IMHxx5C7LbE5iT84OqeFk2utDuWfiC954WiiU0Gpd3AKcLC
CfJJ4ScWvnwF8mLPh60JkpBenf6cYPzsy1GbDK/RobvBlzZ8873S56/oFam4Rih6LOY+snAfXU3I
0tv7CK6Csx0BdAhxTAdc3As8gkFyjPBv2+twVgMCpi96y9Zos99p+fB8+WTDQ9q6pBaMozKe2YEA
0AxG314gWsMvDAoktUWGnUwwGAIsGNeuVB2ib32437oY9BUdXlokmwemXqcYt1DfGhNLQgVvJ0/e
OdxgMYTh+RatCjxHEzxbH5fL62PnB0NmsT0t2l/93Lo3+h7NJl7wMLLDVrD26dkfftV9vtucprIZ
AXdHKA8w9I+q+mrIGAGzvdF9xlkKXrcBmkPDChPeiQ+4dFNk+wPdZhvgYh3nFEBaolbz4vXZB+Gp
SbHVpBconAtCbFl/suk0qq8JMljxdVyWAF5YD3sQ0bdiwEuXVkeLhHaE4AsffS4FBnFqrWaoPpvI
aUcw01FlEiYHTYLGd97bw/zbZEjdgz0cftvMON1P5YpwVPPYRnNVzdbG4TtT8UEk8fAj2C7Ozuar
FaFwPnwExFyf35+9J+oz32QL54caYhLElIdWVHxfccf4iy0M3cMIo0UDMDM1CiXKWWo/PpHzF56K
SjFajU8kSVkNNxoyP3GL/hMJ4BbjfCXwU60MjfdelpeZViKvd4bDPKOGDBBHX1T82JS70lbzynGq
BfLJxhT4E+3Kdb1k+jgAIIJUZCAd9DOI1pINavJmX+FUbdiIrLl7yktR2EpEqjvEc+hDipTVkWcF
eG1oZMjCc76pMeFTTB+KcL7eyzWBdNS6wcZU0BxWTlGd0c+vqVm6+HviqhYqmIFYVAtBi22bya7a
NYhhMRXyfBLfwAf9JzvVgN8Zi3rzPQxObbjCbuwP1YGJeaJ7J5CQu8s0dAtselwCqkZ3ieLwnwWS
0haKsAOCrHOuZyM1BIG77zMlUuRpq1roIQt89WaS/YhImUHqc69qW/nKb9/uCyd8cLQikGLES/ZM
XKzvWBqRkFZuY9R3y92akRb7MxbwopuKlZTN2Q2AMrRH+DL1CCDQYuH/toNcchraCJexUxAAYZlL
Lej9iZSAqQoiGhrxwL7EnDAkK7GQsYvrFMu7DDH2jFp2EY3e7McstBbulbzZTHvLy4l/fI/29dmg
BpaHnwb9swBy+xLvc6iB46WCZJBgOqC4sDaDA5GixtTakg9RVaA9uJsxE3UooQZ3Mxiso5BAfaeu
rv9zOr5MGJljX22zyGUWt4Lbmgak3p9N2vVQnOGBMKYCDGvoJHFbwTTVDqyXePBQpq1wHSxvZvg6
02ffZiRsmUCWxMaUn0uhtRfnaDmxKq5zWuTruLQmgrDV8ofVxTO5Z+1vEaMgjZ/LGSj9BlsilVKo
PlCDKZxO0Fy5TNw9MDe7uvC3rCgurD9rUwG1psLVcjxyitafRT/aZZBcMPluhsfFZpsc6N9W24rx
Ph7tTkvcTWa4wA179aB8n3zs6CACih9nDPJxj7EanHXHCI6p4DTGKE5dFf2+Z8wMCsRdMgX5/tNH
6Kky+5TyD312vqoJK1vz4LK5MmvnYnLG8kJDaYq5R7Cz17+yLN4vTfoisiMB6IbVlhn2x9EcPkrc
lKzEvc5F0eiXEazSJogvFvEqAPhjX/kjb4mDpNt2tfRoflsSgXmppvLnm4ShASAX7P7G5FzLYN5r
39X3bgRVlFeOnNIguhmn+Ad+WrftxYF8Z2bx2yEXIgGwRx0OypGmwUoAV5G5VwLu9R9bq86V3gJx
sQ2HQIoSc/702N80GN6GHM5P04jwm4KgzsGxmPTSJB1513GIkxRurljlhcZX3Rf7e3nisywJIlwz
uKIK26D742mMUSVYXxI6N+nuw3c9uku2sZ11YQeO2Oc3UwRr79ILN2k/Ajw9Z0+rdyNguY1b4GKV
+xkMc2jDT6QrtP+if0qmmTL/2uic5knbS6Un2yUztaYpsXFrTAEvFiYZbUbO0Hf+60OwAQ9v9hx5
ckhqLZ6RaJ6p7mYPFPOWULI6G8kKshHVbUbCcQMjRQGarih/vW2lW/Hv0csTTOAsAOfEvlhcZhBE
1LJLNdkxSyyKYJswuv/WI+TSEXqUxSPyoOOV5d8QXcUMfTdB6YC0MB7VMs5J0kZLBwCQWGOwyiDo
jTl9VVMdlEZQxhaOYXXPKRqfQFPtUZPW4/pricYxRJhEkVgX/UP9AxgZWlirG8LrFAg2jkspSVcS
enzRKfh8VBHSZg/PPkz92XR6ZhxFAVv0TKXFp5W81EsaeX75XAIFw8wUKXPyEb9H3s8LMjUO8yo9
ctfZHFYI4exw/hnwiR1czEBuB0+s5O7O8cm/w8gTTPlaZ5eEug+aUCayPC1Xv/ebIHI4m/yITfu3
m3VOJhJP/ebfHJY0LF9pcJGQTcXahOFWcyZeKq1vN7kuW5y5jaMLk5f1gPY9mYKGu4mv/pm8LrVZ
b7+Q/MDMFyCWkPuQ0nyHFgEgKHLkCozlxGtuAT1kw2wK1ehmDbZ2zpBLJjLA3L7uqinwyRChgemb
VIba4HKml+iysy/CcPtPHnlXseuN+cBC6tAODH3KjygqAEgcLTQUXRmkKnLIgb1KcNg/67Go9fF5
icK+I4DLOKcSah6c8xY4EDyjArQlNa11ihwlwVYsCTIhMcdrPmFxGFiyn3D0ZiywtnRpXT6fLNd8
V6WPjNpmRW0UI6tWfgf1PT+8qZ+pdRS5X6de87xnmN14WLMIUpV+UKNsxgUAlZ+evmOiVXoUtGar
xIaHYStnavtmqAIjriW9U9iH5bmit5bFzbXV4pD4NOy8nEggGNwdOWQvSy+Lsg7tI3QtkX0sAM6+
yNl0W4OTKV4soxuZ6yBfwhulK61hseSZILpn/2eIlS5HeM10vRdfiezYwnuq3E6BBya0XGB57ZOT
mivAnTS4b8LS32tTDDLuTbfQVSTv9Y8apFfYyxKcIioWsytsc1UKxgiOJRH0uhMD9nLeI2E6PDkz
Daz0Zo25RX95aTGiAy+yaFp0dgCHwnRjmjAGn6BDl8K3+gTw6BxwgcyCpGXK97XWGQKVJ4su376W
UpU+EqUa8WJKzxjgqnQAgZXB+6Yb3lZrJuKH8PpnY5RL/h77OkUlSyBXufQdQPFlktGvIJ/Ag+Nr
hLouCNkcEWx/hdfrWt1kW82Lxb7vTb0xVjflRWO+WbuPsA7K630DDUMUESwR9MXUUVNGWnwp/C51
hy7AIP1+p/h/h2lkXnN1WM7oXgdAveSoPlz/NdLSULxaOSmRte1y//avYAgKtmw5MuXTCZBk/ooR
a6uT2fKX6sul3Al4Mwlr0IDJs3MSaMhQkVQjxrVkz8tUngJUNtNeFweJQbJ8Zn+RzLPngQwGH8YW
0M8HoH3FaiD5SEuGdPwtWETIdzRJTLh0SfuepCw4rGQFczr0EKg4OzSm3cguBjA+5X12Cg2IWQ1q
ZtVaLyLPjNx7saxKK9KZNauWNcP5uZLP4AMd9vuFJzSKJZZ+qld1oTvqZgn7puggW5j+HuMY4nkW
qLLw14jpn1w5EOWmU7fiyA2ARW6X0G3oGMYDR/5G+2tcFDodEMkc5uXtDeD16BvlM/E6kJDwORPQ
UYs208Zezmlm7l4EiRywWbvVPhS7grP1tLF9exahYJWxGwTdRviWdSCMve283rfWgHWyydOZXvTM
pK4jh5+P5fIicM5QBzRYkzjmxDuEC2yk6UjpkkxWO8RnnSfAy1E0GZ1ieMvI2xQ6BoAcITINyjVx
12g+dk/Inr+3oSLMCA4LflDCERKarWuqpXAoZoacFwi0pnAAAdYewYdilHYI9k10uNRsFh3rNGhP
bZJ3Tg68i/LBUIP7IpYH/2jf1fDQW8aQ/TGrHjaf/bfGb5PVP5S2UlGV2NClSVtZmjAXVSE5b8sp
iIgEWqoHNBhj1PmL56chcIBPffknscjECvua1H/7bgvohszNmGRcJbzqM8w6SM3qoAPbx+LtPAoo
+vzBhBZUPo/ZWgZnPhawYUYUzahTvlrxa3bKiVqU+a/i3HAXvC6YJapjAHADnYcv4J2DXFkE0NWb
e/UUwIRrnlfwxAidQOkaIN7JHRDhNRcse+cT924sAn9eNhdEKrb1CG5CD0pty8pWCrDpvMJAOFC2
JKXahnZiRpZiW5h/+5V9TYDZdkDQX9T1yummVxFefqWkpuFBnxDu9VCxMzCuLAFu6D2s4GRbZvRJ
5sjL991mXYSnhFHxbEQYU/A4jegHl2zgbcNsUfGtnWr9HcHHF96pydpWWiEwmjZjdykE1B80xe8R
LHg4zsylZ5l0q9y675FdvNTVYLabRnOBfEXcpIoG+DuahfQMPgLn1ox8gEAhrmSk+/kUWBUvOIm3
3/b3p/S2eAOWmX4eYkTeTiBgaJYGZ/beEmgK0SzQR2x1wlhMfnJZArY+2yXzI6A7aFo9j1CAeb38
bMOhqI07Gd9lNfPdoDizhiD77sFBDB+i6PzOrCIc2Umey8vudo4LGepaPw0dqoJ3wdKswCwHprwV
AbXjUpsbl7Vp4yKRnt8ePnp7SfKKirVHundeY4swDUVQE6IzYO9DI5ITOlXVPd3oBgLMceiEsBu2
x76ZGRKueofKj50ND+b6gpuj5fny8ygeBIGG/nNCuM9dbl0+RkQ8DociEKBhXXOqpniNBltmTBTZ
+bP0k8HkxFZ69swzjNxfxvBq18T9CHu9lKzSdbE1HAiUEsMSLcp6+IooQ2DsTCFuVvL6EDiQN+pw
p0/jyWEe8TxVHqJzcfkJHPwD+OGBLmI8wuV5pNt42XWWS8crhYnJ+cr6nB57JPgjpvwi4mfhw5CT
rit99ygNLTh848CQz0w/ZNqI4MSKjQmO7xvtD34wLj2KP6FhoWD8f0G9ovr5310NJJQDL1HK2eNH
j9+2Naa4usgn+VQbkEC4MsjeYa15l3X0CWBVa6U2hRx4ZwNeGVE2/R9/EgpwTrLIrY522E20u3Xv
vkwcln0p72GRNLeJMU+ZDsXJFk5F22UEmT0q5l1uhblXLaXM+E8N6RppVtYod5Tp7WlYNKBwnES8
Dhmk25L/3l6jWFir9hGuxV+ACwYA1TSiEA1HuWUNb+sCN4d0jSvpo5+V8da0a4jQc9VXKPnFFcFG
9q4ZjDNSmCgiBiEj71tBhu+bn3/4R4jW5mTbgAwRpaTHvzwp8tVc28ECYZxj26P5Mj++pqMVEjP8
b6FSRPM1TiHJOormlUUKK2/54YIG76d9U/pYlGMeyu2ZQK4nyM4ekjEsaTZUGe/zx+96iojwwtka
lyXfmxokDUlvxRh8A2yMTEUPYSY00qxbWT8AwloxlTkQviK58ypEztPOWAIL6R+/eAke1B1hZrFx
nqGcGqTW1dLUA1ojEfUZVAcPPep9qjtG5Id9jEZfAos33XEHOgz7qVPLAoXwQXv4D91djXxg1au7
9kG1R2XM0BFYEbjcn/lgD7vC1ADE19FQh2PUX2waeAt5LI+KtoZmCOx0Vxnk47IGUDl3d0XcXLuo
C1RycyVZN2b+8XD/GYrOmUBdZaOM82/xIEdCDO0d2RMTfBs4NjwnBB2G6WZBLzbFvOkvAReGid5O
KB0MVu4uc7hKp2VHtYSjiXOdMcw4GvtW/CtwS7M2XiLAPYO1F9anz1fr5FFC3RiFLsxNI3ZxLTtx
jPTrXDi31VFtxw2FWn3//8OtLkn1FOssbzxNmtSHmBHfzsTBUH5BkajeIklLqHVWPUoI689iBn6T
WqnUsuVAvz8Ys3WfoM/kyyf7R2R6N5EkiWv8uJnc68lo34SimIK4sy2rs8Z8YX5QEasEfkTxzuSc
Gmh18AUtviKys6W2MOvsLup1FmZ4A2imhbfeRfQBT1c3dZAyA+LMehT4wkSEMtuz0LnHuOehg///
SCDHNmJhDsmX6Xb2AF0KVXrcmEw7KuH05rn+IdFCQVFBzymNt2fQ3C9goe9YE9XM8JP4XuOT7SU9
DyzpllmXHp36Ryf1ACV1QtpgxHq8o2TT6c8T17OCdk0/LQwejQ9biiZ8P3AdtR5ty2PKINmNOqqE
hvN9mue3v5Y7kpUatHuSkYVAhyPCmO+ZXWt7nGoBbtkcAZoeH/iSM8Sh3uEpgkYuhYzOltnfOtkh
xxjWw1HE6R6y9Z0hkM31a44ZnNzVX6Jbt7wRMPmjVytFx87tQ2NAd8LExFdu9xKEyrRtHlUCmXgk
wL+E5YI71NBmmCgeVIdikCY3FXmyHEXYAxCWfDphTyAFflI8rfa2kqR4bBEwxLSySGjJ/2d8Aawv
XGHxm7RD9etz3BunXzX7DiuKIWV38hdbzhnZG5O76SuNahsDCmKecpntvCPytMNgihWVrUI0z/z3
C//pRy4g/1jyAWvg0TsIAex0LdjckVHYrBm1WV20zuAdU4+6JPz6aV9O0bavsSc+lESQCK8Y9ZfG
9K0E8A2lcAagy+SG5V7AXiEh3B5fKyzEf2d3d13QtD+8McKWIwb1Ob/8vfXC+lo0lj9HH8T0n5hD
ukuf/z8HKz3V4XxbP7pwwJjcKUY0FZhSUq8z7VauUnGbcOi0yFaDIIDD+Dwa09MJnVDWydUw5jJB
nxrtSj7X4bKPK9QdNxqxkWCASHZBhn172GV7g0X528oI4AkccEYGj3yQruO+m4z2nGDtGqN46I9Q
RdlpooLPPrsJxdxIo/BQsZbZ8bMOCSZF8dgZwOYo2rf9BJySWpoEF6b+n2CggrMaGfWyLnEyoQ7S
qyozDExKe1f3b4H+gYK2B+PamM7rSWcG9b2zQ9SG6Bf0Nnnfsu2Glup+aUE3DPcglzkVmSSho3gM
1V1ejClOmNFOtS2rSfO3aXKmcRd76kJMDKWbNi6eSVbO+llAScx9wF8jn0rfS4F25V34G5HCa2yI
sfNmWjEyysifGaCisvKm6//4YSt8DB1shpr4nFS6WbgWCDrm3XY94s/XfcJEB548Zorfg+2VjgW/
I3s8E33AVofZ+JDUQ3jdEbdmNrMDOmARcfK7b+qx5QRMi5/QFbhie1blFvf33n0tNnJL19bfHIm0
fxIRgX8gM4YfjICUiEM5xQIaB17V+22i2gMfLSMPl3rSzi+107nfrT6yhqoV3t50gOu9BHXNt2WK
ymJaktpCBlssytIr1Hw0l+qTLISb30J+A1Y0WE+PHOke/05UekUUk4odMof7jrvq3f8kx+IBkPG/
T9v8xF9M6BgqRBKqs25MNdjhxVstuNLEXSPAOOfGi2P91Kp+ecRqbuKSUa7TeBuJRXjiowIPsWq6
LjJNqPFRAs6O25xZpOk2CZfEgBHUc0jz5kKEmwWeBMIuAKnAZUyDiCtqYH+87Qc+NPHWuGDGsSX+
MPt1dEv4NvfwImqjvzrF51YYPN2dXrg5op9Cd633lBblGsPNkoz+eUsQOb7SpVUoy57OMQt4GNJf
AfErBALsZlifkuhyu8tBt98MkMo4b1gZ+NvsP4b/xjl9ncOCuKSnubxsKSQX55JLkiierImDCENs
pSXBQOpC/XuPf2f/GQ34RQ/whVJ1O2Fvmp5LTaD3tH/ggnsDSraRzqUo0AKr6+qOCPDSl3U0ii4/
NdObDEfF6R1r3T7+iwdp37fp/R54AdMCO8IrQ11kC4kp6Kj/fMEMtl94vKYXkHWUThQptc/9cBge
7d8vDvScvLSWh/Pgocr2tqIwGgFKlUr5eb5MVCTIa2wSu+b18235BQQqMLGlg59pzQGzqsYq9nnv
G3PHcEN7astCn+bWiZwwj6vVPxlBVlmQiFZ5fBlE7UPmXTuDgc26YdbaHu92PLP7Pkqvdm2Cd1wv
jzzi1vXgubrWsBPdPtzK4bhNl6fLPPSfBPCEBAniJME1TfHLlYpwFHwSMDCs3r5/UQXHG6FPc9re
Fu0pvgu28MxI1LXetdO+pC3kVRzC2qg07PNbHUW7VGWo/eekFDjV2M2qjPYVHx5RNw9tWEfFtg0k
2xeMtsvDaswARmaa0yx+w0L9SfNUZADmtVYJVXyFgDs0s4O4OVoFQmUZBf8m26N6m4cUOVb1fAUd
NwNQUi/OALw3qKZaOvZ8sptZHakYN4zhJ/ftPIXdj04g/zIHXzNbgYE+S2qRgS+44M2Dp96YKiy2
3clCawAZF0tz4rs3PkaTyee+/Zvf/GO/M2Ym2WEfZKL/mSIZsqDPLCVip8jh47iP1jKfMvcoPv/Y
FZAXaUcTwegUOuP2R2obzXJ8SuB6YOyMs6sjjIGv0FWaAffGEs7pLBIVQQ1DCiqoI8kHkk/XitB3
6enLdKlrvBSgsrZvsEH0GcnsijjEDaYrgiHB9jseRo7g2sDYTOVyiuJz9yjPzhG2FllhY1i/FRpj
jZPSTH0BG4A6TMyKvdvfAvYDduio1vmTstEocYWCVDv5D7VLINn8ba/orCS31+mGVCidYKUJXGsl
eVLCmz16HIDW9BMoivgiVV+6vqx84DlfMBKfgNyTUJonxLsBD7Wfabc5hgRtBl8VTO+q1x0IONWG
Ob70ScL0McERdCjItyLppJYGIoiBbq5Uh4eJrU1KWjJsn0P++2wPMPXzjorRVh6VdEiNJX+OsK31
n4E3gYj2en48SH48ZfPsX1j7Vv+h0oubZ4zlfmPSPI6XN8isYHEbT7FPi7z8HTLejyTrybrho7St
sk9BS51zRu94mAK7VnDIFEaNOkfbUJ0VieupINF7m0QO3oEwZzbbs+tDBi8J4xz08CRXS60nC3rN
Pen9s+zGFYlAZ9f5vWj7CgCjlvNK53oHb89h9NXVMuBVKRre+BJt1JfNxXKR5jXJ5GXNU19RLnN9
qXZp1KNyMSARKXXEOLQz4NE1Exwjz5OftTMyK9wpfI6YS/WZpjlSY6IN6qtK5kVC5tOCZ106sBnV
YPm3EOd0FuySYD7RSvVIkFNkvgM0dbzdkceZXuOEE8cL5mqpYyEgKjAuKBiuZeFmCx19i4F6G1qw
4Q6AQW84HH00hNR4nuhbfOoxOKFC2x6Sid7sEPhVNmNP6OQXSw3kb2GU4VvJAJJbq9PC9EXHkph+
i3k2ahIFlfyec+3a+xyJKosLTw2767jJPs4rVPgXa7PMLXhPbJjNH+79F0ju+Otdh4Bl0/BrszG6
W3iw73aex2frH7iBSYbV0XG+1iO85HiaM/uCZFhsRPtP1m6fwGRF6qGR4UsVPXOFRfyG0vdl1qlQ
9pENl7a9YqCaucnBmOLvowoDyvpsc4e4GjzBE5wYgrL2KnMPlc9EqLFf9JoHHlVr36QpSAYM6wVs
pOcIDiB/9Q4lwBAVOGqVprFHIxT1IsV6PPNTzvy3w1UQG5/TsisusVMuqL4HGU7SDg0+e5gZwugP
8OAFaKI3TxqjSKAtScxKBKjs4fmb4/vFMnaaOb9I3wyZqAY2GmODHw/2P0VXmfAFVfLV8nOQaGbj
Tmm5e84dC0B2e6JaOeTnFNasIbufTTZAUAkzjLst6A9jLHcTVhkfFkk4cCtt2fOTDsKBo/MKIXXG
tO+213fH1sX+0CDY2mZTIdGkGzFjxI6WG1NTsQoPI7gfqpBlYfLZkkoJW9753uJwRBwGFkCMzLat
S1tmSiSGtDu7mw3lRkPx8FusqIakLz7g7w7eUXbqrW4gRLT/kYYCk2vIJwgpHpxIO+0UuFeWXJ3M
GDtTLMzuPvtWpDsykldh9e/Oc2bWdAxr128GNTOqU3qQ4UVDg2VrCn8TlMxIlGihLzdhNEBv3O2T
di1q75ldE+4BcBbyS4E/hL9MJXBA3FRnKjqT1uwSyrkRP1cQ4kPUvZ8V8RLtlRT8JuUNfJULrCgd
Vam+B03wz8D6J0Uw9afK7bNYAPuCf3ZEkZukhzrb9jWCIoRp1hNqxNqOt5W5R3PzYj0UTQ60Rgiz
K5yd4G2Cb6/Aoeb7XtzMzZOVCaNItQaQkxIixJS+iVT4sWvo2+1CzERw44FMhHPxkqtX+YYiIzRT
Nz2zDk+Jm4PIjPAVLiBg5+LC0obe4CVdgu4J0jnx2F5gjoKCnw8AMv9ZfCsQD81xMazmvh1cUQ2R
sv2KujBB9VWQAvMMpR3DCGd0p7R31jJgWVZft+EGWTd9kT4dAkA3aag6wI6sCmmejIMVnEeDiInY
gLxF/1JFnVgrMMU7ZN33APsWSJCbCJ2I8AU2zZDlDV+9acusqw8ELrZOkgu0hEh6WjD+RJFXY+7S
NCP0KkMCIa4SlWahiTx5aw72me2k/2rA9tfYM1DDFMYF9vh0+xnxYANV91nUIsRarUjb2sJOhrFt
ZdHUXcjwZfM76+J8e0IIZbhfVywxyx9/2PUp4hDD/PVyNajBKYN/QAAzoFES0dOlcu+wHcIKMu8/
vbpoblhW/r+zmRh6Y2F8dbPJO//Ir6OLKw/Fnq6G0jyLgmOclLwuF9yLyorPCkX/qQHAiBGaOly4
qMVl8ViomucxZoCoUJNRePPyZCmRHczsn2dw351UN2U0EgacGF3wD8DlaDEt4xRWrYeQgANaqcQA
sNop8pFx028tJaff5AsOCQ/guTYubA8ASYnmowrjlAxLqMMcHnMum71VOswu8/IEz8rGq5m5n772
Wu/MtfKRV2/F5IO30NyQoLR6p6EkJXMGDKo3MUs1uhurpdpFXxM6kq9qEgRmNDyx8DVkUNlZF2W+
SYAbJo6Rj872NWGkV2wNQWtioeYGSLJHL75pu2uPpHBO0cpYHIabow/TwnLX40AjymvgIbg4HeIP
md3wSEMwTJH6W52T2acPQQFW/7IsGaxrWVg+SlEckq/JllB3lbeySHcD+pJy/M9+GzLVaNCz8+Tl
4UN8DFu1RKhIa/WhNZfAH9iDDCPywADDlr0U1HN09RNVqL9D7eH4stcxVMqUlrC7NjoRy2ztQXey
wTIRrYvYTaiHAJ+jzwVtRJxq0316Fwj1TIx+6NxWps99aZuxKR1/f/bpQcOdilNjMnOhch5TYxtb
moCwPdic5tybW8G00QOktHVHlqAE9E0umzg3iy0WU0fx3EObYv55NsfnCF45zovhDtVR30JoRLJ2
mEMVONdbhyeJt1A/XDtYsFhxYeK/yD/Dfhw9fj8Hx7hVAJRCEdqW1Ofa2CGXByXIScdbqgJgMgZ3
KWzUSHgVVnIo82SNGzGbUuB+QyYBE2HRoy64+EXkHbRkGEO9UZSiyppgya0jyRoaghtnGkas67oH
FUG37gOsEEcNjpwLnquMtSlGA6/vG/dlOcomDtR0b/ePNuwBweJ08kjAqBf8yJolJ79ZHeeX7IPj
WhwfUctidrLQ664xr9LDu8T8noXBJAftLD/NJbR/R+al8cuivCQizQ5Y93x3lmSsuM7dC+IxkFF1
jvxlDhVl4LzLOAfheiWj4tZ/Klb+zYKVIP/PxJtsWqe4K7xPVmCLDXXKGrnm3FeZrTALOe8zRaWW
3t5MLFa2hNBYRWj1iekklaw2Y9nBec8X0W2HmLkCsorXwzEpyvVqOm7OxJlOt3cCn4iAGCS2IfwJ
+ETFBqELNjwdRMy9+FCDAQVLWNhz7sTMFN/eLcVYxiwAhXlVMNRfA3gWdVciKYJTUdFt57BvCor2
e2ZO/0Ue7WHbNkvq7ar+C5PJux+PfpzvFyIxx+xsYbIlVx9h027L0577EQltgZD3YafbLogYIGC8
fXrh+n1V8EVEQaLHw0gc6ZyUc2BXes09xStId9L1Gu6PVaEEsARIqUGiRIMCzHS3aPQoqMwDKNfH
W8Ve6cFbsH5hzMTrmm45oMJsT9ReqbOPZ4VJwx16f5pPwcqGDo4NZmjmMpGLB2TfCsZZzl83UGDZ
3hpjj0bKHBheVmZCZfTxD0zf6mtZKhY9HOdJfQM1SvU7hjLgOAvPG9JIRcv6xS9uSDTHhEZhBKcJ
7lcQiZ+gjmz4Pk4HMRoHibCG759PoQIJurgARDhA87BQ7i0FX13ClXXZll2nUHCcaMtdnUjWm6ir
PcsCZUMhcs0Ebd+QSG/7/O8RZxFqKZMtsS2bTH7wlbSeSvH0YnXM2EnMtKKAgWOVBO9ZYsQmi5qH
dLLeYybbsVdS6+9tsnEA/CATQpvpORIkaN8ifeyVT64SOqI8t8srYhLl5OCrFdCv6tBOAwoqw9Kd
Y+vz8cjJhJtpWtBCVgUm5gqr0GOQANFkviSJfXOHzeIf7zL606+nY18qN2e/XWbGlY4uSk7aGuh3
0PB06d+vTcVFsSMZ/K78sShuOrpa+0VbIzbQuQEUAiJ+f9+Ie1ZixAeB0h5gdCkjT3gQUpIav3vd
57AkytzD19ai3HlkrT+fZkiuQKMpOBdB52jIxVZFufws2FjNaklPzu4HSU6eKR1WxJ2qyJGhROgG
oOSWljDzLgqXjr7eRShwLhtFfWn20k7U/AfQE9q/l3DmjYnmUZt3V6Qy6QvyXB53diz1g/QtZtny
z9zW/qPP/d59yLUxSqyqbk9XfdfpUmlaMRimrA0/NLke+WvsaYn039EhX3BDVMblWmOEyF7sV5JS
jd17M1DnrVVYusNPtRf8NzpvomtI8UPB+SwidyuhEWKSL/roeVKCjc3qUEJK4p+iN2u8jVORnI2h
zxvDhLrG9WZHHu2zkZJ3WaylaJ5dCPakrcFFG1VsTtoTBFHvguGnxMJOGhccJkx4tmvLJnNEakJi
UwMiBoYqUfx0bRyhfbXqEkudscdOfb2aQCjkGt6bAu4vAFuoHZ5++E0poDcPiDTNtGHoe31ENF5Q
IQeE82WLxvijfCUyEgFs2qCIg2CdCDW8420ihMHevZ5SLqcBsomFA+HZsACOdyzCIjTLynhtH3Fy
czmUkTgs029U4uUanbQDvDZfTC33KCnZtBZlGmXi+RNdtBZjt02dHAyzzGNzmDlIsPfAnbZZSyKL
kihBf+SgRT+pKAYPfjvWGmK+7anqXNjbGvBWlM6g7TxhgyztT8WGrVBkaQKo0FNGzu3RgM3qzZyg
5Zi2UuoGfmTo3f2j9noW/AhTHokbPPG9H23j+H4235n6PgIPMFw+zG6esfEU96k0QLWVyhl63q6P
Av7AA9kQ2zQ2jD83s8RERCj0t3DQefrCxUitxiaQwkDd1zl1djnc8eJQJi9U+oeoqqfgUPFzp5c+
bs6t1mjd0U0Qh/j0Uc4GK2D/xfuRw4PYPDmciuFH4aTo6/Ix8bAcKv5t5LsDAPitZ7GaW6as5iVx
N/vJfPIFdZ4PPqTOQYSHs6CytMQ6zjSE1XpjRGbrAsiFt7nOYHGfRrvw3cJEGsOL1srkHFm0HlSo
ar2vQGDHMB7/2+IOSNGQeTC2AKlhueVkBG+ZwE38h53xMW8ltHWCPTmuD6duwSVRGTrYTRrbgiWG
suHWewEBGS0GXzg3b2YtsUFSx98aQ4fLwprLs/4h5JFvtN0pHw2aMXM5bwr8Dp12YHx9eZXNT/Cq
HBkKV7hUamE+bOFwMhrJ22gBoIXIwTN0ZACW1eQM/IekbfjzyqrfzVLBuP5YiLCuh4Rm0W/C9Jp1
6thX4PaYxw9JO+Qb+jpjN3MK+ZI/+/sP7OfgK4xpcQj2sfrGOU8zITpN0z8Om4N+2cfIuYhwfrOx
RwW5GTDFLq+UPJbsfnQB91ULMU/+PzstcvryT9fRtxTt363x5ddsZn5BAA81A+3MIF/YcpTxFROC
VRlgWLCMd/UIq+bo5vcBBGzaKzGXuc4xuonuc1vP1Mo21br1gFzzTaivSZ/QkJ61bQEFePjWgNEa
27g8rkYV0vBfEDVO5V4VHWvPTXhw0On7MvebRNpibCXTE11StJ34tDbrgjmHsJu47jHoiOwEboFL
a/H4cDEOt26UbFfnRsKjkNBrEBkD9twk3p5xrua2oQ6Yyo0uMJcPqYoOwmW8Tueaz6NOf7HJ8fG9
d0xaRVwH9/wDNzusJg1sCQ+hnrCNITghx6gOrzkqPjUw0Rz4dTljLFg6Bvw0IjuXyJmwrWogUJd7
V9+mIoFfzYTAYypRHS+F0EDaE27SYeEFApLVONlfywmgGF5d8cDnxrGSter4urxq4mk6UtxhnyGY
odXr6Y+GEY9jzVLOHkKRavRBMkuJlyea+rAtS5rFeiQhcMWvsNfkei9kXDggVNWlzqyNXfgjIbtR
hNUt82LcLnmtwJfO9rRBbTJ0eVJE+eK/rAocqoO6Xys0Q1dEShZ8UyMmMOYy0x50M1IfCLal/vQ1
QF8JrOJVXFFvM0gKvWOMBoD3aVqThKEbIOkxTidra2V5g13AfXsx1ys4+Lx+vkKWENRlDInMNv+L
CKqkRSp4wFKs2Go6OYG3rMmkuecHgu8cM7ypTHNmbvNJQqUUzvsyx/l1gyabgMAvaKlmlH/P03Us
HSLT5uUpp7UKSrPBcoOk+pdYd0ZBELkzSe8mysBi4WXSGfzAngbGBxn7aFE7kSRnLPBOyYhpoDDN
L9dHH05xP3T01WAJRK7zGnO4GVM6jDZpWhj+SGvYdpFj8qyzoKOjPN0DSClIvUu8DJAynTR8UnMg
2KArwiCpKkTc4Xkvvh5VYz687VJDRnmYQPvn0G0ijKetvFhIIWJ0usYQlwCZ0YoWPVOyA07u1W0i
8HPJ9x3Xby6XT1DeQdAdbjb1CIMNRnDnTYTlAAfvwIRruZMHEN65VXnMZLRG+S+/XMRCTdpwFq35
nVKKzAsL/IleAQNrnmE6zwNlx8oZZeRmTTR/LdpqFZ62AafW1nAtWiAacku8qcRF11SaPh92PUfo
mkAoxwzIMYMg6Z0lj135XVqGtd8Tq2kJ13KZAxmjj3Y5F3FhB5mK2eOkFsGcFw/rQe/b08rp7HjM
A13wGriI1rnw3ykuIxPzcJBitOsrmlL653gDKcs420XEqWaHV2si/YvXBPZgFUgGQbV8IhKUkQo+
iLI+AOzvjCLMLdpVN0HzCvwRiaWS+s1v5bQ8g+HF94UQqGdnAZwrWGg3TwFISvWhekGn5R8K5w3a
kudogUYSJE5SpcZNSJ5wsyQEU/CYjKgJD2ujgenffAAeBkoHYDS4dGfrhND5lrTQUOYioQRdgsoi
//1/0Vt6wjB+PTKT4rt23CUX2vk67JH8D+FT4cTQrbvm2lyq5QCsAui5+9hYxfDKXtn+HpEqUxap
FSPrf0Lq3hQ14FI1R6NcjhcxWz3MSzzD644DYLcQ/tpIne/tQIvW9fJC0xpk79oNtljtNotbk3iR
1YGKz1YBmlk5yroDYbK0+bPvUWptC8CHRumU5REMPNAKRQFrdnQ1gp6PqWJMWr3pGoXbwEBb3dw5
P9IeCjvA1tOsx0D86gov9OVxxETfO3z165HsISg/ikEzgnhmjlUsIuFED7J3svMzwKSLu5bF7qTb
c0ZfkKlWrYeDVa/0N8F4iQqFpWxcFfDZTF/lHsFZGRcaWfB2SoE8ZycRqOTF0sXvAFQ20H2Avs3O
UhrbZiEzjcefQponG9V7nHbOfkzV6AygFjrZN22SLYUWdZ2I4BkdadyKksxZgZSmQkNCuLBdrLs8
HH17LjgSUyUAVuMtZkzyV+PWzxAqTrF1xVVzfTiX+TA/md4PbjDjb9YtKXYxAa2h18lH6KtmH0Pg
f9U0hWDjTIZ4Rxl3jdE6jmEfZZleYDWjM3vexbDxiprncF/2Ewep4ZGNQyIIsgJWt61ZPBgo/KXG
T5HazIFXH9hjNewVzJlQ19YE+kUwvWbo5qKaqZfWlyA/kSPP/D7PVa05Tgoon7E6KjMSaYHH5PNz
T99qXZP0FY9WQFgN9tWMhT+I7yPalVeantUntpT4UNdf5LjG2uMccqx9lk+1FVJmv0cKEaFC72aH
aHsuK5QJhCY/8xEapW+ya+FFDjQOYwFQ1/DrYvhNgkDDZWPZWvPRsyFCTTVuVkHKpuH5jEd71a8P
sXBNeiyboQnlaNCe/WwxI4WrWTl7tNzyqD2ZUenSBwjxioASkSrp8iplj3Jr+CPpfb00TyasJkYS
53bjMnBGYWNMwCATan0OMxq2I/dai9TnXU4oFWG4A32A/D+AFHvfsyTaR6Kl+IsLAJLVIEb4jhMj
SBybD0seI89GNbOqlhKz6nLCUkXS6u88MuRk9G8QIdJvBT/wrpNr0IoQD3AeJQ6UZQNsQTvUEJRK
Whv4fYITxfIZGiztY85z+oC4LFhCkhGTRtM2OFGr3vJh7qf5zt/jUoomlugXp2nR+3Skv2vufbid
eOL7vl2uAd09eZPIqzKlS2hDqb5r6Urg+o+zekfmMpAb98du2JOuwuBtlndpOL03YMRO9HqIOtHf
4xhbk+GkpWDntmXaMCo3hQQe+K3KYfnYwfRvryuDjAkOi6f3I9qnIdY4nRJDgH3MpmgC2PKJGY6j
75txzPEuTXkj8QQtMWBR9WHmVKWz32Xus83LzcvWuxh8y26aBxlbNltBrohZ1e3QDUUZojZ3ApZ6
H8D7q4NlnUc5/54UzWl4+GO/hYgACscX/jUdx+2IetVeerS5Gfty/Az+EaA/cUwalNK2V1Kx1M9K
R1Cdjg1mFeb7VpnGtM6b3PGXcpSQzbQF/LAjdfU/tdXXxrl0KJsIrbsht+RjMLsUv93h72Oq0cBB
CmoOQ7mpBcwHYKctEo2+U/xlzb3HVgQr9Up9pCpLxjz6pT/gvmKh2DSaylgLE0/rqqvm6PZGq8go
rOunMlchPNJZN41HML2UIKWFYPFKx4jlG/AvvwgcjoiikdBph5xvWfra7MwWVMxfyTDHxT9myggg
2DI9m/gYkBzgTi7hkRtvKvKY/YV/kfZRgX7yOURMG64KjuBgiqQaoVycwUbneQaoRCYvAeNK3K19
FrwX/T8INCun689GieazR2/wrNoFp6BkOwPI2Wj94VOzzwlYS9kF4ii5MU/mAezZqiMnRZ4x041L
HJW8depeD5QE3BTbw0wxu/ve/sTCtKUmtJhl6ooxTPQpvcg4qr7GqfP6vZbIO4+UZ8lOhPYP9CCO
FM26bzDMaOa+jhx8K8owET0lZD6o5FWrJvmgx91MrYtyxAdsuKCBgcD7DEQ028qrH5fBOU3pP0f/
fRZgfCRnlfj+y3XWo0hDG7+4cpkzg1Wq/ePcLWeneWXzrYCtKhk5qGSr1mu6UnfG0mWSL4dL7sKt
X2UK7a78ddxLWN0xaDY8BL737mhtsxe2uYxyHaJmPDEUd0iUyS2rjBfIuPhr/B+b6b/0oUqfjHd7
O6bvWNtjQNZE9mYU1K6bCWn912cBlsVwSKPwt9mkUlrcRWTt2mIvLq+8D7E9ii0+cAYaJVtuOODk
Og2C8z/C1FWfJ267hsDmJo3rqEd4FN/lL66n0THgf55AnLLfSy1tGRwmNecdWGR03/vDtqXwDFuQ
Adwew4uZTdrF3eir8gs10O80xXbG8LjotD04xMwX/QpE9D0Tb5cC/UJc0t1LmihPZziTBVySE8Fh
ysb9shF4/278Iq0vBzzalQ0XhW7GvJjrpxNrCF7wwnh3TWy/o3XeZFvfS7WfKJ0o7XmT2lWSKk9x
gOqyJa8s7Ge/uXW3zZn0ssqVfuxFGjppfWyLBroR+dvnYsNFDpIoRsiKe8qgpCL1WNjrfZ9CldET
Hd63drPvca9h6jzc4mFuBcYQ4qO1vJHzPzK3EU40kqAaUCGlPSpozWWp/x+CKb+FvcMMkW/It5ij
DheaPTj0svBQqLWmNjFwK7rROKvSMTv4xwfcWzfW0eTVoJP/d0envzl06OtCqrVAJp6W9QPvEyPT
KuVLOu0ShVoffoM54DqUWmqf72vDCMMYOcicAHbbSs4FKFVcZVvC0g1QWEPGQ8K52+VEx4RXh3np
YZS4MZY9Db2jtJ5wmqkKOpOD+kG5/Q+oS1hrZGm2mAbHSr8CTlQOYRu6WDimYYVbxnQ+9oqjFdP7
hIi9TWm8q98XVxhzLBqJYnsIA28nndKEqWS6oxZyd7kU+Rbl/G0pxC03JrxANIPI60DxgV9fWXEk
iGaSg915RZRGKG0aiAAgO0Xl5q4DyYJBQexw6ma1piMq3wtMcMnmsQbV83al5gxDPvimATNsmjyw
kBX0MpP//bNGI0D48X3VjtSpHAuSc60IV4fnGP9cxVJaNqrztnKoRTu0FScjkEiIJ9FSxQjn2VsL
NuEDar3Gud7kLHEtC+R1s8FrElXO1lW0sHO2+hLy504ai3RX9x1956ceBWJOX/QvHK1in9+GkX20
l1WUWDPhJb3Bxx+IERNIhtFPXYuLvTWPKrVyCx7GOnbXXjBjkijXrSl9nc+wI9uibAXE1aCMa8Jb
Ooz3A+yXnwVAhyC0kPmiDHk1kEJrSghq3Eq3Qnm+IedgtYBcSDz5MDD8qEhWP898qN5LwYnX4OSs
L00KL8dk8qolIVAZlwJfNONz2jwYZBz1K4x6EXBlI4eDgipXYlV0Dh5CXIIZ8hLjPItMLlKTQzZA
qUpA8bsm+TYX0btEcY5F5Du/8jqQj1VvvfuHCmrkCBAZrW8ZR00oBfO4peF2U0rBCzMGc6wvXSb8
t6f7K7616xvFkdbChz4UWieA5/LKjtOVuhWjDBXmyZgS3S14AcqYK2OBTegGOeuTXzFF96wF8L2f
HpDPd5/RbXOprMq98aR9k/4rZdL9Xw+n0Tf5mS1aY4/HrG28xlU0ipK3Q2Wy1WyqQg5ATys3X/Ek
gcCd+d3ZnnednqgM3heY5RCrFJh5IRYLH8N8QVTopwK7TOXBqRJC/l7+RJ/P/5TPo54HDQsw6TDX
ZF/mIE15y+9tP81Nly006DYyC4+NjAPzJS9IsGLLK+cJG/ME15ygnJVJ8+P/o/WV1J/ia4FFfdGe
y22eoKD2CMgzthShBfBnU2yihm69CPao06JFLokNZNK5SxeVAR9mw8lLZRkAezgftVJCxSuX2V2o
QokucklRw0RldgxX7imcFiAhLIvbVXzKDoLnkRFwm6hF9n+49ABeFyW6TMk7btDDtiRf0qGKVR2h
gPkW5DZThNMo8RFBhnb98+hRkepSjsqcnRpz5BEnfUW+mpuL698Txg7W2UJCAgyIbX9R5PoMQuFb
dsBw6JFyjuOJ4R1fCHPh7pLpPuIPwGAA9ATXj9c+FFF9DDYsfOE0gYCJOKOk/g3Ts4mYhVC0PsfB
Acy/Vt+SAoEL//PiyMn0houbolYQBuUd2AKK+xZDg2rCl+wsDnZisr8NRoFkOG18DSdBL7sBeVTm
jnISc7ePhU4Y05bDYxDoIyq3SaXQKPNblRCT9SPQTs+qO3RNUBwpXL0hvzP/Pkoxwx7HKzEXgQ6H
v7HjN4WrmtYB+i9aiv253hQtAuJHO8SJPT540PVKeNDc+Lc2gE32yvC4UQlza09E7uartJHkklMA
xwhCuIyaslJrvkjQeFK/z4RProUwO8LhEPBv8dS9XyKhYn+hHSBOqjHTDvzpcQ4JE3CyY7x1HsKW
HBLU6MzpDUEDQZHX3tyBfMW8aYq8L4UAE7FXeJuSSK3LHoXJGzp/kfTn8NSyWMGvXvgwF0gxrBnu
bYOa5FpAJpP+WsYKXyzeGbeu15ZRq140VrOse+xBanvYKV4Fj4T+BDKjbiiS8DnCBXwY8rZtdUTE
iT5AGy45G6jTQPXlPeDcCJwV+LzZrKjMEnws1O1Kke5FAP7FGfSCtSVC0cEbokU3+w8nmAX110LD
v4mMTdWvwaT7RqG2bloZw+EwproaU85MQJN66ivlvpv/ZZiy5/EEr1xsB5VIit1+2TfAna19sIJL
80YfS8r4lMgicLn5PDBPjYJ/tTMFByMklDOLxBOaMaQTE6e+Z4AnHTBU8XSXg9cdZDnaFQ6OCtNB
tTOcnmLRcHOLlNxYSg2yl5KUOxGwtK2vY5kkQe0BLslYvYGqyalO3vrzIiEx6e89oj1SlxKZSuT7
5YSnBMUmV+wvyjGH96diNgrLXc9d19GdnocXdVKRB6PIJWG8S4ICC6eWK5EPYZVCU9WDCJSfu5gP
SmF0+pvTs9WdSnj5Qe/G4GJDPB1k/cYDhoXPcHxv8er/TkoWcBBZ9POtnHbmm+zSoMHCcTF3qYzj
NQNq5a3Phnyc2Xq+LqCe+DONxV7qQxplqT/k7LYSqvQE6N8FWaKuV9nRu650g6bpuSEtrqCDRLi0
c3nqjW/XlTBRtiJFkMLrUnAYzJ5vS17zfUvy134lpnLr7xX9tWDIO7lWvWRToIjwa/Q++rJEBBE9
semMOCVUIM5e9t2cYnp09gFPbuX5Ki5NEN782wPokqyS5XlO+HtibJht+9HJoVhRrn7QwdFXtiNl
qWdhuPPhCTwrde6VxFBbSdfEfHmM0tH4mf9aXCb9rfMtjBLM+7CjE/iRufyJB1aQBP7VqD+1Adwr
NhEpOOELvF7NwLDcNQNsEjRNNmonf7MkipjYUYYa/FVZ+YDfLRGEfUxdQ91dGXge3GhmKQTX8mPu
8etPo+RspXHtjE4VkBhlaM8T3416UT7Lw3EdyoVdfGSjbKZ7BKj+ebT5oOyRoBVBpIHWluwGSb7t
0kHPoIgOaU4oE/PNNTYKYSKAjT7Yr1Xb0UIpgdPUUR2dOLsP8RiRdazEsXv8LhpBR0eX9JRrShkJ
IL3/LHobTarCN5GQKyXqqNnX169xLDMaU8lr9Vtfj4M/lCfovagEi54SBRr4lIn+KVx+HmXql+E0
J1lr/9QLxzuLfW0JssxQemGAT/py5/CTpTuG51+1DblDkmgXjK5py3FfDUevlrgieX3XL41rGFvX
M6KT9Qp14eUmWmook+QQMoJk0JWy5T1ldUNlghjZEQPWmYwffpNYX4q33gEV/kDDp1rmnYoEwuJG
2qIQ47dKAmeZPF31vWpAhGhJMjSHftYJVSxHMpfQ8OY7mwt4gEBx3+IITiRgvfXXcwSiKRRpbuiH
qldgKWxbwcPF3+EApWeBQttMmxXH2IRvtxJoF4SMYNpY1tSbkJYuRfIoo2jCtTnXejNuxs+U2uYt
JgFVw04sYrpjMeQ5UeNRbFERlhvPXtDnTRzTSewAH02HX9vjw8TMEOzqoptOPsz+5hqTK6G/M5Cx
oUkzSDIj04bTEMNycdeuw8hYs53SOg2xx1zIeoJDSqxVCQQzYF4GhAJqlbkfjB+OeJbZCjbk2FJe
nP+K7p2CugkBsFviCt+0O66gEA/AcTthbb0ZH1He3icWNLAD1IdNJPFHp1Q8zCgggNN4ZozoujYD
euP/K6is8cI2r2rW9chofF3vHBBzEnO9wMt/pwqRe0HqkgNsmLYS0xEQ4xJ8jd7ADU+rLW9X7oJs
i/bh0t++nK/wAUVym2J44z60DtXQEva6mh5AN/Ip63qDaiOhj1yN5CZQCpQ8Ixr1jPZ3sDaM8b5X
jtYTGf7t+RnNOVUazN+uRaixgWl7rmpHyFTIIMPQE08HeMzC0zBNk2ktoueSG781OtQqHf1C8/72
mDYWe0AjgG/k5/ppegHBEmHVPKlkIa9P8qd4mo1fMm9Fl2Eo/e0H1Jyxh+0yq+uxX4g2IK+ER1FP
kUivRkFcZkpqGrze6k6dbKq45px1R5gKV2JyJlU8NUdIUJLtI9yNbTnoV6GIPwvHnHy+IQVC+9ES
MOcz7L2UwZ8cUnlp9RTz2ByOAy0t43C2PuLT5AnWeFxdqG2i0+CsDLRXzO4iyoSaUIsY+gzbHdBb
0a2QrzL9G3u3DqbB5u5nmMRab8SVS9BrMmLBFN+Eg2BQprKp75qa6IMLcwv1gESOtDttqKtE33v4
Sq8xloWBFLFYk5JUaIKCqiruwkvwKO3tBx+2QuBp4h0bkQgqPlrHLi1qxCaj/YlGCFKZJnzo+ARl
Kh/iJhzkhqh4ZFiLYbQ1mYuW+jOGbmVGn5Ly3E4PQcy9X6nkzMx581y5H+JwJZNhO1VihKloahfU
l5eAHkpDB6azywpN9wfVpOo+WJb1P8gzwE6B+dDW0KCydpjHp/A5FTrL6E/e9Eb+IPz6qRKZ0FK2
T8HyWxpOUQTFzgFPIPb3lN/WA4zDQruBJq9qhh9CokeFfxIOzMwSJ7vsOrfRJTQra4HyuwSupsxv
ne9jZRHyubjRnR28pe5khYMJEQ8bQoJCCIpWou7PElZPTmNCM/S/W3RTcIRnupnKIetEIYwDYVEz
NYCHSSBgNbQxvK2YztUJ4bP3rfQUOg1kerw3ZMEFWlIswxK4CRYyAwLzNNXahM485O0TZLz//git
cyF0ab7YxDpIOMdmnU6o85/1tEKQtMcBxbsxDKLqfcXP47triCySZhsB7h27/yTlgEFhkbKa/iLJ
ZwHdSYyP9QmfA6r/XIjAQfJ6PJ3tKQW8BUiZCOLrGW3i5V1UMaMKOTuzxySWMn2N170vpK6u/gGb
93I7iHYVWCfL+LukuRKEq63YMv0CNtdSyXzhD/YXLGAziok98metQty0n5z+CIbE+vD/6Y/XEW1k
jp/7+lsAW0GIM8LvREns2bgxq9oKaChpJ7/dvalz8XhflsZv2Va2M8D7w7zLCg92129ey9qOidhH
M3/QV/mBUj7qBmqt1JTLvhK0qjImYKReVE1KolK3dFo2JbUf6Ko1hPDYI25A7QdkIm1YgzKczX6H
ISW61aXnB2PV9YuqxrcJD0+QsBkgX3XMzmGwZUQsfS4OtXPuUWqluSEeiFgcrtE84hp2KT8FAgDx
TIiD4zW0QCV79TBVdmiS8PlKQv134yyfr1kFHYN0HetF3TOa/+k8/VLPiEiPe5zrRJ7oN+Suk5Ju
pvlauq4orMCHaRK/2X2zypewe6gcjJhNjEfIPceceBSWLMedQ/mQXn5W7JEc7dd9iVNb+n3+rBnF
TBAPSLBU1U0ncBK1gbuy1hdGYAuwbBOgzGxlKVgZNpi4THwpkCFppyYxH3P7XkHI7iQXIm7ug7fI
QUkGoBS3YTo54oRVbLcmxnQuSFIRFGHZPVpZQhIuqPfGkW7OxyyAgLah+YLLTTn+1NtMkHVMWPUX
rExKXDB0KfWxs8Zh91/G5LRUiqenlGcGw0Sfg1IqLWqluugzImlVAZXVJ3QeP2lqWte9mpnQol5Q
ISRjbLL6cHTc4IUFc/E9CtyEkkGAgggEzwaQL9stS1TcxHsqQxIFLW/TJbBXVKmlPmb6i1XelatR
dzkrVYMwzvDbyfHYfrHAdZx7A5UYkeRN5PwKEpldElmVaUKZP1qiLDPDfqUV3HLarudL/rMW+oP4
F9zUFZyQZcaRsgjSqJSNecwN0xU6mkT33z97FsEfyRT5s1VjoRKT5aowa3MX06vvugW9EhCNJlH+
GkmvqSc8hmPr24Eyki/QqjpPuEabzDQ3psTO8GRu62b0npk4YcLRD33mk5VZwbArbDWCANHE4DcS
lsyo6t8fINfI8wiWSd4Eqs0mWlSNwppXKyO8wfHr3LxhXYE2+9s3fLj7KKlrCV+2F8za+f2ZEA9G
+BdUbQAysQxburW1M2n0lbQxK6s6QyGV08YECEUhvdL2hXAjclPOpm2c0tvo240cI+DRJKf6S2Yb
D7iyGNO8VHzF8JHew/UQvkY6efHdQwwF88iZMFwPGO9hy15syiuYap4pQLdrxX6RFWmj5KPFGN+R
gbJ/F75+nyJJ6mv+3FBUZisNzBZoOHrrVjGnc3/cMHtHHu3TKkM29EQuZq9jUrmgl7telGDhA5G3
FsMqMDgFVwPYnNg5d7wANawuNuijuC7QX603TsYPdEewhJJwTISlCoFW38YRf7WClbQuBHkzJ8n8
tYOgbi7kjtVsX8uhc+qbmUkWzDrPBbEd1wVkJ+GdstcpqZaQ12OPlBfS86qfBq5PqMNkl45UEU0B
jcUiJ5udcxYFc18MQC5faCDwFSCImMLiYItgrBnDcY/CuFYfCVmu+KRjSvhIUE6sddJeyxiX3771
Dk7PO0YP29ltpkdMboeK/gu76jUW3nO7KSlNdzWGLBSleXwKDvCU2AT8tha9LdegRZUsSBUT0xOg
3lAovxSTeaa1iYG+pLmJjM20pLZM8vrf2c+CENssfM5OYdy6C/lGUjq3qjGwmXxJQgGklcs01yif
miF+B3Oq23P99f8CXRU3KBhxW3DSat7qj5qlRqq4I6UlCunU6YRxm41EacfGUrzucEUflh1eW3sO
/IqVpkVNdph16wOVdiYXVPwLMVx6hU49Vz1Xhb0BnhsIPqcOF6cCKNFIRef0lQcuhKMUPe9gT4t0
wurSq6KS+akbLDQ1bM4gBZF+2jUR4iAI3gsGHlDDY3uq8DKoVbJb7mVNzaK2sUvn4ZgTj6oQviy7
5nupvwlOLmYRuve3b+eEK/B00dWQAZvQn6U/Pr8jsTX1wUmf+0UGYmkKj9IBkAaLTICa5ImRqknG
GB1eclYKe0do8Al5lDftgBecpKOgCNNM9pg8h13QxMm2GOElfpT0gJc4YRZwvV5MlzGkaRR9Za63
xafso7YdMjaYcwej8q4+zKuxkz3ly7UXlJuB8cWjrtZQF0AQxdiAbtBMmM/WfrFfGwcFfMpmk/NV
jjRtFWNKEahxtI3IM7oXfCMEOP7lP69KgdPLNbJq1jm97/k8fA0aCzwuw59d21d74T6YU2/2ErAd
x69zjamkulkPGLGsiVqvYIV9GWgbUd9NwJMBxcErD+xLjYfaK3Gd0JlI4c6JSz6mDnlgqq9jCLPn
MoCLGIiTi16sIZgRtGKKEnKXc8LkogcMfmOmfh3L4b8m3WWlVfk8DAW4YtVNP2Mx7WKdoUj7s/Ry
FyrpwDkXhno3equVlLzHJBU+2tQmtGMM5fV4qxUiFMY9gp8JH45OvE7Jj67nFr3n2AHguOTRafl8
uI5hK27RRqC4NztI5qzYVJuS3X4bITfZNZp+tx6my2SEPZly/TuleFdvkviRh0geVukKvbqQFFBd
FhALFskp9Q2i43hXxYYja6WfrDVpRm7JPxXio4xisFojEdYygi8rcjcrQBObk4Skec9tSj7rZRU0
Tqnjk0DSjlzzZQv8a6C8UlJy3BrMQH49zVGg0T9vbS7qyzIZ4Nzh/xJxjdOo3lmTmVYbE0YuRbf/
BVPCEsl5UCPxh3mm9x9ySKO+coZ+TLjlEs03XG0qqiB2PneOxragxcICNwumgBBlchi0AyNc5soB
zWZKW0UcRdkgfb6BBSO3h3ULKZC5xLQm8BV2pmjHVCuvqyhsXRyrv7DkYn3/+swJXMQ4UeA3ysb9
hB0hkDyFjVlrLsf/xFc9mfVGS11yq0LX1lRHJAkAZfG+ycdKTSLQSWnlzB4O6nRymxlYBKXgTiS2
Ak62Vwh6OvEKUEnHqMEHJg39NvaKTRQLfg6jeEKukzoGCfV7k122ff3LxfrnS+4xwXhUDVZId/HP
Nk3/EfWsHxoH0lbADFKEWuSHwyW3fPMTRQep0B3GSYsgEO80p21mlA9uSDznxaj8KnLqew0pgNnT
BQRKhmRXq2E1Yz4jVYby7XjOyFC8F5fnQ6Gw26D4oyZAdGZRfVVDOoO8OhPw70D7CGEU5ak6RI86
gZHybt9GbmB1NunHFBK3ZDW9wsI/3PnggX9+DItLsTtdthYDD/CTfKTkHSg+GtPVNCt5FPeSFkNY
9JvDvAeznoPJis0wHtdxilv2EpvvTDGvScQm6vVZcvn6rSQ0YfuF+LWyGaY4igJ0luozjUpue6mD
KxMLCGKVIR81HakN4P0KBHFi7nDuRsUBQcEV0cusEFw6cr4oFRkXa4mMDquBRMKhu68rlLIn6BRY
w0NBlM8E7XduVjkROCRlF7Rlg9Vub4haXIiJiRAqP2L8oHyf6XudRY1xpRxzTSPxQcySTvhN6zeU
qBlUFybwmFfAroVI/xUf4WsLBLy8wWeSvwJmdCJ4V+GunBSSud9QkOuBKPz8Hh9lj+UltyVUvBXq
NyS1YWgTfacPz9WfvTEkb1bRXg4LZBFP7DFUXF/SPkxgOYQF6BzdA2deV/7WlEkQ0UCjF7Yag6vF
e5eHGtXL0tAhGrRaMAqlMD7fGEhiChH76Skp6sAMCVyfJPQHwXxojvRQTLG2kYaaefHin73ez7Im
GZLa5nqAcRYrHbpYxUHU33tw6s6L/ZFfMiSLjE3tS04giCzgtjJFa+nno7Od+yg672Psm8erZYU8
E4JxzoVwruu6V1dppUZLIosujBksXyMkmB6Y5OKEWyyJUUm/9rYSwTQVFgCo8aCoAd/+kevSMyQd
ddTZWmu3vnN9s3qnFodxywVYOjVCVqyc3lLMliMRyMe4k5Omouy/DnNSmcfU4jwfQfaCW5IK6FWE
Tx1sQYt57vzoSaa5LBa7bMLn/c1qGwIoaTcRMTgASFrq7NpyRRFeC2qE/PkYv8LO0DgIKrkWzHs3
/ZUSMY/9ZopctboruVwyI6/bHJAQ0Gemcq4+aNYHBHZ1uK/bPniWZUT35lfd8hXTqiwjfMAw41Cv
rc9B2W8xuOs92b/UklSotVFPdm/pDDDu0Q1EICbEHup2oOZMLixDYaMrn8PMbN4Z7L1DcN4pAkuv
TCXKImuhVHdsd1C2KrGtpIMW/RAW+MkxGTHCE6iiylVfgku0xFQWjWbbaY8R9CODoSHoQ4mH6jiR
hSD+6H3VX4WMlu+b5m5SEZoKRxnIwq7nHhwTWxY1B8Rxg6eXy7e2rEb7K+fGG/UmONal9yHIKysZ
H/hfffv4wGFTb4SqYVFxy/yI2apDsOCgbLAdxfk3iE14ie+5bhxRU/6ojVk4LA7eM5d7MsvxopMm
0qDhYyU8vfmf7FhqzWFdeGP126I6gMe/IKpEVFo79+mOZhxLdgYbjX2WRAvbbqilrmMg/MnHrBcE
nWb3+S6Ibbim8oACTWsRi1573RUW00fe/RRt7yXncHg3+bu5qoGV4aLJll4Iy0Q20RqOY9ZefVLi
liPe5ktBsmh2ixuG0my/CYswp3AmQyzkI5YafOK0L4C5/RVNYYkNFzx9f4RkjyHnhOBH0fRxXSAE
0RQ1LPOH0WOBlA4vG+fOqrKkeyHImrcydb7PBxfwh9YHBavyFWZ2br28I0v2yfPnaYuwN7TpWfJS
hWpYBn2wjP2bvbEDPGB1M4eg4Re9REaKXrbq8QtQxV9/dH7jHxPiWqC4+K7rC92D8ndZgK9Ts94d
U3r6+q6oBDpbpiic7+IFRRBBmQKxlf7OpUH9my66soZPoGlk26vcQOJgxsBSTJOGc9IdNF2bsXlf
oSzWyKWAClX+A3UhbxZ3FbTtCNmzgiUQyrWqWuUuY1kTtxR5SpFon7HIf84N9SA/EzqhF6Ox80WH
SrviRxf3nq4G02U2GJODzWuopn3hYJgKLCzxNSy9XKK9VdaOT9ivPiIagDTgFSI16cqw8ltgxuzq
cDOVbFbrlTiTWHA0RP/WgHhHbromNuSuzcwXHCbCaDrHbyAexNSwQcDrFZo278/ug8wJiBwfMQSU
n5sgRMw4OmA2NwG/bh6Kgu4tYcMvi3k4s3ZImeBTRXgRIh/2y8U35yxnH+plWa4HE5EKBR/HnjFq
VbHrPw3vH4NTThRN9NaMP/SzjKtnZyz5e0No8njAu59mETWthrxcIACq5E48rKfdjtWea1NV1dT+
MKuKbl5loRqVcqgZIAzxqnY0BVc2a+T4F4AiNT9CzMUeXy5pp/E/sPs3Ux8T64/p0uJJ6DdYhIHy
Kzvt55Efc4YHX7VqqnN+Rhp7DaE+rFoO5ZxXnnwaIO6B+Vjmo9YbnPXWiAVYoJBR9Vd/XayyzJr4
Okk3V04eu1rXx1IzPrQZ9mI7xiQNqL0Wc/Zdh5DyG3AAeZCGACNeBWxlBrDEWWKhSZB+YYzAKlzu
eZW81pGERxpApoq5XZOOMmNJ2MTMh8ffcJTVMHmxYivXaXbVpgqbunVXjXZbqn8/GtVySpa03i7u
e+EPmaQSNcJ/MYlc9mqFyS2W99xRkGOJLodJJQsZ6L5BU7Hs5gyDqi+NXuRfFvBPDA9fyRmTvKJD
QLOuJuy2nsqiu+Svcll+faI8i0aV/fqeI/EKvvwsc75meQBp9/hN37tJ9Cl8gKqAzsNBqwTZNFoU
LUG176n/5ETiYe073FOVkHXLEBEtJ3M6iJgwO17Abp+q/CLPGlA3Vjq4ckUoS1zVCXkRNzV4OLnu
BCtaxqCQ5rFi5dRGtiY0a2QQWseRICORHo7QawqYtbnM+MHc08fH3qzniA/K0FgpqkLeK7jNcfFM
be3Udmj4+AGjBQM/fdjXP7a+CnfSElwKU/FcbJ3LKw/y4tF8eVpz0T2iiIKg4fcjFG1lsmPOhWWu
knz7f2W0BAeAAFHClw5LFdl1pkfsRgMoXoJh9y38MYQrGMDFTFmS7UuSJojGxjE8LZq6QuZrf3wQ
pThJqjGX1ZUbf/GinTdaPh7w/18BqbDCTwQAn5/3fbHQHQEK+Y9Unjw/znMMD5Ku2lvm8KB1xyrq
0D/jBDJEFYGpZcWybDGm4TN3/oLwZntoisH6RV5HBmOCHrrq3gnZlAccqXjVdmRNELxsYNy2OeSd
LFleEqo2DGpk50dUc9LU4oyvSyItcAVPpefIFLcSUzpEPwPOBRpP38lDqqXpUkw8Q/ltVIzNyI8l
3cfiT98OO/U0dWKx0PjhOI+5MFW5qg/mTWgJnJ2USkBm68eg+yDqMVCg+tCVwbL+fon/kiOlkTqW
YEm0f3Y6Pq8SGtb8Nzyc/M6ynfy/cCz+Nyv4eBPzEXELMCCIBrjM099+uXoWq4cSVr2HU1ma1ZC/
2rQfmkiWIqe1y5IUYMLilcw5d0QYdQRiTa/vnnL+hCmdEhMJycNhuHplqV781frDVzy7QZ2xQe6q
llPIjUjejIu4/HzqmVg+MRRAuCdl1tr/3YvN0cC+UFK/zvczXItg8FvBrLXUYSf1XwVfB7Rn0dTX
TC9W3+fRPmoTVxB2nGHo9Om9SMFJblCvszBBAFh/XGAKW5119b3x0Cfa+L520C359zaBG4CF/wTL
S4W3FQPKug7U/Ai8n60btpn/fvvlqH/egxe+dhN1mvUVC0WrecGCulOMZkBFBda0jF6VtMQMxgQe
5zknt4jg/Y1K1gnr86er/ynU+g0+cspQgwGL15umZLMjHh99YSclVWhSn9VdOBvtIvAwWRr01gDw
UCygdXKMlbKdomhpJLGnF2FCfzpg4sfGziJ+WEQlezbzUPhxI02rNquFQY/e+ieiG0TCq31CrQyB
JNHGoVmq7X/Mw06dB5iLBIXeoZDmHIw53/gThZ4FKgzb1Ki1bJbcBJpADNeFz6gQ/vXwSpn1E7Mc
J95wQJuye5AMi+wJs5mh09lam8XgNFEOP1AhekEgVLsWaG+9KBsHWCtfzIB/02lpAfhAjpiXfKpR
E82fMq2+6f/HCJ2UQjjnyNGhIPA3IoMSjyTW7fSrgMWQjjvbgFAfegrsYMf5F6Y+4/MdID3EjAQG
hxaKTUUFNxe7JtCpbwn3OiQLjaCaRuQVU4SrckG5nfUdan2E9Y4KRMNNb+WXKHCFnADmsAnQG9No
1W88mT6z59PKA8u+yOBr7VPlxUZXjlq5Gjyd4dE8TR4GKks0ntDEdjsqDD+6FVTDIJlm55BI6wyi
hsfvOXBkNnnSaXmTckPjyJOdCm5TIoUnCE7KQgT+lUZskRnaluYG3AGuK7k4mDZdcmGPSmT53rmR
c74JQAi9gZGfruxBuJvBZ8ruLWKZBW+PsxoiwcgpIJV/EHiCK1nAjb/7L/sKqnWm9Vh9z7dXmbpJ
N1SXKTz7O10p19NDmJwhpb8J4FMafSVpwtbgprKyLrhgGwTfPQD0AAffewkmimZWUrtPRzXLnoS6
Ovr1eDCgPi3ffpMkGmwVAtLdfLnCOinGEmeQ3W9y+2U9cEVIym//M9j54w/pwAs/FzIorHjGh0ha
ZBlXzJeWp0S7u8WBW5KV0G80oGa6sM5lH438X58GpyZV+o3cBQdJiq8pkZBFwGD3Jf3BOz6l3uhp
7wlG3LAKOPdJaA6fsbQA4WepYCVrTzXajPWvQBRb8ijFFB8AthYb8ANgVOkBGhe1JJcEuqYMygbD
yWoHWkz/NKUGJ3fCb+/V374wcZaIFX7TrlCbNUBNGEjZ5D/KyCboI4nuwLChCowN2sOYXZI8GWFM
/GO0lDKHPWVjC2j+Y2e9vbChKWZ6BEk81ourUAqZtbF9GX3z5mlVaVu/Nl1PXpbSs/w8uMHjMyDC
p6DtjyCdioipi2S55z2t5HdWyJ3Jf4CVajXUoFzd+2VhVBEdv3r6Ypo4oQVj4xmuVGZfLP1lKsEv
ZFGxm/fkK3ViSM9WonyBuWiyvIoqtqIqiio1kBGGgqKegQ1bI6BlSc3yiwpMJawbTfZApJ+Y1Ror
hyx8QK9ouOIrBtjstYJqNsa2VunMF1+tr1outHmxJCHo6rSHfrSJfODAxUjmokt0fkoP4OhSnTKB
RtY3PGFNlCUXKXcjjF/e97/ldKDZtCauZme87JZRYi2OrZlKZpGhRgw392m9WPhjfPAoL7UPNYJv
r6x1NoaXhlsQMGeDXdUzPPdJ9TeeA0T6m7QUxheA4suBT+ObbXzhGhoctojtdB+wKBglWC2xpbJ0
mC2ZBaGbM3bUpvwiTtX7XWa/ZlBX9+alFEMJdiQY5jHctebd/gtWddNiakiZtC6t+j5mOxLWT2EU
J8kyfxW5YNwjyRTvw+lXWIn7q/R5Z5aJHl2Vjyr2JehuArnAhSEMdgmJeIMtDRYOtblXgsE2C2yU
3w1XhOjJ00nF3mySVFPOvS9o9rc6qbxXLgJf/rB6gYBuU7QJodJOh8BkCtFWXu8WadgTGg9BXfWU
gdPVZEfR+bn9zs6fS3RtvZ+NE91vyg6IPpUVF8Nhlas5AZlFzxW53Kf272liLnCuzk1HTPrk06nK
CSXUD5etg6fz/GOjBOi9IJXAoXsK4I71jmEBkdHuSaJFw8G4q92rxtkasyj6yhmG7MCvmufJ7Z3w
OZA0Wz4UOilX9bnX6aA6Qe87nbBz/A/7w/kkTeQjJ/ZnnQlB/NpeSgGcAsTJOCbUw58QEWygT/JP
+Xmumrvv6N3sInDugO28U7yu/btbNIw5l8zBNfq4uJTOUR04birZLYSKZzkTUFYJ5AZfMNNrlJn/
SOzKVzvACPX+Gdvi0cSSq0Qir8MEVV40wksA9CyWrrQm4rU7q8e1QKLOHlnkuOoUwjFMTcIZMqi5
au4VTXV0AfVJ1Xw0wB7OU1U84Iv2Oh2AVhkTLCG0g0kXKS8Ye/MKH12Oj9eWmdbUzEHj5rLg9ifZ
LVW+HrcjlH+XyFiXtFG58VvYwD6n/hI4PLRT9vix9KexKN2j/eF2Vp5rbhiT34BInoIjIFE/jGQF
CxnCvl+dKpOHly6hQx2YFVdMGTeOSAioWVmvIpUhXqavecNesq06EJQNPs6IW5Dw0GV2emBpPLOE
hfhN4P8VTgOocsmDze9REOxU4GrMQ2U8z27ebWEQoRycoal4JZM7KwYFRBBKJbP6qGGah/T2CAGo
52hGsZdw5tfLWJlC5a74coZxZVPQAWZgwVGwOfFOfXrgOYSfnGqWXLYFaUgjJ6j3Bc9SWc3lP5li
NxzSf1raFuDb6b4tUjeMGzAQCs/HL7rAxIPU1OybZUkHZ2JESeMJio2pybF8d3NJJ9caGe8OFZAV
eXJrehPn2wFLhF60AW2F0ijmV2t128K0e5vlQY33eGuSnUK8R7rbkNNwtObK8s7aLZI2lWOgPJbC
9gc6Fvx1i2vul7bk4Xm4S+VIKpryLADJ5GXMdcuktnLSiYwuFV6DklMRP2QjsOO/lq2iOcFrmV7V
zdMBGeeETWESgfh+Thi58/+pZ0DTyj33AVfB59E7Lu8lBPr8m0GvmZww2PMhemjxrUyBzZykQ9Pt
MIknxWlFxHGLdcncqCah9arcvsU2uft5qeO5hox4pyEyW1yoeL8JDMt3x2+n1k5pVs2WCKD89y7c
z8gLs3SXg8jc81JIZyBHVI9+tBeLRGTGSsn/ICuNqXJvCk2xUhjGbjVMpIu7G0Lkle0WAvTpiM1z
pF4zau/4Xl282KXoc6XBDlsJzJiWge+jPVondj3x+GXSZk0VVD6xTeh8j71yefUEKRNmHhKpGDUB
DLcnLOSev8BaY5MYXKBld1U71+px8x9zvh9HOuSk3jfycNoIJFk0H92tODijsMDQG9RApBVtpuq3
8jvjw+WITngOfB/CV95X76MvwQrJ4oOYMYtQpY4WaXKho69VTh/F+GIbq0rcIXm6CNMKddkFK3ba
dPFTAwgHAsu2fpecNAAP63pI/IlSujlqw8xHPRYGK9HBnuDR8IKA9W7P/qZGwfIFxgxEtoissk2o
ZdvkmiLgziz2lh2hPYNOCKNaY9/p93fyHOXVnPynX58ByK4E5pczeyhOldGoTy4HBbBSMJ6yHEfR
2CtGm+OsbJjQHKN2un4Md6uioGGG9iqz40jbMIew2IvX8kOW8xcFQaEP8tTfVmOIgV4PfV6oax24
gpfrkYWlsHZUhkoWH+c8XI0cO/rcEaoRPvhI8Zg8h4mntQ7FVwl8JstG2Qjd/HU1QZa4eFFz/MOz
aYO57/T6LNnvMz0zlP0MAY8OL9HaqbzpVxGofzvllPUO/soxF7+mil2UnAU6noq/WNneaPnT1Wlw
AwKviYxJVAdYH97OWdSYPMgMZC9Liqq+wYvCaJdzAvj9NdFOlcDa65tgTwfIPKgmHJZYF5FH3tai
IX9DfaMyiZKveI7yACKAehU07kSX1zBLChneSeE+rEygpIHnRSKhzndQueyR6OsPc4x0ZpaXg/qI
ehPChYSfUELgvQpCPPRG+Eet8GxLNMuQrsyfHjKQYRngLwLV5nIlb089HgEwu4FTmLb7MSUpVBH3
M7PioevDLlsq+aFzdb5oDAbio8LOsS+uDmwGZciA46Qmh1hzlQMLs0qzcrEJ93NUYlcPKi2NedJR
UR6SavV7SLQROMEE6Q5ClZg4DS4bzoIbVSuR+u7YFqFXbQJgxzILTFxXwjJdIZXN5oqetZ8gnA6Y
bkNyG6W2nvZRV3nmB3o6qx99qNmW/cLlrVyMblsDPujuIWuDoFtEmzzTd1poqrWSYTuFDpnIsxDJ
O1Ffo+QmVDpTs0d1oYGNWPohf62ZiaYqkPqU2PsZh2qLYO1hO1EwEmi6xhRl+8a+x9ZeV27QArS8
20Xr4hLd5FtSqscINNb85xxiZOdi6J6dx2Njx2KI+qgiMdlLo8lBQM87fba+EhucX+9mUgUmRjQg
m53367ElTpxLaYQfiT1q6Q7dBwcPeo6fT+/UO4j0g35TkN3QnKVnKM8E5WYwZ99KUdR9KNUT6l0F
uClABPkq4VWzTFqthoICj4OmHJYWCGreS0HoEcTYssXB5vJfOC9SlPOKHYAh2uF9Mylaonrt3ZWU
j3N+MMrcGEPP3INJuMkzyatiVBC4O1/9QY2VBcyZGDsPYxsqdstrRNXwzeINmtnUD1bkoQjNKTlJ
8Ce0z9ZX9NkFHDC2t0YS3XRPajRi+56OC+RSVLguDZK6uSAzFpJlKHcw8sTJgflt10IOzwQAOlxm
VtAIhh7jxl74rtW1aica2Gj9IpSK4xwPk0jRguSTYatm0WbRrpiEiCQyUrNkSWN4hDoTSlUtpR/y
NQ5INde39y6SyHbeHPyNhGr/semzcEU1G37gLLdE5r6vDss9Z7WxbMJt9ZIuzapLZWJjYHwOa08v
E3p6g3j5uPCXN/r3VxgQoINAbh00dsOFWaLjseYjdA+AlpQOXwSbhoAO8ad3owcmL10Pru408PdX
dYfP2WhNyTBbN+9PlZfayIBhCfc3sju+zsG7WuixwDZAKavv1AIK3Y3/eO5Zuzupq100SaTAxEul
ePoGt/04pG8AADDHU0nGQrMcpwAdwEATeupgsqA2vHC4vt7TdxgmfPSTK55xAXICYIrDQSoZ21TW
dzn1i+R+Xce3Mf0+HV1A7Dz+2XDSNgpM4V/wCldhYHA3Jj2wVG0zTUEvCXQihs3zot+JZALn3aSW
8U9ZMpEDFGB9ST3hqt+OBiEj6Up69rj/0sZ9lhXBYQiAUTR0LLEAolUI22afPlQ4Ev1eZ6yNIr8L
XL5TpGXl4tmL4qjBczkFMpIdbGvO1ykBqzwVyOwmazLVjWrCqFlX+2PsWFfMZs0cw0mWJ/hZpFr3
cQRZjlexON+tejPCdjHq2NprKEB3SCv3eo/77yCKgRoqAX3DLHGR0LWrIJYzMbq66b/oRam76BRM
AIZXTxf0MxOyYtt0CbadlTY1i6L/5ETCJ+VM0GY0BSJaeSQXggsloB+cKgMA/KN5HWDKU92QBeTh
LeQp/kLbSqoSXQNp8O40DjAxKmfJIGreoWD/oGleoafGeFB6wi0HhHLegbs74RRfZxpAmyySX00x
qQGnlRDsanTG9gUISOFpOYYF6+XuspkIHnb6fuqYhcz4KfOXG4cWguRJw6R1pJcG+XC7nZpJYdbN
cxWB9ZetgyEdB0Svx7SPpsnA/MLNh08o5SYHkHW5mLbSRVP/GwHkWL94WF1x6eh3naTcXe4CWrCG
gHnQQU75aLJLaDueoCw6sSlvFMqorNbLOg1S4MPE6dnk6olrpsTaix/YQ/+wh2fwNuDT9Yw4m4I/
DU5ofdRMvstpdPUodpB7M8r1YPfwW8Ib/o8A0nTkaOQ0078e8kpeMR63ibjEfDfU+PLM858GoUre
Spyr+zNskjV3XA6xDPUzY+0h2hF6wg8nStIJ6xs0JYu9zCaRM/6N0zTWdUJqVLv/PFbVH58B+SOc
WcxnfSmP4hgfq8BBprXoQyC4gVOt/L8lMptwB1NqezjlCN7nzDcmf3AuOyfbwku1+m/CM6enrmot
QvMBXOQY3sqX41bDtvY+kbWp8O6XP8iB5pRyKF05dDnXv8M3vM/bXlxayj5Nir8i4Eh20BSWtq/h
bvFcGgdvz2mIKcHxdt2GePCGRXXFIyVotEZDwgddtikbtY9lr/I+fQj2xMJzOiycJa/rBnrmpu+K
LFCMuD0xkan3/R8gHYl/TyATD/8JWHI0xmqq7rzQz47qfglY1Lov/gqCqT05ztdwSmcepj+I6fPs
11MVheos2cxsZqjqKhubWtnT/NuI2Qvx4M8mlmwTzdSpQ0kDndJhxmmu+B0NY91aph7trC14C8aK
Ct18RtXKnIMENKrt3IcqBcDatbpdQL8iXaLagtLSQLVjudHixwSKyF2zHFJQVTZS+0FB+aYBOm/T
WuwJ1cXAYJHshN7niFkdEI/nvdBlI0kL3U2hSSqGBA13XmI5IwNr3vP46Ow+johm+prwj0LlAEAk
s0W01a3qFHJ+GqrRmiMYpmyOZhgpNfSy9QdG81iGTJQADkraCeVs3l5um98bvPv8u4hjpMBQoQvc
5aDxXUeYeevNEuUns0t5l/fIYuLiO1aSA5ZnJb4AHqlUAKhwBB+TAr/lDVIy4xpKdrNyUjVom08x
1v+VTXPMiZ7+fXswGTr5P436gIYozmPea9NuCDHHE9l43UnFShvBL30FSfnPCplRWUnWYRY9C3YF
ytPq3U99w8yKLU56Xmaldcb/+QPegWjNWE6yFbt0kkSvJTbMBub90Lk3NAwBtSyji45o+N91gmKj
AEaY4qQSKDQ77mfOPIqYlh4QwLzs0mJyNsMd3m//YiyZt0iG1mO4ZDLS8BaX4cI83lmYeLP1qIhI
JHpK/VJ8htvn9TogMwHJU6jZ9j6mIfD0cHtLEc4fwUcQvPX32brm2TRAlc5ci342ONn2KA4PwgLo
ugnRoL2O6woMwq6TU6d0+CG3zj7+RBMmdNVD+xcW4iExuID2b8+ZyyY2oN7bhYxZ8P1zEWxptxUK
5f1tpt2x/Ki9HAYhQXoJGzIojah9oeLLDLeSoUx6+N+BnKkZUWbQfaV941Rmr9xPU8S64iK+/4Il
ZT/6nHFYvUTts2nmJK15+OuYcQDC9g2sopbPcuL7Oc8xT9/H53QhBi2ZNnRtIPkLmgnI95HsIdla
EkR7FdD0C6//w03t2qcrJdbj/s6iq7UnbFp4jerKwwSW+PHgljSp5NEnSjxxsOEdw/ZF1P69z3yX
14VohVtzkLuooFIduMtbWSQoOODGqLFOlODE+d7/tfJv/4Ft6jINFLSrfa8SLUEHzZoydvT1/RmX
pwrcGUOX3rNkWcddCk05HcZnQl47nROIF79UezJyKijlHt4CDVTVCF0mGs/G8MlirGJ8tIc2b4wj
pD+0X2CrkuuKODhoIov1EqHDRjhGWwrJJ5NRBpOG1ACuL7WXR4zIVrBzFstHwBpK3VmHOJLq8FGd
eYcsmK1fGv50SofveTd7wa9v4gyUg1NPr+pN6zZW5mPKm3gJOoW/QItgCksptwvM1azCK4cxU6i1
zOlmR8TyPxK6KBjK1Iin4EcYfNzpcsSjs0Z/OEIN4X3b1rueEa/GbDeORBNUjUO/JPvEooSkFFK3
QAsLrSaM13GB0yFawSfHcGxWrXBOacGcrjYR6GBeTVvm6Tnkyil8vkehF+ILRLX9Qkwfcdy8RjH7
a95j+oM2p3t4UkWe26AnlgqyjwX5HXGQ56VAvXBm6602farOnA/gBUyqWIh+b9ukJTqMM7mBz+s5
BmqdJH3Q22qjSGe+TOJCvdzyk1pKPnaDTUp/735ex0UmSQC94TZ8QiS+ATNvo18C8mE3OdaNk2Rp
UfjUWAv3j7Oi9d+TXrWTbcVcOxfdNsFjisS8h50mVqSjLrVfV19zWgBbnuv5kltMJHfMVXThucwY
+WY4hgU1TFJMQUAfT3VhaJOmI4f9hfmzKJdJ3EekaLDAP3dWaPPuBMoA8GAickFYcf9gbfQLwix6
/qJtg/rHXCoTj3264gC/lobvrfz33j0Q2LC61W4pkEeg+UT0fiTqabZrqnRZHg3iIp+TX+6EBryo
1i7RTwYINmHo9t/2RmFf2l6O6HW11vJg3uk+9Z5NXGeFxIoWrOA5tjbzlOIjVtekEyopvKtGN5L7
4y2k75Hbkf5slC2Ip1TVGBr9oSHrdLFp+ZOD3Un9BAxN9iWTZOsu5pjwfrUIkUgGnvjXSmp+9mHa
BNcazcYn3SoxHAANhzfDLxV/JJHJMtw0sC30I5pN9F/AkpnOAib/X/rsnZUTddnYqkOWopK3xxFv
+3o8BmNGqct31qmxSy+H4RGMitUdZIBxbrs+kcb+R4iMJhiCZ7o+8EA6GUReMp7h4JpGAtvcQ4ov
lqH3M96mRjDhXCDwxo4tsHZjSRkRwdZhSd56CegTM0hmiRDHYT3fFB76XQboZsBBUX9nCKEJBCaw
+3v621D2BzXk11LY2dtFL5jrCVFxPKPujVao5ESBKQHgrW/e+h7Qja2YVISFMX+VLbIWUbXdnsRd
y1n8etuFlvG2VHs9/sqi46shSIKu+3UfcuJuW0Vc4WdCnT32YN62zte0UcHhSS1bGx1JoS/fKHO6
WlciRt+yfOyl9xeg4ft8gX1bLyow+kykDXoYFFLkb0IWTWj5KBfB3BnmHJNlAqtdtsCfWrASvTOk
Wr2irlL/tsz8Wfw7t4QPRotX8SS+wR9nJK/9DBFG93e12WxvXAcdqw2JOaAwX8AXOp7TGbCrYUhf
9RTLGEKPm4DpOxBtUxGvkHe77SyArnbrG7wvMIIe780ngRL1QdCUZUy6aFw2IvrwjWdJzYWNszB+
dYIAYr8/bpTBI4gj5Rhmk7maWwZ3J+qqsjVTcOpFau84aFsKIFmG+lHRDQKIr1BnFkk89F/gaZnt
Xpo/vwW/YZ5dP+EF25iS7Dko6Uixulkc3Pe3fZMp3nM7pL+HA98MpEffr3KR7MvZccQMDQOW3dSd
zDBHDa3vvoLBt7U7w5fWPu0bsECpAsifN0j1B1LP6W4Ud+th2gOKzZ3CwWFrbYEItdpcxFO2q7/A
OQ2qXIkvx7+j+vj9qE3S5Oc0XpxKshfbBmH+tw+ZiF9UV06+Oyc5QBpjSOuMqRmvdfDpWZhtitie
xYMklArNKxVGigyctRMh6cXAmcsu1VjIDe5mHdBiVskthqyS2EU/kTBUgI8ShhlkprgXwB6KlZPx
FzPYigwYDJml6l5o5cTYD33PR1/lfvGrCcQsWRrMVCI7Sn+/IYUQBZHrAcRKu03jxAx+J+lsyuJ1
n3IIhKWnuvM6InI8XxILRnZihPo65ewqtBnI0WuXf6sql+h/QmGPV3+/vB/Q0mIAFqT5n+nFEXuF
mPSVbg5KtNyHBsIWLx+jrjrs3ZWQ9m+IRBgTZn/rORB2OgnMH+RnsLUNqnCjeKY6Pt2yaRGniLgZ
5FtDixy8bHdvN+ALdE+kPZpbCvzAFPxv6+7AncrpYGKIXncJAY/aVfMMXoCIB+KutA1/2lumex8T
hbRYSjF2E/He5ob/H2rT6yo8eOfIoot29Xq34U5oBiT3B5t1twB9YkapLvKbC/qqjBfum/0gvG0a
wzy+bpNvVX+iv7896Pxpbk8/ihiHsnPBnuvpfDLHXGRaEjsKu3WHoIikXeEWK2fCQSQjCRBHY72e
BHRHzaPXMiKyQCqfOStzDQeB6d5WqQN+OD0t5r56Uy1z9m3+/hlceqD3mQWzhOyGmBoEa9E/OXOY
aGI4jqfq3eHWcmXAYn12DX75SW/SnTaoaHEBOzNwXoo+bGytKFxiKWJWwxnfhEOa8GtyEwVUPdvL
LF/UcY0i0nQ+nEVojd9bugtueIqxFzSidsADur6WDE2M2SEChn6Y8PCyGSNqDM7ZHsZI6Pxx+aCz
bk4YeidIy0KpYVmWK12NbPrJPa7IZkHSkM2TmQLDmCHGix+/AC5p5UKXlDt+aa1zrim3UKNvmSPA
F8YsTJlQIUCBvjywVPdaI9pebOtO1IYSLtr2SVGZLVTXdZsBntla+l6AMZQZKy0hEoLJEwuHADQy
jKzXYVVCtNNt9MdJMUcsCTWWn3e5D6aZPcyGSdk+UqlAta8mpxI8OBvablf3UM7Elf2Q36d7NYo5
MJV5Lr23jvI5xhzbkQmjiUW+YIZQsyfm2C1TyTUFIt7OdRAFq+oNbSTLQLis4IQsXgf/ag1+Azaj
lTG8yqR3Lyb4r9LC1XGiWp15IGLSXNuyQwO4E9/ofC2h/qfJz5lZdmU353+zTwujqvGKmBa9SaC0
yBfxGSytSPMkqSThjuvxXOrcF90XeTHR29d1nvtIrSGZDktczBy1FpyGM9LfeKZRwdp/JJ5iWRYY
MLcWmub+ZTxZuiWTQSu4aZEbc6uwnLw+PSqfOncK3kvbHnhlWH2AQKAakj4cAUS/dzY9oD2siqzF
MMxkBDSbdV9zQxpSR53iSWOVuY47sPmsCjcp208fJ9V5+XI8BDf3t+fNpic27I7kA0+/IPjvm/OE
+aB9iyQgFMFKEruECbwb3EolqrnqGic3ZKudbHCfPutNk9rtG+ExLD7/ZEBm82QrWHZSDxzw9cKG
uvNhrpUvqakR0CS9HDwhcAjmOOdAnyrSoSeuK0Uaz8vzRmK06a8frY7O/ncsji77O35QIe9axcS3
6cbWUGal8qSTLGtRNDv2sgJbX8ItQVIv+ZJfpa0aRQWPgqpFjTWrCtd0fhbNxzW+1oPR+sE3daCC
NRDLoc8beIiWostIf24WO21mEpFhxdGNYF9gcYHN+iW1iszB4QL/zH8atKzyG9vupHIKiVLucTDC
7G3IZIDy68/bnLkCEY1g5v6wDPweajnUOfFJTQAJIjz1a6x0PlA+Yc0aVTuVrgGR0Ar86vS8tmm0
+tSfAh1hfgQY9XDmEsedm7IMeGMBu31OKHHeom0Uf6W5FXAqW5bdDAr51J2UEgDLL75f01FTiN9A
+dqIGfL4P+66fRyiA0LFYIGX24O9u8I/xuZEniAcXrPGbR671mffLY5nhk/d2AOInPksswc8dUBD
m1pZiFiKcvHNlv00kbq/iaepkyyrKNr4g5ePbUpZJiIYNql7ecBH0ce7tjnqpyj7tsyavkhiEaYh
lIcnOXvJbgkHPgZwban0VU/9C5ohHj29NGlXyNDhijebwemCUhMO00vroB2kGQP9eXbQzI62Wrl6
adzg12V+jiMJ3Wnrpy4C802auKIWUtO8xM19/MB93LVUDPo2NDvnsBAAZVaw6ICRyA98tmVnGOMh
+GaCEMB2Ua1atjsX8e5x97rCD3oUrql8uvTM0U5gWkLWCaM7v0z8LJwbbvDbvBs6vDDWSzBO1JpG
7XwJp8HzN2qK7Dkz1h5WWUuRV4OI3BuPmT4WqkBIpWWvMFOp5Sy98Zj5el+LaOWFEW8QBNHuovhK
M5nEOEaK1hiYzmEVT5mrVdJdexNjUnUGm3L7vvW9x1PeYfb3+cw/t16MGjkuY/6M243zylwvgkMA
9dLhLNdytZPNY00HJUExQC5O8uoSeuMuYC9X6aRx0ShQ5L8Hb/EefoRIpJNC/6Y410pgJbtz/bZe
2GICwSTkaCSKR82jLnS1lqSXHBtAQ5vV0qIqaGjxfx5ncyYBnOicENnJvJ6YWe/P0UQdFAL9aXSb
+UJBdKaSDzjzGDytMhLkFHF1ztZ1HOeC6If+y0YJHz8D+DFSxExtRPR/ibX61cNXslVWLFH3cjsQ
KPQFveo7eITlE8sd8PWHP9Ren5jXln/kZnGbt7B1GYf4QtY/H+/CGQix+Lc0zsld4H5ifFdVUYD1
L8jEJrkAoyWH3+H2froJILSuVY0XqmXKna6PWYJYyp6a6HOXQq5mLqZpv931xGdnTdMd8JHREJu+
Wui9jwkFFEGeZg4hrjdZfMyA3gV6le/EzYWj/C+nyGjGNAV7fRazo2WJxLMYVb3Nv7It6OpCZ/l0
MPjSDq7ynURHNxUO3ZhyqDPKLFv8Y1RNL53C07wKjfcToP0vAKy9Purl0ATqa+1f1Tonlo5yydk/
wgI7zD/lEGKTjptA2f1T+ainxJ6nkvEhJsPHMWrOBIRNEeApqSdKRErJqlxxxQm/wbCKS1UrqNki
AblvOJiyVtk3+MjOZsgkaaXlE9ge0zCp9FPJfAYIzVVNqM/Iwg6KmAesKVvuqHO1orA3gKZXVRhN
IAmZI4vdYhJHt49XaS/uL/r/drlRqN2+I84hmlsLkCHNIN3rbGPyXCzb7HNpnMaG6lPQuC3WNOyo
DqnO66PqBgD/IHa/TXv+qMeoUPi1rBEeaGKCBpUL2k9+SFisgQFeY3qSwj73KREgVrDtI49CAqVY
rD/t1VRXMIYGqKkR5be0Xakgdpuy/vniXhHmvYdQE8pSIMeu8m7YBqGmZkBmtcOL7LJuGLDgMrS1
ZdvlheA7TxasGBvIeGN8/6W415tVOaMgNyDI4kGyBC18D+FN1lt2TTvNqMwHZJbNpANCov2D3O3f
3QNVABQOn8WCG/3INEZcW+YE53wt8Y5KBZrm3V41bSsDVwhGgUFqvGwP3Gv9mMmak9Npo/5lcotH
xguNQ21GroYHT9ABUas/ciPwuW+oOf5LLc0y2UPgE+60FVbYHuE/TMc1mBEcXqfF6F3wMT7RaH1P
EVbnpTx7vUc3bzDyQpkfv9LJYN/nRb/PRrSQUilDk0xiebXWuQnmDd3zYYuDatLrWBoJ4QXUupxk
pU14z2HLySz4mcyPj5+pj3F1Vk18kUHT0G1NWe2S8D9477JTh91PsLkxiLBEYDCYwpwvSIosKNCS
vMHJGdQGwR1DbCkkloNU7w7t3/EBHYsNbLeBpqW9rp93Rn4/Qky8D334ZsO82bOTdMVdSbowSkeM
sd7avUSohqBgF2uhHxVfvlgdiKTiOEneAv99CdXUmbrT21SjaLECw5/y0vY1wRlzNBJUEcaSTC4g
UgZHtmGJw5+8uFVXIv4NeJK2htm/PDLS3TOZAhc1k6cU9MephX1MGc6OyiWeq3W8XczLVzFLA4mG
PzS/qsCl+14gHlhmZzlu1ePTxglkkpc7DwSsrzQ4xiyUslcRGuLHomtC+mVb4yO0yj0ObSyQIdYn
ghd2kWl/+PP6ND6VcRj6b3DjwdFpSfY9DCqPv9ihNITrh06sJ13pqwDCN9Fa9vzgnIDWYPinx//J
TL9KLmwY6ZRKvopNkDVErgvZaIZze6iVFGhuNbbBpl/IHBIYbVW8Ilj90/4YIz+gl0zjgOxdlRck
vlpGtL+79S5ANRrJuZUYcHUumTRG4+JX/dw7K5zD7kIQoLq93wFweO0pPa1cSmcyr6qIxp4LtfJF
4Si05fehQXgvsmEbph8zPBYZusRvH8nBkhbz0Nxqa1CI0DI5pSeR4qMtkJw0V0OiBSbTt2TOnehE
xyw8SZqE5lRMyfXtUY0UKFVcd+dFLsMWBbVuiUn/W5xwQmHUVxI7F9i1ycfLh9LJCIHUhroVa0Pe
bkFYkvorMt1WdbA2bdTELy3EQXV9QuEBUx8h2hFROD2bnrygAiuK9MG5i4pMVbz9+6MN9fMZWL/J
B44qvyBGO4SyQLtut1rEU1Bve4+/GTV7BrEPwUFweMSDOqP79fIkJ/t3NwiZug8JE0Z+TVaVCr7b
gkNmfdBZCFQk7ghk7xkRO8U4tdTIlTyBOGZQSt9uPzbQXyhiVKnqcge3R9tkAQptgYaoV+B3q+9+
APPygCQ7CviQXW4l1VYsMzYJ+xqCnWbQypn7HI2TRe9g6xBnRvxyKohYeGRvjqUNygugyegghBPZ
aVpdZYoaLVMaRBz+fmJiLEEt0aRj2Wkvq/kOb6TZHhoUL50MjpMCfQx+47vSSX+FgU+qV/YgYGtU
hHJjTGzpy4eVojIc/MF1oeUZU9LqVWxsdeaWfDBsnST02DpW1LKYbbatqapiedD+++GfMXaHWUSG
j9z6qdezvIWTTtQOI5FcbjX6r0eYXTrZa1F04ncTLOKEofC4V5gfcLwQYcJzVQvyfdUeW5+syTSN
Bci7+BvRW72rpUwBXRvBCtDVPhLMfjth7seC3Cw84Bwwp4mai7b9BUhAC90vCVLrM/rixX6dVwtT
oF2ELdZcN9zcuMjX+fm7+ainv1+SCGrAwW3pLuYNjioL3vMXUucfM0h9DuqbVGDncP0UkTG/vrLl
tPOWu84C/kjafLpG/8hvoVqoPYNOcj3a36h5IRXkFpRfN0zcQgP2CB66egsvbTCqHubXZ4Alb7+Q
k29yJ8aJFutZOEH6cGCxiyM+LQBVx6Qv05dLwEz7VtDlHWS/vIZ+vmXOdCDXjVufdv/dTMzNvtHZ
Lr9pIE+eYzTg0Zl2jxt46iWskCfACjLhScOlXW3drpjNVqcdZoeHE87fAUyjmqeYXJBqIEjiSc3w
wWYwisHUqmOBs9lMb8KqPZ8PYDiMniXlykDX5C2DhCVFh1YF1KNBhEIGGKFNhHcntqRomQVJXCq3
vmCapPzTlzDVe6l+xB7tt5V00MjWxOLGRGht0j2RiLNJpU98ErJTnYXqODyb55JuS06AGpBmRI5z
hXgOE2yTJcG0m85lTOqlHC5WMBY+cAfE252d1rDiqPguLHrMSNsMz9WIc+mehRxdGAQWjvCjQD3q
jBj0+4r83uS8UjsWG4Psxu8heKvAr31kt/fg0WPJpF9pQiMrBhTevB1cxOafvB+xBrndiBT2Mx1Z
EdcMB0Zd6zvgCdRZyljPrA5oiMFp7O9arGwp5A9wA4JQV0InnXXHcINyI9l6IRCyf9RWCZ9Hlhi5
x/BaCe6S/UBUTwpYbbMJxSxcCDuo0rNDsDq9lETclBsGCuHdbrwLYr7VC4foS+vvlKmYugoG7ImZ
MGma9wXf6Zl0o5Y3LKntdREhY5i9vC10zuDLFODN77X/S8QUFPVNlYd3DZQ+DsomrRIc/D+Ph6+Q
ZCgb1QTdY1wV3blYLCYZWZOLqSoNMtFF1GzdFhCjcTUsuGBQT6vtDzw0fa6Bfxw71TcLX8co2Vz0
JbTtkGMd1NCOQL13qKTqmmOUa6WGi33oiw+Rd+TB5XvycnAmYoe4XvX4u+tzR+DcgNdQMCnd6ML9
H4mKqGAMxaJRaK8OKMCbAvoN07kmGFrjXogqTyQfdWP2EQNZwGX71/Te42zchrNUwEFkMaoFbVfM
l6TSm4Lo1hThqQ868j5jsQjkeeeaee0EZSiAVp3MpZHLd3mX+edMN/HeadoL0mxo1MOjGO0cJ7bo
zAtaZgAy9mAMiLLZEj1xVEeirh7hxPpjr0/WjZ/fnro7mNWx8crgXWBFC4saUXX0RLyfmfGkTj2K
cW/+4hpoM4tXSNh6KuAvs1EM/yG/+iu4QNNukfm/2rooOg0wkt510QdDDm9wD17RWUDpUlyRyAdX
QiQOMZz7T5l4+KExFrC+4FJGX3vj6DqcUOlzf0vOhuQwI414cE3wWQcTZ76xWROCLlt/bu5pvH9n
MT0O3Y5CWvcEh3hGlR0rZZctkgeNng2RzjCUcj7GfgMtj00uh6qEZLxUKaVkFh+rkD34Mg8HOT3s
LkUKessQc0yjM3qJ6IKP7BMC+OW7uLiQTy9/fStBO6l8YV2FjT3iwyDPVlXoRGdhY5u1w8VD+WlP
DHaSf0qtp2n93WZ/X3wZC3S3HrMEtW4tnIYgzXRbxjSoyFHesPKxfpDzaVcKgeM3iUOYcURDO+6l
cuX5p8Y/jT5pXuJw78Ro3t9SabnX/mx3X2lMbyaFtTUKhg1a8T0u7l8AwYIvirSx3TG14HPwwvVZ
+egCA9kE9DxZGM6qwlRa4Dj6PHoe9b5GTJiQy5I3SN523+O4vSwBL7V745+z8Sql+GgpBUTEDP/3
qcCX9XX/Vy40rAen+Gmb5Iuvb5kXHM3BRZT5QpwgchyOiZKsqZfXxmeHLXUScIJOx+ToWEXhaO+g
oThoio2aBPaAmEgcGLdcMwEMMOsKKtYm7vK8IXf0e0hK7WClFYZOr4BP26RtE6mryotkxM/5dQy+
/NMfBkoaM9CP4QmobRwR0CdDPaDTBcBvx1ofGLkajHKQgcsyw9IFCQWNwv0b6+gEjKvEvGHtzDV5
OybFIU64JDpMYgUMXk+k9PsqLci4odkK/HX66F0l7bmnwf4gBgevm9oftsBqFrjqBSCkvAcfcBE8
gH14jemHnJMQ5awmkx9hsHlqUxvk9HxDrbQ5F9khaXN3LiVBPYHuT29vUZBB9sG+2ajiouHVPSP9
dbYY6YmnBV2PgjWaiWuXv1TzHM4GOiCC3AE/c7SL8sUutHOHwcFTqgBprAdj1gOiLblwa1TyAWMl
f0a/988ct+PvO2OcwVYWf3qCj7VrrmOmQtg6Y02yDe7Qabzu8gsGeZmoDDRbTT7ykrx40r0DVtQB
NAPHZWnESsoowZafsTAfkOd9UoyroerzDx0+lQVyt10Up2xTKa1mTinCy4U9sZP++IizyRXG8iYF
jdnuNuvMuytmALXFktFG4/d4yT4m7JYlqNvwDROAQ7/TNF1cSkH6HBdY7EUHvW+UcOK17QLts1j3
SzWvf+2gOOBGDyCUSsG/LKTs6Mt6VB0lHPPyaCTidZ44LBQVTKsUb+Ic14mDwi4Fub/N6WXwenf+
MquqVHsb49J8AidQvrG3TfrZzyXLdTdE4bjRctETzrmNEAGB1Z1qZ0wARIMvf+c3+V8nls9/VaVp
kghZT3z2MOG+WCmTaxsG/lVmenmXzDFSG1YMbFt4vp421Kz+NfG5v081MtgRrXAzBnzyYYUxl9Ic
vq2ui3C70EjtOq63H8z6Agf9iHD1YC1AX8zOH4GVktLeEhsm3VPcXgwaJXHfbZA3ffumL3rD4x9n
fzjb/X0XH60YPM947AA4x9QP27kr8Q+rtPwwus3YWi3hMgU9hgEY1Z2t5ZO3NaA8+5uSjEjKTqk4
eIut/LokAbrRV1wdqUalu2WGvt0gSXObRtTiReU87PfJN5NdzX5CrcUJbVpEm+LMBsnJMBPYAqf5
WaihBQGNLkV7auSq7Tr20veNURhY3KaW8PMAffVW7ewp+Guny450mW8DO26APjoWE9kzdIx4JJYU
We2Q/VWu/tM2TCDDetjmHyf10YYvPzXyI+TdqKMdF1WSxkTLDGmpSmHivWhUs9F1anaiIkG3vvoL
H0bYl36nYR/ClBORU9qcx2U1C+wj+cB34lgadZDHIguMSqSqV2lTi6mIgmYDB1yikxZBW7ojkG5p
i9HXw3+MCL5G7hq+A3RO+SNBl8uzNpulDCEv33jFyFnfNoQ+idpgRnprDDOg+lYdi+jXGEPYDtlk
zqTqPGvlfjYQBfeD5E2Q7irUdmjizwv5NT7r/7e8oSBZO40pWXA/LV9JS81AQBMXprhdVN7BNehG
0+5OgtJQi98muufkWHbPD4wbr9SfHiB1CGvPf/pxLS7f+dp0qfwzpKAR4yI3pCEphUB5WX0YqzE/
jgoZEFpX3FtEAZFjw1KpUMJIvSefg/MyzdXdKqHA/foCkdXJKJ9wzPIHy0aMBoFszx+D8sRxsoG6
CD5o7NTk3MUTChcMuhBPz5hWdWK5P03ocN4e2jnFzHQoiQAVK2D2H7j1SnRkbWpyo27nofzFcQtg
vStwMze2VV/rxhqbnG/57S5y7cUn0vbFT9i9nHuppP6PpFtzVfULnUjp7gupbg3xtRJe+eNg8zBQ
+iIBn6aT86xW6T5+5roa1d9OcCnnAdqhKIqnRsTXNSwameeAp2/V8T7Z3VN8+H1+BqktPKvs3S6p
N0X9hh67NjiSic1rQBRHb+ETl9wyHj3pycR0ErkEoH4RkMeKAc3VqhRNd+AoUkTcGglxeJtwgEZ7
5L0sTkKreqbHDd2853+F+yMj/C3kdNXZpz+PecuuyMjoKCfRwVhKwUuXkpmWkojOkWAN4kdRFDtj
dX6IyPYN9qxPc3Rv+UYSOBL2wtupQQdeQlmpr7wuQbCqQybJ27YYW/iH8mep7s/dgmi4Fwuvdpxq
SpQBbjWrLORu4WwAuBB/ojaUkdbFxVZmPZIKlELNK4Ch6lxsZWL3PNioINhx0p3JqIkVfbFHvqQW
DTTrjwO4TA9q/6/c9F8Us+v06OJgzhjPsL86NgMh7HLYWGwgKYRCL93V0zCBIIyzYf2MOWZKpvCI
sautpSALshM9HdmbbKEzyKPdCnN7HHI0giQxqhf6NvczIoE/BsQXiX1Bjw7EaOLeX8ZNQ0cEbF5k
miZsO/X7A115S08YurCyMhTYyS6+L1pakT0/u4fajRZNcYVjRxyfLpyhE2em4MoHxas+QgRXoCHj
ht3x1iK9IM4Dzxkbp5KPh0gYCPFN6WKeBjIc6DfRu4yuiAMy2nI9thZAQGdr1GJku7G+adlNXJ9c
omLWJ1ANUsvuwCHZ09aM2OtFWZuVUXjUKg9Wu4UWAhRhbtBmrXcN8wIucXfFT4s0VqT4i5meBneO
ZtxaJ4qb3KeAhTuT7J9vvuSQEGd42lJLGcWopDB+WN56VR66/qRQruNaYVAfiaMowgC1wJy3+KrH
B4BHYV6w8mcgh/+3yr04cfcyg890rrZRqYD8zazRVVM8QCAeVmqBBBE4JLYsDASFpfbCMVzXMiGU
BjmsjyCvQS+BGfd8cYkKGiyJ8s8QLD60K5Gcci0KwFDoPeKUk2K0AcShcUjyq7DAXd/m4SU+ZpY1
4fEAv8ba3I/EPNYBZfF5RgIdDiHEd+SjApjYSnqKSEWx2BgA7cGdVM8EZZnwmQ7Sy0Uoz+oU4XCN
OusCQcA53Zwqc6m32w8k+n80IWw/ZnTpEowQgsLz333zjlPR7tFtm8O4T2OvVO1udk48vB1JWo+n
UehLxT5GED/ua7an9/uTlV8OwqcnjVpdU3Q77P+kqTEbQokabZEiy+WMG6509dNZONpzjdnEOyr1
73Mf9c2KBrEXLbAKKq56c8fC8nhtbSDHc4BX0hk9T2gFtnnkdetOZB8r+7vKZrtUd6hlsIQvGn0p
wA+ss97BnWFpUOihpkJBA+F6Gr5j6oqbAp6F0CRmogKw0+zazeyijryGT4weDU4lzcClKBhwc+xD
rX4NUMpEudnU5g7MGCjSj1TBXSYL0MeRdVTCCfr+1JnXdzQbKwfM+aMk28HOfaY3cdQ4Q7alG568
AhVxREJK5sZdekpOqybp30lVcATM4FwEYHAP7QhEcK8AsqpnPp5qSAGF+GnyfPw/A/Be3GLS3INE
ue5bvc84H1MVSIB1ecN9rdRZhmbspi+wUARy9N5hLbTX+A0bVcAtGL2k7qOlqnH+hyo6RVUms6Po
SgQEN/BcQU79kBZBw0ZBK9WN1eIKf6W3RkVAY35Kh72eiMMRSlVGpRO23tchaOTqw12YB7uQRrnk
PAmIpnHmz0TVYoF3MKueEW0N2dcnF8QwoRHvI5j6Vs6DXdplmmNaW4jZap04yuOje9gG34hub0Kb
3zt+gO1IjEkrT4A0otgP6+ecyfa0+as9Por7h5xkSUiwTk6qgv5/basz8E7UB/WV3t3WL7s5ALvE
aL23v3W7LP5suNumogwhHkw7n7GyHcDbhze4F7xpWzkPnB+5gmMD4AEHctEdjUKmOx5NWSzCvPKW
qqB4rB+N143XjbjsgUXn7bfO9pm6wvJx9SUOTQQTEeoP7TEpzSjUljK5ylSLgtBLZSK5Q29XIJSj
5pDxSp72UN7cOgh7ObYeMSggV2DzFukGsFPBS+L+waHLC8jjvDBBy+thBFaB3Tq9ATfM+mwgUz2x
FWcLMJUaizsokNi5L5nK+13B//k8dSurDzhUFHjcyz81u71aC8KwUYMgHySwl8f6zsY5/JznBebJ
0fRDKEni1QgOXl34OHZZoce6PxtADoRkoBSxLMGM7/jnsTcTWNxzo2UnlyWMJYg0jXEvtq1C/OuK
5Eurkye+yr7v/W3g2DDat/0gTSidfulyuXaEb9T3BbJ1SlbkQ/r45y+vIaGSMtma5cTeCO02WePW
7MW6IgsVl4URz6n7rwyBWRjyORoev2uaU3uCkFqo65MsMbV3g6D9mFTD2vAYnpDXpIEYCl5G4gzi
bcQRH8TYB1Gd96xUyUpZjz78UKc0sEI5mtK4tPoKxl6Ww2R7+jErv7KVSaYsk9nCkICMFQ16t5W3
kdYGKxxZu5h0WmIfzHvbfMQLQu1ixra8MyZ5nPFM9/cm6uUvL61BnSrqMGjMNaTp2Q6lMTU+uisw
zW377PIBMaiejnrMNkV8KKDOFBQbRn7ROQ2xoeP6Yc1U00xsLAjDonePxqrvpuxKMNuL6qHzhQ2U
7XU0N+L3ScRNGVDyEyxKcZtQwl4EiuRdiPge25CJqtcgLaeRigOkx89NwHaW5MitIQ2FY3WJkI8z
4zmBlzB3m2KsLLem+aEBmBCRNejgcM0c1v9Y+pQBGupxNZ7l5UKl9xm928VLM3pczsYFQl1nVwQ7
5rgvhj7L22nTgxVGLFyQEbLodYb1XoqOPEjbz48YXxveVYaUk2kThgLXtMEMvk2A+E24LiwToTkI
M852Ry+M0B5SNyNX588ueETYNmHb6BFWHW29Itj90dsDfsVDqVqxSffjONMBIe1Dfb7mNQBg4SSO
zlOgp2b3zA1+23b/K/0wUutlcBlfmtmT/IJWxfmaadb1aIuzDKpIOYidzka7Gys3lzE1Cq5qZrZ5
6CGwclRNtfUhHKO4QiwX/IEIOsVC0LW9wwAnxu72vXXCFnByU63Wcu9OD0/KgGP6t+KZnRKcPXaj
6CcRwBIqYD2SLmFSCajbzifWyfHmhTERO9DXqKvDwZ3zu5LONaN38C3Oo4JXOe+wHtQZbJ5hmDQu
e4sT71UBiIJI4lpLDfkB3sTW9UmRHl2Q7p6Sxlb79UEGVg9ubM0KsfAtnq9rq3JxNkhUwoHg6LFC
+123zTTpOk6LUvjEJmUoJ2sgn4fQM5H/Y/4CRghyJe0T24hhA1eKzqkgGmyMkBj+c/H6alckxnGO
brp0ZfPf3HKIyfNA/VLcJ2vkOwgue3+3/+CExA18cYnDAwwUpKZHyGmYpvwSfAaJuLhUhp33h1iu
7FrnHsiSfXukgRmi9l85pi3j0j5Wl++5pPICJzNM1SVdmUZoA5UvZQEx6ynEdvhgT68kWQR5/4Y+
1t5WTwR2C6Y66BU/+0aF+EIqrn8kseXhYoEmCPDL5ZZbr0rLfUiQLid106rQraHZylAoYZVUJ7Dj
zh6rKeM+qZsoGLAmfTgUpo/1C7b7Jh0vBemmiPb3qc2lqWw3qI6aX95BKaztFLxunLuf6GPuxjho
9z60lL7uBh4jTK0w0co/yvMKs/PIA/AB92sQ/jcO9PtUMFexSst1pDt4ETY+xSR8rw+9CrU7Ab/k
S31yOnFF5MzZQFDJ3pugP2oMszhLI1oipoBVx+odUNVHDi2h7q+y8+M4SfywtxJWsaDiXJjqSdQF
GlMSbMKnSfpEpdDK06eK9pKp7D3Q2kJXXucSfeW7VGI8po2gphrwaFfhaivwbHxaiPD+zIK+zH6J
SMEvnj5meJEWB4/R6t8rJArvciPLMlEBPwkV9Uqebb3SqQv7619CMQ+xtDMTJQv3KZcgbyZRwgcY
DRRUebyij3pX5qlb8iESncqpgWtdqvt1sxkt11mTFQQlVK3nxS+N4Jqqnrop67ZXdfxhjccWRES5
4/v5JlQK4ZPVM3794e2PXvGCsNnL5G9lhun9dczVcVcqr7E/duPsujJeOclOVceZZ1Ko2kEI2Goe
R9lEkrjrxRokI9y3mZdHS0KR+RZeUK0x1Qhi5Qo+Pk+d0RmgSy+iy/DH7NGdGa9KKRrN/ZbrPqi3
VdNLKVSnaNfQUxuTpHvIQDr0gT3R3TXgnA7E0Y0dtgpXDZM7u0mWecJy+JqbRTqoms7FJgu4a/8Y
dMpin7FYwFYkhIpNt/+HYNmuAClo/zSdE9pcJ6sPLqfOgtOUlnwlo5f84vNYENzVuCTzFI1ALQK9
JhAAHjggrvgIRDii+L5ay+b4E05qQEsZ0SxvGzfoZyzebIv2tIf9mAfGFL1Gnnh8cwAM/szMCoCO
XFgTTeJ45VlHWhlnE4PhzYKnM88pYtyV94JP1R26RLECIO+3uHWgoH/XuVfMjL6Mbuvb3D2pZvpN
qolL9k37/pSRiQ2JjFz3hcZkD819OXxCKu9lenTh9DY2I78LusWVXmIHtVXzXHQjf9PrL5dZbCiJ
YkK4DsfBGa31tFwHDpcmvZzarX+ZlGkBXBSR87TBZEpAICqKEqumSj2IaQVCASiJCh/JGGEFf33O
y1f7HcFXR5rH3QKZaoJKNMLIbkbCrs+PZPow6JvOBSAin6q2Q5vSoqR7fRy/L9Muw5PxUkprCgW6
2qqLe4SJXODNxnbOER73TXtcUVGZz8urfExaVoCamXv+ZBsznN/GQYtZb2F7iPYaEzc2c2os31hW
lmkMMviFDLab9a7KdAqk/xV7hsq4jKrU7AyXrVoB9UHKl0WyH6rIY/fkMLchSdqrAPIAaHAKJNhA
XNsMM7L6uj7s2iPQFKGmI/A60i0U5T+KcqPG54qDowfLfnqOAvMuz/wWM0ijvyLJD4KtNLMIrlai
Hcz5XCCSIucOM7aL1n0rLWUNsPzb4Ucp8pZClUZdFnDLiPqUB9cjr4VhOxtbRzEhJEszaRNlU4M6
qko3j/bwx2CDh8cG4D0UuUxY9E/jKotlm+fWqiMiT3TvHxcaMuFy9HMu0GzOOAC35ypHqTYBFZds
5xMekca/d+3p3yYiC3qcFKT0lmpeoODinV3OilN9Yml+mgT2ocMDHkIxdwuSu9T/yyJ16+bS6OoF
i6EX7Hm1tvKjtBX/azCXDpPP913t8zey+QJsUK3Ex40+Zs3eXhadV2HZr+h7bvZDAWap8dJfg6So
FxZ9CqQeUFmP0c3oSaUqmaSu7iTL/sTFUht4g3SOaAs/9KqQVUovLR4CBBzm6SCkI2Ablg7yWnz2
rVHK6ZPn/4qY44dTWprCmCfr7y+M3HZeJEaasI7IZEcaGc7NajPuZ9ndruj0XvhvUP5JMIt2s67/
opFU0d8MET7uBRTEQ+8Ydit37J9pxxN9TuczeyZCimgmHDetfxN3/OnKdHfncUTND04lN4j78Dke
6moAejaDs4nlnSqUG2I7eM9mzzkUJfcH9oy8h7yWKLYikJxvZ9nGEoDoWzAkB1gzilO3LSETrr0B
bGVJquQHvktYakJwCp+UI+818Y59vf+R2eG8OEaqiXcEeN7DIS7NGztIj28CII1f0/6lIlda7eWm
8i2OxuGS2/GyDnNcXwQge/6+dZT6FQ8k87hZED0J+zId+ptuZ7/d+Q00xL7EaEvyj9Zp3Brqw9ie
iWsofjCnIc6toVZHQX+WjeGhJVPDW9foIhMme52IQycYCdR87iGqrs4qhGk1r4NVVlrhzZ9P6qQW
2fyVMaQZCJRPLJdfGidPJqQvUOAySnYeVaxlx/YoK2KRafCCIb/xNfowxEtPd3qn8FhX1krHwe0y
DQBX5XXK76eLbhILDBiid+n81IE8wgoKYzKX+QUjUsJHP2Z52EHbtkIkRgsYd57Cl5gwzLO44M4J
Y/mxId7jNQPxT00hx4LtkoNfjxxjmM5TdpPkVx6Nnl1DJDT/ijr9eDxxrKSce6fTVFPUeQ39h7AZ
bxbM10WrU3hT7JyGkZebYL2+Vww487iPcsvZ2kryX8KZBoYxof6+M+QMMGwaRYw4P3iXUTv8KKF4
PhBqF4ixvQqZDJis/HqapkGCjfYGu2gXtau05ZUDW2k04X0cilvtW7DRibjdC/pOpLS2joYUXQK2
8dJOcGbPD0lVuyp1cG3cRa0OL22pnDGz+ettcH+z4NChvFeGLzIOra9H6TSaIoEz9OSEGnoP1E+8
j6mEjl9NtwfYgSOb6BYg9WBRk2RZj/p4A8KprXcBx5UoZkH38fJ2UTBvOjNjRADZysbBrd3YKYRG
oVeJaKT7ZQcV7IvhRkQdPF5zi7G95CcLA+9kOHPabduqjHAvzvQIloZGPjUN+hfOa7ZO3pxn+B9S
q7mEhERiNKlMFSbQ9pybR1+2T6+9lukZvgtiaxTyCmXGk8qkQlt9cHqgoJyUor0s0pixY7/65v5E
3s2Sca6LLLUqDTDg9O/cZzwA7LZC76/feEAQoRYpUu+wceCykNFzm44Fp9wZBTcSyvrF5IYSQWSH
dtgIgTfowc4AkkXaqzCjfOggga90ftMqMOn0Zycc9snf99CatYrwtWVCh+X9/RS0fCl83e0m0lQu
1fLdmiv7RimzJ/gyz0Q+Yg1qlHTSOAi3rtFhEYgpwWT/NBRzEPR8AdkbRGall8owc6nGxuoHWAV0
Ial/SiCvPGvGgpJN+Todp//u5PM1uKsze087YNw7ccwGU0d3hXtzv2faNlbg+Qv7Wq8o81UAeuJm
DYZx5G7LcKto0fLQ0OvZJ2J2ErwFEkvtKUFLHpVj/OLyYe/N56i2++MaZPXNKpxSsvagLLykQo9a
qPOJjC2AyfmN+3wofcyfvghTnSjgIuIsQda9jxsoovUwTw+eq1nulg3oDZbZ3R632ZcMGHRwhBsX
vF+Sd2xYCtK01pCmAOv9WTvpY4Qn5ZqhJ+Pw9Cg9eVX+1N87WksFf7NAzXXF7lke4/lUKoziDRkr
L8qRmiHXEeRjhwIIkJ4ojf3mNwW1veeF7WcCFy8xWFmpq4QZuv0DbijhDh5wEUNCcxkqDM0d3DV4
SC0HEmk3ZUpNZdRKjDiy0ei6cDo/jmtXAHoIKLL1L03fn5I40Hx5Vwq5q4Fg3hj672bsxIRgJ1SN
/OBdgTb/A/impj2PdNWdXfb4qmXcB00nKULCKwImtA/GIvhzUgOZkD33s9Qj/624K1z3p3kpyBBO
jUTlFY8Y74WHbUYEFtLn7HlNt+AS2x191WHmjcMQNn26S54szXKQa4Yy53nj+dtUSm4aDH6qX8oa
Ehvwlw3epMT4hTw9JqJ2qfpHJOlxn64RovHsh1WRcEyyYbKOSD2SayrPqVwO4opLwC7PCeOSrmdn
ZBAG9LwJrQPkApPdXB4S3Lg9Cd7cs9Ob007GAvcnncQDNAUTIbsVOhpyji3ewrv6iK3+4LPkX6F+
EBgAL6Jn8T2XJE5UGHlwsTieT4BLujUspasuuUoVIK5zMikgScY2N6/l2k8TUK3bL9w1Af9R/nHP
Y84/JH0NlYxDkLW2tYykzKXrFlPh+TT0rew9kKTJk9Uj3LmFUb8KEJl8xiN3z1hanU/iKzS0w3SS
fdagJBcWNbY8he48Iz90f8yyIJ7SO3YPNUN5P5yaJc3doKfLKHQXEDDNmus0MFrlkqnvnY54TrXH
lr4NzLI0+FFubarnr0Gtaa0+FKib6oThwjPrX9kJIaqQHNdOq21dcTWhHeF9ZNAFGV8l7AGWjxRk
MgdBou3HmhauhKQrnkwN0+7Y1LeRHxkcNT3VZt99vbpDQzGdg8TVZixIv+sIHzRSf5+ijxOYMG6Q
vz4B6rseARsDHPVOdkla97BbWH7O8X/Hnms6+IriedinHseri4zRhvR6myKJsjCCezUIq0vaPp88
BdEp7cCShFZn6u4lPXzBltR1IdnIkoyUl5gxfLV6s8PELt0xCZTfpV7Fe+WiRg5vIj2dVrHlL81+
e5DpBq/cCXPGVV0zIhVXunGxZhgVCfCLwdR+NJvSVYBoRI83ufPj9OqJWYXLy1UdD/dbf6c14bXH
+CgzA7Q+6esE/KIv91iR75tpydq1ZOJoByRTFWb0uYmHNt7AaEFwgJPeo5dFRzLF81GOVJnOh314
fQwoNyS+zCvPMrPbNACkUtucbmMbD1B3mWTrE/AtrwsWQlcQrs3z4tgyVVT11nBTCf+tb8L8EfLW
Uu4Ke5FOlLIoH11HCO+gCLSwRfbkRYE0pesxhs538ApOk2U71vBp7cGGITPGAsHY4ERR/fzWfAtG
hTSvIlUKcw4bz2wf7bPPi+Ohldb0WRblsEoweTbqW81tRsV0sWXnQBJp4g7aF8aDgWbyIcNoqfSJ
QFXpw3Gxz+jEmkHpmt72qKnK5yMtQ2/j+RxI5LSG1tccOHjWDh37izj9J2Z78Gwk1ZFiBssH1kDm
Ipq2vQwQuPPvaq8EQ8ewTXtMisjc4BB7PhVyIiIRQgDYdEHY9yUkk3xVL5nd4oWen5Phl+1raHxq
4V9Obkf0p3r9P1Ju/ft7zjZTP7xTVi9258+qCDeNso+qVXaNTCcp5PGcLLfGk5VITlvZswckoBFO
vHEKMncosRIbPdCseXQMGEjvN6hLptmmilrQNiT2/pzXu6i7YlMmkbLYgj7MLKhRO2FrPo5ho9Ho
fvATCX+klhYDyWAAAbKQm9PoKu5tDjPZlzmYpeDaOFOqSi0AzxXlMvA2h7/erMXXRRF2pbkFWhGY
cmy3Iijg0OTJQ7NcJ3evPaZI5bCkAmuEY4NUbHhKNEJBf7i2b6R6GZ1WbdhMuqmhFFywlLD8df61
UmHOydm/nUj7MgMXpZ7w46rJh2rDfrbZGClfr6Z4vdFefF89UChg+l5UcWE7wqQELHNQ9/yveyXT
W0wNphjY4m7buK9u2pvHZSW6fdm0jYcx2RS3zkprGsLLCsNjscCkoFSvX0fk0d1Z8z5FVIxYee6o
WJL/leQ1YwPCRkLyS5PoZStzoKj8x4trqC1HIuLJ43BgK1nsaouP9rPhuWhlivmfm+koKpnOyQcf
XZkE3fScf0A+6dZK3lNRv2QPey6f4d1gP+tuR8CjciaiIMDr3Jdz18ZZILOQzz8qWgoRyO/niwBw
UvHsvL15WMLGQMiIoIa1N5ZDyH5wCFSkubHQGpCqqSy5CMZ4V+FsoEOq7nNgQJV5YNzM+mmgdZ9A
EW/7f98f1/WwLaBT6NFGOUsf7+xdcBOyIkipw46za5f5q6wK1eul20IvlrqG82HzJnCyZ1JjaL+n
uY2iL+1nccoAs61WTFsqSgQ/AWCw0/HP5V3Nq8NaShkAFrryOpiAqV5guzWVGMsbh9/lUuuz+Dqp
zpprEXwXyYtDuRMVTmPqvHOJmv9t+CQApcHRUmTOc1Wb2NVPh1yl4g1scqrwuPDOKQydog8R+y/q
VR3OiQjTxKHJOe9R8ho5oxZ/+7EIC4gAS44VDu3GCW9TrekW6GqlGeIWIYg7Q7zMJEh9z85eyiHR
usons5XHR3Tc9mU4sLsPp2agW4moAKHSwiJNjuAl6mMUDBJzgV54ZgxrmJtSWzKC1ZcOE/P3dxrX
Wlm7fmuXTyIQ2hclEdA3d0qYPB5lR8hq95iy5r/tbhV4BuzM071ztShrtVX6oTVHVIMdsRZHe8Xc
1M+9OIY0991gT6uLgDUvnOw8ajn3atM/yQ/sZv4XkGwQF6G1HaNO1mGS7j12DlU4yCoDscyyxsPw
wgUgwR67VvNyDGYBab3gb3S7s4h8z14mmFA3wcWnJN+t6e/sviJg21LJt9kSgHvlvAa7f9ND8GXc
zid+nV146KQX3VQn+15nSoS20B7BbRW7/hPtgwFj3H6yBL1E0vGuiSPIWMZDE1hgc/LqElMdcO5V
lquFgJD6+8WOpl5OiYpLcTYFllXAc1oROH/zbHa1+8x2nDEPWXDSSYIECiuFe2YcFnzA8sasHHNK
KuclMKC2mh+P+a+xZhwIQ5q5e0UvKSqhQ0+AOFkN+vXLXzYMVD5TjfVRp3XzMDZcMsO2Kmx+QWrY
Jqj55Sd4/0eUxGQ+bvq+B9Xb5+8StRCf288lObPl6UumW0zdv4amJ9SR7nsow2kbtNJXYGcr5NUA
BeyCFybldF2LZ0l/tPwHR4z80hIq06ncmWZz/m7Dnpm9uppB5AxgBS6x85VFHlxrpidUVfzr0RYU
zVrV2z2bZO9Z9IHiQR3cNMJIx8YYR15d8AhRixTxwEbGXhzVUddKwpvB+Etk8thpml9nuzy3tCvq
JlwneC9VcULCTheSzZTs6aDc31FB6cNiQKKOjFXAiuUeIhFMlsXSVfRjySlxquoquTLd319Y4R6l
lEDEo9FMmbpfJzCjx2wYQpbQYgC4gu0lz490Jxa1TcQ/srFRMCg57AFspLPvmJbti+7JbaLSuSQM
GFookBkraQrnwB+b6ldGyqj8fVyskDUWXD8pfDxZ4FA8VaUZgLM/ySlcslblONuh7tWx8z0fQBj/
Q7RzPW+GRAZ/uWxg4zE9bfW+o5B/TFcEpsAlzuAQzfH/+nFBh4EIYONJrLhh4wLvIPJfxDZEJrAe
Fyqp7Nhw1d4FjNewVtqrZbZf6Z+KNhyGpag71UkDUKcRAYXXR8vNtFHxDkEEYz+8lb9hff7IearE
iwX7AmUaQAKJSCglRLO8CGeJFdUM0VaXaOKe+F+sXm7OzOoieb7odhcmD0G6aAYn5JP3w61pMCJx
SMz+afgmQ2oAkDi3orFAb3V8Cpk+CyFJ8EsPfTCAX473zEO9Yz/5Rn3Ca/XNcWm01AT/VsZ+3T4+
dxc9ey0LOgRLw8xnE4u4sSvIUkgjGjF5tv8+dsYzSv5fzH51pYEx3vZsblKG6fTgeVhP3RQ9yfgq
5ANImTQO6poC8lLeobrHdMLSY4q0WyrdEi8DFHcf3BI0h7bg8DcFpg1ArJ+vocieUgfKkub/UjhK
DI1/unygz5L2Ht7V3P1a4SJH3tLv5gmbs5IMFgTY+8qfTEv4G7FaQoiRsrmKIl0j96ZiEYoS1ltU
d6e9rI/qStq/zLr8mxAoStiPcvbz4iD86r+ExJNO12Lp3C+Zi4lQVORkgx7MufLzlqTvUP1oZFZX
aTd98Ik6iCbhZajzpBh5Omm4TebdSVWytPN8R/079JzWTwEArsCv9FdTZB9v7JqyZZvECYu1c0yf
IXXHSvrSpea9LRDRcK54z3GvvRv5N6ewLOBrGrsr8IfxPKPwPuK9i9O6WLGbBuB3SDfV00Vt2x0E
NNn3ARz5H+SwsS6+7fUXQIedvqg1F09T+zKiw5DhPprQnv+0ufYASEuM+6eWofmqELn3+WH5nRWj
m3/RwP8KrM3VcUm4UZ8GMfiuWnBP44cz97AXMkYvZ2zfQRi23lb1I3RYr5rVQDil1y0jb15O1Yuj
tBEk1pKFS/ykdxReObIgHwSkEa/pdahLd6DQWllsFoEx6+JrU6xXzgf7wOzULkv0lhmqEuk4Jr71
Sy8jTekw7VTeHEkygUnOodVQVzIh16sE67I5q7IN7XgN+e6d5RGpRaLw9tp4r6b/d57yyCG6/7G5
cHzzChJJgyEGOaPVX0WiE8wCKbVxUO22z4ZjlOlvEvi5TUSdnDplym8ovzI8DDpzMdoUera9bec3
z7YP3KlV1+W2ITd5aE6VzwqB5Z6K+hjyRfqoCMXAZTgYKm/Me0c30Rx7fUTY/6G4Mq8hYqhqYDHi
So0EKobpJ+wXh6Px8j4jBjhqK7XysJ6tGc7c9P0Rf3Y0mfEdGPlFoP08fEAeo1ZnO4VRCFObWaBE
bsBYXiqciH7joJnouz0sYRMByI2iPZ+owgkMLMCUans9Cvff1NHSkQp90XKu4pNRO27pt8qAJUKU
TkHx5JaO/f8JULMfgAecTI9nzk3MtEGeds27mO3wET90yaI3WiTxfxrWeuYlCrdxr2xQ5YMx75QK
YJWPFx7BlsjxKFVof8TSrbDklQJGW+/W2jYCH23FjI1jI1HFplxhQYMJGwAySAv8H106aO2WC+uD
BXGiO0coo0ICIyAivtTpnWbHMJ1ddhCd+3bxhwQrFr3N+UagXOWtR3ogPIiel9QTE5oNRvAN1vgo
yPZRt7CcLJdXjYM0FQrqYb9UQKwGBTD40uVYf4rhxl6kaNa/hRSE36VFSmYdPsp+QhHCUde4sJus
sgfT9DY6AF+5GY93s9dt9y4y+y8LBI4Rg7C6EwLozIpgv7LnZvCqbeSqdPlwLsjnfrG5oG/qKO3G
K6KPuecEvMMxa6IY7afDW1d/Z17qFdZKqCrdPXjnns6jLjrgcZ+/3Da6Q8wp7e386PHs5V6XOrEt
hCUHVW5bObIQXXhIfFdn4SKDZvdkBqUaQGgVaG6UQ4iVIh5LoCbWs0pLUXo4n7W5N0TM9Vot5bsE
AEEM3k0n/Xv6EVeepr/5HuQfN8yscmVQoNXpRgfEr4PBGA+fRQUu/YB19Tr4kvwfbFxf2o7K/l6k
UFxYZcKGe6A9FqvX2OwhhTwoSPFIbAr2eCM8iWgjHYhOndOVqYSnueS5+/eTF3Q4sk4+ztUBmUqb
yyzhu+JLUk0BEj4xdjocCEjQzobbU+RwtdiIjvs1KSrGknirLojAlTfG+zLD0XwsxZeahPJp5kdj
SQqY/XFcpN0FPxN6yBQ/gxG9UR2IqBE9BTV0w5hB1OYPIKFIaBW1NtD5eTueW+dyS3fLIU5jyMuL
/m1rx2FIFvwt6NraVn16tjHVVMU5DmRgl6RyH6kxCncmb0PoDI5i5zi5zYRuGFKqTTu/m7Px7z5z
U9MP8FO6U2k55fYMVAiaRHtrT7U+cTDTlg7LpPIOUWXjd2/NdCxlCgR+kjWxvg5CXjyydShDqN/J
lLxgwcPLWz5vecIgOsOnKtVpG+eqVpzOpzfzNLcYWyMcfqlk0H1gl8tuOYo6eLNgu9bwWELafXqY
ef7QbwVdhhoNchwySyDUJVUoRuQ6Qu48Yev/Q7M1lLR0graJ+eS4Bu5TSKNqfAsBmkE1vXMP0/jd
cS6so5l70mWJkVj4FL/DmNekn8aKo4dde6PchzJw03jQ8RPiFWGW0T4TPvbIz+YwSn8qgqyUsi+T
0TGMn/lMLwUXOwm5Zvuvmk630ZO+emoEh6rGht6PGSpwjCsSjuiod1u3Ec/vobBuaABzxhMrT1k2
Bpg0qWmwpc7AWfXYMP2C3toO7GBbDo7ut52Q459XhZjJD7Cdo19pzPToisZ07tVD+huEEGGqXal7
faZt1lPBjssdSMOPSmjei/s8f0UiWX5ewtSmJmlir9mJy9qn99Vmehrgd4HxGuf9MhcewGTJ8v1/
NZH0aDfs8yn/AvCrwqIXWlwmCnwvE53cMmbEnvRLp96sGImRZTFwwAS12BuhtTc4WVDlCz+NxrG+
dwAZ0Ii4PjxufuQT4zqgD6fd22nhQTGfZ/NHnKn5goeuEOFpOtFR7WxpBosU4pkTyMVVKkSFBxx4
u6eM1/n+v0f9dkwoZmS0MZeWsuvMVKT83Kf4t79xF0ILpUzmwKoG4opJHtKAec7+ALxsf5fr8y6S
ZF+ku3Vwe7my4rj6ytadWdk02w6jXed+/LMq1WMAJcK6GG0rJ87i31nfDR9cyWBqdSqMs1y5mXy7
k6Md4buhBlzXpUxgLogwg+lWiKDF7poiSrSZx8KW5pUSfIJ9UJYPMZ5LpZPINAmSioboKP8axKx+
htMvFQ2eh1an0vcsYyEtNOpJhWkyHnbvDZwP5Fo4MEcuGSntxHG8rG3Vqj+6IiUtvm8rPLCVnTVk
C7/UtxfM8x7qpxFpu7dG/oFfsSF8+DLZzibTYjVArC6uJFJgoPWJbefSWeujihs8rYWbKJpviHuL
frqJ7R+2hkrsQXunU5ijSk2n+BhuvrjuEphYX0nF9+cdrPZ35Bve+ZiWNJcbN4BsiVPnZN0sxIvJ
Cs63ovai0CnC3kCqD7wFd1H3iLeRm3LTckNoSmDo6BiEm6lbMi/ulEVPyrrF/QTL5chFUVESX7Ky
8hbbmaX3JoLfAW9yaRy+5bOF89KNsTYWSeF7x9HdG/ZWO74qtZG9J32clIA7XHFwZYPbBcV63jLh
6OJ9GJtadsHePpC4p/Ad57dZ0sEr1GkeAJGB2E4wYNZ3SgurEEUl/nlQFrz6zQwRsueIibuFAj2Q
1lnABrb0XasCh6uMkJ6nqMG22netE0x705MO54n9L3Lov3nR8N1iVQEBVB77ISUWAS1h16ikYMvX
o7dPCd+CTJbQgqPVCNjEC4wv+1Ykqr4c0CcBYq0/ZP0AnztYTxlvDH04qludLVecIhYos0Zb6lP0
fLhJxqNMLMI+SiZxscWDzQV3LtkFgUP4qJynzQJ/IyEPGSTztwHe23EdgCYzVDAepE2xLINpaDuF
pAvT4fYn78O3wVvGNj72ay3Y1m40y8t4MEXPTFDj9SNJcbgZ6YslrqNe425QJPRY2LNZxCZXrtJz
68h+b0qg25sGB1KaBMXSYpbDN5nUTyEITrnVJiELvDDQWlckYR4S2XWOI4GmZoDqeqfOfrmhukoe
OOnZmKUE8lvZVmtKQUikMK7vthyedXyOV8EnP89TKcWae65Z/Q1AwXPfc7j1Hjo3I+ulZT6Pt0Tj
1hPHpPwLDDTTuShq2n5ZBl5JGcbkCc2eEc9PyLcVnurBmPQ1z6fMizZQMzPqr+CJklcLGlksdUit
O930VzWG7a//ZA6E89/vFEGUH5Bdl1yGf6tJfB1T41aClb5FnZPYfqKII9dYSM9WjeoY10M+Q903
bb4ri49r4LvfRXzlN39iNsRDjssvnxmAPJVQuWDWgu2e2zg3ybd+GoO0XoPwIv8rttn/fOByRLFL
pCCYeR27x6MsYEeZc0bVhHnwHaW7Y1CMSwnuSgtyhNxld1tW1TtcTNdVlwAwhxMIebwuFbdGYGus
a7pedSVagded3uwpDmU2u+eF2RoECOsmVeJCS525dII5znCEhggv7CFRfQEWoizNdCp+LBKNG3jO
BNC+UJ2q/g4b2/cH4Bs7AmzQUG5GAYHO39iWD8rmYr58o5SCaTEqcZkFF/2HNuhGCyopIbvlOwG5
f3QVjw4L4O+J7GtFeYZ5EJ5Y2V0IVLjgOdn2hglzOZ2sxTdeOhxxv0JlTooFOPxlPpZCxI1klrRB
j98Gse7gXcODOY1a7PvFCB1u9CgcrXORDcEbAA6WddwZuUPpE1VZ1vdz2rAP+Iygpqe1ngmUD7Pm
e0/R0fRpz7BP53UPgxpHFjVWF5aWMpRXQBWDR31A2ShbPVAoW1jD5gleF5iVQS/aWyrEbyXEXn0D
D3FEr8ioCHfuyn2iX56E8ON4uI/zS104Jf3iSMs4CIZTYWkw0v0n/aZ/vbYWGSdht0Ni09lZisyB
+oxhO+cnkYl6hiDqaovJIitKpjGcznMkHJtXkE/CkPQvcUenpRskvEQ6ipA0/6yg1LLqQmbwIW0I
bCq4MlZJWgcvCcw00RNAGkqFYcB/NtWcnGVVcYI/OnArMQS2suQbUdo2WZSXWWhVDnYovwX/GdgM
rOtWSUzbq7ctXF7Y0OgS1Z3sImAWJXaOQaYsmMSoJDX8DP61eEAubvBuDNjO7F2IVdlEONrFBUoR
R/czOXNHfx2fOdjhu1HEYy/w5BP9Kyso8xTZRlGQ6pDCXmK71kL6+6BFQ+03ke2Pn1hVS3m6yrEG
80ZrYppusTE7C77tsk9sn4hyZXaWjwRV4isTRKBQWXg0FV2DS3uG04ld49dpYKr5pDWYvQLAA+8H
tMEqujHQc8NR5Q2HWUXtFaNc3Fyk8eIapTnRrBFccuBqDLUhgEIdJuhcxCCEdntA1kmKXHIDRg3v
S14DnbDJmjMl/V2rdaNR8BhM3yfMw15aYYwtSnPtQlUoqKArfnCHsJhgMa2WvZDXuB3hsougVPdt
1picSTu/WPEehblQEQL3sD1y5D6/ORFqdHd+cK3j+pt3/wt6rFsf0d76X385fyHGhJG6fWQNhhsL
RIW03hBMfEJrWgnHv/D8JJlY2X9JBtoswIloRld5KhtRUAm8+b51xptgToZZRFv1EDHBp7M2o4mK
0X841la7FlguJcQB8ZGsypsmh8yojrSxs4QKwNRVP8BtZgJQRtTIsW4PZk8OBS7l9WSREvvOaPxA
Uj59FH+W6qMjkRVg5RZW9y7Ahk/02kqz//VqtLtg0o02uZ+JViYtOEEPrgO8fZToPLItbTGIyrHu
XEmIB+KdiCwN/7wlbWgMBX5l2ish7UXnnd6Ej2Y3yLncf07xZhXWMC8A2aGCl6Y4/hpJWOUuW5p+
DIHD3zhBDIkxAoIsheLgEI7GYdddKvlcZqyoS9Wg0wfMK8l+exo93TLEsynVxPo5cwRVmlPKuoot
buB99WGD35VC1xlp/OGIFud9yvD28bRixSPSSicYKASxYkpZMOS5reSiWL9HHOv+kCeDyT+wDMjO
1eaS2GP4LsjIy3RFwY9jI9sW0Bvs21e3lbJbYfJtoqr6Jph/UAwummdpDpuv7pe0kDpzwREhtzyG
ID2YYAtaEvNdUS0UxLea/tykxAexjFWO18HCNec6sjgsD4S4KK7zzvO/ztoZefy3Mna9/mH6WMwK
ZiXmXgvP5N0O472WRio5XgocvHzjdu04mPPncJ8lO8LXhMHymV+PqQToCv/onLmTDwJqHFGmvMN5
S+/Fabj7Kgi87+w0v/O2ITmA0+ZMw7j+qBw4LxG5OlMsyTVYDAxfnXZQ0dGMRE446viQqel6mRXA
XbwnMy0ClNyPHiWfUijj00ZCWT3aFuSZQ6GemQGNngp1OtquF0Mc0Uj+2x398juAgT+NTcfBn9TF
JW7+e3ySYtytCjjyZsCEAokCM8OxWgWnuW7cwhzy8bjhVimWqz9piYDammc2Q1wdSESHm5EMWAmG
jkWJL/PWvr+De+TZyYvQTQDeU81gVUOV4izVi7TOb7ioVIWp6D+yr2EqeYyMsI1mCuf2Y91Ajvg5
dsyf4KxAJ31i6VR+ZbEzxe14LJmx7AyEWyZ3868rU9EeCSNCTeCYdEU1GTym/Pf73rXcsV5JGv5I
MYnmwCnokk+ajLLOH3hG1VRiPI68MLp8Q3MbUMph5jqnpWGIe4L8qH/jxY4KtiK8DLVwxcTRphLj
dr6g4Y/V3kzN3vX4VS4V6iu54+QKSeFrkGCnZ62fMZXhjoAwHQoXGZ30t9wDq4A6yh+gOTAE5cqj
TgIlRc0+a2IBdTGHnFg6FHctGHDJvwm17L/ysUUuY+qyhOo4WgP9iqGWOZDlBp+3SFlZJzMe4gsT
qPwwa2zKAVoaAr+w78NyO6KbmkyJAQyfycd42mITUBynsp44r03kG9adnAOoRN7CwrHNGPmJq4cC
RFkuDw8V228OABmYWAMYrVWp+9r8a9b/XN5TXY9aMJDwyNSdZ5u6ErNR7DEXEaejNRZEqWk2Il9u
o9NfPO+GJyIzHni0M7a/2EUbG7nB6CA7urhXom+n+ub+lMyMIikYqlknJ/avZX354DhW134aje56
WnD1vSQXBRRtdKrAaY4lUIS/Q7JL8gDqVCe1xUK7n5AmmUtYer5mPgW7mcBYR9loj+aLu4HQ5mES
+3wkd8mzyd8iOHYtFLtrbtLKLAyYYdhy4wxwca60TVsuIEzJgzQNygNnBp+2Mr9eggjojBlKtTdL
B9JYsgm1zv8VkYfWJnlQ0aQIglTbv/pizf6m76Y8CnV/Wj6yG6FsFdiUUD/O55ZQDQBhKiEYX78A
Wt0YlreaKWRGeSDC/TblmSigHXxBRdFYE/DktlF3MUfrE0Lfyz7DlsIEc98j5gXdA5/fT0KXfJA4
UbRhwm5Psj7OulzESa2scJBGm/Co/LIInmzal85n8oWVYLXc/6h/QP0yMtkIGkspJiykcwQoYTF0
WgXsCGBMfQOjVeIOVQ6P5f8joEm3LUqN7Duz75UfMUqPXHniIGi568R6TrQk4f1yuKAJQCXr5wtT
hN00WeCptprVrmjGGp0hhPhVIBnykv1h8j6Z94udQhw66utevFqMvQEODMZcJfG1KJxCtFAAQSg/
txJAdZP+eTen7zTV7whd1AfQRe8BZCjsVN1r/zmsqJHwxrljB+xzPZvFZKwTam+zkEpP4ghY58ej
v3ZyeYsKtytEYOo6pLOlB0WDweh5MoBJuzmQoaWarsTx0bd8mPLgT+SgnRwOYZ9/WpCvhE6NkpCM
Z2qNb2bJpnyI8NINH37oVsyu1lb5lw4+0GC3pLfhOMfumOp9q0oPqR10ZD8u2Ju9/6CAdDUtqZKE
PMfuw2hZeJp59RtG/us1uflBorYhIcTTAF3fJQsflxca0/1xkhEDVWElVMTQ4TYCrK16833WM7ms
E6J5nT+qitJi7LDt37P9EmnuP7Yb44INDEDug/NC60YxWXd/2Zb5OawFlOkHwjLqUL3v6EPeoz7m
LgLJhr5CY02HkGscs6EKgHMjL4ZnMJkXlbuQYnBoC60Qxdv4jf0uDWlzQMdCGP4KggHUtBgwOzyh
UNAocgQdYIiCnTTLFaCko2QDYTxsLa+0MBdwrKy7JEFGXac/ABo2x3vIoYd1lcpmpwRM7ch7uWju
B6+xdc+awrcBjUX5KNd1dyiaRXZgoUPwZJ9DYEWuVScLABWU1ri6yk19WJKvgfYio/NKDW3eHT/C
0lbNE8F29eU7PEpNi0+UU21Xdkf/kn1T2EQP1+lR4lG5sY2TPE/D00r9AwCpLGvsMxgdYxOBy7Lm
wMRcVI7g90P7HJQivH3PhICuIvKXG/5vwDgQhgD87uZaXzrBdBaYPJBR5zLq9Sk9AI6OhoPVn5vu
6o//UFAHA0WyWJUH2IXQDCv3lumoHBmIbzlN3w2wGrDWOFPQZQwCrcDKcft3uipEBTUSOLgWTR6S
qsptcL4xNEp6fFsXtoi1LI5Jwe4s5MFPeOH8vllt81TdpdNSjJo3JYkueHU8LYC9xKi9r0L95VEx
3/M7ylhtunSMlmnGHIEwXRieNl0Kbr7OG7cTPnoSf0s3SqY6dcbJxY12VowqzWDcBXFAxHcFJDKY
MfxWTqOLQD+3lnFnZZKXxMiJtNVWddi5DGO2Yf7DzuQtevZrVoSqEKY7rZlBwjDda2ICuCXhgM5a
8xW9BP0jjxpIBFR3WIXMazizJp01yZ4+LqqQVf1RinMbfnOuizNJwGToA18DmkPDawiJW1iXxrNh
msFatkeoBLiF5ym/qBAtSm34HFqvgTFshkiii5eUd9f0FbA7B59tvIa/7YR9LYo+mtMCTdeR3jeG
bpkC3RQLAmFuoE/CwFi/u/hSeS8aloL+ABGIxXug8AheHJFvdSlpd/5pVhD75q91NWn8DOnmMLR1
GI9uClLTJW8lmP5V8X8P7WV7JUfGV7MVODS05mRCk6KUHVF8V5eSc+HV5eyiOoc1meknzZRiQNu4
RYjVFKLKsMrOnePV8yusq7lMCfR/KcelqJNYjBOiXCM6mXas4JMaD65n0jec5VRuaWUA4jHvHK42
aZHfmP9Tlw7ly8aaeo/55tr7a+GZpW8DIkkkpOuRuCkzan9WFXaBHQ/YOFi8HhbF//lZFkLmlKuB
QKeSdgHBtyN2OPMNaye0Qnbizni4AsW3tomwZIhg+mnd1A1hyyciOAHCr6bXSAhw8qZsE5SGcFzq
34RxuRLzaMVtGiWrv1v7ZkPSg7vrlGbpCyttzodWDsX1xly8i/zIFa+f40waHIQvIx8OjHv2to3D
iPzf0+IubP+g7ry7GRfk6XAIC5moivAja14/oHN6aG9kDHNL0Xu25GPhiqLNTc6goNpLb5up3vWl
0mfBQZKf51sTGYWSrfAbwq3DhlmPYgEmIB2q3LMXFzi4ykLLigTqJA5n1kYoTtcoXCqM6h7B66lA
NLB3nAGp3tKhUTWSPBtI02JHG35JjmqPslf9ISERgLFrP1oSOJ88yGEQWdjIeX4EIwEAQDJeUwlb
Qhs95xMkXeNlYUvgd6cXgFYJ9uUs1tE+DhgdBP0tXYZXiJXgG5AXN2D9c/BTJR0etKqnAewDXDJc
q/0orMfBTZFSVaRHV6O8E9DM/Rf6MRfFc7/lWYbcoo64qJ3ENeS8jBmw1n5AEf6AF3vCOSJKDKTV
/GHdFIK5sqqXiZGF0WxOpvpgeUSeCYhOatixDhsP7sjeYzCK5KCqmVBfn6/1iLqgwTc3KwpcHH9y
y+GJMAS0oANZ0PWZaziGLwf+lJEfk59vpvINdeL0qXg039oFgIB/MOTmsOzMDsKSYnKU1OHoH1y1
Y7YFoXIt4lGTkF/JJp+Mkywol7pJ62ftGj3e4hrifGisn9SHygZcoPqM4GlB2JxF4cqpr7gR2Y1f
j3mLM7Yv/sw7K4Gq++/jZ0LHnnwD7HcoXs4WFXg1FCqnmLbx6bXtzKZp7Qk8g8O8vWFUhe15SIsY
yekydZ6Z0r/pKI+s1gQq52Ad8sOQ/AyHWNfcditLYiZExV8WnZZYha0QW8riwslwU7t6wexAw4ax
/YWRxI/FtZLd+7eVrcGPV1FS3MzzicAIIDkC5orQctRFD58xqzmru1i6ctrK+J9PR8Jhm98wp6aW
nJCwt2EaeaxSyTW9mb7LA4/DPJm1wmhdrCV28BTNVumgAU+IWeNMMpn51d/Nh7T71ycLlY6DfKAA
cpiYuexByTQ3bouWrHRGA1s6RzKyJoiKhxSObQKo9Og8ZKFg60OPojSnvrdy6e6sGEbA4N3vP+Lq
5zr9oPmYEu/gB7GRZR6nFHWj7qN0m19STA8UxwRAwQcX+6j3+1ziIA599qY3tkGVvRjBoMbyl4s4
/PIoEfQGLeb9QuLy+s5y6kDinqY+CyK1hI+EeZ7FhaVP/T+MDE1JOl7ceKPhUs/8dxwzJ8etQo8h
+r6nysBEwI8WNWVsvw7ZwbHqwG9IoSsBHAMKzxYMEh5qEnfR4nBVdhJ2KBJjblimkN1KbsnG6zSS
gaLcdzj3J7xvBblmg7OoPPOQqwlo6ktJLR7YevkQHzQLP5P5SBfN/3Nbep/9XPBoxOpxXRemOWJT
1RMRPkf9mQtrvrzzmpQtcvqbDFjl/nskp81ea/fAQrvs3ZGz0dh6SFqlGPEWFMC4HEtOReb3GlY5
arE3ul6fcu/JdEEQswAvQ7t87pk/NQnUT3m00nN1+GqzrDSUuXU4UdgXGHtbrpBHaZIafZCioPWx
pNK++KdEDVy+f5f/7Cf6yTpuDcSAO8DErWGSiJW4qaw6zsWLHq3O8py3Ev8GDkC3fempINh1Q+zm
Jn+yVPIgUuk3fJoaA+fZbJWpyvBqkAvL6hi44TUVpMhwfP/WapYHBe3GJhbJRPvdy3mNhD0Yz1OW
NLDGCZo7Bm4bxZ3uT6Lvwx7NMMC2pcD5h8Djn5K4N4sF/hc8tUJdO/S2IntEFeTBkymKb56IXPUl
+qixsFB1HAjt5iUYCqEIIn7PnTHyFiNJ7i6E2OOnhSU8NLKopOhA59wnD9WcUzhNqHgtDd9Oi0z6
WGuz/TtrLaznXZBPkHddBm5dnflI4nxDr9X+v01nnukjytdF5GO0H6k3bJSHJsk4eV2iSB4xSths
IxPfhyZEZfr7t5uVGeVU2hUfOBo0aa3tux3OeaVrcMPXclytt4EqzzZj4IV92Rs78cQG0GZj4HCn
E+dAod4EqQvIp/dnuPVHcpycwbOpUoa/CwQtxzWHqSPtzwrhl+/ENWnR3OFAIGFf4C1TB/iWFrNs
wwakUNjFbMaGES/6rSKvpybU9n+sHrWWsQwf0xAM6z6MV+qcxmt8BDHj0nWxvoKzlu7ub+97Ky5x
qb1/1AbyvUM60V1NerAIxW61Lf8/BGlXE/cTAMLp8U+NhSzNco4u/0YbezCFSJBK3hOKH6HR91sp
ulWU4uEGR/hyRy0h6ccwKYEEmEMpZqvnYaYRvVksNUkr0/H5T/eaQuGtAk9DwcAbZEBWl45LEE8O
7piEqVq388GarIGyD66I4JPMsFEhGSwsnf0LtNXSQ82YlNtXo7Lz7hUePiLGchfrvcw+MzzdSw27
Z+haVE3jK4aYrgyeY7AlaJklUWKqcYYDn23z4SFaX9cJJ1RxvmUUmZstkGayFUY7wWvoxxjtbRcf
RVDb/6bt8AJgThCUuhsoW2M0iXUdup564Rb0t7LvkdvJkVTK8mGMrsMI3801HyvYoy6u+dsL0Qwg
dkR586dVON4Cj/wDPjmquUgnhMNCugkBpWSuAAY+/lYAUc48EahS88hkBSBc+Ivl780jY762VaVZ
+ncyiaFD4ilJ36s6rnqDZoUmP+AgQnQbJSMzmpwrRP6mX1qprHQTEM7RBgZp0N7sCNAg/ZlQhV6Y
EXqnmIgjCyLy2heSNuIRJ9jOFtM86JfEpqv1MGUmtLZn23hwCNCbo6KZaotjXpl1xI/tLTYvvevk
IW1gJa8xHvqPJsB7qyKIRJQhQ9MT2bGa3qm7ECwSKyEAMTvnHUD9o/u/p4aCHyCmT6aN6XITV7qp
aBxiwRQXRu46gDemATHvci1jYr1rq3J2SzFeB316ewHykjNWbDp0KKDCJ3uVJUyJIWqzuU39WDe4
NOOa2zffrNSjpYJsBHrMdU4iKGipLz2UUU5SzSCl8eD/WYfqx1ATfWEHLeeOCN+Y5vitJh9XMgrw
rJQ1ajicKQ1QhEcHX2h9M3VmZujmkF5nHwC523MMxMGGVh2jc7av5lNVyEfmz0dZsctWdF8QTkxN
hyCkj5FaQlO4lC1sW6HqNF9Etybg98qDLow4TR/gtUQO4LIbKqbaKwwrHbtxRM/f+dTk+nhaq9u+
iN47hKzVhmp/W7WYM4DvPi6VxX32TpE1vf2tucpDSxRUchzSgmaHmgW5Z1IiwqVmXxVSuUqYs04U
FSss9icyPvpm2+3Y1p8NB7XK9IGufRtrSwqEM6oC7+QT3Tu0rXZQKk0E40Eafp4dDMxHuI+oE8If
ud4KzRc7r9ssZjpS2TopXR4DeMHdAWxRNqy3G3aB4OpSXlMbaQchCoFCpfvnxAZivCysc9yUJwXz
HCDKRwyU2Y1U3ZkPCTxIDVNolEmB4wgiDIUvOWXbNd3BJOS2H/NMeevaQZPHsVIju7TI8kkzkkNI
H6QOxrASdQZ1oQAP4Bp4PD8qaDIHN1n/pcGkakhhpIxV2LUkrZjr+SDmii5wfU2yqs4U2yy8jKzD
zQFmpSzq0OWw66L3s0PN6qmjMoqi7kvHboCS3081kwFZmepFFfT/KKJW7ITeVadGbslK34MkbqVC
dqKw7kPjSy0X73GljhozoX2U5vpVTbIDxEj2d2j9sqV1VC7GsXSk6r5lXzGdQvJ5sFLTsSLhw+AJ
TeQ2TP+04a8l5dRrZOyIhNghn1YujU5kN/jnEYjSAiRECAvnMI9zRWyd6f5QwJ7XLCteEjsqu64y
ZtTpXAd2qKRYltPwU40rhCgMjL+r87c4pLqyS0mGxerxxVEsSk8YQ/KQ1DJn3DLeo3dLLFZP+7Eq
gcBrbsDsgXk9wXakVDTsMvM262IGmtdb7p0OF6MtfougyFHyjyQp81bqj8eDfseZMDjUmn6CB6qZ
G5EIdc4RonyPXSBsRWcBqBx4ozzv7lgwWonHxCM4KF7fgfB20o/f8ux8STtQyIFzjYEqJVMT2Zwp
8982FTZ1RFYag630vxCnNLuxt69NQ+trNLBMIiC4s4PCp1wq5Zg/RJ5yH6dZayRx88NZ7R6UHfET
yYnNlyXVNWH6zQ6D/Vik54doROoO2AEfAALMUQOU9qsHSHOEwJzaPyv9nUkjpFXJLlEnS2zuT4pv
MFA/cyYmbKS2pcFpuBLGSymERB8v+Rg4yPlgqN3AO8H86L9g0NZ8TZwOseShEdVptm3WI/ezcmtN
GfOcJ0bOythDiAK388Uk5U8YVGzfHv31dNYCwuTsodHg42n4c962BL18kblHeYqF03vKWwK0UVTL
1/kKYyakfrCsjFCaSvXM1lMA0vCE1JNeHB758xZemtVg5PzTektj888hm3t4DsHyNJr/pubgmOQ/
QjAw5bdtb5dkt27FOkJpE5A9T74CJlbDbl1CyN+rgxBBeUiIPrZgIK32ob5yPBZnUHdUcIcZlhF5
6bDX26y1G2iM10susdFnh99/7iES8/fqDxCWnhzCzwlLAtqPSCNiulQR09IEUemkQX8qb38h2pQ9
egek3qU/5M80tXo7mO1nvCZRuWw86Ke7t1xFor2i/8oJwqtCA9hq41d+tXbFWCwHpR8IAkkfToBW
DsP2w+PEtTKPqV4YyD+zdFKg3G+UqJ4cpjn1q5lt2ifaw4UUGKwsycb0+C1w1EmyYR7rIjO+mqcd
6v+X7HBOGtgvfHcwlVYfyQdGarSrI7pLJr9h1fB3qkUVTwTM+TcJTMOCk1bzybMXf0mIHSaxMhrw
bwrazQxwWUnJU2Mi6YcsIv/Yov+RKxqk6jljWaAy5ZCkmeO8vAo8GXfsF66F6pQ28REANPmBA0f8
Y9dpSVIADvZC3sF4+FL5LM69MGeztN5iBVJ8NCR8xbfvcdSRCvOJjaZxAbuxUo54t4FD2ZyCOxAD
8yKZl+OCDHB3CTsg4MbFXF9mAXq2Vd+XS4hF9gIiFrqnZ7BI18wzbP4L9aRvSjyP8v5+9V75Grc5
7daaE+e/GaM6MFzS2STE8qMtVNv2vKAniHNzpaAM9P/D7i0xqBHIIMuX9wdr3xfbcqb4Bnm+S5Iq
nIVwBlSsLS1NGf7bba4VgH6gigORmwx3W92tvCaP/d2USd1OnmemmjVthuOhS6fc/YjLldKS2qZp
mpyhRxlvWMus5++g5zCtE5k18KR2IruxySpmitow03rzS4XEKUfgZf2EGpmN+VSOi8DsL+eGejRt
ULfrcv2OOs9S52+z88BFBx3UGLlogKhS9vCqyzI/g6sOgPYaKtUH8g6+h9g4LzP0eGaKmv3dRxSr
Rtmpo1mVVUWfZ7HFrBSo44A8gsEuundK6F6am/FWDnuPR3yoNLrbW3cpC2byVQ3yvMhgUVdyLPlM
9lpk7QXyBYyGZNmoqt972Mt+fnGuQzbDbcQdZfQbGFydakROs/QauQHRlwH6vaCps10ZqP3ovwRD
rxB9P+oyxtKIC1AVGYpng+WwiMSQiX8vDYdkGnP2JvxD9sw0sGjwtkUI8ipGVqrzWbbzubX16lJK
rw477u59SIWVHSM+HnMUj7M5W9RlIEJsEheQ+V4LVf+10eUp+8XukEE1T8m+y46usYcZgyDBQO1c
P5u+uJY+V0BeSvxRJI+ejs/iwoD57q01Er8Z7x5u3XBEGqsifKepGc/hRgFessz5PpmU2wQZhCCD
Ft3FVhT5TzI0wekzYXDN35sqgwMOVeMjkjYsEZ+Uj9YZtqhP5pY1KeuxCrwTv2qgTwuLeKcrqItm
uR4F6HSqhCz4dCfnipatQt6aczMh3C18/ioIkQ+jkako7xc5jEBxZblDIkePO1T2kh60im6drpCl
7kBjXvEYreqpT9YZRPBqQn9t2Mjb++KZhUf1S4ung4FZlOUosBFvgHdlwOA43plVulkaHwRaxfNu
E5mn9LpZ/VM1Exo+PV6MSuUX3iC7c/kYwVwYVBGJoNXhXTWsV3O9uSsK9lrsEMEHbrSjRRYn+BCk
1s0XC6qiYT/NbDq9nfvvxdJxcJ7mFkUxh/xi8a9kvcxMw6I/gzd1GIvM/mzXeu2ewRDsoWeBLUfU
0qATTI2MmmGaAKO3WtIyiTFRAVnhXXZP6lcqndoCZv2vTVFqergSuIdi6ks0AdErs7TerRI+tRuG
6ta7l/ZtDbYGk4AzmZNvKC3EEjG5jRQeON6ix7ql/8OZFachKaXt1PSKcPdISUoFkjvLOXg3xbhk
KJJSiFPx6+1nqZXe42kUPAWWPxtmeVG/VC15sdfX6oz6zxak8wFlga4lAHsmAMjXtJZWvoBZVsGH
FOmQnVm2fAivXE6oADyQt/kVgy1W2ADgFUR1HI1TunEwZBxti3tfNLJU66S0te1lT2F7v/zW96NU
F4dDrmWkNrSX9Shc/NkBZZeE1SOLWSb6VhXEBEY6i2GeBBQPjdC6MoM/fgAgRzuBaE+KTtSg8Un+
/mxGPI8IwhHR749CltO60jNbznAAPN8DlZ92MCKvECo8TkGoSkmscvz4HjnwyD+kqyILyMjTS/IY
jcv6VEmAfg3s9BYQFuKLCajYtYolunB/HAdGZXkeMZtJQfFit5w2pLEtTqjQ4HyzBqRMnKS/+pFH
U+9o40TLvsJ1iFZ04UP0tGK0eu26I7fJkwq8Jtvo8RwULnx4t3FY3zsQQLJcBsclDnPCvA8jVvI2
7/7KzHMqYC/7U/pTNj8U2t8DCiyX/mIjaxaC0jTHLDxjUPPsO1skJfGTI0wbvoPqeN2RITnmriQ8
RE+zZy4xN3v0LQ8Sx4lkIlrUfWY2eCuKC0ouqE0bns+elK8BzkVcdhw1vd4OjFc9UL91qngBIl0i
DwGe8cEdojc/HqQUGjVkQhiwv//RxHfIufqLq3IbtfdhKXrKPvCKSl8CgrXSU/rAQoK8ZnFvor0w
wPI8NhHR/8+V6rZLBs3wPBNR5yvvKpr41cdPzHtM0t8CXNAtGgJhRCEWqSa7i5KjolNRMA6j8Vj9
/7Znw3wO8pafoZB/EUHbnzoiWmJnndOtf3oV/AXsXRW9ut2Ops1wOtZfTXdDTmSDtr7/fzvMYh2o
NuVEWv7gCiTS98eVMEqQIi3my0uviIG5Hr7u/prqctjo3dQIX9C0pSbxd5yttvaxwzBTBrJlYHQG
WWL4lc8QvM6JtYijKsHEwiehainK6TE8WblVtw31iX1r2USKikWq4NQwotKFkQnPx9/8W2QW6FSU
LVtbuVT3SlfxviolBkTj5jli45u6ZXMmiZD/LMpyNv7lQW25R1VSjA9tMnDgQ4nfzBsJYUNPxaIY
mNBgZb3EQnDfMNi59lonULBqOex6KXQ978AyilMw1vuhjkv8+0zKqPEpzkZsxJlLdKSWITp7u4Zo
Wvu3+nMg54xVB3oxE+XykSCkCK4Cnz6JV9LV752bijfh9g7x05qTjU39EAa5nD0khGG9/pkSlJ2Q
l3Ll5RwdXlf5rwgb7bPGY9CjmNut2vsOa9L6lL23rJBz8jGpKOrMXVu6eNdQTAVUWneQ0kWuIhen
B1nc06Dk3t/oWQsi+Lt12C61+k9hPv6fMk6T2rC5qWrMO55c44r4s0pX0Xs373lSWG8wbmLNWSry
cuNeqABys44cRr9GEcaUDDJqakQTKjrCp6TYmSn1u6d0ftHblIk5QuJe2F/0va05zkRUqmjUaUlF
xMXL/49JUthjq1vNsUyWKt4MhtAdJrpFPDysYQteFGmwqoL5CMRfZEch4+dqsBlOVs/GtzZAHNSi
xiYPsE13Bn7jSxCM5MF6nULn9lqRoNvgWom99i1iOnW1UwP+n3+nTSlud5YR4l/30S7qVTkXI9XS
pM0w5C4MF7KlQf3uKr7T2iMgtnKYA0WN819YexPzUByngmG95SDcIJ3Q65AfwmrWAOYB9+avJf14
L32TiF4opF7fnIchH5slBSeFV9d4ZLL8qeyTUCWu1SSsZ5tNj/MozttYQmFUgrGXSTdTHz+MwWxG
QdiVMJuQGIQ4bXwF+9r2Dvb7+XMfEB2yJm/MfWEuUCp907MkLIT+Ny/Vp4umBxmwbm1B1vkFR8rO
ZOAUIP8sx7HsV0MuyjKP3ElT0/0E8VpEkpZZWv2xn1HzFsQTAzI7wRhrgISyZ94KZ77XH3srwLLt
s4gmIeQZTJ5oraW/cpYL/n6aExKduLju4nE4DVWCSVYsDdFJmo26N5wHrktpoz4G2l5wqOnHZbog
qV5hcThQ9/ZhMCxFYYQn+Z9ZS7AlBE6c0Ej3La4ARN3ClNkGgAW1ucdLwWo1ByxNXet7+1ojcxao
Zqc4ExDDoiW7P10JGMlEIEs+3Y05kEz7rPMBjFnHhRC4K9f4Zom3/2sRKPZVBKFCw7Vzvc4mM9KJ
vYX8bmLy1/d4ERg8yJLIAKfzXBv10CTAqppdObn/Ky+bFGPu+dCUu9AdYa4YzzjdPp4xNTOVId6a
95B+1CavORxkgjrZ6ig1tGZyjcDW/eYlTdqhk6e5JdgL2UXTclyqWM1PCHosK/6UjgKn0wmRoppI
/hvZb44nwMNMT+hLoT9zgCd4QCmKxwhimicICpgmYER3b4tYjCLN1BhgUIGOItmix0iySfCICqp9
S5x8zzK67g/aBzT/lf0St4j2CjhSi49GVs9KbEQHa+ELplVvA9rL8alQ3QcwxS6tEL95uq6BMkze
gPyqKb4ldJA2xzcAmRa5SUS5sNklUL4VnMS0628ntGCEOAZnBUpzmUqA+FCUHcjS3HdgT4DXl3h0
5q95HooG9FiuAsvYAf8AZCQ5unqanJIkl0/rp3ozbFlmM8+gxqo28g3tYzEZ/4UQ5HTYC/iNpIDU
zqXdrWRMDUiIvGsbJr7UtGrBcxIWlXQjxjzKO8m4tbf4W3lwCJIkv7iUgtBoYjB051ch6TOhroQY
EZ42i0yxmSUKvZEQZbZ4XyASXtWCHI4bDCVvmKwxxyi2NvwU7crBGINF7f8W/IStbveyQIVvT0sd
i7SSfVawHrmYFXGg4CIejH9vV14rBYtev+GX+ivKybHHIgp2+OodDlgy2I4jd7hVEemtQLqEt7aM
bW7KZrYA3znB9/uxOQHNaodoQaXWdj9MyR4AO/Az4ZfKJevKmBls3NrDlJVbE5elN2HXhq2gnB/8
xc68CdOQPJbU3OLaSnKDIjTE8aAgtttH3pLbqp3tHYRVikmo/ktLigRIrbaKqhbgD9Rc2/3OU6tU
ohBagt6eX9Mvy6eRxQY2/EACp0R9VagmuRbGXKqiG9YerP1BnGUuUidccmzn0b36iqKN02eaGSqv
8rDyy7R9h2Xh7n3JQrabO3W9WnfQRa8lmm6/OzCiZ+pJbJMtO1qoBxgGE57fSNiORYmSa+LAvnq9
mMMarrKPEwtCf4mW22N9Tucs75mQOqmD5NGxUNFrYSVa3OFrefOrN+edesIvhZO9NYkFLL704jbG
45zPduXeIUjYPkh7Oi2nJrVtFsk5oixwgD42mrXMTO5/htL3n1mKZzulSfSw825INhWchJ0J67cY
aqDW2w7rC0KFV8qbpP3VkWyz5wCvkOqhCcXll1poHA+I+okcFGueZW6Keeu23L4qSWfiAddEo0gj
7DX+CZhWv3q6izUUvQTvIAjtX5yz+348RGslECdGXj/dHwSeOajUpWxFDPU437nnKEU7ugTj/lKq
p4Dc462ppLO0nnlIAipX++Dk+5NRTYF7zEYHxSBxjMaK1S0XeR1liaqzRX1QnSM140n8IvgtrQ27
uzcLwMvl7NqMKCpZ5YkCfaNeyKmjfq0Y4AfnUwjz2XuyYon3kTPJu5GsqKejeaDKhm72PVCipaQf
Ix+tOYhHFrJe3NsITET6ExF6Ac2IbHLbYfsuifE1+6HrwpqR2Ttm3Mvl/FsYxT3UFePlTBcDDpzF
+pIFmrg0xIFyDx4KweFIf1xCwWTBDVIBX+TY3gN1cXv6x+uMeQbQBJ8H9L/DEPRQafqmXyCPpqzp
TpDCKP1n3jOfROFd2WJ1cjz1fCYIy8f+zeMMvdTZhnRJ7WBeZIJxPo8qYfNfXPUbewuf1yllIJ9R
zAzqNHNMvIcJCbeB2KsPZnlVwgMA93hzTEd3XZUVHwzS6NasWIeTOOyzCkdzhurV1bpequajJ/ZE
30CpgHiZGqAAMkdtmgj1xT22yaWiXiK4Tfc6m7JVxiU0Y3y/bWFv0k4/tSQOXXRm2XgOxtWYAxzS
9UsFJ4bBxyWDP3EEMiPdoCr5S1+17vnNYVpHCTlD0OXWBxYWWDM3mTci1+wlduLoKYr3/QhmTCzx
mBZal1Iwg8Ho1B2Ha9mWUK1pCv6jbouQtmag1SlE4CJurxWmmhSPRxuca1eN4B99ttICM113G7AN
OrTyHl+yD1WPW1kdTUg7MVAmJvdQdbW5Lm6hstUrYJufbvNtyCEMQdzetFtpTUKxMfR3fjuu76FR
Ucbj722VNhb95jx1yWZ/9N9Z+LyRQ1LnRUCOKO6MCVqlB9L3gKs4hcWnfE1DwxqzoNQkiacPEQgK
Pa21DTaMyb05aqqmFZbBhLvLW/B5r/ZWzBlzUZ6yGjPuqmLmEc72TBR+z46ilTpXlHZ41wgY7oZB
61xupgGUp/ECECkibVFScU8yWhP6Zf/BF6YdNiNoxDP+mO6snUztmo1apTqJoIOOmrAgEWneLTYz
glwAqN0TaNFNl+OpzzMr8cZkQ3YQohS9Lnl6vUlz43sNfviBHOXdU1hpXblolad6ckXVULK98EyO
1cUz16BSwrGC9XONo2mTIS1FJQlPMzZnU+eSw868KTLQfAmhnOSmuEIPh4Ff3+kkR18404ogEigT
b8BY8r4CAXCrozB9LqkDzqXEu92nklFTOvwaYZqwC7z9gCNbdPdfWNk3byhsWsc90tEZDSxPPkAP
itdc2DSxF3HGG23nwVdycYlMOcFMunyJWu6+iHi27zh05XbuDuR1C2i12vHWZ2D2NPQmRNU8PSei
1P/b7QY+1pTAmoBpiQofeazyIW3HQ3TuyDT7sniu9R9NYt1cEcCtmmIz2Y4Tkb/ExVweNyJ4xKRD
WEKyaxyNuBsUyKX6PIr6KqFXq9FUC0bqlqj+0o6uHlmdvszMXzXHdlwBhe/LEP4zAqsttcUcuAeL
Jm1UM6DtnKDLMetAACOskBt6y6y3q80koeJSpnT2Tjcv7Cb+veCH3bzlEt50p+6jshDDHZTFNm/n
pyEHpOrnEzo4+oAjpFtHnLpI5ypikoCtCejqqbA2oD+R3Ksi0FiYfotRIn7vSyAGMOkJRg/Bk4m6
Gncsjy00dfgMBSIdRg3dTfhUi38NHIkq+lgY6AyeqH/iUERNRqAcV46mEvzOnvz9CefaLitltAlT
Pvfnzp1ZMQTslr16yOlLsZO5obfF9IzISuw1dE4nT3kE73xjxZasZiz3Ufzw80EgwW3r31EXSmYO
35IRqioLg1+DCak6SqQAK7KPaTnGbOzJZyol8ZW6jta93wKSvYnwVTYki7FDLTWw+5fN98rD2iBK
A5ZnIjFpreB7peLR7I9NVX6e8qCN3YB2XucxW3SdjkhEuu8S/uJN7KfsU332PbzH15z+pezmCgPw
g9r02DWb0tZQMuU0nqSiiTGnaAQTBSxoXIQbi6Yx8L1MMX7o7TwkDb6nKiPxOMHhciFZQuRMbeKy
Dozm3HL6DKaiY1EmyV/CEmaQfFdCBAOj4Rkn+d9cAdQpFd2GRuzzTL/B98CImxy3J+pxrtZxQM7T
GbuTF00VXd+P4uez5KQzAazv34rGG9t3Ga7boPcWN7g13GBejDANhEuJGslaiWl0EEVq6jZD4kFL
ny1WqPMJYTcsSvsp/5ejOPbYQ9wmv27E4lw+7zwwD8lDznDCjlpfLcuU3wR86jg8GqtDo8DSXe1Y
cYUPP/IOsXCADWsjNQU0U7plbCHvRzxa3T1SCHAdx73qrPHzN3FwXKoN8KnIlBGgtZh/d5lLIf/P
VgJJYapZ34CtjLUz/NGI2ohrSKkAh47DgCxUAApuUbPWqhXgNmEGBBZGYYSH2rox/fWtxmDetacD
lEUM36EpgDz7zyIJrYKPe4qjkTTlU6MsXj/wISZgXoitsP3GtaRhPLCXMm9Ns08U/tOH1sSCoFX2
c+bGmIhN1+LR3B2on5WJJ5yWZdgKs/+MTU5j50IMgnmX0dwecTTGUft9/o+IejfgKWjvhowc4Qf+
rsIAWzDyxQVrR/7DueMBXb+YxS3TGChKaC3PqqgcgLD1ttiqAsZxws7jqDEgB1wQMerLBVrhZz4Q
wM0x8LYQj97iJVkYu6h5N0wiQsjG50re1po3Sb6JO4FPLvOTXDdCvyzfamnSR/ZsH84W/5ngc2pd
J/frd0/hVmG/+7VEtdtDHCmEVO+bNJI5TALSlGt31POcEzaXgwFoC4PrBtIbp2I3vp4AYzJm9tMh
F4c+mdfPOmeGZCLXin2hG1pixKxzyg+rtofAQUwqG9ZIUc3jgbR4Ce06yd0Q1OnMmfBWQgJXPdcP
al1+9apw5+I7/5jfcLQDK7fzlTFTu34kCK8O/aRQQdKjXHxJ1nqoyCrHZIqlsMHSiEF18WRLC5+P
oBb36+HzcXgLl4KpsChUvfTQ3SUMMg8xdZvvSNYMZN9rkhNYoe73+MUp1NU0TZ5YFLUBf0DAA1rN
WALLzEeNOclu3z9k71OpexWfhXZn/O0z8FqCQJZFo1ieEsZIZIoke3PQWfVPoZy/cA83rNjUtBBt
cVt5z3YeG4lLGuO1YLCJ0pJI4kjRYddV4H8lKqZjbr/+KIrCzHxpGhYQZuUpBK/Myjk9uQgdW6LC
N72ri+EntlCVlDmfMgae0uDbJJhaK87pUz0RU0m0Uu/MH8ScU9sxnlEEWZvSaqY0obrZp81eO9Eo
orXfGXyuZ6TMTHw0rpiYI93ZvEch/4Gxcv9m+VyPh1Fm6svwiiRWvXu0gVUu8k9W/x/V8gqKpLft
Qkraz3XJrYd5RniqdXahDoDuo8xegz/pmZShTdp497M3uwtqj4e+72NtX2vl60iqWLhgjubKqrBD
TzrMe6r/OgEk8Qap0FnNddXfghdC0X/qJZUKbVPsxsLZsJiQSn54Lbss+MY8ra+MIuAIQcQ9LnkN
nslhxbaU8+Zgl16Yd+mVLPRE/LSUY6dDPTWee4IClbW5uTOHYO1ZU6nLJWTXnO2yBNWC45fQtznc
BHKPREPGY69g4BFESEeUa9OnMZWcX/OMCarEOtXsFWNUtC2bmHwOcw9xD8WXG2ZV0R96xiXmsb1K
FbGiOz7xAOc/LtDGuAjjIuWt4vIHQ8fUIPlz2SSduwT2xKxaBBDXTXWOWr6dmtGrSEZ3WQBE4y7k
Vw/grFPoq3LTMeqXgS7OV5k+6nLN+qsEqhHtit5f93ARCrgoI49EwCre5RE4LaFhQync6nNe+q8B
Vmp1LyhfqSc/6d9khz+HQaM3dnBTS9HFXyLnfuCOSKWvAPcNi5QTFgafi8Iuyt3diufXJk2hfv10
ZTC0R9W+/uZ+tU9JV5UgPKgcKnwA2yMZ49E/t4vw1qCWgHI4fIX1nYOuZeVbGgEqZ25oz+6bfnhJ
3YT71Xwqd/Pt/oPtIeITjJgSiftfOwIK4MB0RRkojORq98DqvivJ412z235x9H0ploBNDMwnm+UW
ukoViFgM6IWuw80TokaOfcF5uk94SH1U3vVV8AKnVmNSj7IPXYEssmhESW7bT8H66Vk4t0CbY8fq
cIA60VlvRAgjuIj18020+3psezZ+gr9ME6ieh4VrtAbc0LOk/CGqRcVuAIlrGL10ivdbKWbHgTTx
6ZUAUYhCjSRTIZq7FvvceW/FhfGgOVuLMPdmq6kqNj/A50Z5jFdlvpUk9AVtN8o8vKfjegoaBiPZ
rIJgS8vZUVVri7+WMODPK9AfOr3aNuCDwZcTeJY69MoD1lQe83KwsqOzI7EM1izbOtGsjU4uznEt
8DfoMx5BnVBW2I+iuUn4d9vEwiZ/maegM+W9fnp/0E2bggQPPEnY5gtejnFfWArfg/u+XTDRwIag
7Uk8/TKWv0RQaSowBt6L/k+2R+UmVep+ffeb2YFVws1Az/HgP5UnJvukpLGqxUF3Xmi4dSRBOlpN
uatUj2ONXkfniB2lwzhpEclKFs5ydP/TE5f4l1VSmyUb2t/Zng+mqqxZ+mt0FVRMrQernd6+Xa62
FU/4kPLLwwoGUVlCaexUJjyNEFVSUVO2HruPoy7gkgIDmSDm6eH4UE+DcWiEEbU7slSvlZrWNJBW
Vgww5M6Cn6+6LeauXzIIteANYjx6ZNqwiixNrg43VKRZK2cLD0yjZnKe1jLVHctYweawFw93s1ZH
9iU/eEyEKAu4gkxwP6g3ZxsEUo/hig79TuwBp0sHvpF2/ju7dtvBXCV7NE4NlFD/ZQXeL3oVkn3r
zCaGXYj8v+2xDPIvuOR0k3x0Iw3ILK7fh8rbUwnviis2gnIoDNjGRhPf4VIFgewqpYlk2n0tHdI8
9cGVpsKmnu9DnYUIr1D3yv/GPNvuDESk7Pka3JIO8NkbF5IOiD0kfroz+h55aPLGolNim3H4n/Vr
24Un6Q7Zu+EUPHWrOFGQTiT650TVIxaXouOkdemHTOmltk8PYPz1HIFIG0NIdSBCaVWmUxQYbRKw
6md2ZBH5hKRXshh1xAtghU7GLye9NbHrogQrgOWVsh9Io2bPKRqQWTn3/uU6QuvXrpnphmJ6l0M0
t7AD69VY/keWFt6AgpMCjB3nvn+g61Q/JGNM5VBuCLuOsr/2qtSysxdQX1xFEJphJqZ4mUCAaQff
OBNHlu2dVKSLs7y2JvLYlDDcl9ovc4dOWejadoynKf8dhqCaAcbk/NpFcN7fldb5FupntkG7DiVq
KuNsZnlqCBwc61JjKvE+TeDS/COVkO91C0+TSc3yF1zvW5F0PM06a4d8MFDjPj7qopa0F2sjy5Oy
4MzISh9UHNoynBWKaQVVj4x65rCRSvlPkTNoH3oKBBj6irjGLesrQhduFMSlXwNgyuIPbJ6QFTjB
wvUy+BHaQ9ls1xOZtx3MDwfk+qRTIeK+mwCkdEdN2NfxCZnFv9jIHU/TRSedY7V/5/1aCpZA8gHr
+1thu0hRsPT4yjVQ9UyYhTy8Ll+nqcUUIylg3CRlQT7P6Q98x+4WjzJd2fvnTdYyI9SMTQJWoys9
HGtJWMsQ4QxwiD2ejkCcjqvfMGJaRR5iuJa+htWOMIYuonCGs3YL5ky3qvVNlpajBL9grbLEbLvc
T+Y5efAQ7GBhVRauySPz8mCmofGc+kaeI5w6mi8dxKsuqSHjT7ISQw94jTd1yvK9AAwdAd/Kn8KU
cwM7VVQRn0HxZqcJZjRp2W5gKNp8Luc9BZn3iAGV1IbpyD9R6BVX8tEcXtjdvXZZCJllfQ4G5PCY
v94mp/fUaYiP/jgCivsWEVdVLGHAQZw7j4Smle83LUQ5FqjJfMe0YS558oKXPmjVAguAdKZGsG7Y
oS5GDnaRcmrhvNJ3zX1s0ESXQi1kT0I5f9Sy+1pqvy/WbRQcixpaUBDEQgOX7zOmtBvZYkyxr5GF
cgZjF4fwLYOI3emv+xCnQmBOY0Fq9v77QPPNoXsco7ZEVWU3aukhgeGg4IGt7mbQtm8PGvKDJwWX
u6u2YOE7sNqELY+BkVztsT5VBVvkgSKiiKIxzKWmSSV118lEkiF82SbH8ULVs8PHGiasORr3HEhF
p6Zn0AYRCCZXHdeozyurtOEzydOTAE3FKi3JsOgORns9gsWO+9n4O0k9nKpz+7/gLIYG5ZXlv2W3
riwmJKlZonG/2NzQAkkFx2CXJUWmPuSkVXjYCd7aCCcZKQWNzUtUZ2U1L/5wYF/+lW/BBBQLtLR6
7FiExkmHqfq23vY1hDJNROfvVDqnvXwBEP/zb+Tao71m6EOBHlEKWUfERDR4aaw8V9m//QwF+Dum
iJ7PtPcxR5EzQ57yszQm/I+Vh3pQrkck8X1XX/fe3i4ir9jwbewXI/xpqNNtlW3+CUyFduuWZV0K
Oh/1vb4KAfksfKi/YD4+W+2/L2YjbmeiZggOA9eiNsXppYNmHyz+EF9lxVCWIFs8PolFOj6+QhPC
7fxI5+vfjOY3V0R78Hafi96wLBft4XWXfiXtbHkLp4vUbxcete2vat6/ZBjMN6I/F5MUTmaJnsnG
f5pjS/001vWpJ9aArDIGbYiXPT53zTFgqkMqLCuAFww7bSdtFxYl/L+H567UqSe9Utj9Kj5/AZLA
3nkZ/m3UusnOxQm6BnZs3+CAiu02ZHpMfVQ7E8WTAY+zOoAPThGbfy95JOJqC6e40hwtZRplQhnG
0uXXyP450OmtQHCOkAwowVq8pXX61azU/KgES3b9K+u3Dmm0F6IFY3AE2swq6e6snuCy8mTzH+DS
rXW0yVUOLGfJw1ESFyHSf6uv8zFx+L66VNAdrQ0njurzTUX16/v18mU0ov1UeSHkHq0zVBdPuH2Y
HHEoAChPu2GH3rN//tJTEEtpXr1CC933eFwzapVKSiyNfgKdbeGz9xPxKr/8Pu/wyG9+K94GXaT4
tjUae+ns1v/MOL7N69CuzBD1VzH4IpdYgYimUmFSAz7gU3biZoJGcs7EaigiIo/ABjiSlqJaPFz4
4kOpjcHgx8D7f5rGMeth0UlJv6NJd+ipSj1MQDIEbWMa5Z9Fnc6KEdGbYImmeM9KFw319VUCOknm
x1y7L68U1V6QOXaHZEoZrh3FJhBUY7JyOOUlqzhx8Z94Vx/Um7PSHxofsRG6Zyhh1aVvzURDxK9k
2ni/r9YopTESzFUBrRI9MhZHYyoD3mrFlfPAkXeSAhiVpCuGXchw7RagDWqG2qTJv8eEZAw9/mCM
1HbiqE4XB/XyTGARPLYfaLzXdqSVi+dmD/RhLrJbUYjdyG28NxoYp7S0kbQo55yDVyT608EN7TEG
Rf2DRdJCs0iJjo+vCKCMEVROFMBhTYnfY3H6yrHE4yueo253wmUYNa78F8AqeVfmcG7Zk5anQsN+
YVyzCWzSYA0hXCLjXiWCd4y1SRT/kDsESTj5LH9nzm162WKV+J1/Y0B9QikyPnynrf3EnhNufj8J
lLG2RoMmwe2OcY4M7a4HLaBwoFBGnBJskLjPmTY1zFJnLZwMqdU8I/u5ChgwTNtM3+dRbXYcppCt
yvbw1TTMo+1hi6IuUSJdQdv69XhK/SHBxJ8gn7kuAgJLimWKExI/U7xhWC9pM94ptoVMdbt8u/G/
tV8bTGMqhWBx/6sjZKhbqKKpiA2DMNebr83QSiddtvzRxr7COUNO6nDcmiJWCng76oGDPj+Uht0A
EXQFEOVfOH0lBn2VvragMBVHAtq4AvfY18G5svk9YjWyUXdoCizf9pX29wNa7mchzpSEviebBU6o
8EleEY9ELk9uBTolEZm0kXUZIhxRf7PyMT93ME/Y2DkiomVcOfNtjemvEgpV8cSvd6bQWJchzmy/
FhziyWxJUzSHWP+1sgs8wN//e5qQ2YWIHtR1nb0mZDkNaDB4lofquALukz6zuFipQEmFR+sYqUZh
ocDHneI41gXyv8mGpEwdMzBXRuTUlJO17hicdLmWjtWn01kuBgsu8M81p4IWZ/wgNqhIhod+Lu0A
TNMwYvaIUEbI621GgbhL/0F/iet5oEBWvW6uyr/9Z59Bl9uJRmgmGpce9eJ1cVZqDNdEKJmhl7MM
N7Gu88mVkGW+ZiM659QgOYDRzG13PcFG8k7wYmZY5prbi8zmMKNS5nhy8JqDmW48op/8gT4L6JCn
sWadqNII5wP1ufX9ahQiClaCLF5DR1L3IUlOQWiQqr/hI/drhjCKYoKYcFSTmZsgE7EiLtoVlFqJ
TYpjZ9rF8KpTPQEficPzROE4u6aoJtUY0g7zh8jHPW5TKVuZsAYV/cjsyi1uf7n4OTyMgkEmTDPn
A8pC7HJThdc4uwx2M0fRyxEEukmEm511HvvDtaPnI2xjiJB06DPF0oU0jS6zzqjHFkYoVUT9oY+D
3QZUENjaJbm2tYbZWBDYevFOWkNDCvzvkeWZuHENd+NoWmZNJN+mluy0dtcqQuj3g+OKabMZbOTs
hF/Tj914mZQUU/dxWHLNogh1AkU1s7yYRXuA4ZoQn+35/dSPXmAqVQSz2ixSHWD0xazeG4p3/fp/
o4HmPzirNVql/G3I1XtINv67epbn+bw01GXk9DkStTKApA5Cg4QSw1t9u/S/mcNT1PKW/FE5M1eh
FdyWurlYvJ/pRrwKHopHhwRfWu9C0pRFsAVkaPUGh+ZGkK8hptZ90TUoR1Ret0NKvJRA04BECk1c
JK/vZpZ59WlbWi44N/0LNXcEuLbdr3pQMMgeYwtebQXsd8ZSRrtseKMB3R8noeGtQUaQy7fr5Xzm
scnqbIb39cSLrUDVlOaNqE0jRTu8xCAbbcVCVHUij4FjR6FjJpv7LLgBZs/hEiYK0H2l0iIIGClj
0/czCijSTm4LDsBMPfvAvreOUP0DM1UT6J1T9WG1hPp7Tt2loktNvlDMcNhM1YpERRM9LEnBy2c0
jwjayyxW6uW48U9JDvLn/qTz+nak8ktxaCOOocTrQaxpr5tzj8netPyPXjHr73Ikyk/WXNbcf7PH
DSerhKPfYSNl1+mVG7Ji6mAl+2Al2CXbRQvYIMwuley/aB+Y3L7UIgmPsa8SA2cHR0PGV8ITpfQZ
VDHotJ2mk6JKMiKjryO9EtynnoOxem9PQBG66LFZIVWscez7qj4EZGUhX8Lfdqm66xSoR9DT2j/V
bkuTGk7svf1kYkVNZMnN4tzdPB75kl41EV00+JF2zrYE76aLUMZEFFmwt4AXd1MXE6XvpFu69Srk
beOK/UN3xb47zTRa8FqYT839me1n+eiDEZEVXnqNmD3C1yB3eAAw6p/eha+lOhElOq6v7p75Lic4
KZrJm/r4nDFT9q82TMbCrHTZ6S9+cdBnukgcZtxTfEgxCvREfvAD0JzkMOYz2DFprnJAqlzH81Hh
2uEk3J4M13Z6xxDlPEuLJ2Ox1izqQRJFZjuYqAYpEMVpKJokcI0gVR95TplarUm2Ne/Dd1kBg4Ya
1NhdukkvLq3fh9k6aTG56wAFZTX937chS7wuqRBBIqg1u9wqtO7u/M6Uj3UlglXzi6QYe9IUA77p
fkrsKslwLY3Dc82RRDA4ijc9+s8Nbp4CPjqfVcWVruH2KgOOTu46x1l3DBWTKp3NDfDVYl29JI0Z
tkwT/QfcrLrgB1cgOwh+rkVdfxtHZyZAhNzepf8Z+Pk0B3QatACZdtGLV4/noqGSOWa6guQNuigI
KbV5bFsLwYhrf/HfLPwhOb4rPnxWy9Svi+iQRkFAXLGJ31u+VlzTUi9cKId2fMPvip73G2/puRHu
hwn19Vkbpg8z9uHAEv5vpkCdaEObfZgZ5OiK+pGFSFMVfwk2kx4LqEtU6xUvFNx6KmacY3ALI7BI
t6t8mFNDgUk7icK6i/NrcTw7GEyECqHee2XWszDRkePri0fc2Z21WHjeIliy4Ute5VeGYP22B73e
7NVwW0hn0e/ARF+OYcVIsSnZmutJov9Xta8bPpseqFuhvUicTdRVYImt3G4rMMopdN6XSfM2Bd/b
oIgsLe+RKuetzyKeCraHZZImXSDr0aYJWg7QXNWQjoi6x+LmqaZgaFdCT5CDFAc47PVPyD/ATXxk
80nKr6FhPgSVUstKvT524px4vFHH3VYgmLx+W13T6YrDnxdtiTVfN8QHQtxrHVp+jFKw3E2xGBOq
+qCFtGZHCzwPH++hcunMo17CDATJdYGy0FpP9Nn1Doc5x97GYNLdsavn9ebIMAW+amm9ILYINZFo
qmiUw5/PbOZyZQtZT3aEeEkfSIwWMT29wvhsOOOFt1YynoIR6aSxy4YCRtD2QkRtXJH95W0vjrJK
cDPKgunXHmQhHTsV3Zl55iBSunujiHiSUKARJUnHkg64mxlvWtbMUjdSk3op0U3UmSZc4oiywgV6
XlZ1YKJ/rbcNcm+ytIeUSH3zz5xrrDA2zI1Odb62BCKDoH0CwDeoPQyMMdILPeVCtlfNM6fD/vUW
pVJGSzNFdH7vwqcJRtLUFEHQrvYvOCw+Tt2rDMpGI7WJ2Pn70ngayMVOHgOEihZw3FHC1vYDrorF
EuSjTBdpKYuFi65S5wWb21xnvg4HEH1pErL+RdU8JlgLMUoyrTSpwi+aR3ONS+sbQ2df1pm5xY34
bMyMU7ZmBkV9+OE98bd1UJwwnLCZFX1uCR0b95VOCLSI5D8e+XobmSEWEICS5/tZwvDEosqVn7O0
an4bWC/vrWvD9+Lq5KvUiDOSytm9kDCP/rRvphiRO2Psxv9xjLXMr0m3Tt38EVfFznTFUGBbiGhd
obTHcH8GPOcbD8H6mIMA4bpSDHi+WsuQUUdkqltu4mAxF16IF9dK92RbBsN/uNMtUpA0+DRQb6AV
CvtiYVOyvWUTGb59A/di9Voa6BMVe13YmgK2Tdj201v2Ie5zq6rZkev9GHVrqY5m5kVMpYh4+MzB
Q5KsKEEbFGz66X7V23b5Cbux39wKPTJ+U5jwuUO4xOiZ9U5KAzv7Eak1U9OJhL7quQ5mDC3Lvalj
fHfOIxQgkJ3eUhLrFqYLg3/uHJi6vekwT6V8uKrsA/bXkE/Is6T/FRRqx28kBTavscBVR4tYta8/
VzwbueKBWGaG7yKBJ318zmD/SnDMlal1V8U5yW0za5it4ca3gKokOK9CoBCpjwe0vJtdMYvo/587
7V6twOQwRiRhNKYa43+joJWo5NmQN/pxY3kBWv46cq0OmftPPS2CaCEK1TG3Ar+/WKO2NCQiTHB3
dNRX694C+qhZOcqF6rNbzVQgUTMh8UsIzR0YEAUZUZY60B0h18E788KGZFgJLRWaV+Ckqp1iDJnh
/U4j3/ntCPAXJ7NIQH0RSZS3hc6H8x+XbXl7u7IItD6BGP38wxlBnDHsSGwAwsku8i2TCZl6G6p4
/rkA1F70ATEB7DpthPlwuoVebU28mjwwgt0bAmYNdn6j2TQH6nYDrY835SMsb1+6yN+oCVQ9fS/5
+cbFQ1yDWVd3Z8bOZBCPJfwa9CG3R5+vhwwQtstwtkmPxwxAgXJpSIAbOfhCmc3mS5iR5wAfWbwe
zM9FJblgh3HHoCSfO8gtoJszhzZmHcH1twYteNd3niKudNzDc4z6/XsLNNFDT0RO+UDBvuusKyel
2PDm7ieoA64Ztl2ygVfle91z0KWOTRhu0JxzhogXv1hV1fIL48c9z3Gf4BVslQ3Ts4AR9/Mtvhh6
sXsP/mv734tc+fnrFsmzlhxIOFjeO9kp0wbVBEQIjK4QVIx/5epiVDCi0w9x4BmvX4Jda4OMw3ty
NAwWwQEgRUKxqjSnUS0rfT4/jleo/MnOWpX0G5OL9TsnXqtA7QGf2WTr7J0tRl6KlBgcPCs+k7al
7m1+rj8BxBt2FaIbeWhW4qD2eKE06pU1YB+CKHhU0EXtonoHsZ5s2mI/cg+ypNeG3gsUh+lMnwIx
EwwFKpa4drlSr6heXFdPFSaCu4gdX9asc+tIxBHYWXuuUHU3FLWXRyPCF8JTVyAeymDmeAVRyx5+
EOLyKNpqjFPeGTOfVxh0H+LfdEYDCsM3/OpbGEgD1XeS1gHtrXCWn689aJ7A1ngqRq/T6xIJUcYQ
TeSbC2elQVscj2AAS9U+CxjrBBCO3bQ+bjGnaC8fr0pzdFYbreVTPIBe/V3vODni40cf48Fn+XER
kdc7miTrH+GTXNvsH3WlOdNXAUDuZZa/+McrihiuAPB3jjA+R5W+oOT6Jw1Wwkvql81Ox2fcPwxe
pw8ZoQNjs2rLmT5wprPV7xp6tU2vIT1kU9ZAxIX5QhnAgMlHrqYNIN4EH/TChKzMWb9H/8zGeIrJ
J2mwh4hW2wJQwwjJwX28QluIOB7K/V+JaYgfwP7SL27HD6+EvK+fgCOjQerwfNXzGYQ+GJh3jaKd
aiGR3aEq94XFYYxupqOUtfdQuReZJDOE8Rcf69o/9xxelHag5O4m774pEkPfxI69Xo2+N6uNinPP
GcNChqy1bAIVCzhFxMqLxOhzajAzPLBpGfvT5B9SBR2BMMXEaLaaFNUa3F5MSWnNvcOmUfC+YYfM
nAXYscdEu+MmKgp9cSGrxBP+iXzbVmfc8adXMbdTUK5n1Kow5HHOVulF37XNKxE2Pc76yZwyMYvA
Z75dKwRProuvr1L6y2AW4/mwWlqK6+pd+vvL8sFr50/5n5Zp1IAmpAzRTf13XxtRCMq96JoQGg6L
fIl3BzZez6aAnNJ0U1GoMBzlbSlSUzVgUbJxjNkWNAn9HAdFl/RxkXgDqx89qQ3BtvWNZ07XbkaW
M76f0F1zeHFLy6IZJdXtSmTBXpvgUiY9jeQK6BCbpef1qX9yjE0e8UF9ys3tyUMSA27AH+w2tiQE
w8/nUf4r/X9J9aHEhcFSaaMjfEZwdnEjqEnETxTLqwfGY0a0Qi7Ibzp0OGBqWUfIHYoKkLLNfJ8l
bX5zl/U9VJKqU5tiDbpofGaRa2H8TKeBWWUqXE3AFesKXeMOa5b/XVpkdpWBFusDwBTtyn+4/DgA
qK5ZGHUlJiNn4ZgEA2sbU7aDt8H6Sgv1sZCDhEv0Oq+85nwDTWbh3te8LJLa0WYBHuS8o8gtIBVB
3dCzWQkR3lk05prhDBuOLWmgqTxZbXszxw+NctoDVSfzDwyD3idUaerOof12xjyZgNzqvZ8tE2jJ
9crFQbFsiR3oM9qDpuSCnkAKRF19D8mUr5ZiVXyv31YOuLY/wGx5lCKZ7TGP8v/rnk9bo4TBkAkD
EwS8Eb/nQnkySbVO1Ns+P2P6nXPR7LuU2ao/M3qKiL1o4Kms764A4ASnFJP4Qy0auMrBmd9jgJpl
YDBwhLzQpb+2NKpz0pVkjCT7wFHepQVtpSfD0UuKluUn8cij7VIdcczlnd7yRCSYKWLw07jjgNZb
4ZxldLyxxi75FRWKVMmeKcIB7ZAcSE943wfiCrsZYUNQPE+gbTbhk97ynVtcN8DpthC1kvKI+TmD
wne3ifGGVLL4mPRYphV56lUVCtXwJgEN67SGzcuwc/Ap/2FWOeJhp206Wnvc12TH9on6lczYJQNN
4Oj1V5H6QpLBptQC+9Ct+yPw5wKumUII81r4AxiD8YlIr8yleKAp7K10JVQK5AjaPgP38Xt9WLBt
QVjrIX76RUD8lRIgACcPCisXLeAMFT+kb6w/0+yhbhs8uiylFmMrp/zLcFPlH/kZOKtP2cbwgPtb
oUvc34e3luRYVEjyPcm8C8kBY0C+0tuyFrQa3DKl1/WqzvyHxNEoQDl2BQOPekeinxI8XaJYE0t4
2PqfstbpND7eD5s6xafZeQeOUx4eGk96Ihk6fRWa5bIAQ4J+2rRHBSPkflrAzKbcH9u0egWW6MoD
O9CCUtJwmaYz4De9cxPio/Bndhoy7n3VX/QkwS4Qlb3Wohr0nYRzaM4yPfK9XQpcC63MdL/K3HmL
g5Qjf1pvSR6spuwaO/pXnQ+FlR7xSM2fDVqGPBJE0BhLG5TIfhR9BOAf1z8PuFluQrwRRYJkwbZF
YBujl++nKzHCCos8H5T1w/X5hlfJjKx9qApf9mC5lnmjSBH6tM13Fc1lCOhoZc8P0kHoXMYQJnj3
p05TL6IidSkvP9hRyhLojveN+Re2xWluS/HdX/vyT7FxMby2Fj/Ygr/JBklmmcYbgLXURPAgxDEq
YQ6FSCqUCtjmqrwgjkmISKBgz50pHXUA4Ys7y6icskatBxGR8Go68dYNJCLZDT7OpBwp5bh64NeF
EcQnzGjb8PDtWNdfQO+Dr1nhZWlgpyNaqPG4fkvdqe54ZGhhjEdrIvvDDXLHjITJLWD3hbTw6Zrd
cttvALjY+My/+eMCeM1K1+BfU+I3X9KPwBjCV1wDkjr5ob0r357owh8kCQBs39iA9MJFCBK8mP1X
1fqzbBT2xsS0ZoQZEUTcLSB1JwdLuQcDkvxY8N+fP8hsSRDPcyxcr7S8C84N3ud9+p9y+aP+Mhxx
vbtw9hKdtLMHuiRVNrPK1N2Mq8eLIKU6tmgFfnWDBQ330uyyvqFIuDKASyv1iMZhwOVQbIRXwRfu
mmR/lLaF93wAsPmShSK9eShZjS8C60V3en+C3sXD6/Uqu5lJzHexjLPTBleH1A+JMW9B4le+2aKW
QPeLmw4iBYFC2NtNB6LO+oux1OE7LxWzirN0g0/tIWHMjDCzxoeqYCqOWqvl4nrDZjKZ2XPwhAJj
+/A2toumZ/gzR9rp+gTD6lRJFax82A+nJ/GF37Xe6WzVAu1nVslV+i9eZhjkKMJ4LMgRajLCOaxh
4exY424Nx3vYkQ/Lz4BkXH7hNOM1V1qkNsylfEGIQINi2Ypj9/N2sztXb2cEj01Miz0AWdkeFZ2A
JagVHK4i+y3r90Ewff4nB8p/gi35jzzLYscqJMOJ/N8h7bM3DEyInZ4F/7tL+p818WSzr0q7msGR
X6Q4n1FwFbDNAudBiwtjp7pLMzhku+dncnw6DC7Yky9NSthgoGEycJrXSgsfBSjWC0rouY6fxIqV
uHcNs5OrNqUtv2Jge1xW0jUFfeopwHCFHV3+YilKsawyOh6i99Cx+dr2wQ2sTNwiYh2jQVKyAZke
mkzw+QqYIyQtJGpUbniH3GmCLXU6jziHDqwVdzKi2P2Un3liBXnlfrQTEJnb4mFboQjALh9AVJlu
LxohoChxpGwsrufLuE1gS47RjAVoyUJBjchI1e/hWoohhgfsJSl4LzoLDqftlZhfOwybW9Mvd/GN
WKH/83/r4j2IZSYD2uBcJDWHNIYaFfZKFti8UgcD8jZ18GaVbeQh3MMNUtEQCrZ2InjZVpVpNObM
l8g3v8mf2ICabUaLMnr1ut+oKWN4tpgrooh+dP+DOm0A/VPjGNYkktNKdqbo3csWWjCOxhhZa2Uc
Ngo/b1bb54v2OU38nXBQJUQmkFE8r80jIBGSZ0LqyicOmSUepofqTIHxU5Enme/sJmHTxZUpTnFh
WIJwunMQtrSgghjwhjSAdRp6B9wCbtVLDJ08zu+oso62pRMciszjNEnSyhp7jA9mcuYH1W05sUrr
tLaFZBnqyoOmPEp6bh504MJH/g3WqyWMgfzCelgqOH0fxUa36wA7WJbSh/pLBfdBgmeV3cZ7YeFO
invDR2LtYVaCh1RsiuD2HZ07lYx0vRD5WoFmIBm4cyFqj+g7vhZInFD11jDgMwnn4bU6xB9M/nuI
+As+tpIIXcO3krjQp/btHDhvI1r6YnTNBOV2xs/zEfa4XFu7AnV/iY10LbVl8nBySF3VrLrIYi3n
yMccb1mhbtX1FHFmqIywLobb8hxD75RCNJZKQuzK/HQCNOXSnyLv2Er6zvvBkv4LRzGeZdRnDdWp
VhcAiq6FVhxHIw1TJ2iIN741o2JaPNo6M3D2zy370fQpSkUV48uS0Ani/DvAD4qo9UJE5nDjApdv
Cy4pIe2YGjrwkrSxgNaDENS3OiWXxnZVGYqjHGCjBwXpiXRuX5x0Nk+WsDfmbNXaAUjPcPYzNxc3
3frFZ1xdgcgslPkdtywxufaSympxMLJlNGl4tt99R3SozWQucKpV8fM/rvxDht8CxyQrCI2/9ALb
Q/avSDw1HYqKmmHGFLGFHQKyplWgHgmHfeDU239JYVx82Vp/OFmdpbn+yn6EgKzOnmM0J6IEfSri
YawLiiwzxCoMx5oGXuMaXUqOuMQ/QvgbffL8aaxqRcALD967XmPrfskyPjnPfZ+6/Q2uewjcy5nl
1D5Q6zndcAZL1SgsDBl8nj/fRKZP9fSnGi+5259aWJUOihtoPPDWXFbNyXC3Gq4IAzMBcpAN6d/x
XZvoTb4Qs8I/LP+o5CRt5NydwGDRP7qU85cXF0UyS7PWlc5yfv2FEpWLlOsMsU15CEvLB29jyj/J
m51htjPimPAhnoUhPdLjCaTDDgfI6BT0nYYRIsnD5OMiWrmBlDIAEiBFPXRjxxI3+qGCG3lajR27
3bzA9QrBhDbq37IoKHoZB3OWkHZRqIkP2aSruJIzpQZ1znMZ0n0Lp5+Dv8L0CpI17N4nO23AVXVw
Vze+U2LLw79/Tc9x9eEToQRVAWfW+OmbfDbz9PrgOUX3VB3dcF0CTlybhinLQ2gSIepilFbkq63Y
YotJP8qMQcbWmNJOb/B1YSIuyy+93hV3hNyPJpNVNnUMrbUWzTy+Ii7JefCy8UM/AEKKNdiWAzzn
VyWFB2tm56OwDQRvp7PjZTnubQtp4hCGMtMsToWRKVbXALsRH4cwZC/uG5As8pAHo3+0CROuc/c7
TIznfje8RWqrHQCGKjsUEoY4BO5mh1/mGbuPeBkoLwduVnYq0ZeYdHA7xRK9GqCgVyRmTO5T9h6w
fFwipKJmKrD4afDzpj8jlBWJ0RthPZjvImntUNqTdrJK9+nATh51vcHaEHMDrO3QcYnu40bHey8V
tXdwKyan9nwj6g+PQpMI81qWlSjLTUv808oNmENvg53HO5r6NjeK+52bDEN3yRskZvMK4DMRuigf
EnyAy1XAnyixOLmMqZZEmqRwFntWht7oviFeF+f1vVbPh4pbY2Z5uZ3Yqa134+rD2D8Q8R1qQPky
5ZsWcf/AoMIg/HwiOTffnPkXJfVp1LrGe83d/9y4auewzEDJcD+DlnOH6B6I3J3JLferzXAzq8ef
Vh6ElBQn+qDzdKonHT2rIH7VZ6RQCW9Rfk1whArSkj5sjxFJtCkNayxMPSsrkixbQT/uguwzfOMP
goDKtiqGILby+2DLH0SEjxrkS4lAboL5SjYMx2WgQ7tm2k57pE66vbG5SCcY78Htzmke8eQTx+68
IG7emhg/+PomuHA6XPFxM+OXubV3h3x8ncCRpdlfUSU06yPl1nfxHNtIbXhmDNdx0r9mZnQSG5rk
878/KrWjF1nvlE98WV3jhimJXaHPwNo15FXsVb4JkKZicsT/fbLMDKEU3/JqoH65ZOuphxZiKq/N
3+fuPM+oR8Ld86FazxcyUJpZdoRNulBkgrXFtJWXJAjR7GttClKnTKajPMp3AfsBOXsgxDFrUCO+
+pojArTBkKchnQyz8lRuXeLqH4LJ4fYVjczYPJeJePX7uuUIeNQhHcqxt6ctr5U2eSKdZ1B21Qcz
B7WTYu764Xs3DCH3oetRbugQvxxHCI1C3FUwyK/zn5/JWgbyqLJ6BJ3nLyGyJKUhS40gPT7KSa/m
qJwl3IKPhkRME0rDOcBMrcDDMSNzYqnNEJIdTjSMkEWXAXOyvFvSCHCBAd0cYgAvB1NnjmZy438n
WTq6N+i62FQKoJa+XXpAHcW6As/9GFfePzjXgUz85xhP6vWj5wJuGj5ZQLAAoqzSRs2rIByWGwj3
F11kHubZWMjIF2TdBCfgjPfA8yXqgKyJ/5COye7lMEXVAA5JtYVfbaRnZ7J7DEm1s8znscKRwkdu
tnrx9slYfNF88MNAIHt+KSasjzp8PoqUYY12WyWXblh0XKvnVsR1yo4dadRGyaSdyrJyxQqOCRHL
CcSfHjm4zL/9tZVqSInzKGpI5nlbWvpOllyyU8zHE29ohCi3gMLgQBUjGETMaY0QIpVM2P33qgxy
vJlepKXVr5JPF5QiJ8Kjbj7g9N64+xdHor4fuqTYD6+SXXTmNR9UYqEwHzyuUbPjvyrxCcVYyjST
L1NOSV32lSy3tCE3tieZVVotloDznmh8pSvfnID9O3l8mforN7WioQ900yiz8iueZtMiuV66gCOx
qj3cWw+tTMD2wvknXzwUfDbU6OIgdYtZV/3uwhQkTyQt+JzSEVKhua0mlaerj8queMcQFqbcqqnH
CwDeda75wfetKJWGEMzRRiQcMgIZtpyROYk4dsxvofbr5eCJ1HgRKIiaYxl6h9af+Hg62GsGpK7i
HeBfBC8QZqPY5Uy3gGYUDHRyra0qHhwDvevIIfa8+N0m4+ISwgRVMMYONE8iIUYBPYO8MKxeolYk
IgBY7Ep4zxIRWW1OO/eLrhn88I/rqbft29Iy+zPqdO9uvqABUT3qnzA2IQ/S1cmq2Mm600nBWOF6
uq5gw2og0rUznd2w1rHhGcc5/IKeFnLVHcqguNPh2BeU+wCnSpHrRRSV8ltLhTmud2sj0U6L9QBB
Osj3iowWjgtXK8PUvqHWOV7sdh7DQ6zZ/2pGWlf4XEv/5Djo5oxG+/234XjPBg8qAJ5mb9Z+pvnn
L1wSuJ7Mgy54cKW9jf0gp8W4yblLe75yfV0UGTz1tA44H882v9Cr9YK0rq6GWutNkujuUN68UOo1
gEhPr2wEzvnrS54TxutEmgN+LK4L2nyOzkkdCMCy9UkFZ9Euyldj/z9931dr5PtFg7YIHCe6rfLj
Xx265sUc3pZp8VSZfp9A0q8SurtLkykNkT7JWqRkm9tTNn8MockqTY/52UdpElRckgEIIIZNZBfP
BvXpaTun9hwlLKy56evnD6/OZbH6NGWSSEWWw4oFJx347TbzECEYO5OPoLCRJaem1GromhVXiUqV
71p4vEmyLPxoHEG6sgYBQ4lf5HnlPEErt/xlxiF6ntt0MXPCWqsyPfW/bMy3sj2q709s7hsOm5iD
oEfJJttKMu3oMnRcvO3UhWpSFkdzzm4wHB9Vl8+llQvYSy/dUpbYyxYqNO3sM5Ik0WndfeOdJCUp
l5Zld2D3hqBr93HKaTtzBKKfsTUIxWvCEut4rQlo4GwO59af5KArJhenKcg3Au8HaBGIg20GMZdl
iTo4iEpFAdb/0lpqyEruogPHGZtYKL9VAiDC4wVHAQIWsFUwy9QtLRUsrjM50Rva/xvMBbNUUNYN
bq1fpjnXy5/biioXC3ePPOGcXDADh5+C2qB8XDolZCUTbwpU0N795RPT6L2boqzYoJgZpzutb+12
4yhcyFdiXX/nDFc4BO2iubyQmnJ8D6yxyYKZG1dnSn7d5RkwCdh++tavltnzLZR+eBJgosxFl2Au
odq/TCdzYJh04jAidlKXzErng4fWKumHO8fAwkLg8q88slVkt+gqMIHsTUZvyJpwCi9GjaWk5q9v
bhdpBmU6ZW3rnE3xjnpQ7lfyQioSouknrPM2qC2lNADitmnXP6cWxGO89O40+Ao7fo2POTHIQQII
6z/YS36QsfxKG6tb5LFgbkTZyIoyVVYPBjl8c/rjlsjqeuAwvW9JTQcqvCeTF5FGjBlYi688YAIQ
vEfyYDWB36y/DxJCqF9iHvYArd6ri7TrBj/CFCLG142iVl0X+7F5BZlNNDfwLeoQaBO2bfLQPWaD
l/N3zsoPVxYCBljkkREybDB3GDfPi8DCDvN8vrWZK2a7vevFXBX64pKzFQFs/73SRL2DfLmIucTi
Dii3PrnYM+BogYJjbqcZ0xQddAgmmrTksvvefCN7B1I+JNCeaf1e2/Q4EqJtL0531x+7KVShZxSj
AOQlFuQA8X+nlDtjVOp/DllIddEekbBDvstf/Ir7yGUpHGqVJQyclJzj3Dqfb/QCdAou12tI9Jdw
rf6SyPRpvJpUsf+PyzJuf79Uc9rbpq2fwXCUqKbDq2aHa3bJ6gK6BR0TlncBwKnU6hjNMd+lniKk
RZIxEq/XqKYsLevUSNDsQGQJEcAFe2+8al19r61AL/hH30Z3sZtF+lh3JymWtvHyMJxsE0fcDP34
gonf/X//somtAZKH8xQLU7LquJGyK8MmqkFJHe+Z4cNAa0w3svFzY3t7T1g3TUHgtXB47vhA7+P6
rinkkipO2B4jNdEE9o2zLTARE+l34sgFdqfvUTvLAAO74G6efEwqBgLci5NNIGACdGY+x8N/TtbX
AuYCKz53830IEo/C9/ReG+Bhi6nPnibaNtDWLAr/8CCfJ2smjHEv2GE15ZWpq2X3Ih98kOJHhnAp
jfweLkEUAsKn1DqxIuJ/aSCOadXd002hvXNKni7Z8we29t2oxCyMQLD1fZ1oyvyaqPm3EqaN5ih7
3Em1NURow7GE2sOY9oK29RHaazHlUBBkskPath+7D+Gt3iSLfZNY3+UOERIQM1YX8NF78oKBpy+C
3pULLGhUZea8CGHprrYy/gBV42U8HYFigrQbvj0IVDP+z4TyNiv7aKA0EvqQBV//18NDzWsl9A25
y2BFIZyqvoEORb9B2prjMGDA0XDQlpuSdmQHbQzu279wjgPuOaqB2H6V/o/3azD5htUyJLptECmy
aKMBLIZhdj6IrXwH2uISuXYCqEtmMaeS6059bdRgrG2FSKlAvlOSlKaD5MhNVFYbB9spNfA0ANvf
HuCp41abdnaUBE7qNuJC3XPkt1UueUIDoUAfTH8IDLkOtA4wiWkKfGJhaeNOlBJFU8R0Yl+7/UXC
r+kkjmWxuuky4O7zDxqJv4g7Kzotm33MKHESMuagM2i6H35Yi5FCm1MEe8h8FdAoKHHGkZNxZwat
5KXuLSDOnY6XT83D126t35+mn5IwlO2IGntc5dDktiCVkm8simI/kJbTgUoL462MxaXnr6Nhs9m6
pvooDa9AXO7kRRYkCbpuFZD/nx5+ceD7qjvDIXYrvkoeHcAPUojBJCPxMvPnzuACHWU2/P6PkpUW
1MbTEwW7QtEvWXl9T8vy3FiyyGyEHhikSfIS8UW4TXLfJOzgwyV6QoiYJDUeLxS0pveelidhRJnv
UPUO3a1vlgBnX4gdup3pUpS3S/t8PSdEbvcugExpQzQ49C8LG0PkV1JExmMf2VVJMos/p8T/g3em
pHa1hOKwFKslfI0qxt8hqyWIAjFZmsS8wEkLbgRIsyEjDREWXp7407xYL3gYJnsZMjqm2yxemGBo
vdu0fW6AN5dX0VUXqg1qFEMcTbsP67nlM0by6bO50Ituk1VwquOxnC9ue16gsBBn3dy3g/gPArv8
MqzJqvxerUrI/UHt0Jrz4hgPALnXNSHCkJGhlWfD0jif+CeRcTzJsx1lFIE8KYDrpzAcO0mvINOD
eGqykJ88nErmup/GuYQwtGWLa9SK29onS3vvCMoT3fDhcE2c1oRO7I9lYx/SlJAdEJwhB9Ti3Zjy
H7++tgIO5W5riqcGhtFNVZIoDUmDc4xEh7dxIxGiXFQENfNE1Db5L8NQlxobxcuYeik0Ew0hPhRS
4fA0iLDH8oO1pbYGimtbEiNcPetT57GVDiRWOMh75D8athc9sY2VtEr7IsFuqNCbnkUXY9deDvXK
RpO3I1d1qu9juRmGItw2d31OX6R90jwG5oYF+aB777NCn5pYZE3fCHgF1iisHwzoxizu8MusGQCj
ZJdlxANHZmWOXxJzxMCHEQYxwpe+F16SkYChJU2VjWBgbhy2upOk1Lg/dtis/BC9WyIFhUjSYkLz
mvlp3SQsc5Fgt52g5lrcE9g5LloATQGHNsFrIdDVYWaWaAYuIr9zqH1E3wkqlX6/4sDNjAL4QXm3
U+YsH92eQ3tikZBa5Kzl7OHySWTMusCXdVt4zMRe2UJTrwsh+U+RcdJAdlHt6ghbofjYjT1ocxE9
OT2dKkwOf9PmebVDxQiYwekgAbBeFS1VmMdjDVTc+xBUrUgwsDX9oK7OJ9mFrkHGRmS3ak1SgYHs
2DMZfPyfFhxTq6yQLxC+vh6JLrk61foeEfWMVLw60WU08urM0KkceWaNGE5QL/E/GV7W3DCJLNtA
mytD/QwR3h9WC3vmerldsp4d9TNOyToNl6qKJ8/MU8IiBUq/kReAwG8aWsN3YOxlqbIptHVxyBSH
aTy0bFadVHS9QUCJMOH041iMQkjkkMp/WoVI9LFHpDjGgz3/8Mh4xSOT3PPI87keM7jBAEJw/d6y
hu4fTsFRxAhvWgkqMpjvaELbDWhrGsBP8+d817cd75rcl34wC1Y1YuM+odrWGCb2AP5IZLggMPYv
VEkZsyCFUOCGkqUY40LAEkZjBRyZ+EKrE44vdTDtYC6c4VM4N8FwIsnx0FUAIbuhOgYNnjcTTUIA
mUz52wxHXUUrpb6GKWjsoKukHQ+sofeqsFABjlbEYyWZmyCus6h+kuCDD87lWl6vYRnjzRBSWRAx
L55oTKMzDaNDv/oekK/cWU3mKzuHVLrSpJl1jkViy3KK/F7UHsPU2erVXmzEyrmubHeiOTmAZUld
nLXEumRlzyLmWzi8h68b0moGYPPrnzKgezIkTAtz8IvAW/+U25hr7im6xrvwI6Wq08uU2TqzAgjy
dZARQkR2KN5QIBPfxMfqJky5bkG1+9FD88HK4mfecAfLWjvlh2x+brwthtDJ2jQUSakwZ09C1HK5
xAvOlE2XJ0m3WkDr/94+4HbOTg3u6iBt8WHeJUH9pRYmka/qeS27r99rWpj3F/IYIYrkn6NLeOov
oAZLfXphI6Upx047aEhtGRia7mKMXS75M0VoNLM9BQhankelRaf5tFffYsjgL9XHsfRiAu6r8Rpb
xlzkZV3yyOoR9kGZ04QSiKvK/78JFRKmliLs18WremCT/HE3DyzZkZGXirejWm2y+6SyZ3DnEeRJ
MhTX4xg6Vj3U3uVQM5NRLrkraRXFRwBEjAvhBPmZgaow9Uene6se9oSR1Wy8KHOR0loC/aYqD1JM
vQFnyBfywiEXE8PbTvvN5TKf7QttF+oA/exlp7vyQPKyaLbn9pJKNtCRj/muo9GcSzXrjot2QvgT
iLicv44tN1tKBQvdqQI1aW3v3+poKQ0VnXsNcyqiqqyYd9TQdZ5slJIoYCRwzitu9aOQ7ukW8MfP
WK3C/De1yjZ7+bNr3IkfvaKdkEQf5hwWUWVFq1K06Acs0S0h/3p9Qgrw3yKCH733GtoljWqnLacN
ZypyXsIS3GMvY2ipOGLePutEOj2kOXDcDezl/C9ZyZQ1CPW16vjx8Ly+4R1QNIFhYM4mWt9/G/yE
k+kNaIfZ88txnZhq4bh0PNSSyAYkaISxLyKOcPSccjuWxqE8jL6Cee8uCdpi5dneHShOVozcJSkO
ZqESQ+NhqY+rvX0RtLDGaIwc48pKuQEWNcxr5KQ+o90VBS6HTM0PsX/XrhfZ1zWRjQbIuofhVWs5
HbQpc0l6kxJLX2WBRB+Vt0ci0qMSVn+FvkssvKUWZzmpmY9gkxKhJ6nOgZB69bn2wpsv3q87YcXn
xhNktfCoA5PX/14xWzSGPticoI2boDHxsS63yPdF9FXBv63Kyd6VEl+prx7TJjm3P59+bkx0TK4H
bb1QGwBngzgidPWbjOKjXdM0lx11ZqKaMSk5w26joEYiYTkSU7BsnUc6eus2RRBADUNqyi8q4eo7
pXRouyJdr/6dgdCd997DpdEGCO9AZGS0b7t69og8CLbs45RadFdLOnKPeiR7gYnlrljEBpYnshr6
UwvAsCuUqiPx+Lo9PeIC+Y9sKUqGQ+YzXRNxr5b557xFMEiv1rxmgMR1NGV4CmXuOxE1rcbm6UAU
TfGNcd3cPgQqcy+uZrrF1Cl4wHSR4jdnw6U6wTieEK2xJuvlu34TMp2jDu0VLE5mnQetpPz7kp0o
8qBjemx29ziwydoReuiamBGas2l9C7H03XVVfIJ4ud9N9UxleaINkuxjIutjmhMEJibewKj1Bmln
5FiHzhkehbahhzKa63hFCZVluTap0vCLeMvRUeppZTh5LXjejfPt5lAk69kqKLeeUjxoyYSY8m9n
EkpzE6KZmIVtChMm8gmI95MWHHyI7ZsBX6rew5x7D2S0ntDterXZSBOty4E0Oc7lvPOZHdPAc6xW
OetniDRX61Y0x7/V2LE4YuwG1e9yLGyy3/ZJkzhmRGEoTvqhOq7O8PH2we9KooPGBYyz6z5WBbbZ
4hVsY9aUXSSHNYACEUI6gmyqGjIgcqfVmx5Gf9CQhTd4ZFuyS3dQ3fE3o670p9WERra2v2D09Yxm
d+OMW+pxN11yu/hd6pC5cjNbPWnDyLjUtNU8F0RB6cmRqF2bfIwScfpe4ko+RFt/1+N+u9IaMOw2
UZBEWw7dhgPW+16jT3b8I2eXhCcrx7w0Hx4EHB5NFCGS4oX9Os6CocaHffXXyG5UIEJAgdn+HR7V
HAX92Dedperszm4ZB6mtWiwUMuDI2wX75wa4xvXxMHvQrk8rx95p3CNc9dNhT4hm2zDwRAT4cViz
g6FToYpeIKBtvLw0BJw7Dxs+p8KfWLoVCWyYUj7NvFfuOabUEB3rKxgxYvf65Re+/yVHmYviAKtQ
0gURESR7+aFsARqYzKdZ5A7zLX2D5tocHnn3gDDqDj0eweW4vUt24riTqTLKwJgQ8tCKWxARIhNM
JV/wtOwDAXGaetD0waSGYuniIyjaS9UcfxEUb5kPSMMcBG9+Ht77LZ5zmxhx2gFZ2ArJdWNtEidP
cYbVZ4lzTmlKP0CM8R2F7QRTjXMi2C9+2GW7h5UdY4yoOIPp0uCsxS2RTYe7CKjF7zohLNZgJ8sG
HRZRfsKg/mMStNR6LKtJhZp4A2+5s/znMzKRuP6E4cI3tmCm53TZOZPeaMKIg45IK7CccgClSwan
AA1Oy/Ch9Jawt9ntmd8kg5BKjQaPwsnJr/ppYL/ktL8VOOD/6ywjMBwp/JNUMUT5jETqwiuwZye5
mIYZLSIykrndROZNzBfKwYu5TML6DTCl7SaQXuAC0XUM49XqEWQLs+W/9ohiBBvIqtOGF7sJKXOQ
DqF+PKUnt38XsarKCtWhj+DwKnV4OdQqsLtagLSGQRznl7w7ac0i0qk/qgOfeqw7d/qtG2iME3KV
f78vqhnJm8+P2WMTjFyjRcVXwcDQcXmUckBLBBtcKdM7j9RkE3panT9CXXG1t6QTvnRxoyH5c2tO
1owo2oTlWIT6yRwrhKb/ZNgS1g6bvNVSmG/C4b/IBBCrvSBbVyplLcqmsG1wUfU3KXUpoqxfquvO
+aMd+JMjqXKeMaBY2+mm06sSdpp009j/3E/JTVeRpz45Gf65JjRnSWI560164RzOjpK3l87ppMT5
YmxjptAb6MVizzpgnV1T39xS+8FUw6SKjFtVie9Y9+Rpxj65BUONPl5ErLxkezx6Dt3LqD9QgA0t
eHApc4SSh6REL872QDnC+QVathU0SDLKkQzq3ejsNyjIzOAI9r1SI7+0GWISTbsetxxi06KyfUPR
Zb6Lzz+zwA3YMi7FPZjykppPkZ31HQ7+HH5CKpcsFU1TQvW5/UBGlZDaVGRcK7fajN6Q5J9tAQ8Y
LpemOt8Jg5u6KEKUjHvncorpu9pouxPCS/7yRURiRiCFz2vEXRETZ6nIfiNKvQChLyvi9N0+1aa+
wJtHD1jqHin205Wq5A4n/JbwRwtOjkDuKaMgWZhVOxdCCK6hczyd0ZgG7doPoFn3k/W3lozlG+zI
tm09sv0uvwUYF1/oIGOAdlj4qccpgu5+8OM/qTTZi2u+mFnWn9d8wnjBg0OcxC8ftH2uBtrQ8H28
BLzFzSWl/bqzdchngFbAaVmwTArClsBPf8qone226mj9IhaLnB/nKIM/EF8SxY+PXrJNfCNdvBXE
pc9cu+Sni6by0LcuoKkJ3C22lKYw8QBXYQbsXQt90WXQDIGdfkdWR6tsGqickSg5VjMzphnFA5T3
sLf6Cl/E7Y2qRBQhWcIcI0NgrvO9VvLJru1LFcWGCAoOgoyWZWhyNELfizCHhpeWfJYAPQ1RJl0b
LJeQ/fj29P7EQ0+y1O6bZOrVMVjWICHowEVM7g/86lKHgRRDDo41AEGdAY1tJ4JZS/ufwTEcpV5f
yTF2qlHfpblxMwA8AkjwnQHyUhoxCpuP9BNdmL/z6lu8pWhIWqRzH0cAS6VJTJC4gUa6nzipQJmj
yfuPfDah3hk1C+bEMu60uSfeJB4mCnuDslKc8KfRqy4/VzjwxzxBObMiMixvDLdQYyDyfM8tqMI9
7lX69Yr3ndvyaES7HazfLw43IVKWceT6smx2czvh/aZUr38FDA07Jb60A/Uq53speIMYh0IIEL88
j6l0UUa0oRFbCLB9ttKfJFM9O9ruZHdBs47oOPVpY1Aj5mOodxnSOqhLNB1LNZD2di7/moHUWR++
iSVhMfTYw6xe2DkB95AIEOcnRY3dECTyBacwWeEFW7cz9lPduo8d1OHZyBrLBOfAFpoo8Msa10Ul
PkVV2K3kS9uKaz6N1NBH/UfxYRJBz9jEgirULW5c0KjIvEZK3cvp8qY2cyhnlZ7QRRg07ls1c5tC
j+81ZQ5L3Ug7XIsfe+bExW0eGMn7KDYz2IEPgvjaQkXY0mRzKpaZ4Uke8w+woFvvnE70LUbyRORi
EXAyI8AplqNReqhDu0u7GVBHeiRnTKqR4G+y8ePleqUGuo4BHayPbyGhv98OmoRKlS3XqUAZP+cf
PLQi2JV7Qiz+UKopjQKFHYcYEe+6FczFJBdGuUC0WrdloWYtT2xMwQ7SBAhcIXqR+0auhcXV1cvo
ygC2iqNlEZ6Aq5fhkrcxtUaz3MLxC2WVjTcoUpAaUVEeV5c+5tvyllpg8WOb0OIAMvWFm3gOubnc
o8rlv4Bj+3J3omT/3eT8orinMGSUlKdm8ux3ITnbKx+S8AqfHevcWD1ftona5lX5pgnBsoTBVrkV
j5/ElOEXJha8g6L9SxteH5UDrCzp5YkhQ8M8u1KqEB0IIFhVwwgNR/+wVdMZdNdUaW02mKkM8S30
IcRu6gh9eJUzJZkOp6I0DIcX+rSao9z4Z+RywP6mUBgcsTC5T+Tzn7PDAsozoYBR1XNhFtCeKA4K
TSkSxnWHkvigSgKw79qcqvoY6j20/3cK8/tvXMUi9GTcsPuBLbc2No0Os/PWXuRrocp5gk5FWZJ2
e+Jy8CQC5SnnA73CU7s7fNasuSvISEEaiXd7+BsyqbyWSOxRUCwKtLGZqdpXewPytmSotltmArf5
jG2gNlPSJPQAl56DOmydRW0g+3kuwuJZakqH7tCeT7QoHd0qLxakm3mbzLa7HwLx4p9L+DssYFBP
lWQ/R5JDiS1sTJDNtpE0Rz930wW8YZ4SxG9zkto47mem5ES1Eubxv44pFD2EaGHGBX1sKn1QHcTM
Fcer6q7iEm0jjAofNX0uDv/TTjivgIltIDiCU1W+JnD5rkTNnK4e2QxEFFeo3gj5eej3clA/PYeL
XOCL31I/h7kJc6+ZyJwWJ2usbVVGJVK570ZcsYdDcBzCkMkCLVMd297dWb7JIRzE7X8hzB7eUCYe
NuYllIQzdmdH3bab6IobnXQ3GzyQfPdTtcUJSXWOLsax726uUtjY53npwyIWEvwIYwAQWWt2bc1/
6FO+srxVFFCNvr2eQzDm4NaaYGNgXfmegNsQn3DXLhZGgMlHTvGqgb02DUveucU4QCUbnY/qaxKe
P6gCxBvIq9WNadi3dPb2B8p7oHB7bjz3JBpuO2qBWKIzht2JJFd8fxxHQAiuKMNrDx5UdO/pqEFt
HRUYn1R+MYTI773QXnYidKNO8gyOgQfbrVFSBE4kXBlCSa9UFISpygSmUvsuDc46GB+mb/eYkNFo
m+en8oeAhRZQa1t30FBLNDXXc7nxAGO7RpMsjIZxq7VqrCLNZL3eb7QCYflnuJIMWnv1YnsN+CYd
dT5/u8xWh2O7FZApBlzAYo1FE6EEP9ioaPfgnxnLDLEeTPbi8bQ/5BDwIYQzVuZVZpfnMuSGBcfg
PagWuQcWRb7bFrAUzMj32gFNkifJ96MALYehc8Auu1u+r1Ib/0u1o/EMC3RFCSC5in0E5qc0nUFY
Bfubk3iH4XkKkncBUpon5bhsLT1rjzdhTPlNXq4KYn1hKmGmh6z/456D3yHXyFRM42uulb1A12tz
3c8x3aBE8qSztc55ihmqNuXQKzFnUIqQwsuhyHiypjeO5F0nxzQ/fbTcxxL8scB+XKS1nRVshM2S
KBtnWRd86D+mGPmReQg1J7BsUZfGs76a+wKOwn7NFJ8234sMvPvXFM56pwGMUdpVec74yBLM/SJj
gGbhPnFggd62AyLFaVI3khJ/c9HubfkTgVreMnVX7HLTzUIRJ3QjJKdNjZ415oYL/nTI7m+lyfah
18Dqv6hHCPduJGYjLgdtvvLY/rr2wtmlFZ1Q6TrJ71RXZHqRHXDkphDr/Gldp+JNwohtlDZuuN+N
qfZRI0wXUaaaPconnWZRmap1pVdW9FpGFPVTYfOphJKsnv+2cD5eFow2YumXM95cMxULjcM5mxkp
vEUIkrYx7uJGHngMXiQ2uIM9gaXYabH7LFW6CCISqUntgUckWy0rjqF7hBo/tgdRGH6maC7uPowx
Sb2r35CaED5VnLcMt6YcaFUG8JiSpymRc1isghjfYzz0sZcOe3BHO5Su78Pz+pawpem/yzs7VjF/
7Ldz01oQgDqWrQCADPMQPC85KKibxSGBVZVvMEi828Ee9CE4JsC5yRipVTmQTTfihVQaGY9M6xaf
W+MeZeSnOYDyZVFnmCqafccMYepBEvxMK7WUAyq8OVBkxlr7eJyrj1mE8+2EmgA1VitXXdyf+QKI
c0WEmRCRYHDMBBTUjby/StNY84ZdVUv2IDVMRgTrDa0QigV2/bCOlRT7ID00vdBpyZNl7k03WKh+
QohR3OKNvrgmpdtsMimmvq9I+YFCO0Ci0lOU3fXUuJX/EN9M3ygjTkfTwUP3efLlB9um9mb6ZMlX
coaQG9XFQ8AMJ2cM3ymeiI2XCrrDB1N4JVNj4tfGOi5+f+COXzA5AEwkzspGNYE+13Gg6d25yapT
pMxabTIu7StQXBq+OYKsa5bzrfKX+V8zD9eM+NUvZ6In7h5qpLvdTnOfED7zk87OiiWa9lR3I0jQ
lu/xXNC7tTOXF9qIffIf9H5ZHS5ozCmviyguqhoZ0yhIEm3Jsb+4T7wD0AAMiyhMeu2c8hJ3Semb
9cHppxnsDhMCkVkd9t0SgAsCTarPknPydrayw0yjOiVtVTwgP77c8z3HTJygfonHpNvC57tOdae8
hDu3Y3nlUW1KNxCTU2e2WiMiDw12Yi/d/H0kYrdxP8hWpWk0Lh8v5cioglQIzaTPy2LV/FN/OWLS
D/f6tsSQkbJvMIh33835M7athMxcanvmjUfNi4a4/6YinGoAUOJnUcUWhteTZecSoVIumUnqpF1A
yeHcHAI+2EG+/BBwALjUBq6mT6dKnE3lZLHUhLgTLypLDcoktKjlY0JsG6j2bsAx3nfPJw0hkeVo
VudUq7KNQ4zFmqAYiatAYpSnAqMGWA76h3N0yGeJfhU6ivvGpTJTLrEIPuhTFEwJYMUb9JoBIRfd
6ShFf2cN8XtkAReIfmsunxs8NiWnYlbMtouSs/Y/ERRYaHbBBfyJyZxrsYUnQeeIURABoJgNvrll
2+PrQQ0Zmi6dwvFJakeJ8XAXvuAC20t4O/FHOOdcCpEl5nLP3Jr+AaqyFerBGj6y7x/pz5zHopCh
jlpWFtbpOrbprACw962KHKrxWR9YnSTymaU9UwLV23YvgLWwWT2hJuZSfO/PJwJ5R4dbyEZzCV69
CnWxKwOwMz/s0z9g9Dx9qAV0JU1LwaQfleHqGEk8O5ZkfE7zaay817wO0JBjNNP1Hjhc4yd9QH5q
x7mkcKN5YHBPRxfwUctypyxUl+l3xy/GDau8SL+inCBk2pQGJ2lsL+CL5jd9pAWH/aCrt9OuOVxD
AEzTu7pHmZrlF2mfZUpYewFOZqHRCbrNVPkzUYzSWSyEsTuEhAJ0lSsx1R8a5Jefde1m8NfoGrLg
yJTHFFh8is+EdqAcbGEN2f2u8PIcvfepTREKXJuakfB+D7/QPfkCDPX+cQ/lUIbWRCsJf6BzOhtx
gqMGTW0AEa2FX/GIHwEp/9sc0a8gqtRTwUUwc08uXGVyYvC2PkKfH97dlIdaLVqiEe0m4V0nLADt
sw7wWaJDOhCaw8tdROvYM1PwUEbWd7AoBn7KzXCxXaZu60U5QJTwb7Af5JwPmWuuDOwihNImnEZQ
X2d0OHe85YYsLO/G6/XxMCnlt0r3bLYlCEjEgTDmypod+tp0W5nhN+zVdiZ5mQeCdjuUIz6Y2kRf
SG6OsSRwH9lDHUcKpWLqz43XXZfh1BnABvVyXW/XdkaN8kcGL2Cpu+sIccRCRJmEXrnblXvGYUa1
ClVFMeQxxGafPxfnn1ugZhSqyuwJDj5wSU3dmFKSIyYSwuB4bfTV3VjzrtsSifMZIFLEtZV5j2/i
hvQfcSaEfJl/Oq62iSf09fAKfGTdRV+letaKdT7QA9wWmNTNhsnbTajj7u8iR+xGA9KjfgcQqjS7
gFomnN/jLlZ/RYxwH31tk8qbuypt9HYBw4lpPmkt6lHwFwXMxMHTGxspriEpZr+eUlHkMSdRHIoZ
BQsZs/0N/31vVOU1vz3LHOU7srltGTNLOURdxcnufRyk9Z+vJFD664FY635hK88bJE4Y5YWTFIv/
35ogf9sJTsa07qrXbFu6ivT4Y9J8aX+vrgW2eXF9NljZaBxN2GB9x3aj8bcH2YZ62YLek8Y/PaCc
LeLOmdZpz0GYwZT0rTfR02kJpXqjn719VrpRcqz7bogxR1THthixiYRB8+QSQUUFAzipnniwjoox
9ohIGR4wT3UHBgFgnHyNEifMmuEZ1tS0b+qxibqVNbAqxxc0o+ZlFTf8ZfspkOmDYKNPdCc7rGT+
MsGxk/QhK7USov35A1c1AkYwDgvEAWHp5IW+dlk4ypyQg0R4AQQVPprjlA1KCi0hsep/oM7/28TT
iFefvUb685iLLbkJY4KUw60hi30QT5g0zKyjGU0Gxv9HW1PUVnmghCoSSHgQR3Xkym4qjw0B/Nv9
8Ksn188vSLM4VR9/LykNRDNw6SRWg1TupK4Pmf2QQIbhzANcTydkQX4UgThML7Mfc0g+I3u8nuLI
I+J+w0n+L00K6Yn4NqHlmdR/tsQsK/MyWz9afsbOT/bCcIhomG8gj91QtrwNrUHnwRixiR899qh3
CsSHRt5XvQr9nGinlgDg6sR41TGcmciDnqcLSU23L8Ek8erUPBvXR3iLI+fSvKlotSa6PnXik54c
rSahUTWTm4i1dAGuq+W+pIjzRcU+D4bZ7VyHJGGpExD2p7blla9mywR+7tD0F15jHLzoNBOKBLK+
nL/qN7h/I28qUbF3xfGEg9nLSEeS+KS9/hTw8TMKjiZ8Zvkhiolkk28gGTYfiNh6ZKZwOWDyDw7s
8GBm81ihq3lq7knulCgYG+6DLo5RpPYs9fGv/2zBkzJQxumCFIWBZHX+VqrniCO8RMF4Fg0nEp5g
S8vvC1jpCjQpTKom/E8tGv2Cd2OPlGZl1F5Gf4bKDJPxLJ0r0fs3XdhjRy48jU/73dv5NgwQx89b
rNfXDQ/awIZu2LoKWswl/Nbh+hC+xi0S5efdrz91uvpVDVHcUT7Nf9DuUA+PaP5MPiBk1DPR0nk/
IDnoBpyDZr8YODqkGCKg7QdtORCwQ2EcBZOX1xGWakk9WyG9qYXQlkxoIfxvr61VedHyMfF0YeNH
fe54bn/BIN23bXJvCctNfUSjHz4obZisjJ9hdn6mplxH+En/pAVv8itr/5DV7vTPm2jQ3/5YCT4h
5Zxvaj2lhy81iwJog+3o9m78+Z6hZ5EzDHODso5KrcKCcRsEjTQmxzHeawWU/nXhOHlktGN6Mq2O
7eZW1BXxDWQMwTPHFEeonuKP1a/qAXl4OLzpKqHeSFKm+ZV3ljrSBXOx67B4sjxI7FimLhHKl3+y
elJygoiyFsham/XEJdluzNafIaCzxWry7Vi7NQQ4teq9KWa27zOl1XBovVIhpnzn34abMeEyW43C
UAAHM8TUuR4XqKdF9ksEOwsvxwgI7DxbA37F7Jf5BOkQ55annDV3O9mNMOU2cm74QFRw66+ib/cS
sy7vhotMxnrxV2UXgjqXcctCh8UxQVLvOHylvHdjWyzRiSDB6wiCBU2XxsTgDPwbgbNhYdfHbBgM
KOMaNEjFCs0beNADeyw5I7HLwqS0Q3VZwve/yHcPeUwyHcRFX6gY99SRXTvp5fcMUOGjV5SbwqtV
204XcnRTB7ZINzLfZv2C1c/JbH7v+yTKhUOduMguW+/hyCDmDFIsNaY5VrQ+PwV120viUXhzTgp3
QR42VZdswIqA1+Sl1fqE1Y7POTQ8J9KK4KCLqo16VsBzop9bMBsBQZv2iG1RO9c86qJsdKVLObxa
Mckqj1cuh8zqac4qoxv9BY5JlHCDzYsyheTF31/NOci+D8XUK0NoZqpArT5XsudpQUyPPQ/3Nbh1
Gjyi7YZPnvloa96NFHw1W9RzFYbkPP8308duQC2NXV95YW9SxEgVKHFqiW6Or1NdSBKbxhemBXgV
dhYxVPIZLjsof5LayDvk3K0sJ6QF43t6bhHkDfABeefAi0vyjBTNVgQo4Rl33IcXXNPpppMLkiT4
LvA9+noCKzVccdlaf7ealfxIdzGOBk5J3rHYEYb9nrZJ8kLoeSBeH3bHKUzxsG/DccvrCAyR1uCp
Uuld6MjKLdF3N9jAe/5VdGc1j4j+k44rwMzOgYGe+ff9la/x1UWBk/RQsaAxUD9qsK6X5yy9O7G/
5EUmvp+dsY3NTfVra5hkzPzMQc+Ob/P8titFFjgxR4v876i0E5EwHa5vgVZUvYdUA3IUonLWC0t7
VlCrbTpAn/bGKLbO4LdZyDs8m5S3BxYYbSt3hZrECqP59DIlBdPj/mkpCDUPBx78IBxdhzUNsLFY
CWKVCMAM7DMmp9OrOlJG7zxuJnBRVcdOmhjJyMXI6MONIi/HJLsQE+X1pViXkq0ss/n39+2fimfp
QdNfuwKC4LvfoScyd+XH30ODVprvgBMxftqMUWy+69sZTeprWHM5nYflCR12qEDCvMa1o0PwcEiw
s0tLS0k18Py7B4KC3Z3ODhKcWlb+Nc11RtEMekHyHg010YH7ydtJWYfeZ2VuWPQJSXRGA+H6YvkE
EZyC25O/ZhY1GNloV/lMuM41NPDbzQcGfg9uwTao7+xFlGjZE2WVEbHDbtsU/2i1fRjV/CF9oTf9
bOVeEEc/IqP5IVcVzwGgAEkY9sHOBM0JLfP6jpkugcIn0IChJPCw2vsx4HTI6ELCw3aA+Nuxlaz2
plwVtqs2Aa0AFMXfvaDaOQsLXzd6tHBusDFkstTOrVwjU6YxZ7mMJE0jGtFZDJCv5N5LghKsrEn0
6vmlb9n7aRrBtfz4ucZZE4cjcbriIXtaXVZhmtUlgFZKSEwo3sR8qZhPGnHfxbrXrnZXKqv2ns7x
/AOV6l8a0AdJsUI2lsP/XfOGsoHktgF3DPPkevD7myYtkxmRP5FX09zxwPnSEVv6Ww5dqWRP7hnC
Rwccu1lLdyg/F42am9luCwFhPfKoaIdn7rXBHF5QYgMa52NFtdNB15ZRgT3FO7CFN8ZvGfRIo9Lq
hFombDE7QUYex1mM7uuG+Mw+AYKxMVKsuopxtPm2PNmG1tAfDqXcmKCKvUtNN7lgBNhhprfxZ5T2
mu8javDuFTcXbDE8vbCU3zsqvPUUHr9NkqMLDkFL4Yq7lpJfVrs3ETtKpKnT7Fl294JF1ti5ap9o
M7UKAnKfC8csWBBq0P7yoW7JA7Af07Nh6BvkIyMTKIegFN8WTn1TcB0mQekxFrF+wAp//QN2u4iF
EnhgGs/t+dMP2/MPjP6ZnOoSKfG1AXdpfQnclgUdaFlYHmONOewsJ+dBYbqIH1gxOCCh0V7yolv3
2u+H7ODAvFIDOdrQuwbKiYh7ivCWtkrp+C8yICCPilmRJQUmpayOLkM9wZfx/sX88vPNrIEcNBik
U0cs92dNaVtW4fRFhe5V/Ada8fave39gpUoNCq/ju+0sR4iqhg5H2lZyzkTD4S2j/woyB77+yBx2
A/qFSwm/0JbQQ8KOBLwJolqukdWKzrMfT9DE1DSIKaKSSi2fDPOmCMIVML/eJ4IwKvAWaUEYakwZ
/0rWrhOZAHGTDLWSSuG7chzsqW9DKGTjmUXX4I7Tiufkh3OpKX04k3d30XyYU4khOVNy2svYNHU6
YgCDSEvo3af8HyFF6NUU3NQS6qVN+InYaAAMFUX5p5r9WRhPDj9Dlo/PBkwAnwWQfyjVLb5+LhaL
dK4UXRos2yrlbqwFZ5iDWLgTPbSuh7VJ9mkRDncbL4vqxuxz94dHl9ynwfcf4sOAgwK/MXGwLxDQ
AQobJWyWxLNhmH7ylGuyAJ5+HsiwJhOeSyv9Mc9+yJQoFj0BKaDp1nPndqTYmTM5qL7dT2pFN6j8
lk5llhZG0qOZgCA3sjcqHVYF7uVUZmdaZaw202HRgcUxK/UuRigAMYIwzuY8vjbXSiOpwOsdN8PZ
4c2o+beceWu/4P+9j5QKYerU9blJROw9t2F9//Z52Nc7wGTSFHMDgsM0hr0Gxqi/niFXtuXAIXI1
I1DD56X2cSX40NoA/4tK5F3mNyd991Sr6Be0QkZtEYHVpxGiEhT/OEAStAxqVT8HMjkJ3FjhHUIc
dffwW5Cpw7tKFckdUff4jBI4dBXKDxhIgu7WPhZaTWuD1Eu+xTuvWKsmMFLuYJwjPsJYVumOwtyX
J9AU7cQw+XoYyGPCLY0iCPluNWjZQcmfL1kCaRDb6l5jw+v5asDl9JY53RWPTCAb3q98c+vAFtsP
kjnOUUBRudxsN6k67kywqF965Ws92GTqawhuQyL1GnF42BXPWlcY49ukVMWv4dyqNTH5BqW/6Qja
Ejnx+wnZsZiAg5agmheLKTcBl80rgtsmJFXwhKF6CbTy32v4Mzbt1pTpRncWrSw/GB0GGdTilMCM
4uV1PVTZbWY5o0jIdxyihT+NtjJfxALLQvS7P6aS9gCibqAR8KugzmI9xw5ZmZkRaxo0egK+1TPL
FSVchOx1FCqMWj5GoM6WZ7AyGou97yEq/71yCr9VMs5b1bhdFUqQuw+bllTJQMtEuil7LzzABM0V
FxP+nS80s8K9mFbechQ2h69RDzhe3yW59Pa7StInpjg9LjN8QB5OmB8WCtdZCPGfPyepC7/tIrWh
62UrpVEUAvBVOiIGOIWkA0mLmqNEoJIDz0kfwWEyniOT2RX/Y9La9WRolQkD5hv6+nSunewMcsYX
NRNHmDU6rQaMsmPbjTOzQSgicXCtnVUQVc9815GXIvcY1v6OUHEkec3QxVmiZbCOS+VDbeDGlczm
OVU6Vibuethl+VVd8xxq2ipkdGMi/Yi+lWdO0KG3GFJe7KvOH9n5pHlyLmjP5b6KbmT+4O6e+9ke
XRt+mpuHH5P6SFk/YYL2nTOMLQRxEpU0v4N44DQwaIdGET+F/Okw058BooOrbBfydGBzdnjiWbIn
q4XDymxIEHDSJA7e3aXZongzPXTwpvHXLabzKAot02vs5Csd4dlCdFYtKAVGFDpz65zttQqSGOvs
y+KCYiDouoj/WYQZwFSzn9G73kyq/xRxqb1w8HDjwuYm7fGivgXj71pioo6euN9cMChQjDDyhJlD
dhhA9WNz/YUocOVihi7x0+Gntsy149PzX5Y3M3BIjkXZK/ttFYVgar58Gq+JBviQVCAXNTW1oX8q
j11k/JhcjSofDoOhVVl3bYwtOCD5VdTUt4DcRynCaGfrjHMnboMVwta+CopxbpuNQuqiBzzROilw
Y6iGxvPEZV8uTt6/PzyejScC0Mqrh+g5opnHdZlBEL/tJrLZzGsp+GqY4yGdAxmPDx7LBoLcZoVB
mEUheYcTCpPMZjxrpl5OSVdSOnhMq1pBGj3d93uX8ZguvvKEMhaU+ncdOajr/puhyZV2Ock9Esln
DXqCUpIHqwu+VGtqMKqsCbTydXA0JvFv50tM4nQFLv1iTg2m8NA/X8CtAjq7l2bMo8Gp+gnVsza4
PnZR2zSTGo2qpeEGY4iXOf4wXkTRuQTMFxlNtSlJ6Lx7PcaLb1bwBg0Vj6p4TiPe/fHI/anrTDPl
vJPPRcX1ebjFRM6q2i7o5xSaIWGOhpwhyqK5UfFwGuArbi+T3m3Y9mcyzCOAGnJOi83pMzxwkdmP
Q5bBPRb0Xg+suvilPOsxUqPKtIfhksjSX3tiSq3jfYnnOuK/d+bovtW6B3QCQgOu4tJ0p5P+elTT
9+tbo3dWBn8dButDUpY9bLsPx0MCoinFyPOJcl6yg0IlbNljceKbS2FDNAYI+e4JWJ366PZxFFQK
rQGEqRlRutvQvOiBj7+mLJ0dhl9TfGvvk6sgsIZROcq25OIPnFxG7jbb1Uqop2sb9alb/wUFBBnV
EYA5K8rAgtixNBUp/XPiNBUbutLyuyXGhSJ3AnpEl0PG9TSLZvQEW3FkrcDnfNkXR9XEGdLH1WI4
AP0ZKjPXUQNN/i5DRnyrXGymJ1HGkBFsv4GNceVolalGxzJF2as2bjbySlK6s/SFMKvtYS/JYqWY
0O9npoIms0WiFbm3tACRcC46z4G3j6sLsSETRjtEOWwYjpqRKxR2Ne+39+0Zl/bzH0VRkIiV4Uan
61iivplKoZ18FGZmAiPTSod1zcIxYhuBV4Vm3JksuxSPqa8rmB2JkYLZ4KrMKjfSzD13lahIdWiu
GmKYdNN9D8J2u8koeAKwKdCzeadQWIQ1MEhru8npLNVtrrpqtn/AQLkfv1VxpfUrViLYtH58E84S
fEalpyIvGYLhdqR/AJP5gMbonUSUPw9QpwiV6RVA0P9XqfvMQFm8lR5bZ9Hukm+FbQNiL/1nrHU8
v1RQDuOxUB3+y58WymVW95j+bEolXCM44EEC9K1k0IE0mMkWhbDw407yL6AxF6SVHPAeJQz7kA9c
JNtl17KpFT+91mPk+OyIwFnCJh3iQPHuPXVraAivbsFU0FlWE7p+5IpjdkpDFmLE0P8tRRCWbFNP
/qWanUVCf4/lbvoCZgA6YjuohOm9BrlmMwKKRSdK1sFNouzi+16OepyYWiRMgJ5XcZp3lukkhYL1
D/lUqk34YYECIqSdPBMc7NoO8iXA3CNeKrShjKVY1H+91oTXcS7HUldLv9Pf32rWBvotPtCQxXRl
rBn+uCHOlzjSrqDTHia571ZhQc/VpdxiXqUoAWKx5ETdLW15B8ps+94/ecfM9WaudsKIZJYvR4U8
eyt6xGMSQ8qzGNYQ3vGXHnNUfUrCHv1vluWgESFTr/4KIW54CccbgGYF329XoVTjiu5gqSLG+iBk
mgyA2deWeHIGO24eVJuKaSAqUhn9OY8+iZmxM2buzA0y3BtSX1lixgqXr8imKOaQuKmoBbfKaVNu
T6KhkpGAPnKnwCk1x4hc5b1IReC2tIOWTXd+2eMkEbPqoWE/V5JNM2q/cLLtck0NxqLaGyjvKgjq
dODPh2cMZ5l8vxo9NbPBPSLfIi6LN4wzu1D/R5xwY9rdfV3aKy92pNE38nF1T3sJF0R3RMgY4btd
nALNEaprRld445YE2BOy1bTfDwcVUaSYsdJuTE9QiKf+FFQ6Qal4KTracP3ErDmSeCrc+hChpNd9
9X9x3UEvQwV39Ji05I6MiLTNvn0xiXUeE+1Qt+8ivy7zI2svaTrkJek10CmJVsQET43agLhIqcxU
jX2XlCIloKfkd/A5VpJCS4DNYrNZUcZ7RGt0cToeWjvO8vH6ZjLzRRDAylh35KvUvlOAySSJeo7G
iMUEzsbJPmLBCWFWyBCot0lKbZpEs9hTEzbuOHZcCgvfmjQ7GbSI5lp5T/w6krZOqXb3+ngcyUJK
/d/HHPYQDHF8RYqntKuT1PriB6cVDbIHLfsMGQD9/elxB4btVh/lWTVx03cS4c6tDNQws2SDdk1u
Abh7FVfpwlCcrJdPhju7Uz+cXfKnvCZpseIFevyHJlUxGLGzZZLZEPug9X5/EWbBrpsI6/rjDpIt
EgHAiPa5WDLTB+LtZb/eSfySIPbwm9C9XGobd+WcsMGeZ4aSaCK6lkEbgL7eefSOWsGpWndAWw7J
nJTYRww+95ZOm+TU5kAS6z3qzmaFIOuQy9wU8ms3YlkeiYTFW4SrxGkx57B5D9+o4Nem1LmZPyR6
2ru1pZEngAIUCT55wdjl7bRlCeRA0r1Vxjl0fQ2rZ55Iwt0rkb7QPldLsI3RDEplsYAon0++ivG5
vgP0hfXR0qoPxQ/gAc2E0UBC3/Iq2UqEYCS8P1a4U7oqmNeqagnv3lVMM84Ruy2HHE1KhsMQ7sf9
W0/qIjqt1MHER0/aF+DmGhAHsp2zEo2VxkC5nkxTblC0r90Yw+h4P1iKdfLAzgoEBHeP1rulJLyw
j1HbuKq8QnCSSrYc12m7yEGEB7z5QJwoj5DajR4hwUPZhN0TYuyZHtvvdVV5siRJ3yxCaVWa5FoF
DBHo4zLahedtknCc+wtbfkQe7V5o3s17l+iFu2SwZwJELnDmHMyrzLcYohyb4QHYI7RSrL/XOlpB
EnhkBbyrEU1WW4BtXqG+uw31H2Gb4AUDUbGaV/Dbag8d6McKfLztHfPavmygADilv5YCVXw26jdF
f1yvMQ0kyIdilniKUprCFhD6AVkUdCAQWK1rypg8LafA32Z9nGqY83o8fgQiqs0o7DRNUDgGETj8
y6KA2/FA5zir+zjuFhU6WCzUN7YZYQ3y+Z/zkKIFi/q8N0pCShSXnhB6pKSHk1ulbaIZ7Dz72STa
sKD+A76BdZHYMeZQ3VUyl9bseEO9oDgC7Yvu38gwV5AbzXcLC5ZAaPrtBXh9iFDl7R5SXTxfgwvB
yWtyQhUX/OEO160h8da4xeVRkZCk8BVt5LxiIDNlB1+xJopBKWOFot0QNeVzq3IgaSxkINSuLufY
HerG5dJGb6oNuUNYYWW7ViZrQCva4tIhf8Ntu1GzJo2DGCU6tnkmksv7gEi0uelSUlcECoph+I93
Mh30z5Frt/om2DjZSn+RoPqC08QhKDYVJayiJVjgbzT83Qb9BUG+lvyNmyBmgoyqpsYpDtK6A4QH
LB0LwpWPQETJ1+/Y97GNWpqfO2VbLUQ7pGouniYggQA/k+HZm+Fu90XiYj31xjp8NkXDtj+xmCNn
hKCjdSOTlAzzJ3b+3I6OpGVmmwajru4vo/nKW+hr5wRrWM16dYVMEt/MwiFNCIepZQxN1i6r/IiJ
v6KoLROPjQIRbt2AVY/bvK2FaVToVfqUuUooIQTOZpYOZz1VXcZPAAl2+Qlj2nF9baFVdVTb5luH
Ye3PAgeEwgeilaB6lw/+9DycGyyXHYq58s+QoUiU9VbSTjTqiNy/oro1jYPZLTzg4uAowuuC6Pi9
ICJ0VORbly4bqkeeiN2uiRfAm3++lcB73vYg/dRIzguFelXrPFSLBheePzUbiV5T4uzKPFwOSLn6
4e0sxRsL3l9KVRyiWuLw6gbXzXPa2vIcTvvHRS1Rq+17hJvq/DXGzIrJ9jioK4PvTvEOz4aB50Pf
g8tn8XeBrNnMve+Ngk60lWg4YRuX/PFBi6lgO+Av7IgxtsgJEp82I2GEKQIEIUFko31sjMqnfvIX
WOwinAdQISn/tqMsZ0ODQkd/DNECFHWRtPeSO7Z83oQyzRT6dUUJ8ZXSTMw8xeLqAaG1DizIoEZh
Vgn4J7XY4nHQJKxT9CfGa9tCgcWJ4i0eOuby5tTS347thf2kv/xYo8MpplS97/NKxRvZx5C1Oi1p
pdwLMXGWGVqcqvmqa4dhUjEGjT/Vi54jweB6RJBVia1WfvOo/X67cjSBXXd/+zG7/VP+T30DppLD
sfWXIqx+t1/gdcfP96FHYnsyFotd+jshDU94ZyBNpTV4VL+uDnHiz41PgZg/WCLAUswNlvQut9Bl
gtr6F44hSM22leQ8du4PXtBdzRjP+FcbxsPeUX0rgGKFIOkTsbU5y/slRuecKZcipBYtdr0hlB4b
bBe59T9xthG9oKLCBb9IcUfenv0TZFmt6n9OPx39Zu0bVY27Xq/7WXVeaSeYGJUoGVVdvKxBh6Vc
BOLNdS2q+Cg0RcJmQmZByQdo2XDRwYpx0kg9xWPYQIOry8oDLGIIgRshLcAtvA+qbPo7+jXBxsh+
E3gK5+s9GuJS3eHXlpIzfjktdmEM34L9xSJWFnqopYzizIKsHzfQXmp5rXZFGECoYIJG206MnnNG
G6/uDOe5ZEOHmbs/bVKJGaSX02+e+VRFA+aCoKida88f4Pmj3HKfZOIY1zsfumbue5RMd/C4ZQd/
vHeuOcn4nRUon5M/F6ca93PgIKCgDYHFMHl2hk45ue+aWwaafy8ZV6TLsCoChtUV699M0uQdLV4T
UwgVTwNpMM1uyPM9r83K0fJKpzwxvztci+pb1WJHOuF4m6atYEs9tIdnxVH/6pBEg+wLs3utB1Cl
2RNTX94VVolGjRKZVehxw3TU/qS5lAqzDmaDanhFt5Gx4ZMTeFrfdnoZ9/9XeXNBYVk9C22+OL6H
LJPM1Cy2DpYq9VZi680VASQd/p/3dlNKBGx0OEd88Wsu9d5YnemgT8ClbsdweV/XStTusxjCNb0L
lFyYVWkRIDuRHoKTwPmqSLfTOTWe93MC3tCsuC9S2Xy4QKxARE9vU3nvO+uo2GPxGUNlo8nGOV2y
ahfH0nZB14AYm4p62I2kUSHFibDMgTDxEW3N/jAFK7GwRpXLmimg4iqn8te97dVAbHQ79WlPJMJL
zPDaDpr01RuDhFFgi1W8bpUXRTDcT/+1+1j/M3Y7n23/Q3dijYjPnVFebSWYPdxg99qG/OyH5jtS
+yPZ22aAxzft+kqrJW6XrBCBxVk/qntoIbRPVuDv3DQF4ekvApXzi9pv+raz11rfggl68LQE7FYQ
88ui6cL9sdcrTPHJBp50ujuRLtXK3gBjtIAdZSIN0mZ+HpPPQTFbap4wjB/vHZ/q8d7g6rbl4UK2
3LFgKTVryUAWgbwkKmqdIUiR/kaA4sBa8U7kt5RzptfJOa6ndr20dQekKZqxiyWf1UHiOkELkTU+
TEACdfwY9Hk5w26zWW4KUwEJXeMLGfLIl3CGU2UuXu8RaoQr1A5BidjmvDpppeNVhxmdZXb2yjik
uBqfwHopoETyhzzalL0jb4+YCKLKaYNxaOJbaVMbpLzAqn1kRASaaS1tDcJ8eRwqXejG5FoNICiE
lOFudlzMOSIBuzLwOqOxxPLS19CuHv3RSIFfHjJmu81d2/orq8mt45cH/Ze/OY/Dd52Vjjp/5TN/
wF8kORbxcOXoqGoJ4vxxnVsbQFVY3imxzlnp89C9RgO08xAWDokRFrBOckhHfCLVdTd+yISL7kId
F137dEHKXh1LPKroKpYe5owwaHHQKt6tOkYqzchndv1gFs8AOTpf2MkwXSRX8e5IuLalk7FDCIip
Q5wzm/zKnYQbqtXD10pBx08cInLZSblER5BEmtN/Neep33BoL6U8Yjv+PrOINmI3tuU8Vd7p6Afv
w8QNPoy6nYHuNi178j+o5X7C/0hR/iQFyl3so2QW2Epo82Azm8rRXh9o7QY5Hse66nV/6zInv//k
hRaBO8j35SCxDjAhTktHW+8jf5TZHB5vBpkXOcfS5fI/Z/SaSAVmD1FGTAlmEZMW/xF1H9hUV238
dsdFDmAcFqCm16k6Ua9/NvVlmRhdCUYgiKL111NhxrTh2J+1gQDkFBYSM1ke9Zf/enZrJtCQhHMT
/DmqgqNyRqF3Mt70/wbUE1nEUsDnZKt4tv1YMCkzrjp4+dEfGCca6DM8BbunbqeSGhOqLvNQfAjS
P/Mgqx3WUHLxf90/pd4z7Y0Qivbe+G2AseidNabg0FIaicsDYXbotuqh6WpwGB247gGu0ei2oNRp
R6r9uOJLOgM/GSu+lfno7TaeL390On04wNLtNfaBZOtGTAB4sTtSd+fwio5s5ll341CGfPazabrJ
JvJxXulURS1gr25MB03O4oWnPLcZPa78roODIpNEwaxpAEQVT4TaWJ9iVijhmt/160BNgfkn7nax
xSCVoOwkWzSW9JlNFIpZXp9xy2iWUpKTZX7oCTgatagMBWpJGNs7k+9xnNpNzGna8g/d4RWuSVix
V7DPiWAmPHNdj9oQqVGSqrcCuvc7y0UNz/CHkyJymH6sMtbopyQFcSrRqQZ6MVmbWWvSkw0y/xW9
1DuvbAot7J57MYKGFskG1YsD4bav6GklPH7Od2mTETNd4SXBteZ4sVgnbqyxPp2RsVJuEGq7eAjU
FbFY+D5RZwP3lIdC8BMV1fY8317YUiC6tswnvvuYN2D8cvBJDZnVz38OZIx5m8GF2ta9KfZHXLzN
pq9fU1wB0LjghJxbc9QNAYRqnWgpRbVftmpCrBvXMG5JCY72EX7DGVcRMNfkJ1szGQe1A2I4zmY5
zIlSWvCNsDK8ALG584uIpo2Zbjtbe9EG1bMrX5vP3gvzC/uPbbQsXXKgDH71h1wvYpuGRRcvMV74
df03fjgPluyq8iCEnsLW1CasIm9lupfsoG6gtokkI+hvNslab3eupZkKEukFJCLscG2qwggg4btK
VmD5FVK2mYUQHkzNiPhpj5u1ny0NEPugLwkKcXupPr4cTOLeOzPjV0J0KRxr3H04EXA7D9fCekZT
c2tzMnAWAlGrGo6URjKfeCt+HY5hPz8A/t2ejVdjpjXwoRLvXvAjfxphFANpSBSKVjv0eL1tNNIA
Qcc6fZIhv3ttucgZ8ynyyXH+mTsDGh1c7+3EvNkQ8r7P7k0zy4UMAR6qZYLbxy8bKy1KSYtohHIw
7bctgijh44mIZbywkyyNUwgRFydB9jD6XJZ6TsACNBtGNMD1yQpS/ukQPe4phQ8fV90txsyYfIK/
I8eUxLKkzSr9/b6KR13g3TApIa94x5Lb4Jg3r6ra9WAMFs6JBji6922J6/yrwgEyr/iwCr3iu7XQ
sjR8jAopwWb3XyXlaazA8viuhjnhCgM8Ezb09D+XDe3MqkV/bKE1+CvkB3wKlNjNcx2e9G1Oa9ep
QqPbr2ediQuK2CaIv+4m/ZZcc2heJyqvKzWJggOzssYuO8LrlVYRiN3KfNju1SiTYS5bBD6Im5RH
ZNvgdThzJGQEC1ZR5hdW+7ix/DLTaawZBy0k/lXwjGsc9/6VNcUGcdmyPIq+tomBOoqFsQTzTzGh
fsOy3TUoCrgDSFnhysEgqyQ9cyDLY8XSMx6/uJ1Ir3XX3BouvWvY39xFeOH+dgigfvnLn4CtXNdj
Qz4TGjqZfvW97V7uTJGOhqUe6icKvBz1EMEIE58JzLeJZylYTZNARYQPsH5JXL0Is8dNrMyHYTbA
KTFwEgMNRY0YfmwtcuIMhKSSY82MSxfbcMUTBGoQ9gD++D3JdFs8RYDomYCQnk+dvhSe8T0eas18
oe/QkyVHYTKHcUUq4H5GlTFZw8ATivtQec6ecDopHL3/IYHM1SLQzx8D0ZXZ5aEtC2NPu6nxR3jr
4MN24DArNWk02GgYN5FGmWUUX+K5Wd6iQ+fJTpjCtBItbM/tBie0SJAFkQC6NC3KfFZyBLHZ+j1d
JOzY4FF/TI3k8HuKmpGEit0fcC5doko3IWUvP0BTP1MkLof3I1eA2qeNcVql5nLiTw6aDeo9tl4k
9fVX0AAsDjQ8EGdU8sWCfQo8VuTQGOYgozKATGubCk+jT5Z+hTss2efM8AoL0Hxw/hqWq5prmnrU
334u2mD2trbsMZma8UB7+bdVZgk0Y1o+qQQYoPKHZJbbECycFn6IZE8CHX7YTdJN4KwHBTWmK3RX
n1ZS/62DgjsSPCjdysRrrWfs/xdh31bqMEhFAxDYz+ei6nF/GZEx2t7FJYsUZXwdCJdBq9L1t+d/
xJVR7Jg8Pwa/MAlyz2DHiin2BlIyAztFJgmFqtJMR6RVRadRK8v+9JhtS9iElT0QvyR9f+E9MO7W
z9FQF3tcumsmptWWcmQ3BS/3rzh4n/ib1UoEafVeUYXjG9+WdtWVXTBhil4JnAsqClOFXL60std6
Ri6NhWsIqyv6j1SlTWZh41sM3dQh+eVFeZkMxlCJ2cFZJ7dzTZJSBUwdMX2Hr+1nOjLDU/mfQoBb
FQpB6adUvQ0wCkPp1t3YRRFpAoUQffO7CW9K12Jv5MPIDn/SkGLE3pKxBdyAWicEBiFFVylMIlP7
otMYX7ExhwiEBrrcta6uZEhbKmlHraUCh0ilmv1Yk00iCjL6R+Xws44D+WGwHvTha2VE/eulpLQD
ZJh9vYmzaN7GdMUnr7eHViU42qSpyBkIk2TthmdVrB2t1q9ZdNfPNMLoTyBHED/8/p1kMQniVM4t
8NtSKXcvzocitYgtoc8RwDJR7MRFjUS3n8meeH+97bx+368Xalxd60aAyGFMrJISPHNictOL17CC
Vd9O8LdnoyxNECwIR07+HaLT5krgeiawFSuaunWlXe0NB9wIdxPdgUV5ZX6unSae1gWT1U/0d9EJ
xgjaWaoOMv7o7rPAAhemPMG2CF3kiEIsXajS7ni9GExudm7vI/PGVtQCUI/l5VBRYZJVbqg0GAYK
ZFnAQ5PUy1Hkw6n67FYtQ+0yMJK70Wlkdd5Vp5Q5FWMUGnXc89eeO1udAhHXFUhcTMSNmNrSAwuz
4AvuGdROQY9SqQjgrR2z8SUk926IPm3Zr70o1lYST3f8rUACCk6jJL04msmV6/k3/kYp28w0BvU9
BFmiGnCusjPnvLce8IF5cD+41b0ZZyOZeXzNrhSrPHGwo3ehmLoAZSf1xBdyKW79pMISsWS7ytR4
3zsIJBDvNGB/FKTHiM5QnDv+qh8EiOk294F+JYwpKD+NVfkj+IoR2HuBYJvfsa4Hyz0vanEFZ0mg
aVgJitlB6qArOBABYzMukpsvccoV/AiyVcdp3HPuUCHTBppW4yGDijgaV6kgYjpNJcP91XzmXWPN
ZhAKg29/+jkNbXCCoNEDRTKknGEDZMhw4ob0UEbnFYq9GQZmtZ8Ko/llEkFfs3YIiKc+UyIoqyV+
Sqxg9IZ08iA9SvbsvwU1medv56M9yOjvGk3tg2VUb4iUbUTFEdfQvaU/4K1y8gFBzWEO3VzDVG4g
4t3FdDLkh8tpYPh1/LARi8O3fspdq8VX6nZUpYEtJxWuc1TcE3x8OnrFSNGF5hKYoepKqCahVPtE
VRIkkYf/ImogBKOUtO0/aqeYYaoO+g9jXf/+nSIkts5q4JKueoNa0wUlgLyabdnTQB42slB0CgZd
zmES1MSgESYjX9z++8KV6+x77JNHQNkiOOWTCxd/V9XHR4lOItUSHOHQy1a0yHkKkTDp6JPZ2BiV
FK6GhDjL/uHGeU8G4zUTap4fcJWaXL6cMbfyC+31JkPqtyfNWZGjdtwn4dXVbuShYAqfyuuFN171
h0TnPAVy4TZSJiBZLOuMzd1+XVgAJ9sWkQ7i6RrZ8O/SgkNtMW0aLNsUIRjm4yVB1rJartwSCqKw
uD/kTXGrSennfsekZDZNOMVZi+6Z7ElxiTthXPr87gqi3+EmyKsaUG1FhRH29kOdRL6zwOExlR0F
Enh1Keyy6gproZa3QWe5WB5npaN1bK85uM6VkF9aNt/lxfqaB2WMK3JdRNIn1iY023/mRLrqzSiW
TPn7Fiwiv/EBgceDbBVg60l3SjZnB2qdA4KvgbSpVmXQ9nTEgJbmG/rlSRH91I48zz0l9zDkXwwx
QnmUNzvjZf6OeooCVTAO4BhH15Nxb+AID98k1eLcVBXq/+CbrCa3U8NFgcLB5/1BOdhfVOezKi8j
SET/3E8cfRSlnf4RF5aEAZ4oQh+GCFfKJqmdzv4L4JLVp/em7yQgPJvzeYXneTw7YU+5F0yVzpRB
krwynOuBvZ7hgR2nGoIeJZLBqF8WRwjPuhrjIXIz21q2gcafK625dHl5JzFUVs703kBwHQOepOan
6enU67O3kWjcEYB63usUV0KjbRiH0EHq8UAnbynkqI2pbWiuAiB8/BxXWDBKj1SltZkEr+4n+bbg
zdChdoLP1CURFUliyUdtcP6g9bHJfV6iw4WjX6CNqyrU7xWqKSUSP0k/Ar+rGp2SJwZK6z34ScDV
qY6BY7VxfqqscpXKAge7i20ulhrC57SvfAsWlD7MJ0iKJ9gZ2h29Y5tyfeKF1ImVs3upcY5kAWpL
NCiixzTlDg+36GKD2P8OZsw69cgiDlMLzjER0DrrPimnFFvxd818qy2Y21Ky4maPpoEAWSBhSpj6
VjXRq+uCV+EzSICeB6cWWYDfW9bFrDVhpt5+0OLjbvVwXNHW2zHr/9WtIEYDidcnSNumwUJm+dz6
5RwbLPOXqU04/tEz65tz9CfQnB7VbVwuxIo/zcwOj6MmlJ/Bml5+gVSC7iU+PLBwFrV1q2VdaJ08
fj6YdaW5qLCMpSAE3DovW3rVecbv+566hmvC362iK8o+GGNBBd2c+tssz/i3nwxDVJ2Flb4e27M9
zwfernYMeJTOxGOa0a4KMUVWrHZpz5prNPz5xDdU34f6C06us6NCIU2iQLlS+LlJl8Qf7HlJDF/x
5DwQX6UZylByF0MPcVA5Z0trBvmpVPVOntcTMAxSWL9ZIDYti/qNFdBPMKKASPJq1msSVKmwKIhd
eAGOHPmqbTXo5vuAeGnCXXvCzphcmPwAWn3OAhz/5aTLWdg162cwZrRtsKaYurYhPQu7pX+cTiHH
mwF+yGJpLnF5jOzZFd9CrCQGe2GfcgCO8PHrGCm0NU4M2oZO9yf4n9G1PNb/ZzdM6PxIbnk7UfGg
leab5VTwz8MglsoGzQMNX+RV9i5TLAWXJ99Y4EaroHemQfjGITlXW1Fizb4DD9ttsg9jml3sLyMe
qfnyuXyoXqlCY/oRfnJEVNaZqS42xFnXBcw9RpamcqbNKD+fV/mVnfdOkE8/iWxDty+hEw9ncf07
VMoEzlooQLZYcho967RJUUGFrmGQnHXn0nNQJtQWgb4cdQ9vqzOLWnoQGeX9oZyKplTzdPLPKON1
nDtXGOOaBTScewP1HiwIZZotY22zPuCDMJtg8EIQQaWWk5qjeHMYPVg7IOozt0z4izcAuj+rU7hY
oPlMkbHRoXo4RDL8KKIwRZSFUj3lSyq6aYJx2hXOM4Nux01MxGZt8xsDEKgA2ZvQ5oQyU+01/6Qy
bSQVslgbl73AyEbB233G9AUl17VETdqRAMtKpMnMUvNo7fAdn18SL9N1BACYx3CIbnmWenVDDWcz
wMRYpMZvW/Sy66m59eHOmsEDnpDtXjl1qM55JkiXT5OfFKcOYvgSvGqNtmLz2lqTz2urXz+31IT1
dFwI+OuMGHueBZIM47i8HQMjbCuKqTABfVrVU+RIfz1EwU8dH7yvtaistZpfXmWze+xh/l33QXUm
h407/L4JgamegGkYyq+8FTClzz+t2rTA+s8QO0R5dfkNLvBBM+kbDpdB4Gjg7rCNvNyvc79kOLPP
poz7Jk8OigqC6118Yk5iOcYUegstBpFYLGs7WmPIn3Dsake/8CzstRKRiLcyePt72KQ70aeJx3Sb
ycgYOb+JtYIvyNbff5hAQ9il+8Y0TbAs9qjE28uGQkRVE7j3ZLUa/ccK59bY0VdXS3bwe7uLIHsD
SoFk/WJ2arJQBNIXnlEnaD6cCIaoxzeAlNOV3g7RKQVzH4gIEyN3zOuljzVe4bdd+G8y/P3O6UMa
SUKxLes37BIAGJg3Bka6G25ZBB2hoQnDY99fGXJ5kBVGJDEvqrqq5t5uyRka+56nahKZ6MBBS6ac
GdfMeUS/G4aV/zeCl89JugWEcEYN7PPbom3mJuanGFYYlhvzD2CwrUJ1+KfRMSLBpLlMrUcbm6Lf
ZT43M8r7f8OPw62Ont/qhJGr2chKquu7zOgAZI2KHwhwVPNwRHNqY4lhMjaiN1Shx3Osaukhliur
zMWUSkfVRSP89OwfmXF7sdt9lHqBuoPByX7zTnxELOu791vHb/Yly/i6vxetVNDf3fZxcbOy5jyu
+8KQUld5Hno9wBTBO2fWgnGROYP4Dt6/XjNSs3prtFFGsUT3aIAlNBK8lhi6nuNY/6U6+zXe4cR5
mzH+YQNDf1lfwA4nre7dFcZd130LikBTbm8tjp+vXvq1WaqcKc9VB1P1uIQ3rSEPBFCMqosHc36C
jgNBqYBiUCQVBIkAlxYPEjCyXV3Y/Z9fK/9HVe2nJJo8Y06Q73iSq6nHlpHCZf9E6d4uXJukjomR
nTFul5yXO1N7X1XrxWbK561pIv2q41V4xV34tCvY7v+ryvai7ir+PlVlJy2CxYWjFrtFdznAuEgb
Yj0ZdgNc0mWd7h1WAE6bPCutSHYNQYXsjAs2PFjc0hTpFpFfPL1jrhfFRLOvjCjlFiaDho4kmcH7
fv9MjB3+1UJPaMp0fD7w4SOGmqeUqjPAlNXTAfWRQLeKBEXknwOkIOfq7Ct2n9qnrdExAqTyhbeb
ne7crvEXpcabPE8Lw0SAKoj4F1FreB4CR4P1btQK07cN4a+/Zjxhk4foEsqFULFMwgWwdoJmRiCB
jzbUuKRCijN+MLm1w+GvT0SJwbLF2oAdoB4oHWaJuuCzPuAnZmZJoAO+cyf2JHnsURIKZ2vml7GK
OePncMNLjIpE9skcIM2QY/eaBP0oTwInwOfMW66oL8L3IrSdv5DLVkYZK8PV+viMc6jYefW1HnrE
9TDPaTxHUaYe4S+hMFOZRoybSgBTZtItwfluCgXB7YPo1MAeu0Jno8XybOo2g/9A22gw8UI7e9D6
QDsETgV4kpXoFnew70rMbzraYMGn8hpARlytESYZ+2jJ/81vsTqU0RNdy7TZOH+Vf9ot5D5CXvpF
JhVSFwe8tN1GCYKeUIM3BDaRYkueXZHB1Z1EaGySb/g23bSGe7RIJFaL6ak9MT14uwhQSsWEXq42
33oJgZEs/dCUoqUIWDXYwobHOD0B3dO+mI8mqRz5mu2qcHOo4VO8qLFJS8GSvKpyw9R6VpBCyZ2Q
Ahy/qmMtG+voD65t8yT5vkhRTa5mexsLAb5927nlGYbuhshbAEknu6hDm1N3S0lLxTURoCXtQ6qc
gPvWOYHZANDcchFOl0VJWMCuchTmXvp76vwrrekEzsgKzGpvd5Dfgdtc5eGEOFEgTE6+D19FdoKM
dHx8xzqa6T9rclLhN+ELQIm+m+rzOwWVKT14E+fnMOWu4IjGICdDdq4tmkmRU7mKHfZ5n04FZp4l
GCjguBB8cXa87j8rx9cAo30D0J2hzmSfsgwFDhtY3ny7c/0F1fULsb/g1bdA/wuzvPOnAJKfiFRi
9Om2wTC2o5EyFdixOVk2vPMRLxsl1S4DCg1Pm/G45Z8Z8AvZXliCazPEhlA+5N5cu27Hs1hCn8y+
iEeH1yRHo4qc9nb32VtJzcBYpLthna6eJVzcs0pd0aax3lZb/GY+1OiYNQQrG9RhGfPqDnhAXx6c
jDMHVkGYQMe2J3vvCysQKkrZ3qz8xNyw4rM10/vG1yDpo08tkBMvMhIuDudaeYFsmNWaL0f4rncV
1j6j4UGJAsh/7RWhgmx5gudruADhksOUpesIXFReoi4KCeUZ+BTrTbgnlO3Gk8SL+f6AAlHIWNue
0KJVo7UYnXN/Cawmy5vCGI+RKd8oNd+ktqrDOS6LrdwRY0r7FLA6Uchu4T0NvQomBZaE9seGW1hr
ErJmVtTSaKutDGtSLQbDE89iq5XHZ5rDYPqoQYHN51cVhMj07CQosUA7ECuQQG+XLcHLt9uYwOI9
+3XX99BmcHXnK6ZJtJcuwVxsl6dj4wJYkH8HAJAxBC3+28HYCcLT0PGD+1F+khlxYBQtfLiOwff9
agdJPC0wzYvctbZzF5vLrAG4cdKY7bSgboxDTHiQv/G5mUGffE0YP/hg5VBu2/HuP+OlrRNTDWAT
R9HgJ1o/XxJvQ6K4ABmI2R4E4Tt76KPBbV09tT4+xrPhZzIMGv+0Qhn86wzgKeGoBKP91DAIqyU4
5DpraPFoFU5x+FOySJV92DKIJCkxFqqyB2nDTrxzaviZv4pg3TiyFpmKN4hijh+hSk1t6h5KYIuw
OVgFaShXqrbjfFddctwFyJEG77eSirGxl0J7V5VtIRv/MY55EE20SVB5H55wtJYpxqD55YFPypJD
8OkB+RkP/yTZl8qMLG4hgjEAA1RKhmflN4K4i1BXXknGxPnQ7M8ISCJh3mt324DZPZZo0VwiRerE
vZ2e9ZFz5Hn2+7I+qqr29f77X6Iq0iO9bVkrb87hgna8MIZe6yUh716K9M8p74OIy8L9gBxnE2bf
mvmSf8Beoukp3GbZ+ka+f4n/cAG0DUcWCqxbiuDCbC3nJ5lLv6sjIr5g34JOfta7lUuwT0cz1Scd
SqIumT6Z7bGJ/OojxNL4GDFyE3u14mElHHF22qbw4aEWt4z0IgpgOqv/ZV6sOMUl4SmcHncYzCEs
+2Zv+h/uMyBmS7i84Qfa46ND+l983/s2y9X2DK8PibbXxNBShagf0Tn5+/CaOJZhqbkapmEfp7Lu
2oU9akj+fJHOBFBBHfUbfALAun0kxQflZa4mO7KatPV5wQAB7Q0Dwbj9oqWHpZTdRgVkMTp5/Z7k
8s2rPvTLHF8MPmi6B8UxxJ8QNANOJVATfomGqux/YZ1mH+Ig037C3iS30BJvAXUbhPus95xAU5qq
AJ1PPknKey6aLqQRBGvpeGVirX7xQKYE1KlTs5tniycUKY/85MCPN8fweaGCwokxKIDQo7/oN929
SORgfLv5fvKCM3NwxCtIOdnel4Ii2fuFq29NuWUeUUKQ9lBI8Gbv8z+pK/kOWCdMnDWj+kPeHqgg
zM5CRaK7CXYDo2f9XzvXprFUdgCAJEAE8+DJ9ZXooQc/GpUyD07vHteKUKATot9WV0svOpRsx2Tp
+JnjQRNsDE5Gc2Lja8Ghuq92liBXmIK+nQsRgY61vxakNCWz+Dc86tLjejGgZFlemtYJRl9jBhuy
tRy8qM5KpKnZzihlC0omyEWBEehPczRNC5kbquHniTvgwqTTPsITGrTXPdxU7nBO2bqatU0cllXW
CzLBgEMg70tnv0dCvgFdka6yO341zTwjWaiUGfjalw5XjsdkYGnGL3AhMZWVCg9PLrj0SzM2N5Vd
FP5sOXEueMu9DWabfVwOGCZqiSpaCTKPHis9mwaNUhicBGMaXoUw81Wnx/If1LztIGtqFGU4GV4S
R93WNgDVZIHh2JfgZfG+0WQUsELzv1ih7F5xo9D/Crf/bolZOXpEEWMexOzOBrsq1UO8dylLjzPC
o8TNtnrtOaSd6psBRHyHEI0WM1skS+g15040hO7JgG5h45XduphmxPfqUqxZCBSBbOTvYKnEK1k5
7FmgytuB73RFY2xaEZDeUFTrAUxSAQig1H+L8C/aoQE9K4hQjbN8lMM0RgRPDrIlossDPdAukAR2
YqVEfxhJUmw8YG8VQR2tURPsifcyFjF5k4DtD2CsQTKqa42rv/nduzqN2a5rwwTBs2DdlUSq8Zd4
Kp4wo3eJd5ARUdNatENr7yQN3dlODIvC6lTL4A14KVh+knA6+ZMS52cmtO2SvKnW8wOAPaQenZ6k
1YCyJcXBcykLM/5G8eRMCevzozlQuBUMBX1OCBw4otJhZ5sHMNNLjnbsl+LMYGRpQ6MM5FhGaIKM
XiRqnFZagoB1PvYKwe8v92vo70JhkUUevWbLS+qupXcBdkUYZ+U7svcxrIK6nX2Hdgh9eqaJEcCe
iSsCaNU3N8iCIsCc8Z5/SXnEdPNwd9kg6TLvvqN7Cvnriqsoy1ZwZ8NZXPRR4Hjb9KpFw9sM1qCV
fVnTy2o5i8OxRVK+LvOkHJoNnMNCD6MKX2ZeQHs8ksrWOeqOdiE16hD7Qx2cdd2pXFEvzg6Q4Q5r
cYxkqHrOwnGZ4jJ9v1M1YpTBEFOsVSBCCQo16XZky89g6yUoRlk6qyqJOG5hdHnYwbY2UOPVJftq
/1GLq/iFBug/Q19UywcZkae+z2+EuQGwD/S68b3pUIFuEM4L9xaZrhS+sBndc+yBxeLDxlKGK5GF
AFL2Pv5dT4kfQvHjynpP8QVtcHUItoIcn3WK9bHQbYHYfa083lBvVF9AasUW7JNwSmrIQVjoBejW
fqZqzex/afxuZs9rXrc7vSZzUWljx/frhlg7o7s3fYSBAVA9AHU/Xxdro49tZTQdx8BXjojbnOqx
PvrPBm9CmRdyLsuuDLbPhljmlBZhFbBnfQi5p0hgEEsr61rktISOiEuFpw8GuFO+SOp2LYGndsTf
bu6jH4E1riELQI1V8DNfyXDhFCMH8TucpXSeokZM4Plejf7NX9BlUrGLe6VELML7RwRl207Fd3XJ
20TaRpp7JH1ie64c979bwnUiOII2Mjum4jiEwfwNHiCusCWso/3VS7RrD+17TYVeSYlBT4MYQPCq
UMum9CX5EZI/uxBeXW5Qk/+6EJgXOaPaphD5GfuoN4huKDKpCWi4OsIr47CXCVgpNMZ85Y/R/nLt
WBSvw97NDn6UWXTBKeG5LXJaGggA7mAIzz/nzZlqc/poM+VQ+N3qQrNPgmywWwUcYXwpt20Qn+Tr
Q7V6TSrAEoE0elsOAk7kHKeCLLusTK9G7FZNK+FIiQXfUw9oLDC7BHduvfOd2zNDhGVlDbpsKdVo
Sex0vLY7f8L1dslXtsChfP84yrRBs4UHxKw3xKRWkdCO7PiGfQoA30n3RD57t+d8qRL/x5v7Tdsz
Xq1r+0/mVJPHEWtZ7X5btGAzY6xbvHmxEpVa1Cd7XMWxE3Crk6woLoRHkhc6FWsrEM2DkDcUAygQ
ONszfp/WyWcyYgf7C79CQUi7sePfdd+eZvCsZTtBl6iANYBm/f9/c+lsohesLkwKyLOzVA4eFqIt
YH2sqj66jsm/CFnnxCgTUFeqaXNBPOqhu3zKud4Hv8yPAIqzFJpXBiGuEQyYM71fOcaa7HmBKwfq
5GFN13YslCWh3oO9vlaz+sAW7EaBTRI9ZSseBSJ+hImAqVlDV3cGKdwvDlvkS3Y0xy753zdv5WuU
z7RMulEVj8SB6DDIC2yUUzcE5hI1h82CLEKrMVKENH56NZAClpm86TXskXLe/oHVWHl+kAaHBWYX
4sXHJ1Gh/DEUoWmvYaUWGOTQfvxPpS5RmXgdI0oDt/eBmD3AAAgO0terB+LJ4phDpJGrC6a5oPK8
Flc2cs3XMwdSbz3aWY5lEtCAAH8m7cQi8Z+fEd/m89OEcbiV0YDqUAW3gAmoOA89WPdTI7bOB6YY
lWGz0J3im1h42MOOCHb+srnnvLU6clYkU/35d2I39fuw0z5x0xfN75ycLfKrjbKD28w5W42opTOm
eF//ifH9oc0aZA7xpsxuV/TmyZXXcyf4e7kTq92+BIn0YJwPgrjzbOFIP2vKz/mBCuUPzV9H4C4D
4CgYWHZ9HIkXrME+MKPp8w/hHPPSDzMBWBtA6or9KRjDut7ychhCIMUySSf5Z3p80rfS4NJLoTB7
hTtFORSc+55GFUKH07NUQnvfC9wD9rq++tveghW0SD6+KKTeyXBmFzed/v+gO2l8fiC/4CfvvE5g
6DW/zaa4gre8n8Uf189yhPMMgmtWtQrSTfYdw/yd18HnZok46UfRIODIedJ2WpmLd8EQ+TZ4DODl
+dkFqBPJmvh+GAG32QE6sqBZJVEu25p1baTkFt1yF5Q9IH095HUi+0CpiRLoQUjPmI+ucdSxHCtn
T7MsSLrnDXn3lBzM5wWF5ujnxMqdss15ElMSey52iXgbbDBqAcPQq28kFClsCzF+1lfTVD+8FyHV
4qSLNqqldyDT+YjI/CtsSfJTL1B22w3YSXH0jPhUPbRlFXUoe//cngVqitS/bvqNnY75+dvNjjY5
CcARCtRUdPRZ2jFjD9/qyRCAoZ0/F7Ywao6IAeOvkwrbtTR7HP9SMb42r/gRkAI4hgaHnx888Uod
oaLNvfs6l4K2qp9sYwqk05fQTiuA5Ib5y4Nhf38tI44nPqExOMmyX8bkCWXq7waDN8cpk35O3Ltb
G0EiVDEtefXhA/vuLiHF8fFw3LW0O/iB2XKsFXVr3AsTVlI1DnJu5rW1bq7Kfst8g2ByzwGfiK0S
b75lgvBiL3EIvultCaQ2uSyMwtgWKywhoRKxiBG8aYpc+uKl8UDuDN2bYb2LBdjT++EDjZNxKIqX
Px+1LCTlC9dhZILUTN9XzUwYzQPuY5fhELvMokDVRedFYYgY6HUFaKcfDC2AQEGuu6wZyp2nbkM/
cjGXnb+DYFsE5c+iop+IPYatIkgL3uBnjiLRs+eQYz1CUUDt5vd/XF5E3tbD3ia/VT2pi6rzVWpx
mqAB+FK4eLc3PFxfXOu80k93Z9YLpdgbWcZ1dT6+gUf2hF5POH0Fw9eWBvUY99+OCTLTLFCI2fIU
UeRseJhYVnR7PH3Bol3OM3tO5K01aCuIAiH2/j5kfRlHOodYDUfQKVWLcfRNrGVOFelSF0iM6Yge
m7wNdeBbqQHMU9vu/5+BcoZtwpXf8qUDVXar6fQ=
`protect end_protected
