`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 288832)
`protect data_block
0eB40Voek3XE4QOCP93RnVPhUSFs7gsuZImk0NukmPcoVsXmJhe+9mR0Rh/ZKFkpRupwtPjB+wzq
+iq+QETzGXL/kNGqH9zYkK6pKHrLQqb4XRrIGrPis+mpo0dqIE9Uoct8g8HMTYvEszQQYEBNSgT5
ECf8EDTqrvTtYzBQDOt07EYU7jAtbQ95YspE/r9Afm03a2xP2pXV7xxY2fc7HS0yQGPuLogLx3Ww
XJO5PXp5GN+92vBgC/Y3C1MR+jAR7rQV5XtMaUkd1IkO6sfmj1wyu+QI6d+5z9SSzPev+WuxYUmZ
LqdQOKGEmCnjdp8s6IBITYXjdHBcg57EeRNikeW7qehthYUd4Ur/ia26kwBeZsW+ubMMewcl4e54
UmEzsfnGusrWnRU1yFlYOnFo1pWsZLAK1f3qlQ5qbPKFmx5XVQpyFGtQNqBGj4vC4EAvHvyUKnEm
M4C/GmJx7VGCtgec4ZMzcCXJoPb8QXDOcBgPSTgqxX7gdKLn7klTdSeSJPJ+9laRZShYzY8/cHyC
jTC/cfW3/vxCHv4W7uR4s3UY/+DctanVHkQh0kCpnbQMYLF0T2NUcf0jj/l1V/ks4HesbmFkQiWd
4mqabqnEvOU9xqFJvoy09yWYrw8tTiQdUlEf0BS3k36XSH3O3UiMvjRLEFfqoXassuWEcm9/IXP3
JWsTgXyBSlVvhW55pa1H3rqCsX3dKB8ZQyn5LXoVXri5r6mj2JwRFRphtYCbb6Yh60jXJ7V8MFn5
REO8wILNKHKMNEY5EtX3iz8YWrVCdlGKyPMmIIE0BHOvv+JZdxTrUzp0Ypo2RsbxHT/DbqmUxA2H
5DREmOP0uErGE0AeX0FVnJaQcYdOPG1paH4FY02UD6YLgJPy3LJo6K3MoxOWvzO468z30AbyMbOt
WO+NPvZHG+dgGWTH+KlQ9kZY7RTMPq3tivnWtGqTmCD+RZpe1hxftW1YjepvuWlCz8KiJPbhTAza
ax9Ol9qvLqcKBmrGmUK7FQL5YQkdQoHiedsQ1VEMjbCpdsRMydpZyiZO7J2rl4n8CcKLGdI4GonW
9CJNFf5INgIZdFSoBki1fD0MVQTv7l+wp63HplYtB6CvRfc/bkCDDrgnB6v+KYtCsOYFBcK21JpP
N0FGgekuoB8w5l3k3k9UOwfB2lCNpZCYy8EcbCgEHtl011NU5q/vUqkvvGaR76KCDl5EMeJTeDIk
GS8Kw8VlZCefnA4Os8tnfV/RVOgWhVfW3y7vB4Tcxr8WtGIxLOckI+G59BMWqyq/n90x2fc4RUZx
CBM9rHI8kCaxiBeSAUSacR819CbIrbmrz+Z8pdJi8zDyj9tBcLbId+vD3f4ipDdbNlRqAexGcumj
xTSUH/s6nfP8L0mB8ycGKgoLFf0nFZol9kdEMyhBFRbZA+BawQMhWGrTWUTwfRQbN/lqtuXYw/F3
Ubm1jNlSm6/+ZYPht4UN7hCvREEKec4DwhGcQzdQtt+p+AToB15FYvTF+4JOzAjaccziYa3jvMDc
eHftvL6Td9qPZ2c0+A9BPKlIAhLgGm6SV2Ai0gJ7e6erDdCrxxyawVzBPOTtdwkX+a0Gn4vnXRYf
TPuWePhCOEmBs85dLkWVQVY78XilFcr3C91K4V0dRShXRtzzzHazwgpplUWYAhKcPLHmMydai0zm
Cq+df4DL5r/+fy95TMlUu6AkYgXSFAp2xasgoFwZuI84fQgIG8HQCueQbxYTGWj9LVOk6vzG3kTh
iPZPhPOQ4Gd/qOAeTCBq4paGeGqwV3H24eANnDR0nHbH9JI+L84aYmU9etcQNEBbTz99d6km2JkC
u9LwdQHDOzPHOO2FJP+2CIQ40/91tIgSodLAJnrAScvtPWsIfIcIO2T2ifDv1mx1DFXzPX37ab5x
oRq6SbOGDmBJFsXxFW5ZW8SpaoXAV7xjvpDC6HUIA9PlyYuTGWNcdHtUF1ZU+IcH1Ws+25w2Z0Xo
Vjfdb4pdvAamsb0/pDJ46oEYSF/J4ZWUaQe+RZQlU3sqO1jkMrMieLsoiRSo/qRo0VOjOTRSjc/f
BSwyw+wvKPq6JkDqC2PzoFC/ZLbTTPr4L0mrnpPweRJAyq0yUK7W3rdjlTybQsdtXBqmQaKQtz8W
4PdnFNM6eFqWSy5w0CDOELEQlkB1T5yFSx9ZdOaPldBrPF9TIn6y65N+gnNA9Iz+ReAHkNnvb77t
iAToQKNmLG1hNltC7VR0SF4Igvv3LcDMSn+ZishN9SqUxTLYqzxwyd8G3jv59RkLADfUOj2fGZGJ
IfmhfoinlSZxkLNmMg2KN0Le7DlFCeT5/Ch9hEklloPnTiqe6sHzrAn0kCpshgGEk6BGHc66n9wd
2vRZqyKHMjrbFpfhRmc1CeY6he0EaOZZSMSHQe0IObilKCYUix2lpOWE9qxeau7+TWZ7m704SUtg
7AKmB8InWMZvULUt3cudYbsAeKJhHGQED3WUfmv/qogbM4uR4J7nhN2UKKSV6B9DQdaPO7GLCTgW
ipgzdnwxXDKfzyZD1+a35sS4RMbK+yQtHAO9TsKvbjjPevlk+dfhCddgO9noWZXpoMcRjCUdM454
dS2S+u2XxK78iCE2UJaYHRSR8u39C4V/i6TeaKgVqCwvaXz8rC4pWrrUFNsRjQSdWRfWdx49t2dK
9ExE2UMadsiEFm0IUe6xN+t/RsW5PO+jliQt3L315/8ftDHGFQS53v5Cg3y2REkwfJxj0lAgoeMy
uWFiT4cYvED14Pgd4YeU0oG/qQHH1DU3CqedokEvBq337dXHO6fGYeSD2FB9vm+TrOJyqgpeENWq
QYy2owOWfRGH9atHIhq6hBHZ1VG7ypvKcvUzaua/QNEJ3SJz01DkB2XKwj+3yS4uiJSSXPSJ2CTL
WDiXp5tOUQySoOWVN/HNi2OSbTR/seDyV4BWPTF2umNMLOkclFUEi7Uc1OPg9DSO5hkkR6CybhDD
tBE+Hm4qBmLoQB1YQOkx19urd4bxgRxO66LEAZrJbtXwMyEMGJUruLABaI+/fyXTQzpLgeARbILW
91TqtdX65pm14Pvl47a8lgd2hdX7becE4FEtoJUC9b/Cvk1oksOKxsrHI/7vCdEGJCi/OhLFpn+e
aWpZporW6SfaYCN8O2o4NoXGrbopzX/45RGSq8+HXSZYn27+4lQIXOAd/DhNWCy6grdVbMG+/GLb
eF3vRHgEjrkpEPRxxVItTGGDxZI1OFCOHlaGZhlxuRvcHBORKhWuptlxRSa0vDIpB7BnFc7mvuok
YNDedqgFg2IJ5wn8cy1mDuQmYS87G3bun6v9ebDpLYQg/D67SG+R9lMaLTPXu1fy2gloNGrv1e7+
des4P/SO5qocVlx1pMiVFax0GO3sNtzj39gq7vnkM18ZmZAXQHAX9cVcD6aE4eLTg8BQve5KIWxI
OrOlOdLqGyEPFNXHr9MtKfq24X70Y+Jufegm38dZciezfQQMtseLyg04qijR65WNAa9uK9Wnj8QG
fe8vXHJTEHrPO9hkkhNRZRvlVUP0doJuh5L9btl+LaL2PD6h87zTsyOw/z+l2Zf3U5mJdQpAM1og
s4j6z+EYLsnYGWRrGV882+3LT7R+pdv0uvzlmegm48/EuAiVHBT00aY883rAXzUMkVzm1l3YFw4T
ZvlgtG9++KXm0iYeX/IWHG2O6HUHm+skTss+QZ53Pn5HAQGeFxXjwX4aifNW6WAQk31pddtaBbu/
EyYNciXkoM7iFgBBVdXCOlScoofkG6YZOYpWeSujljr5o9fekk5cYtsBvx5LLSa5FVLsyjJmsN5X
ClL3ELndtIaAlHhRCT6iYRDDA6ig3/+e9aup4fuYOGmpLhccVkp1Fxw5OYaHdV7xoSkmQTl8PD/a
3Bd1HCIHKWC3CvukVyN5kHnRTr9RUaIlN5s8nlacBiDjxiVr0ysuSDL0d3bmxdkQ66wh97etqmDG
wdfTdMOunGppAaoH8jypfxw+y9Cg6RxC7Yffc8rrfk0spPEQzOAG37pdAVSbtgCijMBUsoonzaBY
sgiIUTSwHniER1eHEfpi0mBoW6MtPYDi3BdMu0JEsR/knSKO0I/Uq6FGQZa8zDvRWrhmV8ARThDW
SiaA6P07EePYTalKTHvIl1ww/HnbxRC4Kj/C5V9ZOYNj/c96fyDIXinbiRA0bFmJSURWoOXeS7n3
9m2xbho1pTb8UmMGc/qDUFUTtx5MtZhhS40bfwW4XM6EfT2FdQ3qiZLPxsirwTRs88Bf0kbrNKzc
vcG0MJtKL6jI4UFTcbTykZPkzBsX6Wd1WbkoHMqkfD8iXb+Y5cTRS/WCq79Sxri2FFORt9gf4T1D
3yWZxywJ9/AykcC4Rds14v6NMfKqAaNLPopTOXYVJN4fJKO4AFoUEviVyqbhkeFN+GhtqgjLnoRZ
0oXyR7wXZNO1jS3m/C1hZdS/QkNvkeeje7chpIqRG9sKikXgXyNgNGhTmS/4HszhGy1dwnjP9j58
a1kKHqCnzmOaUwYc/BhXMNqYcl95mwOf9RQ7aVc2JzfEFxyEC5eEgfg58hjaZRLAvgeJYJAeacfX
/C0FGK9RQxXqwsWAHbAbChD++tPm+PCCeGIFfF6k9sWHg52FUkdjD72zbclpRxojgzBIqpWMX4Tu
2iOlqjQQ9WUerARigpXiQguoQbDrZcFPhTHrofC1hBx9Z2GvJ5TMm6p6tiNq9Yd0zrN9ScpBIgU1
7cllqgZJflO9mSCB/b9Y7dKPqfHZuiJKDjLOE/ALiKEwtz0pzmAEkCjwrnvN6XmmFdcwYo4RNRzY
B4ZDnXWQiJcxmVJy8Q7LOGjYt/w9foOcSUkSga7BrKvcjmLMcuykknA+mGMt8UTaXSx/Qif3i2MS
I4QpvSFfqjuzu8unAPLn//hwz5727CnmX/A/fBM22y6kb+KS/EWTxl0bGnJhPJYhr6EV60w5JmCq
f47eWqsCJReawlHpQW6/VkM47SRcb1uVAmewNXOZpMaaeCuaeSVYhrlMofSWQEFeDCG3N18nKjAP
J7rTBk4D+CItcMCEsj8yoQdzl5AZ6DvZqIoSUthhlTFhFkPAHb7D4E3ZS6HRa69T88dvwHLVjR2U
cHy+W4JJUKIOBwv9mRa1RgFHfkRr5uUQWnRydSAj/OcEbRN80SAtTN9P8zJwuWI/NsQV3hL6Wp2q
BSazRnH3F+22ispRlMNPWJirZLL5qrIkgiIIEFkM1S/83IANFzcQFa7TBKdvNt+cWP7s7+BJ+kis
zXxHgi3GijoO/nFZXiy4ohu5F3vhVSn8X0Lzjn7+nbidLmD6v0t4L1K37IJuOKaP/HR/jO9uOlDB
tm4ZBrrqcMUxMv96pjqx9G2DctLzT512oojMoThxbZSRzwEL3aHLxnKSkxUSH7corUnBUWZhxRUR
XWzpHRYGzz55vfEHyaQmt0N3ivXZzU0oZZse9nlPOvssEm/lQlwUpO4oaTX/w99z4erk1H2Wtncp
SSqn4KRYFJk5g8IePEhF5ZR3udAwRotiPK06mFTiL0ITWTmgIfXSOjgzT0LRZXw/IwqzhxWaK7ID
Qhhw+63OVqKjH44v1bVy2gfflMqNxtyYIQOWzZmCUkIinvHYQl6DAYNtsSr8+r1F7IyoJ7rkhkzd
OOWihHn2NEfk1SE+bbRtn7a/9lNxrW5SrDK51nzpZhSfC6GuvdMyH88ITvFO7AK6MMGE/R+w/eeR
oC7xenaFz50G6BGGkRymkuCqZxGXL0aU629It0FfWyx0MAgpggD/ceezuwWIESaPqTqrIwKdsD+8
IYl5YEG6eT6QE0BZBVt44vgXc0IrJ0JZOPQw+oD8pR25GGY1RSUgRo8ZY4Zi+gFOGOM/8xv0NCkm
3ZBiPGV6QvLSBCZ2NjghSwRqbcJEwMa+Jzk3V67OQg/Ii8jFzdzvRmIOJXEZ08uw4rYIKSWOp+rf
YVbtE+ZMMxoJR50qGxHcBcvuL0rHGUFTYVXaD/uHfWOIWPV7lIOYgveFInD1nRRHdirmsB5HFCq/
WgeQ/p9o54EnJiEAt8a2OzEiwIgh46rGo8Lowxum3a5d4/6baHjxEN0m7HJ0q3+dm73JOBQlmE+q
NTnRQc+5SdmvId5bpJaec+a0C6SlFCRx/ZEnjLW/DkFBZcEmvZcHC85uaO5ryp+u/cqRj6tgnSjq
PQkeLaugV3Z/douJQvaCUtTlqREqzcEhsDf15bICBtaMx45666kWZYwPKbVnHEpRS2BdcymSC5Rb
f0BonNoiZOH7yoZaEdK9KAvBdNvZAntNW9CL/Wqyh/j4qUjwQHoFo4+1BpbVniKFTI1QJULp0mSN
aLLcWMkUNjbYE+L+jGKuTzGRsnhsFm8dZmD0PtTq33iueElgM4J6GMZTZxV2CCLFY5QfCybOuSqq
ytlhJNAm+276vplfXdhXgnt7oHYlUPdpdNGtPrQABN84DLa+jWzIcDk6mBJhY7ZJcUR4IFQ4VRsa
mUpopvpT1/VjGG2vSDsWS9sASBKos/huK9mRfWo1YZrT6itaylUy+ZQLBaNjDPLLwEClp80s7gi9
scALlG8HL0kqMb/DSWTvIyt5IjRtxDr3uvtaUeQxdsL0Ig7h6XW0ytBpGDguV8VpLPQsFehCdpK+
HVJFQhJU4o9oExpkPshAlhWpP2m5wxxjau+xHx8pbKBD9QybozO0ZteQmg3aPMt7R94K5RpPqO5D
L1EkST9l7ER+aN8Wc6Wap2SKe7eJ8V4UNqIxD0ci9EiivF5+7PZyBjZ55dRA9evMX5q+zCq9jfHB
Mbc4+9I+A9tFGvas9/VLrJFvWx4EKCPnZNvDVskFfyZjMLaJsTqkx1YRxOvPdkRySL8Q6OBKK8Ju
1EE9/W19xnMkSAr5576Qu9cx326Aq431Jjk88KqtCKoOQbCt/ZHgq+0e669UcmDOl6NpFXCNW2L0
mUHkfKlELylUc6i/JPBVQVE35UYzGVws9AqxcDw5tDxd8fDDavLWsJ7v6kZYyb9bmlY8p3985Rp6
ZeZR3POSQyGnIZXVh3LWOA1678BGFlMABhsVA6jasjv6+BfVlNgWk1wPcBXHfOPfsKT6nVTZ8xla
GRx82w7x+nnxnvY6bS5xw32acCWTkDABALWzZRxZnuT3zBVzQiFn+a5QCV5ESt+lhvOaaaG+y6zN
rbaQ82u+8T9HeuQ/B/jf/i6nYGUggAhROBlst07jAcbyacRdkpeojf5yIJcCyy3DF9ZUECFMBhbl
ALXrI0Xzhd2+2B9V1T1EWpV79CW/2pKtW9dZj/7PZEDTs9bJjz52+bzjG7bxKHabxHVnF16fsR5Y
Ki5gramulHNBaRrjAyeCANxlCNrTn3zmrHA5QotUykTy9lsnRpjKvfK83wgGEGn2R5mw9WobFj+I
XQQiK3/Ye4MyeE/NDm2ENTnzDYXakkR9P0OZ71L8sELYi/GeeFEPmVUQu8yin9BzcAMvO1FAYV0C
4f+iVe8zdfDobVVxnav67ggaE7FLFneAf8F8c1AvSDusBrhEuMLuRS6rpmBUFtjuo5OkPg/hwN9S
rvLX7JyvX7zw2cYSlsptBfql8h6L60lknYcd4wblQTy3gqcVwU6T5EI6GwDKRQgovIm4ubu3+tow
2ZZ0fqokViDsJ3dEe0nmpzKs3BBPmdQwZEQdZNk5RhkIFMBfsvYGkxv3o3u3GzWf+QkMQZAn+dtx
tnVpNZ4mYSry3C63FUBOT6vFeFHZvkRANyHsGSg7VroYwUKc3leI37Y9hrtXlubS8pSE18cMBbYF
e9gfCoBpuS91vBlYdC9YLZXDSPAp+cIdUOM1EWisD+tYjMGyNY5kieKwgJjxT+C74dIOTR0fwEUV
2LqcR0Kf9wzZP9Q/bQU6yGmBN2eZR2k/lKpxn7JhFpe39PV0GKU3dPnsA6DADUmMgvukaJVF4bfY
inP/wDzg76MMJLAVaqoLB43RdVpUxm3tb8EJCkDhcM+CPOli/qCZ2dvbbSkM4pylXuFqj1RQD3+y
359zp3jeyj5uTi6cHAhf7XyRmbVSFvTPsgUKiH26h/qyJrHp3MNMKgPRYV6b99vYmDzeQTtIU5L4
is+3WAkGQzRNyVg+oMw5YRky/xtz8GrWdKVoF+CsEFdxiW3ELzfVlB8Z9VqrOPtZ1T/sO4823zjx
AbXfYg75IQ0DofZbie0aYnu33EloiBsPe8itBxOL59h44rW21JXO9CWzIh1UuHwze5NQQQ6bZwzm
jj2xPX3RhrrBQK4WOT/pNkg7wxO1QZsiz4Rrvz+dNa2joigKthPpgeKcR/SfC556pKWZeRh4MWyO
YOVWNo3Dy0cDSxUIHfQ71dgEhhjpfIJ7gINROXpc5VAt1ndGBBigYHSUyRdEnP4cURttt3Q+lfy2
ABcze2e4cJDjx4WBqDrZ0+/kndS0Wha8Czyd2GqL6IbYh4aelhjcKBYpUtVH0EHDgMwhZ5oK9uij
GvJ2g2V5GiOZkK/dQXkwy9w+f0D/jC6ZhRZ8H/2gCMjhyYs434I/KIDID3Bs6VjQhhCFsRBDuKSV
qNSmGabDdtjb6MW6hjbbcVtrHpwHJa/0s5Tjy4Q4NIYZoQAbMQsVfk1RFeavpg/XGStKYGPqWyiz
/OxHMpTwkXnwbt8MqudUyfmjscSTup5QUNaYoCBHpgzRoM7Caud/2enEjkFT8wIa7H9/RSTvGn28
9GZLotL6gYnFnzr+/xx2X9RTd6o5dy7bwXRZLlv8jNtHuEXoO8ayCXtnFGzW6GnsU7Dqwcj9c0fP
Fg6hNZ0tRZQyqlbUd27obVqwixrq0tp9EtKg8uSUX5WZ24iIfoEuyh89XBxZKpXDXHMOCFrEdozQ
Vz3j7N/wUKJmZR8Ky0QOOJjeYv3hCSmVWFAUkDrCAkGmU732ZieF8MAWN1A0JcMjV1xrEbMFj7Ld
jzzyeW1lVRVhBSXL4WHh9OngcIEJNEH2wk5bJO+RqZbzpoaNOAv2wC1NfGcaa7JDe0qKZuPrC0Bg
81f1FgJ+ahb39xlZsFmv40D/8BpKtUshhbyXs8QK2udbiE3DaAtPEvR6k7rP15M1sQOEN8mx8FEF
fBvMx1p/dL48Nc//X7hrKuCHU8sZUDOjnIYdGp7X7AVdPfnlgHQtXnh+SvK6cLi4vdjUGpLCLVwE
FRq84f1w7bSMhjFfFAmW4CjZQc9H6aQEvhSGjnLWiKrqg+LPLgiMzz/ctvVkZrrzD/bk0gdQyivM
rSJVGTNI1dDvsCayavy/m1GSp8fINbjcJB3El7yIWmqOIm+KrIt1gSwR8XZ066NbifrEyq2bxn0H
8AONhZi1KlHk3tiqJy9TjYlRYqpYYdUao7g8kUJ//l4jkJ14MZkhefZDul4OvjAY5zUa7lTQJ3vv
GddcY3S+AexvLPiFclveZGrY7LuvjS/f5LDPountdr+7XmaB6PrXgIzGrXAA7kGkvVJGNzr4r1le
qcnqWjOU1rAyN345E7H71FELnTFnsfkzl8VbRabYGPzcPmTOyUmrExR9l0WbLF83rcIt9LqmTbGh
Uhpqr251uznfSiuztPHydFSWoQhyCi/wjFCCaodHtW9nmMwO/0QieDKbW8czey5aIzcT/sOh3LQ4
BeAryceymoEEGk2qU7MSyqIruIgIG+HwyxAAbOBE/lMpLOR2xX7BZuZYwD55ZjTrKRcI2LRPUeLi
FlXMnAtvRoOXWyhJfPg8oOPBfLoIpf5RcQ9RJr8EU9mzkDfo1om1aUNqpL1rzROYM6YyRUrNa/QC
dJrL7NEol+8xOgDvYmUBvmxar7Ty+4gQSgB2mk1s4XYtGFu3XWM63aB2x+2aJ++hLfWgspn/9xNt
qAOFxmURCoHK0PWORhQC8hQAcBjSIwJuGK+5TqaKMczYee/EFIX/6CJL9xSBVLhFO/1H1pp1VuBz
tpJk7voRIAOb1PkWij5ZWY8649VVE2m37HnXpYqGPlmgS3Y5WaKFTOfch5eVmx786732lq4waQqN
sywgfOTtujiqmN2VJLw+EvExJRHp9lRWo27c4JtWw/73Sx/G30UxvlDqveN9f8KMF5mXXvgwLcif
/PD9q9TH8nzeynhhz/8sf8IxdVmpkeftvJ1vWPz+vvzkBzeIk2uRLHGSHeJ1DPFccAwPXvKTii/b
ok4Ysoi2D8pkEYb8hYXyFuMHOpB9MnQoE6Ajp48m6o/JnJ5mbdL3DAXGXRiQ1dzJuvRyKfWImhwd
GXOVi1ZlV74kE5/p5q/1qrLf2Hs2YwTdNdBMDO5r/Y6yiJA4mrTy8yyryqZmzfLJI3Cj209oeSTR
lxu7MRKewp7tyBVoyeCIq1ejcc4uxZDiiunIpxsgYYwbJf5hk+DeIcbIVUAsB3RSLMb6JIRK7lbc
GOEZMggmvf7E+ec7Jzsbs1JX3vzv8DUOnHrd/BDqc+gMhtCDWDhxsz2tIpTuAXbXjv6yVfDak+y6
kB92SkmheHiNKCog1sIEv6p1VKtgtjXnUi6McE8JZrA6W0q7Q1SyKDkOEVPLZMyVmGKNpb2vpkt+
/Wvs48IsQAPHNHXXLBHhx3x5Gs0PWkwiG50MzcFVk8GiAkZCZhzyQjAAQRy2/JgoVty/+/2eRZzz
Xp6tVHdUTREe0fRDXABofxklzOhBxcyjRl0qeFtRz6zS3Iq79A7gtkn0/DQvDF/Ljy8ZebY3QLPW
IqDlsnjJXinrukV+5xokVfgVDNqQue7auLcm5KNGRLjh1aLDX0SR0qclH0Hmqg5pM1k3uLMgtPxV
TTT0rFlTHXwpNf7Y/l/sK/G+HjP9bWjfy1CCZ4iMYfsVOh101ZUoCy7bAhMStrjOeWp96/Rf1CbB
qOnYKHz2spcQbfufIfFz7QLTPjpYn/tvZD1P6Zj274Bi2CyIOITb7/vpdWdkitJKwOcBTPz2phqy
pXpqdqadorr5H2xsC3FZn9C8PJxcOW9W7f55KmxbngRiB9hB2+iKYpaS8c7Zqt6FZWYaxQB7kpOV
oNRzd/opWbOaRbwN50STL9FgrpvzE8D0pJRH4IUjw+FV1Es8DjJPWNVrfoPIbO6ORqNnoFvAs3TJ
hEJfpQL0K+tG450WEeaxRw+Kxj+suht+rBPr7lg4h9DnB05vwW4iS08eka23n/gVADnORKpp7Zrd
WHuE/+UenAnizarxQ2NOIDtIl9Fbcx4IiPJ7lTRDVdr1DDK2oq4uolJ3I3amdRMO9LBKkeIaUaT5
yVfJu+1ZmJDES/Zt00ViTCXMORaGCkczn8z8bxIuIXiz22ghgxu/eyRy6atVaV6vXkCkfbtOkEKv
ZqGBFRlj4ousgcQEIqrb5Mk2TVptO4RUT7cZxQo54+KEvwSRhWM+h7bic+9G+u5q+1q13ykDFWd7
iOgNawM/NUTbrDNktVW4BneO7GDf5aX7ngEIxWhb4w7pSzRXqbAhaJQf/hkpQRbEJz8EovTE7bsX
GGrsm5EqBsy/DBt+t5L+nMnJOcue0eBh2SC50AvKIDmHHwNf0AoHuQHINdupMr2zQTtH6QJeg7Fo
oUqBAhQM2WqVR3wsSDPPiLMRp4h622VI2sMnu/we9hN2lEJ1IbV/feManPuI/DH9sekr2xO0livp
ssif8H+PFNe08OLty1qyGJrj4oE3MHT/gzp4eVHDoT9PqkCq11cXorEzJkvM/SEhtfJMGZp91os4
+AcE3Ccnx62/KGovsPH7eB67VYda3T1Ia0FWW9yu05O+ETUiYRwhMTYljc/dHkJbVGJ1DmYf3Ds0
5cp9a3aQWXx6xVd34I3KQL5CLpFr70BvS97USU71tt14Tkzvy8ZvsGsxowNVALwc583+QJbQBY78
SnXoTh+SYW9w9tKm/o4WaGmSIkrpmij9cZx4N7ajlrdmGM13BWP5pt4759fwvSnRxKRcjnsoPqhn
5azotJuPgAabNNQEPMOVLkHD0dPCb8+ELaY+SH7F4zX8rVgdLPcs3xdfPZUYmZgyaZc3OkAoFKqK
nUclXPtoT7Bv+SA/YwKc1syrzvtnBA2Q24gjxWL3sUdrB8+hg2g6wQXmU00KecCoM7snrzmIIE3m
ZLYY+ByLmn+ibJvnc7NxRIIduykasgfIUL83SM4LauX/8QMWNduq8/972OyrhyqkS+Y5j3fjNWQe
ovepZXGAb0LYQsy0Vl/5gq+ZOD+oRvdYoYjJelG60ihV/mBNgAkLkIhZWm98KTq18gfdp1+1Zny8
fEmQNNUKU7JXtTcqUCXfFYBJ3Mz+LoDRQ1cubMyT4ieLs9FKcCg5M3SSRIfsSHnKGrVrTjmvk03d
jKh7HbYoala+M5i2oVKUlDN5qoOlZYRr25PBEE4zPRXGgmyTIaIKGyWKzA9sS6QcivodNewpEXFa
sk9Gpb+k+uUcPzvm+jf557261z6U/Jm7zLo0fOAv56e5xEp+BCX8UsWApoWahfHvGUAc+uZD+mWW
MIUMrAaHzQLCn8JylidUDzS48cGBfL4mBe8J1Fm8HbPAUYGK30iQRFjwp41O5IJwIeibk4CF4ndF
1ivbnQHwK23GeorFmnnOHWUzRx39ljhIYzgMvpSn3e7N0NHt3/9Ewg8p/u9fPcr7QFVG/X379xZ+
74xzg7iPYtFpx3eJ791ikuKJ4jhw92y+tqa20r4LU9bkgGFmcqwRHj1UZMLxqWEph5VPgcFxPnJZ
H5MDU2Io5phDDM9RYnCw1IpU2EqoKklcF7/9bfXFGo12T5fdodkhxQWuH/8ruSH5b+VPwisXCPIy
6t76TCk9We1gebNf8BOpu3WH+RlriF4rNarRIhi2OpQr2hN1mKNja4xUeMuXnw5+3ZTPkhLOa38A
mFA7HLL5vGdTpgniZ9QVMCy74MOAsNIEqbv8X4KIbbetSWh+OGigAwxGCkQl1vNGSTQewWgv/1W6
pYAkSG839X7ogjSV76OnC2lEoUUUjd8AIHILGlGLAH62uLr6L2roin1ejz4dWVyLus18w6ObmUfa
23CPKj+YVIYjlvUTMn//sv3FcdDM/6DxlQ9jsqfKo/C45YN4+1YeLa+L8M8DeyIjz30iMqgMSuX8
YxU+BLYKIN11eMGFSdOpgAH4tQODbAKfq7bHuPF0030HVY73PwVX6dZUE8rcBUnEX83GADIXgkoW
Ja0uaanmrHeYMwm+xhQFivcLUHQ3RaCaZtordGAMYizi2bbaHwXNGljsLBTQizkCLc/SmaL6EKFV
pipKyvryyCRuybLTdrlB6biqU+h1eu07xzp+tAfXlHu+M2j1cAr+8yalF9B/p8cbAM6w6EXWMfid
RbynLpfMflW3Abyd+9QsdHDxznWLonhMBavebxeHQtC25uzdsCO5Ocb3TH+x3hITDvlFeKVa2I2e
XK/unMiwGiSWwIF+s746JZfiHMIfuPFW3DbTRn/joaPf8kaXems3tVvtrhG366XWoS2g2KWXmsQS
FzIoUlGm/RTXuY3CYcaFprEfQlfY3f2d9fYShxDHfeqaYjZUfi7nmvgCaQNu/ZeeUMcKxXQdg5lD
QeWDq6R9pLgfsKvaVjCKnfrSA65OALW68lCx+D6brF4Ynu/CZ8B5VyFCTMYoGm58JMWNFtqlLNy0
MczLuEnkQFwaJ3xEkrKww/z6VOUArF3MMjSJR+pVOA/cVSalq2I2nKXu3lvNniCLY4fyN0MP6Cpw
4cLboAe/0eu2dz1Mg8HaqW2rV7zGK7Jo1OQHYkGwixC3fBxJS5Xy9V8VdtFOKns+mL3FDPgXCvRQ
9zwrlsAwVDAj7ShL5yA7GZMuqO5Lhz6aZq0HfzasEkXZko3Z25R8Op6JtN8FEKotck18EuOU4DY3
SnP0sOW9Ydz6cHS1o/UB4GkhxRGFZ6iSL4o75dv1U9nDM8mEndvXl1pa+4c4y3/uSKNhBTst1hc6
eOEcprOvHic+WkIt3eWftQZw6FJ8NteAZH9CPA2LLWJF5Qucbae/0LGxcN2fzo44IO/1QGgXsZlu
mrcJ4SW8BvfNdoDdILLXfGtIdg6AT5XsMpux+4uutEl3BoV3SAuWxXjC1+1Wijguy1PAxkb4lLsz
pCahhYF1Y2iyGUDsKfzE/AcRPGVtTcqY9POcu/Be0oBz9mIvCxXpelb8Ut/gCWeoR4U+oJVcqgF9
D0+5C2iptikqih3OWfUfOTm0Ur4D8BKYGyKcBe5s1UVbu5IX1qoqtjlcTN461jH3OZRfziotmb7h
9rrnbUW6/Pqtj8YueIkcjVOTxbsoLjZRYCNrAEtQo8QAg7SNKh/qfibmHl+z7ct7PGxK252yCe+T
IXjAbtc1EbaKNvqQm5r4XGxK5YAyIPnxaual1Ezih1AtSFUfFGEjbFoWWPoI/zP2OiEVZo0iYw3K
7pFSMfq1sr/CUM05iT5ktoJYg1YUeY6C/EnagY+Z7QrsXkEqmo54iJRbHCSlsGkCWAXvQJZIpQRt
+OW+7UfVHpcShFVVOfz+bH1+BfIck+Aa2t3jRDQUimOpdXv+UM/mxmUvzw2WQe7LtM7bR6rTTNUV
tugwHo/1I9U0FFy5XqniIuPwChYzsM8EyX9mrDThDpzyxBLTEI/P4E1yKijCVce6DZRePDNvZML6
IHrazvaUbF/aOzsSdwpOp3len6/nx6LOEONgy1cQM35YhNxP0LNLgHqoiqn3e+MGBBuf+NzwAJBw
HRdmm/hZoib17PvwtPQX4IfwiN8JwQ9aEG8f7JhETwVq7nceEsq4iKTAY4Kbe1B6O5RaAHmEBiJF
eTf+1aYBfH4+6SkkHXyTD9/2NtkoQHVi+mtHHCrfC/ak8LKp9iNTZFW5M9DxyJcVhyv0cn6CIlIu
jt+ZzCsci9pKVyRVBzQtRK9YP6hJ/6JTmC/VLR/lSGYa4BupbZC9F4qcV3p2Pj6cRSxnb55yYvFD
hezuSfZiQ28ujXfr8MJzlOoj/X9h0SvBH0HYXzyuIQMSsGBvKDH9NGKHaGZ6ZnW4L3ZRSpISfR1E
8S5zOHHTRGBhcRh5I+QnTOF1N6dOGnMOKKAfTwPHnjglwm16cmPDEqXWmf1amF/4LV/U0ilPbWEv
DEL0Hgb6CHwoYqKEXhUqqO82ck0nUi9sg2Mh2yAjv6XFlOXEXn2mYrrYLAlg/eWn7/ozybP/QJmo
T0ZKJ+w/SQ9J60O6AD+wtNG8BLiMEpXjMB2SK6NR+jlUVV2HhtsdhG8Ej9BugO7DMuYz2S45w12c
B/A7mVOEP6IT7PksT/aIpJyXwTd3IOn1r7eGeyrgn2GxLiKLaKB165VEMD5LHTuoMRYfO1itdPoa
QmpKS/J6aZV4YFZGYTMtMq4XzeuoCFBRntRlcGSm4Lafb+3q1UE+I1GlcXuNjIc4/HtsUSJdFmDi
tQwt4GQeBMZgcaPZ997JDRzPgTd/7WMJCIWvSkGWWDewZX+fQtyc8UpxQEVo6ZAjEqwF5Q+6MHeo
wNETOFrj6OqbfqpIS7MDgaGw83Xi8BnsmuiTy+zjhrqHccDXb+cM+gkMbu1V9IQT78VFyIHfx41/
g62VmOrZrTpBYWKAjH0srLPF3mrq5N8s1HDKc1YMRnBLN3kCTYQgpxLmRDLvxPoCrbJP6wqW5O4Z
zXcTeF1X9JNyVNruuhO4UwNx6gkIARQEHL2JEEvZd0MHF7f4WlXMsNYILBr/PAHQu/3g9I05/wHk
9NCHbpaJ53uCh5qA65dYr619qKpGHGzMLpBVbLcMgMH5WB1vrjfZJr0baxywEh+Nyy3rw++Mdi/q
JsA2dIGqm51AVeYM/zpsJYvK02+RV+rtrPDUNgXZGtWPaBh+BKk1/aONaFRmD/cuJquP3GuPD4QV
Y/8A7ldB2Kmm+gqJpiK6LTc+iW5CMbcbtHq00OOdDzonvjQg/kNiHPXL+M1DHvAzBgCd6n7g2PdB
oCagzNmIfdWIzfYi2cwUO97kLQxwgjsZ0+z5zgBK/Byx+rHP5e53K9WmEKNs0eHg45WIDkr5OX4I
J6kDXzsHlltva4vO4OeFGoWO89VjJCJO1ZZtWaDxNPyjGtSq4v0Q/QR3yAoBABj7HUbs0tIdBoLh
4duKXgiGqhkF9VgwS7xNnnJIwxU6nDT2MlPvw2tA6PVJ6GXzRLR+b9z4Zr6FABe7waFGmFg5QTlc
cXXOqp4MF1FSm4XmGdgy3epzYLRbvpWZ31JGEsqbAoBSRIajShgl7g0qYnBB4vilflc4iTK46f5P
FL9JYbT/5l1P1fAi0iBamV/Jt3TqLPwSrIk0qmyyowxp4kkEyiCLGYOA0td9osYD9oyo4ZfDveCy
9RR/IoPGSj5KZ4WXZ84QE6gDiu/Z2qTu6jGOU/+yhIOoe35D4iuq0T2mx8OPPi7NJNGD37Fw29mU
9bJRv+yeuZbLXjnQm1+hwMgtGQQT9vVrc5XZXP7eubHpZJSszEJXdFnWEi2bdl0xZkgO3A5PFroh
ruN78T8GUgsqNT8ReF9StV+J0w9u6L8g9U33MCVX5iPTMMRbtTI0QcU6cdnUFi6x80ZBkTlT/mAK
l9wjp2DgB5uRdgZN21se0hqHmzEeQR4N/Hl4lnLcknw1eMlARxDupRBH2pxS3nMfNpl4H3gacC+k
btQodglfcwee3mPNTOi/Orlv1k+uelZzFic6JJYnNyLi8s7PVwOnkxM8lcBjSG4E6mW1+rMDJgw7
d3uhIiZ9Tohg8fzsoNEm2QCf3baY8iuHUBavLKM9RLEOgQS7dcHor0Z4+fDxCbsf+XV92TqMIQLD
XAQIQyazUlXk4hQJiaSzEgnxTOA+6cEoEFj7wfB9Y32w4+Kgsjen+u7GAQUuP0w1B2foGU7NHNxX
15bsO7JUYxghft8UKf7fX4cvB3WzkRDDlGFbD9siqarMDJwOyKeBW4mXRRJ4+ok8ANs1xhU+7GDD
0EHm+oC1vPz8RdF5kyRa9HCWV3Tm5CivlXXEIG4M6jtdUJ5uV7ckWaP/+pGDBlbz81zv09XU8x1A
GZaeFEK3Q8nYTOSVFzmpGSvo/z5K03u2iS8mKP0g72/y5PLRNZkCRGs7q9eUi/+eaOwblB33DwZ0
pCyWHUqZgwtOwXEfYKozmMryrA/Sv7YLWZ+TERPygI2XK2Tn0UnpLMAyB4dBxcpTOxIXyXIMiwiC
SnGAtc8aAI8JxHBVUg0w90aIgCxC0Be4XVfy2T9NkJEZHtvLyohYQVlXGRZ7sQFNbmdYD+VKeIv5
QeU4XTPOipuN//ucRv0lWugzZIYn+41O+g1Oyo5eWHMKMJAHRarn9jz8BgFG+Qz3fQziSXMHNxxl
e+GEUyPjhgBC3sGGPlBxIKHosNsa5Q0eEX3XXgwT5hXJ+EfLxbsTBVP7O91y/F/k6lKZf2HemBMN
9BN6+CYlcMAkS95vRV+ZeSTzEW8NpW6PKjpRqI8vlVShrrJpuKvlk93/oqrXJwKwCRMajTUDIOUw
iYqyg9XCtPNPdBZS3D60VUl5mq8BwsVV3Vbg9CPU0Gm3LyY2AV/NkVWtojjPHhMACXu1SiMBc3Ns
rNU7XgYd0y+MxgmLpHF14qKp6nduLIP0lkABiKAE7V44M/Tq4jeVYeSnWCwmgyJ1CZp1J+sOjF8J
CrVJQZ0S9eJHtCi/UAi9nUvg/VKybjOOfK5tJgmq/m46vMh0niuz+g/wE2bRA9WZhywpdczCcOqq
fk2C33bI+P9MQPyCLRiyqlAaDtq7gxlaxxRxlHP7A+FZ34B3bvHVsrZNfu/uzIVSvHa9HyT6FQrW
ZDH8fXTuCdIyd2fQI9togN+FgMeRlLPiekmd6kmu86prVpPIfWk4haApaKTZK+qhr7tg9Kb23BnH
xbepzHcxDCjE7jGCNGc+I4QVClCshgk56CZC540csV+rO57y1E+01OUoHJiVwZG3UyFT031AA1SS
eJJZLv/+3Rwtlw5+RMGYo4GlfQ3dWjw0eusOTAw/gEEVxYZUuXoh5pZbBfv1WzaHWNaRMMab0SzQ
5oNE4uA5oB+QjrdTRXPokNGHjxoj77xs584+xpS9k0CU3oaxF04aLi8ZyV0dTL07NQ1TkXSv69S6
1SP/PG9UpWYEIbhJyXwzUvWAzbz95Rbv06tpH0oJjxs9vhdN3WoAQ3Hlynw3D7auaW7Mc2+Uzr5k
RuJNIjj70kcJaTqQvcYkcmrq1EWnx+TGTUzBzpK/CGu8xSOhzfKJRNha3qeElriyH2VLgobt9xss
xfl3bInG8oFCB6UnyKwje8s3t2l+hee0TNAxqNg15EN1XkfD2RwgZynBPH4CH87m7e1lE6+ihmc+
67uLlN1/kVx4EWXlM+Re+1JgkmkWOaMB1oA0f74mCG+Ju0T74Kr964CaG8MdyYJsl8YkTnl4nW1A
5uqQmF0kXKE22E1KQ/BeJM3sh7OusqbyI5pVdZXQCMAHun8anAlpHPcsuGDDaiTbNAfK7rBXRp1Q
tPvuR9OP9cEP3jC+aa1rXEfg9ZUWW9bXgZRsJ4EHdZrX/Ch+aYSTCBtxkc5ORLjXROdEvo1Qps7K
9AmsqAmD0YgRWdEzp2x6esG6UuZyh4hPF/4bEjypDjNUmTmi5lGQcu08/9YfWoHioUw83ZXIpUwR
5WhR1Rgw7zfujeAdw0+NjCizhel0SJXcVky39bcutKv/yMjiKPcnvUGjmKi2V5m/SYkjSw68Q8jC
zQXtsUIWrvcd9eW9ecYhUqcT83fESMc4VFjwZpz+I7t+6hGv2g+p5QlPLCylIlhx8fKhYX/qKUkw
KGLK4gTjBX3Ofi6zeL8ZA+MXNjAuLUNyCRnzPpSDaKmCfVI1HlU97KsDzdf+TvYTTSv9Rxjp/RX5
xWnQ86EYhBzQBjrmKpD1VcZrSpAUXlls+c9Ln3rUZb1rAxKFzE/GfZW0lHWPX9Oo0CtrAxrArZV/
v7FOYfFHT1UjNzgcWDk/pYGm464zEZSeg3PcNdAWEjBLg3Fkmy4cfqKQ1o5ZInBhiS0JoSirOM+q
LZia1EfIvM2kBLbpAFFFSgtHs1XbI/du0MP/2ykWLPTmiM07sCkKP2F541dcdtAWDQMocQuWjbIw
ZZ9B50zZSdTHRFQo0M/53tNHvRxF7ekTNIY0Y3UcDssuXjS1xUBhddSwW4NjLbQV4z5Uxk2bmgaK
PlzC3QWvKc39o61FUTuDGuolqVbYHLyCn5eNKDbJGxwQH9XcauYvgwCvhCjjkMnRjogxt2STvK3r
rJVwX3Z4xq/+8nbWH1QVM6stXj7eUd4vTqCDbXkt4aKkg6Cy9mTs+QijMC0NAWjiABs9MA18b9mj
KnjUybaWWh8Dz1jt62MPEmHtGjycMD23pNmDaCI6UyP0Czz5G5q8kk8VDcBHN58yjejtiV400x1u
IT5OmTIVp4X9a4UzsGYS6C1owUAMzUwxMopjNmMWaZ+1xXOK9rQacIFpEWCMTMmYjmGzZkEP3t/b
ArgaIVkyrvk8hqATzU6+No+8foFC8XMXqcstkkpeSoto2CitMa69pdzfTwEcPrpbsiAJ7KOs+atg
qy4EPi3xfxmIuQoLAHK0tAZFIPrhVYSCZy5tRNBo+EoORTbvbV3cbrYULcswURtRc22sSg5SqSmC
XntjYYDtdk0OyIsMu/2sbgYpFHUW6j3OOjZDDBJeVcGZmScOVfEAzeFydQPeszbpOqyYB4GasAvv
+cef4BuDdWC7+Umazcv4h6iSOJKGYfWL4pGllw+uSy+lmK5aYv3AlRlybCTNIuYjuPAPuFDgJmmM
ItPTzoRQTTJuasZ5++h/N3nndN9QRimsfVL9N7jM+SrtvhNOChnFkdEJYsCrUc8zR3u11h5u6Mtx
Gq4YadrNGN+K5XNiUFBEVL/7qNkTiJU6sQRirUDg571BtCNOIFrL6TafkN0TNc3dXqg8S4+NP16z
IV1ozJ6WGy05Uqn/zK69AD8LXATHcIICDSbCRJED6V/ZYD8Gdh773KHsiGOt/7rO58ftY9/K7zjr
viIewlhBn12RCqFJ5GmiIhtqy3lesc0HCkELPPwzBoQGs18O+j2IFE1YSYIQ3pmV4hbRE/OVRSad
hcDrzM9Neg72+sTOsZoMirQpDFY9f4aR6p1iXsAFy+s7qtai9sbv5erf1497rnyYUsHwCmlw+/Vk
JTS4A6K+cBotFJE+CMOC0B2mQ+Ki/1As+D9KTujORZnQTEc5tCFVlQOZYC+X24ER8cAxOiMbQg+X
+vyKULw4ADIm+vm360q/a+q/kmC6I67Uyh79gXvmqn9vyoav2qLr8+iL/tIABXHaNiLYGeSrcrIV
og2SJhdb+EK3dVZ7YcmNuaqotDvmxfbAFuJdCiqB6V6Narz5ZbtyncLEzhEpgqSH23ylqlD+U5t8
aSKtP/6qTtOm66xyWFvfkSQUipLv4PyIK41WwkC2hnU2YoqBa6Ikp4/ujM6S8hFeE9O8F9NEvdso
eQGCIgUTOV4Ked89tRUm+Db3xZ+/pSCRdMiOl6HswJEH3b+IqpjftdgXxp/hLwCrplTnWEsJz2FJ
91OFz95aNXP9bAEz9kITcNOemYEiIVBYcG2c7iz/iki85rE6TEHssZmt1YUtTiHX55vj5l5ztFLs
dKwrTqXA4wcccXvtGiD4k9lB6ij0SIn+rDMUBRzeLxly0s+LW9YOazrBTsJRr1XmpFM14S7/yX2n
P/iHnnJWWoGsbs9uXHq1JtfVPTgWZ1FHv2xaW67XluPWmmTQjeCciA5jRpn5PoBt7JIPGtz3mWx1
Y8PTQPFd+VyTHtPicEaaHLDIUxzxvc+LJRNQiyWy2BXT5m0E0UvU7khAZ1ywnribjebV5WCRROmu
lLMxGii5M4e29CK1RYwhc/kCeOVbqd8LgquHlLSHz8FkBlrwfTwG7R5Eww+vff/usONzRxXYYzWm
5LFTW1tRcz2K29dJHZBP+4BgxGvHbqiY/wxwxQGDljK5vQ9iKnm/dqZqLADl4+M91wrlprRkaSsa
JGS7CZByRZqhEnkvppo29GObPVEGBKP1ma01dB7S9KKvaM4VdYLHx3OuQz3ndW1NyEE6dt/Z5tjC
cGak/vOR05mGfxq6kaQtb3JCK3U8bI5/5yVw1Ru8cgE3PE1qcZ46AsJGwxz91GlqKMHHGt4HDiFV
nUCVcIydVSU2A0ZDy6uPAgeMnrMZNWS5cGeOMh+u2NIGmRtifoPTmC1Oj65lv0sTT9ENA2/jyH5J
RlCkMLXfrtoSPjd8teqyqByCz3RwcA3AN96IKY7TGTx/CUR41a/q+hZUiqd7stbgdLYWrGHp1hZP
glKmC2zwMbVpk6Rlrjq98kX0zKezhdNjPKEHBfSKzZJWBapWIiCgcuucK9K2c+gTOkR+bea8BG2y
6k9zHWg9ycvqe2RERBvUZxvz6ePoLMeysBfAIVP4iTVCbffdqjdrpHJuruuQaGaqcujM2hI+zZ90
TdKXy8CugOxLZSb9iyIA8IahOIwxQV12CWptNrOQKf8fMtjebqmI/vu41Xg7ZwrkOSbi+PwUSnib
TjiIwfSz+UCAn6Zs4Jke4WvOnqeq/f2M7viB3wIwcw6+iUY0ySvfMvbQdhjiVmDacaqLmdgnFo5E
ttIc3fmuZbMh/0jj2C6mfekXL4TT+f6PUi7/42Kk//oknntRfayIaplof9V6k6M1eAbafoh2Qp/X
dagbTq0ulVSrkGcv5dzQ6ETlyzTSkzpAEGP43vofcOwv84hZlYDacbs9lphwsH2IDNGF2jj0KNLb
m7uZHOAXUbMn3bWzS+CobZTkRDcW6rcnaJZwdnIf7tXYCAhicGudDzH+eb5YGHtuSqxlYT1+tr7m
DYVw36H8A0S+2vkPiheb9POLTdA0TtqJeBm1UmJExLhAbZZM0xDahhEHgU+HK564aubBL5lGMoe5
uq9QdlxwCyuLbYZzHpjMlWRxBk43DcpDNUWs5I12NvuD2Vd0DG8pnnIZ5G0MiE4dVzu3dhN1y/CN
bLbXXggRX1lIHfvczbi/CZsH+MpERdk2+McRr82Fgxq7g17fRPAUFF2seNStBqbegnabOiJCvOvG
rXGA3sy0v44TrQzQw7IVCema3SlYYZYv4yWiFZpQdZ/kE0ov9W5hO/Q1u7BWggfHcc+E7bHM0IQQ
i3VkixooWmE3NJzBubSbnbW686Sse6D1j1lKyuLiWDqZWPCf+nNrxsJJp/1FjxgUHaMzgYEJrrn/
9KRPLLVC3+VBLgdxHdTJdUji3Qg/Nt9mZK5XkyC8YF+L3xejdjMTVrji7Q3W+/nX8kOP7qZlKc9I
3EbOzxCItCzip8tm0aHheCO4tQ0uNEcdiebxb0SK2DCxuopN3toqQXcbuLqqS+T6EWM9jdVZvlWu
GJ06Jgc4F/4NwHumEZdHPZ2SGExnTYNpeqSHNs9b9NeUyCqbMwofjleKzrIlQUHN8WQxH60qZZal
mRqGJSh2FkVN73a9Q48R105FK/E2pVe9BYax13pk5fpad3Os2r23tKwfJhRuywYn+Q69XobdpwRH
GMKOD9nFHKPiIHsnLbcPnfLxkDYzu3ioJbca6qYU2/UMrtQwuiFTdfxAQs7/RKSuNzInfa3+vyao
RDjTBN8X3GuYEOk3U1okDVTiXo0SF/vHjYhR0j1JZuqzH02R3Y37ZUX69zLwDZkG5rpU3dNdEDRA
daWbyYLUcKy5O0SksBKq7/pNUIhzA1dtPuAeSDZyvhryZrGQzHeXJZJcf+ZhcuZbYgRRvnJq9mft
581NDcsdqW4WRs78fJkuXmzohea9vPFFav+HhG45jrzecEgZiO26g5pys/2cB9iHveoQIRdHnkV6
oQks4v0jTAc+jrgsxRapCuETbxluvvDIO1PMiZksC2aOMEesaSbz/QckmFMxnqS/dyXgYS1Bmy2U
MWccNOz6CeX53TLNxx3ltazrbP6Fe5foageEGs+auJ9ZkbixFeVpkivaXI5tXVJpRUeMzSgzHcB8
/TN0rIgkzNCXiRdOcLNTxSUgII5ghZib4wJceOmYS5bQBMldqh2dhvpsLu1Bfc/oBgPRwZ81GLoo
pf42B+KG44w0HmwQ/URDmJEEk8r5Iby3KQ2TgAf82nOTh9DhFPK2Hyu/FlqpXjZW3aiFcfpSWkQE
4LioAM+dJqL+HJJzyO80OAUj20nfY0wJT5yJaEa0h0gEu4DDAAxGDiCPREGpQcR1Y0g6G6+pAbf1
Zv39fiaXo1JMPvsiraHS7sMqDHKfUUBS7sEfiWdAb0UuaeVmNOqHyANkUp6XK1qOCVirwQuBqUo3
TQ1qS3T75a/2jUwbdwKwPTyv0Ih8+Am2cIDv5H005BmxlYVY0/eycbwmr8VdHk1/yLIpdw31buNo
hKjGEoyXcmYeJrHyN5KUETZGXTR2WJ9sSTWxhpbnqlJpnsCPV6Xc3kDVERoU3NwB7aIu1EmUi+Gi
RVAZ1qtkXQ+blv0VSYcnpPepWoTBYChb23SJg/FRpd+nz0oby5zTp89X7cbvVibmXbxBmwU71ql1
J3vVjRAwPvAODCKPCZJYL7wzzwhIiuEALU+xU633gYXE+LEA15EctPoxCxpGbl4U+/zEONbn27ZM
8yY7/071TMmlsgbqPEzDnGmlKuQgPItpH7z7UhDO89qSVdIq0sRrO1JnBgn1wShpJns3SykQIdNw
fITlaCQySi2UnvzKPLlr4EPqgP+OulRo5EXXZInBL2bLEGt/qaAdB2jMX3TUdWEkaMiRzSVy2h1R
GdOLgXl93rQ6amFN3alZsYZz8vS9Han149Ni8m3Ie4d9S5mDLf5QRmb2LZ4c0k2xrCYWJU2o9T4Q
qX3loM6iZxxxaXhp4V7BNbRutLvExHCbYRCVV3Tb1D2n+1yDeEejIc+RKtroglH+7kYt10FZO7yd
8GQoSRZo6rIxydPJRk4DLIp2gJnvulYaRa2uUftJJFb6H/JM90JUuf3EmuHV56S3/65ZtOUzRQwP
M35qR8qG1u7S1UmqqFFohuvD0Z2Pp8jsHN3YyBwP+SCJDg1v/6OvFtNJyXQcX+uR0Sz0Jjj/5sse
yHThhZT0wITmwUmCGg8rY24aaMkS5eyfJ2dYMIcZEVTIZjWL0yFU8BqykM9CXH/kyR0z7WWsCGjN
QKf+Q6fMj5lk5yM/nYS3R9CN/uraUBJT9SOiR/mQPDw0uoXV7p4giyXxBI5MR1g47Hb1BNoh0Irs
xI7+TEy95CT7b3YHh4Vsf2YcBr/kYSYKr9yvzzhLsED1ZtOVYcHARqLeZEY1ZZdyW4zfl1PlEbl+
WJG433t1VqRgnEHoJJ3YursfN+ro2harCSEmnBE4YNGEIg6QfNdSzX8go6iuT2R3XajCtsb/LpEX
Fv1rgE91jkip1SI4nzY7PB3NlXP4pQ7SZFIbQh/lw7tEQwpX5DOg93L9zcTETgmhMxT8CLSdC21x
1+WmC8NxEF2duJdIDeWinAFWND6bksgbl5LJ2O8b9qQ/U0TWs5ePLGl2SjDqBcJctMK+jEH/QTCW
8ViJdQe3X4u5SoLT2+EwvpJorkdwYoyIayE7SmwpFWvScUnWEWVZdM507U7K9GrU+F12Ag0sPQNI
590XqIxUAbzeXTrdQ4cFPk9bFTPaKLl0qyYL0iWWBdLWvheltLOex7SJTWLcr5jjJD/383Zro/PW
8pIMj38iKk7TSzyRmAENO3XlzYyjuNg+Xc3JAe7tFmthqqNJOdSXbaVKna2rvW/6Zxxkf7ewFbqJ
KhrIHaOQ0RMP8nGbMc6BZ4SWD5+Fv9zlr9nIj8nih/Md1iez5O2bGrJh+ZgzV1Gy4debqzf0xPjO
blx3kenyLXxZoXqLe5TIwUOSpattN8YiWvehA0dLDGCV0c2omDtPVsnZXUGm2YDrKtNquRecY0aI
p44Z+8x/lCfeDHHZXZBXVUXV9tXsknZl0V7XRQH5zGe72MIh7rsiR33BTOYJ6LQm1BwoDNMX0FBc
p0/5PtSKAPhxOjs6chI1qQ/gxYUNxG5DElZu68lgEAeGsRfRjS0UacoBguXewsurtDk32vXxvHAs
gVhCI7Av1/rFsPouDBf2XXhhzZ6QOFwWrDTJxTYAoeIy/fBdFS3L3N7P63ZlGoCoE/z5Jo4eKkVJ
Uv1BwMm4zdsODcYkWnGW8uB7X/oq4crjbJjR2/KmxqoyRnzjD6ewB+Gvf3aScBumcbP9mYLxGyxn
euDCvV4Kxuv/wVv5VkCUS/DXgn+5VwE/pftqPRpKNyYrER3S45123YRWAEk+fX2GrCgZzCQ+f+/d
MEAmRAoo+DI+0xJxT7fFXQeGRP8jkxHORf0Q9/++QpW863CU3sWa1Lwm5cjHByFMbOopOHaOLAf7
sqrmhVGdiGzRffvZ+nIwvSAIu/cp2kFyYglxix7rTnpQfA6/U8fkM7XRSRfWd+VWc4peHpgpOnaD
MEMYk6JFoCrR5EhGdzAqIp7JQmFXmIl+S3WCXWmqHiMzg5vX0IIUfisEjD9Pzf3W8AfcSR+Hw17l
bEfnWuKnL00oW+OzEI2Zt21HXCmtBonWJN8iSPHOWGNmOW5Kpk+r7e3oIZkbz1VxP1LLg0bztSLV
XDIAGfH9wbzSlHdpEHRJ9gMIrmwQpQL9HZ4J3QQpRu+TJ0o+gplTcxla0KOCHNKRhY4kADkk/rjS
YTlBZnvLbRn18YVzRkQIwhSxMuSz99F1mIfvzTSAvbakFQc92HmchpVt2KLIHqEzscsllNsOvAdQ
HoTKb2Iq651uWB1VfB6Gl7DfRE8ripnUsVNFv0QRO7y6YqjION549c1yfjthaWnvNBWAmN9MnAlj
wC0GxAbhlBj4yOskhynPyfVOci/JTYlnCgxa5rIgmPdvRuZegA5H+UYFeSmES3zT6aK3wfplHLxM
BfNfKNhf1KsENQWfWSz3a3sILnowqOsg5viFyeY5s76XPdm90bXyewx/Q1DD32+2hYXNw7xwmsBr
jeax187CoX9U+nY5bbIyImLWInSjG8kixqfII6CQvnG1RXThdEiS1YagXEi8PztKcPCGJ4vZi0Ol
IMRrBuxn3VL4MxwBhAo+j+M0daI5QGUJchYR/+Fpz7GngfoElhWbwDzWyE0HBhvY5dJpArBiu0As
XtzQAQsxPexdsITW8atp/1fipAPGLp7Gzqp3zbz9yWmEmbpQKWAtaGCaX/q+LdpXOqZiSa/eqYez
HqKh20+32nF9lrqieNdoXJS5qjMjuINPKNLUeQQfIsyrKpS/wVV5xQb7m8hH/vmkKhL4CclaGGvc
BE2UkTFLnytcXAeiFGajub3vlhQXJCqqQ1U7tCycrhlBTbhMNAVFaQlJpn+9CZn9Ha5FQ+/tq75H
5kTuP+wf829TUYx2/rlg2nCXsCvNlryIfdgr9hwhE7ht8wROKya+zJ4sgipuaJ7MOxabDUqeDzHW
6P5CG1kg07tqcaerIzR/zMpk90GNYztsDDqGaE6TJ+dWysvjlPbG1tMpz0CtgVNsYXzFjhpBbcNh
phHaa4OWkojIlK5cHdkPjpwmlalFfAKew5koo17dn9U8LRB0RZ82nNchBm1WpfnNbznvGXUVieSj
JNjTZPACgMkjufA2VMXR/hyJseq477zGCA/R8Me7fYSiVecw2tqS1GoCSS1Df/xMtQolvL3+iq9w
a9zhv7+XT7Hg7lQ7w0SHdeSm3UskLYP1dIOiKLBg+Rf+wXtpH7GxIDYul+LFVw40sObOeEMm6XLk
vxwWjjiU29A5OMz6YDliQi3COi3XJzd7EAHlFOBXlhLV9ZV2haB+/1hlkp3rsUDt9hGfP1scdF+N
ksE3PSxthDEuVB2C2QZPW2KvM2IJvVL+nZte7UyNdBLUT6CLmSIKx1n+9/b+MllGQW4SwM0QmkVz
e+A6AAsVjdjfkbhg9/SxTTe5c15BKDxWKPF9Ox+9EAfD7b5us/dDwJ6sLCNfUmGVwGSDmd5E2RXx
IQhybJ20U69UkwT5VAepm93/+wbnW68oSjiTZRY+L8UoCEBl+vuRsAvV1P+2FVqzzU2JttP9QZU9
Bw3MpPTzCQrBBg+fAWUJ2PjNr4wZFJ+AEwMAIroU/8617H+HpbSjCoYafcO/E9V9evKzVnK/6TA3
XSPggyx6/mIAqOAK9J5cPjq7Zto4IcnQs45fyGA8a5SQT41pm+TxEVmi+zqYMB4QJwIvzCEj3s3I
1zZ2BPBHL9pr+l1akVYkY8i3U7tW3FNdvOCXAphBps/A5BCzw1XAblnw7VQqtNIG3hEmBuMJBuNY
hMep2jQmKLycoWc+0+GoiOCd4FR2aXbC4QfD88BjEdz+7eaSy3jxHGuP5U5nyXjtnb7l8W22uyoA
wuKLySuUcvQ0xM19+0IdYKCxV/HyLNDye3ZueGquSsMF9D6JrwZs4q+/OKGswT8h+2KBMiQxkmhc
TV876ixtO+2lQOetyEfPgvTNnCBWUiI/U5jPQSGyRNKUXzyTOrDia66N+KVG7ai/f7Q6ovHPRYLu
C3PO5nFhWU9kxHxN4aw0X0tWJwRqgw0veuYoFGOb4sc2PqHLWMwzyMmygAteB0RMBdfEjZ8uDCrh
ZzhOAeagRNvqU2/v3iDL6R4kAGh8mwmueaGf8V3RS93ApOxuBv/oqRh+DLPlxj4u0yIJswec4Qvt
0iaKYplaqbnfFat/IrxCp2HSvfZQCLr6xMwbznQnaH+uhX92oznR5/V5hqnsoAtK4qMvcjr/VCn0
4IStHMUZvAuD8NjhW5iSdRxv3J/BRfFF3C3XFirGZwKDHCYAbOy38rMReoq2WRgwDUuUr+g9x/8O
OkfE2KZT7W3GRv8XXl0ntyTM7V+65dqk5EaeaQsc8C6dpTHtLFvzE7W7XQSkl2yUIdt6vFodx1jj
cTsLTY8g/+5JrFBW0bMc366NzcNancHkG3r4HDjYjZWZG8tGdaWw/wBgqk+yV8nckx4g5r9Hi5YB
XauOpvHv9bi+ipiO3SGUb694+A7aHPyrJWuln4mLT2rJ4r1TapBKPDJ/nlyjdqMnhsD2dgEYytcd
EvyPrrLM95+zALSEehgQJa82fN3R/KU6qAd7ok9auIfXv4/adkpwgYjfoxkt119p8MZJk9kn8oeM
dAQtllCoWlabt3nCv1ScP6uh5TMeDa59EcT/VdRZEHocaabhmZ8G4e0p1QeqdsajzD68m98pHsQN
KJ/v6+pWQOF9xiRczLNytPH/ubInIpmsU7WGkGa7gFBvgsuspLX9TFzMvUfJ5M/ZVuOz3leAgKFk
Fj1e3ji+aDLfMvgGFsfdbBeiLerbQgl75JRBDJjDynZN+RfS1cqJE+fw6+NipObi7lW2amVbuVac
d+ZeTAAvW3N5ouSQFnAfTamLZaI/zeLRyJr7xNxRKr7a7EJp8dgHK8Fm59VC9S6sLrHqTwpQTPoO
SUC9jVMyZ76ahNiD34GEVup9vjdJ/zCO+z0/gTigsc+rg6/QSKJXBs9B8b2772QPhisdukPzoR68
A1PX7M1JHr76kucFChgavWUeWrY05tGTWJKHZkaq69EhqcmILo0Wpv/jI/ZHfTX8ahLWmwahbRZG
tyc7zQ+sKZHi0g4jtVFwwxiOEFskwydowDAfAN8TPq3EwsW8fOrdeHS/2ZB27kb3kmlHf4a9FZUf
ljOmkym1e+xfnJ/0hSE+Dhp8pw3Lm5Po9sZs7rPUJkmm+eukOvS/Z0cRFSQeGwTvzxrgZz+7ZmSv
nS5g/7IjQe1s7HCSc+Hqu1rKKR0xIjIEjLUKsgVmjW5BpEotBtuM14P1T7qeMu97KUM9cj1UioHY
ejG23PCnxiAaz0+OpRij1+dBxcoKOlNYb22tKzNN752YR02wnDc3+MNdbNE9z/t+NNw3SG4pXjkR
sSsrSKkVavTxMpZ8AudpZLQe0uRPSHB7Y+LaN72HYIREoslEGHWSNOXkNJhv+BHfENUu3qdOyPzi
9eD1nxqeQvcQmhB67YV/OC4FNDNz9LgqwTZ/w/T/nmAmxosgZjKpBls574NdEc3l9KYNVI0LkdfK
BBSxj4Vu1m6YufAQSKvTuDPTWpBSTyk3V4ZJg4bddYfqndFle/IIZPr/ZdjHOUoCLDZeOHL6KN+2
2JDhNvHkyL3HoJ4j0wwk1QeJb3pgwZH/JUfC9CCuAUX5AZ00UuQ9zxiqpmJ7978JjQruPkmH8AiR
/V8fTC5aGunJgqXU7wNDjuuWyJBrn/IiJugkNE/FjqsVX3OQRg5b1ONQqhxzPCfEeF3dJmQBjlCw
Xq2hyqhfhpabVANiFsjnUPG5GUYk4Lc21Ta6iR7LvP31vF4PNCF/iD92eUSI13QOE3tR6pGsY8OT
JpAGG3nhy8te7MLrHY8RSVhIQrGDzVwtiFXztm6D+Y1gfUinEJfsJdM0jLN6weAh2c8yUKm54mVL
68+ypyjLvirDymmFyMMtKLszSHwyPa83j6IgEPtXJuqHqKTELITVmCMTgDIxqHlLu8CqXAz52Sv2
Lr9bqgmWzKUjAnChVgENS2JvZl1TuM2j6oqmLzXZgDt7v5XgZFDe5YccoNp2heqspzmMYAX/IvhT
TTQDhkM75nVb9Rl+LP0GL08SRKuy89K30wkrVE+MwBXBlWmE4w7sM2mvDOxK1XL2gsgAm6Lyq62R
bc0ap9G2uCvfNuod8e84JvOMFh2qSImcCs5fOHQOX9NxMwiF2i/Q207UL/roC9etjRDiuDH81pp0
BacAE1J8EzlCDO38W/AexL0dl/prcYlNsVbh6vt00F/QDSaX/nX7rCqo22/cbP/dnEnBSwF1FEvL
z1XU+/LbIejzaNJFfpUQR8mK1waBU5ue9sSWzU+hLAI5Zsqo39hdQqrZhDylr/H69kIgbiN9ID/L
9gCzQJWbJ7Ey8UKf1NMFgSf0HnarUbPKrW5xkDrelGAphjUciqQC5OLCLcevZh7p9P2yubAE3WR+
WoTKYLYG3EPZ8FYKljwf1JpTpveyk9Uj1wPqJEgsTTyjLqwojxpdBM/VySfrjzTWolJ8KPPlbn1k
JGuoME4GvAduS6+PtIhoI2LS/7MCSVmuioEVv/8bz8xeh/OEJKRmdNoZXzAnmjsWwys8L2fCtlSu
4cW6fnw+C/paVUFiPEYOK5Bt0K00GsUsQnsW8YISN4CrEVNUj7jBmxiC8WlvGxYqRgZ9UJtwql9l
yzKpVCpQQskpDeZRGstwKhfd38v1uh4V7JLPDVfsD57Wx+WhPc7tL+goBMlIOg1yClP6rD8ytFH+
zisrO8waMkhTJS4uG8NpHFAZL7G/CLSCb/qV8ModX8i+JO7jKKhuhMMPRwV2YTKIaHzFgrN7oe7m
86hwqcGzeHlobuv1bUsykip3VDg8NJ5vQG8pbQJZFwNG9LXFoN82WwYFeDmklRVkuDdOVCwx1zTy
T4nlnAhHRlIUTGJUmmQ7Oro/1xINGgBn3SrPrG3brEIBccvNLfxjSp3a8QlmvPiXHJ6OOApSDD6j
QsBXLJ8dEKvpdgB5WvCihEmK5eB7XmjdWWzNqWYegoohYEVzh5E0ZtD65A9nDdIB8GzE2DJrT0Gp
/eCULBw2plwk4h3EXIPsF8thH3KB8e5PYO0o1wUR4P9E3bnAnFzS+7CrqTIH7aF5B4iHP4yYzWw3
kIZcDnASNR/ZUZ8vbpBp1WOUqZwyVVRF7xI49HXahVKGvpObsMaYS+dVmM9MhGA16u2ypkc5dcIM
ajqm66j7CErvtlXDwGGdH8WJYHrNrUyEJ15QfLyALuAWLyMch6PlU+olT0dEbGo0yA1jpsvPYDtq
Y2eh/jaAAiXvWc9beh5s/oCnsdFikjf0/jE4MTi8yeHaLkDk1R2NphtX+hlbQh3yJPs21G7qSbM1
mg7NINvfsMqoPXlhJYmhuM4nIIodZZBY0csBtnN1Uf1ZBIJD1uxygbwnXw0s6ocyTO+yuiMIODHA
19mEu66q9uqEQRkk5Ur7CbYgxU/JWH98w9llJEEmVgALcjiswMLuawQzR+6NO2e53VDLsLpYXT0q
iRpWWyOJPLVyBiTGdscirx/bY1mnzdWY/MrP8cReMNSVnJSULDT1gxsxltRz/naSJepJZlZLkj7A
Sc51iVmtIPI8AiZSuiupMNVLeuUGW48tU/aVk27qJitNa3jSHTspkktfFNvEfmjp6D5jJ4TaOWRl
iJgnHCjKfnsdDd66ZFsvnSVSWkMczqXPt5d13zBhOaiR8pHMWB91UGdIphsSrm3XLudyvg17d0xG
qhxW34nx8EjGL8+J5D+VxNQzvj/OBTZqDmehKH3jJJ1Fg7S9uz9wtRlrkNSW2Us1CaIaKdo1dN76
JRCMZWLjIq4fZTgJFcXBqJpUQCNxX4DUEhaj/n4mj9kEmYxvPzZV62yPRC5kiZafS/mxKcmciDaP
EMEqy+sGP9MW+0wkoLVZTXmrmc8nl7dSPgyFTm4XdlVyBdzX/X+E3cfOpv4YElmuExZW5puwmM2L
raBFXgJ5LLq8Hu0VXqgWnFViBIdahuz2O8BtHjieMa+HChPZNmMxrTsAUZGYcCY/CvZanaep2iUU
Khg2Lr+3PEpJwIQp9UwwfgCuWdQE5usEJ5MbAOHPAjVrazyKi1erVeU9m1tXwkb3AMNsG4LFo0oq
E71SYZKVq5kTxf6Rx9m8QOwT9ednt9AVedJ25R0f7gHCvEAXKxRUPHETgU9vahe9a+K7GGrmYZED
59s0s2CBJu1UqintAhu4pl37sK0MoKyUvtTohnWngKCKQbabb1aNdgaRN68NOgl/MaIPfPkWajGd
vJk1XdwdexTSjUggW1373iGPMFA9bPilr5qJQrVZJjj/wXJ/6GTCenDLETiY77aTz2hVaHD8x9UA
ED89PruCKghlnNtKy6G8z5UaMZqmPNNTqcuqUIG6Ri7tjn7vNZQ5EPNZwVMOVaEzVfEy6H5MrUgq
mFoLgIFbHeKmiVSG12lpqvS9QCHccGi9CsZQOvV7wZLTmSmW8IOGajQUum5h0ti3piLgppMfIhxd
Yuk2ufPXxrwH7lol+Ud+38dG8n4DTIh2fNXp8EVgRDS/EyV8k/6VEd8WaotnfveR+ZA0baR5Vw7t
dmXCUpvMHbtAA3hCXQu9hCE7PfNG2/zch5KvAJfOBBWFK6rcncjjuFCZBOc17Z7oQI4A3UY2RKaS
vf+nHllLqEuZOcbzE+5GgCF6FiUDWJFNX7jae6XfVmzRAPV2mdk8Dj/gZDAkYDTtIUzOPV2w4YSr
c9Nf+5jxKX4fFOIDwFlUG016aZMzf/cUGDz+XDeFm38uzDBfkmEfGotVbXU3cjxLTkJlgJbi1KcW
yshYuXBVHNdfhkpdjqJCcGStOeh5YSa7OvqV3jyF0mxu0+SvwB21zNinl7zBeXcxEm5kXFWbKLa2
BO3WmsSzvR3FS6wiepjrAcWy9vrKt6ouCojWRawZMw7oviNffs5gtRarB0CfytjkWWkP2GtqKjH3
mq4JywRGteXfEyQulbdnKm3f582qOanQ7cJCQplXOkuRF7fdAge/ApesJ3PKjxx+8ilBof2irgGr
U2FRJgsYtT1jLDur7A+/2CV13IEWiYPUCNeJF+taLcchNnW+w+FcuQMrcmksmoT91Hj9sGXKI3D9
AVVHtg2QU3D8GBCVXBSqsCVHWmmOgUQkpEDXYr+mPeeEqlRZdDuVwiQcvm69IVvk0tV0exVo4fQa
vjOB41bAFl7fUzs14jxTqZ8hbo1tj+ws0rml/2kne8cmThISGTlQA7C0MCVxblrLcWA3MDiFiqnG
IcckcVQf1n1briudZ19rPvuBoRNKaVVknuejwjvdUUT/VGcl8xr+iWVgpJGlzx89YkDR9t67YsZU
CshUMzJjqo0sB6gcAwm4aB+qv2rLhBMGotyhSTtJmmdnu+PKlH/ZUTDteqKeP9Ve9Ca2vWlN6upU
EkBHPkDSN9Vw0C5+ZjfY0blpfHolakwaIMEYmdkpA7qQIC9EMM1Jam5OvJ5Q+B44nw/usYXQbwzE
6xB8++9bzvUdint+g5DKuflWVg8fkrAKJ0GtiGiBuw9WR79cRp5zD2th5BCR11TidnbPJVNYtZur
h/jdvLJKjyg1rWBTCb1En7RHRlhoTCjESuBrhOdeU/eEO+acUpVc6ud7sAEy17I25tcvISLzh6cF
cNiEQZad8jmVmfspC/ZJXcDf/QqQMP00UQA/cq+b8DqXvSxRCwkGQf+0Wx9U6jsEkYhao7k7FNxO
Wlqj8CQ5IQ8ipPONYEcubM9CvFoxm2+xkQF1zzTnxiN7Hr07ndWS1TTFwe1din2p7IOGD7Cp0mrr
CRghalY3pB+PwdBLH+KSsY/+3+5qFdQcVeGglxra5bp+YqqiWFmNoWnb/uPFGmWV7lUQW5sEJcGY
sE9Ig0LhsGa8Ltthi6grwLh56rdiWUcOxXHZwD3pQxn6qCeX5hfnWTRqGVO1r1ZVSTptJNgGJYqy
Ykl5K177C/UJ5ismINsDgKP3GBbESmLUyR0ZmhqoSs4OBAIKMZgozwUuGbB0IIGwwqtM59SloLDm
jBlKHlmWdCdFhpkD4ctuTuB8Iea0HvXWsKV29B9Mz91ZgLwBYXgo3qNXCbbqsEtY9b9al7BuSQje
XEkc/9R9mwA768lNVZu5rsBSw1ShWQkDMoVX1kKdlVN0YbSfzil6QEdeolAGE28FyIP1m7WJXf86
fSuVtGvwlGCo4auh5rzmbRqTAsqtW8siW3V3V6E53JqXWRPcFnBTKTFba4e/MQivk8aCHzBOTTdE
pFEBUcKgar0HDYOj/slwrQ8G8jK0SR5kxm9nmlG2L2D9iwOq6iZoN4HoUonh9txUXeTvN33Te3AM
jaB9BRi40CJXOYsyGOQ1BDtgQYimAzHDenVl2/Lm6KtFkl2UL/sShMEKuzRsa1ra2zU3UOlL52Zq
uWdrzgUcqDge5klX5JITiGveDZe60+6ksjtWvVSAreoDw35LTEZGa/IwttGxVD2U/Yyko2CbMtmO
lfPZm1vxoCX8cN5dzROOQMZIwZAH82bGXhBtA3DYzLQirzSmBjorRAvDbFYzfSv1hBQWJ1Xv74t0
a83+lmKOkoKjmtsO0rp0JXGLQC6t39SglMcyxnxW+y6ExxT+6i5zoc57GinzTlDvwf3NaHqfXN3N
MK4mL6PxjGsmh64QpaGCfLsKdyYsElMZVqJjg74N26yBm9sPbl35nDhlfohs6tyufroCEx2Hcw5R
HS+oT8Bwz4uI8ssOVBOgwv3Rhs9xbjcgBalzlfiLkE8CSeaaAJQl8sCoHuA0OcSxhfBhOsbUDLv5
lqwVQa/YMf6v64ADKNs8FmrnkOMJ6yTf1wsTt9Sf4Rp70OQA1B4b/sAXetadmWQ4tw+m2EHLFOaM
J/ce3HXSBjvzggoAAsoR5xU5DTCAzPPzUVSTcac2Ehaosu5dhy2QA3uvGELLAKzuXcVp6iJ1xRbU
zNtp0ikhUh6yXM+BWYmPm7YPZhHztr5R6RAiq2XlnNcMsHtHZ5gn+gxaG3KbucznmbQF7WPYYm3k
sB+jWgjMd0Jtu83LJfeL/YuzJzcpkQbu5Cca24Jg3pA66G+t7WCNscosh1I5hv9Nw1mQJpIeO2zs
vOuW5FGiZLCv24n7pxuvOcjP4sknBienIKik0LirhWWJ85/T2MRe7ZRqOuN9Yn9GmPaVb/RaUXKV
p8s4o5TRxW9Zzfrk8MG7KnoUL9yzJgRzxnok/PaSX2jYfqOzgapXUkvyMiC6i5nlE3h1D6x1vtZm
e30nLWXlcVifObvpdPrm7JoTdw5Lt6sd/XfXZXs4p7g2xytw8HqSh/AlYoByr9yITCbe6IFZBuxz
Yva3Bqmd9cq7n2CBSQ77NfORZCpfXuGHGdrLIC1nRW/valDpJU0NqwnArP9rHyMd7rQq8gjM7QVb
E9ROp0krwQRTXh+23/wOahtkKMo8W2lnCPBsqqoUdRsi3WHs3OhufJM8hnjp+4f0Y4LEYBR36AQX
ChlZ8Uy0P/p8Hky38PugcmDWfzcDinjpMfeRpbefiiMdQlTKCvzg1VCpEY3vQcpCohV7MbbcEzFA
ZHKXi2IurXzOy5xBLsgXOemxQFCdSaJ8daVfFDy5u0gFJD35DGxYYHfYpkzSq3fwioKg0aiatlwv
/Y07c1Pe208baEnaHibYDLT+ac8aX+CYfZsPFTjtiTE3grgOExt7CLV8nT4QhXXnT2+IMKNXGQ6+
DqFIZG1aRlgf6edB/Oryi9YiRr3vOWN/XU/4OeDMjr5225qcF+2RCWUL5PlByx0bj3OALKoMYich
25u0xzhLBHnXBovGn2aRMwLe7MNTFpESo00nhRpJ1fBdHCtanOOKCespliX2VvKPYGhw2HUiVJBb
qyG3OErFyxOkAX8qVkBsQQr6kWWwmeEpmUDgKnNrhcyTQFSJvjzTrarpr5RE00M7w0PE7bAIhnQ3
J+OIPR+PZN6iPuEu2WY1o0eOb8fLPeW9s6eWvwgVBB9rV5Hajp3T9cPhC2wtO/snGrPgnJzLfMBx
cjLvTHOXTMw9huM/9a92x1mUf38l/pXXwopMBpcrh6Bh500e2uM/lpUI8+UoQHgnVRmW127mzjnJ
62QFDp9TotRzpHLfcBoP1tAsOnRwaiBrekwr8YdOaMBF7NpbMwGDPvZd068ql3LpgceFfG6NzSVJ
ADsR37j3jTcmkqMRklD8PoIgKV8+BMAyx38uFhU/Sz0Q2ZY4dec0myhLHvoBcPjFSLYmmcDIm2E+
XiOpQiHW0rDvDyBXDspRCn8DTutAC7I+HQrbtWxaGCyuQ4znWmU+ADD7EPIdGx2l0HXw3oXaiEro
QjovP1xgF1byT5qah/zk778anLeALA2keg5MRV/s43I8Ntmmlwu/IN+UqvA886oGtgiMrZyu4/VO
nIEeP+AZaeKZghbEBMpdT+GrDG/vxYVdqcvhiz4lAtYiOAfWLibfkyQelWx0bBUJCDvlhMIocbV+
rG1KeiXSc2lM6XsRR2H2Vr99iVNYtONoVWo1fsr7uWssJSPEw8wU92tPog+n3Y63LJtLGluMT2Q7
uiXr3ogljsi6nwPLYEXGhUAY2RCVVyBCv9A0OJZOfWxvDntRU63e5GJ+cXdOFy41f1XPKFHuaRAO
ZgXtXF8Atb7socTrBVFW33PkJX4zi3ZzrLi2lhsmULZeMwnCvtgbDWtEyTqB861JJzqr0smoN5C0
lC1Uvy/6Bx0WRSDHcoNK5VU2n/k7AyBxGBdLCXc8sYZVb2YlpKxmfcO+rsqGvktK38UjXDJJaLpg
R02/nJ51HJwaJjIues7rbGXLlhiFKuvp7wV70FWii9AIy5N2N0P0fkhopd+GyVk9xdA2MeNz04nM
WnfER2MGCnjE2lsYiTXpKkoa5C75taPRj94MPWwVe5gkiEBhUTD2oXjpqMuLnJp82JZGilAj/89f
6DUJ/T1PkyoBR4l1QTr01br7kK32o/giWlMChSxFF0jALBDQfybUD/lDM2usstmHKI9NwQhk9q62
OxOcRkbd6Z/kjn2YNQDDNbOfDU1Qj3CS7WthOm8/I8Dxg6n+xN64X2tw3VljUlp3AsI4ecRjZdef
Ezisjlwr6yEc2dwGEpPTrzPD9B7dTPmLaFVpmcK+SqvX84Mk1vuzAklz3ar6+JHHc7N4LfJS2oPk
/VucLKH8Unoof0nlPJwKidMbA8KauOTKDZOm1M2rOgIg2DE97CreXv5YCn+1m4eK6VkFL996LGt1
ciRsmNFMggNeaiWZo490r0fyrqpqEHwy0OT8IhNPmp/zM28K4hv2C0JeB6puw7XfMII82pHtk8Xi
eW816XpBn2iEfPNtTTeD097X8+BdGJR7lehSIpAjS//oLsWidPMEtPZefSzjgHshT8F9cF8o+wHs
u61/cNh1RVRyJcIv13WHDJyw5PBQW0UrDSWDrkfWGLhMsL1/bqQ2EDKM3s6f5Ak25cEROq5IvHOW
FcArrqVX+8yP52hjRBxARvWBry6aCkMFnTpDaJ4UqigdGfmjk30WqIUaB521o44eDRZKjBfC2Wlc
2B9sp+JtjjGLZGyivGDA0zWb9SfPGqG15KM//85C+iM6m7u1GEbzgZ8HWhI1Fr8fh7dfuGJbGbIz
TTOZ5+NyPtZJI5MwEZucl5OUDL+sVvmOuf2jcAxqAqJVb1A49lk4BW78T3UQ7rqZDEQta2Qc9vDD
+TFsASx4qAy39NY8H4mYaRsYrMU/Hsc3cAW1n33PQqRGrCPdkimozktxq6qWjd6vTaC4ml5S+MEp
GVqupBHRGPyyvEkUCaoQ8/maqU/RgPwkEoFjHf0QF4anjOykj35e1WV76kNzz2MciaSbJhF0A31L
rCydr4kjFlkD1FGaWfz1Nd3tjhi1KR2UaTfZZU7ZjJL4S+rRRn0DEGnlC5uz80Jc6/i1Jrsi6HHH
wq/mI5/qgiy6ITP6dUYH5rKRkek6g01dbFKMQ7qDLHwseuW7/ALZp1Yls5WsjF+PqxI1aQ8hnixH
1+B07nLeM0/tWcz4S2+ajzBuUQRafDuHCXQ2GFz3lFjqMuFBFxYitrYaRSI0b5rirMyruEBElU9q
W5D2utIOsqZs3rvQBlE920lqcM6xdjxCJ0ryaTaOo9Z6JhgX8FnuQV6O+wEjReXAWEF376EL+ZKC
YcV8zExRWy/PYqyWr2V7vjW4jiBcLhkfaHyRqk95UqUMr3FmnsDQTbfX6yPRdk4XvHiepEAQ7NWl
gXU/3fAkjBOJ9fCqIVQ52wEsFRWaTUh1d+jE4N4smNJXzuxgod6qiXOLtJPlGPVMzk4hG8TAKJvE
X7eQ2ueohL2o4QC++FxWDArPIi4EZd+3oy8CWu3aldVEtup4BgRlOsOgIb5Gk381EwGng6BahPDT
uzkA/SZZQ8b9sG1fDJjYkpX2/7rEWda4k4IoGaciawP04yTosugyg9T5xy5kdCh3Blt2SA7Du9Zt
fg0UZ1hNY6yXbaOQX7sORmAYL5HQXn7Uopmft0RUqcQzviElX6QQ9D/SqbylR3+xnNfPdOZWLES3
qIyXEJhzy+jCt8qVN/3uDAfyH0hNGAYxW0EW5uzYE2le9cKcYe7+lhujOFYP4xY7CxiI4MeBhjSn
FQMOTeWYYc3TFyc9J3Ys6G1eIh1w1qBXfT0oYmzY5VuuHraLYoFI053AHoan6AB1i65lZxL6Mi4x
Tn1fXf85YjFJxK1JxiCABzX8I4SN/Hfxbppp1Nvl85Zx1THZBOCwUS91bSnrAKgv32HCXa3xLyr4
o5ZxLAVxOpNdWFDEZ/FoM04uWWKl9iBFL1J1S0xZCi0NJ1LFUsGfu6CjXDOm7dsbEGFNx25i3a0a
0so9kWWIgCYAs2JjmrOqyQlPpVuU8XLfyDNmHXJKXvRqmd1vI08fWeMd5pEgrBNiTsE4DG/CkSYU
bY7KYIjZx/kb6yqWCT4GwoQCE9w+14Yt4r52BDcCj+mfL/Dqdm0dothODTlh/xDIe68obN/1Yt/E
7uTWyQhphuQCZFmCnQTSsNH2EAn1DyAT7+BC2LsDcbKuEr0z7OT5jTmdLzNsxMQPnAoGD+tlvIvh
uq/9fu2HLXMTED5GXpb8tvw3rf9p/5JARf/YR7AsL12lQxSD2tWRLnfcDmOUiK/i6zxl9dmCbxLz
wPPDTpWUnJohclIdmBPkvE2tErWsVMgLA/cJJ2JPKZPzCgS/dADmnExC8BojJDJPeUG1L2ZznmtD
R0DDLzFzDEyFZ/DIQ7ZP9YMvzlwbH9SX8B0EeK/G3PbnM99sp6QWj+rSauwBuodC9GrmSmH3FS5j
al1D5FvpVmC1jVtlGSAKzr4FvnBClPQ/p7A0x+Up7Hl3pnD9k/I6F/PwA2UDVNgW8z4L7r7D0X6s
tu1dQeVzLbtdebVTH2ktOq5/E9K4EC05lgMolDQ1AqUP5UR3xggHIC/S0jlM7OVxqeAfrIqEAniX
sYU1wXvHCiXwuuvM8trdvowkHmH1atybjUvgHGHz2SYWF3avhZqCdvy0nCjCpmn96NnvSKQGYACW
KOUW8JXwe1s4M45kJ2+yRjw5XkDMEW7BnhkzQHhVdTLVPUDRHWnhxDORqe/HluctAGZIuXHoPflp
R6udVVciiSROYIG+gZpD4d+Nt0KvtQxiYZPcl6zfA5alE6bxGK0S6IsSZ22YQdIqxK2Wv+AaGo81
TKDPuHn8xPpr/HmfJ8jwpFC9ebda5Gogn/dI6JNxyi8lsRf0y2v9RERUyzGWFRgaL+7jRd2M+If/
9KBDgoA9AOD+oexHC+/NpVa1EIBVEIpZpKvn2RsZAl7FsKcRSWjsezCc5vzkDzhngxcn7AyXCaYb
YItZgvakE4bgUSKCcPoPeCRCI2fdtgEpo/0XPla0VBKqTi3KCPMIk5OoVl74a2MvDRXc2sXb9W7E
kJVJE/e1s62R7V4nDa0cuYtuSe5iHB25GhfLcqBX5CdmJLEdd+o+Ya4i3+edtlV6NKgPsAOERAO8
vtQM3xyUcRaj2IVnRI4yw8X5KisXHweJ1KmBjLCIa6c0n5VcCztQ9ijLjCDSMUho7rmqCuknbiiW
LTxYKM/8UwmPkSnp/TBHRwHWE4pKTGLJz+ESLCSMOH2g1weg2UFLnzUfkqusSaZKNcR8Evlo/w+Z
ye5oz3Qnlco9OwQQj4Dw+FXDv4E87ckYh8azt4HXbb/irXO+uVGS0LK5bXRGVcSB9tnkos+1k96J
J5GmHcM1N/bpfGkcEPtUl3sF5FNNv/VnCPyR2yIyoQ/d7GvYLm/42X1lJZg/Dj3APUvf5JRN6fG4
e+IqSusNDp1qUpsuhj+Eric7lp/3oCPq+bNSvAkGmHmyZZhquGJIkzqb61D6mLwwpZx4WUhvAZzl
v4fKB7fsgI1gxbdSklh/qxunX0iqErk7brvQkclO4sJ/Ms2JwxnQx5omcI5qL8ku+jsx84C0GwdF
3REsr/ZS1ki3C+11XEVl90+O9DErMFiZ2ZLyPi5L1uIb+qLSVCnl2bgHSUDy4A0scS/OBfCGKzyM
y1txufOzFjO1PyM5qKIAzega/IJ7zSQYGXU6Bz/kYgSY938IAKPLkHFvL3BGtK/dl5Uijmyx8cdt
YfF6CGCYpw2Ygdr0gPR1Se1abG5SB1OVtwdGeJpceLGKOWSxztxM9zVYwfDy5DPlPIbuUeDJ+iZs
7LA7qJ+2x+duJucd8rvXnq+D/HDU8ViWh9/W7zaskEqhc1gq1PfyN/05wtHuwpyZOkyZEWwj33nN
tHh+mW2j8uEBGBYDahS7ZTi7hof15Nv82TIwWSCfN1x/8KRSaO83xyuLTSyNr6nHFdJcemeBgaYM
desQK5tcHW1yhXnz+Oln2nSrGlKenZW6MAJUIYDScKgiUbPnKW5HUmmDCrzEucwgCfq+NIBuCJ5e
rSl07hhCCB4iYPreWjw6BrS/sNSo9yVMyH23t8KqVqXdVnGnhFZn4MvQv8uR26YktDnCn+0NQwhG
95RerUW1bq09B5PmbiTmQSpEobUvjiJTnp/3YYpzPJZARHRSJhqbjzJ1He3ygi7E0fMI2D9C++6j
xXAESF/Mjq+9OQU0WlIk38hoUZqCz2AcpU6pAr1czZrwsQXZIBrCfPZJCD0QySnyEuNL/oeqTqc4
Ubdi/su2yfhIEaNHPjB+Psp01xRztZR11STZwNXPCBCGrEHfTSr1/XFp9Qsbto9BhreKq4qBe0Qn
yAtnOK6JvNJNeVaZBA1ZdJFq1SL7pRimjZ3NEoW/oY6l3Z/h2tAY1PRxQRqtEtME6Q8o+Xhv6cl/
DlpRcqXFiNkopQRMt2snXcC2lRQ3pDzKug+QqAejxVihZfQ2hmA0y6/OCHYkvD4c4NFqO8D0I+Uw
B2jnsFsaVMmc27OQ7LyyzMdsYlSDpHkbScTuAts/Hpl/04MCfHWV0pYHYgrSeU/7NTansCfOF1Ng
3YQYhO85ixFAzYvwEE3DiogQYnSNggNjEldlFIcKScCaOHYpGhJc7Aw22MTwg3AVzJZwDKH/5cCr
T9l2KkCowBLgL47ITVBKnyZnk1om7KMnrv2apU/B6N9T2SjfeGoxuPWMWeel3Sz+8XNk20lN/hhO
lGBrdUskzZNKp/WMr4secN9ZQiVrccbvY/YTT6Fa/qldFLkFkAVBAuXo6V0VCMTmV6emXk+cau+T
knsdlhXRqIZAac29XeAVKngOONTcyyGZ38E3KKVbpm5UAeomK5zlu/lnsRQVsNdjTfjiKzENuSLZ
yiB0HXnL4BWCJdJCFbU2ASLmQqK9BcKvOynkZCsscpFDSp3kXUvFgCRnMUuFLuDhvwoWZWfdVkCG
nSwo8MNzOTY35b5Rzc8di2sby+ddtYIj40sMMlBqExPLZvrnW6D+b1a/kSap2z2jZWB2X0m3Ng5V
tlWKKncWz3vFQIpXQeb3zaqe/7vRqX5uC5P4Tq5nbY5cKcFeCdCQkdwcaYWCnEa4/jVsZnk8f+pg
EVj+6m0El3Met+7Gn0ZA6KClyTdvWLvQom+6dRaXPfL0zhBkJA69t5KAPvrivqJ9XdiXUeF8lBBe
r0KgueA0P6LeaKYekU2KYCI83YBJSkFGxo+6sQ9+e2uwR/eOG0wTeAYfCjJA6j9QCsfxnJKA4vIz
LNqihzMK/SSiBsWzM6AmWpRp3fHcyJYAB8MZgAAueFwEn8l9R5a0CvtTJqAS2jCU0fTSNxE+aVsE
PsEw7wgkLmi1a5ccSLtZvq0Y1fCp/+8iLvGZNzs/q6OnYX08JOdkfl08MpspAgrEpPBa2WydgWPn
r0rYL9/US6b/CDR3Eu8WouIsbgHcPXFsn4D+lYjMubwUUrPm3n606jAM7sJqY6LPEhYXc56+G+Tb
h3bGjr0C0mpQuzdr2y5Utp30n2SvQEKFwtOxk0rO6ePJ8taPF+UkPwGZZkt21KOovmZmRfBrggNO
hzWDIyeRpvgpMujJqW/6P4Wm5jeEPAmbhscs6Cd71p0G/eLXmqq6Qkc2+ljmGtf2KoMYA5qdhwms
epwGgGQz+ZehffpnZdNNWEeCSNh+V2d/5t/jJGHdkO5W924Sai/TpL4Mkg2u0Rs8j6EqLhtKexf3
MDGuLLB6sydKzCbiziLH+mn+7npTKfum5rw0+G5Sx5EK8zfflARKoToOd+kL6cQxREyRtg/ROMwt
7e6D+rdqJGZtE0fY1USXMj+XQklE92sRJEnuskPg+SrsoCqodVYJxPqnjJLH/0N1C+dbJE34jhis
KyELfFk8nYgE+nWlExSYsi7LF5lnzasAGoHXxWhYv9p/c9AvHvlOLdgI3Ei4h0UyuOHyFXffHgxS
MHPYlt+C4s7SbdtOsg7+OhkX/D5SQKv5I8h9gC3rMgD8Iou5VssM6Uh8/vJiTOvTF3J2sXKGNjQ5
Lbx97g9GmlE0F0dZ+It+pDGxq3XFysRbLfwNHOB0OTdHDcnw0bAVqqqPUZtAy/pCK/2gwZXYh6pN
SNGLZgf9ukKTq2soZzWd+uL3ccu859D0Gub0D3/h0iyXJ/VVUVH4kXnvNpBZfOKS9JJwNNZECRhx
lI3THI2qrAbytCDMJYLHTnpeSg+eFuXrxxVYLvgaztdk8olClQkmEph51/82oXPurEmo8P5EVQGN
uCy5gtVdfOck2Fpscf9gq8UaC3tsKgnQqNypPRicO8dftzdxxNAO10BBSLc0SdmFLjOPR8NKCahX
qqf1vPGR3knz0mkAMH9IEWcOdqqxQBDwHFkRNONg3rpRQC4DLOvdTeu5kgK/UujGG0hHK7/RkePQ
qtKSa1f+vUb2LhJGBG51PuEQSNsuPU3KOf3fdpwV4ayWzelsCsdzKQ8QoWsjHk6Fkkhb0gzzrvOq
mV3Gmnz0ufIMc8UoiwTElRZ4amuHUGWWTRObMh4kctIQTAOOejqyw57pgOwU54jrnxVzWi7bO0go
sneGW0WQmsBPzFVf/J3Kxy9w0NxZD7d1zN/khFAAxds5ZY6YqoH+ZkG5jJOh1DrA8bTo4xVyAgIV
FPlq+x8/KaLdzDxLAzuF+FJojDIAtjNsSDZt72sev5W8lLI1SH37DlPnB6bvGE3i6duIVvOUxF61
0sMJd3xvd+1SmBImQDx3UykB5l0AlCzYAuVgPap4VzWTrJxpA4POYZCgBJh/ERGw5/pDXvlChBhB
BXfNYQGHKYvh0WVsvuYdd47cMlFQp//qQeuPrr337bZmAjLOHe4QDyEfJXcjZJwRycP+9hI26Zb2
0QzDlVSxkkLZYytHA74tO0PNlmShhlA3E8Kj100QMlcuIh0h1IS42kthFR+cRff9cu/GcKV+5j5o
zGdss+lq3iZ7vVUxe5B+RRC1LJA4c/7AX9pGQgdsBTgM4Cq4vPX5sEtxVnEZo/43vpKI09n6a7Tt
ipl6m0Y+HgnjH8cqrc6OLOrO8/yIVXg6ttA+EO9U1BaQXDxy4MBLi/fVTVTHET/oBIJ95+K0qwNV
pw6Yq1IpJTfDsSLxSNQVeANoRojislapCMcbBuEQ5hxp+4YgCGXJiLIb7t0BUXAR4b+OkCWKZ9pD
VyO56S0e/Tmf1lj9poF8n2Qt3iNFAH+PIZXQxooOvRm2A2WfGxPRIInORNXcPMOIMLD9LQiIVU+N
1CmIXnuOTMnz9lK+bEYypllQQE9R7JM2iR5WF/8Kao/bFgSiWW/N+5OQZU4FNQGfg7+JKv4ELyxl
fMY4MAL7Y/Yq0hcz61sysw8QU/bBbmNkwuQfOyvRXOeQlyRwNRTk3mvtfDd8EYFqfLDcTqHSrTmJ
BsocuPrlJ1ioL/I+fq+OYjFwqzLAFb4drXExYumO6B5Yyd32IuWWZBPyJa3hbU3sC2ZQUkoNT7M1
5ZgfzQgL+qfZayKTzE9WfVJ3KXqRPOKAnsPsFRQ5syD8PCjmrGp9LdvtJMxRVhx50MBHxCYTErxy
sCWO5vKxJ4ukN9xDyD0fCtOrZ3ftBcA3llnayOzXBXhil0llV5QF7C8j8YDp9FNn0KvMR7Xh5/9U
kwUWvGN/SyYSMFte8ly2ta6in/Lawd9i4M+WrAXQvNXwxWlkWP7U9aMM3uGFnlAzwF9ZMfOD1FF+
HdAU8u75NrYVohxSVlhjSL4vUELhAbef+5xf97j+yJJ21BN3jGvxSW7+SVRi848ikyMKTxHvyiK+
b2ss6wD3e/Wg6EqjD42d8nDiWV/XxUcwVxAG/g35567NUZj9xqkelzuUCDqvQiHAuoGfr3jdsgjJ
ILfq9eb1t6juM9wquz4mHmLszA70XYLyHs6QICOUIkfyPa3+eyaeIlaqBqj7Cb4SubS/a1b8nv43
m2iF8Sc6J0kg63iRXh46bWAFP0rt6WR0T0Fqp/UkoRVa0o5/AdIh7x90nzE6GPB/9eVu6Yl+uyis
v/9yQ3kVrSahtQvP3qZRS3Ld9QOPzToSxq2FRFcO9051x6rt/JeoqWFhy5Fy/JT/snmDc7cE3jVK
gJTM0pCMsa0q4QVKScXt6gcOlMCyBuVgJgNvcQ0h2knMWaQqEBKJ3lDiXwHxGE6Mb3L7UH4QOFU/
gZp6rQty5UFktkNX07T6BDMCzanfS0mEHmUhs7nsi1Ra487NbFTi0WxDZrpGaLVpagr9qxIzcWcM
+JPVOcNUVHKNiIU85xHjStH804PEYppbFR3VJpTPFWeyw4NpMBgDDKY7TnjO5nLrYqKsBC3bkPpJ
0eIOusmenraOonEs/GqPyG6X+YJtjZE4B3KaJlfn4FqufRwQOWI1UhdQFrZ1zgDXGoZaypKj5fI8
2kU+Zh6TklW4XClEoEY17AdghC322zdnNhH3iRHHcE4huTk4uj/tyYlEV+SGRmbjCwonyik49k9p
rLb7VD90+QzQ8aQUxNvZ5My6bHUU54ZD47RT1xkaWwQFvZv3sQkPkONjVEzRI88Ghyg7EO6CwRiJ
vCocefbRrulJATFURd4MyVyqFE+VkZMnnRfOzZh/HKezdXxd7hsbIuWvrhFQCQRHer5+45vDy3pr
BH2OmV92Y+yl3HF7aQflKYZ41EObnpr/LAX9UsgUq2+mYhpSISu5QGLsWOFVhCMROLeMdd5CRhZl
houQrtelcPNRSv5TGUjpDLJCaRFjUSLVfp3+Pf6tAck7IDdt9L3UgsCSuLX6KqSXvlzYYkM1zuJi
cM2esIz6eoygilrzP45phwCnaZCQkUl4T7DPN9AFg6PN33p3Vs7V4pFd8vQ5NWhaQ9+m+r4wpomi
C6gUcry4TBHlevm8SPxGl+07rKPRQiot16D4KnIwPnyg+rZChGkAQfMdMR9sLWwzw7EtAKVlKHo/
HeD3Znqw9WEjHZxhOEVykr4wdDCeOS9J6oTkoyupp0SblADtI+HNJ+cV8NI7j7fLywE7l7RrG6pC
BcVd7m55eciVhFc6lkwGjGl6i4Ke3dilJ0B2Ikh7n4Od2E4drzff8qZ/cvOV/0zMEXyFGjSeTrMZ
rcA6T7TQ8kqFwC/Xn+FBLu9/EHK3JJUfdirtqVdIUMyCQXw3JYtBbsAfPXhpCxNWwlyRIcYWBhXe
4bdQrAOFEqh3J9wilOj59+XjW89yozq17TOGuQseNqqOb73FgadiEE+SIMdGQT0ymRbzwIUzP7Qf
53dxsByeDsvLbyhy4pRJpBWxVp3Er4mJmnc52NX8Jbn76UuHBWSPSrp3nQwJLZix5teJxNEas03T
vWqvpPkKJBVjJqGe0X0zTkbG+zbGWAik4ItQk1Et1kedBbo3pC6brgwmF7pBbcjWqznqlimSr8Sm
qIM/h1cwTcvwDLq3u2XE3U0boZ8CfhQNyX0XJtaqcUmMbPXwn1l+Q1SFxGV0Ipfa/Y6hURv5Q8cX
5fQUt2oTa9gvCMhPPvcihW6E3cJaiCpQIM1RKmX0Xl58ap4l/weh86SEJF7B3LGKm7Y+WzHTLNdu
lrJeD1n/UV0ufTzUdXtTkIFQljYZM8XerEiQURsA8oanrjEzrgXl/9WFQxOU0vZ1iEaoa9d1q/KX
0mwjQ7LqJcU0isirfIusoLngWhC9zC6+qk6TKwB7OGbKVrQqT9vseirKVQCKTfq4UXBJZipzWSt2
EoDcjT7MhVgCdUaC54WVETNCPeTtCdzgDxSS7YMQp9b0Q+Ccs7w2YHvNzhmy+MWpQmHfwEo7k4EO
ESTbrTcFUCqAAQV6n+IWEIqQHdDKhpHwjamKaD5aIp/HbX4pXn/AnZ5vJB7dfM2S5b2AU9nOlK4o
ltJaRMo6GR4/iBpurfq0y7AXsRGquW3rxigTvO2DisLRqXzzrtGfHaH6BdCO4+rf3jYuwQlBW6LG
HGkZR1V6IKroUjSJQMzHcgRY75O0Y/r4UjCPC+NfNNFNF27WPE+e8X6mVOHxMQ0zQ+sIE/Pfzjin
3WP5Slh3IwOX8c/eKTvYJ3S9DdOZrVw4bimAzE7RpAuwwZf8yDXyFrcdWL+wBY8kUecuKJNsOzhc
L/+h73+ljhqUxTYHUx4ZoZ/GFqfDTnXaEOjLTF3rchTDteLPFD8wo+htcUr2O1V7Wtgm0wXskRgW
UPO8xgIFytg3ze3sgMTzgsoRReL0obrtK5osnZnNtSACIGZnRnD74SdrkM0amn2nbvEtjX6W1tMT
Jy1pv5QQWvZiUL0C79m55+cRh7aFoFsvMh6l0OtT9X132lXWcUnc+CGGpszfVb4q5cM0C7XXvRj+
dHH45UdX4J5+nzD2KLplSwNgD9KNdwJjmHoDnUYnB0K1HRz6MansZVvlBEkLEvC2/U6st23TL3Fk
O5V1OuWqnTz88QskjgZWhnds5WAlSF0ESWB5GlpwdkDF1QTxmwI4mqyFc9D7kbypZRT6x6guXBNO
kzUgzgaqtdPkRQRo7c3MYkc99nGblw4qSg2+NbUhnlqa8KdeBEr8bP/PPcOe+0kDEvA4vLpO3VtQ
K6hM++nyHhsaYtLnGqzbRoV35iySFYBy4j+xmqaDHJ5qpr1MmHEm8Pq6qyI23SjO9mPCk3GIP8JE
8CITNwCG6lvfRnkLEVR6LYSKEpFT1TxWZ9E7JMuQ/X2J6lnQQ+HnU7+eziMEIz0xaBHD1uwQpruf
r6H3fgkz0en3ZT6duO0aChjOKufuHYdeTUncX2PD9YPM1mqu1k3I8+KJA1UzKCgYb6UJ4QV+KbJP
MTtaxhJ8WmRZFwyuy60igAMuJUhfWjvgzGZA63rboueB1eOL1rmGbjl68Usny1rxi7a0NuQFqzTU
aIN2vAZykYPF6WjELwj8J6wFh70bZmDS9qoBxCQ1yvWksH+X6uCrinAjEhL/5iFs5kYDksfJ+cyJ
rrl3pu4KQYD5cSM5vfBy+0QrgANHbG2oMrvxglNyIR7Hu5G4CvJjssuk5R7hG6GbfYCglnKKwach
3M3VNgFMHti2NKL4h5N1N5oH7VtbkOwWNotpmzKhzZRmRZ2YVgj5b+WTuzokZjo/+K2FLQIPxgWv
UUWAwMX2JD6SbPpYd4uQ3vX1LAw1yPLqN4yqKqSG7NBQWrcxxselhAp8oiCefksWIlAYeEnv+3db
cDb97DgUZJDil8r4VB4jqdjl8Gf6WKKTxGZvKwg1oCukmtf6spj5wQ9pqiiQ4R8PtogK6zpxnsWT
+j53hP7FIwiGrkSVyZ7a2qm3xoY86Uyw++GHUrflHEOeuqy/ProsQuV/yU4kW44kop4LpbhcWake
vPv6406uG/9twVsuUPcI/nowzZyrAuUk6JBRLR4JO95lFxrxKuc9ew5noiViD5o2VkbMqwQRLA2E
pP2+KTEgbajtXrQZVDccqXNhBnOpVk/K6AW8tqPLC70gTJa+xqQS0s6Eq7kOrmf5HwH4UsBl2fMm
pJcoFoJjeZkS17mPqk4mnt0c0a5CCijI/Rs1FHOLFOHP5iySfMMB0vpEir3a6lU1gSlttKgdu33D
UMOtNyqniizde42PSIly+45eBCT/qOBY61petMpXPPl69+XKWRhuWlfaVykAmU5pzWcJYDG4tllo
87OUj3LlcUFhgS/m5mL4pLN1GmPasSQ0AjwNoCRmons96uv16gno0Hio1vAOVlG4A/oKR81kPzve
zbMg5pu4Z4cQ0XGFEicXgMfZFPTrjTgusMqwXVFhhtYCy5TSRklTHSSbGUQTzxse4ccNCo2laI8r
QRtpGKi6c1jRaFVu1H35wFCZBcX2DZB7bDBxvfagI90CZKxbhvmoShr6BSrFCMrHPmaEfCiJ61TK
ytfXzCofBpzY6VlNAKXt7pqZzBDMhe9M1isX/4/2FzDOclBA9cU9GqnukTdbr9QAagPV7j9CbcR+
kK50recZq6vfUq63o7Z7TnO0cbHSJSyUz9CiIX8EXxrhXY6QdfsRMRoKBhtzgzNsoPMjjOO35XtV
aXgpyqJDwA/tfksupI5Z2hgJhzqeHoIP8sKftos4ylAc/9UIy5YkQpalB2Ajs0O3J1ymVWYNjlpy
GoqMfKj+YTvIGS53ais18PDlFmbeAK+EHFRwtLFV1mPoR4+3FhD4Riw9eYSR38JlIYQcrAElvdOu
Lp8Zn6DmRJKCHIrpZR/l0i4jGlXy12oXvWz/Vco1j7scjmYAWX9Q3QiLQ/Bu08bceN2DpNEfo1OC
u99k1IQB7gw3ZN6M3LSkpe1iGSlLah65zKmqKpin9Fm9/Dbx4oKY15TawNhC6epNLgs7LEvqx1vD
5wGKpTu9GRR7uPb9lYl7BBhDK0yFmhvgDdWgYN5gRkPNIpRTuHfB861r8HnsolQd6wW+z5fjpkCQ
LflYcS0S1xz3gYpNFIZXykf8UX4UNdSCy1p4C9lFi8R7OZB2cxXpp/gexLQwLYFCrv+Af3jao2Y+
V/9Ge3z3lOr6FapmERcEw2i8iTVd98Gwiw3EEri0jeCgvA4ecPIXg4+j9O/XwjzPci0QTAkhUt+E
wGOi9PCsK0mfGvYvaMlJCHP7Wm0PNqIne+k46L4ry6TLxMybHqxtWhh8xgYOmwOmaZGQ0o0VAY7o
9TBDod6A70zONdAXnc5Vw32Vdi2GrnVQUxdu8XmYeensVT3BIFeUirILof+97wGyn4wQDxTSfKdP
CfFDDljgx2k3tFF35p55xOJcXT94gkRaBNTfUS6ObtIdyiVf4MWNjN5X/+f7KtuI55svHajcRfJ2
FLa8si7QBDJY3d7NNbeesRKMBkFcvEFOnVEcwu2FtX8b6dhd7uzSHHZI0WfkN6JsfBqK3sVl2jrw
MIiaq/3xckknA3tqxcmmy+U6fpNq/V8STQQjy4aQENFpbra7tb2FLDBnL8wVULr7z3QlRQJerBNz
/Pa4XobsqnA3Jkq+I8Zsdnm0JiuJ8a3/oosfB7cvud71IezKdNrd32P4sjQYpsl/emHKAckIznUP
zFoQDLcq6Bpxxki72/yjNnOQA8ABYbQ/X3EtY/b7IsW/Lvpb7UfwwE8oGh65c+Clii+7UJk4RF4+
E9icsvJQWRcsWUULTAG94ITN4cQON3DErDn6+1d4j37/3BrU9/JAHVF7aFcuEqfJYZA6bjnTMSfK
F+HsFMbUgwM0Uf4IqNxDAQptLdvYAsrvtk9SyjPJndLmGcs5+B5DUlKiUil1VY+TAMJ9xGKAkNLm
SGI5K8q3opnolHgg+J98f0UY+IECRMu2DBsGlyT+9S3Cp7i+pXauwtElfZv6hB7uVJ92yu5eznGo
wl9EnhHGN0jzl18I3w1zzEPXg4afB4WBkdLj0CmwSGrSJezD2eguOM9M4fdC0R9o9HZW6nzaE4gF
QmkRzl5Qpbe5qgUzm4e9q2S+RUsbScw1a/S45oTsWRxFhUfxTf2XSQeV4tmmkuTtCusJSlP2HdgE
NrWiy4BVsKfwFk8nfBOqV6VLBikBuNoFWorCrpo+W6yTdFvUm6gS/+Ese5aBVkC5xWsMetKOaEAk
PaZPVM0UkbDm4Mz4LVl67y6wN1ecfaZF8yzYCgmDL2EVYkyqX/hdIAmE44SDLnluIU1LO5Tv6z8j
9gi7m8MT06n3Nj8TDe5oyjoCgeZe5AV0tvsboy7ApljtR9KwDE47ajrbvau1Y5rt1b978KIYm7Ug
P59MmO6/qzDreypbWbIzbvSOgDI2fa0iL8yKPFJIPD/Nys7oztL0VPPv/5Jt7sr3EFg34XYCkzsX
So4nLF9LCzggIXTRqnF5yeHgOrZxLVtwsHLHhJ0MDbKFn6JMUZFQDCtT32LT+qHB/5mFRhfowD/B
PXd1+yHdhaXFIXk2xj3CeGJzV+0M2RXB3JmlkA/vjgAQw036KXhZuQfQ6xkB3Y2E89r9uCjlzCAF
ZaNJmiqSoquU/lnEyRSgLpxwlsHNlRKSehY01+oLNqlJRLuOowVkJUiDkG4x60ylnSZlPvsKg6+Z
BxbR8pEY4OGzBTDnyu5gTZxcHtoE88/ecCZJsaDkgO3pgBszkMx/+senmXBF5dq0Wn6p/dyVJVNt
IZj2qYMwySX3k9v6e4sc1aZSbHHOW82M0TriXI3JrVo8/oovhmimGxdosPPj2pT984nTInWYNDqo
LIcV4m5QAz0nL9PMQs3quzneG/3x5gGtaQXRBO4pazGLqlbPubS5Kq+/OksyBqIEfQCIkv3B4Kyp
yMi3PhngwBzXmIos+pKWO3DiQW9EK8vL++256/hzuVL9rrdi6oyNTIIlo/qoHnNQZlEmtZrjDgET
n414V76135tOjjiuUkQPx2mTKkRfqR3xQK5qF1q8ziFAWMFpnvRoTkYMNZdGzj+9YAVDcxHusJnb
q/bMLxlsjs4XysSdB+yVJJknY9lo6vUZpNWUvjbeWyMAhFrQ2uu6MXQmzf3yV1UrmRum3lWQIzzh
bLcjKaY+Tf+DiA+vCOUSTlGJgMWVENNrge2jQaWGFnEa8iz61ZlGGcaUazqddQ+io00fKoMbSjeK
Wuphq8da9/AKPPF6Ne+WmuFK6JzShBBaxwxtFQYpAm6yKt44iiHm5Hh4MEDMRH+RXtBJNDNyiVSS
JiCy74/7d1eEepk4NyBpbXpn2Ztfx0hZu/H7TQqjhmbz82v9MBn8wZltI72kKJzo1CZsByCozNGO
Mp6rWTzLmTCeZZ0qCRgWrKM/N/yeqXMWhmYFCH+JBBIwFcS7V/+kbxc7KqFYNqEpwLXO2Svoa3BK
R45IgWlVlNYJl96F4yjK7CuU6rke6Y6MfCF7cWpVtxSVhn1N5Jian9xgPc5I+Hl2LDhg4e97e3nO
6KEl8f9K5rXuTaAziypRZve8q4kIZ05h6ejTnzFWC2z9CK2XG4uX8ZoU08GWCxMXAfpi2JtZ31vS
hckfvAY5zoPZiRxmAOgPiWXrlAh/Dp2w88r/yfyPdfC/Ep0NyaEIrC7YjVFVVMWmdz+CpGp4EfWc
Z/1hSvvuX58/IyvHsG/HJHUNT7cJfrxUtThSDJbLdkkc/pWrVfinw4ZYgROMYRZ3AU7xXkD/8aVk
LFPh8ttJiVHRztUrazKeXRHXu76f1pQ2y7gJi6bzyt4bgJ9E20ExQck3ftPILixVQ8unwhEmGA+Z
1vmYXdBEB/3RddLcW369V0O4M5vDz7DoTJkJQCKjzERf+tLbQbtY5fz3aZpbAkG5YuQGfBHGWyKP
FWu9jzS1AT4qhv9XyP/VJTpLTFd4/+BA95BsuVkNapy+rI8KPdzmuq6o0b+XbwZJxI1JGAsjE2gx
omql66/K2kBR9mkuLaYTdsPsIVEmWfR+CxaalwJLr8GmlW/tM7urt1kNMo6V2tQeVbPC1UfsO548
QkHr3PGdTG7PW0R9YKmjfQj9Z7Cp9T8j5GwA4vHpf0o95RVFqLKwlFamnTVnkebaF73dAq1E1TWX
Miiyvx7DHfLQmYJCpWVoEzyclz681xzud2grqkqzbB4I/1ad39WG1FWsyWOCKQJODzeXQHgj+/AR
dm9tBKPH7NaXpEdaRr/FUVgAQyqkMfYwuy/JxQLYUgsgxV9KLwmXeyOp6nx317UO9J9+bOcoxN6M
m7EMYwiMFDXgBvacssp2MGmISxl8P0egGB49QElDjgpJ6NJ1Ah4fRJDKQhb4xBSY1JZdo1Ut2R+P
fljQcIO74U3HU8aAaE8nscKcACQvoEjSzGF15kt2qqF1GHnEP03WjuY59Ymf5kPT0MtkBgMXlsfO
CeOS1cNrzh55iVsi31Hk/8mDvBBKgcxUqjr3iPFPpp72iHHR5VOrPgJORYxvLhnQqOtDF0dgnDR6
Oaj+DZZWcxthlsGm2S0GXdENI+BM4L6o0fuctGk6BQaGA6yo6fHbg0P51eaEdE1FEFExo0BCvzgJ
BgSEa1osNStQjDAN2WzauY1k3gpuRncCUrMfKU8eiUtl//DSIDHXG8xCPQC/qNEGI2rgZPvZxJTz
KBnV+9u6BmYsREZcxZWOK2fEF/Zm/KWOoLeh3KPGRvqRtEsLFZ3nY43+R1d2p6hjCGudEbEZL+yQ
fzyI3wqSU0BJh5QM3ZpAtsdA9QSOp8HOoTY/8AIAhIZiJQWcAaqPKxZIW8KVkmN84EBeOhj3Zk22
QsVed09Pf9mdBoiK71JwnyWUlSvP0dndL+Gc/hX3LF1CP860Rh9ZGyzfkKhyNWY3OLaqEXh1roDL
CFQdmWvJdnJIvd80KCuS3fHq38scaW3cg2DwvPh+1X1rp8hYlWmYV6WycCHh1kUxqjzY/CEoBn6L
ZJWgDKvmWObH9xPXNhq9BrdD69merzz+NdoAk+c6mrKAV3LqYtMz5VSZcL3paThIjWjOJSv0XCTO
0ixvPf90sSsdamOMNsKCUMFA+fFwBi+qT1h1XeZMFpfRiBsT+HmPqrc7qvEMPpACvxj9xdWnY6HD
z1xOy3TsCzJITgChyX/GdVLZO0mpjj1fEbbVmCk0ns2k8kFoidrZ0wsrDHh6vGJZKKHu8umq7OMZ
SBpWdpK7Y43ag857PHMy2Enkq1IQfZZiicUQxfoEbLjYLjCai7yOnjOaJhh+GGzqpRcgVWcwc5My
gH7DnWUbcpOsGsERpwW5n2NqORY0lxqKO/Le64dscycUhAnY8wT2XGQ+6hFwaeJvo4p/1ZBruWi9
3sHN3rKl7+jYK/cQWxQbuy8wokDHNW5DTdGDkF9TZA02eL4YQlDxN7ZmZ2eJ1AZdEdnD/1NPnC2A
4NKa1j0Tr58+dDYiEI/YHafaxbyimosTk5eufJ4oZ5diUUa0N+EYV3sOtkOiBS69GbMTd6cJdhsT
3ftxciCaFme5EcGsPtZcGxXSGxsWnk3r1MX9OD3csM/1ufBW79mmxf4REWf2+r1y7Aahs2L1go7c
KCcZAUY7UnQGpGkKgb7f8g6QcUw/nHV14qPu+5EAP6djeuBmXwBq4rTcYhE+QpaIz5DpyYDBa7Jv
bUURyt1CVEdig4QvGb0HMlWYvtr7H/VJ/vx/Ld5k1hCtJC9qdeVHGNr5V7wzWoMgQuyfzH087Q1d
3fFkrg/HtLRGI84vYB9Md8MbqGZofLIJ4jN/4oGsrfqcoqCPsIjinKv7Mz7QODwzmIMSiKnNJn+/
wZSAs4/QpQVDZkX766IyHdqnkXhRsGWb6rf5rpg1gJSTjDx5D8SvMH+/rih1xSwQJsEIv2ZJQ3aW
/B5QuoAgGIfPhC+QqRXfr5Ma3LCTmnBcadEJwgAP7r1Yw4tNBOj9JC42OK7aclKx44aAkYBEHfQ5
ysDoc/PVV93IIIukgSSweMjC2Y8+WR/DzsNZyQNJom85a1LozJFMD1T3WKWJ88woERobQgaug3l/
4zsPg3hxawa/0udomwBl9zETuGXZ2Kt18kK5ahObIfN/aUDlrTwPYBkPItI3knJFpyNUpcD2E8El
lghx4zSpJrct+3ln6CTmryrdpsR//ISjkI7NEUeSIHnBLO7Fw+2dCPc1Q7XFBPro35iNhcamVzyk
WrG5cpoSLRJ3k5C6SlqnjxkjrkeMDGtfoq9+a2CNYMfgCvW+DIxSW/ZRFGQS2i5736zZ6C+yFfEb
TcSPaJ7AfvEOSloF5yT98xyMzyXwGc3Tt7MMbXIlSX0nv+7A6khzP8UCU0ttm1DudcpKZZJzaL2d
vISKNUGyiFcvwq0I+Cz98D4DF7NrwRZjIBWcsC0CPUU02kCSG3KQSTE1OzhovARUNIR9co1RCHcO
cIrCp0FbDgzro/TdtuolU0+rDAOF40BHQ/91mgI1R5kBAjMrPqqdEJb5HyboadWFQNj4QG5o36vG
4vj9uiLP7vxAoDYyaGn3tcljkVl9vFPLcCPLk53qLpERLwpYHBqAsB89/5ASddLIyNBGrrJBmApO
IYFU9+zteHutxQ6n+r98gannpMdAHU0z6wjYp2P3c7wZH0vlmAO5e0i6F3bxlKIXKiLVRrKlS+mS
iIpk49bp5ZcWXeaRRbrWDLF/u2iK7hJgG9FXQ/V3UZhACqFh33Q77d/edQCyXgr6TooX3HE1DJ/z
xoaRaOAjIkLiDJ0Q31OJKBFrM6AA4k1saUwDB/L/VDVpRYN4dGU/nOT1/f90A6rHDtYWG6eJjAL/
4Hqtx2dR1qLjKvrxUYA5vCNHkzmXMo6MHxqib4ScgTI6g3y7qp2ol/PZhZgTj9LPDv+sLJCbA7A3
U4fhlbNt+aZA8WFVBjYwX12ckrUXdPBAa5lKyccnh715L/6wZGtWpWTE/SXNxN8NQD6hfYwn4lbX
5G/POG/DGxj3UM81BP3QZMsNVsf6H7LU9kEx2Homhq53c14U7o45qVilxOB81M+DmfyrFVtNkSeY
ULnpl6BHJlmBEMx2IqnI85sWhM3q5tp4YtnMdW9RAeWRvrn5VHsKRcpgnSPCjpw/WN0Z/kZAtLEj
gSwMx8gIEit5SGj0+nBU24P1w9VoKwO4veHt30EbHG5JUq97i66KkFdTJE5rs2E8YyV77Slzyn6J
uyGVOcX78GXKBmxog3b5G7K3k61Nn1r0J39Ky75kTclqkxKN57LH/YPQtDPRiXD9GPKRLZcEaX4b
/5gdGoKCwN1Nw1LK3I9ezePVPWnbeyAWeqGL007LSJ3EVLMRzutS/hPllBRA53MF28VnXFZe/FSl
c9nKa8n4XgoCen20Mm+ipO2ARDhag+jBjqXnEdGME8XMIHg2oUj53iVc/LXR12mv5GjiPiJ8d3dN
cxob09RyELJSrzUEJZTMaptaKLovrrQp/Xo3bzOOhHHPJjT59cRixHQNshlOu803BApH1rRlCfNP
6ysEISDQ6ZMTt/vGNRkG0uXUOl+PuaPLNz4D4zv1hwF6AXWdr7EiH21ErJqq7NGd12EVFG2aiaOu
ftfTX+5N64FEw3e6JQVaPaicIAmZzVJ2uXwCCaaOxRAflJzF1EVc1G8c+UMvljFly7jonxW2+UaA
7ckr1vTiBBglcTbl8Uh1jE8OdOez4XsHuvVl9lCS1vStJB4HE+FQ79fgePPyxJ+PaRgLrO4uDEQX
gR2Pk08WM+TZ5J5xl6cyW0KYGJ/m5pkLCBB2pg8ojNPTrTHVFfvqrT8T8N6Un3BNiREDdvqerDdO
ngacGFb32vp/SLkoqHLyyn6dZSCEINksziB9m2F6o8/KTeWkhNG3XT4+m3u4vfFJ2dC7jEJ0tRRb
R2x0ch+k6HT40p1TlWh0jRLj1Qn91wv3fAwjyTnBRqieLegIKOuH1k84Fq10dFT3N19N4yLuGmm6
6OI/SsweNdBowSFfoBhrAN6c1fh/wksac9b+eZ3lG2ss2RGCWr++MaFztEH1VQu+a2rulUur8Q4E
V6/T08jRWlRbWkuB3BlPQEwD0IFwulA+5cshlzFa1N9Z4eZOFshkQ7Q2IGsqvyvdUO1R8CKjetTN
fdI2GnDfFBjyhs8UYp8M2n+lX3xlkl8O+Gbi5JqVJimrt2yGP0KRZY94qm8bw8I8iseW58Y9lAD/
uQkivqJiHTC48D1+JC0HX6CU3OiWQk27mCVij0bPF6JUxqTHwb+HqWzPJpqj1ddywS4J+RU1tLkF
f0fqETxapGI17LX8jqC11ldajJCmESRvP/DSTnVUzWRWkpkomDhBpVydUiHg7p9Z9Vba2/Knf3jA
6d7jPGOcU4p7Oy9Km3sYrpJJjGyF14Df1t9EA/DBxs3WkeUpXkI9ZhV1kXgXd92HRgEMs7CRoBhy
Fk+wRvTeXDJiwyJNL4BT2OmfdrfuObxMm00wo06veOdfM/WuRiS0OLjiaaGxevO7DE/eaqwmlY71
5Lm/wOPWJmtBa7I0EhCs6EUU9k74FXWhEwXoqscR3UrOqPHIPAvUKvvgo4KNmvRCIRrSvQMuZb6u
mPH+MBSxHqH0ghJ2ntAM6+wmD9aLtr4XqNo0xeKR0x5ZxRofY6r/79nQWJiBKwebo5vgNY+N1Sj8
2ckcac/znqxBn5jzqca4wv89xOscFwRafqL7/eTiQ9uvP+y8Fk/xH/BLsvAqM2W9/0uimowyotlY
EkpHbO96tpBNR52yyyD4AYMSrDAOqINHnXuwVots9NdfF91gSXYvx8ucaVso/ZwOBTfYTR3CevtU
J5/5C3tCGMVGA1PEfwe+TaRFhtXAMwVXauM3QCQCI1C9kMkIyACDYkl1HaGqyCpcn7CdCSnQbjI0
rbCmlysxnrJfSfGdb7/WASBTdJeqmF1kerPmtKFfpqRFS4xfbwu27cORkwTSfelzxop11kKSExxv
WBqt3xjKqOu0hwew9SybkwbbuP9X+cYc0doGeO1FJyN6Dn2sBsA6c6Ow3jEuz101bNgJ+FuY6dcr
bI/+TqCMlnusQj0cnp3/kwJB2hMcIue+MzpD1CFReQYtqrRP9QeJ6Ir5suGj70NNJ/9Pwy9yML5L
TgBPJoNzWO7zGNuKk+COLGp4Tq3bW5dQTfh8lCyaTnbngNwrjdRuVMwVkKd8vLD5KHThJdlI++ZZ
EjlYpHh9aj8MAfNgNzhwyy1w7mhM7hGkIW4yES2BBG5SMbwso6vladliXi12nZFj4zrNBTQ0ZQKz
g8pNVo3PByz00EiSKIhLstL2uVsGYPxupK0qwOjBvE5wQ8PojvAjEMt+qcCApI8ari2PfQYcX1BQ
o3ZfRAwt1pyHSExSvypmuO7hI9BL+Vp0Tu4Q+tF3gqep+JF0dM+Pjd+5vbjoYAeD+vlsMdQ0yaqk
aBZ9tV+kEkKTS6UPir/r1LnD4YadTJXBK6j0qNe4CbQipTmcPKBBwzU9scCpHG7+op7MMjN/Qiff
7ESkPlavQHYqnG2yzEDmd1G3pZfo1IyPVdQXcWHy01qwc4vdCGVS5i61YUVkJB1yU1PbI8vDexbN
cpC7GXDnhoJDwPClEhWMXteTig9BK2xnrRSxL+xS98cBOzAYTOz4jgJghyqxxXE50Q0UoleEsBOH
GThxmJbvIdqlW4DBbcbS4SOGwaTzTERiwMuVvF/WTBYx2hQz46/a3C2k2ycLq8YwTSEzgAsBthoi
2dPyWOpdrnkzo2EeKxeo34tftOXCrRDJgth3AVXOQQoY7XXGSFE/tcmMRNGiQsjpIGcc6FtOFH25
xGiWnJsxneO6I5RIIvlFtvabP/pS1I6z4Lg1mEHhPp6d/0idLXa1vztd9YZIHckfKb9Sx5GSQyY3
NqD0XnlpmktDIkiLUcrmjxR9VvkGONxeidk9cmDzvnfy9FMEftkiw38cr+IjMqXCTBACsqbtOjNd
B/e07V/h827qwAPvvhsezWlcsHlnIn0tlbol2U9l0XTXq++o+06EflU3DdHzBYpoxHOmxye/+Djr
b+FiAn8eZe/pejUx4F2Iez4wuDs5DSb2pcKlzHNehCMkYxoOPW2c2GPHqiLTB/Yk90VUOJSwUJy3
ER3Fgc1zzYuj4aDvQ43j/yCWNHnr08QPC06pEqNHaGzKrLyMRv8pg8Uol49kLIGDYwicn9ydcyqs
U1sk1pDNDNzkOi7QSSlr7c27mcuuXyI8J4kezV0rSE5olKCZQTeR3XI89xetpmtWe7tMc+wMM7CT
6pTY9zLGjTspsLB9pSYX0FyTOjg8hhOoCiZhUhq0e11ItrN95HpeKMsi55J1ommtHQbQIB+uBigx
2vwjn642sps8bBMkCk0BQH4nIukEWsTf38vcUG4XcNtaNGkAla9QZ3qRN1T8PBSLBdUPB8REU/Hs
ETnkKcEwc/Oshr8fYVinN+aQT5B+6Zi6bk1wo2R0oT6wN8yy9umU1bYw8amjeD2dDZReXplD5MgZ
PoJQmqYTdxL2MFdsDwSvhCcPLFS+n3JoVFzBALIchJ6NTp7T6VaI/Iz+pxNOueicLWIKQsRhQte7
yBuAE/d7shGDWklsUo9T2ASBmIVwcaYXbZOiK4qR/12POa4ju7so5tBlEkWaVX/BgLT3J1oqSrda
Zl8Wd+jfij7IYw6hYaCldfK+V59Bvhexq+1DFPuU4SftjfSaFh/Cc2uBzfJuIHJBZtuFB/o+EfyI
rKW59OyQyo42vZ3f+kUrLGAIqQgaMwre7cn5F5/yqmLLg+FNAVq48fG5RRYWmtzkJ8TPI0pFL8nG
uMan+yKqwFyZ8MCHvi/o/7f8RhCrxmuVQcBdW+BZ3FRtGJsbBcsvYiPJrYyMsAjf0vsBR/8ZC2Kg
a1v2rhfAd4gJh2yfo1A85W01wEqCPZQvIxaczEqgqCUYQyH04mUsCtir2CC+e2GSzztkFBxsz48M
g1gImGBQSPckzSNPqeXNNdTvMN5KEiXt5S1hU3ByYwPRMSqVV3552+Wqu7StTVvoAUym/ijJvbRA
HP5RWLe/m4vkqac4bcvADD6bVvc88wEXEAqXifDvRtnKyIgwHfKsLYy2SoGPtHU3zyM8q1zKwg7s
QV/dQUky4sd9g4qh/UWZkcYmQRy1XDLBASbFmXLAhIRYdjob7qxjy+0CGROvxXeNh2hTaxmdYvAS
zqH/1Cr5cLCDpTKct7/oStR23y9u0+QZZYaPjUJtvYdf0z21voLKcmoiD4tYt5s9Ab0yjydo/zif
AVJkTHaHBTM248yfrZ3RpN7O0BurLJRYNr2g9Avi7jd0aC+rbWcYHAQERPKJ0vV9YWPU+4X5iMFo
ZyF0nQiFybaQJLFe72C1P/S+flSDK7wX4DqZ4QF5N3qu3Vt65JKBZ8JqElbKV7ZXeD8H+HaysNeB
uJyIe6XuxY8ZHIXfHVzA+M7YmTsK2WTowsSn8ndORMiuaQ2Bpvn8V3xuBQc8/ad/HJdsUugPguNI
Kw0TAMMC2/qFHsLtwTA5iXNfntlkMfjG3G0o8pzSYCrnOiMQJRE2zW6iDyM+kXxtq1Nz91WqAW9G
2Bv46PvD53Ji/ptDHEXQ5WYtWgKZaBdteXE08phyXoDytcUIX5L/8zmYudBnvg4smGvJRi53u07D
edK44sNGH5Ow3YNjsY1aDwV9BuuOeLU82LbbfITHlKZfmNn/xjSy4CkS71bI6blNWuzW/v5oQwKb
TdnY04uAcq8knlbBnS4rpZ2qwMfknAEclL34dOmXi8JKTZYBuy8jRSedN0IY5K6s06gSyMqzTSvJ
D5EkduS1tUN7l+WHdE/2xhz0Cx937+k5a0p9y3lhycaQqRE6ZlGZy4/O0/P9uSmYUrjVVI0oOwYj
13u8SzeikgksdiZ2RRPnp+E1kC/shSj7ev1MhSTqtofBMr5AwNGNJuLO3/w42z0UYMAgejKeDcyL
odnnSLCIxgyKP9nCaOJ5F/mwWvcn3Q0Dx8dXECYRjBpkz/RLtgKRO4e59EtaDfeeyaE+djairwxl
+iQ9LEkaSutpYaNKAgX+IByTT55nKwvU3DyPvXD7EyCvD/i9H3soPa+AxjY1gNrbCnRONb8GpnRz
LOD+Edz9tfQ5TSXgL4K+6WSXkH5G+wJZ7vZdcC1d2qcOQ+BiDRTzrw/UD6fmKp/KK5/4WJcjg7T9
EDKBlke7amR960oXRlNiIGPLux/TTlKvsuLzv7OXaomLWSl1zjIpnK6Ct3O4UO62kJGRKbScB4z2
RUdo8svfEDJ1Bjp6jTD2YyKBGV16GkQ7Sz41DZObxt3h1iocZQCc7AX8NWvDTQ7Y8AUcoS7FPSW0
mC5yQrMtIpQtG5zdbn3F2D3zbscxTaS8Gs4jmBD1olKgnihBqIzZMlxplSn4YVF4v+h8BAgEYs77
ztz5vK0mKvhAoaPh4XyAH99QhHa8F7imfnoyazEg5NQflh0HOl8oW1VXmCGuDys2w7c2PU7bwikq
//pl3OzmYncQ8PMaA9zwEOwt68NkjtWi/GNni3ZVlgi2pyOIsNNlE2xB4Vuxln8S2Ns6YD5i6GS/
fMmo9wvC/bVnV6VwSpSDz8g9UVGge27LulgN47+Vrf0P4iHxf+FPaBVqWcANGJih7HO02yI8bnWM
JXhBt26NGgwG4UOQEpf4ruVE+4ZYqXWtxj0NaxDZrDu/mj05Du3Rm/whE5moafL+r39DXSVOJVUu
R97aDPM1SYT85FXlIYfR2nW+EXQ7DEmzm9EbiUS8WQXH6xY8RxjgLffFfn97hDiGLVtkhJgTM9e3
BznxnSmMkAsvZfYknnsl8OlHrxRjDuY3DM496OT7hu3X0WGtq0EuLeg98jEinINNRCp8MaVFwnIb
fFwHoAGILbNKM1ht4xC8k9eYNTI9jgPza6cDZ/dTqqzVoD5gVfWKZpaO/P3N6Rg1QO6TAn2ZkhcV
bnsnkKgOWQzvqZSvMdeQHS+bvS4rDMlUitLRwvrd8ITd4BEvNBMHjB1/EHRMaC8aQbFXHZ0Z9GKM
UjgTRUHJqlDDN7kAx1MVbwg/40aF4ccAoCfH66KT7IFTZFV5ux5roPEbYWMrPS6s5YXP7dF8F/Wl
CRQVXmBlubi+g4tDYl1FelaC+TnQ5IDPvQX9n1Z75bnv3sZDcrcNVmt0ZsX7AeuTH6ojYzl87AFE
YngcrETlJgYwhD5+hDLxRTRRmdp5SajbMHYXaw8JJw/0qdbTAZucgtfyhdsxE1IKPG9vcpo9qgc8
76fnaWU+Y0QFS5um2Wkc8gsfg87djCL3xI86YwO8lo5gB60TpIBJJpkoK5gLgFXSPx89kDdfZO4y
9ZsG3cqpG0F7Pnii6Kcd4tNxjDxlYZ7UK8h85n3Lbv6Lptrp0vHrSieR9AEYMDwsFoDMFRrx+TfJ
PCm+Doif8vFBPOp2y5CjtDRpiE7BU4ktMHo+Gim6yMVWQYElgltcAx9niCXnCYdcY47VjfZ5J4Yg
qwykcp6PXhraiaVB5HSO8RkeTn4ICe1I2yY1vGlOJW2Bz9gnozJXokU/ThoypnReiqhw/DpJ6uou
+pGqNlyVwuzG1+RaElVA9KFrw8AIZ8lPY01OFpcanQOwAdeqzyE3nBZtuCE1qsrBVnejhb4nFzV8
Fb+EDRoj344O1nMfULP2UgAi2RqGNvzjtkOQ75/4EU1prm1sJDwSES+mASkBsNJ+WGCAAcsl9k0p
IAHZcnRUz0+TYUERyQBLzFnJdQhfxTDHDRN1yMTbt2pATCbr1poMU4qWmBCXYKWl2COTN32zlHNs
0gv4yb0XNbqnm2V+zT6Fd3LbDdJNFijDhbAkxDjuOFlI2+jAJ3Y5FwVmnDcKGHgZIPtApc0t9+ev
WyXYxueQ3DWn62ll4xj8rNIW+EIm3WflnztGjEmoRUknsUqgElB0yHOT+znU7TJEDpGVvZ3n99yj
44Cs4RpMbwMKzU7nhopefleqLCzC+lsIhP/uGAYBRrbIbAIfjylaEXBnujhxq8aTBcI0G5j27gWC
zdBe4eBDjoR2M8M0W/ATUlmsNrvCRRMdfRD865CXrXIye4cjj2sppZnKW7rzwe/oKA0pmSnzPJ3p
kg4iXQV/ey2oPUBKKsiCxKPkoyjpzhEUBUuyRazPKSAhtdYuM3vn4Jb+EywzxQxas4oyiAsbb7Fx
EtykgUDd9DHqcsRPWfNooPKexWp5VdSJLBObjZZo2AVGNCsxV76dDfVxs1ZVNtesEGwZcHR2ml8D
f0nr3Qm+ORd9y0eHx6PJQW0Kc0FZVAFm3zsd1Uxg/IaAKPQ24wNp/vwEIFfE/y2jXvTcPouOJ08Y
1+DgYqGv9K0Gzl8T41JU5j+SmUSxrGSsFib4H7jvzCsFQYDMtHutVRJK+8XG0bgtXszaLcVVE033
+NWocE3MBveG8x/tTbaQdXmQfu1PTHDejfrd10IGssyr/P1+7AkFfrsTTtRB7u13/AHe6DVSC4t0
7l96zbhigvmidMluESR3UdXj+oZV4w5FE8ILvrUXILwIIHJ2DIoCwPoh43jCb8MJFzFNtquq1s5g
pQ/iKwOfdKpDJFf0tA5ANCqj5RkFEyOY42HtFUjE0gAo7DJQMegsggA75e8+4fdzknzPp6pU4Pi8
ZPJkxnItpWroSTCRD8Gc1DxjE5vG+UwUO1N1ElyrNcgnJUnATqVsBRDGXmfacBoEfj0M/4vgwtsu
blhnaTZFuYcOMPP45dhVu1AOyMXsbZwW8qK1gFpjlgBNcqlb9lPrhajlEtdj1uM+3BWY2Ad865jE
PoFGMe5aPgitsPFgghA+Okp/NPVXtRdnd/gC3rZ4v76SGLNS2vLQrMMIC2ttOdX04vhUYEBafywk
mYVmGiwlHwEoMyPNX97DQewiQuvVPpj+Zu7smBexDHRzOKC/0uzwW4DUSUr+0BUHouwfNtehKO5n
kAPwsztU2q/Ef8kuozNG+xZPWojiO8zlWOK1oitTdeHHnFSbEeArt0hrqzziLjCXuJnJxXvhjFRs
CXkceXwE+/zjV1hM9cQCBmPdeZF/uAjvV8M90r8MrIkWr8H9l3/Rz6itfaTP6QssZVvBnGt9psWY
4y+Au10jiC2sDml+DhAFqpWlzZEHktz/CH2BBi871QqsmfGcWKo3ige1IvvWebPrn4Ryo3PxQG5+
5dtbl2WJc8Ar8TQVarg438hEQYrWnY5heh4qoRRLLBAXWx/K10wf539SlIzJd5uJE6NmCR7l1jhU
66YvEON3+M/7LXFzGYJDzR6iY6PMts4Yixax1YQHbqnuaMcf6Puj///PBfRCxDwfDCFtniFc7gdj
qncArntX2KbypuQYZ4ADSLK+r+o4jPig2CUwWSAHmwNWCXGQcppxUGVuuj5Ed43yHsCTod/2jMD2
2YatMxtfuRffCjr5YjCR1WU9JKCLwDSUt+CsZPjOq3NltRb6diWBim/zUDp87PoRqZsl7+NZ5gYG
RE3RZJdv/atxgCM9H7R4SGHMASA2RDJFM2YPIh/Bu6c+M3QUWrd70cLTUXhi1AXzRh8B8/Vw7R1Y
qCaKJExc6j1nMQFSNqsGCCwa1lUdO0g2SbT5+LnByIMwZdL53mQG+MkaxxNid2b5YGFronEBbBOT
gVsrl3QMwNWMpw4hunIF4pCH6xcJA+5HUs49grq/WuPsxM9CRX5oShzxlafX26eBXodOETvQeO/t
meyP2vJNxoyeCX0wi/10OybIwGDQdqQNBdpo1dG0wYuSG4ePYLiBNMfqRPV0bMQvR1G9PbSilthb
FwR6hBddTCGlXmG4Wp7fREV0uhRM1XGKrquCSMIEQfI5a38XmgZlXZ+cg9XuuTVyCGQn9Z5R95fT
AolUvsf0LFRglqXKyMJRq393QRWkT0E+hg0fKHSFxgX9xt7Z29U5vB/oyo/XeaBsCJJHC3DRP0fe
2pyZwrEpPQAclfr2JEnwHeCLzRix1I2cJjcHTEfhNA60rAXCvGaJGfWlTciNPDDs8iLWXVN1Q3kQ
t9CNlkxEqeZLAi1Mte0umDYKJPTfYeJShNUQYotK80NuU5a2dJ3zSNpwjGlaeY7okL/3n8wQAKZS
6iHmBWMPrvMANLqj9+Nz4MtoYd9gwRd0+Rmq1I2EzVo/gr+F8ZpJSBt0P8UwCLGWEPLVFWNm8jBj
nBYDGXSpuUTq43E8KBAm3Eb48kFUq87LGdwKKstEZYDod3Xlv+7ZmGLtmx+n5vusyygSPz/RTJta
5skVcucqYcjd2ndpzgyJQGn9Jra8gwMimsuewZQIP9rnavXMJy5t8nYUn0DF8cconIVijK8Nkw6o
emMjqveg/4xhOBhprTsRxc2kBflGcdLbCu6PIDjpHozVLQOrjlFX51fF2WFsN2qbbXPH5lIAYVYD
WF02MhQp3QSlpDAjaDi07eSvrhqOkm8VbsXB5Hn9ulf4iLJ0P2YpiKipFFnvCXQWIjh/bcqEujY0
o7/s30SCrSQleFtrAAd4Fe4cSl4H0fJvxESJYiVyjDz+qJ8WQMleI5nzZeU9B88EMFv2eSCnYN4s
3t3l11v7V7XxZm+KiwX8AJfmQjKogcGdBSgsxTjoaOkRmuXAYxrDjsscCjSBghG1txFzlzn5fiCr
pmBSKQWCc5LtF2BY/j1dYMOUCERpfTfhyxXdO67AhKS71rUvXWUcCIY8MdB8CHyn+HYm2Xo62ec0
8EJ1yE4C6mybwq2KnW2xDOOQ5IHjze2NJZHhDPnErwCprOun5VnEPzYit7uXvcEvhRpOPS3+aVOJ
Oi0Ho4s2DwKKct0L/YAwRqT4CMClOHnluq7CkFFerh5iwmmfRs2a8XuXcuScsbnH+NSn2Jk6037R
kTFf5+FNl6Gld7XFyWa9iRQwi0MaU/0PN+c97bu1nGLLCZJk0xE9klsi3sp32GFjMoCl2SkUIGGS
m25d+cCLIeccKhnUqyoQHZ7OEIVGfdDg/lasvkW2ZGc3ZD0MGKGQEQT828+rXJp6lEVmyu2AToII
RpmoJ+5YEjIOaDWRh/soR29oObF/ve/WcoA4Zcd6uCrncGC5k6TcmK/rKZ+IXRjW/UJ+O6tarWsv
g/IEXiiL70aqQrvcWwLyqX1Ip3nLg+9Gq4Lu+1RvV6QehKeVEi5vzGsVaxtKNNc/ZvMoBRFBJ1C8
BNJ1U1248Kz6Y6A+U29YexRJ2nqTrLT9wI/vm/aksP34Hz3AIWNXYz36mzbttYhjBtgszl11OAGb
TFmcnDAEkouLrDY7Orx1CyWqjk9ICjAiJcsO9cUkqUE2P/hqf0ApObqCj9J0CsJ3FBFpr8XJiJCP
uf3OeglONmto7kBjvOl/nyXp/UDeKZtyJmkRQbxn3v4BI94T+P2bBwBIILLSwYycj2YQNJ8aIZ1g
w2T1Gacdq8cH7pOgSmc0kjtqLyNy/YPFUVmETmCh2Lr3c4HEiInllmouHt7Mz76hdBN9UxMNez/F
YN9aGhZigdEymW3xNYVmeivMGfX0YtLUZXD9TFWKMA8dbI6KHfQdcT2L7ta5Vrv/eco5nigeFGuU
6Kq4KoEmTvwHepa1mgeMZLMKjEZvQhodGWhxz0Mni9edi2DQyGZAWb9VITrbBdj7mCXZ+GJ9LqNN
/haqi0nMajdYj8JlqSMs4ZB2VRDOaLr86JNegw1EHdoHjLXeY8E37s2BS+6sYS13p72SUJ5xN3XH
tzBIC+Fkk9ciQZAPlfsnEBH6d8EmkF9ylYe27+MrxuvJtlB7hHSXDukpa71V5mpn9cl4it4SsHqK
07VWPSRYSnuMIl4EsGzrWpQAg1y/I3O7/EUrZ5yG9CmyhwA9fyBRGTocttnw+76IKqmARu6HaOcU
yUU3DFQRJFFKjN8t4kN4HLdLAI20AS/+Q9+9xiCKXcwQCp/TyjHMl+Ez3hK0rT941djZI6H7YJk4
ctyfZA+HkD50xuI2afeKOyFzn3546bUYS4SET+jZHUlM5eHwf55/4kjBLv2VwhNQ3R/LXOb1xSZh
HMwuJH8IywwW2IwDW2+MnpGWzcg706JYziKRSf4+bkwqubTgnssjuoNIgPtrNzRi+jtfiMpCP0ob
CT433r6u7P6WEQdV/+6DRrHV+5rp05OYIZqYVsrz5dKj34xM1yt4FiUBynPZmKTa4yODsqh+0QIw
Lze1jSCoAByHu7WY5KfBmnc8bD1NaOA9v8aBxfEd51+BgqTaY/PELwZmOl9vcPlX5/YBoRTe6hL6
4XXYe25lz6ZJWUpwFb46T/fcpybbrK3X7VSLFqcjvRuoAfmVQbtOWq/Vx5yJLwVLUxpViPb0n58P
2wH/riFOxzinh3FqiyutG3yft/C8PVU7tPFfHa4cLBwmYU3Y3kcBZeqZbLhmEAmYB1L3CQsEKCJo
aPMRXKeavaEthAX4kPLUbcxafYHA7lrR/NywmD4CeaHySnnQ9MJacIf8zWMAg4zi0fG5g3wnn/Ba
wXtFjSSVcxgToXv5MvRgCwmyBgnJNlpE3zZiUeiGFabHxGcwA3e7BTEwiLy3leODxPuXR4BpjIQR
x2LfEtPkiueOh0KtBf2PVREMXEvJSBNrzoz8Y2h0bG/h0fpFWvJlK3fMy1mCed/EHicrqT+aR/+v
EhycjHiFU3Ytd+bBgjU8bpU/xaLGuE+eKhLcqgMM1fLB436mWEHX/EQzSG9IW81ZKNm/2JEwbMYG
dd8Mz8GjzHbUn7kIpSE8LT12nXHVBgvvbt079GrGR+zt7ZggEzKB2gej9AYW1qwCrjhWC6u3BFVK
PTFU/UieEafzNltL2BzvNL0hecPnQS7Q9LFUrCnWUG/aClA79Hzp92tb0Z2yZL85DvzHVX4Z1pIS
t1+5jLXN5eo47dXCsmVqYrgRGDGa4V12dtLJWcpYPRCqqI9PpGZbPn6LaB1djowCy4n23gFAiPDT
9/IDQREAbZseQJ95GTNSLrjEBlkOZuewo8CdyBb6dPl3DCukW7+wyjfCByRwk01tCsE/luggHujB
nDphq78zLKBa+L8mkgYDgxvWq80nCq054/GWmy708601OjWGpICnJ7a0vkybQJseT20i0btg87Xy
8GC3wxgzvQxhnaccwgcjcu+frhMfm81UNcWGNs6gMEH5TO/657vEhJZex8KxyQySqaewarAurdEL
SyTspvf8E+WoTV0xNpiSg4CrULGG4PFNTSY/WYmvwr2r6+BvDb648SUnHHy1lZ0zqg6XVa7DKlZv
9t1i29LSGP8ZXiilqnLAJazc8QgRwkfoPOUi9GZ0bnERFL9kBc7MDZ6LRIL/5LCC6O4O8bCcHvAp
wSyK2YmyT40wp6sPrmtHK1233SLywCM2k3kQVtk5n56cxQ5pLI6/MjqGIk0KVKXKknY4ohbLXmlE
YuDRn+MJ4Fs/JUtkDnrGKkRkC3mSz06lR0DQp22uFrjSRqF9yrJSPYU8/Cs5/U3pnDH7IeJ6t+pB
vpAFthlbbYlua+uCqczADJlblRZo21HYm51DfS4m3Q1IyjCe4blLTV0J46FR/27p3Nx8W7/zFNYj
OTfZ8gI813aNJOPh28B5ZirX+YCf4c2PgkBtmUJPw521HrQbM2m+pKMw0TwNXsMRkvKFXGbI2gCN
7nMDfKApw6sKGo8aETKV57LAQ3u+A3wfksau3KszbeB8Ki8EGtC2d1Xs8ddtcMoDXJ6WsJRfXxRQ
zneJyZ52LtTWH/GRxUuSrRFq/3PRUSt9v3+zOMi7YvoAxl8u5/2OZb1oelXSFs+Dm3dgfYbH7Kyo
Nhp2otrH8+tQfJj+S98ZAu//cK4tecjy2R2Xp4wT/hzJNKNDIUmw+yEO4UCmokMIzyF0zRnBAAAe
6uDgcnDpFidgInFmRUx2KPWU+07WJkXJAQKnlN/DnZaNrJr8CPaD+9L2Da/hdGV4LIwJVnpTmZPT
3AE1t6J/YTDs0RaEXk/pYMz0rnY45DRkc1iDF+uo2GBz5VRMYJhLnE6iqFf9AwnVqNNgwb69bcpC
Var8rYHsrASZwE/Ph1OGNqMfZhSatA6PfSU//VKNydFMEVw61WkYCQwqUmQo/il8TmAN069WETx/
DSskmmSaoIX/lO6nfNmYm12kijH6EeErLelFPLdhG5hwLQd/TCQBqYr73o/kQpsJoOYTQ8lEzVqG
MgN8pPj3MOyjD94XJalOtE0L1lpBo0s2ATG8yBylQ0XjpclI/itrTbpNpXsnHqCre1TMC88L0B/+
YMGwDW/GQmilQEqjeK2oPRxkJTx6qwcqn5NJXgDQdtYAwN5P8O+2fqx7gr+7bURuxAt3ttiFvWmK
ZEeguG9GUs/9EGzljLp7SxYRgAcTGJHecJXBMt0ov2AP43T4tAdFF8qXABZcXTxKl/qqzzm/oFbs
E6xOqu9w1kiCZaNDf5FkfNcIHFeoFAEYWjua42ZsedX6R4HTH2uXbSld6xg/PdMctBdwxjTRYK7v
IvJI36nYR6pWlkOs+Fe95z6jHob4lEEK6OAeiX9PkoAVESXlr7CdqTpQ+H4evu9XpfJOp12FWbIU
y7tgzBFKMWrHqcBDvsdK/Xb/vKyjMAdXlQkCGbZ6kH/rIHb3rmjPBLSA3LFBuYxBmoR1Njpvr5mM
lbITZcuuvZZ4EyLIuVZHo8kbEdmDQ9/CfMk45UVjuUO5kNFJNDjvzObg+oggbmnoDnW83+wi0eZ2
tiGX6zpmHEEiltlj/1ppz+7Cqk/MvLXUBa7d2kjMs66zo7wI6Flx1NMa8V2Zshr3cMjhDYbDjWf+
06dKlsTp40ztQ/zVGNxQihA+viriSVCO8O5nDNndEwXa2nmxrse7t3149maEROMlCG104/2cVPdY
WugUwU3Zporc+UDZrPhQ86cyu2G3a83Ocl/IdMJM2OHuoVd062DKMNIPTuil3ghmcei7zjGz1xXs
SO1R7AGWYQCK2xK5njosNgpSshGyl1Xs8ImZJ/QjauK14cVoZhs0EX/HEx+MQvH4i+wfrM7ZWzFz
v/93GpP3+CLfHvwL4a+a5D9TexLHn0CvluBz9S1dD55WWsJNfDqn/8FtlCZYJYKhKpHbQfu0Td64
dw8Hilh+LUWH5FC20B18gTwfYEU2spzT4Dvzxi5eMi1imzI6GihMQyanbGZEZqCdDPOe1YT/hSow
4NHMvInMqcDaD1A03UNS9Zk4y/a5gme2ukJyjF5TgB8nKPJlap/NWrANJarsZnlqsSkgSi7Mjie2
hny7Nw55j4d3I4R4vgpdlmADHeqYuCQ8ZK1pmCbVXbIHsflaNo3xT8yDaUvthaPmrY20AI0e+HC2
A3rlTt+CjtX0JcsxYwLdXCvmO4TfHb/F/UIgWivDQ3w7F96Rp+pCtuRdVC7AgLVJPvYRDJlrbvdc
PMyV4C3lqg8EQOYYHnQSeSfyvwY5RW3J5QE4HVXTPPga5rkaaNWvSBB4LF3z6qWCYMUjxHGldKcr
4i0FAkLgaIdvpmJ19h3qP2DWqis1XkrlVwJ8zHX1JcqFVbkjvoJ0+W7r7Hf5I9Mzi0G8/xSHWTly
aIIoEIqt+soIxDE/hne/wTP/t5hiGXL6oMIygq+PNTCtWwbRpvui5nvuy4tON1vINBgphugnOjPl
WvIFd1TWQVdqRjbI8rRU8yODAdoISHWAq/zSSzoiejymu0ygSR/B4RgUv+Y1HINK2IAtefJYdM/B
6JQNyyf9Z+5jofCIVzjEq0gae8GyqNErAqjeeuDUz4e+n0VaOBK6BiJdDcKU5+FlmB5zOShPA534
UyV9e8GpgOnK1KjqiIX5wRkHhe5AQT2AbwkSPyjPYi2koqdNRsH+UqIb01gCr/h5xxR3/YgmsTHn
K3sG/E+pyWv9XdU3Z01nD1qQAcA6lQH1ga7dKBzzQ0Jge1D7fjgjSJHSpDVo2XDVeTJ/MGFl3e2y
qO3T74nD4E+dsyZ7pe+16Lm5PGa5Mny3DbtJ3/7sRYVotUP73+ONdvNMhRPUD65ZyW8huVpHl5+Q
5kMFVhkYdeJlCuQetTlCGiLd/EHU0t2KYhkoQxXhW/RZax1qEL+OcDFpVXnKYGkZN+m069bXDKyn
nCDggazaHPOjpA66WV69uUazUKVlhSHOhD8cDCOy4G/tHFIy/+r5yjsB/Qt1pwRCQ8P8reulYfOb
X1W2PMPUmbU7no4OgUo3h946mGJ3ndPzqDHDL5c/Ywigzdv2YKU1SZ99jeLpAtfI6a6bfZ7ZPTlm
dd39lUnPaSW+U5NlVy9SxkMc5XVHYZcBXVihH7pr8H8vXXJVKSbstrr3q7lkmNXgq9OSyS2L70Dg
K+B9O4UprAS9Lzfi6CemsEUAm6TTM0Rajr7n/BfqmSeLF5CqNgzFY8WlkOqUBtLgx0twO6ctFA/J
OqeGR8obvapPkLdZcvlW9EvZSUz6HxhLpaRcresw6CSnOHXP+eVjVIAe1q5G22ts8XjOUhtAsGIg
kLPH5bPSD8FD14fPjBki5Dbsku/ev05Hyk34b7u53vOyt/ivwIJ/CxSSeu5IRIlUPt+qv1ZNiRu4
HtXCueGDdaIbPcXm6ZwXVnkx3dHcffOp5u82Z6e+5Iwtv+baVjsjYqjyyMeFl1Axibk30CrlQJ6d
AuBPHT/ZFIqPKQ2v44Q3zL5wjtcxVwV4i9CtkWdz3jZ5eQrRvN/hpTz7Ihfbska/NksrvWJWfyWG
40Fd8weRHKYjcEOG4XuRCAcwbS+knJoLxJsansFv1WumVrXq3JUDDoKzkKTCvW44chCsutL574Ux
1q/RvSdJQw552yRzQUCjoZm+lTNJtjemRc3vZGmASDNdbLRvYJka90F7q6v3Vo4vtku3HBK70pTF
1obS7nU99jqpEFtmK5ytlBVMz1SsVmLnZHIrJvDS967nf9ngM6wrjaIKSvWIflWpYZEGQ9Nd7GPr
797NtSXkI1cxilALb0HYcQ/89wlYVnmPTd8Z54yaHIKFV8MvYeOU2sofxoqrYchDoXtI9K79Jtru
s0F0oCe5pQ4CBMZm3eioF9xJjXzFaJlfp6SUE0gBIaAxMsqCRHQ8ZBdubTlI3RR7nn83pTj0mkXC
JXodwKkG4cbgN8RQOLueDbD7uhCQnK61RT6w5Z5XAe1MY2zfiO64a7iroOson95Gl0Z1j/Tqt6c5
xYrrFQnEjQsuTUstpjClHEsX3WLR06ouarQHxUOBoiOjOeqK1lKp3+93u0F3e/rY6EVkFRNwfdlW
IfZL8qTMAIU6FfgeBhsIxlGwOJwADeBYLvSuXCt3bl7z4RWAv388lFMTyh/dF6xCFlUMhEPwRtgi
qD/e4lefw8w8aFtePcrNsCbH6Qqpr3vmhldF58S2bM6ywF8PbI7SvhsadVs0ocIQ9dIL5V31+Zbw
azRMni0jtLngjPsrBtJG++643cqrDWP3IZuJZENJGl7/Qmw6pe3lyJrtZ/J3QWh/QU81F9Ytu9Ub
p2AhK68FtR9Y9Dzn+rwRtbNFdzFFWIR0+89z9zhNgO5r67eawVCiuO61b+5wEki07zxbs3x52V+z
dm7O2F8XcgnjjI9tcfMLU7eeb6pDn63h11znrwdGA8MTmtRa2z5JUPRe2+44DvqPWec8Kk6ov5K7
tha6Wb5TGn764uueu6xMvrVBbrBk9e0PCHs3bvUSaLNsa6Rganqh6cnYDwFpvvmNASNTllWv05a+
QrVkfJt07y1OvCJoWW4dd+Ja9ziLzREYbok177rKPOPBJLTDyRkh874Ny7c0ih8d+XGIuE/XqZJZ
PdS+IdfJlVROo2WoPf6Z3UdUJpFYQWXPnL3FPc1+UDlqZcp1YbdKeee/I58qs+WYCqyBOsITeAdr
hYqLmve/0UN3wnPT/e5j4LZPXTfU38HaaQmQhHGrE3FQhRHqU8/DZehawdu4MdwSuvkoAXUuSiF0
3izyENevz4KxlS4iR/LOTAPXoJ+c0Y8hnVdz4rSY28rZjmZGcVlIEnKgRATY4OVBbE1nPlvPmlGu
2vLAQJ8gSzGLelAD67w9uSMnm51GDfd5nIZo+cgpAp/X7Gts48XfKhyba072FCz2R/WhB1rX37kW
+o2Cs4a+xw/JXqh19he3poT++4/V6vflDzbSR+eNeZd+PRAwbtJLwOEeZyy8sq9q+TLGOQbOZxn3
iM3NP9WROJOPXEiQpIn5s5AQQDGfGm9S4X4YF2gN50OxZ3NOf1GRXK2j7Ox05uJ18kWqgoMHnAqM
d7Z3aBumWVJ2wXM5QsDXBenI7ZSNpAThjxQjySVz5ynD/vCEx33tPDLHXDIyNkc99JRhLxFaBMdU
442neEHgb8MHZDNXz/n9Vu8E1xiri78G2786cZjSrQ6p8HPSyp1HOXwp4X26tSE6uhu+aCFLpiV/
I0kWKs29azOlFzIfv+yO4IPpLBYxiPGxBVhmaoJBWuAA97Y8/I+TXFXWSP9Rps/jBxOT3mycjG7l
ne7l8OqEeUREPrC6G/YUdlAHKIXIDEZ6/Pu9DCA0XPGspemZQqrqFz9Ri60sCV8q2W3XVqkV8n2z
tRnPny5+AMmkuPRzJCcsAdRvFwAVIXAJMGOnWiQntEm93qfmD11R5696+ap1WK8YzHYFgyXcxRFq
Q4WnMWPXAE5xMwEXO9Yzz6Q6wnqiScZBynXxs8YHpE3Z+qR/OrA59RmbItoZBLSjaOzUXlstiK4k
BzNGegeV6Is/M5VzS/3UM0yha/YMoQOIawD38J1/q1Q2oHjD4r4pLyM+QqC1IOeax9GO0sfV0Vq/
3w/AZRZcXEhtG832otzvHhise0kObbzq+8JW7qmdNLI/6EZpm/QUUAJ3dA1MzKLtwyC/Cu+o/Njx
lK6NiobNla2+IapODNxF9Z+Cpl3HY/qQKuVonvdSQ6cXp+KzSJTAUET0lb37OSzrLxpQnK/NQbIP
bNLFtEKCo4SUQ8NXYi/ZXN/mGlz7RyNjRkk84XYC7VJVGHVxND+9CxWPZnSzPcgDrUxbqZX8NF1N
VhKkihektCW4VH5il0OJQfDtJPHcZNgwyUl+3wCN/X9DCRrSQ85w2K38z8vDEaay4FZFRjFuAfUI
YPMUEGGxmCfUDgCKQRHrP9OjUN71DAnPHevJiF9gozlZneaeWs2wBHVE2iCT23H53/cx3q6z2mhr
/t8PiY1vEq14UfjUXj0N9xs26tTBn1m3QowHs9JipzDgxMkYu19yZUuTN74xtfj2u+gw5WqP3yqV
8s6TIcTLcxlmZXkFlS04I7UBQzwQql5NciishnoGYLS068ZS4fEXAYGvwum8cJXeQgk2U1K2HEyZ
PGckS3I85vIxq3JQHLGTnTqHaTFWX1cMLLYWUVXGXhlhuDjf3Pc+TaQx5VTeWDwwF7p9m/FJYdf5
S0uF2/SLWNdrOGHRwi8nCaVPxjfIZTX57LnO+zWuXrGxIA4uKTL/fuWMoDAVBUNkiSigM78GWWAK
MAwO0sQtvIlbA7ZNCDins4Z03mhUslWPnRcywg3xs1G1EkDnQFhJUdl8Ecj2cAZsy+HNZY8xBg+z
cwtwH4T5ZFoW17vaPLTOVQOMqaB842Lm1gbs1UrLZU3hrlYCmBMHMhT2LDCismatncauhlE0m0Mx
wQsmfMi/UX107tBvbhO6XoNsLO/OdVwiTTgCrAa5fsVOOeSEoxcz/WUJCgVKkDrTplWn1YfaG0xi
rDGWgMu357vOCSVUTBIk+5mqbVLxu3I1jBsNeyqdDKV6bRIlzmF2ZA9RXN4kpRYC7Txm+NhASkef
0WpVCxL+YT5Cp6LAMwuRC3RwSWh09WU5jZ3fKkp2gG8kQzaPDBD3y94RQ7+MvoeKRnEATDeddVi5
Smr1aDuKgBtzaP9fJrimduGd6lCKCkYJ+0AvuhVrtmwgMd3UyJ+rt+CTqwimWZqIs5tH0Nzmdjul
vUYgaj7UuNJSKooFA3AYUD6T2Vdw7h27p9EF3H/0PDGHrfRrshHGlJ+gJ/oIx6c37PPaeQu5j4QN
lFlcDCHzBLecVxM9JJ2tJ9jJylxvbJKyFXHI6k4Fx0tivNyPZVF3przul9TsSvuYffH11y2OyeUi
2Yoo7QCXkcFSsapt3j8iiDznNj4gSOHsHD0YwP5SNSDuaJy834UtvPAJW4BXvrFMQ/eX449es7Bk
MAv2x0m1/kwMa3m70lVQ05iem7WkINoPb0DTuN08XavVG8oFgTe954XyLREsIhdFSuLiD0R7UYFM
5Y06vup/WVo0NoK8Uk/qJ7W9BGMp+0FQ5X34VGRQLGV/vqPD6R2ksfcGwOVlNFC04UPKkiD7Nbqd
usR/UICXQ3KlS/g4WpH7CVcV20JpuSBjsUlTno14x+m1P9aFcn7VCwEu40fd91I7IUt5mHSdOldL
yswuhm2EMaMwlgFfEcaooXDkn6i4K567OTsLkmn1d65csxpYsKKqATBXsa0h8UuPT5ipmQOtd2I2
IY3Ey8n4HrFxXjKOq1al7wvPP8M9qZWvDSEH71IxMFJXaPLh5QWL239A5wcFIWbL1CIVC7Cb0tHS
biFwszMjOq1DDaTsqbTtDo7ezbxdSO+gr6x5jbpy0qF2zsxLysAk4QAzY9DW9PqDLQiTnikChzTV
vyUQ3u3M0r/SRsJfM5Vs4uOmBJY9i3G2PPYqmdAPmNYa3WciXSARVlSbwyreKXgeyQoky08Iy0xz
Wm0jAZhCuyfL/oU4WL88rPXKsQWe4m2227wQptDStAE2tQzFUsioeeQAKqsDHGNd6ix5hi1ZDly7
Gju3ITK6oWUkFhAjEygWVv6FwyvDFSp67EOn8Mh0Fs62Xr5tp0BFK8upzSStV7Fxv28DA/su/VUS
udOkBtvvM6WHUfdXAhP22RGQ28XbV/luRR8l5vdWwg2MtPbSlZXPHsVQo4/ecThHebb18Ea9M3vB
kJCf04OSpg6wBh8hlzTyUPI/8goe+KYjsMB0tTH7fw6MF2DkbjRsXOR4m7hWEKbrJ7iPQ+MDUQzs
hGXVBQBQnvE7r05SW6WEoMQK84IX00YG9EsVWz0pM+sVBF5QswuIjghAr5JKwdchGd1VnX/Zyhsk
4I2HAqwEu//wJzoYyKVtR7mbQwGMB3EvQsStHusavqCO5m37tYmzsVcvScbMGZNtCsWoj9OZ3Leu
CSlKNYBQWsEijxhb+Yo8gZCZkWgT3BqNFmQTO+hR1F8WP0q4omcBKo8JkiUCShuNK5sM8yn4kjwi
r7ReZ0lURQL4L4VeNFOoQOYFeRpNcfh0hZ3pbcpJ7IYJ7Tfr9fvUzdqGzEThLWsinEz8eTX1Qqj6
t/fszoSdC7mdti0MuF3xEwwQENoiDBgqFeeNXWO+MYBekWwPOhsQuVzXYG6/tAjSrqmO6CzOYwIo
3lJOuiVIpi5mRm+OioJrHa1In3fevUjBd1ilaC/8SFxZkHtxFWxb8JgtPKFM6SCYIvZfz7g+pvP0
zEQerBlkL7miWKCyjRq9OZSeDYy/8zMB3hWo+nVXc3UeFDMpJRZlNJlrAEqbwVl5HfFXBGY1iNzy
fn7xRJ0Ye3WX2BsPMj0JSGJhgqzH/sH270C89H5enl8PhEniBomETx//nVTri/pULO81C1TYSbqN
sgw9g1u3qPBjAgh1keeHQXtBco5CqgTILaDfUEUWy/DhiFuoeqrg1T3j7yMH7+CwOPuTOW0mHKb+
We3OQQ5/K9WTsYiF5pJVOX9nb8UVPVz0oy2gg68wtDOd8qC+lqudr0ZcYkr25ADdQs2X0qurqh4e
TVM9Se8aeoyVmnJ3A4vm+XWlKn7yASI9RCX0bYE0Txa+J5LM9Ddll3rbkHs+LDxjEh0QNfd+Brkg
tpfcs1jvF2fH1I0T3Q+xJnm2ib8wUMfY8WIcPynzdBBSOrBX7LxH78sgK3/eGPJ9a5UgLw0zFEAN
nbEydbGEwSqWSn6qS12vKyVwON17Z2I/KWs3Z3t7oqVjL29U6l8X9N8ED4DkDbCQXhqHulWTVrYW
tMw/9bCN15ppcrd4EAVT07LPs1TZMkFh5itds99hTjZ8nrJmFprMZoT5dafmOBLoCD8QX2B2OhS6
iw7H+2C/2T2NqKC1OYQKNcqkjAqXcdyB7DgebvHXo553hHev6ggRYVaOmoP35SjUvjEYnISSIcQi
FGROcgRUhSDCtFx3Iz+4AI9ZSAtYT6Rd080zvQms9Wn8x5WEmpRkmrCGx1rZGfq44hFIw8v7iXTY
O5gskJ9LvV0rgXgFQgdEpQi+kkRZFcqgC8qTU4cVoYi9122+BN1tBpUovcu07I1zGCEbrbbw1lHY
8yA9tNDXH9xdBea++RuWxkxERRWdzxXyyY56+jHLBRF8tFaLXMMJRzNJwYwzV7bnUnf0cY/CNtC+
vwrhNTGvF+U/7Pe0au12L8YLcSnrqSQ288BydlutAwoadymsE/nvmJpcPWZ9sn8G2HfaYY4mi4aC
k1KIPTsCKmqyN7XLybRElZnVplXcNLoEmC/A/FJOsS99Ixp0Mqnvk+8cbenz8XXkrlmjk0oSW+RD
Y9vDp7PZCrOgQmWCssP3bkUU/l6owqOxY8jTrE7aWcZ6ZBU8QzwDaQSgOjKJAsOPkS5Doiq669Ke
OYHUtjrg6aFxnKqhNUh34vRsXL3NyO4MO7uM86xClsPLj+ktYUTcO6jOxp/1Ta3KfH8apK7AzGjX
CGHZby4qA9nyPxA3VrnySOL3q7PJFITlojjSgA4lq+icdTN1wtlEh+ATHTfQ3Egr72JgmgZp3n5C
X85qTqj1R17aySCQfk9VLJHzbKL9PrMjdvNZEbuHE4SRmbsar7ME/Hvl1z1CAzE+Ce6Sdbv2eFid
hTrqEGXd0kid6hw3MgX7S1HIIW+vzBkPLA7dtZpWZNI2wa67CeskXLRqJKo6c/xCo4i54j655oFl
SQDR7e5/SXthTOc/VenPVSGV3EtpMG/Z0O+FXwfboPpxGE/OVO1o9PlZWwNGM0Io+xd11Agt0T5x
uHlYkhoSSY+PLmP0fguvqbswcP1b+94UEQ1ZPRi9HE4ZXI61K7coC8m6+Kfqsv/BD8HwxIdlfKss
ylpad+tTM2hIZtfOZQ1cebU0CeKIuQ9s+VAxCiJ5Mwx1zC+oX3bXi5syl2Y9vlRUMf7oEPthaoUr
vPu4yXunQvzIZEiln97W/zv3IdxzxrrTJWgn8AdOGN9qeSDgsIf/doB1ma6UHHJmPZOSPgyar4yU
9l8tSYUmvc3O0dXBcjfvImv3E3b/KyDSLeFywpNpOMMHZOimxjt8Yd/00S7jXH/OH0U0JRgo7OdC
D5bEY4IyoxquOo7yJH9DNxEcwYQOo/is7OGAF8CUYp3SU2UNxnZ7yM3d8PLsY4Si8KnJKvxu/viI
ZtEGd17vWw8HQYeRHDjKUo1YTpvdI+fwbFHnX0BXCoqFFrVYvTeE2T0UAR1jW0jy4FtWl1Phmxng
MhXvSn0c+8GY8cKEKJxVLJq3lRQF/bdi4Hobj2rOxiXnKsBluCVMqInDtJi3ap1IIdaYmDTUpWll
Hv+60SnW+puljCNVVzt6iqL5+35Xan54iFfIuplNDIYo5IFA8QynpnQlbaAjQEW8JKscf5VuA0SR
FdDILDzxabM9h3L6lFbGJL6rzhr2lztPV1WwMolMQ/vn0FjsVLYp6svg5QT+y4zYg/0b5EI7rXnH
o8XCPWWQln7KF3Rlo8XHcLj2zdJFbLHM5P33xUEOM0wazsO3NLhiswUKNCPDAeX8rr8DI8DPSBmF
eYxs1SSiRLFVF0/VB0OCgH+0r73GFpcHCOWrTIT/dQ/7FaKzGEVNBsEqf/2QpsW2ybd1T16cQLvC
GYQdTZYfJ1IBWLAphLB730dzFn1RGJhVwtu4tKSPjB7CEIvqKQGSPrXj9NFlg3NNnEfz2KTMv8EP
8Rrln6HzqIaNnnRHouGkixU7FZaIWrWUlxxGQ7QDnVNoGVDUvFN8J2/Q3K8oi6/mOb+tZzF62UrU
Li04pLakO+XZ6g+g4DntmKy3BJujDB/DLmAPeL6+WNAiDzegUqsfN3VmRW2uWYQLF+vLjxb2MfQp
Ti6M3g9qnZl2VbsCjb2LKCWnwe9d9MSWLYXzG4KeHyjCAlqqoLRKiZgghDsbVS87JVrga3auXvK4
np6+7sQhwB6feOubNXozFb3OTiSDBF5aCVroL+Hl+ZI17EKI1Jwwv4xcAPayK/odAaksdtYS4e0x
AMraYhtpe9MNvcn6rt3gWAJQ3xp3vWACogJ4S5XRo1T80O1UJ+Qb5qlr10lrfaj+1r6R9qPQxLDC
gclEX3FMNMvQwerLAEuQOJ/Afjpw2LTZiWq5WIH7tvtxunjEdu1cXbEfq7QfGvAmQ6HFz2N8f19U
aLRXd9l0QXBF9AOr13FR8oN4EukPlZ+KqZ+Jyp7ViM4fJYSuxg3L85qwPl66RRNBaqQKV1agmwxx
8hoZtm3bclswblE9VdwZdS2Z6YIzr0S3Ef3HDBOWVJIAQIKiFXR6G+/170g3TJciHV5ua7gTOrsY
jLHENQgFlMvPH2LUgIRv1TiszjLy59x8TgSz3mIYo7A2RwLrMRlgQbRYu0l957s7Uo10hCn1B7vo
SOunh2I5G1D2zth0kzZJclAwoas6DM64425J7Vvbk/Tz3NZFjakfprvZ68kDnbF6VN/SRol4ZkHX
13Sx8UjQV2aofXc6gjBhLRNqnEYl8isZZhZYd7hOAuR4j6dSpZZ3l+4Efbns85agrpXirkyHjXKG
vFtYKYg3XGEmsc8DzRm5NXxNouEwxDM5iFuWMxa/xlX/0/e2q24ZaaC/1cSx12+FxTbSWxk8nlr+
Y4iQHj3qB5m1Wf/fDKgggcEWsgwpr41B2xzFbHZ3F5xYVNOARKyaCFXl9GluTE80sstaPqoI8OSe
pOwuqhJg93025s9fQYWTl1V9j8HI75fSTvuy9RYQCPXmsL5djZw/aEZyUBnDYmleg4AenkM727Ok
8/NIHgG3ydX/24hA71z2J5rZAUGTBMtwb/N6fKzHNBQVbz09PFRHO4FeH+MigZWywkbD+dsV4tIT
N6+lrNl2wCKtVt/7ClOael7vAVvaOIVKu3tt7WeeZbFmKruZ3JaKOpaXrrmLZAqu5BEwqlv1yjnO
nKzPk5Mlb96fWlk9OROSrmJ+qrQ2rYTYZwXfDtkLPtsDrivWX8hbYt1nbODyjbmt4VUI4bnFdonV
DWuSzDW/pZnOrCwf+yVqBkGupt738qIBrKRvJMF1W+QJwd8AWfrfQ4l2U56m30hPRNQuUd6EpuyO
K5xwsxsmZ2jXgPF7GrwpkoVv+zmKBrq5RUbjmHxTjD1cKT1/YfC6ZMsQUaS+wOv/RtSqIi0pA/Bs
R/MVOgYiMF/b+atfVcMBQL6bKSbOh2Ep8twrAJ3ACcWhzUoR5URVTioiu/W2e3eQw/AgpijfKxbL
xT070jnkem28vHCjCvStOqYvReGlgT9IVQ+L2gTG3nObNyPq02vyUkf7FtnIL1+A77ThdWCx2BvT
weIHZnnTr0ZuCo3/Y2oHFNDygHopluioA9TlYutJ3nzl4NtqrICSQdtMii5PQO8OcDppOBJG9vGt
MOJbAyQUglmPqTF2FW3oyEQOKYQGZ6uUTOZq2uFqfv27J7kVOQDGwJjINhnBuXJBuOVhW7zhhiWc
1MZVsbDAWFgPIW9oz5bw/SSwN5DXHm7Q8kfmCWOmJX1M9xHLZUdPOOqfQ6Kw0k/LJI+d/vvXF1NG
7mvVh7yfntRjUZwtVIEGveD1HnEjPNNv+JXMlXU1f/cNkCQrb+QcqIAU8Bz5A7JkMzpFf47w11s7
TLelzRC/o+Q8C+djcZwChR60U9ccY3PETPbBc48bRYD8wNI22UUQfNJXmUWXb3HrwJATQ1wxeSIh
Te/DPGAK/xLB1m0ou+OOOwa1+bJ0sMrigcSr8ymM1Rlji3rchoXFL9cSQ9Ov/VJczekFvg6y8gqR
ZnHwZBZ4o3WxTU5MbFa6phar+hLMwcA5j7SAsBLFsrlzoHAnx778cxyP2zHiSrblFlpFe4hj6357
mBVLdiwcAjZpezsa+NOxza9/cHE/fU+pUa2bw6KDGlPE2ZFQ3CUQNmqltBP4IEXpHH8xPQ0hpteu
s+EQWAz7BFEdU3I/hzkvP5w4vWGRPT2CVHm6VQJZddUZmwUeuts6GHfM8Pd94xnb5EhHHisiudV9
haGZ2FhawksDkYKZvqtbzpN00zBQFCGkm93XlNVljArcHrLYWaX966ncOxT0WCIlyZjoxSAU+it4
Nzapwvb/j1zSt/8ZFL8fnyzu5Xet1cqu7VFii/fK/7qDvYh6+Yn8seK/B+CroZQ0iEH0klnPcOAG
mnPNOnXuNQWhDgz0E5G5B2Our43aCz7VHVyvURXPtoy7P5b0WnSiRPbERl8u6GMFbVdnYsOtnjn0
/gVCZza41QxsK8zL6dql5pk5sWJBMaSLCLg6G3gBSj6VnJLNVxCHWRrjcQ1Yv/AUxAQiXGjF7L43
SmZR2h375nWcwMlE4pUSWXrtrKYTK/FTCmwhVjFct5O8rO8mdbeBv6toF+aZzUotztqYregM0QBv
wTGBGgDm1A1fV03nmX04lxozdy2FDYO9pPjQPEEiM34OqnjC1pH+iXdBNQSHnoOgYerUH68JqnPn
tcKhYQod9bQTwPYXnNx0sXHTkWgj4c4JfzPIDGyiq/bOKfjlGqExnduABjFFUEw6YthmIZiTBq46
sXUAt7cjl2Chxqwsj3xOc/vBbSFIhOBJMlWWEJrTyFApawVcamM75YVtCZ2babRDoR6RowpCpaG/
iQp+uysAqLw7KTws94uqYLv9cuO/HRhgsxgKm3g54MIwXC6+x7HbPjomIEB5MNmcuBsI479r0j4z
ayMs25+2gAi4NxfANZ+pmORDIBT8FpfKxD8JqweXGJ3CaTgiRYDys5UgWm2q5aYTKIrpJ7XR+ltV
Pf9zTBAOaFecusj8uqSBDTK8TPSr4UqrH9URVGy8oI7DnLcsP1IDmqJhHrLJIxQtLmk6gFweD7k5
pFfiEvL6jzlPS4dY9esf6P6MQd6rj2U/m/W7Bx6qGLjNc8h/Yu2tt36llDff2gVEUR7atXzPdG69
G/Xpb3WULD7D0M+qUk+pWFM9JbWXTLNfMAd6aUFhbApFzZtRMeF2COXIMeDkmfHGWEyWw125ZpNs
tgxqIsjpTjouuxejJJMEyffAyskgUT1KavNqYVaqM7cMs5omMoCAVUglUYqz8cgw65TLuqElomS3
F/FrHE03cQ2VLPtbkP4qLZCzOQFWDLCZ8VsLx4PX2R24O7D57Uq3nPnza/zdqZjmiLce6pKZUxCq
Z4VuFGKDe/SrLBWAdE6A6TRXo8nzk2bQW5wsaVwtV27fdg+/DyGNo5sa7sjZblmEjUzc1WQ9Tc+Q
tWcA0vwe+ERRzCN+ir7EC8UYg4NutmUGLSEYp2kHKKbMcRmhKKZyznbJvv7z0ZprJS7qxKPBIBnu
AaF1pYJxZmc/pC1pCf4miweKFglEeaTvCu+F7mFiIGGrYoygTbisyRkDrDGtk0Mu6yM225o7jHk4
a95Mbfse6njWOGB+DEPXCER0ThP5puCNzlA8K1nrgXSBzu9AF4auTletcraY+UwlCB9Np8m4CZRa
hbIWaHeCvGkneYelcAtIfAWWv7I/a96lAKeT9qAV2rIhgxfohcAqcg2eZam0SMFHQvgjXld0JQM8
Y4J/szZb4tPqtbgaxZosd5P09buiKVObSwsvBgszoey7St/oq4WItQMcF0CCjUBvbeR6W+zn70Sk
zTYN7xiJ2fzNeig3J+6e/10kccJqFu/zFIUyfZa6pHUDjaI8BjMEvWdQWSSFKJqih9PLAaSeN9OP
20VrOWH8f/Fv5HY7AYAsZ7KDGIy2AUxf8efM0u8hRchEjzR2fMCy8mkS1JD/Ciq0o9DgcyPk4Z/M
nqxtzsOxjtS/AIy3F6fX2Y6hp6bVMYbcYIHTG8/vmTV84RsRp8GerHVdEp2ghXN4/es3gnj+2mPd
wmPLUejaMC53BKqVJn87aVyhTa/2d0XnBIFVufiNTZ1oiagftBtn3yp1U0MysjUZocHdxGecw1RR
jz7jrmiolGMa56oAwkQKfLTxeKoRVU09xFO+LfVzyxUlqCqgb7e5KcNQE3sdyAJDTIu/0g+Nl2nh
co5nncsU+xgToYt0K/mByN9wFqCiNhR2gD3qFKhg22Xi3n6x2M7Q0WBfl3iVHKZOISQvKxWj+AYz
Dru+6GWn6wriqBey60SuwRledGjj74Er6Ig/0nPUDTp9TDFbhIe4+/QS7p3ECDt4/e78uqspTfVb
swNTow9DZAEIzj2DiKdyljI6yxw5n7a8N1imdAH0H7eMAywJ76SGh3lG2S+kk+M+us2I5wf3FgxV
clSlQLTeRgHvgjXSozcedrupPdBIwGD7PgsgZkctzzUd/1k7Zz6sAS0kyXJ4kQJYVamfdXY2nAVZ
msD3dWD7UEKfteoau/LcThukR9McriXQE6j0nXBJvsFyyzDqNtwYpJBpSn2Cjqry2+BTZEEqggIA
sw2l+Uasxl/4RMw6Is7qh4ypeoo2IsG0rmWMmFFoEOvZHyWJkYnnuyBwpmtmXM12JDqHLCjBPpv7
XgDtU6lU3tzx7K+uxZY9v3Q6DLPHbeadzBu0v3TwG9FT5fh/YU/JTv9yjx+lnW+LYYbggxxlg0QS
xW4ctQ8o0MTEDWPduDR/tRT5u684Xg4Twa+QYSvZFL248UusQigCl/W4wFfCiQUdEEYsFCAfauKr
zuwUEImqUg129ptwkzSBKyQleeIN3o0YmkzcDPC3PWEkAZidAMzIIUP9AdU7WPa8VDrEV5Tz83P1
e2n4LSdYQ0sHVDjF8oHxEVuxG2WfXU/iMFkN5akwdy/SvEOcak3LsIencFd3lrF5L4znHyXQQ+8B
dx+eAL3ykj0JG8dTDvwxDBxLnvLNGQmapKJGALffsKZirAdGWzL34pmQGYI6DFLQoR1v4n7glK1s
ZJIVuUGWXQ3BgqwYbxIDXDiUt4zsFS+RN7MDqXPUKbg42HyELZ8ThBrl0SHwJuILY45veeoDb2CN
Z9LGW4ySptSs5wgVQpZGBwCoZ/GHBsgqgdFow6pwHEqxPl0ruADFdj+U7eoief2qPuTtjuuTnCsA
4G1ygFIZoYn4u17s6Nh8jrP6cGcd0t5tHoS9DkxLipCPy5iQrEFM0aCM21yfkYSmS9HWpb7MjQ1Y
CSRXLJ6EdgK25vcD9bqBdHquYjBL40mFMC4umloqTLoD9KVRhvDFKNyonPDLS7yziS1Un7R+GBNS
9i/J3CigC4DZELrmb9xcAiU5cZTAFXD0eJ/YP6xypPbZlpv9X1aMFcd7Rl5G6JBbXlRwDWru8bQu
PAJFxXBYcOqS9h4msNi7hsU8tPYOp0A6U9cHSMl1ZDopqCWoNPHdJeV2EmWsSErVjWExljyEFmSU
RusTHqJW27wnJQGmi7teSW5pe89lCOtKJ1Ofa41TJDgAV3S7IZLYMb0qyT5zFe4KGdQ3qWZX0MxV
OLpoucGkt/zBUKJVFgFF9irnrhFifPNtI5y708/Yvpq6sOiTxcNJEF3CZ5qgLkIRbk+NlgLRqsmg
4hEeMeCH/+JZPw+86Dbscz3lcwrMRHb6GP3k/321BOGELyKooIBDFChVZ07KPYbDMfj7d6PqLVbN
A6bP/hRvHoJmkDzSoCD7+Aes82kokfFuJUlCQ31q3flZWpgce513HZc9tOJP1Qr0x+0kq/Bx7B6s
WDFJ9fYJa/7csrcwNP5h8uN3OSwQ40HgLF7Gs2yHpGnXzrQh/AjrKmkITvc0/u4s8/zPH0bGC7li
Y3pCCZ/d0VJiedGxm0SjeiduvIWCgJjSIRNhUd6w2TaKZ7qjwXqgpp4Qxwt7V8nS/09sJ/fQgRC3
bn9h1ZSIX3eA9C2R1BCMpBYM5jCer20t/zobSslTUs5ELM+i8In7p04HBIltT6r4PXor0S86YFpt
Rr2GtdeWRvEWBEdly1VdalVMHFpu/fBPbGZIZmCfymcxsaEd5dR19czwyDU9PVv0zWQ29lbjzwLk
jT2ani0hEDX9c6uI4igYn1YwaJfc3TqG9kHokE//lw5LIqqZ1+hyyL+itKjF7FUS4bqHcCL0uX5V
G1P3eAq9RLU+yEIAW5/6GN2Akrgh3qRF6eV36e9At2JdCDL4djqauYYmH2dbS43MCShP2CYJWcfz
54I0HFBfVxprHaxPVLjwncRLMmd/naMHTnxuImUSNNhzl4Wk7EX+pG3GuWOnDVZmZy2vDqppe4mt
G9fF15whb47G75ChtIm6bp/4Zx47r3NbjHKctXc5H53JuozmQGFAhbJcfxmCMclbayYNStOkVWrU
0akAeYwG58arbsxMdbXDOt5/A7QPrrPmS0drSaZdwky9X+kywvUNSK5K4ZXFJZPyQwyGFX8ZkSlc
8yIjDTfdQefDJrTbzlvwAc4c1GqX/Zxp1ryMFmF/n0baz4k+T2AWLhn3WKoGI0+EzublG/HZqR0x
jrRCVNnFQ1VIcPYWqmcKZeWIb96P2JIW/u+J/5f154giDIv8vXoN/yNdUQQYWD37w4CxOtqRwmgy
kWZXXsK/Y+Q+WzBKQ7CxT8KLgIhI+WfX0YyjmKu0ngfGOgg5vNXy8/kv7+shHSyhkkh1SUhjXNuZ
cgmVYcgJlRq5K2JFSv+1ArGBta7Hx/YoEo81i3/r9avAodtKlrkdgtFZ0MmfrJ8756SWqUUF9ZvA
U3x8aac+6eFYe4ooWOsqveYKFrj0f6+Naqjels3jboJmrdgv17m6tTQByWHjdbQRRZNtcI1HiRK6
iIH7i0qk5vIFevBTcEWLdUqDwrMh+25xHjw5lzGItNVi2tHXoIiZ6G2Ztj4uqStbgGl33eu2BJAP
O+fH7lZDmkVjXELv5Gfqlch5BJWxm+I3usRpwCfkNNCa/jQ0Qnhk5q+FGuU68fHc6bpXvmWu6VRn
J29WXbpVWNz1HArNRY28mHY0Gg4LrppYiClltdL2bqTPeaofeIed5Zy80KYBCghNxaWE+cF0UcBs
ej6SJfJ+wHQhen4rySi8RCYcLzV1wSFGL8I+IJKXNmhSm5p8lBrjVSYVbWLBMlNigCHk7aNGHgse
c9RpidKMS4ufZh3sh4E8K9oBUKnjXlYM1LsCsxt4LaA4+gLHtV+plL+ug44ExJ2lbyr5LZo6Naxh
W8N/k06x4Gak2NjWX19LGa7hg7jhqoQPufb/POUC1YE+52X4J5dsjYsdhzIlvR5SwfC0qpTzUvW1
FnXT8zuVy3mZ56aAY+FJaJmjTD2DfrDlAI7VXWgH/8Fd8mUNwKAH0pYPQP+gOkbRUjanAVP/4Oaf
+OHmVCrt/bJa8eCHr5raCvo0QgOM1cCBs2pj7fIm0HqSxV1EM+1EYDpccUGKODwJdqFYIbbwVG1i
xbYsBrPHVM7imiJY3LnPIzFWGBAlQ6UfDEz4elJEgSY5f0MdbwYS48AeHoPJ89iJimy69ztGjZgR
PJGz+yyNM/dt57zIhzzMb6HbP0vuO+4R2k7+ZJwdCmrmFNgDlIGJyYqYO5oSa2T6FOG9okr8TuNo
qwkIvf141HX7ItU4WynRgoP1b/IdR2MqeJNOzbGyAP55iZvrWXiUQfLBKndP/XUkpEgDbvNdWOj8
Jg1s2EsG8JiQ/bxvPO3Fkzc/DLYz80EoKkrXhjRlBKELDAcJZhC51ZCgBwWTCwZyc1j/YYH8i0Ag
PRtiNNNhtnZqC6e2Obo4zA0uzCVhVTJPGzKzb8qJJDa3JxMbtuwEOL4EWijBX8l10uXUMetTREYg
nTufx5JEpJs1UohOgdFTB87zt/MTjAxEopFKB5v8mq2rnI0Ng42V/yFvAmXmAGXv4mlni+Mr4d+3
bEe5GZH9NzlyXkKf7bl9mPtz99HYymoSIOK1h8ijx6WqHZ12E+JoLZwDIrqJzs6bomXWvRYcbTQ/
iAnlP4Ai97zwNBsEw8rmH9t1L0RUBPt+gDF+5Sd/l0UFXVz1PYlCqu1tbU4B7RsRNH1HY5uevrZa
Sceq/0LnsTV5cMfsjrbCJ0GhrxWFsdOJihboqi1zSTOqcMJeWifzUFWjOd1YNWfI6IHcCfxrnEqE
/QeiC0YZo5Y13ZeqS7xU1dwymvCmJwPOi8Pe7trBHN1owmbExNuXNRZ0ZdQ4uN3w+YPAkva8PWsy
RmRMd3UAbP8AaC1SmGN/S/qP48zY3741RhGnHFtAnJ2yYIPCwq0jij1JyULihMXQYmhxHYtpCqYQ
e/ayiRnQxIzrs061RAVvr7FE4gJD98Nyne/rZeXnEKC3RSQDg5te7MHUk7y6ElhQzA+wWoEXDg75
GJ72hbLw1uEOByba+/s6vrDlPQWEqbixjPhncXT0aM3ZQBHHqUOLUkpC7nWZWc6az3mjDdHJkDcA
WlT+cWWeGyEDoMswsxdoHyZI3FTGNBJytAvUNibogF/qBrTn6ux/+jgo5rbb2byP2kJQ7XDX7Fw7
FnogcuYX6nmi4FNNd7MMeryMMfcGhM1vSgeKBxaLWAzdR1MUusKPPX6UTap0Bj8pL8Ba6ud9hwz4
8XGVyhSENnIrq6J+Pmd2HP8zcr+w2nwgRz6qq3d3Gdj1TuFt4l5dFigL86Sr/RyFM2/e9TogNTYF
hPuH4J1PhK8hadWjIy9i9srUfCbOx99HZPW6RWTgr874kK5QL6lhKj+sSsHbzQVoXJAEGOoydSHG
DBQM5idaIRBnpsZKjHTTQrbeWqTkuACV+JjZ+x19TsMKRdKg6rX1wpIFCeHB4f+jk3EcxwnD7cha
eGA1gYvQq/5qZgRhjFf5hYIdRA/lz4N8owUoE6WsxM9CS97YkbUDZHEnVgIAZmKVDDHc/O+swF0+
isumLq/lfNePmsOcW0rCbjy87MAr52PVkeqKbc4OTEVDptAsr+/0H4UpsxhxM9tft1Tvi/KpmIzL
6Z61nyEvBL06Yh+Wcj/jryL/IJbTIjaHSaElB/qiv+m0kY5AE1nL9PyEpU3W16nMxmG8+XK7E4hl
X9238kkt+dOOjtdpadgvX1eZNQl+lcqlnIamy2NYv1jkVSjCwOjef13HdhMw2R/z2m7H7slynqM2
6YN9g9fbifBlClj9M9yTGugKFJd1D/LpTWjA8466MUsjggkOqhq9hcYRPddqgZUZTJgnjp9cyUNZ
X5w9T1eQEOh0aPJod0Q1YtAhM+11+tGUNkuecJjuCiuHEedf/LdMc/ET3gQpWyB144asZIvocnHL
slRSZiIJ1cOaICogwqDvMTbU+iC2G/xOIEILAkgn/ZwoRyLZEUuLqhcfWHIQwTim+sDofgdHbfi2
cdGrMQVx5I+nyq4hNDDqwvj61zEv9cUapAHbQzRYJr2nZf2QfFGX8BauxgcVIH0HT3+dim7z0ydE
tm6m6VHa9eyOJ91+pES6JaLjJAuBCeKdUnPMWjE+8ShffKrK88xSCuR/0+GnseirV88ih6+7gLVc
OH56JEe4wKTjCRKl71oWYqPm4xYXuJlNlUTePmykPCgGuDKac2iuxg6u4XZqbeeePP3E1o2oJM2c
M5PLbuhE0rjo8oQB5JEp53SyA/CmpNJXgawuME65y7iFU13K/CCMRs4Hcy1gRMxh1YqcdTf6nXSO
1MjNugT0mm5DPB64M4FVJT5i91PNIoWNRYCKHMySvQXurJySMH2BodRFwSU86jaFiCBcB5aNQQHa
ga+EDMqg+mXsomC9bLU8Vsacrd6n57ZxvKXoiQ9lD5Nw9kADTMITOl72yj1mafNgI97F5HV5rcxi
fp9911nBh/RUN6PVQ4QuDaBzBOL4An3l6R/KBTOFBubxh342hiam/okjPYxRGWfujUDzowxyYrpH
rcofjAzHugn5UPh63Hc57tQEmeQNSkJ0txiCdQp3hHJaE4Xwb1B0IgoEUTABWpxHKiHogIqxB+X/
zD7IXdLhk5r0DUkSe/4ADzjESqWEjt6ZhZcyc4kt11GG2O16xKXq7j8Ait+sjk9DTTknJTV1/4Ls
w0yTtYslQBKH8DpXf9b1r71ZXxVRkUkAClRYBB/JdOD/SMRN6OoR83GfzOh59QjTZt7RuEb3CRza
QxhGHw87Ls6k4bVQLwh2+rH91eGubmZ39/BQEQUVElJ5bZCzqkDb0/Bvyq0YseFdSs2nRPi/gRFm
OMrteoUm+C10SfmZTHcvKGC00mqyBUgFK2upVFbfMqdJ7lqAaaNV866zHYULXCgL0+TStmeLznVt
s+kr03tTGcRRPAv+mlk9DjkY3nHrY1YTembqPuVlHta8ZlURfIEkUAFOItzvFWYvgmJxZQ5OSz41
jHyo2e6yqizRZEpcKwk/Sbn64v5s9pfOqu/cL9f1XdgAim7fBYKSMriMZt+5bwX3Ef6OWKD1sj+8
2o066JVV7FCLCIWDSJSGhstBas40ainExot5kxhjAggiOV8Rz7o/7D0mqswoBLTivSwtVqy79dh/
XmcLuBIZlWggVrvrqD+fVDjZe+DEZ9NHjuQIbfa0yk0TOlQjLK0j8iLPnpRncPKOgIpFMjLWYt+x
hlM5QvYO/+6eUi9tbVTTKcoB6afnLNubjUzenXPmMKJGpf7YLpN54JjxGFztwZWtp3Nmi+vg0KuG
e28jBJvJFkQ16RythJTVumrBs+f019nxpFbnKw0xNIsHa5oIvWR/u+zYGqDUevTXGDiU7mMOA68i
Q4Ddw8jMjVxtw14E10OR+i1NeEHsPxOaG0X8Rcd4xzXgYqthrHh8N3KZB1Xs2kdsx6O/5XJFNBoZ
k2jxwKO3EAu94gHQwcY3pI11k2k9z9igXhwZW+QcF8KRvHBkxSt5GyfBggDEqbA7nlrntzpb1Iym
noiFLqRHEB3B39dhunvg9dPQPnSXue2UmLChl8HgNem59usz5oj1QaO+OTZzib2441vZ8Ya4P6lO
02MyTWdwE5FS5vOYbLUy5cJYRTAmeiQ7aqzCCypdfnH39KaIczL7Yi3VhKt4qzpmJu80p8WZZgjL
bGqCiD7BSzzSrQLNnCg+1PPSPjqAD5V89EXBuTb5Oyy6NxYY5JvSJvKwVGHVy25xEKWZd5H4MhOi
fOXLGwmvrwK41CYF1R5tr6KRirnQoxIEVzjGwlUF7/93ZxXJDWp0JbaU2udPwaWh30onXs8svJPo
SZwjozEc9K/o436XYE+xcianeB6YN8HEL4O1stX8zd64mRyKcGjas2yUk2cFjg6l/+H72e6PITMr
00eFUBwUmmbP8HgAfqkD7hr6q3Empx8gJoueid0FPXtbIWZAffh25KHDILBpsm4fYrAbLQB81lU9
eUdQPALWSnJtLI4zvGXSbVS7Ra5KCF1QVaIUnaCC9SAr62reuxakXGYxJ2JgiHutDCYhPlNPsIIE
9JbmKNMwPC3Ilb8Q5u3GnR4bOMKHGFML99/F16Nu8FQjOxijXijk5q3ACSqKRK1IC86SflzuSAr/
iT3SBViH6csBJNdV8+xJHwE4KNURuggk0VEvrFR1IYmzpX4CnpRGxnjNDC/2Xuc8zJPcFNzL6/kL
pHTLwfGqoRhcH+bShN2ZUCjsAmyPJ7Nzb8u6jOXNDuK7ChWm0ClKrDLe/k5BE3DivsgvQ7qFSNuJ
Y5dvzTp3/ZjAmX6Os+Af5kK2HerCZCNyI1eHWHpYRgKCIkaL72wDEr080UHISrDSXChVzAakbFWu
GSWhLtAYb3ttwakpJGRipK2zhaFmBgjOxgSO5uqSCUTmrLjq07zWqt17/HzSpdXdFp0IPyvGtVG8
vf58MJfV86Melw7xgPjNj+IFAfNBS/AIHgQWCwrkxv1R/faaRMGRXVTiVd/EPeKFUL/RjqjYeLuT
2vi8lyElsBAh2GpbUhidGyWs/+C9v7L9/TkEe6Bpeid/je+DDa68aHSFwRpRUkHPOq6Nm7Svq8As
rpO6JNYEVuPjqXQX1EH8o0zq98tn3QKf2V7a1p4un0ktctwvF7kbNCyGG5M/0wu/cEuLO+glt9tl
qdz1xIRboCcd7b1kJJYA/P6OszzlrnIn6LbOmKZXXb8Ht1H9KYj3vlg1vMQaVu+0pl7G5UOwhiA6
tXNGBkKOdlTual6unGO9dpQGGnk9jdBuPHXbnQe5DFr+ccG2di0kvH+mrWB5uThCRIV4rZDN9PO1
GzcLBtzEGu83CJUYa8+MAySRkXr+IoypYPwuORs7OH+ZFrVhgG4T8RvYIN9o+ammcuCbJVePDfMY
JPgm4GpFgoM+CSyXpd4OohqK1mxILDOij2+xIlQ4PUdFxXkXr9WnQy0aQSyRSYO9ynjI6pfE0g4A
Nqkx37qQDABbpucQEGFJLhly+6mxi4u3DYfQMLL6hpHzoKjRR7R/7vqm3pT+uWgBSeWLRKLiDsj8
WaD5ZWz455ZL7PspTPNYSZgw2GqCvhRqBAyw0IPFK5s2PDejeJyWW+KOfQ8Xav8eE/nDdli2jkp9
Qr4B1eS6mJvqRFTrLw0OVR+wLPBZSKgLQu34RZCo/4211OLfCOyNe475D6pGZWFWcEJywddI/uPR
bubTeCKUVUMxHVqq98KctmLsxAJoioPdvzxI9ObCXMJw0hDiROjo+ca9mJHGsujvzxy6zjDcGJAC
9kwTsld56uRKWRYrkoRlJg/1MU1W50kxEBUAmoeSlQxhgqEyX96DjezxeH3PpbkJfR5YW6viWP+q
UBQy0LUjDuiRHMTbdJJv6Zi9BOj90drUUfVK/pjQ/qIO1YNmQNkDre8aSNpCP1HzapzRNO5Z1e4q
2/qpLoWJADZrp19eut0ao5hGFY7haL5mgvGe2yLH/NGqpX3Szz7yseee5SSnYct3VDoxrcculxSC
13jDllWRGfN/dAXBIs1l/WYPZHAfFc+T2IIIdx7yVyqpehd9bL8WG5hXQlxWmsjmYVn0vUC7oE6U
mGEjXdokQC8+3Zd9j+FB23V5xo89UvFxFRcC03inGQYN7xZzhQPEmBmzLJue0upuL9xB9EAHnVAW
dyxbWLy0wPPHqZqlTRLXmrySWZa4t2YANhUBDNYD4ymsNZOGkyQuH6oezIsve9+e74rhCkYdFQxU
XTFORwCLLesR2A9B+YzXgjW6Uh7N0Y/R4mO7r0bGInHNc4fmia0IEo7qIM0qUKW7h3EuIANY639a
LFHTvdoIIHBbn/bMdXWrK/kPg8k5rfLFCYh6Aq6fh/V9GhDXgymxDOLvt0e5NLqcn+xF8jKdciQu
DspI6mqScsLuouVHYAXqt2ojGr2zGc/UZVQj9CT5pIYzyp+jYezDtBhtG5gaM7WpAr6DBTSs09cQ
JGo2H74EW2g0HUF/+s40JcbRDEd1Zkhbs06FgtaGox13O2rQ/EA5xqKxv4chwKWqLmRrf/on3IgF
wRBBQoN8mFawrZJfNu08NQPJkgu5Q4d67tjktFNIghFFIFFKFGmSxrDJeD77EDrjc1sFg+82CmuX
+8PrfTG+o24BX0WjseGA5WNLy4DUGBOjbhoUoKQXt8w/P9bqfz2G+PmBDXSdgy2nvuv5rRxjjzZi
v6FKJoA+xHlv3yYvtabXCiUfzuwojC98Y0LgskPTdCGBjCPZrZlrmIhE0sDZj6m1SspJlxp61yGW
d3uYEkxvp0ypBS9rqPJa/2eBv3fIffqthl3hGBJabTRzDi0pj/bSJmTHteZaVgz+2tRQeCXYDHMS
xARlvzsxOHzTv1O17VgZI39Drau9g4V5LE1vHBStWUjjKKxqEv0P3V5gWkwI/dvF2fAKZFEb2Omd
I/bwrY+rEY4qERXlJpqQU8k1JdLBPpOd7zVJadKHLinW6HphKzTW2al0XoelbVefBpD2oj25NdUb
vT7cDXAuQsPNq/vvxnK5aKnS4BJiKQx/cP0HYsIBuFRshegfWK4oYcXDoS4GDRV5v4dRifhW6bL7
pCiwoe6LgOi6Pu7qFScleOMeSx7kWOTZkEbPCX69+u3gsMSBw0FQcOGqrkc0NoV4dL1DmdSBBkSN
zWC6YtRdzBoA9kjnYp9kpnqnfTSZzTdt3HbnzKSZJ1Wy//7cnFgpteB5IGp0+ILdKXMbLurqreUE
nkRN3wG0hSNPE80Y9nhyT2op/j4Yu7DPpX2+8ruwmAFf21yoJbNePWGcAcdOYu/uvQuUNpg6inCo
6pCa1mwsHtc2dXV54gpDNrud19oWr40kpL6uUNnlcT0WvLo7VgC4PX/Vy0WIr0i3N/m/na94DUT0
WwYoOE+GfQsX7DObuULnByk3Co4UbTTkBCkJfoYoEnO/G8hfUxXFpi6KORtTpmAZswOBP7VuyN45
Q7WvvdgS/17/RAwwIGPic1cnuwf87ZyMbbfXL9Gd3TAVpDpeRqswcD7JdjezwKxxk/+waFoy7PrO
ECrEhMHbZjsqweTpK40g5NPE4LDzzF8PrVybw0ege362YIAEJBuNNh5SR8oWMcgnUjRRnpAPeHLa
iNRv0WvnVK+gkeXYBgW+aH1Z1R+BXrtapny+qY9X0+EBocNem3JnQqduRv76kucQ/7FZZLNMB96n
WJS9MAxp4PJqIqrlsWxFyY/bjG++FJXvJsAuMhUx1auRerbVCMzFpRiZC7a2qCOcUkOvcUigVtUN
2iSwgdeSC7b98KIB5ts7tBcLibPg6a5xGF++4b7MjCoOh2shb6uonGXVmYcyJmQ101U8Zx+bs77O
tsLnskrt+iR3yl3Bjh0/CKBfPjO3LHeRk4FOO+/pHN9bOY3gwsStIW/H4NmClyFeVDL3gQ9mUUod
1IS1gWm8EaKpO2tpxUEuvjliiIN//rVgwNUzImKNMdSMzv8oD5TckTYZKlpnznWRYi3enyJzFH7k
UYTUOsvfsF0kubHGtECj7XSJknA6hgS6tZ3wXzGbkzhOJLkpQs1iMyJ/KF8Uzwqd2RYqQ+FjQMQ7
C8eH9mxqqrplOdxjf5mFXtpFN/YLFX9lU+YzD7z7gnHtJkgVX72m8arwwXxIYyivyuYxRI1ar49g
hZI+vDwCW+ZpPHA0weasf4gvZMDhCFC4uVy4VubMk/CBOnb7Ha9DBKwo//xeuqeRlOb6QMaa02J8
pdJ5EoLHWqP0x/vB7qBVkwW/TT7ViBdZuRE5qFODoDV2KH8Dk+FWPIh5g+Lik3JHiJQa8CU01ULF
5Mfgxvlr8sjNk1fnW4Z74tUlyza16vqTtAFmMnaI0E11mLolPGGNnMahn0r2+dI0HWFnd5aWmzvT
ZKQfXqvfUr4wrcPl8OhFfg+LNqsP4Uyt9epjKTTCj/L9XusxzBLYUm/+WU//FRBr0XWsPbzphEPP
+C9OeS7g1AzCrYAfSyQ0mC89HxMRqukVyhooU4y+HB0w8Tc9xgaUr0jisM7EyfBvTuVLBRvSIsLQ
dBFJlNIrO7YKHdrt/MD3f8e22H8XaQfBXMRyH4F5ToaVoovG5I7Hg/77EY3lxsZS2oP+pX/iWVJK
Tbn+B6hvXJudV27vrtIxtT1lw2qG+4vV+tCS0npccWmxFb6FJU++FOLlP/knkpIL2UyIdnak9wZB
bfnu7PpSj+ZZnIal+H2HaLBZ6JnVt1VApjcpZQiwlmmboK0kIwo9ISlGLKD2uYEYh0Axpzv8o/PX
K6LyWi1rPFECQHSonM73wszNAiJV1O7dtS0BldY+Fd1INJEc6JD//HpkTiRXDVdUrccZJy14r+lw
Z8wu+Cz7MDsqQt4YH6sMoMk90RE8+WIpbzFNlewNbBQ/or4Bu+E2arTp3wYROwQgYxYVeGQuTJiW
8KdkRsjluY4MLqMca2Nj98AE1TD3y5t7S62xTpLLkJdWkrfLhZ5uhCcfAdEVQU3aBIJjLQMuerv7
/GBDCTuDcPINdaKmPXKV41Wh3zCT+EKUikTf74ESBEaaDfAIWXY40yxSZYapvt8o6tIht8PmRm7h
6aysjIHFGnQS1CbugB1nfN4aX0/kUQtaVh/HZHTktdiRVGEkzj6eqG+WMseEYta+6WlQkTnqmFRh
Nh8i+poMbZ5TvthuvxQO+/gOiKVlgrxDvshObjPE6SDCPtAbh+35Iv1P4IQ4U52A0A3Ma6f9Zp6W
co7/3f/Biur/Kkq+HW7UaRGwgt+Xisc61Hy/5+z0rmAw1JW9fKjy0TUN+uXawIq3rSPcK3xXmuC1
4teN1esyuRubBMCBgToYOtYMELXoTkl3XWaxr5Ci2fRyPkV299ERKnvb4Qusoy+grsnWw6d4Jube
uORvtydKqshhJiiyiGO4/rJdhVyHH0vJlUq36++LBBNEFWuFVx+zOZjfqgCaz3Z4mECwjZUa/pzg
84caRe08RX6VA0bBjI6XMjCvPHcBywLJqXCe5s0dEzlKg61VlPc+9cpe7U1qCU84uXBOXMBUGir/
rq4hotAzxDdW5zgljxXVilkyI9PtSVr0zmJCEqx0SWPq0oHyvlF8bdb2airBoNpxG2MLadOVg47Z
h9tojnFWzJ60lkbu0lSqFZIiQuHkgSjTHAAyJvl4hm1tBPfFFPWIhujzlH8ldhrRF4/UWcN27dsc
81Uw2vsMyo7bT2N1yVvT1xTJdHa2gxoaBk3KvraZaFgJsbK//YIkjz8Jiw6414gcFWcpwsh6IOkr
DWgku1bCXC/UqN4Vcp4RKx6fVIjRF+7STNIkaPYMsEAH3Aob/JOfYHn8Jdhefaaz7d0rgTx9A73M
Y9kqnK+HbZOdPDNI56f6uJYIcDe/K3uMDIYMCoSjC3eI5v+RgoM4Icxhb5NNa7TXnJrlKUR62ZUT
rnTuJr0lKg7mmQxvouau+T05g+SOBjqf3XWNGh4sfrF++6PdYa40RimqhxO2KWvfhQcyNMQ7rBmu
2J3VaJJuxG1r44Xc7T/zgxUc7Ov9DxxD6uY0jty3ehjYreH6cqi8Ywu++WR4PJz+mGxx2djyCWAX
E/9bZt8j3FbB1aSxeQa3DSGRFM++537L4FbNAE0WwsZ7olOit3aEZJQeVRGFhpp5izw9R5mldqfC
ZNagK2Kp942Mh35JBGCOryg05ExxjFPG4orCt2Wqp0YBgOWzCkFUNw7Dc4yJcF1eYjqWB0qsYjmd
+DyIsHZe2x/78icRbPCw2IVJADxdyxzn7dweR+/OiQVGHh1ganLU2bJWOcABeLNO5p+a9U3rHKUr
DCqCjg0n4rVzcI4qe4EtfOsxgD7LYAut+IoWvWVcfchsCVCVAQgyN/Ui6m4UA0mHKwqcgx7VMtpd
lFW2VnGoYgOQCCu93e2sRvWXFc0hgI90amCCqj4jzVw83LNuQ9yorKs3nlhIuvCxz3hz6rTgypXk
G2gnRzWFAXyufY226N5Ez9XbZN+eBRF3cN47k7AYyMuH3pC29nuWunjE3SIyKZvm/ecbq723xcXw
RaRbwqooYvvVphUWnk8gPYW9YrKpk0eZngwo/YAYnfXJOjIrC4TvcRlpQPh+9tZwW/lNy+dBcV5n
DQLeOEDm24ZK2dmY/uWIGoa8t0eqqPJFGPwDmZUWcBxCMdS/vprUSxRaMTVcZVdTFtcNFKPsrjTK
EFhmf2yRwuruk5oZd16YXBOxGy8YgGG7nRI0ORD7v5zDYGARApumOmHnU8dqULQPMUGiVd1G4Pui
iqgYvXqfpzAfMnL520c1679TWOF3IXWQMeKQrzUqbVm1b3bYZTyovEHVYEdi9yR39hm/NJ2KV0Y4
zgHgwaxZIhnJKKpMlNYni7uSkvEwuvRE4DNwDcsM9p90lDoDPBI+mDNZYElODbhJt0Dkjx9P1J8s
DhwvrjcGJtM/Tq+ZU0O+Fh9sv5wv8FxIjX804/WiM2s7ZYhlOh6NKh2Zdo4Eu3oO+d93Nh2pvdHY
BP/ztFe521HrKXA+BUL/6NACV7tXYYwpukuUWG0GtWmaPngjzcItwJZhWdv480JPAGmS75V1uo6T
OTgENBZ0s5dx4gaM3sNDD4wN+UMC4pQ3XVZFWSIslujv7CloEY7iB0jCjKqAFlE5idxHBc3pcNce
TR+mrwexqSQWap2Am7FDot0sXKb1qTzPKzCGQv3CH/nw5/rGXyV+pNOc2lGzoxtulh0zaIjxCkuR
9RaLZU8D6VKBv2BYdTtVEu+zPo/3FQsIGnu3xdZT8hIntlFPUj8eAPnWbQJkcvVq/YIn7WXhzLod
d+tqDVlRky6eKqVYCjCXbnG+dUNBxoK/qvF5vpMy3zDowCunvPc2r2d44bnOunziAA8dT3eQZoUC
try6SdzjG2xTRNWA0BY0ur1UkdhQg3FezAD6w1m+86ad1x86qO7lyk4hs6vY0yz8y5C1AixHt0DJ
saB4Kl1AV2EHeSkmHfAlsfCr5OtxGgrJduzS0pzSAIcGm4RUai0HFFRf2juJSblYNYKLdiO9lu7G
E6mIiM0KNfWGZ4OFSOnl0/kft/XzXjl4p/SMrju/FmTul4QVB6bsGh2It5jn5EomvFxxr3mD977Y
hKK+etJVkmqt0mGDUXy4inmlbsJOqheoz52Jv2v5V45D4lx3KOSM8QM8NfJyTcsIfw8Vmr0tnzFI
Gbh1sXFs6LZWAjAjRRqpGgMNbY08v8jk3WGL/pRvHNdG98wO3KzJ5c/Hhc1/CKAepoxK7meybkIJ
GAvaE75YAxGIrF+FG2QAbiJdPfARhkqkGVRY8JObE49pBbjaDIXkyWtWqhPOmW0W2LRVZWUbmZJC
H223bKJ0MqqUMji4c2//+MZU7oycmH34MUiGWU46LRBlwOOG+SSfVZucp25/Gk/LCAT0WQEkMaKI
/A/V92sHugCFrcOND0iXMBzquXqSrI/jL+CrAuR3xdsqnzUH+x5iycBxTK+yJYAOxdn/Pal5hq/4
7yWUC26s+bCc84yrGNncLb97fWKRhSDPRZbQ0yStfSmBhzzwVl7q/Gh0oLnDF5Nk8E/Sj9p5hWBg
kHpeT/zt59wdg1LPgDU6dLug+Sn32Akr/O8gglCVJIz1V8UXmmk6v7wvCvUcrVnGaBD0/MVxDqxO
EQlEwDgXYwqbrWInsTqG5Z1aLx0794wD0JRKAg00qdsufemLlZxuRklYPF2wOzmAUhILz64iLQKm
63EgurVCzB/q6G0bSyLr6x2ng9Xd0ffvh48oS7PdLSy8C6P5SdkdslhJNnEgv0wi/tZgK7eWinPO
aGYpHx52srnD9rYBUgE/JKlfPWOC1jCUVyt0fiDzvmssZoBlcQnPmFKeeJQJ7jWZmFPg8AqM9v/I
s6tD628h4nK+5/LDuHTR6PHgTVurl3NsGdZX6ryJDAsGdKHI16IqL9/j4nAzFfu3hFc94nT2zFfC
Yp7k4tM4BNGjVGXO4l66E0FszdPtENAwAusT8MSiAtdaFXWIfX2vpTwLTYFtQOMwKUDU8S7TZTZi
8wM5xE8v81QEiDapVhpIBMli1i7fvZRt1mYO6ZswY1i4axnYDcaTnS+d1wtEYzKqSObFA6Ls4NTk
E3e4JGJDoaTp7ThA9fRy++Aqni2f6FEMLhVREqnnK9Cbg7ugfKVZC39oWs4J33CF9Bm+hfpqOYCq
eNfPc3DKBQBgQhDvfnqpVb3Vpnbqtb1dQ8WNj+uyOvhDCrZ7CfMRa3o4RrTvr0Gw+nG7rWkGxT4Q
YLQ9nvRBCqSB9P+kpjX5L6MPYxgwKIufMv5r7zKrOT2PY3QxHsIVAgRRnli0/ZgWWFQKC+EF0vP7
9WvXIo0tmXNKZLt6JNw9a/4QsUxye16y+GRgzzYy2zoExTyBJpMHkc+vcPTQolgs/MwncX506SfV
527T1VUBt/wo8W+jJVSLDeq6X8TMzOSuVYWUZOYWse4eStr8Jt6SfHC6041hUMMZ4yL9NJmKnTII
cQP2ipGTQqKayH2oGmURwjStIalROusfH1f83fCuJF33utEJRh0C/mmmySyYuIDgHSOQ88o6cFU4
MoNhlYvI945e1doMdhoMVUy8AHOSoUo7hYc1kEq1yvfMeKlxfctE4xeyzvngNMt2WmuzU+NPCHs6
YlidBnVUTXc5hOn+vyAZPNdvlK3Nkdrq528oyzBS9S9N1sYeG6edu/pPS2eqKMaZGGnLWBfiXhfD
SkXHnQeRQffhkIKb9yA84VJut8OZ3VLQTNlZVMcw2yA2E/n6qe/+prppCmLXSbFGzzAtDLMAvi41
C0FG62E7wuQkOXPO6OTGiwLPFjmxuzvYCS8C7JObYxbxj+t5R9h6b//RVoYv5s/TMN7NsTsRYR0/
dGEDGNKtQxhw1fOT5Y4JLzSD07lLey+4ytW7v1um+5OuHKFrt9MOBKSApFA5nF/azs4RpthiGUlE
6vGZ9fZjad92rZYuzBP0K2yiiuDyClToVg+qq5rwY3Q+p7vUw2Em5r3RCNZQy9cpfNALIls3nciN
5xCb/EmM39qkKpgRhsaRtrlHlBAx+tmlC6U7/RVPsvqF6sh7FHSNn/DFPtaZzxuhiSA47BCYm7eF
Kh4RXjj6NgmMl3BUZjwZae5+a1m1dzPPo+NwX60yoTPVX9ZQgzaNcGtTD2wsgkhE0naYVDXXUAkD
Q5AjZUqJQUVbCreT4wodRp9ML5Us6FruVRebr8qiNH4kNfNiWlxko0tL92fZ31wLeedrRXsszz30
9UdwmRu08mmTiCkHrclDK6060e3m9vHHoOH3VitBSA9ErEswLi6wMA+mGOJ/zzXzVQO0b7SVO7hT
8RhoWnOymDfbZu3qYEgMNA6TuutLDG2hQmFGU7wKVmvUNhpCXOXl9V7+TbCu+G91HfoMiknRORXu
XMz1hAFluFltG7MKYbwUEcgWm//UQ8Zkb4c5ko2RtWy0B768fX0y7FrHTlrxy5GZYb4VQ3V2OGl4
O1NwqEB8t4DfZMTycSQPk5VEnfcRS367+riOhak/46u4bDTsgoIqWOOv/Lt1IsrJbtSWjVq5OjWq
pu6c+52G24SgTlfgUUWwLNXEKfaCv5vXGZuILSWRyftEoVS8q77fuiRzRrypvVJpOLeX55xalaCn
9+CxIKkBKilQjoqC7jYh0hvHLjsQn3Y//aVNL2jPJwKBKVbgAIG7fQS292uZXlacR1foPG3STvqm
8vbmcGYQ5KwFQapCTQOQAUdS2xhF3wE0TB1We7/o8fMjuD9k3BYF6koBgrK5Ik3ckFd/1jRKQQsj
mZ6NimAqCbub2Daj4m1aKEolBCMlpCGnTXAfh3ZwCGSpqbfACJbNXLceGFy7IDeoXBLm3uudw7N9
GI3TkOUQhEqXyrfeZYokeJvq8iznLs7dHsjd6r12Wu3Lbv+fYbfgIFgSUSMltmJ+wAiXKXMi8y9E
bFK9ShumFdKxH6gz3orJXVJ7JiQngyf/XVg6yyxIW2z9msy/0CGy6QhERVYY3rpAtGZxS807k5+W
o76jmHlUX1y4Xbuf2GhoRNsuZ8lT83SVSDqh9CIi5tBjbTg/DROlC489qfSjZ1JJRY4GfZiciiab
/fGO7Y5iZekgePze6UgGcQqFleJKCOP87lDQDyCyKVH62COIW4Rn1joe6BOuUDiYkMsQUO9ixVxW
Rv3ASvriVCa3oUFi8IvQrnlLOUraLvMrRcPJ2wnCY0T7nJcZQvlPrKQb8odv8rDj4RNDPMqpnqS0
lI0MiRxfI7jyFNRK7HQNGFVz3q7qkGJ4ifiE0m68rnfZs4cngJprn1o+w/5XOlmPxLqABY9ydrYB
L6ojFwggrPIiG3ER7F0Y9rW5MGKj/aF+k6gPvnuFoQ8ukEDJ0ZU/cMJkf2MP19HwAAJYrtTE+C9R
YJSzwqAE9mm1p285/YhloMmYMICcAM41F9VUttIB2VxIKOnotTDy4LxjzPb5w4X3EevZCbzWv9ay
473FJfjZ2fO4/4kdcM7DNGwXw2vzTvzteNcdtlCqB1QWmvlLEoC+3ASM4y45t8LvTvYJwv78JP8s
NRhtWgqR7P/O9R3Qaaq05DwmbhGlcyVu+Y1J2CsC85ODlIQnPtBMV8LcyMojTQ683PlfHmkjMJYl
T4tSSEwRIodsK+DnbQUVYckiDxE/WB8hqQqewREp79wXB3AwhZovOc1KaHYz0yIEBwXwEzN/ERnE
wOfcw6s8oMAAScJRd4HluuyKaLlYxQfUqm4zIb7/of/WZa39VghyRXX1KiYcj+hEUmLcOVLl/v71
kk1PzCaLHTqrSyba4dWYsEHLAK3Z3hhTVn8TnupCyH0UOkUBSoHoGJTfeedKxzFWw3FEfGi8TzY5
we3M/9t6pNv/4HcoG7ZYJvqErEy8w0uFRzKExFgfKAuBToy6D3TmeHG+74BpawPT9pxfBRHUJzMH
bT8Qtp2zaFVcdzIX9+gVWC5ST0MAE3Zwynb4lWjyJMxwTOmxHmiujFHJAP5Bu0HN4nQ1kV+Ygznx
eBUp0GaTmqDk7qax/znFlMubPy/+FezDw13Q0ig3ihp2qPGbSHsE2kWd6Tlu5ZoAt7wszTMNqFHT
y+SxCmvlMekiNCEGem1ujH99dmPlKJ65afDV5e9vxBDDm+dbbCZ5D6QORKGoXjaWZ5wFrUd6aZqz
OKyW8hWoP/SGRSwVyJV2AfP4a/27jeNsO5l7HDEvIa4mMVmsgV2JJtLBN0JnbTnkLTZq0CGrBxPi
PTZ0LMs3piSnajUKtzQHs9QRRm7IA2PiAfkPVLdWqrSwJy7PP+gy0I6uCdtFDRybvOxXTMGxlxwa
IKZZkWmdizs4hGP6arDGxQC51IGx1eoomMpRHn/3rwtk+4zl0h8hbWwCpZLzUVqNSVTJ45307iNB
Eg+nb4ROlovV/eY7fKhhffpyWfCwiTYzPZabT1HJiPen/dvCkhCFM7tzSYLFgHoNfIVyNXswqecd
QoqvaVkrw29EcCLhxTC1ezkUZGYxwdWl1O6pqaINL23alPUVckIFxb+TJ53NYHVKqi4xnKMpYAig
wRfjIrWMWJGFW4N2GTl9OtxCwnGhroc+HsEbFjoKJXz/mYXzOWF5wYs8/oxGzY7+bpMVJfxu30PD
dS3hJE0JPqPz+8lC3IVhl8P1GEC9o+qTqY0kG1Ukj2INj+GymkBkg7owWyeq3ahunKNzNND8rvUt
28NtY9/LXrjsaDVfkSgyj+8XxaM/auuahOCOp0D98CN37dWJVogV6UlNksIIUcCZAKil7ymNMltD
BJrN+YFa35x5w6J3vPPoh+IYdXsasI9JrpRLT0M/EYXm0tef0tSOTdZjSNEsqanyaj5aJnBnnaUB
we3GMi0zwTseC3tIuhsGV1SJXFpMDrJ5KLtFkmwePYeWmySzfyx1Zz5N0OIf0itfLjLEPw76gaa1
glIiI1u8uDFJbBwp65bCbrIhIfzikprcIgXF8vIhaCAPQ/jg8MEYLfNs5znVtALNnDQsHLATFUts
iDCKiL3MNofmrD4hDgMYpz5kPVdx3WaPy5CNXZZ21j0jP7Q9/BMajX8LKUpVZTyFWTI2mlZpWUWk
bU+mClKKp6HJdPgGNWwMX2caP8iO9JjP4ns4evXDPOe8Yejq8c9DfFMnLyC67cnxr//09rRvyfC5
0OzFv2KfxOJBwXabXpmN3WEFNzGImIJv9j61qJu0b7PIS7Fo5cNeLGcJng9BUq9LhmjPiXsNMjue
g3zEYj3dt2/iBZQkwk0tBdirQU8iLvBUhvLMyqmBpy93dyFgrzRM5rRe17rzM6pqCclgPZ9HNml/
6LLS77fzhzcoHXDHunmBa8+xcLa7U2E5DSyCVxUuOtuNU2S0n+56tACHaK6qnfx7HQhszYBpQN/7
VBVJqyZRe46WBIJQ7IrePeKCmAM4eLu7OlkHCr4F+ZIiyOuOxbimDBFHlYcdBYbylgjgUxEsuBJF
k99O9SughspJQnWTN75JRUNJOgpFGnOiKaQx5XivlQtz/SKHPxoFahT6QBCOVkWhF0xNr3aufFTj
kifYjb1PSRzUeeaMTeXmwuuW1JnQ7zaqWXmNdcyJr/iTBErryUWJBe1wBj4NXclE1EvyxOY6n0Br
v1nwfDpHsMViIf9U990QR4rb8rlPoYdshaWRIXZto/lxBWAXWMXM+nde+aepiwn6Ep5d6WkrzcnK
9pgVnn70eRNFIOtoH8aU5T+cm9DEg29KkMCAG2EWj5hKcNWxKZVjwUdvGinE0Edf8uOzPqvpOIc0
tdfG3i3bVE52ipDL7yI6oVsfOBMUI2kPdkgW2c/zCAyo6CNbJ+EDJvZsiW1swAXyLN1FM017zGkt
1IHzYD6JwXTOv5szQCv+a1spIljLI/72vR/coz4KAmEcn2oornRJ8ElLLfxfrYFnJldtuHKgs3fA
AObE9OCCnLaDekbygYLZMF1vZIsZ7/SNuDRa19WzZCKQ5dthzXUeCcFIrMtvBirAy6LHMn+yf8kG
XBA2tGLnGOrFLuKF1iXLzuAOK/YQeLY/zz2iBluvQsNx8/bH0W8t/F0+VX8vSG5UV4Elm7PmOBjU
qcOGP+CZRIFpGv7yrzoFF3K6S9U3NNhRP6kvunQw1HWSGXYYTYuOEiChSkATFmTSOK7BaSUACLAm
+7NGe1PkWHrB5j1CzNeQZfz7Y+FL255IpS55hP1xzyaYTe11tL23qwqptaFAvOaAGhaqbQCphQnl
TG8p9an1k9cFuomDDiKXwo0Yb1DrneXX+4zt16eURZqe7ttkVKPw32H1TG3JAPvY6ynuJ8S5ozaB
Dr6zSzMthouaJrzOjprSscuUUs6fU5cVnDXbCI/DBSOZAPKRdKnPK2SFP4NMHNBbvfTXc/QAkt1N
LF/BIcyXCPXxstm+Z2G/ab9ndZhS0c9TWjr5Duye296VRLNil758LzkoODqk8Rp/18AnwE/U0HRl
umHQjA4OCiAALpg96qLm9+WJKAClTAV1pzd14fhqDdHPvkbEVsF/mGIAMb3bKvj+65kLh2oqz4vd
0hlAMaNtodb9bSZG3PRWp8k89Jg4m28eGW/RZG73Oi10NDFKt26myAsD4lXu7192opqAWR3I0Sq7
Xap8ckb7cnli86os2nDcPH8ijTupUgTlp6+Y1ozgCYeY0gtX5lPQmTASZSA6eENSNt9wuXqgedOR
WryQ0TbBUb8rfMGwhzIhKG1jvLDsh+o0WAJ6kSK/bmCcTckX21HAACdut/ndBPtYqgUBcrp2WQkO
GvZIo6tVpcPi807FQF4VhI728AInZPAlsE5vYwGQcs8ZplJtnJcKRgm5qNNrSnKtPdMofC5fEjIg
E+RRMwa/DNuqBGz/eWQTe1GvVslXaX20HX2Kbp6hOTVgxW0pMtYDVIlyi8kwQqWtw4TiZ1Kx7JMl
MmXOZnz6qWbIjexHWc1CUY7dGMtJXhl8lO6aAYjUFIdeOnRcFR0OmfPvNH+L/j/2d4eryTdtFzPz
vlvAtFQfnQQY3b2cHxOoYZJnbatnxnCa6Ak2CghoF9+PbVPAeCbU1b5oEB9nT2RKEUShfIFokYmA
TOZGowwjLwNuNJ4wtGXRh10vWHr2ZsRzYEzcUTvbgBwyQPO2+wLH4sCFeFAziaVi00+GAItUoPBm
gpMkTQBgxi4AQPH7UU6qiOhuuBknLKPwfX5AEhIo8F5gODlqsIJWVG6n1jc+Qb6RTEIrCu54hBBV
UGmNdkKb/PZEr68MU99ftulQqB+RUxneDYNgGOGsKSrsO3A2BcfllbdAb90tERL0q2y5yAbHhomI
jDWISZ+dxcfTBjCMMochx5CrB9/phrVEkPDW4U/dCA0+n66COzK+mUPctdQubJuIANMBA3o7tPpx
vtNOkxu88VbjvMTg8+MqvagrNCn7Wk+fFMup8FM6+ca7LisPGCCZWxlD5xzGthAudvJH2ZSue+Se
LSp/S5Ak70HKC12IwswI5T8fFu3OkSC5JBIgsUz28RKldRC7YnJ+BRuGEO4Qm6cNGhnjkB66BeSw
RzPhrI8EEr0/x/2ktXk9U+wuTuUVrJ5F+oFBxpXwV4Zc7jg1vj7Y3YJtaaQ8F8FH7bIG4y0TMJ/Y
Cz+1H2m3cGcdAVAFodQ/HV9M+HokAEYaD126O+zkmtmDplrdDnZ6xJjzaeG47VEmdNVpSKsTxqCr
qD9yMTaPorrbQ/UeTPP3WHIq9PVHyf7kZ0v/RjRPRNLvoLuJCiB8GLmvFJhbRCTVWprXfxId2lYU
VRvvPxyCElh2ur2MsBduwMDU/K23uWTICb5/kZf0F1zMECj8ttOG2Ua86vht9rr1XHrS97sGXEbT
KVInKbc6+3AHCEUkMEZP8es+6nKyh5NLFy1iRNv7fmqFKgHwKryz53Tq+EIZaRxemPNRWGhTqqRp
YPcGhC03XX2V4yB4QADUwrQXIdLWP9NwDp/14A8yWS3evxqbOMiu5lW2X21Fl3cLbsiBD/Fy++Ys
gS8OejTbjddn0gQvKQ/y4FacPNvzmwYFQQr/B6yBNk3IhOXOcXIGMM0SgIeu1LC7r2Yb6skJAEMn
MI9oHUF5rVEACyKL5XAbYDsGpHOd9DSGF5TCs/p+bMkytxcDixjd5sc3+Y0yWKdvVaSSMcpFhCJ2
lvOHOWAselsU6NV88dzWTfdX7tWwRSONPo+ZSUh8Qz4+c10qY6ujaSt6HvgHzEg31H0JsDMV4fl8
0BaHXvBnAVbMpYqzuF3zLi55wL97A6cqRhWMD+/JWF/nxbHXA76DrfAJ5M4GWPKdxOysHdGUpr0f
Sojfl1GRtLG8J+zJvI9rZuk4DrbaOQ1VPxe9cvRqd7xDX3ZuERRUFBzRA8aVA0Vqn27ckd/5kl9v
TUdw5Mzc3Pm58y2QJ1wN3FMDo3hZW3RsGqqAIoIvt0EmnbC/Z9iDhLSV+OMj7jLrFuopLYnKcHTS
OdP8rFrA5CFex+W6RQyUEMTRisFIhQRBO4fzb5XyI17Et0GbHkNZH0rTeMSoK6MzBtBKothmyxFj
LfqKfQfudxRCQt11JOOBn0od8+3QcWN0VqokaYSt+3yqc3c/CjNSIyuAE7pShjCiBxlaN4pQ/pqa
jZT6Aj6uqsMNwaUIS+plLd0mI2SPde+uF5I4TguiP2h0UuStQZpyf6wPfX4ekskywi6NOGHv3XAK
fwckp+UtzDyc5fNACuPxxi/sVU2un4h9lXmMAZEK4BMwDm+yrHTN7ueUGlI2gh3rJDUQ93fsBQyY
VMYEyUdXQ8DZZg4XeT/w/97JM8WwHDFEWHqbdWtIzNtlc0RojQof8xz031dgfKkrpsBkEH9l4MDD
yrF3NA+9PRn3ALfxJHRg2hwK05V/mhC1f4HMnJZzgdAQvuxQuuH+ryFzbMTzrxMzh9On6X54ZBEE
zv8tofxLTnyMcqNhob7py/S68WeWXKp1jflCtIxc/YqLrszp6WQXGp+8Q5ZEo6v9LcSeQ6CSn590
kAK3EyF8MzI9tWntZfb7vQjPa9MS4TsefFwhzwhwcrZi7EkvtiER/+nN5I68SofrIxHOvdNDpgbC
xv+9PTXLyUv1OTzw8DEDtpUQsYoBLxm6JrZrS0IQ6fE8DVRcTkT9Lgvo32dOUW2/KmI6Yj1hWawi
vc/umao93X08htdalZmj7DyfYOitJxkpP1j7rEUsov8SlW4Y77t67Cj80ZpnrkVO1thAHjdAcVyP
xPGw3KasnpHMs6zFr/zqv2iUluFf7URLbh4jbbt/igbyEi5X2364dxx4fFdGNF3llJE5Y5qFQrNX
OuPwcd2ugZXwrf56nGbTwcEieBn3kbXtqvkY9Rpga581XnBKLOy9l5pqIjFVZYBpfwPMfhGBb0on
OhDAyL9gisuKGyeq1g9DDn8XhXNSX+BZ/Cp35jBuj4J1SHbB/gngSmsz0Ph5I37njtpSSqw8N0OW
lZNyNwEnPuJ7XzDY3YD4QWXHgJzEmkZPi8rKb7IcON3p1x7xrpzqdL2YNVfuLZfRq2Fd+8YeZrSi
ppllGw6OzZFVSptEdp8fv3pptfS5CIOB8cbrBK0XvLZhgw/vM1+DbKCJqnt0Utl6dOG63iXwRISx
zALdDA2Zx6mmOas3OqTpKW0Pie6sPmS96uT8TUWO4F3wPcvuopwvvqMuKyofN//sItvz2NEx2NKI
FKqXlD8XrD7dxbCX7lEsY8cbfHY+rUK+jLoSUaTHBVxwMLMhSEv14jPTxtE/RQEg4RUvBiYyX+Hx
z688mfZmpsFbzZqC8EwGXPYEgaHtYdIa4pqRz/UYz/Zw8iNNbGi0hi9HvuOOP6xT9fkyazHOUCg4
eBDHzxitgbXNsRqXS+hB7AZOPKMw82JeXi+NZXFTIHwpGMzOTtvg6ALiRPYJWBFn7D0dUD4qtwyD
iAJsi4DKTX1wlzBcrZ+UcyRYOknUKzVYSfRKydKyNnHiAfs1hKq5IIhP0AjGznm5NBXa7RYvrcVm
s566CCLcAB1Iq2Wh+aamHI1uYVsJkDgbL4zsT1eb36MjcRiZkmy43eSed7mc4+fkbf9SFI8b+gMX
N78x4nvWtRCQyCHROfpptUepMX7IOTf/Ksi8J4Uybe0tiG5kxmf/7LYeKW8GT45CZt8KUn7LyQiG
dLq5YbdAkUpaKiB6ADWiWd7fJxmtkR+oTJPvBqkvVaKt04Zb2rIE1i2yUvrNxeVqYd7n6nhd7nHF
aqnC7tcFkVVVUfjPMd/j7ncDknrH/Rp4eu9o0X3O4zItp+X6n8awMCR0Wx2hREdoW7xbhicOmydR
f7l6OfDwo1IeG1kXgGZbdtm6MbIqi0fWEA6N+9CGibaRNqDlC0krzyfZkVnYWLG5Rsp9mT7/blpD
22NR6gXpWSaZ9/Vg616l68q/Ee5CaiMd0kcw3lFlrY1I2uapDW8B/yyg74Qx9jNnNO1QFLOIocHt
R7pBiqBojqqGRN5dYkDNmZfUG6o0WCmsW4E5AgXb+OExlJ7YHU5wjx2KaTDUZiaqbS5ZBdIfHDVA
wKHnTizyLBBsFIZS2g/m8yOc7HYYobCVLqimm8RuGvKtB2uxgAY2zC5Cc5aEkOaWsCc+iOrahyYg
mgKyyR3asak5kxeL50fJeS5ylGPDIE1VryIK7g1qoX6t4nXQrd8QTE5TRAzTEwDel6iOuAmdXWMw
s+3rNKsV4FVc2sm6GXz/pxGZ6KAPdriKrfEUaLNJZWCMnwcMVtmLy1GbyTkBRlOovkL0e2nLdMTX
foHTweVUbZfKi/Vu8eMyqRBPCid6fkJXe+1l8EvaZa7TO4fVNjBfReR9lI7kBUvhabxcSjVDVDuX
9hjLYxJu55L7OSaQSdLmljjtRNycXff1I2cIIuUZkWzkNke0KRnpgIRJb/3GMCxip/0p2llnXBdi
JVFLk5o4qtccahMjEblv5CpadXXTlQmGAma5smDr/srZlVysvq9I52FrnmXoLzytMJdNsudN06ZR
8NFXkY4jXt7sA0Ytnwm/Rj37OcIjvyHZ0NRmdDZt9H9qnHf4v22rwKMIJAC1jXc8KhDU/W6CcikS
An5O6mRP+NBDFL2/2kALLQp8G91pAv9pewP/Vxt/8Rpkw3S7O149XpYv0N1rk8Bj0YTesXSKzoJJ
3SiFry9OoxBnI9qPniI0qfedWjJv7Z8sFJCD1eZIDikG8ZfTZkrgwbZeytxHun9aIol1yPyu+Vqh
tnkSTTcLJ8+X9zzVGTo53JjFq1nN2z2AUOIAW/VcsDv0Ktsw67dgRh2or3m9Kksr+35cZGe3DjNk
ZXFa6xZGB/3pjaWNAN7SnG4J3pGe2XJE0AeMhhK9ej8vvN29TmSroN+GJjhaM5EHjjiVNSPauLLb
4l41PPmxb5vvhhCVeM1+F3eEJNNdcqtfdPpsM389nIF3/J92+6YBdUiRlHg7bEH5yQPgQK0McoKq
4YVeFlIoEV+YJq+A7YsKMPqKOZA73JA5RUR3lbE7mi1V0aRriqKdv/9zSlwJIvBWImhpeMfX6R2E
Cn/zkhZXusRh7GennR8u18g7Du3IdpYDPIIBOG8PDyPqFAVcMYBzRmpdUkTupD9tVBcLGE1oymfT
iYslBN/WdjSb2a73yxDHvzuyq4UnG1mJxL7ae4suSkpvarteMEtAu4wGCvEMoAtD4ffsReUPs0Ad
VnIuJw8a4BI2rWPAlvv18A/tNypmT8gZQBXAC0GjkyJ5O52jyLk0M/0drxRD8XyvwA+HVJf81p1Z
BdjIkw3UN4UIXTVXgYVw+x0zX+ZUUtp/fNUO3MIs0PBOklvUDItjAPtpaQVK4kMB0fCRuiszgOj4
BJzNpix73nNrpT0oRM+H1RypzrwYYKPsHlMNVjt2rvetrqF2SKkO74N6KIZ36rDepTqMkZcrVVTV
ayue/KPoWYyVbym/uesk3Hh2EpS4aqgcpe5PzzIXUKUN6+FQNqzzm3QnKyDG1xVxsRpqNpi4Xy5W
wHBwMQk30oViXM1wIxUcGiU+mf5LFZC6HULC64gd3dGY7k9cb7tkDhKD7x8tgKTG6eo6m2v6gKcy
nzI4Zl1PrgaBCGefv8KylHic3jHd/mJ5v06p5ax8Iv9XnCthhdmS2ICkn9jQW5DYsW2PwgfKnsAP
T5qtkZoQUB50oT0jo4TgBT7d/KZFUb6qBM2qu8fT9ViQKkLtbppFnKOfh2rvzryLu6tWZx8+3qrO
wgd5X898iCU3U7q7CX2q/zQDlKjfZz4rSs/i5ilabRZhV3gB5GsxcUlRb4W+mjL4mNh4nXbywz51
nGK65+qUPW/ZPcFTQ0yErTmCetMvIvgJSU3hZ1x9EmQFwWQw0LPPMvqSupkkC7lxK3tCH0aK9uED
Vsx/kIQqjVgUJO3Ee/ITqwkR5Yip0jz72nyujmXzeVfqu5OLSbn6932gL4oWYuJs8rdo2SEsJo0o
rsj/OUcTnsM/TY5yAbx349FqeO64y9SGvEdobsO7JwK7f2pW4Y0UpX/cpPExFGseRQpbo2wADilV
wSWuI6AFfWfOZSG/jUXgK2ycQWy/7dBRWEuyAhjipaEr3/PYXYgr8BBq8iV19WLUm1/MJUghcHJG
reC+mKg1obD1dttRIgDdFccZuobJMnRLQRq2zPDLHT/tJ3TeZbF7YxbAUl0fpgj51v5k1UrzuBoG
5uoKcL+ZzJcgLqQbRvPJKHnEYIlXYAZv0bnkNll7pZPmR8pTxKtiaOFQBNNhW/7TonffwXE8TIQ1
eCH4Ml5fMMVoDc3Ewm2tKYlYeW4YmDSHQrI8bWzVY06icd6V3jzUm1AmTIG+WvbWbmN0d1BJmnQ1
NERuoh+upg3EZ9p2OQvIVPVdtUJilF63XvI8ysWPdu/oQygyRn6Y31EKvZnnqnEsmsz9vglvyp40
Un8En7X1r5Yx8DqcPxLLQOuqU1S0R/b5oPXiKvHp/YlNLTK7lqIbvrMglD4DiSaGCE6+ITXcLOGd
xRqydbNd1W2qdLPae0Dp6zsavmUGQI+2QGt9kANevOGoDoXcOCHeQidUwxrJuD7vstt11Wpn8CgD
DirskkwzxjfLuK9HUtMcoefKvG1dzhKplpi+vuanOKPcwt29RYX6M2CBhnox812f9LOggZhI3Pov
i9lqLILlZYDxMN5ZELocPiXsC1DVm6l0DUGFfjKm75vc/kXyLfdYWsjtI/36eAVckHt6yqWQPz3g
/Mxb4erGmJhaVW7N9vD0Vs8GrUjq6METnKDpfjRdHLdvXAs7UloR07sHW/M66VGnacV1cmojGrTe
ClhITdk1ZFcclG7vbSgppiAufw4vgfLEv+cb0ajb2C1jn9nRsjr/yefczqULJuYYbvKkW4s8iU/O
MbKpnMRPZup9bquuEl+Y+JS3qUoIHBaPN2i/W2N8UVmn0sZvapBeCsKJ1ehm26ypb8WJwj2/qC8a
nybDmKgHi1H02gWaFo4j//tCnzcjj5MnjkUk2St+k9w7h/SZdWk9vhNNCWVUPZV5Dg8cScjCtP7a
be915vmqoLrYOt1wtrDSHkcWHgdy3jKtBAYkWYUfNaay6Bz/VbHm1rWZ98Bj/Jv44GzpqCuXy7rc
4rXDScytcUPXeWFJOpxfsO4yUZqPbkW1dzN7VtbBWZcX7OYm8OYJSUthTD599+iHCWZOcclGaHOx
z6QxAajbdoimVAhd/JUL1fYOb7NThoyLeXtXh6gcns4xrZP/PKLStJcr5rs0QmTAX6f9X156uZuu
gsfo1WoioArUFtNzrawEBt8jGin0M/5FQnU1T7CvEbnnRY1uF9TgdLC3XhCuLcM4SceTGobxDnbI
m9Pqq4MeyuqTiECfFzjOOrEcxq3X1qA8aUie48megK0OxdV4e6fghdSMjQkAFW16xyhTv7tarDVK
DIf98fQnG9Z+O+trP3Ez/ink0F5tjqPgdq01y8dwsKRDifF5Mx0O1wuVLzhjTsK6ISJhWxwY5+Yi
xJfAWJela+LBH5LYaSvKDOAd68btBgPw68OEd2ytXmpw6AinXVJHVTjlNj+d3xLknoZDM33R0YHt
oSt0CaRC8dNUakMgWxqxMLinseMF1Gki48BRV9WibE4bYKb6BL4aFSzUNM9vdL6k0Jud/kumhflr
fWz2PmJtwL3sx2PoTc5uIjYGZ6GdRSlX5ei3T0d90gkzsSO8ZsqGKYB9KjFD9BVo6PqUqeZYyEyg
THLRca6H5sZXj6DYiHICbS9eZhGT2AAukapnXoQ33Jqv5elWxC5xxMXXKmqWzsyno7sN79PNBj3t
akhs6PcWtCs0vf+WXsJqVjoKbJXcq5OTKL+kqihToQ+h7iC1fasdr8e9crvTRJBbafkkSS2sTf9q
2OWLaXcj96bsxAMg+/5ockgSrkuv/MnWrrzhTgsvLjIeRZJU24kJb1VEv8sJBpiIbQuoUKNDnIFT
LmSXcMbly3jWzY4LmsMAZRpw55IW7D1UU84RQrkPMCj7hQQMRTwfajawHH3TTXoOQwMgcuT/zBxx
ZugjaGyC1imCNuAYYWdJLy7Vem0oJGaPPrpyhmFlrblnl71NfgupzcFyI9GNwG5Enr8pGSJ0Aq2T
W6bitMYTeBdciOIaBaASn813hF6kQk3Xq5qRbjuQSc3hFW2WQTHAsP15L4afZh1cvFdd+abuVMOC
DKiincH8UlLwOHgcIX7Lw0Hh3b+xLIFFceNg3Xv6Eps/cufaJxIlsBHIOTTarpbZJY3v74u2l63G
BdoCH2oUHLpY6rr/eQ3rrqz8Gl6G2Rfl5QIHQQa5w8x6JBL30US3Dk996bHybQ3/shfQloreJTCQ
s6EehTMGBsIcUHYb+QZaZYW8s/8grQS+wSAzI7o2ryDya6pbmXHzBRD1OpwbFEfEp44+H57sRfMd
/7NHDz0r11JSJdLu80vIQLhKyCC7M+FA5RxKhR2XsDeSQ2jtMbF/nIoVTQNKQsH/SPCO/gT+0zQk
Fp2yrsAqvT0ptzF78P0vGgUCDfE3hOPrK6jgYLII97UlHnoO/4rstjemzknIy1tybBkkCFI5kBTn
xDK6B0zJzKsNn22uexEz04lFQL5I6K3uD2NHcPiiGYc9gdkN0ycRGe1aAm2ndyi6GdjLcNrvwoB1
d8vDukxlvJ67hhxucXQ3xVrIsiM6h2OpY6ctR7Yb/G7o4ZxEJRYi/KOpfOTwB+3NzNdYv3nu4FEz
pX18nIu/Ia0HD3WfhHajvycwCbTeTIE7d5C+mmLYGEwQE626YXK/afva9UfQueWuTKxnJbtYYGvg
TaDnYBOhbXCgXn5+KvqcHZ25k4aMBlcNk4e5fYhBkJBkOAauR88ZTDLtpBdR0Izk73IJErdw1E3X
WfY87krjloTw1c5OQAeWiJ6k0/Piizdyxzk7W57gdvgk5+fatSqon+xcdhoKA7rLiO9xwXm49Cvz
b6r+TCbedcpjpKbPXa8oz9J6m9WbbSVfoX3oZV48LMFPKc0ut4S5+goiEgo/qcHY8QI3jdMCId4p
HO92u4vZGdDfrUcKmJUZNfXudSDapRoWCrlwUfgiwHKsbxryCAyT4Vz8vOwaLFmWUe4AJHNLwc/i
mBfkrATEbfmQg/meU8lCWPJmbL+3PhTSFrSRjjaY7cbyy5sBnhfxn18agW/2lofUi2V6Xn6XQDi8
iko41ie2814d1jl6Z0heti7ltsTsTAxPE48u/2m3MDNRGmIazQvqvfmVwA8pmGN/obg+Bu0rCPRw
drE97bE4svrNuIWH9MW1/BzD0ztYXZGkSPKlm3wjBzarW8krdDu9x+0/vCwk0IvfIm1dcLnP2pK9
kyfEksXs2ZA3lF1DQXybBcSORs7FFsKebnC0nn8+nJeqtqoyCC5gkcA7PCXSfxfLKRYvuzjRzgxG
y0p5ZA6HGxgtvNxlSidITvkczani7y3llzi2Wf8vo0+h0lBu3p6S+Bwn0q86IkVtz2GIPdeu64To
hIQI2viEK/AIOxaqgdwpt8jKn87UmewR5bhnCRfhG0oXuUl17OInHOffnjhLNmlclVBzWpD+9W90
v6cDCqAhfh2x4w3IiHrqSNCFCZa3ZgcgR5h9GFltjxSPTngAhv2dA0MQqfgv2zfiEb/RBF35aD7t
Byc5AUedsc7dK4zUGBMjotQLf2uHHeyWIymFerHV/X234fPxKJFauTqrvrX0RKIIs73wmpJ4Kt6k
HHxIooADQNG5vmbBgaGTZlIGXB+pLBkyiHNev/ucWqzpONpG0XRDZNCoLS/BawWruj3AVQ7C1b6I
EG3sF98MSaSZCdYQIcDN01lHQiMQUPxXffSrYbZlomLFs+1VQDKdsT01trFJnplzYArXE37iwtAA
pyDuvWzDatONeF7GGoJVSPCFp+i9Du1G+CLxqy/tiYORZ9PyVmu2AGzZKw7DhBayn5+MLfNlu8de
LqIpGSlo8VRXc3MGubHPvX0ePvjFb62zJJJLYK2kT/h96JvubRXYu3Hfx6zAaX2SpBEWEMpWuNaS
luu+7bEu5TMbOQeFlricFUtlkhsh61DcE0OgL/zsZfb3QHaszDm16rHqvHJaQlzv7/0MfFWD77El
INly2W7j7wp5CoevYxuYVMZWtstXK72YMyVqrLzg8tdTjZYqwrIqwwZp3yb+BfpQ4lrni/YMPJnn
5O0SkxgrbNAsGgIWKzwd3EbK3jpKbcJhDQrs6LS44SQ3+43xvxRDDACtcr2tX+55zV5H7U6vUXG5
efygjhWxf50SGwjscmJrcIPfuZrWsgd7eQxqK0af/ipbs7mDQ8nJ+btotgufvLI+7jBSen5pxo5X
uEAU36ZKTEWra753d3WNLAF/MaYNmw4skiinuDIp9WGz4rKzwG/A+YyVsMx9JIMnmKlEytEdpafe
/Pao5um5V1lzBMTQnob+ku5ZQnq5+PBvFE2M83WFoCpu/ttH+rUEIuT5/gpvztwbWrGN5kPcvhod
ZSih4ve/ZAJl+ijHrz0kDg8HY8VYrjAGR6VsLN7S21T4ktsG9jO26E3Wh9JeK3eppa1R0rx+urSU
wqMbvC0+KdUoovOTlplSXcbUn+PhskB2aqxhe2i548Ov0+phqJWgXS2A1FJT5yS8hfMUVeZdGfvF
BVGncg1LgfjeLHFKATPSKg+6LX83b5RCEvKyiIftpJ6tBjmUXJBS58kFIGl43BtDDUO+GKM9PXzA
29/6KCKpnb7Oe9Qb2Jzcp+GPfdkHm1aRhiPKA2uuowWkYGY8lZnjlJm2cLEDyH1ZbGobmvSp0t4I
EGZhEzhV8gyCzBduUHGJjCX3HyuzAlGw4Y4yX3kmJBUf++aqbSycSRFn/YLz/AYvuOJpXY0xEs2g
kaPOvLa05djSk58c1M/AQ6ry+KMOyJU6zS0m+qOyCxb9mJdMBTNq/C7ZGqssoXSh3SqcDTCSyHkV
wh9ZpjVsv+bb1IWjXiIZ9wLBS3F3MNHxhqeXNdkeLFpkc+RlbzjBROtJplRpHm8vrKYpJGODzfuX
TYMkVTyjtxhz4WqNnIqh+pAe8ILPgeXctszegv3uXmS3vcZC5VXT5nBlwIrWRTpE+ralicA3mxmn
Jnt6dHokliIiCBqEaqi5cJCIOfguF38ZvyFCdIW/1Db9z25oHXitcUcISeOSwDCkyt7kEGa67ouy
XzT3HKuFZBXWgC/IToLVFNaBXlGD23urrBNf2/aYKmtnevfmXIg2zsSGOYcyVRHDNzUpcJmotiWw
mW1xyn+O2NnBtEJvuUjA6yNGxFsJDd1MQjEw0hFa+C5PTsnKOw0NbhpsSZrTaBXt0ffPdF9VFrJk
Xl6ppTrd0aGfzchoxI8sZPtYLG6fMBEkCCrK3hvHVAiFIKh2Fj/SQJel0JHPGNclQn4E2LYUB55j
tcST9D7Zh7ojxvw8gLrAi6Qw+B2+CwiK+H+L3VkpXsr3l55VDNTCmqaOaePUskGhjY1bJdWQND6c
uDGQ4z8k1D5zu/6hZF0cnUwHOiWo0UCPGS1ZQC2rFB8uthd0bd1SaO4vTcSYJb9XcYYz5POwA1dT
/WiaOQ/7q3llfuCF7NTByCny9zBrbFNzWF8rDRS37gaFAmFUt1ACY1CNX4JhS4xOVLiO/IyD0YJD
OlbNAJhCdbMAu3RgulEjdD/8pebVHPrU0J+HFIE8bRoqUygR1Ktto1gm2WDP7VXXY/MALiHTsP0w
u1Ufzn5HPr18CTf8sGOBFKZZHmCynQRcMe8jtUO+dvTamQ3hi/4hMMFd4JKaBl8w71ewnvW/BJm2
tqN5hOxuvmIkw5tZ4MMKqAM3KYQr2NjPSiIJ8FdMkDgNPN+7Ywb+Lm96kjpixF2SCP2Km6y+zK6K
sKirgV39yS1FL8V/61LL0jKrnBdD9GUM+1gWbJMfCZ02BpWlNTH79O93rwaZBgKJ3LxfVGQChztZ
kKu9h1U0qeysvWWXSsSAPkAtyfNC3rLJ6X7Auu6TNiBnpSMzxylHEHiQB5rBKlzmZFapzqRRESPn
n705fqK5TBheWoaYQ9TtGzHijO04P8g17MH3cgKegKZ7ATR5dVsjfLP+AgiXHNE3qZZJ84oGmH6U
ctvVafNF/V5N+Agn0LrJsmauIQM2xyx1KyNGHGqss9vwm6giiLs2YO0rj13pS2v8mZFU0q2b/hhB
9XjwFrm0ypAQkP94418uH0y/ViBHO6yiR9OsVAHrN1hPwEG2wUnEFOXjdu4rsQr+tm0UvTmcx2ot
TuT6m7hAJ/Rvwz0b23G3m4fSlvzodT9W9FGb78AQ6FdL4fYpXsWkXET0EBHuhQrDNaVkEZp3eeJs
i9+MRvo3k2N/dSXaMyXu3ee9JcMGWf/KuM12lNW9izsP5hjD6H4LcngTN20r5IL/l6I6m0NGEiR8
0hqFAnTfo0Pq5vtt7A3xKTeHLIFRLO7rHlK9x+gNqUdToRWrEDe5e3JpZ0BmTannpL5Pl/E++7Jn
4DW4Te1IXQgr1xECDhJudLApTLx/C0HhzGf7ifs8PQsa+pnkd+W9jSw0cYY1MEPPOHYPZURW7cli
z0j/UQ2IIZvx+Sbq6w8UU5pzS24ykYBT2uPI08Epl3td1YHpO6hOlOy5QptZBh5pIKJLfjYDltxY
J/LX2m4dIz77a/Fsy8oSTx1W2aKkSBRrpUhQ8WSl5R4Mofws2ypn7YObeMoM9UETNaLgDOPu+usx
l6eqr6desCBKuF7r5alibR7s5PqYNCkvgSyZIuya/IzMqDoLlgSDfhJb5VTycrMLDqqkpvRdmHiU
bvX2+4vCdylBRlNPL2X/tdvDOpfd/C5qvJNQmFweTFqA0xoGVYUNHvfc+3CX3JBtO06onvsZXj1X
KDq3GR+dtu9/WSjuZaxQRywZNd2LFHnvqrHroJm12kTg608gHP6HrKkZxL/0I4cw/ueRaAHpLDy3
moDidPVSjrRkiU44qWkqhERj+EeRzrVrR6N4hadS+/wjHMQ1dV2J6noLlhdLYprIIbunzAaxb4vx
+AT529Uea4prJWLMM/n0MsfJp2XK041IK5mHkNfbqsOregA3rwXyNfz2gadaBlrJHLEl1RV+k1G3
qHXCqQDwQtoag02VEpsY+eDMEzWELCzSj8y5QWSC9krv0R9DqZKdes4sf9dZEtLU9AKZ0qCDB2PY
JK3Auhwfrewu6qXUtfFwwZyJjshqCcvqN8chg3FGx7yAa3YoGfj32c77WmTKTPE3c9QpmFARRAQV
sGYyyjhiCw3jOL7iibCot3aoeWGNaXuIrURrjd7VPhFRGoIfjhn0WnqaDpnBagDGYXiZ0NZ0TEPA
55pcaCpGEkMbP0eu7la4DnNslrqTuiQx8FoE+/WiK6p7WG+f9LHeIuJg3zAW5TEEIhQIR71bNNKE
X/M5hyX5Utni1iROOx2jFFCTvTCMffxrFRuYQcs48LDe5BzeCT9whUB7ow1wItHDj5IF7fW9/fAK
IZGdizvigkQi/QNa+kHLaK+Pn513gp4wa4+gGORoVsdJk82BpQuctpOS4SNcOWQ18wFZSKuzKP47
04oIg5+QJvfEX1AOBdwHvuofwfk/9mRsx5q4LYN50MGtzinFgc4b8+J6D6VNUUpyuoXGbtupY7Db
ro/SVGJVvScs9xIspBywid12S0n1iJkpf7e7uMZI3Uekyd1WUUH/157pB3PAHzedS8qLZDOX0Z7L
d417TSmykU1r/MLMYOG3Cax3ZtmPqPL7n1SR/GSwQ5FyBQIYrAwzJgzw6TqAu05Yif5/v47chSR4
SZ81rZ3KmVGcy2hKPoQ3OWBgLJAvGbwO9Zbv5x0OQxOlklbIYHEdMv228YjTA2YUMWkWlaGWBkO0
DRr/i7TLNMbejWl5iBcT5CO3hRNmJRSH3/6LBrtoqLMibigicNPUD6L/nL762nUCf9mKhfb9ttW+
DJKVJo+0jMELrC/rQFyBwpNMPmJPkQ+joXiLXDokmhXVVe1ojV2+lD5QBwjUxylqj1LhzhOZ9Qdq
ASubNUQgE3rAFeAc4T78rL2iH3RWoTxBIoAkxPfKFHnJ2XBeuCL3A9tVNeW+4dusNZDONqdp3eyU
FFRuBKtg1hBCUaM4zdeSmBXJEvh+xU+jbHYKsyYDXbRTWvMmdhRSb0Ya1MOPVrojB6ndezNM6GaR
k2KMKoy68wzyGcGKGff88krbBj4NFbxaBXxRwD8/rdyhGtKuwth4wzPUBBzZTuG4KzpQoNFjHT6y
Gp9PG6WU2xUt2HvDww5HaKMsUc7hvS81n2IrTfG1vZtaPqLicLQmju6FGenilfFvjFPiV3G5lC6X
BgJ7yLyXb9fCKoh12ZV+lD/p/Y1chfnpnP1aTZEvpqG8HOb8Pm1XIl53SbOr4YYRbEBct6bYkNTC
P81cMhfpUCZNj4XPM1xjB9hkQU/q8ennUfXWYZeLLjA1szHwqAVEYT7i/XOm6feZIlew2ktjcckB
pAXiAp/X2FcL5JqNFripZGqyDFkp0Tn3jjyysQa6aAUYqOvCugh0PzXTJe8ynpKM+P89Py94kFle
j0jD52/zCB+YkIcTdFHgH/S4pLDT2bdDsDwCcGss7+POGo5cGRciva2Hu+nXPj+EwjNrAaUFKqHv
Ap4c1j5YgCMKNBD2FxoZt4GJfHf9nkkAg5Cf5JHAYKG5l51rRQfd8zrXRPYDWoQ9VO3UbEWFZ3sv
1uMdAUyCfb4yRvjnUfOxfYD56Urn0X/5SwHiUOG4WcK8Qhz91HC1irPkzt2XK1jIEfn9d7EvYSXO
UjbiNj3OjBwXEs15gZQSELD+bapDtPOutVBMsxYDjq8UvgEPcXStlpacUEbjGrLehWytNwly8o0I
ph1iAbavOWvlr7dnsL8ro1foixBYbcIjpuOUnnv8M9OLXrpNCO9iQUTq1Q+i2Oh7HjPT/OnmMsUO
EDeytmhNRX08i9eWUMLlTKEdk/fzrU1xTExnJ0Yfcw359j57SI4/r2u9htIHiZyCzeqerq3sRmfq
YsUdgC7hV6wB8kWuqIevd+n5Drd2PZsxeKqWqN8VUv36kdg4cQBGG4ZLppKOn+HZVoSI/a+ehYeq
YU6h++XTvK7Wvf/h/GcE/1O7QB27llwdoGXNS+t2FvExdHNXUXcTygVb09vq7lqfk93JEk7Of6qh
XWgoPoGNLjFU3gYQYhkBGwjqxwlWlsDsRFTcaNY8lYmEpfLzgMtFjtNHbH7inecRGyEgpbUBKlj2
G05kPWEDjkUQftZZMD3kZytl6Ju1BAhezoqQYHdpuwlzO28CH7IHOa9jZZIaDMcWXEtu8d145o+m
zjF5Sa5PXkRbatsxftm69JXMqXz1ISjE1NRuBk/jOmAUXyXtoH50gkwaxaOZ31p/+Kth6lRG+RBF
81/6fM81hxfZfuUwfc8PFQFoGZI9ZndwuD/WaZ3mjOmmQnHCwb19HQeOArvl9/J3HYK8ILBCt3Wb
IRL8Yj7N+DnElCZUpgWWiVcyio8KCXRKpyAUHffqg22ar1X6B9h7U3kb/R583pueo/AYkS/8jNBL
CnXFnRvf1lYe1ejCeOPDKu86VfvMjxmCF1LjLONymUyRssFIK3w8RgtlBdZrH5czHhq3FwwqlnxV
Ak2xYlRWgEoOPZ59M/vBFzlYHXJlkczt+JqEsWhRw5r9KmbckfQJKiIVfE94zRvV3bJUx1LyuMTz
UukFMc0CUSm72ObgxAqh9AXveIl9gHftVJ1zdnh4YRmO1ASAlL4q3oGFLWPDDC+Dr40PgVaF49S0
k2nzoFcYDjKq+WPn/9jMNeFW0RPYxbSV76PxMEl5YYwa1enz2FSZOJkAntRz2UvXZFh22gWfz6H9
MjLG4Uv3YD+JuprmhAwQXIDKVF8qJM45NHnnwNS3MMnC1u2to/UHUEzY6apzrAYyuAO4ueVh9JzJ
hBA/zEQ3RDOjoAE+svmtujt0YVb5Tn792PPtTt2ub/RQ3NqPvyeyfp+WgP3SVTukxdjfoSst+JXf
miwSEOZha2UCM977+jXyh0pPktm6KO+zuV9YpF+ByZ5UCZlqf8e/7mXSUw+/N9WlGuDZRgCXbsNg
R+yKMajVKww81gJaj4DTB/6lwByvTCErBAanY659UN9EnhHLpzwNmW0xdnnr3otsGZqQ+52rOM/M
dZNFdgYdz+/Q70wTc3e3IQKnht153IcAqlGnMcZS47NksLLW34f4CaKRYuJBoB3EZ2ixLKEhG6pk
EyQf3DbiAXLsiEWE83vgLsedOBVFclfkU1E5CJ/OxHaP79rf6clgM01DRVN7vfhrYA73SMEdKVaf
FSS+ixpGnyAJ5OgsEViyv3P9zqg9RVY0WNKk0bXG7UbbySqx1Ic5Rr2LhKWcQ8wPPODDoLGpxEWi
OfwqYaMXX6465ZW2uGSa1+owhln4HRqdRS0WrT0OaxGBEie8GOfuPSsGonpCEjPss6ZofkPIBjMm
dD90WLL02uKvMToIKmfrmT3F5NMoT9vH0aAngknRL4H5tc0EaUI6cIRNjb5aVXg10vzlkeYzJwJj
9zFRfpW6k/Mz/VOVbrQo3EJ/cA3rEl+G3lkP0jYDgJb4OSyQ3ADt4mJ7DJ2hVVSYfaqvdLayTGlo
tG8qj7n/7G0xNwQ0vGclhfv6oujn4Mq95vqcngky5RmOuf669FJMaDDbKU9Bhg0PL9WbgL02thmF
F6D0pW1OjajQRxSCSFnZH4W8qvNQnnyDnkI6E0DXoYNtevZJIqr94S1lZ1euXaO6n312C4i8G2/Z
WusXOMIDf7my9KGpItK/dKShpYMZCf/VjWMzT+JrwyD6mouJT8Uh3JX1NrXp3OMHdihkn3AKe32h
hq2rNpwe0hDxdLkMa7r7B8Ni7Wb4HuWAcK3UZ/acyh2UtNTN0CKU4zdCUN59XzHdeGLbZXG9W6J0
56JwJYGgX1W7bowA35/C/qt6U6zm6lvP4sVcJXyaJ3P5ITu+hZyj80LiRdJYrKy1LBzzThTshAaT
+mRpGyfVQ0+KHBRjWIAENK769K2uEhGjloH29QV81KapVyQbi4tPwEuZbYyc1vUNOskRvYqq6qb6
xl131gn5ENVHcPzQWCA7sJppBQIZsSyVG6BwWWKDIJ65DChuijHfpTYS74hnLTRuLbEBsoMP1iNm
A831AN7EvKKLKiwx8vYfFbseU0ObDa0LtP+ySlQiOTMbiL+JdhHWV7xoeARaAFuwxaMfgvO2LAXi
kNdN82FkTBT8CWhavzPgypqkNjypPT+vXkYvcokqdy6mAftpEiYGSUyDtLPqMfVpkCKY9vECsWOs
Knhtf11aK5aFxWZo6xV3b3sr+/PSVyC/c+sDAGH3j7rvo/1Q8OV7UTIfEMx98jG/Xotj7qZ0oohp
7vB7VzvNco1GDsD4rP/BDUEBsxiyc7TE1WLB722676H/IqUuaDudwRYM8c7equ/RMvq0JSZGzZdj
sF/p0EFMxfHykulCOyYyIHcRH0gHm08WEjrZu1JbjH/VUCtx7LQcVovqXmHm2qM/Ah1GvgPJ0RHu
JeVy5U7UibAiXRBcnl+SH1k4tUjjnPvLhGtd/dGSYpc/pDeMpS7ahlvK+42tzqQbettjAVhygK6P
uH0a9z00oTjDsdCA70XVyet/Ne4lBqjILpeOt1O7OqRsI+Kr6gD0sYktMo13Ga9XaaygQn+gZ60P
WPkDOqfLfS6PCzjaRRmbTSf09ti3/zPYVCVyGnw5nbbCReyDf+ckcZIIA0RZlDoogFuuDcMdCWDl
+y8JbKzup2meMY0TQWtjuSTry3pwQSvHaFZTsNg8RSqRtvsJIXTjXOPVosstRbnu7QhW2KSaavpj
5kxSQC7sHkAm0TJWwkloB8Mjs4iQ8khtLWfS11YWBoLSSnC24ELVGv/QILhUCWZ0AowQ2QvYBRsI
csUj9y1BJhli3wRHxzWDiHyNTWSDc1HmBiwUKB8a0WYsf8s2P9ip2tZaUuCwBex915tMs5kYVJQG
lENiaqlwuwHV7YlcywHmZPzsQaahcRJf+dFHRVzJAXev3igbJrnII9UVymy1EDqWm7e9A8a9blX2
sWx5uaDa7HUGA2m4Es+2znlBSQDBKvj7uDQyNQfS52AKv9znVv5NMrZRzrv3E3hoTIx5VPCh0LOo
42FDpZYuziUdDanSLccDT333dpyKxYY2dfIfieawP8icX6NhfKecIbr9L3mf0F6jMEYP81DI3z20
Yp2RPYcje3kuWXt8vysh62xqXQRGn7KuubxKVGzYwm143Z/NA8DZddix1ohPMaDJHeBS7w7FQ2AX
Esb+4LW35uBDnseVFMr7yfeWjkngYH7K2VjSEa+SXTsE+G6YCMh4G7Pg9vS6QeXHZ52/tpvFj6bn
MRrpdsB4XxlVGWYV6A++kg5L9a/PmIg8cAVBW/a6rnXHpkwJkkIjNVmIebVKCzWNlGcDPwGWX/N9
xMhETAJlUwFnvyVqu4E+IcTfxNZDssedsHj/y1/xFpeaXnlTVKb/cpfPq6aRhFgRRWtdJuad6ke0
HLIsHlGVYAr7Otriv+zFpiHnpdJRsVuN6GCz40Q0pGJic5A6DjufhNpUSQDoMHIejZ37XkDiqETg
Ip5UL6OKeoBBsUf2HDmUwIQ2tmi3QkpdIcU1RUqkYjXrAzOskweXb3NMM9gFC6Bx0APffFy4wetr
CEqkK5S1e26Uq6GjAHoiirdBeZkIchmAXbikSVSpr/3ubInLETwCzxhR8/Bz2mSoSE12T6nn/OE9
1HAulXQSAve1r8uVdnsCA7NS1VxGGuiT27hpwSg8oNSmDUvzsiCYnzlfLt++4WtF9ewyC8TwMuvP
yGzOp+cZx2OzuwwXf5yzIbmyWbfYkdMJFFJeixmmZCXwNpUl0p4Ie/DmZCL/IRTZeGSzhuZuK5Ve
QjGGYwjXs3AAw122NmLCIKsBKOPAaj7fzCC0bG4ZJYeiiV364PS6ZKAYNVbe4KnxvT7mZ826cGxO
+ZcLShriPaXpxC2nbZ8v7+6YITJgNkmCswjnWpFL8fd5JfSc1JHoHZmeDxdZQYirvQUZARUXSia4
vDWVgDf6nQf8CY/MPjYBcm97XuO86TtqD5qU2rcPieHsQ/k6lkjPMtbuZjK2Pp4qC5KyS+RnLtBj
2kgCmhfMKcbyOmOlJTMr+EBeTrFvrDu5FnwdjPokTe8U42rpfQb/9SIXw/ScJgwHmYZtvEHXKiDi
qwaePG4LNlXrqzXPN8RZhnt2F9TQBUAm2W0pBLF9hX05zdl8bhHQB30gtfkMOS1ph+I/r3Y3pYO/
nKnkwgb2k1uvPHsAZYTxbp02lP8ngoPbMUSiYPKMDbz7ssN0ZkfAz5u4HqtsIyKOVkG9ayg9L/am
2Oogr8yIrrGWpJE6GubhlgxXCZ2hYyojVZs0BYICXaM7scbtrLFjJ0mMYpYRrauF4a5eZ1mVQjaN
1Y5Q9RhlnPBMOlzBgpzDAbAeJGA70iRL/61AsFBMeHWaA3hYLKelnWREtBk2vJ1FgMvbkdkHcjyr
Qf3dkRicwrJyfH64fqdA+QkD/BfZ2c3Mj6T7dP8U4PJPT8qAx60dF/1SOp5cnyp3KnhOvIWG/Ah9
FL7v07WNuDxIfY6tYA2I/BbjeX8enShl63RSD9F9Ncn5U1oZVRJ9PUHZuPJkKWfbUUL1Tt2oXqm5
Ny3yJXnceS9XFTvVhIAhSsz8+mc9bToCev2yafA56lxvfFHGIFjIdPfVgZX3IH1DhZQmsTc2KtbS
T8HDDxDLv1yyLObgWxV3W/4VIUUfrXionGgcGcTS/uqUtP/Q17xF/0cPCRDs24P+q0e+13D7rznC
rK1MI7Qa5qeZEU7z/tyWvG9xXD8jK0er9qeoOIvtXTSsr+mPjcuKLSDCK2ZhreTldbX7v0P2t8lr
OGmAVuOrsQw9UQDtnHrodW1nj34JrrfvXt7zqk6E/Al/6VGmybEuZRCNlgE0Z1lhkmZCNmCTip47
MtmEsZpXpeYem7prxknQd+mgLvq/Y4w/eVJpLSjJBbm3vfhLsin6eUDvjnqCR1wqcSSaLZ46UnhY
1LWzjRX9zWgqElRacnOwKPsZUoSmW8F6aWhGYL6uwYKjoorHA74faRCCJKIPigGIXD6IOOU0zQVp
WOySajwQTQLSiSYHy/0Czcj3k8dPhE/8Sf61CaIaTdzLynHirhuDws+m3jCPx9qBoYRG+DR2jINz
OXx9RBqskHUeHy0Sx0pD4CT7hnO3YlEjj2i8GyOCr/DlxAz/qCVCIh7w+xuk3TJygD1wqW28OWS3
WeGaCikflvUcIQ51Vtho+qKWVYl5BbnehuN8uNupmC+zKcCbO28Kr1TXZ1Kp2HvsCZeOnmvRDSEe
1NxlxLYcnThnANbNVIQgj9rmM06zo7CrmXjp6fDCKqrHIid15c32/KFebwzvYbwn+4CkZhmKkria
XNuAPG7rtRjyzSWY5xwG4wvX6dJNapdm3bA2LUeXGlWxXnMTPy36Efgoj3bDO7pCkl/Zn+4LWm3+
2aK55HGyG4KMR9Em+Z0lQA6HwIUMHNIcsomDLrQBFF0BTL654jvYp+QE8vDDprFCkEdolByfrrKo
uCgI9Yq6zto9IitUSiaq4GN30pmOAF+v4C3JFvVIbWto/aT2hbXHAWe0bUYiInY2qccH8uSsX77u
coDhjXZRinvHZzLwbhYNFt3k45C44f1y7TPAs73wE9LD6ZEj7R/sbwNtB0CKLshua6YsA2PlProw
/hYFTuVaUo2wpoTlC6yiOTfNfUxhQj8qzpIus4MCX/ujQPGjYFASubzszrWHavp/CLkV1DrcoicI
VOdwQynpMNRHI6QKSW4e6H/+CC+2q4WoBwqGe0ayEuRqbCVd0zpFQHcvgLxgMduiv5zRqI9cR0UQ
owDjRsc9x9vs636cAKupy37UosmjNyHj0WtqXQCsoIoCs3mA4bsE3oQt9usXBYlnJZQLHVqHLce9
pNrpbDZAdATOsN3vZIMdmjdRDLJcVN3D3/8bGq3TCGcaZSDs2a65LekFZ589owJZXiAe7BGXqW3N
u7npS45kJHeTAmFETL5IGEdQMAv52FmWxYom75I2iEHqU+jmst253hKIfbqfED2modkgbv3g1s0O
sGtfMf4Z6FdGX3rnK0ySBUJ3CFe1rArRAx9aEpQk9+9Z7p6TURMl+A21POhuLO9HJIP4PW203GrE
1jRZAFHuU4tzWp5UAOx4dWX2V69OJoPaSZnoRjLKuUySAmRwLZ5AmP6wKLGPap03kZDuiq0RhWgR
uiIv1+1tZ4OTHjTMVnLEpnGHe3NW7/5iGF1qRK6BXbL41W1Th0n01VOK8cfq0zxPpFne4Acvw8lY
yZI8mbSfDmIy3wVrJkIIpQJSo+TJwvIZyOXQqtgQQTfRLOGCf0MglxajBFwpex9N286xjqDh0hlX
XpSfAz1XthTkE+BG2yl8vgXiTzIwasvBCjN5YzMco7Wvtvei/lC20CMPl0111NRGC1QIM6zFv8E8
dC5qc4omEb88jY68+dXZmn0URcr5CeRMo/TvHye50PfsRykmTY8BWCfn7ETBfirBHNMJj0xNjsug
1FXA23ln3mVaDhRXh11k60tUBuBrvoBVsNRIQ7+vehPnFPiDGjRCJ+BEjjkahtQcUC0VEhrAZkuE
BdANsKEXARWxCjgFJknlAErJoQBd+odcj+Nyqtdu6t7/zBkbncgHYTpr1TD4z3mDi2r8niM/fIye
lIH2n3HsNKAAK2D8i3IxTGujWEgCWEZLQzH6ASDjd7PYJluo42SDbHRVd0BlWvfI+Mkppu/+fJ9M
PPLI9OulRcrbV/kBCmVwnn5wNEvMCesMgtS8RfjtG30fDShkELf9PGKY07mmsbv+wiP+W8PtEMba
Kzp96qITXPRLjkn942vGAAtKXpa0CUNSDIzinnWxDDE0Cvc6XIlW9NHwNE2K+lt7QQU6qOuFPg8h
P76yztk4dHthjZsTgYV1HRJOGaWlL/VRJqZNlXk+HPacHHi237I7SnHB4tbquc/3gEC/A42GnXTQ
S/6oR5ZHZ99JTfEI840fwzswVsQJI/L7ICZ7cnAOQGZaQe7wOOKaUjzUMlR71TObMgF1uY1nH6xs
geWufJMXi6y/lN4DVz6mQdTs1Km/7WHO4aRYiyO75DicJYqTSszHOgnlSXMFz+G5+2vLsso6WBgr
HxrBIGNCa39LMgrhdl+ikmLuxDyficg0+3qw2FfIXEKqo11uuyh0tfJtKaxZmkSQUjDqBhikvuXn
XX1+KmOZKxZQesASL0pDmf8sN85u5yaSodJkzgtBaDcThdWsr3iARW4x/MpCnVLlVNw7YREuxVwt
V+FjXwpbQInCvE6ebMLrOBWzpibZ/+rtiQlSKtbyZjm4msun+3D1FR9ptUkVtBUt9tIFBIW3OvoD
WSSHt+vjvtkPqFxEgUD53Fhb6wEQypcsNQXsWuRUXHz8QNDnBwk6qf+aP0jTPuo74SMP+/PavN/s
iqkONQ8TJb++3lkhDyVWRN7Xk5T7C3GHFzrlu6BvAlExonnGFBv8ncNoyeKlEG6gMvvnnYtW/Dhz
OqMxTshUd2tMK0OT3U/lwrrTiODNduKFZov4ZoJdcngAy1/baSq915z483lZqlXEuxz+yzozSk+M
JcwXwwpTsNESh0qcQ/QmVmxf3c6YWiTvhVfzGqEVJdGVnZ0mP7cKyyuzMT8AM//y08zaNMo8wstB
uNn+Xsq05Q2aUQi6aYbCfp2dTMzgbUFrfvUTY5Bfmv58JA4fEulbanHg7Iv0FOlWZI/LvVPA1XvB
eWe1WqMcOoiam6epeUn7Ks+tfABVpoA2bW+0Qqvk4smj/maXYG7NZBMvvi4bzNNL7dAY082yboli
sbpZJrTMQJinZh2r6SMNf2Hph7xcTX8aJehx+JgrbStvKevGs8LyCsJeHjjOTHqXWwN2TfxkI4J+
on9oNXVevMFXUgbFSH6Gya5fslJvGHKiErYANEauRc+Q1aA9VdFfYjDtVexeGAfHNrGbSPR2LgCN
I1UM8Cv7/rUFMAcpzxgOkLJ1nZLdjc4t5+YCxt2nlV2gHK8eMYxa/x7mmBekKFkFtN5U89EZdTUL
NXxcs/nVwwI33u17wvyjY7gyM61y3hnqfvJjSotRtOWP3MTxGQTgDHTqarpIcNugtsqpmRVM9mIz
86DJvSa5nyfO/gLhnEct1A5Q9ruy4RYn9BNh/XFRbTFSVVGd5sC6Uq+nxnVc4UzHya8kPnPQ2RGR
Cd6/VMXoMMOAG7y/4nytZ4P+1YbLcNuZCLK94RllAB13C6VUswZiKWVlgAnx+cO7RXTmqF3eJ4Vs
H7GgOErtqlLtmMf+tEEfrMSdpMHaarkCxUqtXF3uZr1nM0Jw/6xjoB037Kn5xbisZj1rodJDpEAN
EZon6h3v3vaaAGki1w+CN/R1vEyusa1O9atyh45uI00GO7ND1YrGqsaM2uW2FGbrHCAQ0RHq78PV
BJMWuZl6Q1xbkDwVM66uR/Pnbo8aZMWHWAtgIf7t1otb4W3Hrj5OGYU9iF20ONiGnvMBOe1pBd1m
l95Kgh1H4+AduinNLrBnKju7J9KiekqHXx4O2JundNWwkSRfOgyzO0/FBL3SWIzingCHzGkNKsto
fJonqsf7XwigkiYl45JmWgkKly4/RSuJB5SHEOCrV9PdHEAcvxCl4MH5hKng1ELWbHXsBJT1en9R
Ls3s3k92N2l5Y6JxHTZYLWQXo4l0Cxqg2d0jHhuuja3TQHqqjqlQk7OeabSu13a6lbheCdOk7XQy
g1ZSICmdCcA3TWOWU+h/v89iVU1mikNWGuXfnuwpN2qihRR/ysVNVYl2PtjuB8330BUdPQM1t+ui
v3jXht944eCx9Kb4wYG2ruzAmoPRto5i1VrobCm92L/qE91qsynOEkICtNLWx0wzjmEsgh37rND5
bmRPPZYl+dACqEmYvqn/2LWF0DYB88A06zA1pxLSWu7J6uz43TApCJt40KjqBdJj5CQ5PbxeovT/
8YXSy/rvI/MuS1f/H+XbO0mda7qm6B4z9o/mqLR4f5+5oPrCnyLcRPrOl2mYx2YZgNPllUg8zsfh
L4yIqwilZMY7N2XWaaPpl8j3suyeU9OMsgY6nC/FnIF4FAoa1rq/ZsZKhjgp7nhkmgJOGxiDfuxA
EJbc1dN/ejJT/jS/L8vMHIfsccWnXcV9/k33BQeBGPiMghvbqm6hkg3uz5MIE8Q+IDjF+73zw184
7SwZovzIF80x+NS+/2c66t2KA9q5DavgoTm2pnnrXWNjZn0Z2CAnrwANnQV3PzHaJ3gN95+OAMNE
6/uYUPPUs/DTPkeSdFm9xupnBukthErUqXeEbo2Ibkfhv/gdjpvKnvmxavt5tSUxlRjiNqU1oBJp
LfYAfg7bknAY97cAPSrxpOxjVoG0YKPgaHPpApVpHe6gA0R5GGmH+tplTfeAIjoYWgHKtFnOQOzY
pMNKgEPgy1bTJSHNzt+n/nm+lEZQ7Tp0nJIuEVDkB6f5zagQ+2RFoNMqkmDXq/++vMx3JLn37pRN
O116cmGCAFhYzPFkkyeU6Jm4YjXRdnmeTYoAh5RtRxxI6HyJrXk5JoIuDulu3HrMI01kOxjyjDpx
XXct6Yc3TIs8oh11G8/uy35akDywnd85khuoHSTCK7qJAZjSJ3/Gl4rAvZae/gw+3MDgj6g7PwV4
p4qcB/jcX2eod3VBxlAoSXXBeUowsQtfPuDRIBNPbkmnfLTxy6OGfeLsrrzkZQBhejP9QSf3o+h+
r9NUzoxTF3U32FvvymleP9VH2mByp1b2nbRlukq348XkIM3jvfSDqPGzlmgJWvIwm7U9xq0zG656
hEdFRer4MKCvlcVEf7Eshyzfx8Ny7Q88n/jTFIlcd/Y/Z18+RH3T4DdcGlOH+i4hZv7GN4re+I7N
JstlrcwBmLM0KX9G3auMRO5iNbZoHcwsW/p+2fSqSVFK7JcFgKIuqfXW+cGuxK8TAGOczL/xpVGo
OWsC9effb+wXfTNhT8aoMaA5ImPf7mUxyuTsctpm4YE9SG4mkLIBOKCYeA/o1fWg0/sfWDiRy3Uh
C4y8Lefvqrdzgm/lOpYU0kwe1vp8k0Dqbt7xAz9xwmLmLwTyevIAYcfp/o8p0tpAM3ZN19Z+9/Ef
HSeh7VfFbRrCSFOS+v+ZwJCtxvlRgFPP5IYe2ouC4ajUFNyBh500CT4r8q7t+ZbP2FspE67E3ACT
gKdair1Sy2GEx1K4SRLCflAfJyScs9l0/U+8/owYDFrcQPKs4R4Gvv84e02gzrXJfPuGX0agPLhb
H73UE5ReA/d5kANVBKU2IS2eHiAjxxA3C/uZp8YN4KU4MWV8n+EqbT8r2CaI/jWhB1vsoeWwU/so
78xD0J8lYdeV6CquntUSKCvHoQpQ5YbtPPh2QuGRFacndvDfhgXmhRs+ApdwrimJFekfhQ65RJtp
Q9dhr26JmSvuvUZZKHlmgGA8x5n6kdHclTVT9KIomd1v0qP2ncWawBeOpwTFuOEjUkcr90e/sUSP
9Pz+R5lQ73HMzpGY/1ugOC1KXqb4rJrO9yHUZijlB64AZrlvmsvRfGzhuhIaL4J7PzuBPjhuQOSv
n5rPRZr7f3u0p3NQ7TY1a2N0WD2nL/5t041uUQ+NjYplXopn5ezgWn3ZGJkH4cVZC38KcsyNxpn2
pbrL+mbQq00XCBpLgXEYE+kly8XkPjZ2xC9jdPJppLW5MDtG8LkK+jxpua6M9mo8kfJWD3zTegLf
Bz4Ud/i+vKkgY5gvzT22yw4eIK4EptA4YU2ZBzXY0/XYNItSGtOboSGnEELYxGbDjGClGSyfwSeA
U59kuViLL/NdIFXK9K3c54x415LYleR6ve4u2wmxnbOjt++qfs91d5tSSrj4NfzYdGKu+R2/jvfr
cnmmClPfTuHMW8tvmYT4cDnsDvDHaeTpHt8bx5FrcTLSYCY9Wj5juc/59MC0C2bzIMm7FaplRnW0
pEj7pDCUK4Xw1mXZ1akmte6R23kDHQ99YMP1HHp/1aGskHYxUL0VR4bs+bj9vWl0XuukQsWiRGiu
1omL4ciMC8Vnbi8VZ9tnHPpfx6twN4Aq1WicB+wD7h/obsX8zZfHkjzGV4kAGd8AdHKOxnWhATN3
pzX0NIfbFOaWGUOltQCVNyZeYlu+HXP4aLp6mp+rOFVCA3bGUAvszXhQf4xWsWILpOvTATj3H4C3
J+XQnxsjpQZliAq4sdUnF9OlQTqnRPexLX+Pt9VOC1kn2bR2snS0BldAYx/CA3r7Z4Tr3gEzIivR
vN3LOL/mBV6wFbDWCT7GEt70R9LZJVUDOfP+09qpEjHW4mCZzFlioKMP96d+HlQAGHIJxTQ2bvPP
EZnY7PE3ceLs2wd0p2Yjb8qnpiobjaxnOez5ZsUfm7F2pgkTObY7CnKWjiZGC/Ij1EQxDUWc5ggn
JRCdPBEXsohdSn/JIYk6Rr/J8M5TyyvNzBACSdH6NkonYuI/LdUVLLAVs5eGUR7MjR+w5ppjuXSI
ROSl1er9Jtn7nRJ2sBVl1LHXXds6KUG1GuETbnpr33u+B/90TvRalzq9FuHC4KnT4G1bcK9WUErW
5woHG1suyUMt4gvSRMpNkhXYvK57NJNPjnIEJkBkLAamsDd7qqoS2I6gb5KUIYfYLL15MiBtBbeU
cjhb7PEhCVZG0OWh2T7Exay89bM4OFpnB8cQowmR0MkXyTh8RljKtfPMslZG5YDagr94Dndtrdvf
kguM16ZLLKjjYrvCNPhpScqm2VrpZhKidph1fTaIQVB3f1xeo4i/fHC04xSHQwdRZjaEHlZvCWzD
tuezH4PhnuoIuq4i2ftA7AljRPJHT94OHOIoBWwtyFi/TY2cENmucoOkh4DymK/F2CYRTbo0sRfc
Ioq+AE5yPi3JLIbCOxT8yJMI4rnk4aKv8I+K7mAw5bUsyKLzpq7rnuh1y8LU3uIs6/F8EoH9J6vX
q0DB0M9Jafmg5UrAVPp50DacPrr30f5+g+xSbHyVeAFTl0cZFEYqMii0Z+9eI4WpEQcXmeBduqqy
+ve4dLPd41bJ87ZZwCVE7Js7g7FOYmw6Kg/TAI7RfF++lrCS62ARhQye5gIenQJW7avld+DWnk5u
iJTDEUimpxQYmwcZRY7p2EahynZj26Kco8q8VIle13E2CXQQTpYuwYVS1PDBf2FuuSITYPQ9doTV
qEYAhyW3EYFCEa8Ce9kCWjqqVd3sZjX4Sb4T86dkBwR1dFGGhRi288cY4pOtjELtBOFSJWfKSDk9
MJwGRE9vX8szYBlnZ+2o3GzA6OV7c+Cr/QwjXTeslD7Bu+nAnTYPs/CMs69uvPh3BDT1GJ3I4ujI
YrLj06FWUTCAseV7njUkdku2AgIpD6osx8l4bX7lr0DziV2bIhHgOo/fncmIPayFixK9lJdoalu5
ubdSKg5ZXQQ+pyOWosAqYShJO4xSpLh7JDzCiHodLA2s+AkWiqAT5pcPVf035BvSAFEBYjrjnkDY
ro0MZnzoKiIUSfZJlvR/DZc4JNpNL8s1I0R3s5YvEqHWeA7oEqP9DqrzYxSY8fW+qNY0FvNRDWkb
ykumsy2kmifgQ4WUGt/8bOjflicYorz8JN6PN56znWW0ADWoAWLwLQrC6rSBFh1iESyAjhCFaRwV
X0WQdq9vvsDkX+fqxy52BdPFL0KuG8FNUk/zh/6Pgm2jl9tv30rlyEv/PGLyRDTWKn8nMQ0O/HqI
tY87XrjZ4uWi85COZpALwks+8dYaPTH/mMUPKYTsPT+3zyhBelHYnP8insmqpNsm79FzRVhW+94a
wDgl62AbRRgZqUt++jOKdz7SHVgwjApCwK5HbyETz8PBRj0x2jPMUGaiX4CEV/FoZdQXRvIVtnN3
D+AG7i5Prn73jg1yuq/Q8J8R6GU9E9Fa8Z7Db3Jx5Id7HhyaC5uTOm+1gMT9RcUkKmYjFTNste+4
qv463g28dgyCTldRtOnt2QmeeGEaiQzZCJn/BZ6Q3gRm2JxD1dmN6nGnm3QvPvqaEjwMbXIFJZvi
KvW/m14PiR3ekEbhul0BLxf8kY+Otnx5DGRS5ITBdrQmjR2Bq0WF0cST5MpC4SF+fbTxjsft+2Tb
9O43YaiNbTESLPE1tQzIZawr8p+TOILZoQtXfTqxo+w0qFPDMGBFLGQfUPam3AfIja+Q48Vt/Sb/
Nx7qiURkwFG8eYqNqyv9LlT+H1WP0QrlTo3PQlWwroDQel7CDO4JmVY1qXsajlciZvsVmvX1Gjbr
9v5tbpL2PrLNja19eoIKkY9LN02/IC7ovo1k71m0cXhsyjyOt83aA2MWRzcHDPWMLN9p1Gfxj7WY
HhCTMSJ/Ya3rGwvj9fv0DOOKqDxboHY4L+Lv9GxeSAcq+/C4WeaRAwqygiwlzlZ02J8CrFTGdzoq
NLJ52q+zPC/4J4hdWY3V05q0WqCZhczBt9eKtpe+7DgJPd+ZD5w/4Qkj58VfZaRzru5x3R17LShD
lDnu26xxzJcx8yZZJMuiJOo2G3IejljGr5vmIjjGWuW7Gaa7G6oZGOrc+oXLbRrjxZa9eLXx8J1j
JEzJLmf3tZZ/APQgjQTuTnL6Y0Rnhz6yiCwxO/GpgayZyCvfJJAzp/6NQ367pNRllYYD8UAlaY7o
+FebU1w2lNActnYKWGX6xASKKdXCbLSN5XyM62HpLGxgMCN2borTLJ4ApKdVnV5exQ/VRRF7Dx5Q
VSRLZpHn3i/xFiTymy4TRMhUXJ4izAH+CdbhJFHwD6AYFrXnRwSuQEDuzUcw+UhNV0gvrJ9AY5Pu
m0ERqodPe1X/xRVzZmAIuvJe451JpuWIHwgO0LJgrWB4xxK9BwSzRnDcV1nB/OeDc7A1JnD1Zr5N
sa+3L9vIpaeYgF5lsf8I4I6yhNDHIMHkg//0XOjYFEwT4l88PrKUCmgJhXXZQJ3/p3x8tu2aUM9C
s0J0zWKTf2lcRXsmCgcTZkwcnm/Satz/flMxROxmHvHCGRiqbhr0TpzyXpl6OInGz/IeyesvpDF3
blb3nLRkzr6koV+0b8SNiUXaPBC7GtkzeIG0xXRVRpbZN5nj6WMDv5sue66/bkNucYzRBsaT6SDy
040ZC+Ma8WkYc5q1KuahfMv+W1aIts+mawD0oipNGs8CxP6M6BkjVBQT9mC0eJNY67vRANwhdx9g
dG6JUM7BSvhRMcasnQ0pWxPLAsINPutZkAXP8DjLcMD8HR2b2jJ0BF+6uEBIupokxVgX5seABJuK
yhpIAIxCAkw/sqKPd85OrBOcUjoFoTzAL+CBIFcyLzwnJUt1rimLmpYyLRqALGA2UReOIU74h0k+
fXrMWfMi7k9ubuyN9C2Y/sXn2PfTfY4P0HuxvLsjIFkasPF/0xum/Ae8TijnSQOClR2PwpW5/kmD
1CscVmvoFjemfMr7s7BcBPRlVojIvHn/AeqySWDiQmhByIWFgCfeYo9QH0BY9GPswAvg1T8K+h/j
mUwXovZV1fAw3/Y5o0+PDZWvvjDna+36jhXIrQrxanrlJbqUevCGTxugHsNFpLaSvn2cLMsq+ZTS
VdBU88+8Cza4Jsp7DvxKbqrQf5LzkejDDnvS6sMx2htzBt8MT4j2jdG2+zVmE9r7f47vPbq3lHwv
ufpb0iT6C5+1/2FOZxogwl1wbgOwM7DK2zW3gLf0Rn/il/8IO70RzAxUMUsOU70eUr+PLtEbh4eX
FVyQsrBSlqW4Ra8n1F1z5gn6FUYMdC3Y+xmurCMzr6UUx8VClvltPklE4boQtv28LkjdRcTUj+yJ
/pruSERCGYgnaNswYPlrvXK5NdCPbEBnIczQTac+kT9ySsMa2aZYcY32de+BObqs7Tia+cZ20k65
BVtX+7L1584ra57qX7+FRcvvxQwJvQt2SCPDX7/Q5RFmKtxpaApIt/tCah7KPcEv1JCYyYvp2pUZ
PP2zXkUvNwM5VvFPp2sGU4TtdGwtKP/AI0hp3ceyN4V2EQnu2sK/+6eSyVDWa7tvzl7KmS4Bc3df
J7sBUMmcwNlpGMYpk/OWOcwHIj9nczKBKgy401T7F4YhBDFTc5RBRhpLjxckpkjZnFLZ+HVSOxYC
6taWcLen6bIVydSv3e/fgeddWn/G8xZNxEzgfpCt+7xlLLx3gv7XHx4tSZruinSfSXZ5qwkrN8EN
+xcNYGIgZLd9oPf/kxrSfAIYJ0pJglrYB/pQ5/zDhTWJoYIaU8IcWTyM2Ln38haJ6ipT1XxJYp+R
er2Yqle4mU06e+GdFvGS7SG6fRdAunfQrs9jjVo4dqqPa/0uER+OEup6Os6XFRQhsUB0+5JEHyJB
iY5urAe3qpU7wboCzSlmc6HD5BDmOXGb5Hegn7XbBKONVvSqVGFjikU9An/9CnexyIfCMCpaaZVw
DzcIKHBeN7cKpsParuLkmYyJDjHlDCdbNYK0FJOsjlsAKJkFi+dVom9gFKo7oZ4i0sQqRPgTearF
mQrpgXEDoqQe89/3xsTBVxbJwhRqQOdWQAEi3zFJ1ta74LP58t/kozZy7HVvZHKoEbLHEoV9k+72
/A9v05SInw3rjL6OTWQ2QR59jxHSQNg9/GvbUynYQKeD1+HFtJ9EvkQOqHtJF6OTBMWFttQh7xnk
k/N11hiNCtDZ9yw+wHbxpmK14QYAvzj0OwImJUaw+e8+A2npRudajUFlbUtvgprTkm9shmhb+nFH
cQ4P4QZL1uxWfjNCv96MF0MuLag1xBAPfbrrWLWZsAweE+X4zOrMJwCSztH5XNd7r5OBezXSm8fD
3wDKOY70Rn+tj6cq+VCHi+bzr3JrzNgjCnCf7pd2XRDjCcL1+ZqM6oIzKi+PMuvp1UQt0k6M0ss8
z3YBPw2WWB1EwPFqzzYZtZ7ZPnTxiANvb+fS3AGLoMHpZqM8zMZ/nvBwi8imQMgJLtdwx7BOlJYP
xbM+n9+JGn3CK5N18Bo+SYmPU7rwecazpCHndloPqkjW6uP2A7jOYlUoi0RI4vnNChtPL9y+h0n3
eKK6qYZVUCxBX97BAcsq8Odq9lAeGfkOlM6zTNtyvQvmGTiYjagm1bZg5sXgNhbM1ppXaU5/teZW
90mB7eA/jFQJJgyKdcvnRTDDlPkVTCC6m7kd+H/GFKrov+iG2Nl70PUAWnyMFGAuZGeqWvo9a757
/o6UKawT4FIMihAjiy205LDVtWK0vMIPWFA0ieSyV4MWRT2BJW3Bo6zGCyM1vwKj/LnDBVf6tfEw
AqI7cfgj+NF6bTUZlc7hlfaSvoR8nGNwyabMvxfKKUKPu8SCPeMVrAKXCCOn+4TH0h8DTviF8wCG
cyzyVkplMiXHqG7Aml9SnZLvWsn+jLpJbD67CKweMXAUynfs1vX9Uuemfdn83QWx6YMS7NMjXz8C
SSCbch2ee2XuM03G3JoXy1q959TdZ/175lSkvnfo8UEDuyTv/BNrkHmPlCRvjA3dISzgRO7G5H+L
t4GyCTN0JqIJexyBoZZnNcGpegpdwEUKAYoJkBic/wBuq7G6y5BM918imsi2wVSUaHlAqKAFUswW
IHkNWdKPcQQAr7QifZeIIaUTWcMPUdjxGpqR6Zt6vPrzN8l1tMdlJsp9DVgkhRcIdCSn9dVE3JfR
ZNjKzowwNL80TLiV5kZ6FQuK3dGR2hYiK5iry25MiPdIp4nkvLfOim23IAybh43VlbmBroez+aSr
mPDR3D7hfM6XZK2SpOwyfOSXgOg9SJiWOVMLoSTaHfS15SkKh+I62s1aSS/6uEgboYIc0heaftvl
OKV+CiQ90u2GCul1hIgdLORruNYtniW4DFh9BvhaEB3IY9HeIsrs9u6+/2WOUOvcvO/IMTyoeLe/
YOtLkmQ4ZjRofu97Lweti8894VZZdzJ2SlDsdEdMzX4SxHjBZcwwOYawEyDwUHQhmmlDgReaHME5
fE6vyPVB1u6XQH8p8/aLiLoUzySfD3pcbgA0Zrb7wxxNzTe8k9z8ZfzN1oJRSZWEIpy/yyPLEH2s
SjeEmkgjUbGxHHdVZcvLZdmuhBrc2h8h1eibpg3XgRFsNkOIMGKNUy5iyszMhWI5d+RXYpr0c9hm
T9CjFDpUqOihSKeUAiBeGjKMFcCTYmRaFDgmE6OBYKeipjzceNigTWT9i4U13kBhdQIuQEDly2/x
gkTwXWSKU7QXdEiHf5tt/4mqEj6Hs5ymqc1+xyVZIUHdrVzkbefSE2Tp4JZQ0fp8bsrUq7hMeF9I
t+eErnCrNvwUcpJumADwgIaSeySBF1YUADOy+s4XPHyq6CWeli5tqxiM1RobMQLsI5gQvvF8dYwI
wU9O+WP3Kmp+4jMnnolsHger3VEpJQlTQqaHRGpJR3Kda7+2QDXX7RCALuch6lKHkRH3YArJu72K
exaLnzVOMRAKEnIFjX+ELdHSRGbvuOey+u8nA1Pv9pOI1Yp7ihYge+Gn2jCh7Md+vXQBI+ijCfQc
vTeRyddhYt8s7rISsNE5Hi0pJyExIkZ7d0OxkPm0Vz0nxEzkHK341gTKR/KWCF6BDTDo0J2xcG0v
i4gEafrruXYe7DNnABHJ63XfStxSS11RDQGCQ9nrGexHZioxej085EA/ULPzQyfN4U0DvUPMarr4
9hDzDf/4uIVTvUHPbZz+ulJU0BuKOcVnkuB8Ib+7Y6dM+KrDSVOwqVAHRZrafIBProCQQO6N/MbG
AD5Z34/97MKIdmambphWj4S+f7MtFhhzO9YAJJInVeB/5EMuaZoYPqzXhtRzEQTbgyKDvHJhw6rk
cVthrTFlIkzz+GC2bh8h8K4jX7z1AIiEsEE+UzksLTbo+bMeR966X9f6yGyvpAxdqCQoKvUPSIA0
QdNEWNVr772OCKH4CdtfVGXAPgQYwiZ+Djq/tj1QYLNOqvOnaMHb7XNbKG9tB6TK0tDm/UNR5pvX
W/XcD8SCkCYtvtxY/yuQ0sx/uynFmivWUs5SrAeH5eYdXMrNm5gj7dBOgvaCmw9fsxzxjoCDrusd
cvPfNb7l8BVY3Ft+o/XOVifRG14qB7W4o8Q71h/PRd18ZNqVEx9K6EahdxgKl0DHJ3LxZQ/4P2fH
2ws8giLLqXnJJpfy2URRsvrLq/899hv8pjHeh6moggx/FnKj17lYl3WH/r/SXqiuMwlHBWh/VKTJ
JJ4Jl/h5Gm3MP8TYwf0oQsh2HcGOxv3jUju/eMGfgV7JyXbY3RYkx6oiMy7ur7z2V291qCV+lR+h
WQpe81bNKgBTLAowXAhoWQtjbz+zwyj2/tyAYhMyvrtoGkW52YjyoFS77xjfC8kR/zkIbzXkNRS7
eKf0OQTlTH7pujyteaCE/nQ9s/BSWF5bOK7y58cHN+toQWeD4StgP98rXd5XjQV4JqzjUpRSJCU4
Ombg+Q9ml6LlJHrLrK0q0RFism+qr5w+nw3aKyPLGemBTpwd6k0IzguzBzAKJG/a3gTaNvH2Or/s
HuYcVkt2puuRPOrGzvWdhjMx6E8EFSKOlswgPpdy1TJk7aEDnCFFG1RVjKpTPI5GnKvWSlUnGctd
WJRi5FLWePUA6+FYo3wTnu9My47OdF+Ac4UtM1UdrESc7jSc0P0EYr7oasDtPpXbis+k/bVFfONr
UhxQNb5pfslyG454DlFLD5nFv5bKJucpwLD2hC/3lmHyAfi+BB6OE5DaLlIx5EK/5/9pZXXze34H
Pt4J9PlnRsyDx0HHiSexpZZ6/C2v2h30v74Dxsdy4RjoubWRsPMbWtquQimwqrMOGW53vVrsHIlM
KfjCNdvi0qLIohW7JHP9AT8c5Fvfr6DWPPop367oVLzQ+wgJLqY3LYLjhpzGxdOzL1/lZivYW9nt
vV3F4jS7qjgD09+WMX63bWiaHaLb/kWFMBCtovhgmEfhz0lflRM6eD7AIXZL2OBMvxnBopzpczAR
MTVMN3A9zQp7tC15vnbhcljHStWnNZrGoPopqNxlwyzCU3AMy2uHl2C58ZEj/KK1P3KJjD/k/Fnj
5YLtITKcr+8VolFOngcevLTifvs1Lna2SblhhkBr+3xERlI0Z/lxdWfrY1nsFl0nAvW5ICD0DGh5
Eis1P/76tqSp/64iwIlt4DdlGEMGVQjIrUTFDvM5RcfhZUzhyVYP2fUMhZASvBkoHnipBR8hKWJl
wB55vK7GKV7kkgaWwtpFJ/VuBVJcts+SKoi1bock+VIUEs94CyTX2nlDMIfdVhsbKjh0gcLUi2Ex
TKVlSuQ4Rq1FabRRP0y4nLJF30/p6uiR4858r2XqdxbKid2YO8yJ8jvVsvxxddJS1jSw13X/zkWI
zySc4CW1rnr2bm0kD5+lQHuXojBTPt7Ob2BufGXFgFqNiHbXPhFe342I4uM8IcixGtdXQk24ddhV
p4ixDccQ7zlFTxp1MEFF6vnMEJcc+WR/5SWfFeenooJWWMVIndMZ0HKG+Mhi3vHKQ5EJFd4RJHx1
vEyAdeRSvfNrqYvl0PZzJRZYiv0w3k+DUUFeqidLAysTXmSXGgbAxfmX17VIHXRW6QIBaWnMiEKC
Oru2hBmYFDDf/r5xOhPZTnIs6kYqJ8EbAnuz6gXMqs5hmSfULZzm4SVJcUb4C8qJarL3/HtfL2b6
CwlNjO1eiszLu0LCppjbTxKe1Bw7ar9aDHc0QjNVQ/prb89Lyjx5VptwxwVFL+j6XVH45s8/eKkj
4rehNOL6Z11+5RInz+tZgAtYfh1sc5vUrQpXQeyROszTMD+V0s2aOcoEYTLfyAw9xCFpNYHJ+YzZ
cNRVqFsv/zKajoKw5NVQjC/o1juks3wRwl3661EUL+y84r7NEDkMUMtFm7cUZASwz5fRsCn5ArkR
Vh6IvGBYcdgJPvpdr5kbz4kVsQZzN6tuvwDxJsvTT9lzN/43N1oOvlhE4IvCtvIr13HMIUTUbbdl
3mOJuYYrNgsWcOreykgiI14ToCaa5b/p9Ecz1oYMa8s1Lo+0E9wuK9guxwdhWRFaR79gT7pDA+ck
HmJR5blHE7XgaZPISzHYucpjX1MFAPC6ciXf1+7NUuXmEGv0yADJXFodgim1LOZBfgtRHm9NB8mO
sYEpXPvr3k8rkYujitx69dcZnU8XNATS3o2F8waDxLAZoNyuWIT2HdP+nz3aZMLiJA7gAOMNjDg8
VrmrKG2g7zZy5yhilMx/JCwAXANdu28aYPis0DD8WoF5N6MroY6tN/jeFYLa/siJFPiJNYcyuynQ
4Zr/cSEtuPolFxXZjfPqu7fg+8zGjW7U0u2E9wjbnbZQ2g9vN2YZHSj+sVtHgbVSoTFKmqmA7QtN
hy/0QFn6EXX/G+/Ke6aQTjbIfiEPBV+0vzYNu3RyugaqN5Q5+ET+VELl+3wGzBrB6qgSVA7cqBk3
6AEc34TGnebnXpDAVp3b2eznmljg1AhMermSV4jY4atv3s6VCXm25ZF4EWnSKnVqNGfkR2UZO7Gf
K0Jf4/kwZb2IE2NiWSZYS3DC/UWodDsPRjSS+X9K1KBTmCCeTJ6QyrYBmLqxpewroSYr6kdbDDqs
4JlvSSzAuIuTBu0RpBHs95bEp8Q0rZu5eWJ3cFiNGIKg1JWjRxdf4PFFj3kvjGxmLJDOeAMVQ8XE
KsSX8tYwdS33QtMOA6ObrZydn/OxSmxbaa0y1dKaTfolxumvyqGWvbPu23Dw46iSUJNM6Bf8OoT8
w5d52Efhs9515m2BjfvQHHnzwFkN32qJfYfpxCJfmel7Fk9zBBjy7H5AKTxVb8iXe4duCk2ZrlkK
PNBYh2low2PURyEvpGgDyjn8adpBXCa3xssX4gVQoafV/pAj3uKg0RZrJ38YSnR6zE4GZT2ms1nD
gnLtbBCP38OpXRCJkToYwloXqSdzF5PTHcW6A5dpHMtSL0U6l5KcepKUOGkXh7ihy/LB8lhCdmWu
vn3TMWqFfsmx6wJ7ocXZ+z4opaL5MBwEeyFsrOMnwMm/aBZamYggSq785XNlc7mb6ogYbAyJ//WI
cpZlbWXYcZhWvsKVPfVDphm+IJlJleN0DggdQBy1yZrt2NwDb6lTf4PBvFiTqVwqBsGkQgmzb2wF
cnQPN5b3mBA7Pv8tA1zImbr8sLluJ06CgsLJ6yg+CSEl3QGXasscNHIAnUK/352SGswgO0o14OyE
JMlhkXjg6vKcYE8m5cjEFmV0/78DD+/NO/+/D1cj8Yn8zYtnVkc6D6we6ZU/KqMjSFHmSwEiaGpw
rprICP2tv0RKFWR0AroB4PHa+5SftX52EcSdYUxMWhrngkL4GJLLZ2zbF4ueiKe6DtfCqAdyHlSW
Gj6S1mAzjfDdRziXANSj4n93ZfEgJZvp8DgFU0FbOAAXLOgyRsrgCC+vXl6prrHN4XG4+XBqIcV0
aiLFf+beBR24yt51GY34hpEa9x91HhT/hI+JYLoWAsf3s6XoODxiRQdkcMDmCv4JdFGGzetKKqI/
WdXb9PHcsD1H6jt3iB2psyKUr1NVoCgbUE9K0zAUiq5f3pAfcoO9cutHfd/jjmnnnPpoCBCQfaT0
rd1sxhIUitN0uv4S0nCemrxSC1vMr+DwTmrnukx8o5ybCMYryOQqlmkAifSse32S/SPdPBUv4mhw
dh0tFDuCDKRPwwkzE3erEfulyzLGAMHsorJDUw5Nq/uaUa/LjoDOBgDlK2X2Wu9eWBO6ZNkAg009
miPzJiKCB2ObKefYQEUjgcCUDZ0mfv+jLM2miSJfw7C+7n/eyBCp6UEvkLAD8f3ocFEyx8EwYciR
TRof1a2cL1Mqs79aXoiJAlOC6iIXF1Hbza0aBoLkOMmJl6T4/Nq4hCkwNOhccT0QF/7tXO6MfsdY
7KuBO5OKKzTWRyJMeK4M+ck2UqJlkh7iQhrsc1CqNT03wET/xU1L/LGQoAu0mtWVetnvH325gxON
1t8m7U9Mu+cJs2pDJsSbXndhWve35m4kjQGhHZ++xY0hCS+u0HOPDbrbqU8ZCggX/ilVJdKDtys/
/cf0Y62DQ6StTSgcAM5+HhGgX8cWbKGfip+Ltjp2q14zqVAuhRXhHBnJTgT6LSuGPpB9EwOGgcsG
23/y6BYj1t11D3D/woyiXVOUKPS6AVE4K0m9deZ+OnGt1T0nEV5FcHmFk50w8mRlAWGKit8m9dgR
Tp4Ds/RbI/JIYtgCPrM6CsRVSumBWe0mLs6f2xoL4atvUTyfn7CVEXWojjCA8gm+UPCOx6C9uDnT
THM4ju+nfv9QdqVlE6CAtKVj9AykKgyadv4kjynE3r0yapLM5jZwL4OcJMhnn282BkqZEmgAh04c
GKn65tlinwrLFpTNFRZQpqrXwW3ooKS8yanC+FjSpfm7oFXku246FiZf9jyPxrEby+S9QTKH2fZP
bklrc+wEF0KXLZRDaBO8bij9RVn28I64KptwdPLG7wZxngZA99dRVlFV+b7iA3xMlY3s7uh7VJk4
k/KsdmySYR1Yv1uOfz4B/5E35L7RdFSfdwMrwJH89dlVOYaIyyEDwjlOp9/GEo7aDzNMPfee3lPh
+ApuxNrNN95di0ec/hggz+HaD5IboNVbfXd2ZytFFXFFhSNaCKt/bYVxNJAqW+1s5T6ghZdakzro
lW58raqt/BlXR/gxFbu3JjKBBQj0Ai3WGes1Hu+7/4UWV1Asd6yZUncdZa+8tQEv2e+riMFi0kge
b630JSnyVGoJUa+ztsDoMU+fiSh3lbDL275/ZpybmTDonNztecQjUX2fNjFrukxBawvsac+OEYgG
a43qLPfn9NxTezFpzXJnOvqfZmd5qUG3z3F+OlQmA4IxiOvvrvU6bNWZxTyYqJG6mlr6sRzNdlyi
kZnC4eIcJw3jxuzg/T5Eeea9eG4iwvGQu70oH4gaNqS3Ibz0kjIFou5FGKgNpg1DuQNfZQNfksRo
HkSmAtVD8UYTdQ4KqMlDUVvWqOR8KP+PoBXyJwtfnxAql4s98xrE7QRDgAxrxs+LUkhLpxC5lA7j
d0rsUrTqD214jIQTRMRYqpcCpWod+ocV4eqsW0ACG89iH8U75rrEXDN/pP4YwAx3BsPVT1uVpXR0
ZkuvngHrYbGiMqQeEZR2PqJ65VRbF2yrJj3XSoUKTGFHGt3xW4FbhAr0OBRVGAd89R5RN9Rdk0ky
QrtgpU/3A61ik5dkAFFPdbOgO4T6GwN6iarZK9LrsVoXkVKPq/0WEdmSSWkVdQnUYbUT8tMt00X5
Xq/ofNxqDLrV1PvdVA3aMW23nF4ozI5x0VoPRGFT8etOetqaZX1NulZCLYgxuGxAA01XlFbYWUoL
FXKZuNuxyMVxY6nFjjTtu8f668s8+G7EkdM25RBEex7g09ahbfY8FDGTe2C6/LZPZ//1VQStwU7U
9e2/Ku54JMLzqXBWbMpxA+xHKKX7/ss8SJaQg74/ZDfzXO6EcNSxBb/7kSf1PGSvkB08d0Rq53a3
5iCe/YSfhGYhbOGPjFVPUnsjpYGvfXX3ARXT0I2dZxC+tx4SaIw7j5CqVpk4umpMPq9HwbqvtRCk
0EBl/JKUaDSGx5MN8ueqw4q3QMM/T1A260wt1QMVclOxpE0od0GFB1M19o+Tc9M48KzTdaCaNxwj
cLxkxFYv2mPII0J9e3ySUArE6rIg3lEVU8I+QS+Joi+7zEVuU/6VlImHsgB5H9trn3/xxpTq8ilo
Ql+pNnOxOT96MoRqMEOlRnKgu1Q4nPPXMxtZJmlEjXCtuSphKJcjskoyH1SK2nHa0ky+6qs+9LjN
ZxtyNlHVXKqSoj1d/3TBHS42P1RdeIZl7o98rTm3uYt4SAvZDWA4tVcWhpnVgwWobWBvUFiJCUtW
/dMPBLEttC0fHleg8hlykoZONc82cXi7XUPkxFHSeoserNv+gHInptm9ZtZIMJa/JhnRRU9IC8K9
nhlRKFKJGnY6ofwX/N5Eyqi30Ug+czvMiKW52kvbNzFVhJKQRrFztsEEEgFE4wDKdYQ0eGVRjMZ0
ZQTCGfWhboZxHLF283owLRSmi495X/xPMiXWqf5nKel6q0lwYSewAydRN3lJl0DuuAz/ZoWiDBf3
IERdeo3H2I9P9ALg9EtDv6RUr0ME7zEQyrLPH8h/qG9mDm4A+dgS6srNVZ+Bq4ag21nJpQO2+HRp
VTrOCpJnW0T8/tQzdk1jbbkGzWMt9Vzqj7YLyR7l4Umf2EItJ8REWgEfhoaa75ckIuHnBKng4nYn
AhhTc0jsmybRMPF+vwuLZax7wHEzHrdqMeNZHYLTJP9XXAcWIAvYh4rw82lLNQ5Bhf3xgN+h1ZUW
XCFQNKT9kJuE3I4fSyZeisyhFCjU6LXsgHeswSNOafcJO3MyY1xMi2awsU4511yaXEQBQVhf3TWq
1iwVD96DnROhCV4j7Vv+GjB9FJ/EjAj64WKy1Fvjswgds4K0Zcn0rdPTuoCeu/mtd+8n1N2bVNM1
QM/eE4vjhGKQriSQxYVLhE3fAb5pe4mRSo7WR8xkVAejolO+PWcBwkC/VFEY46Qty95mQCwl3A7Y
c2N1nMjR9cxE3ExVVBA8My0Oi5b021mcJWNpfGx4ltMAcLzjyBOZ0G+eyIBV9c6T7552e0pkI9TL
k5D2umaiwMLCBNQpsvOhsyE41WlKVpH5z15+Jn3ZleuAO8g84V6JQm9JV7uf7jEmom3E1sSwqfBX
kN14PIaD63rGwBZX2euaah5VzGJxsNjJjVW0m9gfTVmqrs1A/OdqvNPT5hBEJQsxogbqBaSBpvxa
9Izu6sDgCIjH3QSNVhDMCxv+JVqVEOwZ8fVSPWM8cBSoxkBKTiobQ5fm0JG/TK5A98erNy+5MQeP
iHsmf/RG9Sles66T50Biosu+DrVVnbyJGZEERw+D78+zBRXweZEnWz7E3qwet2Aa5mdifOaeLlTg
d8k0okAtC39Ii+cxeh38UaEMPNcU6B4pzzDyw+9c8s9Gl/VOluhkcL4RtjXBH1IJETWaYJaLiGhr
H86351U1DnO3ZPGfdUR9vF2TFNwAeVMO8dXn4oCzHEMb0F8OtOXjO8WZQUohu2XOgmahCeIQv9Hz
Z7DFwj1Vn6JKtA/JSiTa0PX8eiZ51n5264BO4F0Qm5+o9UXizv54wwzs1VXVghxNr4OE3A7CKkfh
J6Ome7oy2XOLRUwTdk0C/FDOXZGVkEY+ELYXldFwZ1sMPAWrg7LM1VA89peTRkq1077GoXBaM9Kd
eMTzrHbsF+wDxPkBOIYiizNnmBiO4QlU2gHe1GFksDMRnnFM8Jfa4ewv7JsibP9eyRCMPA3JjyfS
Ql2XWrj0/P629s9kxwh97ZgWE0zvh7iLwyHICxouN/88QuQmqyLBonOv6MBSpvmAco0U+Y5Ch9jU
ehvk/ww7Rju5SjwpAMlhmeMjcoD5oJQu2bM5sHOK78O27HtML5ofzZcRtUQENQcX6F47NoQaHacH
+ruAIlOc2vcCrYpl+540cRy16MEabTZ83zGMU3AAZD9XRt7DQCSwcVtCJa22vElREb3Hqm/ys1Re
3rq7x45TbcLcG52DZE+EO2xcFwQCv2vhasTUZEo6m0tPz7HoCsi/CIr15Li3mUOFr5mlufxI+Gaf
PwJtIfLPECFJXS9l1rRmkBUkqde64oMZ9JId/tKNCuNXDaQpl0cZFvcnna/UU6MhQEIwXU5zEg1p
xIPgJIHkD2SM5xXWJTcUSqk18f2ENlN+kEXGx8lXiWUxGeeKicgd4PO/pomTDbgRzUghAAfETtwT
b3a8FW9/EEU1tjNAOnxj87AohSaiZaKJHDpHPZTMmtxAYyNtkXFkcMzeETJfJ2kthjOl/CwKWgRg
fhrEAXApi2KRIYmbqE4l5mE0YfCZ5PckTKS1bNvaO0UWpbp/E6Hspm6DhIGpulheldt0ki/MlyIc
I8cRGyL04kt1lt7W+p0po7Y56UJMM2uXXSH362cAFsQHeX5sE7m7nC37nIzJGyhTkGp4ow/kUzOZ
wELnDD9u1xIlofPeoHEb7MsDaq3pd4Vxlinl0N7Dx+nzt+UrWeH0zdZ5aKqok2bknvIbhBO8PQJf
Tnzk+7VHnJgO1vj1N7AvMEKtw1bfHPB5qTCFtPq5FDUulfEfuLIHkWOnitRfhJK/BAylUAZMbGdU
kh9icq85EF2NvFIlYyH/EKTT0Q0HBOaPapZcm6+nl+71shE+m+dIkuHoufn5Pu720lHY/to3XCdd
Ahk7seJDx/lv/l9f4POup+fxm1mk1yx2WEKZAjdvq/aH7Mx0tChQUSjgRzPRIVox+S8MOjiBqnan
5xDFeKIZZRiGfuTwOFPJviNkp4W1mTqZDaIRGgB33kWZQCVmncCbtOYfBMFA+eEdBuUjhvFqfLPF
AVvhQAfbD/HUy9+UMO0gS5vpdNBaDbgbFmkluvFcltEIbir7UOBl7VX6hRmWnZxVH/vt+HpuIU7s
8Px8C9HHhiL+ecE82kdLy9UBJbu5qUruk6EyJu6YJ+cIKGruiTb9s71OznOBX1bn6mrFb5U0nGo+
R9gR6c7+whnLal4FiOGEaF+14UFCKbWMFZLLQDP0fYwCcNKiclHoNvZaw2stcA0dWekUtyv4bXhr
kkdtzqTLD1dGrCtDCYZEVktYC6uvEpwcllfHlia3Bpjw4M5nZv/cdCJmhc2jEoQ2P41iO8GLfR3k
eLu48vwXkvM9BIKO5TUYza2gd2rpkG+hpN3mNXzbFQlaL2GEC+ThXdrT+ltRx7QsEjfveEAoh6Y0
H0v2/ioA91W0cj8XuBnzsFoSxupON7Yl5MKdQkJj+w/u6JEtUnkkBpAdUvKQkqa885te8EVXAS48
XfhiUProBiVLZO9vVKtXZYC/uVu2toN5igVEvz2YMDaWZcsDWowS6lDALGQfOTX75EpR+UDUwads
Thbdpopi2d9buUz4RjYRbue/786Xq6dTC31itJ0QouPToHfVEiEFeDfhuBwvEL3IN5RsTgtQl7Ly
EEhycmWwRGSAMTiwicNLE2BQwAbSqdZMZsjbkoPK1Msi8y0jrWm3UfW+ncLmdfFVoMqbfjX8jEU6
xg0PoYoduEs3Hov5LrG6M3dKkOCy6sV8HG3lJYZQX+FYKOFcOMp3GTZld4Z31cNufEBI1rVNp0as
qiLg1lTj7puUNypBITGhEZL9MGBscnl1mLFWVdQcZ4nCEMNrHMeA3nznujFmjitt8UhCjJoRqcql
bDfts+/+grPP/UTTUQAUPdk3tj5G2rglzOom4ZX/+Ed+JoTuoDn7/tDSYxxSQ6W8dHDQFUeEa/uY
YSYFMRlodGvbg2fvBYrlnEt5KbGObJp7pQv3Kr279bhz8xVcUpXleCnSykd3fvA89k98dRqz0I4R
q4Igo6dL6rmggN/sDskqeAhWYpkSdPu+6F9s7Dn4BLc5bTAuHiTZAlZfHo3prscm1ANRRy7LDfFp
udpg7Mx/lnfqvF6LfC+iPAKvNQyVgGfeypdjMN7LZcJPuiKcN5EOJ+91CcHb1LPCr1cZ5SiS62y2
h07p2tfXOjcTEg+RtPJ20870dyc8eEbYxK9eXex2dN6Z+ibrqKVqjV+2x6FjHZ1IrOW785LGs7g8
ZqnRaJPRoVt+xQe42lZHGu+cK7hVnEIX5XRmUhPRGvjVsJ53siIfBFGboqOcIH3DQz9WwOY7mMsL
EpqcROmMCOctOf+jef8KFMynARx92uoZMNIjNXjWC55PPzTVQiwfyt/KZLxRdcnmZjDSLlGlE/zb
zJRHCzNdNSzUljgWJeFsF4lsui40pS7eM7FImvFnWlJp2hU4i82zD2qmfe9zDirGdmsz1aQPy4aN
gNfdpeUSZJvi8/R4LhqeghRuuzwSdojwUEQKXU706UzTO4QG2//InLkPk7JU8VgPFJ0C5RqQznM6
+P2EVggSGqfOlNseBI1wJ7Hp+fUJFCFtHSlRwP6++HsRa772JxmCnPJY5jv58N0+acrm0qpvLbsQ
9EpPrNBw/TkvXckXbUKGnNOQgary5vZDYKvSTg3QVWhKLqbPeraeXC3nc7V14ujoDtA7J1mxd/iq
p1sx6Uwc8hErrU4Zwk0zBRij93eJ51asWMBiB9FQfwJDTv0puCM31nXEmaExKbcQom6ld21rM62d
Kfa61sj5xQmOXjGeIDg9jcdx8mbAMtBh+SDcPbtVxlL94cnuARRLzYtl9qO2jQX2+hi/oVvwPWpG
z+ov9ICCp7s38SS/KdukrXfwHtll5eh/VL0lnjBqHd11jrJ59KCeTmllifkgKq8eX21FaK+F1EG3
3cTNx2PiAr1fgNqGvUY0Kj2D/n4hNgP8Kr7qlVxl0vgkfuh7dt3UbaUX8DLLh6i5PzSzgE/UU9oo
qHUflzdTZyu3+tdnuL2yVckUY+8RWRnI/LCDDI+vtnMTovzn1BEFXtvE1GD5rVBmzuR/xbmaDZHq
csYuWZjBpNGI7U4BPI8F+PCr7ZiPGfEKtMOFfmci0Zvktp6n1novzhOQgmXC0dsq4rAl5VZboiJC
2kKE5L+FxO6gTyEYWUFcmSxKRrghZUnnPnLBkaiIfGpzyTOape93s/oT1VMhWlU2KjGFWz3YcOW3
eRb77dk1xtqin8fnXth8+GlZOOPhaIVjuOipzvaFHzGfgYpZFolM0cOTX1U1Ihf9cAciJrE0ls6w
Pe4vykKklNFdeEv4p0mFWXPdCV/sB0KmoDrZyAGfLck5mAtx5fWvtDgoorqd0CO7hPhWtKGTIghn
luYTypC8MdAqyAL9qXRFheFEWtKEFikGhCCpOAB/pl/68sh31RdRTepEVlFm/ds6RGtNe52qO3vC
aU9oqTyMxhA11pQYJ9CpmmbNawxBLZ9eYpg/xv2WkTsl6vDxrLr6In2lZLTh3m0dXQ1eDGeZDpI2
4AMc5crQBsoTzf7eEHFM1ef8cI1UQdJmCHYrdZGoxVATM2c5NJ/FAMVGFVJPzfd0chmThjhPtU7l
UgMTURYqAiBhLRSez9pMPXdkVcLDV3MpN9oOrqCbsggc9Ae/uklkwrKWrEY+7P5hR67qGCj87q3D
/L+dqA3+yqnVfMFj/PMT5NqJx3ql+2bBQ2y/ZH6stxSCNkLbSamsPBvkxjpax+LUBkPU7ZwfoVIB
vvYhVhnV06PZn98WvdKUgoWxO4HOFTqcv8X3fnu9OYQ1M88WC7wOI3r+uxaJoO0rTYbhIqwbHom7
jty275G1vPLXjMzGRfyP9sgjpwQrGf28JxBomS2CHeTNCAOvVogb4P+vW6XL0uMqI13dsELg3PBd
j9GYqz1xkQmEv4/Zq5vTYWM9hNHy0esPc81ugtXnr8rtDb0TyoZz43F5gq2B0zSJBRykCDT5gtyM
9/t1UNvylGQMSaBHEGM7oxHMzVXAgUQmCKkos6KrVNsVmaG4qOace/+RRE3/5hNpR/+sR+nagYVr
PdyzLz2uoVwozZi9e2tP2kZBouHlPGx1j7urHrGZONjiYtpVeP4OiHN3u0V/ehEo0EgIAza8YuN4
3SonnmVgTUgV4KjJl6dqnTJ64VhZNjQ1AbobgbsuUvPUYtpD44guxw2/BXN0xKiOFl5/9wF3s3rJ
+1Avy7krNS9PiatvK/UlA20oksObFcNVv+SmFwj7K+80+QummNPlHnVhIbOUCR0YLSujS8yaHIE4
MtNSJ2k8HL1j/D+gix0XagJR18xE+6dJxeLNNBZFzeCRnMzd/SFFcgQl4rh5f7rovB1dhlSKPpCJ
tKkWQnYskikdU2NySuWjNgYCYhqsH83C4Rnz0trKjJg3pU9/vWUrUgVLWyFwEwJyNaqewwl2izdz
q7eq6IXPRQNGZyNki7ulxiaMMaVtGoi0Up4SIiOugXqLNSccJj26S2u+ofLbi9GatdmQnDDDdcXN
8AdZST/COhNbbe41S+nWXHEsQYpEFYipEI7//Xu6giC00kliiavRje1kKfFnN/hdtRlyrdcGBW13
XbkFLUdMXFP0ALyqV4GxfHKZSrL90gVuQW8N7/Cb2JTlijcwGSLHN8j1prl69y5R1W/N1UBWcNAm
iGXTaSCmHZKkhJULNEEPoDRRRMGMOX9bRLdfvZZY5p6+RRisPkVYYPEjMXyQKc7oh80ekoKKG5Sz
VUDCVP+TqGcZzUAx01pBWvCtL2hymriJV0V5nroGrU3LeQeGGN1pfOpVBRJPDMzDfidCUIK/tI6a
aySz3DcwasHYf0yj+aHOIwhqPwISiAH+2ToXx0ag3tgSM5qBgR+ef7N7OU565EQ3uJZJQ7e314PR
WunaBYC8pYTPoaWNdol/M3vkqdATwDwndJrJO2tPFILDqw2DsTFAD8xTileXXX/fMv29BnRHQlAC
65OOLhQPkZ8ORl9kc3/IXtNz5ulvQ5we+/MFy4vK42M76iSgwiJXmqVlOD1VuE6Jia/chF/Pw/2T
JtaixMu8U/fhtpY4J5nMWuvSupqo40Jz4ofk5vhm717zllJsSfRFFIE1Qu3dFX4wbUai/OZNlUzK
jkO71Qb93xDuMXvHd/u1PTOVBVUc/HgZtWCby6DNl3fPsKotkAY+0OcAyYvNQDIfupdFpP7y8To8
oq8LdPU3FljddhwTVty9rk2D0ScaNPDt/roipl9AWJ05pCiZwd/iDncD61FunqU0AOJ17Q8PGBEd
Qahvn5TeOtCPxVCQz07OruDXWTLuItvCC+phGU6wkjdPlg7unEGZAo6xZLMmumaY0zS896rNlPyJ
IaN4VuAlnuYFStdS89narCAvc9godHUH2lfei7+4jKFSV5r3IzqZBUNBYiYltJKIl6nxuo2AgsT7
k9f9Iu9uSW/9O1lL9yPG743157OGtWtcgRLknrqUejrpoVIlyVIDElU1P+sTX0RuwE2CAH11c2mJ
SR4VndcaF4Fvs7NcJ8wn4xeT0+VP2sOCbiohtwWq3uNhhwapIKly4eMphE2kwhv+pxgCpzlBmnO8
DtdRdkX8utpsRDyvx46n0AcJCzk6XwoQSvRB3x84jAWi3XG2xx77dlwurNtveNwCccfmUKcZGxpS
Zr3EWinBX9pO3KDtEqqS2JSKv3tYDP/bytPyHkyzgf59HaVhnc+keu0IScwbD9v7Y8wvg57jGIuX
1lewb3hBrq3Zn5PuOb66fHZg2CnCHnhPcwTgf88/owESAx2Sgpex2EcBxcmz6P0vU8rrtZ6IQ71A
nRxx3+QIIeLczk2oWrjNdm5g3hO70X7tHLdAdaccGUF0JnJyWKMImdpON/pdXOyTcmgpt77Q7ofb
1jKD0KqY4BkRT98CetTZZaZUntDt+C4HbKE5Y1kWHsOotJHVoj94XsT9FJZqv5OyM3cmEL1kaQNF
oK0QegXChpgS9ftjBRQzAMHo93Ukv97bx0HoXKNyMIZk8xPfLF8JuRoDJTVkDcMh8LPLMttfRE2p
egQ/ybUbeX4eInNpJ+4vDA7rLHkAowsYJ+oaH4gjNKPKtk+fdUAkcn4jZDTqGPEqGEHEU6qo4IQa
mne6qt0kFyp+K8S35ID8L9DITocb7KrbuLLcp8mUYsekBHvB0DZsEFvgkBYWASW6hAIR/9vL1CDY
vAIeauBn4DxURkjtYA9yH9vAExgHw5FQ9jYsfhCfChiB3LHW5+NGoINhxkCltJpkbuFhARPaPzRB
l7NXLX8irIxO6FkyfwxV7VAV+vmOCxMZMhEFc6Z0GToIpCp2CwjrYRlyhMAiFZEGjdg9Hlmvesff
C94CENtKCn1VF9Yqxsuhmm8qz0wEVARAivzEJI+rvK20ox4v/4zT992J1nY+XhtSMOZGtyPwq+lm
A4lu22ryZhI+CKPoeXjqZYVFFBoTzHNJpfarDd3LreGGczMVrWLeTg+nuGBsyuOlzFi4U5PLmZGt
M18KseV6oecjiGTidDVG5U1IxOcvzlg0YzJRAP3/h5GaqPQoUIvtyYyKAGp52GXygUhXC7TZpM07
UIyQ3WGTvvbA/pE0iLTFDmbWvJSDZeye/d6yi/xzrncPy0OuHFzMTCvszydcLwnXKCtfg8pFsK0T
rZyb9iCEECJqUStoIqVQKssQYemzAlS3FkpSjp148ggexcXwwIKiaKMuYJP7Si0q3woIBQXZxvIh
6w5FKc+2iTC+a8Sy87ypJvzjX5N3JrTqnCRc8MTHrIS/Jx7O4gTzPZMal4ri9t/z3nqvX4uG1DPO
vDVyDo22YMOYTmRXexT8Ds4gXL75i0ZCVvZYzBXtd7d+8pQHl4EabjMefuCxKaauPGosBtdjW5pj
djTqkJYqbPK+1uuqktrxCwy0NBp3PTMm1MgTlY0za2xpQ0Ge1G8V+Db53QGMey2q6A6MtaSw5xdq
KY5zU9WMgWFrsZxfA2ZQXosF2CrkERKQ91FG0xQIk/NZ926ykq3VHZTrXfjKxIibPyHGCqzK1J0Y
7e6Eb4kNNi5COY1dffrl8KcYJ/7NYCQXyoZD9tDGpj1+wZFiHaztu5XDZVI6Q7HqqJCpGG56QfUD
SDEnAkGgBgt62jIbaY+B3Z7JFHYWVXsLRol56gmBB+cQlJsuWe0W6HTxxflVz2mb6sE5Wskywld8
U1P8NZ3vz7QowSGFeVu3sQkiETl2XelAlMQmdYNDKHlaydmvdGIqCkloBO6CjyUi2j/zDpz2qYFN
0Yb35BEx8Q23jUUXQSDh1QRvKnbNKYaBTz4goMRFxixLcz8wTaubjfbWrUwoyewfWqzgjarxuYtm
/62jYrZhetNd2HVcWthG+HNswGSAA1B7S1DSyrY6OXLBWLzltlO6qr9w8kqApTUPi6TgOz1s8F9q
M+ERgElfW9eA+agLra8QulYCBqzqjonnJ+wl/PAtqQPKBTtZ4CwUs0jYVoCOYUD30+DP9/j6P+lj
FslLVFAKEOqdmTm3orXJOqv/iEti66sajkzRCC1qmKJ7E2zY7S0zvyI2taeCSHtPbaBrrrIxRFvA
xWC3TYltIVXOdzSefY5y+FOxXU/oPE9+WtirHCCDIKvzism6vqE/OWdT2wK3YiVb4xwWy7tselVK
VVveDz3Al8oCPQ98eJcj2NMVLJzl5STX6IFjRdGq8qPwHumQpOPbhKi9elyUWQBEAf3QZZcKYqUm
QMVKpsIvZLNAg2SyT4UUTLSQjINqWehi+rtjXtI/dmNqXql9KNS8asVn0hzE+HGwGhFDAhK6kzXx
2gsNsxaW4Vf80yg4DQXPX3Zfkt/MBoZ8gWxAzH1wSAM0clRXRN8t4xF+QPzFJllcrTD2E7oIXSXD
uuLk3o3V7jIHeHWyfCwiEBGvlJk0w7hpWYSuYpQMVvQpYm/RRW33y++ZgPNj7nn9tK1+BVfTE7uD
RjUA+VWdU1/wF1V6HN0ZzrQFJBi0C4K055XBYsain/nifqL6mnlTKtcV8Qx17o9dkErHtHINYlbo
u19wonal3cjxW4vZJqFxxJwQ+gGjFreQ4Z4OC206swgLxGB3m/6WXQBZQmmiMV6uxv4FPaS82rUu
nhYSws2hMNpo9OAVs14c9kLivBm0eh6OfLK4x8Vha/shoyVAxuJ1InzGwCQFDpOXrFeyPgvd/TcF
LxwyAgV8s4P6zwGm2m5DW4FZCIAOqle3GUsrYLp6SQiPbuNKtdpdlBT29Iv7RXBVf9+wnbQnYY3/
VYInDR/2UqrYGJ/4qHDLHQbLRYN07Qk1JA+N9YM5PWiIkl+ZpQOj8I6AqW0pOwwK2VZ/kZA+0Q6A
XbtNBNy/a+5XHnSDy3bmQ7Qve4meQyUAbJRUftW5xjbpx2s56/q9lgn1S5p2mstfpEzbrUZ5FnvC
MWrSA9dLaPw6sduCg81hkHyuQGGch49RiynsUl3zactKQb9hJQpVmiaWT8JGeWWFJs8jFKfk5fnM
q76tHxCeVI2DIhz3ejbD7HQjoWN4dTCWsCkrAc9d7lo1QlP4KKUyJEbtvj+mMmHuuW/QjNs1hQ4m
1QZjqpscpZDZLhcPJL2qQ5ipAW86wTeSmJuwD4J4BJGdTmrgs5nZr3QzJ5VZ1yeE1Oxe8m7uZAoP
7Z+r8y26sNEHMz0DqDiIz/EgxtkUCX+0Lq44iprtsKHGbn87shZ9WKlXOiwUMwIsf/gR+b5zXHQb
6xMNFraL3bI8LUUO74IJvKM2eaAr206PMvZG0y24gSLBy9YPH8sypF7Qk1TlzLk5zZygoFPVocxn
YXdRkoFS88TYM+dkF6aUa4rWqw3RgsmAjCJFS/XPDgJTwZKUSQv5LEjosmrliPsAb8PPBFRFYNAz
3n5CaEyf104eiG5XI3R6eX6grb8ZPsj9//Iv+CLJrS0k6qqPKRUtAw2xeJcBpLoRtg4/6WKkaUrF
p+64gT2m+PWZkNrG0TaJSIS0XMwWYYHMKG0O6nNbIIRml3OuJrCAOZJJqmzcsVMJ22WsIlwANkqt
6zz+dNExSqlSsh0W1RTi7FYKS9/hgtbRRfh5vdNAhzIQAKvt4741PAamH18Fl0D0UwpSXOuw1rYv
dnno4ZxVVQhSiv36xINjrt9wj1GaxLDlW6CnYgqsGQAN4OYaKCaGUMIiYwwQwYXHRPNroITR1/Z8
es73rDcKu3GkTGXNOPexn6np2kRnlLkqUxOCw4FwMSO74BeW30UpRJfZr/Xf9EG9ObPx6CdFVbE6
s7dxpzfLP/ywPPxHBpgl6AVkujVhDjZjEqWMN32KJSV7IYIRXj+D5uLhP5xMVxkQV7DhY4u+8CSA
pwb1fyA4WzIiPdlorhJAS2S65me1DjhgJVoA3FzwcexgTZh0DiNrvwUL1EZ6YAyG223T+DJZX5Rz
PuI9ALxar2Jterse8btCV8UGnNklLu/ENDwOXBbBH8Rp9/2ZUBQ/EIZ3jfsMp5KsgZZX8dtxsH74
msFXvmBWF9ez1nNRvi1jdeIUyDznmVCn4c1SUXBirL7tVOg8KN9su0DWLid2RGEVALFFqR4UAdL6
bnAZJjVRtJuoj3xHQxsjP2n5FjifyynV4ZX5wVPkZy9IP0y6kEbIcwxridkVyzv94qDAohF50hnL
1RDpu03vA7dpfoECT9RjCc0mfBSENvvTKd+53st6A7jfBp4W6EjQcw0AJw3ypaWCTW1pIus8EYvk
qNenCzAk6H9QcGLr/vvN+nYbrol0Lry4th8LTR28D7zyb/EBNAFjFIfubiAA39T591nw6PpcObhN
MAdQMfvNUuTxNJCnC38Fq7E2kPVve+O9XLzT8YobNO5KT2o0a1oe/PowFUwGsp03qfqcByf4U7t1
Jyj57JLNin0tfXSQaC/6kmkTwS5q1o/virNIyvJHb3m/Mv8tIX+p5360KhNff7rIj0KxRi3Hf+ZN
2pNnpZkb4fvuxJ2sMktEqmB+Qnbt9bGqksDqMROBs0RLbB2w9Lvoiy/q5VghLOpUKsleDM/YfKAr
idZq6WdledTrRN1JHR5by7bX2zJBqfpUGwFucc5l7Wd1dDmVxbf7fDLHpTVavZ1exv2+rCGfSNKL
iG331Q8f4Fk/xHDcFipmwwGfnD3cREwBu5DE9M0PJKWrp1Xt7iAfOdX4z8B1Gt41nj+CCOrdZRVW
zw1OdivpC7Yb2MW7TwKA4N3CQ05N5LWFYy2Dcuf0dlVoD9Y6/sQFRWCLPFAsbcbqcEwvZgzzX+uR
2UoWkC4uq62bYfz5WepiyBwuPid1DMz8b0tEbNIS7oo1n/sMe5Yp4WPJZW3zFjGacBsrJHU42xy+
BagSOqMtcCUf/zvPF6xy/LLcSqYDGtd97Sx/vrPYLrapOBgrRbSHEMizfTPNXt2ccR2SqRwaF8EG
Imy1SUciyxU47pX+p9Q+bk6gQ3iflZEIRId+vlCn86QxudZZMQstXJEjvAN8CsO91qzxZryslNAF
ToraxC9rDKLYIjIi0ZvtuRNL1aPKFS0UMT0gwe0bKrvuX3HB7nkv6agcfY3fcLt/7AIpg12HLxw2
/aitVdXjGVT8o/rw6K4QRNbZ4ILCxqxThi1pl8WlamrybZXziW1vhZtOCvNHMDBl3l41aKHFIAm4
A7AMsVLxBdG7sVD2gP5EUKHVBW/+iMzhdFG8Zys5gznJc4qwAkidMKl7/xlqlJKTN73crnD0ADoc
Zk0jMsiu3ft0/WNQjV/w30y7xbL0x1K9dbL90m27v94DJlvc5zGfvJ3YQR+Jt7V60zSuBFC84yYD
JSIJZ5JP9DlBLuthcMCycrRDw1uqf6eZo80Zy9twbecj0cUufQlbXRK3gUpA0rMNz8l2PfFutzOM
0s4XD7AJP9ZcH1xs/HovdTxPoRf1qzPAJw8g5ueNIQZxlZNV8Bif2a1EhBrKELe2PZ8KTWkSHGwH
aRHGTZwyADAvnGe68BUpvLlw2kmRwAwBktb157jdsedUlQ8rxfKKH+yMk3s6GGWbPZAhrmZac9vz
VeWrZ+xEHkcb2BnNavDMjV9QrLsK/nTLRNXMMWqnMukr5ehPTKTY3+egsKN4bSfteX4k/t4e1Uev
C2U1XTqMd3bGnIhT5vdstrr3JkvVduq+QKrnVZ7szP4BsNhaEgZ6+7bdyQVECfnlTjnsKU9aUNIY
mqwkqkmPj7K3q0uuW0gvfClWt9m4xGffInqFsbOpZcMqh1hu6jIHLj0ttjqLr6dWu1B0mz8MqOLD
JIw+43Y1c9MMLuVbjqakJWjQJntT6PFuWfp6waHrHXAVy8A1hyjmpPLPlv4TWRYwfCDDBIM734C+
HjaRDgqxfAWasxtoxfLR7LTqhvTqYDUu6sCnXMCCmwzUs2yPGeOtA7INE9E6EFINCBKYPx3yKHs2
KzeJPt8qM9Y+XdPSdPOiaPa9Zukpl1ktYhAwGBwykUvC23W1omVLDemehbCFk+n1UKZxlADByLUX
ju8czFz0iUpR6gfOGp+aOwgQtctdbn4P3VhWFKD+jD15l81ZYeucximt8F3MiQSG92OQAnp/foK1
F95RXKJrXQ+wf1LKSGgMHccaO6swsco5NtMQW6F3xI80wYL0dtzfIqKuiqCQ9PBleTs8dc0s3S3Q
la+nIJSgeC36boZ0KqT7TQz54fJ1dBEn7OHC28ZOsBxisAyCKuM+LO8U338hrLVJVMTpTBfxJjg2
pdizfFDsCVglnhKr3PiHeQhEXfajsEQCByjhqvNtwgcjg8Ruj2L36QCEVfmUMtwfCR/96b/svlj0
9PKh0T7aD+GEiZJHZNnmuEhA56wBm3EN2BKMqP1nGOyPd+kzZ7hWUb9inDRpyST6hjKlcHhhrWE2
lF/csayEvIr39dPeGgb3n+pOmLadq4erQuItyb2w9yoy0mJJWmHTQv7DT6qT5i+WJQ5lW3nsxJjH
C5Z2tlim9x8aqEN7Ou+Rib+z1p3N9C5WTkNYGis6vVbGkEXHI+TzSAkHnhORvPpdnoFi2/MICrWc
Wz9IXjJ2bJxobzyppl23fo6upNAkTGw3UU8wg1MwNAlFvthXqpekSk8IFLaet/MtCwmevPzCY9tt
9JuYAJOlaODuUS+p8KcZO4HNFAg7+sXHdOgY8YgrVP8Je/Z0ySQ8QyU7k5NzjdBPAVsA77HYTB0+
Rt0/GQw0MXgx9TTaxbFqdaPFvsMJyyx23kgiIUANWd5xRo6pE9qEoKaxp3d2BIxuXjcmcGpatCCz
290hr4UzuQa9Xx8odfhDq/eiXGuZzJ0lnoRr9Gu82xlrK+cxsunAlbnrcErgG4tmq2UhW4jjbCnV
Lggz0TX6kYLESvStuct4Gi2UaEFaHeUBZJHXUm9Ec5IA2biS+PBjc2CipXdRvFZwm0Ra5RAo1hEI
H4aWBF3YVqWUCGCGYD8Nptv/s1CX4AXfTIBKfeAgcNuAO+9BTsLOQ+1SmdgJ+/7XMLdsDsrB8wQU
y1Pf+2xrDw/9GHKM1SVbAnCPJcpPh7PfQ37wZbZPwY7MDiTGgUIb0OSBm/SvuSS7XJStVRjg+Y3b
zfBTQXQjNYA2spyGbaiOTAEhCYkWc4y3WCY56V12XzYh1mwzehDRHL0pBi+UoOryiTxECS0DdVwY
VtilvRFda1JK4jMWlzZULwJJXdxwgfNyqe2r89lMzvNTieQ0dv6hduNGASyF5pjVR493ywXtKD08
+uy/7eeFkr1+0NBFuZck3e0R3SAKE5LFnPluI3MXFimfjFqBhSm87OVrSx2EiVTIic3LT1UsyaNA
vBWdN5CARoxrGG79/iYJ/F56rBL50bR5T2Y90dtmlC6oKJJngV6IFza9WHAg6OW0OcP33jbGYiBT
0rpni5slN0sccbqSVtNR303AGpJlH4g3V1wlTXvIO4mye9Z6yIDUyXsxLmb7wlB3pKECsorrNftG
dSjgC/c8SSXxka4d9vlIvnP7c9Mmi4+bdah7vZ/sot6Vc25QRBk97EbMX4uu87HLlT3cZ8nuqr/r
2ciknp/dKynjBp34SR44mpM+gc39M8I5YVcENUzAg1jJ663qlZx7yqrLrFH7jWei/PENt5zMXBbe
vBSj63YJu/tn8jBSXSQ8742hpNvdWA8CONIkA/AP1V58GEr03Eyk2kSY5RP5DoBqaYftCnEMnYhT
1eb2He/49t1GxWXkktm6fojYTwNqndXObQTfCiQ3LAJW8DCR00HWadx8QbfsxbU9HruY8lONzzW9
QM2QRGJxX4kveG6ARGVKAlXXvteNcK8x3HYWAL8VEm79JPR2qM3f8yrHIAqraBRzU57wbwjyvElv
HORL+h5iFCs77JpQnKxAUyIO8eE174+lYtRRt7f8fnKk6vEWcxf2pfoqrrNmy4yPVgnyBxhRvvT0
a3ZwobAMnfl4CKcdZgAQxKfTeBKYzoicT0JvYurLZkDjcgy++URTsdrNHC+jcnJTSUMt+E99egJd
r7LB2+oL/1ce43Ew+XqSjMyT3C0X3Y0rvTShsahKr1XDfcPmR+Af4B91K25mWR799ostnyNdTlZX
eF6Kas1RB0rdv09PVUQYhqAbkROJYbvlwSWqJ8NcJgJs1RZtXzoYqnZap46AOfACtMt1lDpLLLHt
9M5KhmBgF3mXw7l8F1U7pZ4JuNoklKKg+u0aowrtVHX+7D6D19qxXgRxhTSdnsFq6ei67ll5U5i7
LheycjCY1QcsyZginKGp2a54+YDS++WS6p+o8UBvYUnNVA7Xqhvz3L295NnL8VfEr2BZrRSUSP82
/RXmDMhr6foFWxl0L8Rx6iNx7+voFyoUBEGliTXtYtVzdcA9Fv2S/WALakMXZ6176X/ef5wZsA4+
23sdN90WH7Hk/M/L9nZhrK8/1jVAEL/H0/VpuvRzc/5YHIzcF1BrXeNbTSIj5AbJS7QhsVJOeBky
Jb3nB5Alssx4nLGQlAfNwo1xeyqWJjBeI9Lmk1b3/Ayos9PMTp97pYECxuF8Y3xishsPTcBdt9ax
CN2LzyU5F41YnA28FbPDXYKl7FvzlqApNIQrLgLtAGhDmFUMej2N6tvaTvbo+fiNv1ZGGGYL7lNt
AtmOgxtwBObXrTQ0Wvi5B2c02c+UHzdjRu+f7jbsM+D70bvGb43KTz7ZHCLAl2xV6p6k3Cq/sga9
u+z6Bcy1MD7/41lF5JQ9UZYbibbKby9ovQNv5lWGcCWEBZiPO+hqeiRBwMaIvnUB8zWZjONBKilT
xiPn3ls/bZuyj3HF3NIqEmpfq9oJy6/bYHIRold+2U+ucfFiW8Qp4h8T3KQKAtJtFcfd+1Iragyy
Ak/bAXTwpwSWg3OjTTRu6IbbVS494TxXAhjtp4epFvLzi4cthKTyMuhzGZLwZVd1bZd+cTpzEK1F
gzowyN+c52oOcGfRHLLSpQf5QmLPfT/W/uKk9OdHrDrDVIuprCZZV06BmmGOny/eNUhSCR99972J
eNkC1l+TE7kyab2JiOEcPieRKlaKh72eCOdXOpb/7wpjUCV0XDSBnP/f1SR7OQ6dfHE+oBehkYp5
92KaDbR+40e/R+Flf/AwlAxOaluWvMovGkjzU8KWdFmhdbGKUsJP1mQgwti45W229jPICydlWHwl
dhUfSDyXWfhtbsuBYmF7iVvF7Uk9o9xl7YUVASoMg+3nfV+2adrDBbfT/XJRed0Uwc/HzIRV92Fy
Ygs5R+8/Om+9WwOAxQ0ZPIW8MNJH1zXSwYo31zfYdQp/lizgiIRlvDK9D+8xDDKqX4hOOVvSTNwk
JxlLY0z8SmxMm2yaQuJGxrWG2Qfl0f5UsYgIW8vqHFP7weUs5Em2U6DWfmaNysbIF7W6/YS5sNkg
dhHb7aptEMDzBmoHkSMLG6E3Eepy6/bot8P1YtiFCvlJezu3tjtJFL5wXr/8XtnWkTgELiya6xOU
7Xo27aZ5yEM9Btd2jbX2LboM1J0IXtE89M5LmJh3phP6KuupjQ7sJ1NmC0eBz5IfUGdxcBech1OV
XW7Gvk8/gXIO7XiP3CsVqRFJtHmH7kOdOvpjNjlKFGqipuYSzFivJaB+EHk6VIXDssbV8CYt0jrA
+EoW8zfel2MfITEWVYhjdPewF+2MjA2Iu2TTwEc8MvdEJ2+VPYu748rpBj1Seu3U8LCN4m7cgNHC
dMuuqmab7BKeM5IWuFfZz5YfkI9dgtC3t6ybwi2wPy5I4ImFCCd6VOCxwjLl2kCz8vmwO3UtK0Ra
DZVN4mMIoOh31S+7Hfx7YjUS7UCTEHGF8lQOefyjynqNU2wgMlHbQbqLwUhXq14GYRnmUnnlwK8I
lyHh2weXNGAjXZZJW89ZqP2F8/coS9+/qBWFPKwu2DPtRh9D2ZnAO+Zv65C+H5GR3zF67YUt+bCu
zhYj8Mg22U/YK7qgqb0a4XPLWHhkJgcA/QjcCQll++jmbFwUWqoIT4aCKO94XKgOKZxWRcvxclM1
v7/PUuzvzEXuM+QHTV7hMFdwT1L/8ykIqqj5UaiOmwXsrFA1NjpATV7CeODjCBhQlMp3O/LSL/cD
ClYcWbuXYsqrXrABc8BJTuHykUJKpGtucdm2VQKdxPRkjUd59j+UNRR1BiI5Vt/arp5LqtwxPlZ1
13BMLCRXTxOx2MkPzD9qYHo5zFJabGZPd7rbsSHjCloefz8d/4gXTiYEGXofeWq8K0YsAdIGzGCa
ua9W/8bQszuNL62byWLTDFOyrK7ZA6N/C2zVxyBMbqg81oqpioirReC5HIlz1n0wjNIEGhch2iLD
IL5AkUHdnr8fxSMzLw5uUYC39D/fUp1DKNWxEp5rF6iuckkiuzcRdWu6m3cIytFjsguWM+R95Q5+
5gziN+Juk/Y1yy6etMumrg1JtK15pNhVre6JPVwmu0qs4HB+B35D2HZzeU1z5uT89Dh/UxwIQJmC
bTg8xGSh0BVhmsmCPdk0ej3hMEdWfJZ/OdsXYH8z29hkup3a/Pde27v8tGaQ3MBGwREyQkQT2o+q
uJ23qdXEWE+yhse0zDkWG5d06ufsxfSBTH+vTeNLGOYvMj3UWXiqjV96SuhfvOfI5pQIDCFjKKpF
LiFvEXmtjG+Sil/A32UokCpiig5MsRfV+VYWQwFskvAZbRQxQDbDPicI0x0e1PNTelvy82LiYwvW
QoEdK6Nu57yOOZ0QPc8ARlDh1HldhqUacjgG0yiIpqX+0IMMzhBhsDn4sj2LTdCfxIzqccxesiNO
dR1gZAQsfVUWt9N5Dp/TeRaB0RCmKaxaQxpt80m+QOnZurx/jaLHSCgCvqVthwaLHq3a5CMhyFiC
SoJ31fNFlAGZGmKP8NWqmeC8COoZxVoBVQZENznUjrzC5XhX6Qbh212bwCC8u+PtXS36JmuO2inx
j5NV5nymANAssiqwdwDravEO9tIoDU0JSTBJft/mmpbBqRpeRAT8mpxRdL2LWwDDL4tjEK65n7ga
GsOsbNoGjPYhTJSupQzUwUaRCSjKm7ZMi4GiTMoNQ6tVYtlmjo1rGpkih9J3NpB/yotWp1PeTwfx
R6uxS0Pq13OPWqn5iIs37Hl8YAhMPT5XiILC7SVthlnQ+1naqWGpuC5uhbCtgbRnRg8WDs6QtOaF
Q3F790hIHLzUVr4ekE2xXhUa6eK/Ns7BrTjR2TSb+xoHC5pYPsXmDkDcc1M3h7nTE+SNjuYJs53d
+qNZ0cWOv5ebaXQLiVSz38rmU96tpjlakIO30b4A+/MqbSNAIxAyTVSET3dfVlb5aN3YWq84cg9x
5qCeeZCJ5vrYTW2gS9SKyDtOKjBs3bbUfFX9XrzhiMppbOE2Pw+kwdGfSqTjbU9immVbaUuO6zT+
/a1IPl93IpsZIDXL+0AnllzepfRlwyJpx0l0qMA/vE5U0+00tbhz3IjlntYpkRyBSCHJLz4dfyEJ
IfDskruDYy6EWYSiC2tBA9LMiGRGifk96vmiibzy1WzbycERQ/oXXKbbNvt/aU30ws+1oeCFHrRU
5mSMoUxIkchQkm0ogPte4B+9F7APJ2uy1yatvIVO3YNT3H3rUh4DwRDcOVf+025UcCT8LsPJiDg1
B6gVY3nS8XbMU8NdnjG3fL9HpCS7LUEmt4Svua7efk68jV4ExMPjBeMRmSXZZO88uQjKLfSU9hDz
Ht7MF3Ybb9PjTZVAz/5pCj5FYMq3uW+GiA2cgR7zX8sqp4iClCyQy/pCqNtdLu2KnbvEe+5AwIzu
cfvW14b2N3VTpQklPtMtWVe6OexqsGzhuLs4T3HDtjiVvyJmLkjeXSLUNgSzaQL8CfCgKCPIVfim
KHtBsJ+uYou9J0DYDj+z+7G9JUyqmL3XfjzUxsws4/mBs5ODd0U2u1n29CmuN+c1qvmI4eY96U4v
3mtCIBurrMNWafeQX7ZhRBOCEorYaEHGVQshFiuZ8cFxJdwcUsFV7RlRtdv26h6ZgGw+lAUGgxXB
DRps+KmAnFaHnOokEHsBOF2B9IgutKp0Myqw5TT2avji0ErIZmwwhMuvU2OfeTHQQa0s3w9E7uo4
OMCtTbO3aRlrrrO66LSa69bTScY+warFWI7fAX90IPgdoCAiEFEIzLbUhzqfjZ5imypavD4UrJS/
Z+NUexK6v2nASkkfOfznjsWyam8Zh4Vs8AQWAuoJfTwvDVM0I1+Hk6vqgctFd+5Yl/YJ07+KgJsV
XuE+GR6E/Zvl55Fno3Bpn3S/vtCgIqGf4LhjZt+1OPYBQ3ocuvuZ5faFr7sjO54JBJN06Xs/dBw3
CzoXKIiYTe7Kos6N8cGQuZM9JmUi9mCKJnduZI6sUgTKjsfwuBKpTBgQ3zztwSc/Cm9OBGKSeyum
NreSSzGwt5QFeoR7rYEo1cfGIbqsR3/teMWmV77kX4cE8bQrxsic6+nQmazrjSuIbdETWYaA7re4
/6XujJm72JW2kx3ziO4BlDJixRDPsLLghxyoUKXWps2pBopt3zX3YOuWoH4iHHqPgDe//+NVXOFr
22G3wEIB2uo4sxsFoeeBQyVQcgOUwm7L44t/97tPt0PZqHv8htSPFhm5OSQmEHwiUip9lz2CYm0r
HdvX5Kvt5IU9SfJrSEmCjoR1tqHG/10sEJDrdzsRfBI0OlC34j0RpdGb/upjp5CRcBtFlOanYS++
gD3xAK7oGslk740E+WjF6BW6OzSgjp36iB/uW6WlHAmr37bIV5+VevHtZDjoa3aJ7UYYK/4L9wAy
MeTlWPP29Ep6oi4uB8dgmHvW0i/vrjAynA3dnQL9QcSV/siEA0mIuIg2BWHURfZ6C9fs1J6Jm5o+
mYcWg1ikPIl5Cb6J8wkUiUjwOhGUOpAj26c9kLReXzi9EDA4iwCn+wAQ37qPD2i0a03IMAy2IKGT
5iLhoqEJyDajOsg7+wW1sqjtMC44Aq6pDVjtvBHSYLgCyUZaQs53Z+1thL5qmmu4tssZxkQg+58X
MTrP2WY/0KiHjfFKtFy/3VEqbkGhanKT8pn8uvenE7ukcR9bDCd6qherhcsXDzk0yqCc/pD1wGi+
XFGUD9Dg7yCLnktXUjTlXOUPUWraMmwfZgzDPxWWcJYl1QldfFTVPXK6MhZGJvxQWp1hCcdeFzYw
zaZZiWqZ42m6XjFNe4A1o/S1JkbcHsx82abvmrQWdBUAZtUiRrgROCYFudjbn12iA4hVbBVswcCr
H3Cs3luG/meLcwtRt+rMDt1wYnXvlP8qUpKHNQXmggdif49E22KhZH2zOdDO+ePYfFRyPRhl5Dn4
onmkuUaP4aeKnFs5ujNaR0q3AN+s3+ER+fED5wtfXY/kxSfWIb8Kojz7DP+I/lrjR/zBKy7NvgDy
a1e/LQnepfmrWP/y4H1dxu9hblmkzbXAB08RR3nTCZPd9YySQ315ZIqOzNgaviJvvwCwMZ90Kk7z
O24KsN0s5Y1SPoWhcQijRYrzzVF+v1UhLuyIX3qLZ6vfUosXsF3FWIY41MMpuMyQox2FtaZpJJM1
tWCuWJQrSsPokTA3aO+priCNQIVwBT2aeHbv6Crxt1wXq69Aqu/3ltkf3TdauMtFH+ybD0c1XnKl
1TO/w9QBq7yteWJ26UwDjCUwAevbhX03pycIjxmq4S1SRD0PE3ktXnxr9/tyfB0Z4nfmqCJtEaGN
OemaAtKC2N7DCdIw8UyiDj/MG/4wRv7D+ZkAJcE+HVWW/0JTfRO69VD1rALDDxBoi8vYUyolJR3T
BzdSlHr9IaQ0fJrzQ+zA12HgBrtGZQieOpNs/BXB0RBKpB+NkdbBoS59WcUflmsw/EkMnVdenWRw
TFbsYpf4lBh7b2UIugVfFLCQikgbRUwnZIPE7VbmPQWI/eivKS5Wh+E9+XHYV5/c6qrRNqDEqhky
/34rxr2QBaL9ewa3tBGfvXxsmrSh4vmTDRAi+b2rPWY5/h2ep2RU51MfeyksiiM2cXbPSQlv8aHZ
FRgYhEcAg9XkLo2t5V8yDsiykV4mR7sP9uxP6We43c58DtigSx2rbxZBAYqd4OjFYDm7QV0JHpGq
nceNs3y2nI+8sJrbE/BSxKr03ikDIS++KH/uH3R06UNMam4RF89Tw5KyCVSYljgvm2Cf4Y/yLNXe
QrIfedZm9eoN70qHDgjJC133Udqt/y/1u9uXd/sRW/lrYo/iTyq/zNGAte8cQZAlfZ1Q9RP3D79Z
oiQ421cxxRAUmbBWCVdt09kehX7yAzqmgkUdayKX35EqmzOyLK1wwspZ2tlQn1YrZ/zZPGNBR+4B
2jVvA0RgTdjsMjpH4tCNNJJ4PY4ofZYK95EOMPtLhLL6YaFuFm6UkA6qr5FJpLRpCwZhFr7yiI48
SPeDOAWZ2e/l9Wz8Roq25iGHo8udWZfIJw3mZCKPKb58RbyoQir22F1OgeNkk0ptgtUzp2zlLkfN
NsBoXPfL2DAaY175WYk0FnoyPJjHCqesshz9CGwtsNajd+/cJ8JDyl5pWhvFidNRzYv5/xDXNcHa
TB8TYcKqNh+pYPESzWBc9DoYKNV40mzIPWOFpoA01uEmQJ3qF5wX7+hktXeO3u4qVCP9JalTtt8l
MiBK+i4h4MdPCp3lDAWYVH6t34tkcDkWO/yBCJ6kuB1hVxdO981J0whbJAYny2eiO9F30dE1R8iO
rM2hwITd8CmRDFA4r4NKctd6HynCmrU6Lytw+uGIGYZ8A97oG6H3W9CgtJfINksrIN6X1T9oJqwu
GF2UncVhA6Zv0J6qMPfhosEtZnEo0/dLfsHkyxitwTVdh5CJOXP9EMypc31L7PWedHuhFICxoGze
Dqw/AinVYMWmaO5Eb1pEm1acdp6uxKrs8+HaKpCqFsWmlPlv40n/zHYgXrkyaeUAup0LxX8O/soF
dXiHFJbN9asjme1E44w3IZjBVpbQZqkLA0nAC3YBABxiNJXOTZx0b3wvChoS3TaauISuHk21mZ1M
fj8ZsOFDtWRZoEIr9IT+SS6bZ9xdhdz48khQsXFcqrYyBkQMismS67eWoO0G6fvVF2dYCOCXzzTh
ABKzp+cI61Nv+pSI7usU7xxe5bGI7h1XD8sYyWOYBdKzsvbarsrSkHE/EoQA4l/X7X3oDWra/JCf
SE2nrNSq1HzdppD9l7TbpzX58khBQY6oKl85IzH4EFbbFHF7hQBMm3ygiuORQ7jlAATye9/0eJF3
hPKdl4mLPSRLgAUb0oTsK9qS8juh6dcNLZSUGEba+1zsdS1VgZPi7Sx1OjgtBZXXp0yOyLOLlnRA
FNYMdSeMwRR4FhfRsmDE+2NHfdxvySBLkKxNfsBisaMZHWGusxJ4P9+JyoDtdb3HX4rPBuuMawPL
cu8K807C0CpLBhqI6XcDET6TquXKmfZvsjYH0DsA7N0pxwvObiYc9WDLZlTXvhPLVovKim8BKNDJ
HEgnx9vGL/i1TlJoOubSN3vioPD/W4ze9+YHTR16dvmWGVfvp4LyqCym2JdPE+VJiMTAbNPVCjpG
L20aOiR4f0rXCUtwvrf9Ep48ZSYCVYAMZKJKXyo+QCBbiur2HSbrpMYxD20fPVRnus5GIxNQWNd1
2HKDv5hhm/wA4QekyqGy7Pc+VpBFdS3rJ+cFE1Mksstevm6hIAzA/R5vMhNkyd/hVRwHQruGknOk
X/TLfGF0Hs4EhEuntlrXTq2Wna94wl/kFCu8v2IYDa6vux3+zghG1sOhATqkLwtQgeFt2YhLhuy5
vs5CQEf2Wh9va0YYDHOQKrLI8pQERih1bEN0UOmHc5hyrc97xtUbUDaaZOvLuPPLIH9K4qMIKCc1
mfkvbhfRKw0sLhuRPVuYVjTh/QQql9HhMizk3iwjHNU2WofjWzpXUWqnnrD9cHeqh2MN2U/ikyhH
/j5qKAiA7/4DOlrx/qatbofEKdR57UcJgvSBFrqxvAnZlqdAwMp6l4tEjH7vj/RVlSDg1SaBEaXf
3V/ur2tEtj6JykRlIPPu08yOf6hbEFDqe4l4VupQILOvXCiIuYYVH3p4dINkPmnNy1NSCnYaRk1D
YHGyZFA6lw7KDm6jcCpFM0u58QaUS36g1L8meruWmSI0jy2Bs9AfBGKY0IAZElcujHEjavRRXY3i
rK1RSXaQiB74lDlGvez1LbhCBVMHDszkEX9vS70KUXpctXfuIvq+qWX1IxLNiq9dXowgBCquMGe0
CWcWF4c+Oc8o0Hu+QEdCpMEzZJRDwlSuhYAR49QEdWXV9gLMhD2rgVhNuEvXy3Pbd9y30ZQCcXuJ
basMU2BrJP5Aez4y5H6xxvPYhMctlbgTSMoLtomxBOIHb4oI5AcLHhD5GrTaNczosBb/AR1+cGOX
kymruG1yGhTVCStJmWYyWQBKOrbmRFnKGdsDSB1pWpl7Bn00VXv1t4hOMDXFeaRinDq8dfU1Vdee
e7FM1ztFGcL1SRn/kBg4HIam16Pjum917eR/fox2XczoVwlPOfmfMFjUY9H5hLtfbws18SDoVv+0
BL5KJYeExZ8PTT/0FFs6s9getM3xfzZE70YnW4bXgnPwee5oWYKffTwTngUA5Mrno/ok7NLg33XQ
1z8xDY0uNGxdIas4u8fQG8vU1odlXrE9I2cix5t4j2eYDA4DlW3Q1q1wTngQfhFl+PX8Z5x5r+vx
yMqVaGl4zFupW9xdv8tuRZwgDnoPrrsEQWhIWQxzIapSD5OxCidd2dJxN1t/C0ac9lRGkSs2j5Tr
tu9H6DJzobEBEwOjTsONBRl09nlbt9hH53klE11TOOn9YKIEcq/S9PaX5svhl1FTNg3G3W4wbg47
XsTWbRgbdWc0bNwm0eNhL3q/03empWT/wirNnC8ngScThYt9ataXqjwNbkGAZ8cMlo5RIBYH9kT9
YDC1ZpkgG+LA7LNs7ql/icvpl+Q/Q6ca6oUZQzgGCX7gTg9apcFhsM1pYGE7k7KXijrz2Y+UbN5C
FK0qxlyQrW9eW7JTfxoQldqO/vGqfV1Rc9vZyRFx4El/ygoruStSaPqFwJi6FVCDTST40fVf5l7U
dtKn3TLvPzCSzpiW2vz2hD0erJw4fKGtjqwJQENktSxhfiu0CtBCDceyS7xhDxPLobS76CLMVRYl
QdbpWAWBjnSDIYdg/yODuZ2V9eVHYs0TR2DtOPqOfA+nwFrKFDF12wus+mbbCLctRNdsYv4G+VA2
2baYLzI+y0Wu9cAkVux2CNGy1QaMKrZSLkTN3oHm2C+Ds+zFERT1B5dfYf5svf9aHGQBpvvy8jyR
AN55apZ3dqy8Y94cP/gZqqfs9DrryNTwNMeE5MXCOzt6xNbZO8khud8MDvFaPYKyyana/Qn/cuL4
/sMhBSEVYW71C54USWpzNlgOiieUz/DDRIB7rIB+mDAB3z7jpwC8o1Uu9HQqJiCLDdvAtzATKn7n
zezZlaXrId7f/6mHuI2DSIcwp6KXbZt0t+Qw8VPXaXcflgeBou8E0POBL/2oJPymUG0UQzyR4ipo
7rL0U1LJfg37VU01s7U8fmvy1sHV2sJgHOq91tKsMXBOj6J3kXL0uX+G43oKVQD+UG7pb3kZQvof
taEm/gvFFdZ3pbr3uMg+hFEEyY3QK2t0Ynx9xDUWkMoI6sXET/zHcy663L7olp9eV2FfNvDWkrTZ
utF9HyDhUKW7YczkSJPjKZF8G30YhHNS4Ny7t5GuR5sxcnEi2lGF4WTwEg9rURYbJIQm3vLWwnvZ
bzK0720ljYCjKOd3CPKswFsRLt8tHvgHVgcFsMO29HdvYlyCbKd0v5PpUwPXif+IIl2X+2tERQkf
r+AgPj7XI3P/+wqEuFQwhxHLEYf0UugnSCIaDfaCuCY1f/HSeNgCSmP4HAHOWDCyWR3GcyVkPzfZ
rH/AJ9/7VCszELE7ZBtW8/anAhMNlmMguCffU8fw+EucNLYdH1Gn87s8KKEdBhRm2Y08OTKagHSN
foX56BfoCRyP5EPoJn5YAH8/zp106C8MVHbMMQrLhbmazNVvvjSUWVjQse/UpHd+7guqts1ej45l
QHZHGQ2O445mzILAQDy4liqCsZv51bYXLErr42gnhh4Dt4gLZ4of7mLCdNZErEZ1jZOFUyOTDde1
Csq9rpJdiS8Gxz5bjjk4jnFWkrEeKe5ALpo7qBbk/5/65Tzvi29XBf4JcARRtZuXqHGnz1JFvmbI
6OMXqFLtLB1vpWnVhHbudUth344xRWBFQ7eQgPHr8yEpZvajGds+gIdgUgmwskm8oOQ/PT+Qjeyu
x2P3/ph/K+sv0j+USkvNS/JKneVSb3e7sWyg4HzmPxFBfcqmi3iFCrbBLFTDinA/zVi7/O3MCpm4
z5p7Ry8DN3l/DEw65ml6i/9TJM7dEJZI1ClrMUGsTGXcIMbiTiWnh2PpPg6mB6xJFN1xEuwu5t/c
3Uc8qQgi/4imh9Qg58F2r5qlkbZCeLrKBUdLecnyMVlMbnoB+INhWqF0a/V4VmlO+85ILK7Elulb
OtfQ/g9+2RVf5YqNjdA2DU4CN9YR69Jf+/Un/hLkhzQgDDyiLwnPj7AJZFlnIibkcIOUYzuPIFDl
oEbhCDgNVzv6SIgHBgzEcHgaJUOHci6wW03IYZcA3Y4DCBbjsdU3ZPqhR9mmXYY1KaujNSAZaO2h
01/B3fWJQl3GCmY7czvv8PH9YTaTeIJ0+9CENCfz8lFz71RMxPjLXBDml+V8dSoV11maqj90OsFU
guz+oOKdZmBBx7Tl2Nk8QOs97WGbOkRkbeDH4CHdunTbcWpGFxr11+VDtuUk3XsW9PPJzSoBVoTT
iJRZ9my8mPeSftwKNE85wHWldG1Tumo7dkKYgB4T3puofwRZOZ8ui6xm3S1VhZn+f9T9kXS4VdgL
9k8MYKGhBpTtZNtjf3tgqsY06D6h0woAL9ZEzBW+P6lpjdBMfk5eokHF3yTY1Z65EbFfJxlYpe4l
QsMLF0R6Uw4Qtr19XwXkpd7UJOdZFFTm59W33fQdlARXMkuzMYAt1sKTwVQKHDEPkZApnmOJ5WSG
2ReUbAXW/OVhadHDqm18NQFizEHFiutzThOzCo/oua4cws4Ryy0h+L+ryQUflCSnqk6n7CvnH0Po
I8a/vWry82/yKU323oA72pyI5/UOGe2W7EaX0+H/Fwr01qBe7tH/mAA1aYLm/SrfBqYH4c+XWdTg
5A+eghn0/yyXOzH6wSo86QKTNzCMvOAlD6oF95rbYmY9nfVgyHn0jT+YgmTLKbN/Y4T0PEG5uCVf
opk4NUZ9+lYK+TO5iRfZtS/PD+rC3A0AqR9m0ltGvT4PrFv9GhJfS7Uu4q6QSMVBTIkWl0Wlr2r8
1LBCqsmMZlhIM/tgRXsTXw5CvUPWt7KDHOa6B46XjCafTZZyD7vpR09CRwGt5iWOIxbgBAKjow4U
DbTQZJeOrhm0FNkf8pptHpkgcivjnoHVnOK9aRfu+UcVcLi16PQnsUl/CrKl4XDiRrlNWAKwi+EK
ge20W7XX6HBAp8iCCQ5wpEocDKjD57exhB2nQhA/8ujC6gyMnA//tig/ysjFSb6PL9g6bJR3GvxF
uLkME0O+2GloDKreE6mFqO0ffZyXlLGBz10ymzIkB6ty1vQrD7f6RmiDJD5kCnOfJITx9N6OT458
dHm1/NXFURnejJn7pWGuVM9GSTWhElyVWwT2EdKctqBh5dVaRKwB6q78IuFGpq1tVTXOS5UvX2Uc
cxjnBms45TNMXCVfwkIjFHRaUn84woxyZnVcJZ2xwKWAIVdxxVrINdlCgkF1yMjUQ/WH24XgGfH0
9bt2DQ4zYPdkc4P4iriJfw9oyRsnoXgLMIxbE0vEEX2dtoBwPsCZOH1n6RmYMY0B9Co5bKtSHuqe
zWaZxSohi2kDZWD07wu9fwQ52PtwUW+BwbVFhjtc/GaDp/R6QKPEzo/nfwt+JLHFS2UzVuZIeygN
tjHbGfbOAXROOxIsHcyY1Rp6XQbeO5EAIOaEVT4yDMBB9uuphrSsx+iZmd7Ck4x3ewwqRipFZ34h
ukRSvrFScONlOYK+Jms5xmIuKkh23E4uRh0jE4EJPBSxD2CGSCk6NOyAjybqU8rp3KabCsZEArJW
OUSPahY/qyjdcgMz24NPleaKB5ZBNN4upOmXtYv9Kn8X3MofvGbEeHfQAvcnf2nqg2jlL+Xj74ng
zMA38Zs9lqCUYHL/1c7cU7SkhfjXTSn/isXOfb/sgjNeYjeQG8oPuYqwypa4fqGBqkjgXH5Fw4E2
QTDVO3RBZuFPz5sKzHl0nXy59+IAKSLXsGqlK2VFNZ8S4u+pqSLNqeBpTF7EbVtKBkdJvkE7oUfG
jaotXlMgXUEhokFIIsZk+r8Ub2WPrNu3Yl4KretW0oWSn4wY780F66ltBRly+m4sHWXv6MFxlPi+
8qlCeQUb986moziG1SdGL9VVOtFmYJXA+mJyBfmLUPrew1CKYE53jY728GgG/JNGO5B5aIF7xtx+
8DDL+smsEKlw92uywXR6d6aulJIyiE3pkVYIC1mq1Cu2yK4t/3nJzd6PZAMFID/SYE9CuLWIwdKW
HfJr1QZHdcah81v7YtV+ZgCZx9N06yoDQhHPYMHYH+TdGchvowLG3QAGB7x+ncfprBuE2GFNUO5e
ZLUsQb87V1tefriYKc+Uks+5+SWmPp9XFvshtxTXFsIsz7+pVnBV155/gf39jARCEqU1uba82JmW
wgnD2QVZQtSyxLELnfeFklk7HbnmC4hDVf+qPPIJYIBj5YJ57SASpzOsU3exiBy4mL0mZUFe7Six
FwI7RmhqvNuAF78MtF21tZydMHLxwBAnTOTWAiUlugYM0BwbGBbm/6w/U/etWkVR+VjxyxVEBmRU
MlC0iIdPr451eumg8YbixWf8E9GOvfoRJob2PhjGyFuAInr5MB7HK80oUWBreT7oiaKMlxfPdr/2
PTYRvV/PLiaST/PHMUKUZnokjKRCeoSpkxWiFUbLj9Kpy4B+B5UU/nZ31hyisw4ehkU7k4xhA6l6
Ck48IkwJgg88tfYOdX/WoQpxCHcsjt2hDw4Wz5OmzzjARgebyjgxnfcP6/APE7JGxKKjxCPNZbYW
PGSyZZ7yKy1pGsqHcB7OgjqhjtPsgp0AKvBFX6ln1xK1y0bold3YPKM1jvciGcB0ttfSYv9H6EOL
r1LqTx8f0kFUs620QSOlzuIHDynOYSFU+f2FERVC+wvV3wfnHJ88VI9iyijbzILpPdPYGMRx5ein
I2eh7kVgJOy0GECunhl6G2fMbfgcYvhiVUFZb5X8zepNLo/Xo1zw/XaMlaROQQBnz38PSGQ0qhfA
K42Vlq20QL+4DG/jKmzAyEU30nKlQVLp8uKLDuT/Ashl00IteWqFt+v3vc/H5sAtYtCDTN2ItuMJ
GhmmbP2iXOjXSVQbRo5AZJVjKj+2shzRDclVUSMF/EtSGHjGnoJiWQMUG+jriP7rNC8uof/dpaJ7
Ze7jc2d5p1NXUK/Q1q0QnADuG2StL+DY4oORWA66/hV5fJCkzeVhQtuN2zcT0fUCuR74aa11PggK
pbmTVoYZnKXBg6s1E27JfxzReQR9QX4ADLmWwKUZLNRdlN04z0uuHHaok4yjfjtt+rk2eX909fr6
DAvxN5fOv5oMfQ0odRqw+LQptwUNQpGQqC1UeFhfHEQo13i9dJQt/DUchZ4/eX8mpNKIdt8PvFoH
xWCUYBnrXyrRohMqX9Pexc5Y8cB4FdRDluPW8K8CuKeVIdAZWhg1aL53z0R5xg+X97GYhjBvTKSx
l0wzrUaVYSdGHUy7vVi6vsNxHoT4E6radALNrl0jzYLMWi8XhDvM0ReaZ9zWl8gHMEdRPvLmHQiC
ZFtki5jh0KImdaimlkXNDBVFMOckInnFzTd977cAmogUrAF2IlFX1nvnSt3K2TSa8jLpOsG4E/Pz
BEbLF7/gtMPJcJ5178emG9doBppqZAtUe8W1JUdXYXIfafDB/MoSy1DW8CHQDAUSve7cN/QeS3xj
gGimZFQom/XaJvpwzWAFTP1RKpPhFxpniERgovL2Nl5cn+gwqWdoXMainY/P2wYvbqg8OZQ/UuB5
XTVX1+aFgVc0cVS6LdQ45/ZdiiBfaN/whfuQhjE0YjqwkYqrGuizDGqYcA6egCptgt5GdxvIoZca
NC3JFWhitBOTkSjVlPTKDVBZGJDf5hEiRAIfDe9Wgc1w2dGvOFKa95QvV/O7jFndwq7ZZEDFCZdb
t8U19PhdreH5Yf/gMBk/YsWqdq6d01UkUz6AbfJ7ud/LH/AsG8GQZrM+hWaoGXL7LXqpztYUX8Py
tnMwbgTqu9ynr8QIp6EdCHU/6efHUArof8vwx+L4g5yiEFR3zk3HzTDe5xp5pICvMsoqiLfWroyj
wOTTgTRxCaInmYJmVA3w3F4W2IRocI/Nvwn7bO1h9zNQIV+d7m4dWODhnKHGLCCHtTtX+GRhBHXm
twTSTz+1kfQx998CTSX35ZBUu3k+jbccIEg9MJm1dGX7uCUwj84N7W+9dv9wFehlfWTG1kdhO927
BWIqSuAlDfZ5ZEYcZxALQEEy8WA0kjv0NVYgYMnCSULL8FkJoHb7ymeMsT+N/yzSrHrqQhPBf+mb
dikktCDJFMaCNbH2JOsgWEyEFzwb0pr9Gub4WIZrVAHmvIy+4NGUIEpUPvVVzIZH+ESGOgolx3bb
SJFLju5hi8z7RFO1lQ8M4HFHoWmqi7/3W3n28BZBv3XPPICgtt1FNbe7eRyKvQBIGL+Jtn6bSzYj
b74HwFXKzKX+1vRtrWkNYCR7fGutzuqHMP3LCyieixV7xnbJoDSt86OqluM2lS0ESAZHKm0eCYN/
u+qIW50cDZnbNQQzF/X+NOKG285vVmyXnvwELOgyzfbR4OyoUx0wRvxsUIOgxFLGhH9UBKIVBKcC
SxgEr1kEPkAp3r/Wm4eWvPcCDKzYdK5fH1qS748HkHpM/CTjpKSCyFUJjnJi8MvI9f91q7CHkFdQ
XGMahlKHy5IGz/MtInmkdZO1HcoPmDixJcUIMOBIsO0ml98e+MgSiXZsg7EJp4Z2YIqBwyMpCf/C
b5Imht9LQkCSXF4JEdhLy4CYyxZAJ4xHtecF+LD6GCvyslRbhalHoaqXDdUG98LDSeYy1GuGRgbi
d36nfF610yp2voadc9Zztk17WVZPhqKV41T3GwX1xC7OblA/7Ei4Mx07Y4iVpOhiRqxvHrdUEoUn
vTXcenq1x9bE7qzr5P57teNLVE3B29pimYgM1keQfmreSlJ77X2j7m/ycyUqdWgjAQhCjmdUZXXk
VcKmc/dEGwVt1ZTKxiF61Y+v1FZjvGLEj2o+1WffU+utiGI0RqWthouNXg33EguLeDpshjcxjMuv
WthjEBiyxtVV1VdmJzSbJo+0ZyBU8tD4u/kXijpwWuL6ck0IYn3a2Sz2C8GtA9626CN5W1OxSldC
yyocsS9YUOnhVj/6+QYgY4Qf0XWrDESHY+f52g67HHJXhrxl99xE/Jb1YIkkkbIe1ZbYiyr/SCCk
LpzVlXPUJ80Q+IENo99O8rhqs+HVk5p/qrEDDkuFY6SOz8FWlJgnTwFaYIpy6npijBcxCtcMdBTx
teULx76iIYwHD8Wgz2p7CXyIgm+dm4XU+9Zt+zBIbZsNeVjHsR9TzDuIfA48xLFtOSPLk16J/BUB
d8+zisZaHvNxbM3P96l0xIKWWhINJhP+sOHAtdD7JFCfR+kvgjg/0N7p57xaEEVfuXnd3Lpf67Pk
DFlSN9LzTGAzMffD9841L11HMKoBqQ9sr7tSu0QEb9bbRMJ3nNz7rPVN6dwEo/FUmvbGI7Yc9EFz
r0SXRn7TWdvzW4PbErBqrGoGhVL1Pfa2N8LGcuOPfnbWlO5RWZszzFsxXm6fw9hgmFjYrx4MvMWq
LY0Pv6RXMJwYlHEwdkVKq4M/cJY4h1I2jTJmqK765dU/ANBpAFX7TAD9F1ZuSVGO0aCYXLYjcwul
d90IRuYPMQhq+kGso3rLTYNy/JjcY22/UHdtzo5lVDwH84qNzCcP6AryiPDyZ7UXh7oGK7ODQkAa
/SzwYG29wkki6lNW4NnPWBv76xkhFlE/XYLhpQBPXg9wTeQ46uv9pe3zXkWcBuwusPhqKh0f1ilB
Cfa/Wm/YPkWVgg/HENqmPpqCblA25iHj2XDKD/qZAXoqnseGEo0j02525wDxFRh/l9v93C5VXA90
ms17NKDTUP+tBNg/KRVM9iVCmd8jThvpDIqgOsbbrRBlwnP5PY0GB70bHrDjDTMTw7R8z43lywqY
sDXD+EnRql5LkYytt0e+O97EYPaTd/++kpHMXPgvtNZR3qCTAkG3GXhXLWLrwJfFGm9o7GphSYqj
bs1T5r5J/swZa/BZWWUsz3nc8jsG0nQiGqxmOzjBSR2dfb6ugfBVAvP5daEU1uc+g8MjJZ4X7KT8
Avu5uYbaHyq6SMlBgpbTFoAYwdV3173JavU7+FN4Mdtucgv9spIp5oMeihlMVds8elzSsnq7z2GW
RrdMnyBgnm8jHmARW3BgZTFn38DUWK9+2Jy8ARXt9w/YsW6Z6H5miqyjB02v28wPT8kxyb6s2NgR
bUmhTayrhqvfW3LBWwXVsy0sf4M4EywpF+gfC8F+klxaNsjchJKdLKR1CjrWqxnQMGYmClqGRBQf
7v9Te739KNegkxRQT4BIpcsn9g0vtjMnzuHvcM9/UqP5vHTPL+VkaXLYWIMKh+EqApMlBvCEucwP
4gvSIiYFMY5LV8QjEH8L+BMIY/i+HJ0UADb/nehqsfVrWywpQfdtuBHssPF7jUnbySKi9aCG0Zwf
/hiIewe962iigI12ct7ENNTW7iUfGqQHWY4JgGhkF1tAZhvpAePHuYFCvxa2MRnYmvO+V7G3WsV2
76KS7Mj7lbQpVZ0yYIhtfjmw6I5F0enxeYTkWA67ZvoXVqMcXXJWR0GrE/9R2Q8oT32EwroBxqxQ
IDmMB1Y95zAPxIOEpN+BGqiKablfl2mNg4Ic0xsqPveLuLUjLqQ4hLd10dSRSwQIBILGziJkCQFK
OUa7O6QzzYkSZV5MSoG2CHApai/myH6o9uKpA+pRXBeaOKLJmu5RiuJoFrbqh9/5jSXP95qogN4S
oGq918Z/kVEpe+YckfS7WYbJ9GU5rZNUtnleE+VIbvlJflf8vZL7QFfGgS4hueSF/bn/Ikmg8WsD
pEtI+qRF+eoN12Nf1BcdQm9DogS/uyJlGZRVK6+X/VkmshYjCwbMGe1FcE/GHsivV9JtI1+prmDj
6i4cwcaUwmD6/GLicmAuoJ4j+ueXpGdbxZMi4IcwNniwBk+iH69NNAdVQQO3UIjckCJemobwRJDD
JgxdlcW1Xtv0KtvTNXSoTaqCxzp/NQoMSB26ip5WNM4QDk+ubLE+NfCb+pq03BflSChJZVElMQVX
yHnMDEMlfpomjY1oADVXB2MoUwoRSQY0yWUQfm/74149SKz9/6kImPb7d9jd4C7Ugtty6kwQFg5a
zSvyVmkcuy/c9FTNXqizQWlTg8m3rRsKcCVUN5TWCm3x0aS9VBujMiOyHOne8UMUdvPxj+Tlw0at
Cyfd49FWHKQmBXpFeNwzmf6j7tdD4NVky5mzQ4W5JBNDu/mU1bSfZZT3o3KMuWAnMvKuR2PmMt4v
nTZFXs1WCr5Tyd+QZjnP2wuezS4rGSDR2WOutxSheb4clRvGUF1CMhMA8IXlVAY1tfhwvWitxNuT
rZa5NflPXfT6oQfYEtacv0Af4GEpLbeCiczRhQiuDCe9qeRheV661/gvrOD2+nCSAGliTGyNkvrb
PQDokcFtyrxnSa3+pJtdG0dE9QXYF9r9MjjzZVL4xfQ3zzOqdavhqZ0gFOBBaJZz3LMv/AcYJOCP
NGAwHTOysiMpB489BFfAuXNFusz70r6uADBJEefWj1pljXa/9coGX/KDjvBmeyVQRHJl4TuPIhJI
Pj5KJhNb1C+nMVFu6KAbsl/AG/DvdEYDHvTqHTHSoNyzCy35poGVFPGVqeoo7kesFYFfwvOVDh9U
bSZFu3m6aQT9ThQlg3DphfiSr+sNNvgjmxCpH59PH6lc7KhF5VlbzBnute9J2Oo/txipZzNcQjz7
oDK/4UuR13dRmq1Y/alFFEwZlve/mFsJszNOGrFKxztKG70aZJLTNKuF8qawPYdNi7LUaxhyFOc+
RlwglVdy2z2boBE8xMCFros4qxr5j6X7j9z4eOPCJDso20TfCLvuZsgBL/iVA7mVdNn4eJOREydP
UAoV74dTJ+uBjY4qK0Hngox13sc2a8XSlhzKpufYcAJfQC51OwLB/WaqgnFKiB2n1Ag0rAul5MMX
+DSs3VoLgrTHtYS021PAHQKFFGn3ZEdpHNf4+cP0nd0PWnA21IIF0tHVQGO7zfJtF+MRdI22IW6W
JvP36e2vuFWVVLa9JIrPDsSlHML/jkFu+LD/gFTNcPrYpoRRD32e/GU8n2gVI1349KHQ25CKRxHt
8PS7xK1EXcNMsGUpmWAnoEKc7L1WF3kD+3rJY8qd5eZRRldAZE+5rApa7jpTcrvsJdC85Qxmc3pZ
q5w8K+iFf6IXxmbHoBqOk76NPJsZmUgRR+aLqOfMtmKFtvQVQ8DwklVs0lt6BDb+b+Zyg1mUdC3N
Oq2mGvuzH9tX2w6CZT6lifzAyPm60WTP9hhw+LyjD0uXZLsA1+cNtWvCM2/pqJ7tmgArzlhgmUTt
g8b7gP4XWhc0wbVfeOCAV4tWhNkmjxYCx2n4nNZ+6D73SVeKKleO/2x0oKMsiDDOni5VZyWC9mT+
1l5CJNYJ5oNTN/SWjLaDujrFabRBoeCnYK62jOtHE9jYy5Ds4l06p/mqgr8fBkt8Im/7q4hiQJ8r
anF6gWyRm6V0xe2xrmnIEkYU3gf00AhHuudUNQ0XJ/gjjohXw6cWmSC317avueDBo7eJXavciuys
XozkRLJJ9LFl/DP97pxsn4v7fnBunZU2cuKl//ODKHUBofhj97JK5KJJ21tqXCVnEXh6VVUT/gLE
EXi5Ctp+C5FZWGM8i5bg+YA/pWEWJwL1p8ok7wnxYq02y7J25MsbqUbyXVPyFRcLLDF6JwYpu4Oi
a1skJDFaLEAc0tQglLJs0nH6pdSdwpclqipbM0an32L4UauG13x47W1u95MLIWGfHiJh33PGinF+
jWr/esyhgnyBSy2n3sDPCIm6bkn8rMPauP3JEKKOXBpfVjuI9ljHdAuSKvSvk7639lWAW5Ew/OjB
hklX0cw2yivgsOb1+ewmgkBJsHXJdPvJ6CXz6uvpJkkouMznIQWqssT3PVpzqxnnS9byTmWqyj0d
En7omukgHavy3jfl6ZHgQ3JMEFqFzevyFaNhVGgv3MuQyvGHhZDMMiYnIaau6XhJHS/RotGMUNye
UCirEsRl1brNXmkD2ZZ6NEN2O9wHxngD0L1INb3Fcne3LQy7R9/cAPkUZ6a7homAFwEJ2xtcU5Xt
jrTqs9qlfu8kgJpX6S6FdjrxrQx41jRaewgVt1wuzHB3PL0Fb53GyIqozlZaIE9SGh0COLJQL9EY
cjfUDtwQs+XxaNyzY6de/WfX7iwFGGujx35FfpMcjOq1d6xCAyG7ct2N4Hpact5py3mtn1Wo++dA
rI/qSME3uaL0GHUvP8fDrDZqlsl4xMCfoNzmYcXo3LaoF8sqVcCZvPvsJlRmCj420KkigzeHIdut
JIL2IuPj82hQGMbcNDWfjSKj7QC6C6lB56aLS1HwNSgHGBqPKRjH9wWYit0hC71rp6GguURvdxl5
wdgk4tN9ntsm+S4B1jh0EW2KDPEmMLhBmE2CEcodot5IFtpNOIpwSKd4Zd5MfUzVb1Tv3BsC71iV
zoaOMeIwqNYqbHjjIphDFhRRAxXNGF+gSpyMQo5fhSRnVmQI496QSgxGYCEzLjEmaaIA0frVXVot
8Cr7blj0X3ocidwpaK1jhozgPvPdpkrjeKeYkJAIsLQHhFNGkqDa24drUVIQxVCEed0aHlwxVf9j
mgdJRYILi4xAu8YQmAr7Xx+Yr/t8plakdvgw/jTSJ4oo92zKDVPbOREQPfPsrZkK/2GNBKemkD9u
ElUb6KOrqYT18rkD+cptVGxrkDpU7mprsqM1fOP4Bscbn12o1aBFKVjPMmOZICu5lZEx68mhhGKd
v5g2NSlpqaqniqHdWhMPp15r+ZCYzeuGMJRu8UvvFByP37wUo/4b7MJ3dFj1THGlteZ8gUpdCM+R
h4coj6Mmbsc8rdIYVPPmunLMS6Z5BhEaUkLDd3jSG/kc7ZSF81m6DlocSR2GHDPSCDnusj/erFxN
1G++qEBb1eFvWvrO4uTJWLswtpuhVFGewKP+nmtM4eZnvCL3bsO+J2zG9QOpJFz2r5q9MqC4WdzO
oUrfjJzbALfgkIcip8mUgYVlKoM2cRzmc5lKGc6ted2tqsvCCgME9kMhl3oiNgQkhfk65rLjgpSH
cwRXpehRW8pMII3GdakKDyyHbcTcgVy41K2audmcUF9ug6/wXbkJfLlNwEwZ8Tg4i/3NZIdkqDsE
c6VyVGr0Qe0ejwFwszpw9ue9qPSWpqOrnvUaOFDZhc9Ki7SQ/ydIbKuxPX3WkR+gYzpf0MeDgapI
x4dYRKg0Hp7mI1skcs++sXfXqk9E5maRlblKtFJT3Cn21/40n+5t1tyh4oKD7kgoac69bjbMLgNp
Hm2Qi8YqnOgesBNj5qamaC5yvOVnEMAyRDp0cBi7LegTlQONBBWlfmCD1eEInlSE4BgLuCtYKomY
gA1qa62CbGpxejjfT54ovV/ftj3HDHahwJ2fA7cSA8al5SJISnPnvX03EtsquFoNyI12+mM6ETyf
fYl7K2rAS2g7WRksHvLEi/V5fdegap3nJT13v9RCeximgwgUbF1D3Pq0WCDl1pdljESSD6ZUM2F9
Y9zPQ9wr96hi5DVsUF8Qejee5gy8tp51exA2DKJP4noEN/q4Y7iLK1vyZw4r398qAyAzsLwM9SSc
MQ49XQnGD+r9O5XT7biX2wCQ2nz4GAvueifu/5XRBJDwAKVvC1Buy58uV/awEMAP1Zpt2yqT+eu5
ELGR6iV+FlQ+mS9XC1lOLldbbWCPNpNrCFERHqDUPU+2AkfdkGveZT+lEPKgIoi2URoXYJfu4DzF
Yw63D/ynxBb020oFhqPJXi3mWjyDzcAoiYogCU65ZOx8y1CyoTfA1lq20F8dr4lWdTznbUQx+Oz+
lLvvA28JKgHXHldm+1Fuaj9nGbcgBCBEBnsZLDfAL1jWtQFzwW0d3VvraTJFz7qQ4i+TXiRzNFx4
xakMsX/QQwbK7Fgafx8jRHIxe0Y25dUp6WIOEyRvH8RyqIBQRhWu6iRbSC4qZVDXh+hoyTOxXp0P
n4Xxq6ny9MC3JBIxjeZnO2XmfT70eeCjbHXDp1KNt+aZ1TXkEgc75zEKx5i4zBZEqJjlQBzzNdDe
71iVm7kU5F+Wzc55CNI9iDFLkmQzHOi84UUePEV+fMebkCB7ZXwEISuW2dqiy09sYKteGgygaunF
17Qo59WaLagr2V4QyjKv/IgFsruqKC3Yj1nXCV3Nthy9bdz5EoNVDeQyq9/JYXRSR+6sJezALBc2
SjCM8ggHZUI7V80ImbMcUX32nBJYGk1lH0KWgZqqU9sRcemmi6MF0xD1f/ql7eBvPJl1EGhnfrx0
+lIc+8hcYF0qPKRuXA7qC9EVDkBsuxgFxowpTjGD4kZCFOJF/1eVs/PxZmHhDbnxCIPLfBUADKZB
mafAdLUv2tIjrGHB0fOQV3Qr7mh/Q+oOAKnOCjoCPiZIitYjotX+S87v9mGxxXW4DmsXGpA5w3yn
bLKZ4yaYEcAYfuA4A/x/A0GG73ntqOTozJnjR6JDXsRa3rwHqxKlQEWnqeFUvgsQr37cX2qLv4cS
tWmHiTz9/C8m7/Ps3r3hD8zxosW6P+CkdtBs6oujtfzEJ/TNrZ5/UgW9PmNMFT4sraSAHlhM0vZc
8jhj/eGXOb+gVvz47F4LT3laOqBBriYJBDG/ETwTbnuM7ZRIOd6Xbhtueh/Ww1ZgVxl6Vr+CA6ZY
aN5b4eEiJBnHavvXtL88T74qWKiouqcFTyM/HaGKHBZ3a2PYNYptOKGMPaqqLQYUMXOf+rZHUJwS
kHV+6prnleLz+MiqNjes0cI0HuzPdhNwaRXnKSKFD/6rtWLKYuF+DPP1k2lMna+kpUgwFNw3+hXb
BxKoSMO7nPsQHVUDD0J3tt8gJybUVg3qgW99L1reYCe7K0bRMYVqcXJHdu52YXdnFZMoBfgiDF2u
16WJoHeOECn9+7KkGycO+tW20b/Dyi3Ps8LgwKdpHxOFVshjw41ziQCOz0cmKfintUUvnoGk11ec
s/SFu3Dz15nEBlTJPeNEmRcmuWPpQV14kzhLVrJvVwhvf9gyjItLiaZJmYUiewTHHumAyLRakN2A
eN3+9rMEv20j4wws+8Ln2DOB1cWiwvawGYnHL96qXlzfPcxce2tyfkeuvGE5UbBwEVV6g61yieiG
dIAFMx7R1MZmrN5h1QseGKNor7hW3Uox8wBEGXIJQNfLf9bSZ6LgNbPcyuYkVqUquk3KvDbxMZI7
8wGLg+NAZaSgHQnunevtqGCSG7a4+9qHIRBOpg1HCSMtQnkqpri8uF7GFVNmYlMSuQ7FWSXl13UX
4aIG9dQwlADweSRIhUfDONT2E3rIf/2SxJN1XjJlf4/fO6e+fQdIOsxxuefV/TPsWuK2TAiUDn2Q
LXfUDHcVR8j4gxWys/1nHWj5zc6eheNSogVQNh2kPoX4QlRh2vdj5F7Y8NnoGNjR2TXZZkie6Q6W
ro+1NXJnEWyur/BuvzEk8II9cw6pFH21+JBGlSk8Z9xyMayx4MHR8I3k7wzw9lO/KnXd2Ga9yASi
NcwaTF/3lqNepMm53+uwLLxUhbm60/oTfz04mjFcwwzjiGGoES0Y1aXaY6TxFlcprIGLV424HzY5
/ww8CQdpt/1DwnB1pxO4F3YiU0XtgMB2eVvzBiZNY7WCKndV8jmK0T/FXACGi6s2R3ZRyHpVbqpV
u2Vb9bVsoNUdugbUCnLJd+8MCHwAj0XDvMJBYrIeoLSglOVWdrqPlyvo8THQVOh07LGvBuw7RzKW
VLOiWhe2s7DQIo3L/IqX+E8YnNrkwONt7skq4W+/a5OhN+oPyskA9woSScCh56exuEIDi0Py3AiQ
goYDKAzvGaT1R5xrCRpylJbVjMRmNE6yrxxYECYeNFvq0ihXVUMRjNEvvzPwoP+9+0bwkmj7e/sG
MCplMXKYHgP8MYcqKJnk7Ne7CDDVFTjLw0gzNVxTcOkJe9PE6PT6Ch8dtGUSmY0LjIJKKxJ7ESx0
O8xGQ+woVH0AB0zTIGsWEEWJPK6oW0SY3jqspGklsoUyUrfAmMYYT5hYsZbhD2baG7TqnOutbsI3
rdYJy0maK8gZHRDZJ+hsfbM/XuTfSNGtlYEyWsbLJDV//Rs227lLr/02wEzHroaA2lPTYC2CMZBa
5ZJwCNJfGUPe7fTkzlTdBxrpKedcsbbb+s8moxrL/aMlyYdWTAgPshj0QOfb1AyPB9U9p7waH8IJ
u8DkDVTz9ncIgQM2TIhs9H7g4Th474Y18KcqnBBsGQdTeLqcieVXaoa1wq64yM3bVJ+I9bwF/NIq
CpBt2C2jlD2a+GMFvrWkQpnt2pJzTav9u2oieEUhnt/85SPIl8eLmfWOQaDxEqr6zNo498RR77s3
Eq0WERbpbI6d4btU+0LiuSut7ewm8cKL0T1uI3VxVfUzqv9whS2X9+SKTjx1yPQ1JPi6q29rZJyL
+sO2NkjHgcHJFK72/u7iXSZXQmb9ab/n4zrSKQIzR3k04NKt4ryJFXusppys9/LSsWJQsK9tfLnw
N3ocfimzIGTpyOBy6zDwVlwhXglLOZ/JYDeX96uIgFF3uwerNPdoJGpyaHVbvqxrilpFASk3fbZ7
az2D36qF88QL17p7avbO43GtRKJMhgGIbyyuXrNozQrkrX3qwiM7cQzRhmPlIcV7OsRG4xoMnxRh
HDuYl+WKSbBe6aJIsymWKq0yYdsZ8JpZE88Z/1HGsc2AEbbj6POBdNHNAQ+3IXQoGsSynz4Y2dwt
wInKX1Fc3yAT4uIJ7ltYiRRp/JV69qVUtj14lICSQYuva5O9moq7YP3Noi/I1atlLMRbeV44HRbr
VR1QSoVO93Ei+6zNQpEj6yRdAsNJf8zhCZFMOftcALpKZd4xStbxKW2gZhKZnsYZC2nPYJD0wdby
RzEzt2DYjVJreV3fqfHVqj3p1tj/lsrn3EiZWxgVwrhbuv3oQPVrq+pm48RUsVzv+Ef/PEhSXRk+
vcuWGWUROC99KCQX5zpR9U1lGgn76qQfST0jFHTugoCo88uKLImOZBmyUNr8On9oSGphxrzvq8fJ
hv4J4LcOAhjiG0x089DSksd7tShTTS0lUjq9Iivi+HVyqMpNsdMQ6gwwY5bIQqQyAjbtEM74U/6j
o5ELD9Yz5seCGfvUC+cDtyFmxjdY0KN/Qd1Tj+A4fLFmr0Fl5hiGT3MeUOtw4BQOfbBwnl8K+dsU
cUxBkQ1eymVCVy53do9Orh0vbSk6vVS3GiuGWd2PIYmRYq3G92CZ2tsqHErgH9z9aT0vQNkH6lFz
dSnNCqFErRajYA8ZVNK5Ukya832wLCy7TaGbsGTp9eqEl5eLyRBMjxu1NN13AfkSXbUK2lYAOxLO
mt6zgHfIqQ+bKaH2Qqp78ECavYm50K5MJftmCDfo+20bjLce9Ingg12mthM6OsD27DmOLVMPf5BP
5XoKSUCNGmlSFEOdmXbrZ7aYn5q58OFmThfb1EDnK1B54l5oN+dM1JGSx4i3ch4r6nSvvKVnZCbx
bO3a8leEbTp19ykE2q491JQxkMTHWumNX72pr3zjff/5WXYtT2yj4UtEoMwHwet0XH4U+etI8TJJ
0Y3jbOFZyzKCBASGuglsohzXCd1JfwM+wVlOwlABcRwOSSY7okSHCCHF1Au3h/3SkgRWnKKGfqGS
BAlosIHPkAeILl4j4DbrpVmBk1BwudQdaKgwpgN5Xk5Py0VM1580yC5TR1HbST8I+tWtJbALWjXG
0VL181llhpbGXnBrXNX6C74PDiDA/DYFdRI/yjXxWk7rbaFXmLcU5NFdLhDXOK244aKGhozKCePt
6aNhiyECBOl4NAmcW0edyBRJRe12/RgsCMAOQ+wW3Z7Q8lsTy12rYp5A0yXW8Fn4enY9M7STig26
3v3CngxivZId20mRVjhNw1WLNcXuYsJ52sePbns4+/lNeV3MWyWbSLsy0j/4JmbLhExRMARZaqWc
ZFQOiF9Hw6T6OBjrBHGHETNSsgnWk94OycvsrHQ8ogY/hR9FXsXiwF+0B6kgsyFVLMA/nIPqOLcw
nSU+HtpECaAkLbNBi4MFM5eeOYJQjOSASoFYiJoirCUKPexiRuphgoIS+Phc9lBsQLc4G7C1YFVd
6fDbMu7kOzB/EUysUfxGqjgprPg/1KsCBwFaLlMNvZJH5W0EEobfVfZMwK/Yk2+txfEe8PsIprtk
mOoPzT9vJXXCI0QEul6amkQCrcFYB4eFhzPhcbWRsM5RZqJDyZMmPS2unnIPqb9ZcbxAwEd/rBkm
aOC1xIOeomkSNGjduzMTw6AKkFNJD1CUCAG1XHL24gDfGemiXJ6xqwDYOSApPvyDrSkrAZQpXe4a
JWpdtK3NKQ7IGLRdOT6exrt94i24LKdE3x6s8xbP+QVl/DIH8q6KWvcCgKYNkYD/ZBcWU/UBmiHg
eF3ubUKAblB3amqpW0xqtDpr8wECSUZ6U3rGjNxdq/GL+IakUbiYsur3M7soClrxi1M9q+r7NU2y
eN4qBgMm+9pSuJ/ahFvlMcZdz6A2ZZ/+DFjzviUyYzL46Ve5bZWu74r/EI5KB8B9ch8SWl8l2blv
sL1CGD0yPAVaQ3MzdiM8Y4ylyxr9tXtQPzTWegm2LpciZagbr0L8Lu7xnkgu7kPTBFCgZQM2bjVE
bUNs8SPj4MZwyJCCIVah+sSUSgC4yJs7Ozv6mKFGXgD4leWDdmbAIQvJe3CeqUV+swRTA0Fldj3D
QAR2GfmHJjR/LmDuzw6T7tV8R/UkAOURQGeTucCqyDKFYNbPKjOOuJeTSeKkRWVL3uOkU/3ZEPSa
MjKRx2bvxl4G0JIpqY3ivGfF4RTNt1fHaZdcSQBkp2Jxo5XWX2m9x51DFPeYG6+syicK+ajyaP9R
xJLbbSVzG3yxdUcVfr2MqNiXwM5ngASJaPO8r0+Vg7rvTA5EeJ3TV4yHKdn03Sz51SrVow1Afam1
/+V2LSyIIFhW9hIFj5tfREnpQtxzmhLSHQs/Ox3K6Dqh4QrW7kJfjE/iOOIoWBcpCr899AHdn6g2
WykKqFsNw9BnlaUSLMk3cYQ5OCbJt6QpuU8s7fFH1husY/Bkl12n0CbtGcjoyfjnQSNgU8i1UaR3
34/kKzWrq3UdSsS2FHmNftg4oZ/Z0nAK969xqQBGiWfBZaJWj7IfOp7T6T60+l3m5DRJqvXymZmq
gJlLJKVFhW4/vK1Fvz+ogz3aoKE4Y6B4cTP+PT1RuT2Y2pvhDivPC7EqCeZLjEtXQ3vTvMJm4u9K
2z087Dj8ABslnc3Aj+eX19lzXIOueU82mpKBk5QoIK54f3Olzlyy7ssS44fKKyam8CivmX/rtygA
xpFJbkK07M+6CFK1exdSZNNthpE4PFSSvXDzwOJeyRIyTmCz0tRFFMutB33birQli41lABeTzNSS
LTrEOAiDKq42h7tu83deFjErWJaljv8C6jwwFKGB2bFVNw0ZoH2wzuExOa9hWE1xB5BeNhcDjRpp
EHUimKUjaXgHy0vzhWuQZB9tokGhKeWqCuNwRWOfWAuulTUF91QnPbyVUXypyIFSVFvEHwpQS7rt
LECHG+Dd0yZS8t6QZ6P3qFyjVFrqU78lO21AVTBbACXxBYb8W361RErIyPBgncmbFBZX8EhTAOQ1
Q3fuZ3dO1Y7STZ3gUZbTlXUVPbEwmkg4Qspleti7e2kiDpikJEMciUjUxF+aUj/sXeJJZzc4RC3+
MtKJvSRRsBW9r/aTQrv1azvQ+Dl4a0TK2yxQuuDOgTF4ra9UrGrJxXYpsInpojzxepV71Wgk5IER
0/64UQwKzyU8jcCsEozKbMfFZ+rq0CGrkUe3l/hL9vWBGCIXiblb6F3F+YF4Xg/9aienlbJH93xJ
NrhcWtrkLr1D5X1OaNiWn9yOgejK0HcIo6o8ESYxHDNgA/iSF6l29ZxFgNg/WvxYj9RgJuVyI1cN
eYjvz0mIs1SkL7isIe2l1BgQerVve+JF7oTLpjfmU+RJZ5tkQkzpBeTuV7lVA5PH4N+at1pQpcF7
8TbIHlQ/xRZszEMIrzo94Z0RdsFROn9CX3BxC41yU60W0qxuCYMZRiKonP/5zDrzcXm3MchmOqLX
yx7ROK3jZABo7HEeKx21id3J4kwHfbNHbZOsbsgHemiW49z7SY3M8m7tdEKHURYOe9wC7FPZnI8Z
5dpSKiqh3RAEclb5twR8n3C30YmofMU0p2FemnWSv6H94TirWpSQlvoK3UFZTS5ND7hRoxsBuqah
QurwWKSi+wDy7enY8OPKvMkS+p+IvU3Tju3t7wB9vcFA4UhgiHMFdeIE9Ex7585weGg7VO5JJyA0
ORLLsZkRA6J4EM+8h4nhMIfQQhjUEk4jc8dQh6JlJBHsF0qu2e0P1E5V3k3/parZb+93RF3Xaym1
U3bQnwZzwW/3Lek2t0ZYvBTP0k+0jWC9HKzYG/ZIBBbGqMrOnTWYCIE30YLJrOCKwDU7Kf3ZaOnC
B01jLSDqGZfUj7ssBl4FVTnu2xcmgXN6yB9Nmnk5qLxNMOOebfMty+gOqNd+bJT0M/LLPB/eopXq
DM4tXKVpfrwfzG0h4DShowd+8ua7+jHPR6ORMWgRlIQ8A0+oS+GE2gIhFa6fDcscD72xwCqjeUjC
n5TXL0F1ul6XEIZYt/7kn+vJ4WPLgryiVa8LL6DFeLi92WKtOlF1arzKKkaap7TCoofFxEjQhOs5
7zSs41BuEZrs0BSLZhqXF1Np1Sl2ctoEIZ8PKgfuoc4gUXeS4abA+047zMCxAwfDtqK4BNlwjS3l
Yw4cEGb7pNJ0I7sxGcNE6P1vP9ndtGwt0fmYA/1jpyqwlrrNNZFgc1Npi/Y9NbDvgJdPragENJ5T
gQxPXrpU3wntXeg8JUlKz2wYzzLjAbEjMmZWAegu/rKAxdEf7IB0wrkFG12OPswGe/jh1bx+l6jy
nouQOffdvIkENw++qRUyZebQA8/p5CkpqEVChdHxc8QrEBhlhxMCO4wGrqMxN5tQEXrfgtdK91P0
SBaoSn4kLCzRM8kRuPjlMSTjjUou1cOJMsyffX/8rwv0Sr1FqgESUxupUvdohF8q3xbpG5F6T7Nz
864AsqqTmXfINSuXzvYGVVynymtwZlqT/P1xET7mv8G4sASZ/ZHOS4inGNfqDn2AeSleD/wZ5sKm
iyTD1iCsKxBBIWjz4UsIqFbRTDGZPNhVaFlzHGEHDsl+P/uzK49jJqjRj+hh7WtY+AkrE8SfJMhU
ZIQrqNZAA7ilc4uMZRTzO67kcQ2pOjh4dMgwLM3gs+RW9nB/bHXwifpDFCGnKZUJ/i3McdGJ38I+
aGD8Fg6H3ydKIp4TL09nlPLdBfEjlmtRrDrrfgdLhgLLWXW1LaPcwWRWnhPR8F4TsfoegzdW0xJh
Ytx9zqasQfB6IERoADcLj6mifAx/TooTtAmrcm5KICUEyELPgW7nZUBS5WmMqnHN1jpOOx55Y54s
48FwwRUn2B2ApbRgrgR9OHy6B8KD/vPS86mjgY1VGG+IWFWA7tDnecBz749KHwRmip55ObBvqZk8
oxVndls6e78WRD9Vlj5elEkdZImEOSrVeBKyxDL+2OLqJ7HpA4skFvLoTOL6j/E4hXo3vuJ4Xszw
vIfAVWtHy0Ax0AkU6jOuI5w85WsWjpirf8RFF/IvmntVBSemeAY4IX3bG2y0uEBqst2zt7pHC6Hk
ufZetZtsVjLk+8PSmaXCGwsKC8QHKAyDdClnKs7EIs1KSbr0C8s35e96JP2P0ZoU8EZ5Rf4PXiMq
A7wm2j64Ykq9UCXuNn54BZ3ec3DksPeG1Ow+rNG3cXJjf9ckvE0oZR62kBE60/JNw0N4N37aIfN2
DTjrx3r6g1ANjS/8rja39mK3c0uFLGVlBjKzf2fvZxEqK8LDJNUYTRlV/5IKEYyg8+2fpUQLmtfX
d63X5OegMrKt0B3XZWYkn+CC7KH5kEnKa/TDlYdi9ePSKdwSN04TDGm1rYB1qatfKI5qbn2BEG/k
ZhtOiatyV/P9DwnYq2OeU8nj27B/GcAKGriRuEUIf8ogPDWqe2gWa4yNPH+wKdtqQx8EQ00RtEyK
+M3tOEQWLtJL4nlRzICfuOjz9c/Nct89+ACgvqjW+hYVwcpV61DwdsRyg2D30rIGO+XzGOXOzlM/
FvLhI7qgNPf2OXzwoaNqgkaZwWbJXJBZeuBF1gFz1fRu8IfKdJ8i4Pbl6RLWxlkcI92aItEDblOe
6IXtqkcdQNnOzt+2lmJsNfRFNlMoyRF+faG5X0SE33LGD3XyrHIjED7h72SnolZGpQ+c5DZDfjny
0/RzIzE8l1SM18Aqx6O+ay+JGUP98G7lomn+sS4ZYbmgYsZ7Cnqi+2BIcgm4WQ2WpoCU0Uv43zPO
IDh23u6BZgMRvaQQn+yalGi6u/JkGi+dsEfHhT88qxwiouE/8xKt1WM1ljyJwzBgdzlA2PDecT65
JE1pmcCPciW+hG1gwpyChL2SeUroA6picay8YuZ49BOZL/54S2E2MykyPHrbwaqBg9ShJQpU2MPr
0GYvOqnINJ+X5H4ELj2LEGayBFfu63xNOmV9Y4itAWPe5IkCMqfCJxwHvE7EFpui1jA+5FzOLDNx
pvDXaU4VeNyiR3AcEzlGqz8LP98QdV3omoMVyDypPhxSXqcR/zXp2JbWoR7EdVSJ8OORwZJq1j8g
6taXGE8wJ7NNXI29ZFa1M3KwFAEBJrYudPaC/PFMrzbYZmjjI/x+OiAvePUyxOuGJQSw//0a+2ZI
L6JzJ/cIlRt5lZPffOQvpGxrygzU6/XMEqhmBIx3TBz1yv4qOBQQXKZfY2zWI8WEYwXXqGtD1vvS
EnCUkMvP5LXsSUhleClan+6y/HRtwldwdkxqrUgw77mF2mDpsMYCIjMDKDxWKpq95MA6PBPjN2lu
rnJfSFF7KJEnQUBNPtEnEMhLNlehD8+CO8xSshrVveRNIaGPQLYl7tFIXh9QvhLd6hYNB2VER02g
7yCaZiJGi2a4R0uEuIyjLOSTh7u5ikPsURNzo93hh6OHjpitUhrqsrodoakPu78pfYugQoMivdVu
USvHHtsohc7PoY08VgJINzWWIqYnWcc4Q8QkReWm5o9sv+f9M3dlmTR2XpEn73naGvmJUlosjqdG
r+d5cZGgVlsbfq8XsKggsEcZb+FoCd6sBJemv0pWGYs+zcfR3Aow2OsXeP0OOx62Bfkg6nBivzCB
MxkOq7mECHcUkewS73HMnJsfgFmgy1AUfgR8k20UVccsBDEzM6LrLlUWFhSpo54wtbGdI8u+EyO8
jC0u8FLwHHJ6Pg4rJoC3DRfEPKfeVpeH1IBk5TyuJkQa8Q2SRH5PTH0cQcPw65dAlca/CMm4CHzV
zCZjdOHMkjbqCTylIXcfgEXloPJZuyRpm3vEZAeF4Om0OtjqWy2s76LU84Z672gCt+8/aKT4MgHI
SMJe+5hsQwYKf415KDY1hICtbuQVgh344ljiv+EtlZiLGBqqrcFUz1erWPJQjBtKw0DyuMUb6khT
iN3IPl490Q/vfRp7DXEZYyly+cD7FMUQNarg840pabImtXtimWkRWgY19rMarnNOyBEtuYlJ6lRV
4vJ4tJsu/RiROA+Duw5WdcmtZoycC15HCFj5dv1XcKAsOpzznqz0mNh9pF2b2jekHNCbaUrQ3FYS
RTrEhsIDlW9oDh61F5S5IFKyoh7rrwrSJuqY4ezcGhfYbu0IYMI6KbHUVabSPjA12n0CO56VNGKa
3fnKWL8y1DLj3QxB+ZL4yCoh3AWNEAb2eIchsq/4O1k/u7iFbnNRbznY+td4xpHeEvFCWI5NdN9T
APo18uv9Cu0imfCoECo5WmTtbPDBcaV64fIj7XeAe8gKKDG8eTwgFmLjvkLTWYaFDORjtbAO8a7l
MPEYmeE4ZzdyOLqFS+JSATW+igTwLPR9kyv0KiU1QesLbPTk4uLhID/lst5oy3bmJNtz9ihrv9Ie
aflEAmQ83ddIs8oK+DRP6dBJEVdobH0PVHTeS73kmahc7QY7Qzy9t6nk9ZY5jqXFypKvMTPKKyp2
9eIp1EZkQWMUvg1f1AUUfMh1jy/kixXyO/hBsc29TAUZZYwk28VmQKe8/qDtIDVS5cL8bIinRwHW
SwifFzC5QIq1i8/4o9CIy+DB6bntlIP+YcQIqTvIyh6z2z4VRIyqogzfzjwxfQ9FqZN2zt0e85cU
QdTEfUUK39UbsdbSch/UD4Jjd41ofaugDG+q8V5FDlbTnWB6SFxgRzp9iMisxZmXxvzHumTgVr95
kDY8v9KJmmMZkzjaIb/wCoa6LRBTtfCgzgw2Sl+ECF/8iCsyEHlyEbF3xpxnhC0U56Ztlvn/cGxx
xRGnbVb3hYyTUJ4dta3Aq8DiCdAttq6vslJ1MaOEdOz9b30XON8t3s8qKbtVqwJ3rCD2ntVuhwB9
jgn9JNJEVzHmaQuoAbRwtmCsddiJivYhelFfl1D2BNvm21LWt3ZjxiUX3OntJcXO9DdE28b1Asg+
W7Jok1XNYwd69W6XKlUfCo+UAP5SBOdXtSkhMdIyzTdvdghOejLXKJZ5k39kIEh8/WCzfF8WOWQm
FCEYZMQXP9jEMcwEGLkEtFO5/XsDAaSSswj6zTdKHJgpIPfEZnb6jGkppp0G/kmL/Qq9SmdzCtXn
mnbAFV9XFZalgeU7BW3oq6yLUAQcEN/ViKH77v5FFmMR3rlB/xz3iP2tgy0YT3W4P3+SJzN/o9On
yZ4yZ1jlHTzXWXzyvdG5WTWQAPlEOKexPjVrGY4A/1PWcYo3ZumKPcywQJDptZUqogW9EoNMQVxR
D+0RliDuqVyj2Objhz5iV4gxvHbZPoSSnR0CepRvWjEzkEuW6r5Dz0Q9rBSOFpYkolTF3VEE/3sv
XQK/3anmesU4byzsNbOOeaMZV9+2VXScKAtPZe1DD8XSQ6NbLXWKdj7aFyYFQbLWq6s6tDEzTkWG
xVLp4pAsdW4Uu/Ynqs57/UuTl/hACHgpJ5r6bzdR5toRCsBRWr3g46CMKRlrR19s+NpT88valMwd
TDh7yxr5SxkjN9PYQKvTTo/zuRRuazLpGS7LuhGVT6Axpi1I5IcBWK7sAe7otvNB86lAWdES419W
lea3amk258lTwBWDZ/TndsfkMAaPZgCficLDbPR/Bc5S7B93omSg7at6yLIfNJYxgIMngZtbVdkI
IBGZUqHX9kC5RUgKAr5gg4Prsewl9WnFHWPAuqaQkLFQTMSmmXc0iVhaACOj/Egm4x3LRcmtnKv7
QkMkloJZq402lDTgVjY7pkk1A9F6LDOgO1LepksWR7r5wGUcci3le8/J5/Fm/M/5G7zmz7chN6GK
MfYfDj/G13BE0FyFwz4j/hPNb+B43ti3P1BpZvjIS9nieHKE+4PDX9xwKH+a7lDO1fbkcib5KVSv
yvvQuvu5GE33CIFwIfPOOUZt9anPrhG3i5OB0ZyY7i9gk05ODPmUW4KyiqQ4YfmHiZlkA/Nvy5ph
EXILqgL7CE/Rn3BE12zSlZ/aJvyA3dzAPkoepbzyPShTNwZb4LwMv56pK/KuOzkiRUwURkMYBLpW
M/u9MS97W7orF1vOZt0b+IR0w6HkS33pVrDchEE3eu52pFyPG6PUq92aIMiKsJE4wCb4QUrb3WVT
BJbfCfmxZQHt3rvlXJgLoacV6AmUEZ1Xb5ADR4XNpSVymlRTR0mN+DJaGrVS/Iultt2dLiNHCJgW
ylNLr3G3yTb2gpS3i4JMy0P5WwqXA87LYbJpDwKpvEhJCucw90ozuxDUUgvMUBEoJRDNFXNsJduR
Z+gtpFTkqEqYyw94QHUztkQyNnguJDxQKiC63IskQzltsaYlMNeh8vrFHIwkRGW6KX/qFamwEcQr
g7hBqChsCsUHY8JZoCMbSCEdNP94YtlsjSuo99N6hjnZvxuqDDCSCcE15GkCnVsYpDbjF8HluP/O
F/bYHUVNYBwWzakK+xFyKgwmZWd58hCpGtBQfqVWpy4Bw9z3FFoFgGusjXZSNBb+dtqO4Q9UBr6S
6EkgL8WTVKDwXbDXgJ7tCqP7AIL7GCl0Y2qN9x1TqTY0YzITDfBQoEiEQxQKJ+BEyoKAkF666g0z
zQoqI9AYv8jN8jphwEtLsLcTCRNEfxx3naHo3nJP9SADjhFqaamwY2yVSivEBNdoo2ZTRcNylGBA
d2YtIxFostFXpTGjppPd/fqXmn0i4POilRpyTlz6tdZK7j20h5QQZ4A2BzbFNxV1Pupgx2t8erEa
oPdlxD7mclYlD4//juj1bN14FgD67UCJBCUj7EH5MxLHJ/8yXhEMQUChzf2RTtIJFXobmZI9k5mx
XPFoB6I+xs5nTA2tu4TUxEoz2joe5ErkvYjuJ/c+hhNvhGa6+05uLnmWGIZiS0zJiWlZLcVQBB/Q
7WYuTbFvUmGJvHBToNXyhzm+jcbeEIa0Vy0hlDz+aE4ij1IRp0KHhs8iNX3R7uTKdTPIZuX3hjUp
gxYjmphx7wczfiwFr1xETA7SjtRAJyV1gjd3fT2QBBq3tHF6wVZ5y7666NdBMaEgzf7dn7m6zwHa
LOxaQaxQtiZq48oFefIOR/ARsUR39Z7uIpN9lXpREPexjPNhIyhYUthWlCbhhTZy/i6fwC1gDZ8w
yGwwBLUyxwgCEzxFiNwFWXdSVdh2mK1rylgDhH1zhk8Vu+MWxauugeUz+B0JnwMhhW5Wnuc3AH+K
3AKPEdt1nGRAiGB8l5xyhYU+dPqZoUIFqO7U1H4BH0Jhg9ORb5ywX2dvEjC7j3C2zHR18d2hQNnW
IDLxFLRBPQH9hJn1zi7QbwVNtVt7xfLyUUJYJVOd8mwNzepfFttt/Ngn62KrGfpJrWA5mf8LeHzI
MaOE34k8hf3LcPyI+aX8IZwKHPe51E3NAWN+FeWrukksSKZonH2Bmt8276+roaDWbj78CRJikHCw
J6cDn/C56oO5mu9PYMWFsCJ9zTts3nCFcSm3tFhNZ3AQ4Eu+AIqm8gygSlZEHlxOj9cIuV9Pwvsv
Q6EeGI3XWIYONQcNQvpzcXS25Uii4BIFuCkVo/yx7OyHyYA9PZsJN9ETN6M+M8yGMh0WWTEH7PY0
/cWrwCj36wjxf5ILPWB1Ak/SbwBRlLnVRidZ4sHV7oaI9g8cFiCLIjzw+jx2xjrKDrgPpnYwbE4G
lyBMAxZRcrHko66zpuxNPAgEByoDlr5zU/PSbOtUhJnS/npMN7A6cfwM7TjuHnsMU7w834iNnlTY
Rw55CtPHKP8nFtelbRmDjB7OadV3tncG8VlemG+r2ILGkmj6j5n0ABP8qT0+t+MzgTWWGrUrkEOx
KeIqJ8UFnEURVMaQD7xbb3of3D7UtgEXXJIlZDf7ZNV+T9HV9Uvi0QwEdsgSlsgqt7kARAQyNEKl
jn38e3+40mnqZeR0mCH7/1s3LFzlSNXwVFvnvH2FGtkW3TfAUuo/d+i2lACeTbMaUenprw+9aa8y
PxrZqlIeqJbLU3XfxsBPbVkUZD5MHdnyxurqg+ZfLpKo0sMH2hIJFZbHTrP3HD0pjQu+kgSvlMZ+
LVW/jatq8UqSqCRuR2pxpJdH6F+8jjRFnAHeAXMKHvbbe6UpE/k0kXSCTaOfSumtkYV9VvD4Vtew
rnHsTuPdmr7KacEoSEPl+z6GIvYD3aPkO/jD929moQ6sB74agBleJbO6tgvwnvb/RhkBlg166bmc
nbYUUPYeBUS+uDiT1euSSBaCEORGQPApWxA82Sx7sneGAq2k4H9Gc5F4v86+z18UryQe25uWT43M
U1YJSMnqMMuadbBKCceTD6cTEosAPSxqT6WRSCH3hsnMM6DutmF2IdqEpZeZyWQASF4QtQVlG0Ub
8AX3jsIsVkU37eDNlk1V0RI4B5S26BqWu+MBrDScY1oz9rLvODbYn+TEaHThX5vWkeMJcH3ZIpG+
bB7pZWLkpQ5khkkSpWwyDkhgf5W77ehop3xVYUg7kBr0Db38DEatiG7o/rPK5Q3+su6NLEkaYh+M
jAS4uj6a+75Q2F0fcwfEtizN28j+CIEn8YWhw0C5iMH83ekqNPJ9uiRjqy2pwic8q8oqoD/B5ldO
wqNq1dvXAKZcNcyDp3opE+l704E0oHhF60U/OabuoNDKqBmeKt1oH0PCDtfaYJDb84IEp8N1Tl2m
3kiFBGCcVSxbb5/IIG9/ux30lOuNBzDePuncqDhhq4/bfdzVWD9f6o5Zfhphe1thHIBS22uwwzx5
dlIxPmnvgQn5yDt7ZYqey2SfyV+KPXPYbP6OFZfqdBsP+VeAPFLlIvyu7BgMQ7o/5ujNE0EOrcTI
MJE4Zy7cQYLXg7zaOLHS5jvsdO875CEMIAAnc8N7aqEwX662CKy00VpvLgSUwiiINuSg7oeilUie
YMkAneFMQfn+lXYlJVHEUZW248mrKJmeSrCOsGdVvcD0Egi7USSZiZqyxpx+0ILp3e2JUfPBWEsz
+C4RScWFjA6CR1HwqUu5egoTcYllDKFmDbsPdiyrc7dNbcBnWfXfSaxDLkoXABTweWNyaa7nTZpV
95c+110hVqNXiftyAHrcZ2fkttAbKky9llhTrpL1BqRZ+JOORijIWL8LxE+iax9J5WwK2j1Xs03P
XOCAvNe1QTXAyqzNOlBF5bA6gQwJMtmZsiEWOKo78oKyBvbR5JmczzbfNhkLy+0wtbaZRy1804Yf
k3zDsRsqv+2LsbI8vidDcxBJdI/7uQh0ZdamUAvCNnz27z2XQJKQWozPDsojqyf21rrKxuri+Giy
bTZ3+ueHk0fTYv5/ExtcXUTnkCt74AIULnJtYp5Q+H8E81HakJ8DvUAn6q/JndEBatkpL6Av8aYG
4IVN9Kra/+HCI0sXcGaXfWInjAZdMwH6ilpEBgVuf5331CuJXu6Qfg10HmEngoIa1FSAb9QAxgqV
S43QrrYzFHzmjnq/6nn1R5b9n6HjQMuEMXFgyW3PioFuaAIPHN36bCgyIxVB2gqIfWkRIHwk/wLn
1hI8t7nKpjpk+Nb5Mq8PMYTNWauRAYIxpT1QXSWBQ4u100phmNPLvTKvFFW4HL012uchuVRGJ0eR
Gc5cT3+IwyUO4AtyQs2TbqIjaes2KZGzLR+9P2URvX6LxaHeZgHvavNW4uXTNoCNMEzNx5i2kDek
qkPjTPvSHNIfrZ7moxALDqkjzYCxhFsoohvdsCFdA56KYYbmezEIeKeQ09pieZ2VCutJRf4qgNgl
OhpBq9HviweAnMSdv5J++nFgoLt4jxc2KCGg7iH6ht0BNEfH90r16PJNkDXrFXE9w7BvnjYx6SEM
XYH8v7eCfRHXREObkfhlKKTSslYSXRDBRiIpaVbSPsWt8M92dRLGAesDcstO3P3iBFwjaqvUkwuf
4u63Aao1Eskhj8CUhRBxAsRG7Q2a4hTKOYLYsekhyWouInXEm8mB7HtYbwOHo0eRNg6aMtanNnzi
N22lshiLMsQf/VZE3dNrLBFzMCuWUIpY5D+9U0MZmua+xMF6nn8aPOeHi/lkDPpGFHzdcJ7qU7E0
UtTO4FdAkaKPa7qznZB8W2k8AROx9zwuo3GZuU5qgMjZ+A+TMcOBN7uhLDYB0drj9tleQpDOTr1o
/Pt6kM4lUPGdsSTUCsIrL9lgXoHPhemFbPe/if4vFD9aGlu48i/35pBax7piRZHvaCDuXDnsePKw
KsBgi7O/0NEeDNEh1jc1ynQZo1rmUkK5D4e3aPDMg5DACmo4MhumIjWAhoQ2maEnRX43ijfmZt4P
8rg8miDndMtREBrS3VMt6k7Wi0AaJHZ+DjM9jgOPFAvc4OR5tEqOQzsyDwXI4FbpEv/H2pGle7dm
6kp1vSE4mu/Qu5VAVuVJzgeZVxw9TJcjUNbTR4vcILjNAHNO6lQUb2apBzcTQDKLAYRDTKJrfOTG
kb7afIAR4y8DilFWw08UR2SwlJ3UDlVDXk7PFyR4Bv5v7zHFEDxYhvmIf31v7+tUIP0jSfjuCsio
FZNTTLODfTK5+GlNTPCXkFe1L1L6mpWVOpK57r/wgQKGROJO8NDYMDHyydTMSvdiIwm2W8BFdv4H
5/rYp8m2DZSPxDutBTrcf4hLgy9SXoW5lf7B9MdsTlqfvX3wJ4i+ctjWb6h0JMDUjJV4bgAAyi+V
afcP2asyFZJ21R/EDMcCrZR5SdotXd+wiXEVTUx6zgMfIjUMwOBcsfCwAOIaNwuAzbZJlYsrUGGR
CEBkYgzat3O8t4iJf0WFbWaimNEIyGpjVWUsFObNLBeFIjQ8V4AbRPs07QPtr62ubBwgGWuS6I2I
fT6lJuDrYKcZZ+uuni2QfZYufUAaEEQNqJ2Avw6J7gCAIovpKWMIoq/09V/Kc8Aro4B6ybokHzgf
x7hqSn94UY/OSfevlu5Y/O+v+H8vummrC4npX9pie2lk6sXOO4YBpOqXfF2dOwOd9KTD7+6c3yuh
Id20+5SXjKJ/X/+LPlTix67f26+x6OCF475qKpN7I6X9ejkEqP9WyuukMZ0aqPd0z1ipveXFFCUf
lCQiKQ1LSwN4U74v5pKzDuU9PJh4jdubRPw0P39BUwckcdzR4QLygq3TcT0DWDQjSKlvylvwskK9
qiL63D7FeI65rog957b3N+GF5gKBoEV/zOwjYXtaUzMw3W/G6cJcQ7l3u9a2hDEQP6mHeqd+xtyA
wd8wZ8yJZu26+lYl7R3qw8KemR91W+kbapLMP8FK+gVvWFHOf6gkWRWeCjSs4JJde9tisv/KkkSy
lFy2G0t/kAdqZYXwIMCdOJ02uVpfskGqTXPngeTwIhmpQuy4YdQJWH/BcLm61rmzND03I0tksKUy
i6y3p3RAgNT+9RnhXCnULhOMInDON3ACMOSnXpyQxpCAk1C9Rcsh1GlbIUB9zIRzIRJgPPc5lVGi
iTeMC/6sCI7toT97eyOirx4QjyVjrLZ11Zt4b8VF+kKB0ZmFZ+tqjCnMqVkOVSWqeCawwsReigl1
jfKJ2WWChqZyaKBAnykRyp6ikoGhqqcDlasqEvrR0kz3WoWdExn6XxX/cIq/hTmPQ2MoJsBtDBgi
63+667fH3cGckHPLrfyMuOgfoEZxAfKgLiTmi8dQD1ldcqxPb4iOOHiSQEBDa1E7Aaj0ysKEV29w
ae72PA62klqk2FjIscOnaJ3XR3jvS6P8c5EHtVNC7b5FVZLeU3sXVYZlpsHO2hCB4dr9COXDu33U
Yk3iSzOtn0lswgammrXUcZnzNGsj/CxdPLUhHKVCpHmDZoA99xSJ87tt38ooyrHywVepSPRplQSI
XvSE2Uuv+W6XkUivfs6bJyCzqEarE9FRIquKYNE7IAbKFHApY/icQ3ScvuHKfO0tNQS969c8iP8C
Yf5rKN1PSz3lpjibrRcZA6Hd8ZQM3XomnYdOPu86KI5WdudO3tvP0D6fQcmuOaYY8NmbEw6D81mK
DG4kc47XVrZCCFMa9/g0PJ3feHh3KFRk6dE31HUZZcvED8XwqLd7mxbwtCdocqjpnb9g9ZOcYFCO
yH8zE/Z8tFj4PJYKJM72ee2fGxSuCrQqTKhDAQTbpxX0GhGii7mm6fbcto0WeD+6dxEqIMhMifXz
8D85tc7R2RM9ffk+1ANCPQkJvWGkEqGuX/eVr4kVSR8vFUMQgvsCmLxPULof8ymzKmw9VLn8T+Aq
jYH1KyvLqASb9VSttkalr3qRW9bDQqjOOhwtT+vK3uvV3XrNaw57KZg8+Q+iuu/bHcggjwwo/nES
1gZjMi5RWhqoguTGpmLyEqeW2hT0a/UyC7NnlYdwfsPq3518ZwSPushXGLOgRPsAF2d8LN1cI8be
eS8Y+9pG7gC4XZSEUdZeVfWVTVn32lqpyo1Xeexp6OMOxRIjrfQHo+cQ39nunuhph5/2sbowXiEm
m2E4YwXiTvzJ/K3EpljWanPnpBR3AHbFyvaNliVM0vKXnL/uzlHCMDZkDO4M5BB43jlpm+hd21Td
IS1lxh51b1S+ebUTBxm5ARlAB4+XOj14wEIbB00dcjXGUBSx34INVZnVuH2LMVxs1fVNCTFC027N
lLioIq/xzynixPyeYW2XJQR3QUBv56qeQPI28maY+F1sGoX6RyXGpUB/vt9mC+vJaypBJl7lASyy
ZnN6Vh+LKXkvFg6N2nWz02G0dzPhown1WKXmTL+cVcXgXa5axXisG5gTMZXiys0s/cEQLvqp92Qf
5iC+iPILCDG7SHF9e/o+gP8GvZAO0N+yz8mV70ufGw4aod6wzlJrKpvd49tZ1QAvLdIWwXStDTSz
E+hfjb0I7AhK+TWX1AWOd+4NvUHbcNyqtvqUA1TJHb8UKCtEXZ2nz97VHnKdJ+b6wqs0pL359ghF
O3cRBN2RuUXXJLQl/dRyZM1MW9mfeA31QVPY+/f8HE/lSaboTHiroFsaZc7/nnGocKw4KuGs1UKm
qhGDTBAEVz/FigK96cGjURQnmfAgkt7ZyEA/7xhQBQ1sHTpjsqt/t1ldNwt5ZDM3BD/I2ZQsze4R
8+Evb1/OTrtYfCIp/ppD67X8jr3v+MY7bALdD1y7TWgIzYRvF27EE67W1LZMWBgtMCpGRLybWS36
gPj3vsg6c+sZ5A3iprSjtfE8wfmMADMuLxzaweH7SOZIVZN4eRpUhXUvQKI9xluS6541l+2eY/FE
tE2B4xhkpDG+XGy3oZJPtFkpscyjGwRR6TRxRKnqC7u3fuVzJnOglr+xGl5Ld9guzj/o4qXBqqIH
kXjrrJ2e4gPdMP9OPofRM3GcFKxiSWq7h333q9jbJ15f1AupZLu+cxaFaFde7l9SJYstITkHpb7/
C1VMwaCOSy8DVXO595jb+ChJKINQiAVPPajh4Zqosgm+qy1nAbONAJs9UCumtnV4osVlJ0RYLcNC
tw2JbfZ1UmU3dMuNrYgOcjHR2zXr1wYqNNKmcFcsV/zDj8//+wi3fp4QUguQmGd+MssfE/0xzjr8
U68qlUNANitwJCRU1BiJ22DzCDlMLvoh5sdHdPXAtOYdcc8u3O0O1abSQeJmpxyAfGqG3L9rx5hV
EBUFk/juCAc52S13NX9TD4aMlnjAG4xx5jGjOYb6QXx/7cRiy69YSNf0M0K8N/nP1PMI+jXzF7B4
je3V1uuspcY6lggOc1CKT2mFLH9teN1lSStrKH00g4SKwr2u07omKD2Ye+om9eOoU/EOofYQ37N7
PjUyW0JTAjXWlArYIz50SMfkoclWsK2v0kQWzOril5vOQM4dLYDLbUOzKrGOlMfq0r4mc6FOHk1W
V4cuIDC8d7w3Kc7O7utZpq1Myua9+ftKhgjLDWY4MAA+mSV35sn2T8RKRQf7b9GDl7n+hmoKX6m8
FatwbuoLjrBAJp8x6At4MB2pJipirR48pl9tcfXnaxvSjHjIpAJqbojRm5BkEpaqH7VeeIMhLDLu
eaUNBm618oIUzJ3WKiVadk69T10PenCEaPQwbdJFJmVmyqNLHzetmIFlYWQyUS4IX+oBAGUfHWJs
uCfOhRwa51gB5L2N8BmqI9ru+UccKGXO3kSP2QpYAtAW3l5fP7PcARgEfmSGeXrG1zLLnMRpmQPU
dInSj2+YfB84iQ5QPNVhmQbgdJC51YSXOyvWGw8t7wO2rbVN4Qdn4OnE8/cKfvA/G0JcGTGGNX2u
Dd4OCzONDzNwwhusFuz8YNuSKAElMbcN4lkLaq8EU1YMpcE4/EtuD+VG+kIdbmi0DoyI2rLoCZSp
gykhw1oMzHSasbhVhHMeYzPXwU/72onUJenlpircc6kLjErjxP0XAx0H+ApFz5ZB82zO70z0TfYl
dA23LWnk9+JX6WDvQFqAGwHbljn+lNQPVI6Q6Wrnstq0JJQvz7+lb4vEKqqXoWQqDk0FBu7ObRwS
dWqyNRmUPDV5R59fEY0cMwIQs8ocyLLIxXbkULsFocrxcDmvMaHdyuEM8rjbS+QmKBpMquQpMgM7
owWmTkit2LXk6xfEaeBP4fxZjOYzbR8HWlW3jLGnU5mhdiaJ7XHw5JA3cU/So5Y/0iFVPyc+/uKR
rvR5fIV3Q525N5DVWdmhlpnIZEPvJuPNB0Dh1RgKXQliS+1U01r/8HDXskkXuDBo81C4ykp3YgsX
3xMFGUv85KtK5DAaYW+vIBGT1V7LV/6/x/s0+iun18oCdRnNZNhoiRZxAlDAoU6QGVz4yUC5RJq3
W6fAP4DLqbtIeB9HIyH9rTWuLi+4ZZCZiLorSxu1ukEyhE1+QEmv3MldM2jnybZqGteIjyhYXJgA
8dTE4792M0QJhQYuS4UiKfgXHKm4A7SA4t7w5JhF+ffZmLzoDKG4Hlsk+wY/4R/DfVTWZbHHFghm
inSmv2y31B9lkGtKCdLMtX9whPuM7gqhkdbjZIDGSTluJKwJcCbAh4F1Nk+Z6yTJBIOawPMcVtvl
bpbO4/+pBH9h2DD0BWlw7oLifHDKMQccWfj/q7Qf7F2k2s186jrrQkHeGZvFV/TZUh0E+oTSVzVR
xDDnTs9+pzvX5cCSxlmjWXDHC67o292N2NMOmFBUOdB3is53tkc/OkMcLuL+YrBWp8742SYUyVT+
g8+r24kxsGOWss4F0gVffgrMUKpuQQ5pNymwZmAaw80opDcRhipn39NgnuMGntRXLTHGG9+LHKji
ss6t7UG8u1fe6YNmXoqxycaZhS8Z3e4AvokP1ZM2jL2dKwnXDrNHfJi5dQGLnId3wN+qEnnCpXZe
30i3HqydtvJo85xAc7ThQ/Jk1XdeeUlhOQVai2KzUhg+mJulbCrz0EVHnqeObb2X92+iccITYc4m
BNgq7l4HZEeIW4sUfjbr1gO7PZ2lFxsBFzyHFH96bB/obrhBPsPa5+PZUiA678PeX+DiOg1ec+Tn
D7DC9XbsrEvIpb9GhHpX+aR0IFeMJ1UFsYVSIbmBSaF3Iv7QfapsrO5V/Wx3Wnk4q2ExblDCoRiQ
3R7slSZy2F102BjDDBEwn1kRFCOo2sLJqR8QUtERJP+lp+oJyjeWmaAWhRlv5xdd0bVM6ESRqXgO
YqGhJHFV7swC3szKIVsLo4ypZk4ndBnviojxxxu2+vaNA+IZsNMgvMIw8NilEpLQUZ6qfSBZAb/r
2H3AF0GR2MKKjqkoHTWH2oAj5jGJRJ36560if1UrtVfszV6AriHIixdpfkM+FJY/v+lKhGbQOsj5
DK2OrKMwD+G8mm/Zf2TYt1zbuiyvkjV37FsZcE6Db5cXQgcXRPTJuzJxe/6fOwBK3tgb+kg5QZRR
nexPaJpyKw3ZlqATJed8vwaKuKKhkLg1eWsc81Aq72XCPaMtM6qBiCmA9m9X8K9L2TY+ZWQwGpYP
hyhDt/sJrjTnqRj1m67hNAlncXvTJ6T6dNABqnBLlwtbl0tzqjKmLMiI5cTqmAeUFMKEYaMrcpAT
Gxtp+w6PeF9zfSNljPrNoVxBxd7oofM18jom3uqlZ35eJHcEmV/1A3v84VRw3YFMRjW+JYjC/b1Q
H5clydmjWUZbJTma9m+7qvdXfOWVftRQZccRDWODVu4NysFH2I4/ljScqjN9eEbYEXwonXjUu44q
5ExTifbk8wlTu9nplCQpgl5B8vlbDLW+f9G1+IYCb3FlNNmL7qJ5oaFQQNk6UbNFO6rK1JCUuze2
fXMo4768iSfN5YUtzEMRI15wJE5+GM+ugccLADD9gMvu9gQ6YUcuLvvs01jlvbcOGkujN/dRvxRH
y9BQiSU2RovcAVX/L6M7U7CaqufR6roK2EEhXjVEE/u3WuSKuT9BobJRD7rW+RP6bO9aViNpfICH
iWPeCgntQ9QhdgaMjuc80SlMVG0o0ioW837PJxAcjsqiZACEx/hOVt6NSqT3+LjBaFrTf8MlfKcX
wQ2UG7dC1zx+FctnWIwNb1SWNZ69p5Lz1JS+ugB5ZsoW1Ij0koBss6B5vDY5fV+NNOIkVqd8c6l0
gA4bpOSNi5PBKIjiXO6FkshaQA4rlzE0V9kcoAshWJ7SnDSVNpfY32OgZenmGFkZOGvd7EmKXcjf
/zw7jQiPdeu0hO8sBn9PmI/HWKjReqIpq5WnVXCa+NFoxitTrIPyrKuj5/iXgk5nnZNmfxajQr7c
UZOWlqpKX8cuMyL8LsAyoIMoEk2uNRt9TW2P03+bawo9zBodLIl7PXT/g+gYaiMhrVd3tfp1rgaC
frUL8knLGClso7mIdhWVR1C+Tr/YMq5q7ctpKJbKdyRCwJBIfcklrSRlBaQU2yqnidyO/8/He1Vu
3xq4Mp0IfDx4+zgyWAQ+wFMveMg03s0Y7INzCi2Vmflqa7lwmpQYQoaWKUouqFOcR1FK9dx4MzGG
Sn8e9R1UMbZNkVAwciseM21fRjDJPow0Kz8yzl3JrBGxY1UDKezEYHtU2zHdWoe/4lyoxJBqlIbp
e9yVPz6qe7/mAxJd+EnQSy+eXMFfCeesbscIqjqDhLjQlouPwHb86C/Z2M0nMKJwy1lHLD58R3Fl
bdS8khcwEPQ7uv8XFX4zwPGoSUmBDl7S952a7F/NCEhgHsof03ZyvaXelIQK6neNfs5iUuOU2NYV
V8z+Jvtg5BpB0eLFU4CiaEAsvZHYZzhxcQiMC72QMfWshihzwxyZQzP+Et5WMKFbCspJLicwLxp/
/cJgT5jtM/ToZ/uGXtVvjDLMMZUXwyePfpL5QgI07RQFsizSHALfAoNcHjgDxIuGZdbguXmUe3A7
QRlTvuHk7INYvND1UUtiIGIpDuKQpaylx8j3Cq81Ipii4iI7xtm1fHNSCxeDzuE2V6vMvsWS5/Ov
sFUP89sK07x5TrMzvpmQnvcI9HvMvx3tImIEWdaNZxiuWk8O+UjORd/g9LAvEghJ6xoKbJsXil+/
Vl+n7U1TU6TrXtxNO5Eis4dn62+8MB66fBQJsCh6xfO+XWa7Ny390gcRMpXreR+/FoQ4vaEcdEew
ZuGamj1BjJStodp7QZGSTFawup3ea7YHHb+kFrAc4UryKDEXdW8NhzVrG5CgicU6+P1pCdgeEYXM
DbScNHc+ECaovG7pBA+ZA026b9i8J1q3iJQvIN7h0j/WA8FkbWvqTLQ+zGqxDP3q0yjskRXY/6mk
/Ye1/3csh3qwAVk3P2IWmz3z8ij6ssKtXE2VO9SPL8scFsZOdSaTLRapY20/50KG76P32/qm9lo2
k+P1SwP5gHWWLPYUbw0sCURZjaSMtLoaUZnbJeollnvQZtZ+4Xl0F8OZ2FYyBA09QSIef4pYsZsi
TWFnyxvlBeFJnDd9PIAZ6kefo7+2icPlg4EYHeNIZX8+GzxrrOtI4a4hG1cnVo3BbYsr9UJNQKNc
K6lgcSLW3qDTsycBdfhIKIA/fxHj1gQRS6px6hVL8OWwDtUrcbUsI10o9uE70SLvgu3mCtmxcvss
YhPp09/ie7NjVsEQ9mdBNOA2kpMd96gd3hKTlRpHwXPt8mPFigM+oqExfmkkPh1VY5TjVOA5SDH1
X4oTCQqa0OXiuH6Ap8MNpMTHELiigoFg1dxMnF0ZAWxPGjavnwBZ5CsBQKqTLPy5Vh1mQF0lHdaL
7ozWJPyPeNBX4ZCXOpSCIFo/Tp+P84fF9uDk3vEKEgM7Yc2jCi3aOGcbma9ASXLOLZ1+9nu5TT1C
RN92d8EHSAcOdonLQcoweNhBDCQiXiAY92vPdHXFCv5E8P9lX/TAPq/jx2WTMfhLmpUPauICkAFV
VeYsEs+VtgiLReCCTas+K7F8+as+d6O1nT6WE5p1Kuma2OdAvi8YtR5jFdfL28E5lbJfKKb+0aPQ
8HYX+0d7Q0Y1P8LXNM7Mgxx1pRpEGdGCndXGrcCAEoASaVp19yPGDlamwKntVJX5QxzvxRQc/pgP
w833svkvWd8juikOW17J9parR5r1XYm83ycHvF3LAfSdSYUHBHt5CpXx09bkn4gBeFmygD+99qZt
AZ9WpoMmJTurnGnCFcoVI/8J10+Yo0VYywu/5p95hy2gahSm4FaAzILuh+gWppCV9908bD42jeaN
qcYXHW86THJEs3VKtJFFp9oQ1WKxPhMszz+oseQpS9DxMK5xQGGDSfTnp1YCB3pnAqYzAwGuDJoX
sUGq6nuoT1rCmuhnrPPgZNwIqZUV+owhdWjhVrwB1xgFYyzBV36R6wLqfEbESRjiCpRgNLitrIkN
LbHh0H/f3kUhkiAJDESwJYILWnGB7nMvgjIAExIs5jFfc2XDtH9NWwHd50S70v5P1pRUrgcb6THv
mL5ILcRhkaGk0yXpHISpgktgqLTXHCxSBj73GpsWfar6FRGH5cfWRIeHgnAxGoFQCJM/c25Rs14b
FvR4cBYDKLKQ/443f2s5euDfbCvF6uQZRrEaluX/MA3atJ64BaFQAhJMFFcydQgzKOYxUR39F7Cf
zfau3kpQYUtaBjGeHQzEVPImU3vRc+hfiZzK/j/Z1xKeAdraFL1CqABDTFtrkreEg/RpHGBpWhKT
vwNQ4Dz7T1gutdJsoNLC9BXeXEYceWEU6oNLsCTwWxWe2+MNbR9R5iYSl1+DrDJFcxG7wjzssjWv
q3DvvKqToIbn2W7rVykciq7dbREeS+w4sYCEmlaxIRSRTtqXL7SOSqxF4NwDQUUXWPpSJc2rBtIG
W7mwIdgU4xsIyEJtxsTRlIIJhY3AbZO+SnoXD2mQGUDiDq6UNpzd0AZgv4DfXROaCSB6QdbVumbI
HC+jlM2ZrsMNDSXOcL0sP81lLwQtAHk4cgvUxyr7D0dPiYIM43npozf12FKGxD9hh7N7mcSpQguH
mRisj/HJOeGRb8fHckmfyqd5WeNRgT0ouWOsiz3XXXmxsISLtorQWeivy32fjXDWsk/YAutuHoE2
2S8v1ADe7D4u15YFtK1HoeyfsPlMgO+JwcYLIZKDegqZhscKd+XP9R54iAV4aoHH3Te3abgdVKa9
LS7OxYzGtH+QH6myK91xf0QqWsWsegIYcHjM1pCrgdxQ0wi34JNjg9SsuICyCADRLUkycoWcho34
KIP60j1Alth995nI6pA8Ezk3ZCs3IJ5xh1R3aeZIZFiD7DkHmUYC9+mJI6i+4bFfubd6qFJMp728
NsKLkWE7IELF+lkt1jyu83I0dTdan9QrgYbzd28vl9UV6n9oYk0KNi0w1/kyGygWrI2sBEiEU+9U
lK722d1r6wTmuvIWGyewUKQO5wGDN/JYX4ngQ1yevUKvQPRO/5UpchoHQ75mzr1ichssJ/qQglSs
FIp8Vnl4YO+5nJpNOBNsFM2Q022kyVw3GVYDCwJb9TVROpGf6wRWIQPYq8JsWpFUV16G6aXf+aob
RoAAOIM/1stWL1l6ZbZ4WtdOkiP7OnQwIBWb3uwGZmj3MtFJ7LTvdjqSZjvviG8hVGkF7T1NcpTI
I9rlnNvxUJzqNH15vXlDFIk6I9X0R10uHG5Cxn5jymICaXj3RWQpdx1Ntf26oQPRMMWkj9kMpyMb
oMr1IBAwq5aYQdw3gmNGRQCLqz+EOhqJsfnglvz4Brbkt+JA4MnSN5RkYSZXWFEgu4CBpHwoheXQ
MvxYrj8H7WrXr0F7njwc9bWrMQWlSEwSFfOiac5CXoPHR3TkBj0UD8jEl3HcCiSKrHH1hhG86IML
VIFgnjFI1kP7hrxPgnkB7n033Hu4eS8AVcyjHJb5JvzGoPoJkSNxTWBiIumPgoFVAz5TfXH3MN09
oHUWntD/439KMw/kFRqXQIZ23WlWCwcVbr0Jk16uHG+alkfUElZ/1YSTlL0YI3QKcy7Bp9JnL+2J
0fNpKDFNQ5hFJ/aFqmkDOvAJaUcEqljUMboQHA/vG4xX+ruQsezi9EBdm7X7rJpSz2aW4rkF1poY
SyjJ1JM+NIHbM+j+7CPUAw5HBc6jUxYVnz6pEVboeLSGUziawCuNGPTJ+kRE6TSmQuNefbm1dRSJ
vkTMyiL34PI+mU3fE2+0XBiAIC8dN3FzWI+HmzxgE31ddYBPzNScX+0GQ5OWdyFKRRaaRsdEY6my
ykIt0b0ap2102YeE4EcDijhtZO4ybOSik/hRP2oh7h74aK8aXFL0tvVGaz9vIiDEqPFWYSCAo1s9
E1OBM+Bpt1c8cLo5FvSFZjuQfJaR+rv6pyd8X8/gGFYfLnlxapJG3mi7d+4s+3avy78rhPCiQVgw
sQi9GuAoGW7r2d1Fh5Oh2j4GswZzmhhN/EB0w8HsCoFYq58X5WQaKosYYfmoLL/kB/XQcUcCECSr
ZmZqlw9gFzV9cCWD5g9jmZfSqeLKpIDIk+oUSuHqVAbryD5c68c2PG2fzv/eUMn2wjStTbr4BUk0
Kx4stYd592oBrjgDViOqI9e+yQhHG2eq0E5K1l8LAXrXDgV+Wq7VuGznDJh8HY4V+pL37Gd3XDu5
kXQm9QmYAgzXSZRBpPufs3uj7Amv9O2xifeQV2U2ru7Kx/MOulU2o74QYRoaBAT3UhX60UX/u8gT
eIndgsmTMtzD1xOD+v8S8w0/aRIEsS5khTP8oWiNCeaf/ym4FHrl4tait5V5aipX8uU8vP4fCVhz
cM815gF+cY6KGQa4XbbBtmo1K6JU+hhOCFPCRz1y5BI7UvNinPYAM8Gh9h+MvuBZNhk1Q7sWYSnf
BwjrrbzfYMdBel7K+uI0s/Wn2D8bFDlxJgq+NwVLIklsyV+TYcvkdiy3RBkIToeH/C2nSerODB0L
F3zaNhKGI7PATy5YLsxzsCsVQ1KMsiR4abuNkm2JT8onq+jd7GVViYrWARKDez6ga/4GCyohJhTr
pWhk5d/KcWJXLsjr7ptw1y+ySJK3mNJjT2mmhy4/M3/QZCpvG3F56nxwKXb0m0dExouq9sB+j3Ek
8itWRa8ZG0Z6hjzukWa8jqofxXM3d3UrQqAlwsmCMc6MAWP6ejKlmBiFYwSZIp8g/C+24v/qQpg5
6bV3b+cmilk5R4oPl+h389qn5RphUBHtefe7Ogj0mtmULqLAOmzu09MFs6oihN5yrJSO2qyR24SU
yFVYwOL1UcJf5eOG+FbipXzsxuyf3G7di0qXpSFYOcN+j0nAIOM6qUF4IIhBjU+2GgPeUliv5Z2F
RIvN9ijTT6axen8ZFmaQIDaK0Mf0Glf0ocQ3PLNOaZJORYz1Ripu6bl8fDvZNvHPVvvdS/8Fu5HZ
oMpahj0Cn/+22T1D6wnyuJzMFfMpsJRSXHe0nNZrg1NlSri4151Ekm6Fk4+sB+5nEb5YFmS8XXBU
q/0r5st4xeoW98rlbuMv9rujBqMbFGZiT1dqs3nc3b8WwQn7QIUcxNm+gwDHH0tdoWFaDIcGj/cE
dZHn+TD7ruYdDmWgO3DUGq+A4tC3ZDJkM7QLm6mPhTOmKk/8KwiBpL4H0sXixDsuF3ZD23g/u3n6
qr8kmQxalHhruW7iz1Ged+vcXWcmRK8z4BR01POCTObbELiIFUra23lGgysql/62E40wbctXZfrE
ctiI8gVEkjpcKJ34Y/Oas4tAvGOyGT4zldG5wPK4bgV0VG8q9b2GSlIVsT8cli3k09tBLyE6c2+X
7w+qH7osFK4Q2lpM/dMBS+pwdcagySd1Ia14YESAZ/DKbc5IeXiZ/kaxlOZPTtoBa3AtGIcDCm7Q
SzsAmr4u66n9J+iG3rdQ/OPFX5S6Jgbzh401Mg+H97vnddgGqQHHrnSzILPGyaQxTygxL0//KEdZ
1JkYzSYsMMEL6s0GfgdkqccPKo2q8jqb0/k7FHozQEIKKAY6cpetUt/82OXUU1XmcUOsE8qtgOcS
HkXFeIsHQGcoqfza/JNQv7lnbj0H6ymvCgrEnRsmUl/iYmkbqVr2jugeUxuatYahlkgMzsF45ROq
WfU0qSQDTTMP9jx/QeReV9KVVpwQHrK5ckkAPh/H6EsmJ+h4VGd7sK/agxVwFlru8WHYxj+lwJpv
XcG7GIm15acjj6JGjCC62JA7YovdP8+g3PaePirOQwGFuWAANetZRTcFX/d6nY8W3lZf0s99nTQo
z37q46I+sXnurKm1HVEL1hFCF60sB7W5FUYVGL42KdQlwLifX2/8ENWB6AZSiF7uMeGKJykX5kDQ
jJnNL7I4w7yzDPa7CaZ8RwfcXS2E/KPwFlR9XZ7ALWsscWTmrOZCIwvspCNyKu6wqrV5FS4lh3yN
y3YqZ/e7N7mjpQ0IvMn+d7/TTkycMR5sBMo6W0epTdaUduwgIYqyjz04y1Vde/+FrWL4HpaRLLhY
0oyU3rFY1MxA9SNuVHSP4uEGVNHgOG9kbG4DetFnab15AveP9QeLCcJQjmLzFtWawTxrbdh1pPqy
MD6USgxhaFG0ENkx0btFcG0sRjpM7ZoYe6tCTNt1K8jsMODKQA8EydI6O8FZDWrXwUZ7oED17qma
B9Wm3iXW84UTh0BVAhkvbm+DDJID71QCB/fyisenKqqnM1MltcR91JIKOGPt8KIqt9Jh5OivfYen
M/1Cqqu34PJ6K1WfqrFfnr1BdhM5lMXRzeWPlmZ4k2v94hXau4lJqKfYDfp1IN1Pc3hwjDZSPqXL
NozD1SP8J34zNQ9gn9SKzS3GBuCkh8P2ZwyKZ3faT81zKx1oHlkOt6VlP9yZuPnU1lL2zfIgfD/9
nEW8T7l46J8SWTDc9f8hgaci1neCikKJbi05KJKNhMG6FEqPPlUzmbbN65OqKTWDto5ZHrtW4FFL
ElhEDjW1lNK0cuczObHN31yMH5EzbLvOoARjsEXNIIuWlmPJaf5e+D9pNRiw4mbqvOk0303glfQB
z29wgK2mZLkeuTFcdBTszsf/yamiDkTvxzEEUcZtwEF82i0MSD/ZuQ23cmShO+4QexT3YuOgq8b1
9yrhO6zgs0t2C60V8jvxt8nL/hnuB6hv/6Do1lwUBEYI/MPXut9wxepIz74TM4M7cVxOR7qupW+p
0QKJGow9Ywq8tWQ8NvixAzVhBURsve2R00n4ZBg7R5RlmYim7Wc9oPIhVJd0IIbZ4HX2DY50Lu8j
Ii4S7bekGVrj01wr91i/VFpLphqc+xJLD5eODIJz4n3EVovMrNuWw5qnsVJlEFpeIH4/k6VDWOPC
2knIGN26LqZjc0RpqyzN39iuHp9Fh701KapCOOAX05lGV15+TV1qwzRUMZeSe3rt5AbZ+EeCIas/
xJPEJmOX5ICbmc31WYWK/vWqwlYp2ux5N+Mcf62tmlv4s/EPJ2ztntGYJhi3B0zfFrN1noeNQsDe
aT4vxHUpeT1me/oheFDJI0DyWfxBamhVk0KiJ/0F4ipag06aWnumZf7OptepNtqqdrefLJ+0ghPb
pgtwiYIl0z4DkDEWrMoArpJVcYT6wsSuHp2Yb3ivmtwePU4f/BLNUOF1fPsiUImG7AihbtiGKbKd
SNagyd7/6zreYnT4D8mjJnMUEmx2zLO/oH3+sua1TMm+QBlzIr/yJcb+eFzsSinwoT85smb34dKb
u9ye9d68/Iebag60//+O7HDi3g2xeel9ezUMoWtLIGN7zpRuKN8dRxiIZsC2cOTb2N8fjjeTzD6U
0Gmtkb4FXDGrYmMhWngwje0sPqY0NpGW7Kvt4cwi+ejbQIzy8fXQzVteumXMjk2Qoao4DiEYHlZY
hCCs5cArEEdsIC7Rv8BOEv1UDQwRMxgCQWJCX8eOz0FBKyUMCxC6PLw05yhaXGHVbwIQaDtY2lWC
TN/zcmTkNkrrfTwWI2mcjE+FhKCQCR4TxLt8qb9JfrOXsZW1/yL59dCUXyv/OBICadBvZuf7Vosy
3r+d9OBuI8CxeSBXhNNeYamss9MWKskEXI9USnxQ7/xVKvZ+zQRZr2CbDduTn/1YtA8yUCjk8Bo3
vlq33jNLe7xkUFi3AtCmrKFIeG0uLHRvBGzAqE2nGJINh1IGIvO+KOftFwG2esOHDb6gX+51/9IZ
v4QTliEfJxtWh/aISGGP/goJPH1dYs1I6Ne4VZYdGcF+UQP5hVHB7fYEQ8jBPcfzTqvClch6vEnz
vM98ep4OQaKqv+AGMZTgLn/C142a/u1ZOkO8JJgpaeifMvvJmz9P1T2rmbqQYSI0YQ1K9OF2OxWD
jK0eL/eoXnv5cNBQq76GBFzbmzD/A5CrozBKLQLQB5DaXx2mtNmHRsOmqBH+NU7LukLUO3CHFyTf
g0OFlTViYAyz1DtRkHoyemEhu4DsYPZbVorwCTt2Bnc4eBr+FScReT1palnLp2jMHFm0pceFVUO0
rR8IRsf8lOXkJoXhOmSCG305SDFxzXumwKQExqWJci2sUAGj4AAfHyj/57ZY4b5p5MR74Q1ovfAB
rFiYUnTQE0aiVXYs8UWYTBPOve7JJiscJE3rcCxoUV5ZgmKyoC16iTCfGFoitSiwn+9jv0XXUs4t
laAvH2/TklicPctAwl4CGCEbEt4BNIYLqCQfzIbMXFDrVw5Ako6NOiK1c6XvyRiSCXY8otG2ns+z
XAsTiPFWOEqUFc42XnbU5fDGINjXoZpf3OK6xpszHIDgRK0w80n7PK3GJzoE9nHYz64RBYplMwHC
e1jg+98xcO9aCIklCiFZaK9hCdGED0vzftiX5QaONmiDy7eodVSvJJCWRU1V7MVjhPnKexYoiede
ciflVVesNLFQBQIHoGSdWfApbaIcmAx3dVOtfMIRQRoBwiYJ+B0qHWb3L6JULQ+v5PnYAFnTLB8Y
JuTCQdbYLSstRaqFG7YVvhKS6kJI+FbduOHDK8S6S4cIFQpNlJHRw9BFWDcdgvZ1YftW7ZYGRhyd
7lAnHlG//IqtiTzbA84hGqXe+EZmi9iLH0Z9s8kbvMDGHSyN8uLv3+Mx7FktM0RCeo9+j/O37Wvt
SHlVNsYHG8C1X7ZeUppQATektDXzQQLV10ymYD2kSNb4Ge2dy2K4hop8k78Snf1LnAPH7bAOpJ+T
bbiD9fvspZaWn5cRA2PvBqjdZ11qoSiIqUXZqoCZW0B9SA31bFGO4LDDwRlQlTcqYM4MahpqrNmq
mlGy/OGShMKHh6HDZfzyO2fDmNSRh5zypdETrGzP1W1TLnFUwDWkISUwGZB/G0Nxsa+hq9dh/Gt8
Y3WgZG5NOEeqUdFNvRDRhycmuhpAlL84J57AUE2qSm+6Mc8AGp5S6/AlZ1nCq+tUANk1d+QXJkct
jQ5kWvmDpbswESE+euGTw8PKwWfCikgtfYV847ssfsZGJjvX8NBDSJmmWu6Wi2F8At4g0gkKFiY8
qZ+AH5En2yM+YGI3UtYIIbFw4V/pjoD7srlqzbcOlN5nPMjtbLSLqV3GIFC5YhBoprFMxtRD+5Cw
ppL54Pm1/AXC6VemV4/SkO7A1TGOMdswWX8wx1WEiJgiqixpzV1McFdmQebW1M4Ysjab4xedwMp4
jfiH5Q5Lf9B5O5ULLqbdTx1lOvQ2Jy9ysdrhN+uWcRwi6WeMd+1W6Ju3y2N8QFl6Grug5/6Gdmx3
zJQ+A+eq7ZEcewBW0dUYiaZ7s2YQSiIwgUGk0+QgY8zeP8VbrxCNBEBI4PaSJNjaF0GFiV3SCQdg
kDMi8x7qYj6Z+d/qdydu/10iPMjBKSkupgdf0FqLIzemY7fftCmkV/cSNJmoGxHp7VF2FkppLkLx
BTYUxpKQZPRyeIhoTiS1kR1x+LmjfvB69Ql+cf+34ACxCEkdScHhF6jsWivyryF3osBfqCIZtLVm
ZvgZIOTGchj1oC9OMd0ImjpWRC3N5yV4Ias1Mzf5FITdmYwLZgHT/c+QTSqBRoDcX1FuLSHgpYii
MnVZT2HAm/LUPW3s6sSMP5nagBGI8Wt+lfn7B5/jnUD0Mxek2pQoi7K+ppNkk7E4qSx5RxR/R18i
CoUKohRyK4vHX5SL4oGH/SOMiS12yUV08aFqTNyc1M8FsQjy0HuR2AP1gjZVNrHsdve15g78AZbX
u7PDj6BcxG2VNxL4/yu1JOMrMGpfFTNCZV/yqKNeZG1iixM+GCWEjv780n9Yi0hvaI1o3ixWKS7Z
TEXMZSMFDq1vAgHmp2rEiZjbwU0CTZNMi383Bdt53Zx1y1ATG1owmEdAHr6kWEJM5p/C+Bec8GxM
kgrUvXfzAwOECSBKkM4xxtmZZBDEXjliBYh+KzDtxm5EEEZB3UXlg5HfTWkxrF9YSNUqItF1mzK0
tHqZgnmteMo2zK4Pxyxv6tOBaPERI9B8EZ2W5f7OZ56sH/B1NI3FDuvXt3ajYiRss5fGm0KdPotk
df3J0vcHsgBY9Egp5+VSaUsi6eFd2apt6w52MUxA7SZfotqD5GAFixnGFx1vfTQPNZgLIBBJbs2X
5WifTkoZDN5G+w6jLlLqXOYorS4jvFrWcTgxz9Woe7z8ZStBVFBuvLFyJrjnxPVzjfaLiDlgQ3fN
uoNfbvNsFtLDRj0QKsMfpM4MxqqQ6m21QPYsEG7uLXULwpHRJz6eBoFsxiGRiVLNEQVVE/6atWnS
msQG4bMtIHfYwxAH6NI/QHJNJ7zSK89X4FJBo/B1HOYAEBQ9ONxMIImH27MDip7oFlosNicitiPc
dRH6B98+yciRUaK+caGd/EVhzModat3lQDIBh59EPnn2ZUCw94tUe08X5DVMVF42w8d+JBScDkPw
aUqeT+wbsEXWyaqccohXzx5QTDP0GFUb32otxdBzAmsIzVh86o8vXboH49mfJsDZ39MWzmna5Ypp
fxpaMYz6lJqaSZVGJ1zWO+HBEJ8L6IjdZTXTzJBAQHTJlcya25e3RiX1FNnnIC6QW+wlMIxNzKbN
bTvxu30LmQdKtkUHujIHnu3gi1EHY0YDzBRd39gjG/L9PWv6dw9/dOJUVNYgRkvDbZMjQvcZS/YG
WM9nuSF/49ZxGTsq4LjbDc00HT55ML/8S6932XtVk0NCLO3bhOGcybRZv/EV7kQTkn0AVU+y3itF
X4vbNW91b/9eLdJDtp74gYuMOhGxkdOE5xQWmqK8hkTgkNeAfKQCAa/C1AgZ6rBWeb0DbPnkdM5m
WVBsEyZ4RP9at1MP/yt7Hqac4l6HM4IRNnhcSqlgmrKOUgtVvXY/ijIr4qzSBk1p6YF6B/ksTsKS
v8qFfgufupQXPGdblHZl1ybJiPuZeAdB9zdU/PZIx8W5CarP1qZOvMf/R/Cgc5E6TTiVzO2zsNl5
ir0ElafvtIktbeQWIu4aq/hRzyo7JZ8RDQI34DQRHpKJe9n8KAK6j08aaFPaxnacW0xKYOkPcNpa
+FORBp0+pgxj4PuvORnlEWg2LSfQnKVck2vSp46x2/9uhCJFlmfFCM/wnvlBpm4ki78vquavdNHc
LYDSMAXZSDX/9Wnng74xn75J/c0egM/CgKK+aI1irZJTGz0qv4E7Ngi9l139DV8m71yR8WRL0B/x
mSjFoCos6SukUrlLpaJ64iW1qH3YhjJbzRgV5YWc8V+0027PUKypfs6pzq0v9iZPH7ueGv/nHhNe
zSDT5h/DPp6gUbPLAX9cquaBPuqk16UyzUvOMgZpInulKQMUUnrfYkeJrrygULZ0zs1zg3TnSN1W
dERwqt+n59S130hFS73bUOD4arZRdYU8kpqf3ySDTOtTO242mqGUPjywUu14QB3mMHsK+Ni34ctd
+if6tUoUuZ438kOTgGALjbcHX+KrTsXB9bv9FT/EJ0X6Dbj+m5vAbQ/brylj9t6GrURv/xfAUE8y
H+wrfCXiwSwFZ7mFNUMteiy4lUK3B6VS1Cggsnj7Guernvas0ud3iSpMO3Wz4FUlCWMCinGJNDzx
vuZ3J/SQnfxX1Z/yamqxIJ9uto7KfX2FBqWrsMK7DSQYGQA+BRaGOaKX40WEi8GNiIoBwL5aDcFR
J3PHkIbVWhHG1StEBZEL0JXojbFmkRYDfPIFFaUrRAPrSbNgGMLylU07oMUJrww19TeFuuKVYS7q
9tEbwVz2Tv+cQ/YfjTTNnwWwPSoWkQUyelLaYSvmjPzhkAI71jk/hjJr+hD0PQJXK0WpWRoYK884
+dPTY0z1GgoDhM9qK34ateCcb0xkQhjEPJ4+PqA7wtzpUNzkbrU3lg4uZrDpm2ZUc25LUcrK2DPg
RAclejLgrp9Qi07Rp8ofrOpc/WxH8OePSnvPMl+Pz4HAXRsoz869rTnKSAMKCsLJFKO7/8BmDEWf
xJE/H+H4m2f5wPdGOdxyLdsqsqrhg80xS9tR38kSQurotAb64VrtsR+Xh81ccwbesfDkVNmyTFKQ
l0DgsdRxVFjgKLmnxe2J293dcQfmwXocUVlv9pH/FCi4ieCEOZ10PcowofiDxE5tMQugZuY8bMip
RBZEJc7M1p10DnFmgpN64JwlnptKb4EbT2va0d8ghJYTuHEVFR1kCTfADsHv0V7aopMkugx6QdM3
pWSFjOJKq5KW2YW1f2Nopptg2AU/cAC6zgqo7T5rARVC/ujtEGOvMBAvnvXnIdiISELuKE5SQiXG
djahcaJxQd168AMRvoG8BL46BmKqbv5VP1zxJKRMbNC3fRfU9inoxwxpH0sl2Du9f8a/7K1rmV9l
jqMhkgJ+C7yp6G3yGwLdbLL8WUl0qW9wducaNMjbUkLpgImcgRY6v1TSzFmCmMwUYclv5XzzM+7g
U0tBfOzKSS1qY4qbTjz5CBl5EEZ7zclpO2JAYtOPH+Y86Cw/JuBsFt95dvAQPCScm+IyMcaRExXD
HlWQPXcpqnWYqtGOtMl6YOqm0dQtKCPHTwQ+mXpdIqf6vPO8ssRCTXRhesv+lqJMr4VqbY8WSNTO
bG3wTgM985quubZWrxV1P5krQrp33jSY3X868VLv0jYliXknh3F94IErIGPOC7vB6MYkSxZ/PA+s
gSB84ghnELaP4f+ZsWmtdMR6TC+qN5clnOm+PIRRzJTHkWdaqT5CjVTIoFvg+YDYZiymNEoaWHGl
lK29lijHD7XMSeB5dHT7gM2IkM+bl/bIMWezEvAlCZFGKASJSY90UqTh1+eMQuMo36HT1awcGrY0
9qSdcgweRqc+sLsTE2xTUGmG25A1kM4D0pJ0VNnWmNrxylp3JugsLh5oOlQ/ov7NbNgXnYG7/kSC
By4sjNBxZesGgKK1IMvAr1T1FgOdAYeivCtPsR0FMMG+hGcXA1ef0wEncURkfhY5lBMJJMRmzZR1
i4hQdVohBHn5bcYCpvwV4Ot/+hg7bpDvgoMDUOQynVosckFuIZ3G7dBBRzW6uv8HZqaAyJE9Gdfp
SLkrpnrTNBZDeyBWjsiHVS/Swewz4CUcCEGPsjDueMtqy0XEewNkZzAG8ZMQF+3fAFNcwz68ZWrO
itX9umgf8F6HMSDtCyY19+hcx0jjDFYqLcg+CsnrzH5Q2FqE0osn1kYv/QJYq4h6Qxd/Sp8mlfJk
lFx9tr0L4D83hi4WrPmnwpaMo3JwYN4IWR4BxR499w58Z4lZxj6zieNvzmhQWfn+PLALqmnZ26MC
xj1RvUgCt7UrPdD8F2boZ+0cM84zA/Wj283Xkgb90vQMMhFnn+x20Yhmh9HhpbJwGjysEwMPpFxC
dBqMreV8V+fEowsu5nz9Fu8yQtTBjgtF2hIGvM3cXAIl0cul0czFoiTeBTxz6mdZTgsDtSA7EGz0
NxZ5WidHz84UDKTw8c3JSZY+RB/92ikebexk/XvxXHx/QZ4r4AoMumqD27LrILA+Hewd1fzn0CdF
UhAWMVYbq/P/ZDQQbM6yI7t5qUnb45thtfp5AhuWbFDhaCWdSNpnZHL1t92sa9jO5pzgtIa6CRl2
vQQ8DYgkOKWR9qgh+7ZfKG00iXJqR2xhi9uj0stLH1r3kNFfx9h7iyyRWkw0hq7QBzcP7d84RNNe
8HpBq8BZqpx5ZdTSw7VQtI6n+5yyg8ZooMKURPBOb+4kuv04IV6cvmCsRmyo0OOu/Ge/hXXN3ioy
JW6SK07qJvmIDPPKSvN9jsONMDfIrrU+JhyfyiJV9Vf7OgR2Gw1a5gnjVTQmyMzyWmvuM4lWk/O7
+ogLms2e7d3o/QFnnh/NJJ81GmKMgtFo4tiP3aEjx4qJjhqSllKmR+o084tBjSufnkLLu4lk1QkF
9FcfcbH9Qzzs1/P5R2gYteuJEy0RQK5acH1SKONrX+AWBfRkuIMwbJHrSZ4236Xhs+sguIUl7s/4
5Q0oj/HAvQRpKq5BWKkgPgW6M8QbDx6N/vMtJpSNI0CL72Iyqlz8c2IXId56Diaz468/ZfhSc/5q
p2w8wqjA+u9dRX9HDlc95H3VGCmfMsJjI6IWrl56t97JMpoyOxbQj3YsnpyrXVxBZ473zGWMGPWk
LD383WSId7fGDaamkLkIiisFqmE9AQyHOiqB3on/uIcOQE9XIu7K++kro4eCUfi2HDZFHE0FjlCM
Ab3vGmm+eIDbmkauTbdxMeGUFOHAJzFTGLgT3HxhOyKvTS9sIGK2x3caehfnWoHfH/8HAnkNSK6r
EzF5Johq7+vlK/XcCy11YYiEsQmNBwtyXQfcOBZME3FN/qD1l89R7f5OCrzuAUhEjKkspfGqu+59
JhCGag2NGgyPjVnZWD3yPZuNkrdGdKD60RHfa4QRf47Wrv7r7RtAwxFPmm7y/FvURBJvvXSQud75
fRqt3RXMvz0dSFVw7YeDK+0rnpmkL37AzobURoZFNRYg1MrpXV58t33zTTHUOuVGuowNOReRYqLs
iRTHTBU4/6Izk0l7Tu43z7EWM7s2kQLU3WELyJTkyehxJn5i2zkWVbetMwUx45yf9OXTLfm4381i
/vV8ieva9lSf3e9joi7C4vJoyUPoY/JmQVfd9ydMSKC6nvleRiHwa+KuPI2kR6IX1RrIs5Qm5zTr
FN3+vjaYvCNuDuRlOS6kwXtoQdckedRodg9OLnJioSZwfZCdfrWlzOpxOUGhn9uSCBe3oy6D/cv0
E139lk7rnCQkyAfVptt/E7yrVd3aAKdZ4jp4C3PbFQ5XhXqzR7uv6/0P+NvQVD8vB3Vxnb8J3HAx
TxB7hEUlLfF/7OBztVFXRoNMbTZ7Fuio0BY9OjebV+LS/s6qgcwS+dAEwrrpfgfmnu6lHqGiVUED
cvhrl752jHsm+HWWOH7Ec4zwILG0BUP26s8wi7oNdPRFGmvHsTenpr7iEMlsK+WMx2d4sRf747Hh
QqXybfbwAu0Gd0BCdLf9YRnaylGnRV7tmkRPiJczlrJ8rZhRFiG57iSyvsWcIt2FEUJjM+rT/Cay
X1LC+O+Np43nnNbVyiSDWYIoQpSLMrOY7PHygE8uLxsmI9P1dnmfLBthx3MU/aW3JHiBq3RYla4y
0dHLxRN4D8uJwnuwZE8dJcfwLO3EBeepvMJ0dVwXcjitkJYe6UZTvZYIAR8a6Xd2DNqnqjuDRT0z
vZbtH4GKePM6lh06DqRcJ6TJYlw9nA10X8NicrFaA1aZ6ZWNjFfrrbRzb2JdHNuLUPxpflMGcdjf
tN53NgIq4vdIPoz7PUz34HMfS9RptOn5xBZs1Aal9kq7FlMKHVjsFu/5ukZcvPodiyE19q/hsq7W
b2N5TUZF1V0txMfRv/FYPCPCAhFraFILDppoNXOErh6WEZlRStJyVySJYRaFcgC46/0nB1z7lqLd
pAvB0IeS4dJ5sX/I2yOcwHr9E8qsqaNW7QrY32vhMt4W870IeD1nlsGabqsFKFvWbN3xkaeE1vMj
d18lUpWClqfQt5/+6Fn8GgqBf3TPVOoTTEi0BpHOK8Qo1qq0S5+9VMPXz19UKOlaQ068e9VsKonr
qc9PY28+65rmGQcJDdV9ivI79yI+AglVybH8AZJ0GqyxwrVIASmhjhCr6CcNghvBaw81KP7OAHKr
Rxv1aQFe6AaGGvnNVs2/pHrOHWFMGfvAzJdUFf4WXCXl0TrKU9adEEyYxC9MbKDoDQF51lpzb4Pn
RXekM42LJjlrXVoxU8ir5Ps/LTOrQRCtnrqRUARRU6pbgDmiGIe0AIGvwcHx4f6CcYxvgDoTx1yV
NN6ns/5vaUZ6gNAet5W8nERjsVBTe9NlL341vf77Rj5nyJBLIucdjexk7cpI+sU2UyyK1a6GV9hp
yVnDvt18OTBHxIDa6mXWm7DqR+QsXMZM15nDlvc7g3jOSLIDmB75GTYFYv2JSwsNratrUxkcuf0X
/DrjINiG33DUJIAtiHLEk5Gl/MfCb2L3yKrMenu5Gp7JC1/kdRzU4Uc/tOvbbuh/g72eCNygU7nm
Jcy/68ceiKCTm+lFpafNmO4NrFbzolEwab6iuyU6El0Ic14Exc0UvPfpGDfSphBExYL58vVnYWd9
pR/IFXB/+An4NIVY9owwAHnSmsX0y4KiH7SX/N6L+ui0I5enuDxVBiGr1fvYSUXJVwDskwcI/glD
viNMvd8QbTH+Y0HuoaOh5AxFkdGOPiZw9XBlgLnL/QMNbnHtDsp1O3VQlLAycFrnOUym3wOqCxkp
TR740lzn9dY5uGTp5hAkjDYBP+I/4YFCPJPZKfA/cq4Yib1b42zcC+lBmaQ0HrLqSnESfribqOdj
l0DUajoGS0fAU8jhvjDq6sL/aSXpLK+B/q6u+3fv4s1OvQ5CxKJlw5tj6TQjJPE7X3NW77+Td0TC
MOpsvMGJXFE3pYwvJ4ew9Z9yMNDP+tXnskALr8y3rYZbecZ5LY/yv2KXWaW0GbIEBhvGijzJVKqJ
cWfQtvhd8L0xoX7T8Rbadq2s4mocufK8BzezI2S8ydBqpp2yGOCFWNZYYvoNfGjKXDwNsmr7/vRE
xs+uic6w1IAlnUPzwNO7zUt3GZrJWR2qKbSIQtzRV/2awDUKjkmkK5BUCrWo6XXh0L2RgBMDziS5
5cpHvCKZbO/dUhrMHHbZPMoPIKYEWrUsgsbWc+baVCDg229F0quAK60dUdSwe+ysugHt/I1B4563
XIf/FNJ7wUz0rDJgz/sOnTwvW9Va0uTABRZxikugXf/b+QjU1GK2Ct3NUyCRIdbscMecKWsUDM+d
qr07rdgRxx3k1HztrR8gs0V7ZeXmm3NmdDwLCS6qRP6pWw6iiUuYWnu2oZvHewQ/pVkKYx1ItmNP
k11C9cltq2YYrOqZSARqIuWgsr9j5kkc/PUKws571Nk5PxtuRMOs9Tjta8KXWBZmWYKxpbGlxlbI
PFrRs+Inr3gfxX6Z4wByMPbZ1qj/gdyBgSEFqwe7hwep4lUjNUyLP+MNIYEoXinDURlebi2xG+fb
HOcWRN86c0XQJDlP035+BD/GniHTN59OC/L+bXTQK/o2Kg+u4s+twNe79w1qIM/Pzml9MIlJuGLh
ZeszFKpJa7z+LydQgDCCghc/HeLKYWaH27wcXTOtfOyO+xpuQIMHEZ1oXokVWAjixzRb1fQv69xP
yF5/WtIYB22YoWlRvJC1akjNFuJ68RvJgnsaYMKV0vcM2zPRxRKYvRkFNuVcdRgJaoM9FXeuBYgH
JEcMIkSgOnRD2vP8FHQh1AzAdSoJ46AscMNyrHgRfFovW95oadKKAZkQWbXYus3St84ktviW6K/2
ps4/eFSLaeSHeCN/3l60w2bxoiplMi45DSzWnaAtclYK5R1zFUL/1YRDYJsE7g+1ZM4U0goEhLPz
M9r/2//boYbCmBjNpjJpTT3tWu8R3ND0Ohst8MKdTjKYZqQoHUJhxb3aEeovH2+7b+ACOitVo4L7
Um/40hc3DDzlbGK/xIgs4t1KIwH1j0E8bw+vnWki2tXH0gcxlzHa9r7+vWS2nSIJ3Mz3Hlw1oAXb
Am0g6LjVXpbBgRY9+0qXpc2j+kwKuR2LKRdmtu6NtQJFX7+zJIFD+2JykLWz47U3wBW2FV22hYdT
mn6r2GIyHL0Bu9Ad3d2WYFx5YNRpa8uBitDCHoxutLe6WbT8pGjHH+jHT7rUL8eb/uXmN1MSAf4N
a9Pfzp5pOFszNPMUMB+RVhU2qeNIZ6RLj2r8fuGClkCkpH1hIHL5RrZBkipmdGTN6aM4saGVMosw
8EtTsKtDSKmC8WJZgOCnz5/eEjpK7u7DAwJylREgrtHwogsCdV+k/CtE3cgKgAu8sAG7+My0QtmY
lip96CUvEJownu6qry3CDpT0V7wd7LWhEhGra3nPh5gn5F5jyLAdiRkPncKevZRN6ezaHISrh/NR
jHEK6HCL2B5ctwhL2UXECc9nwsGN4xHwoLXcK38fjNwXQnXyZPGBup914D5QLb+4nSxE6yagHnBK
U3jSC4BTXZX2IW9NL3nYcIcv7ti06U9+Jy6f14s4cTcsSqfU3TQ1agkhJ4b6JK6vcl6Vv3JZB9TE
m/b8dOg5fzgd5yQJwIfAERtZR3MEKNytEdqiKlM+nq96G1zm2Phwki+fRagrmLsUl1x4UBI/an/D
AbI8B0r/cvmlJTorDx36neQrq7BIWfEFKGzP7SzJDFbbXZ8/K/Irk5EQtY3LUZVEKyFwngu+d36r
PTjL60e68UDhT9F9Ux1CbEmhlFiYGxRpQ78GD/8Z5L4QI+WFh5G4+RedRsqGY4dX8ljtmWvgvjbA
2BW3kqSp7EwE3jyIkCyAHYQX5jwk8cZ072FBjSLffEm7XgH9xNM0V3NKnTr3xq9rJKQVQn4uXzKK
8jZrIL+Lui+IJP1PzwI5fbd/OVpPJZwNdNjjEM2sHMresQfRR7eoZUy6X21P3iBA2sDQa56go1gn
20B/qq4QsLpg3gSQ2rgIPGm/oU5kV47NGNJVmIQd2ScRkZKzDZCkELBPBgNfp7VPYEgTAFd6B/hL
hCtx6qhAKJyS/HK8LFC3MBvvFXiYk54uCtlWK2A7Mijv+brfZg6pX9azD/ykEBDXDnoI37rXrVXh
AR/4ZYV4XjoVvPkGdB72/ogaje/LN6UXunZCDa7ORkT9busvDx8GDKBtmPuWxFTnrVH1EZ3DmJKO
RGInaj1+F2xEyylFI2joOZDNijuEH4QComkG9nNXG1RrzXojKQ6nwuxQziFNl+3oF9sm/i0SlVvp
7+Yt2mhT0nrxZGs+Gn2hhe6uMFIodqo4fLI09cM45PMBMPuJD5QLNioUFiOu1dw3sKvPmofzpf8q
k7g3gBgXQjH/Fbv3GrSpdRv3qcH0tF3wpqUk1nRnyE1yC9vPwdRa1slRNQzFlUJo7Oj5Jf0elgpf
/HIlpWsW3slXuGmvDxTcDfrHfAmCV9v2mDcl2akgUvx+thv34ilBSzeOLKi+gvTh8jXa2phCGRdk
xuQQD+/9YmMeOdspi50VTeJF0ortAc4haxVEcDyBzX7idAD7x9shOWeBzF1K6WIyVFf69fhlgRJg
M5fgMUz9D3kFaK3oTPHa6jyXv1B4QllV8QS+vZdQlbQUnDECGgI689CQegq82NywL/GqqRObESwY
18YG6zoXpJtjxQodj+gOl1HRZbI89prdvv1vEmc2y9N/IRCrvS6WFZFqz/SYFwI9+06LFuOxLU84
G4+7KpD4aLNbE2iLuMxuiUvhLPOPWISsdwuqCGt6edOrM6KF3R3RCgVh49gcAEHvzXXR4xV25N/X
oRpcWpVnTNWKFzsoRbV2/XS8LGyuy7ZKy31wWRL91y4zwiMfQYg5MJKAVZlQo7cFF1eGoagCCwk2
iY8aHrB5j6jMXpzQ8S7L7GzxPe/1PuDC5/sfFFiwjX6KJxSvJ9KyBYXmgbcCTvhflGXP75LglvGy
tQp0Nmu7osTV/JjYzEo0WQBy1XQF85WM0VjkOE8YyYqv97L8/KSQrNbqjQUu77diTWvjmW32tLiT
7XE0t3zMcOJYAttNMC94bxcDwOR3ffzgrnkfbdoXm/LNDii4rv145pGZtDIJeedoPDf5w/f/FMJ9
UR5i1mS1cP81SJguaUG+PI2fx9mlOsy5LXVzT2vw41NaGvZOK1pqm4iPud1PzG4tgpFi6Uc/eubA
l5Hh07hJvUvh2YaTSJgizsg6au8Y6knuD+KaIY6bv7qkbii09P6LG3hWoGPG/nojNOGRaUZeHEz4
HEz/8A3jc1rLb44f01SVFnZWjFQlPQHHlDhV7QJWZ9cHWS65vMIjtcxv7l20/RfaxZ1dySYJbB0/
Cm1QSX+548SubTSxGXdrzFhnneZD0ZkgAgvaTeqjhy04L+cpZB4y0QqN0S6T5Gd4QX1ReYePL2YS
oaA9zQ3MfjtmYjumLWKRD+i3zCrduCsUxUVRwtttq1SIBxsobFOva6Xs2/wGFnhVi2YtjRr/l84d
DmSxRA2NTphmr2V0QT1NaxBgSsZ9hRIvUNfvuCuPiwvzgpH2024iNFwnr0uB7997KAn/56yqAKIz
5uO+QmLNlSb5YWeOsulQ6RpGGOr9hT+hFtca1jDTmlovOHS482arcmyQ0WTOmZUFsxSsja5OX2Fg
H1z4CCv9rHKG0+KWRLlZcJUSox77sjEiD8f7PJq0TV/WZDCU/ws1skBxa7HT32YsEdnZV7Jz+ui1
lkNuQpuXOKKE737sogBD+xSjCYkvdjMrctO70+QSP6QnG+Nq32J/Q0Sg8r8UKT0SW00Z4wlDpb1D
jA4svG5jCvucaaBnws85UQmeh/HRhBvKOzKMUwrvXZCmko6LELPiJRQ+H+nwfLAAjI5UW0PMqi6g
/0YxBZMlEC5kMJL2VnIMH9OFV7kWFtUWypCAEAuqxPrvP437YKnG0tGJkKxTgEJoCzlm0+NdNMyJ
7MwsrztSM7LMsp6OSE1W/pVogXJZl1gsgBnNMwAhDLph4N7GyCv9t+8gVWy8rdfzSgOJJfLtvtSG
VWW9nnesIC9YWo14M6pLZKcIflrL8ar7fMw/QUpdbQMoI9ExOOcqVaQNeK6Ra/l+59ixxsjQ5vIz
AoXh4j5whcqAiHRceAUAP0wlRSOLXFa71rIH9dm6DGcUODZpZU46xi/+g59SbTDJLCdElE2H/MPY
S8abX6ghLNJS7AV7WalsbHDjFjmVO0Js3p/n7NHRXWcz2WT5UVIwbiGmQy6RpUWIDWCw2KRcFcs5
UsSk+V2o0MHU+1r2Vbgh37LBDK/GOKVikxt/IkTAYG98hl8K8knGBnfVJN5qKaPWyz2ck+3Eu/MH
277kaRGsYXUDmnTselJgprnhsYKliVisfO/uh4ST47qyha4mkHWAfCe9kXihEiPkioiUTsRmf/IQ
w3J7YBROouri0Scfl0uXpDIDVjA08hGZ1qE4JcmNhnqEmu+AlTB/1QM8krMOOoot6bAvlJgbsav5
5wkOE/NODVH7OFB5MxNcEXs5W7D1BWuSQkGXPAPNUdWy5gc/4I5qv8RhdGYyXDvHnAjGLOqc4Sym
mdvVH5njtu24oHahUcI8ASRDhTjAOl/wKI6DjdxMsOc7kdtCzKMVlCCiCOfkCMqu45cuXLUnh8HY
/tmYOWANAp82awhEjNGZZDnZwI6fotkbIC4o/q1bfNHa7uGCgxDtBJT1Q9ETr4+uI0bUS6XP1s4H
5cDcJ3koomcOnX3PPSNSVE/hog8WLmbdYX5+tGR7S8YKyPbRhoSGgBhh498q+RwAnqZMWb0epLQ0
tgrUeJdZSUxALOqQKFbZCOFD/0auKI2Xmf4Y7OC+UWhC5IOh6FxVRyBQWQ2DQWhA6xaRIP9TBgRc
YuuN7k+VvkasakLJXXLSgiVOPsn7GAL4c5bTotM5zafObo73QvmiskDLBJ2ZDzaDBjT9iC0aBfzW
pcmlxUWx9Ws+AfNS1BKVisHviJQjOfyWeePfCAejoYJ8NkQ1CsDRPF7gd4zp6rhDnkueOY9JDwPn
JhxMqzkPiEOAAeetBWrpX62skbg/dPEvmKKU6TUySSinydk26bixNAIwQ//HmSKJ7A5sLBbAk3Ck
l5leStZVh2n60ORvks49hd8r8cChZB+LQmtnD8VlMW1Ql5NBcjGotEHgFqdwGJId+7pELwhR/4fa
i67w44yzKnDnwPkgWouXuRat165AKqdNZUujd03yrwU7pxfsU4Dm3sIqboSLaR/dqVTD1nY2A7IF
Kr8u0ZNNCCRPY+DwjdkTAv2zJmKok1H190piz/6NFajbsPxB0mLLdTgUw1YESWq4YQylGXKLd66/
qkJi7yXVL2iDM/GYzvykuG0dNjZIa6PKHFF9UJmHh5qqTKkb16cOq1/D1g+xAjZAaFrGkM7zYnCM
enEGp3KYFsPmQYTMQiBAyomtbdEz6t4qhuTJGaECXMxQXmgHgZtWUKHutFh493zRGKVmsDFAtmAJ
HtUA/QKLX+liSJxL4Nh7iNCHOZEEFoH4h6n+39GkHGBge4qEr2YU4EC0JXPCRlY02Z+A3JmWZB/p
R+KsFVkQtayEiqJ/DoEt8nn4AVMpN12c2+x66+hKVtBlTXdnc8ZCMLddxndnLoMjH6wogV+SAtiw
x1eOAgqAOvffTr45lRQ2qoIyexE/usOaGs024f7cbX+K9dLZSfkv+a1hqGyaEmiy+Y3yQ81hout+
HJYO4du7x+ywAWgOO4xsFBT9Xx1eqNpwjnnKZsvQbP7cOP5f0zz38G6vUTE4daiydvX78+S10e0g
3JzsU7/m7BWAWxC+je3pPLSXbt1VdMGezQcVCUxoOM6KxiWYfYptY3oLceO8MqW5DN3EkE9CerL3
z6COxmPtMkgVBvuD3SkcElfVrC0TR+2+rZSIaxWMJdGVu1f6v/EsGgM/QzY4yOJrRjhNNO8u7g3f
OkDDnx/VmF4D5DD55TOdOg5UFxm3t1jHDUbFpNNueNN5z9Y2y7E4jROMeGkoczDyKlxsX8wR7ZFa
d7zVRGZQwKqyvRQu4BF74K9Yy1qsUNYtzH9O1jEu/XnelC0N92a1pMQUlXAhMy/3jdFsoPgv4Ity
3Ahl9UFs5DUCSkAMO72FfmpTDeRSVUXc7dEDfv5qfgU/ycd9fSBDUHNw3TEKCcQH6AFEMRquC5gK
IXiypkMivLhruc5L2nSSrk1QmEKlrOeIKZhtkG1hPZj48+Mlqb9e0cytJEtHONxumLTSJyYui0T7
MxC0z6gGPYkSo8BydxQ58F/HJxVVIgAh/ly4gQxgMVc0NixzRB+3dJUDAIdy1Ocie0fo7ff2ZCDH
hkECiEtWkqqGv7denzsDAZqlRBxcvxKQtcXBXeciexzyz4J2QLl9t24vks7twiRKnqk+cewdOYul
a/pXkHsGd4ZKot1A3h++QPUsz72+PXnRPoghW9zG8LESQNT/iR3s4eMMlrpkJamnE546Q9KFWr8z
B6JcWct5IuDLkEdRGZNFS/+e1TP8Go+ENve+WT4FRSxNSO1oB3WgjThjarMbv0pQF0LRrIR7OKT4
wpYb3IzRQt0i8UTaAtjurL7v63vBihWwQ2R3mCgHWnL0mxrjkGfMuJQDF59MEI3ZqsopEkiGQl7Q
EvWipr+hzwusD6rtbBcKhDpKHNcfZQnMbybpsAbBSgJbHb7d2eYwJ5efwkETaBdEn3BhklsgJuii
fYjbUJkIGC78KKJ3D+AerJ8ObOJw0t/v0nPMgkvggxPZR5lsUw9pQjmweYidNHTil4TUaeEIHO+N
kqmDCofImryE0GBc5lz6vG/WJDDDmdE8a974RPSogz0NzYEZzdZJTmmn4we3e7hlEdQSRjTX0W1w
zZSBge7ioyccLRk2Tsp4PPXG4CqWBdfihJwxzddhLbpNExY0+q4mr0YfaHrjszYTN70XAMMWt40R
mQP+7Qw73YDvY9No9GqCiK8BETi4wbUFK8UYAAa2MsMSDF2TNqz4pKy9gTKlviCrj4LYoVy8XaNC
0zOz4YvAX2kfott3MA11Hoo7vBhQMhhAq9kxXg+zG7kj7XCFkyhjXh3rtW5WtbvAJceHsQlPcCvL
qOA2nMV4W0D682uFSxA24H+OymqA/B0GJH0LjDpmAUQvPBtR9veXG1ws1gWihRHbWDNFOr+kLo4B
2suOHZb1rYsM2JEd4ptsEoVJFLL0rreOaPhDF7WhmqvI+DEW+hRa5RMexUAFDoO7pnCuzXmvvpo1
Vh+eBQo0xAAhShRFMIS7qQngPsGSg20x46V4iqOSa/vHHFbFUHSeueJedPUU+I7AzF8R7mdx7nJV
nEVkca8y9CGPVa0HkUzMcs4skRhslxzkA/rAlNcJjxXTP5De8+ptEoTp5hcYhjjYlMn93kdUIqhE
cJZrFFJODFOHRXwovrNsZNo7HjiPUHG/bTRnUHrBmUnz/TDSyMjDcMA4jNpKYNQZAJMVqvtygUc2
aGRDSLHqIytKoAMhei5ioajcgVuPYsADPMTRcmbTfoQpS2r1X9usRQGzMf8JzDxUNECV0RY1ccsp
uc2rIQ94dPfinsLSOsRM610NpCDzib5vv7ZNJ5kecWyM+dbw9tP0XPCfIVlsKrNRMqaqQaP/9gsg
lEUrLRGBHD4YRuCqglQLooC0fvVw69MCGu9ILSPnjA9bd0wLoZ1L+u1nkCfu7kDhNuqA1QHIsONR
2/2dEpHqAkx/9luQhJKiW8eBqbyBrUA9wNS7UOyPi3/IhUwWEKBGoqUFgFbhq7Et/ERQWWVPzgaK
ZEfVXCYGo8hNsaysNo2lR1bQWWHq9eiyZiPqirM2xooOfb/i3XQrv0YDGwk4XgAg9lJGMNx6J/hR
ceOVnDZXUfO8CyEr+8HvUU9Vhl9H/beeftILGQY3W0cZ8EFFOMO5cMOMW6bqT6R290gTkRBSEPvw
w+88GR4Bmxup3JUOW/ddJ1NvAqMn5MSf3vjk/WzIRLv35EsGFWHn8bYu6tYWVhaLqQ86eCUVQwLy
1/ohQ5aCeBGcVhSFlWqVQ6UfOEFhnSHc4XumYQySvaEtM9Z1gyTHpxfwdIZSrPbIIp3UV+IzlpSn
cMeomaXr/lBbiGDp0UyfIjw4SRLd4urFg6KRtCDHbdNXElScPbu00l6neinLaqB/SJcVMXpS+oaL
7bmqyEgpkyqwaaBoQwlDZgm54+YpzL+/KQsqIy0ITMLuE0S1Ilv40rMUw2cMHqXQ8iJboNlpWlOy
OPcw9hUeFPE4P8YYVkbZApfoSe83AalbL8kXIrutVHRurRnTaXZuhGDhDHbuZd0OzqvKMLmF4vxl
w16beQsapwuVf0/WUv6Whzv4dFQGcX9xzXc7S3TTjLZjj7/ra9Mu56O2xp1jXZFIfz3q/yBdRcIR
dxwKq+y0Lc7+Ns1dmC5CnOKXvRbt77jfHwmk9POrSQADt1rLjCeEWNtfOCFbv/uruVV9dekdOnEP
MKPfJSb54ZdzpCGhOLrRoK0uaJXZyY8vmctLMs8uVyLF+aQpxGKJII4elfTIja5y3lA08ywuJODN
0PpwqWgSWOBnSD4uIblsexVKSuhikm+Q0mYjhUXxbpdDyMiyrs8/TWbboFhfzgi+sPnBlW/ZTZBj
vKkWGLyMUQ/zMgxsf8ViuE2/yHWTK7TGT9M55KTVOXszdp1jNvq27JFpPt3YKPycC2qz6biSeWkx
yb1n54vbilQfPG09jmTBGsZVb24QWU7iNMxo6jTA1aR3MG3WpfWK6qZR0pSCQEDQ/u+P4bREavMT
5BEm+HLFnHSoJ8Z2WoFBVWZzrHVzzsTUqc/sD6CMbytndw0+06znJvMmUDkEDZ50bcQ3VctHMsEQ
alnhPJ3D92wrWcNolGKnKGZFyaa3l0iIll6+dOlw6jJcBGW2+FmGJGBMIeRPnvAacG+Ug58RG8HU
GRooWFXyAWk4kElxmWcsfBlXiG/sOqVhxLRXQsQ56FLvnRfi5prKCitNwv7YovNVBWuXiOpW11oY
5F8A3VPotIyqx5zvGY6TRsjrnO2WVjvjMqRcJbBmVxuefMqiyAXYMRZLRkkkjP2TPwWbsiIGDeRd
n+LLz9uNDxxBUMCs61mRD5DsEdZZEPfYCCYrGnFtxvI/aUpqzriL+Xy6vjBNtW7IKRSqsEgo+Qba
RaGySjjuxgAu3GBF1EiRuE7x1VOaKK3DcEf72OKowwWvfKBMRJfjpUrehjDsbZdEuDBG4lLEeazv
xt45psqnArYHq9nkWe71oIl3+jJpyM0nF1spePKVhARBDJO6W6cpnM7k1gWaugUvdx114dh6Menc
pHkMe72Pc4Wy2Pfz+BxfGCoaobFSEjuTeZyADTrceL2HkHProN9N41NF2Zlh23erdzan6T5O1UQQ
pcboRRSHeMVddOUJxl5QMD/2JS6YQ0y1gihsVxdI3A0rYJ4l1/AZXRr69ncYI/2yhYNEmfcqemGY
ujL56aoTjk66PDAqtty3t2ID6cRowPnNZdM47qUn0i82BfyESmLsI9GLtGqo9GbLnPc1xxZoOUSq
Gah18rE317USw8mRa3U+uklHwXRmS9s6TWiwKc5Kyaf70WbpIE0jHJbK0mbDVIP8RWQm1E1ybjAe
fXVT4H4+J1BQksEmvo1EQbRzijaviksNsRUWV+OBSYajcWrVukuhUvDFtJ1+7a+UvwkbvjaxDnaV
YVmYq57Sb7FzNlZn5QHWEmjHXOwc1UF7hojZC/6xR/RaQxQhILVGZLBlxkobtbkQ/j9dMObDynp/
MmMrh+4hzIuHToZelA+QGhxdTE/JmH/Xu262ZcAeav3cN6u4m9RX41lh/CuyQh2p89YZRhS0OHkR
IPyGD/ypaw4aG8nDAoIpUEkrV5sjRLtJA0QwhWgVUSpqkKncQf4+TGKoYJCXMM37YIRFuE8w62+c
VU6HpQKJChyXdoSErCMuVAZ7ta01lSDFolhLESEkhAPQMPa4/Fu2U6NMk1BzW5Rd4YlK+oGrS0uZ
4rHghFYc5uCaQ0f4YQij8tm7KxlRZY+CYMk/WxF4NTc95Z7u3OYEZ0EdWXGnFqaao0UEMAeTtN+1
BJ+28zidalEOctEJYLFNxhB2bCgxnIjjMnKKObEEJNhULw9beSkMVBPXsh60RK/QpoLUbSXZm5Jq
qokYTtK5RT5hi3adu8GymlCEQ4Y8PJh/HjP/+YcDt8aAMaROARFWlPERfr4UQHUiezHCFXrNhP3n
ByEJGl2x9aTDisiw+aNnE8gC3BW/gZkBCZdv6xDtt6SVrn3d0Md8sj+p9rfbhO5zTTzDGURbdGDD
YNgQKfKdN8jHykMuntSqFvWu3bbjFVd+DeSmY8zPerP8ADDCKNjVoEjSnTMCrPjxE35VdHGvUk3O
4zFDcG4H2qyXwxkcXJ5vHnYrYnLS7X8wlS35X40s8MTIt6FUqd5Hcwbv4YRzi/JyoWl7bmFbOktT
PzASw5dgPwQMh27bZ/4bMwQJYKkwHruQkSFXNbGiPZ9GS6RY8ee7mWpf8t+ZQGLFq9Z2yps1uBjU
hfd/hD65sXRLhC4M1Krf+PTAoaWuqIZ/yFkjqs+hH4JtqoJdPqWulXeiXDV9K1UbqDlp+e2dc+5n
hpU38HfpRBguwfeKOWgDkuHCqh9TcIxMboAIfJieKFzHoMDjKJk1Dbv4k52e9IufPL56QM+qZkKF
42WYkg6myHpT1Ft1niZpR0ibTtYi9VbuspW2DFzo/ShiKhu+qAx4phXNFpW3iNxKOGGg6wBA06RT
6jtyniSK2ROJl5TuJyCckF0Z8Bj411LB71fZ7xR6HOdAq9J82MsXqhZD8Z/UTJFUqG/RQb+9hRCE
i4dOgPvMptk310HoFswcn3hWic1tXuN7LyH8ZPLUEQjMFeciy9gcr9cZaHckK3gejBuYJBZqRYxc
9hqE+YFvtgZZFAGEWmgRxq8ItV5w8r+RKypkwJaofR162SmBk+IXKdg1hKWPlDhPzyFLysP+86PN
I9jFteFQjKAVRqM++n4VoTTuhB14M9nXCI+RLFryu7wdhfT2HCuzxBxQuP7c+4jYY2zxedK9xbXq
pkreBSd3EJJpevuofvRjqwdF2TIRDfepYaEog9P5REafz8zpkFwhPJtThNCcrEzq3yr++FnT3S2c
9ElOc5EvgMTyEbrpwBWaUX6Wqi15tBfNM5sOMn2cRl6oaT24xvhii7GPx5eLXo+cRN6+lbi7DkRb
0hOfCtyU7D00U0lVvyNU9Mw7XM4svsoUtBQkjvIINApOjNbx5ZFTgAVv1qKt0W+3A2LTbB/azjaa
jLKRHtfLpgCVXlUUbxPhNTrS+hdwLeOkksNDTTJbBb4xEVRD+8rIokbXfMkBB4WpJAcSJBzDt/+N
nQHerm9dUDQ8oAQL89yT7DRqrt3qca977TWAlJ+ii4cwfyaFtw4zVPlVN+Zv5axY+KBz0f34ANVe
tpi1KmTz5J9eBTRxckpczZWElkBZbJTeoGQa29txscvNf6RC3hli3pZohB/PBjW8fp/6MpFN+fQE
IKmHKGTZZjbV0GX+cKu01S5x6zXZS+sqnDQI/cGXjPfSZVjbg/LRs84mZGiA9ImYLqTR8CD36O6N
ttQcvWoytLViMnrxCnnYX1euRZpiaJZRDbwjoU7eTWRkcTK6nMkVTCkelzlGHxjBhQF24IosS0Ii
rGBLO3mnDiYWe92WlqnMoWZjm2Mc+c76SciYChsDMV4bf+iPH4+LUt4E2g/55RrXDvSAlOql+GNR
NFkcu0tcOXaQGXMi79wjU1r09ScTBXGfzXYabhgiAnOIGowj24aVLKatcLPAbNwTm0mldjMs98F8
slrVzJ7HuRkTklS51+FU/0ahOUouMCSwj8MxKM3M4X6uVjQy4AKiRhvAd/ZioPZNrx3t3uDgUC2r
jkDGkupLz9abCrOUA1JKgcRvUEH2yLdgja4v9J1DBmmLo7/YG7zHySJygYZIFjvjYuu6+Fj1FBto
Tqao7WoMcDHVTc29C0DnOeZqEBL2TlvpWf/tvGCujN2q3ERFHwc2OVL+fGYCF86D5IL7043A7Akm
+VQCSEKzv1K0ccMk19yWmPHDtQ+/b7jZjBEa3tXGrD2G6CYXH5XJ9CnsAL6oi8Wp/SuwIM9ye01A
tTKsZSJkQJ2QRKqNNG/gIv5gXR3cBVhWLjPVFR3xA81i5aGfIrEKhjx7tPxNRhb9fVt6mPWcZj7p
4HCd765p0Oar/iIFXrDYc4Lx2K2r25bZ2RGyJ00wNc2zFLC8G0/pUEbKhPyYYOpkKZCOwHu/oR/j
wJmwEIlAwurEPflY+jqK57kyeI9q3zQ7FD+HRjXHqscDNu3R++2heXbTDNSZRaRCzQm77eE9kGpa
ULmAM2sK0S3JCiR4OofZRhhblqZ957GnizH+62XlWMKgvoPoQ8OTuWoMuwRxk4SURQcXDvIgfFnS
kW5Pe5tVototA7xus+P7fglOk4vL2awbnc+DDUncwY4MrX7QL3aHLAjKQzHJBbeYxG5ncOFYnzBT
xyk/KARpNX8tG1JgU8VourtzA5WZUHiRq8Z4GAIDMFotm48t1ymq6uoJUebaO0wEi3Ph4NcOfh9M
8mPnur62iOpCTeP5N3RBjGsVjQRxAAb7N1aZJr2+IBmh9L3TIkltQrUG8Yv6I5KPh3eFddY5xr1/
46mnzAMVLRijphMQzJgTzz7c5lpeqpP5LRlfXzuTtyiRT9KtYLnGtUNWyOBOTNff1mqk1MJPHL4l
wT3daB9sGuBTSUDBDzdD6fgvjgYiVJoqCJ0BSkgDVkHYXLwj6kjvfpS3MlYIKaoGOSoYIPZrbpUw
gVoYeKTkjBywTCduFtbntCgLO79ZtOe+xgM90UlewxjS8wgCYD/HnCRfjHI4ccOm/lSUja56+Uqp
DC0fnubMtVMeOCuowflXLHFL5QL3FvhqVCl1bOs3ZB2rU/7v1xHPB7TLDI/Dt2G9XANAM7NPBkQa
30NoVmaLfyHe+tyyK+OOgF2NCOYNCr9vJJmrHES6fu7msjg+aku2x8ujHKYU/1WtB5acPY/U9Lfq
TkFRKaFSz/8NuEeIi5TqL/ssO+YQK8SZd3Hdshz5N+Q5oS6BHYV3OM9PmdL87NvG0wGlqLTIRr0E
zYT9hcWOb7I67oWvHeGLkMSSkwFu0ZagJBZRIjt/ED4mHdnuSiQob03wvUhJCwf4rW81B1vDabN1
8xJ9bQtOgwG4yXct8LmYAesBerXbRVRcl5gZD01pOjMbtPDXcRdAGIVWJxvAxayNBdbZPGCPeq+y
NaDSPAqXHCD/NgsdsfPTBtKRCjCLZ5iXBlx00045XDYwyv2hplg3Y+HeNzwJql71U51adH+1Bbr8
isduu4uHZ34YbCYTwkO6LtTFnKxug3mBTAtrLPgNr8zI6VPOWWfKX1jh8DoWsvBIgPHAPAclMg0I
1392zB8VtZTYkHYvne9GeQUf+Cv6F/f3M8ybrq9NvQsaceNwwgXDuwXONIoRyd5cXXMGNqkcGGvb
Ry1m4oBeAtG8H2BBV8K4IJX6IR86kr3RYeMy92/q2da7fYRBuBeSifKOulwaf81PGe1cXdQWKcD6
VA5M79SXMF3H9GhH4yI43OSeytlSdcQFcStN6hfrLVIKOrWmPpPB4dOk7TTxsyvRBePDmr1www/D
YWDHvDvw6UpTRVf66PWTqkna3gN7TiaOPzPDOHAe2l7Guj+07oyiwDDNgpAKPVo+vqjOyQ/ziwfh
L7hTjdGqlC98DSsmikSKQnHk5rnz95P4L0ooO5qExWgNMczpjR68rxYiHRF0YkptBec4tmCrYnyO
XlgIDIjQhV5no7gmEJ7DVQY+7uRpNo+HwcMvSU69XkOYQyaCiEimCiaw/Q7831f8Z3/clrN8XdMR
RVjU8MtOMTeqWQm51hcMlfK7IxiYxwBBWVDTYAYtEkeYwu2PyQYfvX0SnERNRGHy5RkSC0eKqvTA
wo6ojqwFqP0eTCMNZ+igvUOpO6CJKEOlXbVEmf0YIp7HyAU+sPIDHv+ovr1+dXNL+UX2P8x0dEKD
Pcm+ZkOpl2TtxTuntUbZTVFbkWRuIzGNxjYAGPTHThyZCZVwdBk1PhxamWw2gy0dAuHWg7lI1fyP
3DSDrC7ODMufihKl5bHUbW/6b4pCb3uvJ9W9Ne67CpQP0MHTALA4RnnwI2hA1zMYXBAG3SJPtgBV
FFs2MADF1sKnpy4W7b2eELNivuc5m1vAsJwJf+ncOPE12YfQxu23Y0imVTJPQxa6UQ6zz38LBac+
wGIFcaje4nQWA8GFZj1hFffmMiIfxMPz931+xRMizcHtExV8EJ3NJYaVz3rt+3AxZi0Wq2cmqPcp
Lf2sGgRFyKkuvEMkozFGpFpk+9+IMqxuuG5b1LrQ3IaaKy0FFvpjEeQCun6LHuxiYCzQVIlnsCY3
Abdp8AV1phsFutgbFlIUBUk302Um8ygx31kvrRLnDiIXGXvMT8qA9PkAqXL47wH7Z3KiEfpMRCnB
X7V2cZYTE5A+EPodyRo0T5CiRAHYvYGAmiehUCtzaZK0jY5n12oUCOGOC22MDt+rexFq704ORVzp
sOVtDTlK6tB06qWb2jOfPha9jI1ce9RH9qamRSp++oaqeRwSEahvaQ0YL8vlaLcmblA4iQz9Iy06
JRhft0ewt5IvJeTBRMa1FlUzzSoiqLEsG3Ulou0nVWT2CC9Wt0ib6Kjho9jBa0CNUKIhZUgYCG6+
SFnzsqcFtqxZoLUy5tX6I9aDdLhujwkp9WRd2mgAfkcjQNWAR6RisRv9iFe3g2i3Oj04kTsfqzAK
+EJRbpXINTZjbnqI8GmfCojpNf44rxR53vzekW6u+hOsasGr+xl8MDXQ/asumWR1bnbLckycF7ms
ONAPMUpUxGkSNxPlfULfLPSZ/Il1Sngr+S1l+B4SaNkzbuy8bjUANZYy5USIQ8i707uCE8IWeGAO
avyZTHfUPwlNvf1KUfG5cOhnjXs2ECuvJRnkJNfQLu9m1OdoI93/kYxc/vKDkUHT7cQ8lfmk7NHr
j22RDezn8rSrhypYDvy8FogpX1rpTf+SLTTqT+s1LHx0biRsumD4gcyoRC2OpMrBM07Dh3ghiNTE
BbkfqCXVwkFZsbY6BoCxCNMp7o1Fj02Hy/cdNDVoam5JU9Xm1Wr0s4oWamJGPHWVrJaqo4QhASz/
C00U45xDJeKNzS4ZnW/ctbE+AX65JWff1VRVL/bRzbiFNNChIPAMq83LXWdMRNhCJlxyVwjtS3dl
kYsUVFSZjm81hMU4UXSTHcH0totguEFUZpgL5PQvPU85BHZcX/1IOVUKjiPujST8er2UJ6EHmqx/
yXFt/+2oxNRTB34t/tInICP10xzmf2+jUkCaVDYNe5Iw3Kl1/WIygZbLpGA2Uvzoc/VxcaGYwTH9
dw07HmgtIX+alw4r6PIDFkhBlHX+q8FZy9suptd5dHdVsLdcgNtAFF7VyU0TvmFCz5V3PE7CFcVL
Ltl7JvwDqBskZRERmJD/lO6R6LSowBSvdUR8okiActD7NwzY7PbFLb7Z0yKFBRYwO8ZFGR+KB3CU
m2R4IMkEVs/WkcvgCWyhI8mgtm7iFEm+uGb3qcAp8ODeQTfuX0OyuBNFD2j1qHDOMvXuWrSkReHU
h26McxyEjKoVePF3yn1wCpZxaGWhU3CzxHwAH/CP5/UJJo6LS6owQlA7QFLfFX/aGye7Rtimb5NK
yd5rRmJeve587E0YZS1dogTs3jihlZ7jFZoWJBsF4tBCe4hTR8f7VXutUiiVmN1OTr9fA/yL9ozp
502jsDWTzGHj0BoJUBtY8nA/64xUIac3NMwyf6txFaCm6S4RgysuaybtKGDIcnBxDDL0jN++/Akp
bwRM6i9TAZTV2yc1+pACcNtzFux3wT/z7eIw5MeX5NQJwXLRCAqzOAa/OCvB0USbkCNfbZa5awcq
R/FGh+SjwXsRVVdBZut2aqa/PfG8YpjlrlWHbDrvpq2jyHnFS3h80n54xlLhlAVC3aMupmYYY418
oM/hZOm7EM1HZ36wopUh+2SN2tajSrI6VDcTu2WFuAj+tMCIq39SEP9rNDPoc/7c0ZmHlA6BWIBP
5zOHd4XgMAmx8vwt886JwBdro/9W6UFadOwYr9n8L7i5ebRduJLZDJFJNlP3iKMZ7GbBOBpysvsW
FD8k0dqOLo68V6ESQtIm/il3l84WKUejwaNthSpXThdt1hPq012GZbav8pC2rYgjXH0dw/9WjR1Z
yZZDFGwMNFjCbb1t0BaRyl5HagdMzyNsEIHKEVRBpvE/uMc8kN72sgw4rWFl4WPjQm+pWomqtBwu
WOjvqB5JHLszJg5rdOgfrETVncBeiKGEoyHy7TyqS/WWoAcjdwOESIKoNBaT/jZjCa71lMPPlDuO
O+aP3+jmqSd88KEnblDX6O8oGf3YtQrXUEFSErshuzlHTPKLgJ9DERKH1JxyvgTCS9NbYgkP2KlZ
ia1qUhdAIi9l7cQdQ7ZQb64g691Myz/ce7JH2G78ZkdK7VuRfF9p4CIFOZARZqRpeQpza1sK4I+K
YsFIIyDw+M84xRFn6GBNF+cAsrpc9i2KkDtHyruil9WbTPW6uq9ynw2I16ym5mKqLdcA5imgpVml
U1O5OQIT40Rzi29esD6OvkfL+Wy2Qf4edZ1CRdpp9JzP92rg9iwApS43VvdWDYzu2Z3gnBMun2nN
nWmW88s15wEsoB6BEwaJU5/O6GqMDkQoGXdgXY1ulB4Lh66uEFGT06IumTqS9kxfxcdFyBBMqgri
GQdwb/UkUbXGmtUBbZ5Q6Wlu+ve5QBzx8ySz5fAP8e035lVDV+iEiSayIxZA68xVoHhzLbDQoAJb
pFjcoCAj0A4dxR4RnF6R2Neo4GVZ609Hs5Hu7MEyzG/bI6i0icGYNmaAxOT0T5Um+q+AgEwc4ezj
axT1sL+CRSkCKekzVENDiuU6itkqEyTcItsZfz/E8WLBepM3pRykWk08L65VIy8SY6eLm++3VJ1z
ZBDFLmk3Rm6lA/AJUs+Sy1dmBw5TD+GoofvPtD2NxwsgjJi305xv8X9mOsENfN/hVCVmn3vryuzC
9Tt9kdoIEJOi8lE0X1Jo/swdSsXCpx0msQOeacwn3H3U5c0leCUGwG2qA2G/AmBxRKtshHszimNi
LPXAE/8H9fKAX+zaq7bOAZUJ8cbF7F4/D0dQkOdU1zAGUse3PxzGcD17eLHROBlSnMkqxBDsffmA
scjR3tTnp/xAv5iAOH9Lwua4PtzfR/le954W7kT9GUuDActJ7lj5Ab41cfQfyQJBmFMW5Z43y7Cf
NwQ6nXPZ4oLYCUZBCTUtu56Ea3FVxXrafgetPCgEQMiBHjDVEzUDs6EtP48JLuZJ7XAOWHNyvQkw
gXZ8Q6KEsRh0IoAr5jnp98Qnl9Ll2Z8Du6IBAqp6DJGg1ScV1MvGxB40fdr5hMop3sPBii+siXka
ZCemOylPK//VbnbeAH/8HlgwUFCWznITQusZIaqDE2yC/atEeIZelCpaXNqfZJHFhYqNNHNyWX6p
oCiSO9N1CaGz7QV/1Ut3JSy9SEFpuGz0PahRoAH42vmJAG693MQNdjvGSmOYlxqsCiVwa/ksNENo
ToVjIFAMMxR6gvro/ftypplpJbwi0Nlad1Oc92tTHAr/jminqAu3O1Xef0hadEq+H7sQOJSZbKq5
sP+cunvsKHhFHeqdoXZiAh4vFesBwom6MeXLerUGbxvPgG/xJawhB9f6033J8T62i8X7mGhJXWb0
9eDmZD0psUXURDCAi++g6NzM/aGtDFKpzH+eQhnNDHUXG7gYN0VfWbn3Uv/pjjLvyYvZTNWeHJ+z
u+1XipvwKelbIQxHklgAaKG+ZeGJ//+8nzf7suidRajLItMx6OMNvqBU06g/mERp2ccSDvgyanZE
OMaN56Gz4M3QI1Gmq74Qe2mYX7aLGXUxhhv4yhd2GWGwo2FpSoEVVRl4X/dbT1OeXJUMRbWL1gKH
8dr+WlE51eDbRiBHL490k8vdAmnFnkhvF7rDXsqKtiteVDCasTntByhyWm9tZZvp6YWBRpbODrHv
nZplq2vsupcLLwTm87JHxzQ3bGg+YRS/W0fs+ymvMNog7y0LG9/6xpzNVYUeEKFJe3y06D4L7MhR
t5bQkQhtGpKFex7BYl9rFt2mMz9bqxlWysTHf6tIsqumhTs/w70MP/LqqMGXegoJuZbARdlgTabh
DxRUpuMKjy7nln4tdba64kA5eg6gnLIx3SdTDCexkuiPmsO4L1BnGqlthyPVXTnuVownWuOv3F1M
HBbYwfmhAHKt3LoIxc32t6pXdiGpjpr0fifo+ahqT9esiqRqE7Mmlui8wbdnNayuNeZ+AAtdcUQU
0i9nK+syIVAI8atUXsb20INnMX0QLQbWd3gbPNQTBfN6pAV/r/1uX+xeYa43TC8cftu/xRpRzkI9
Rd3VxYexL/AJDR6A3vq/vH6t8qEhEl+4siTtu1JCIpKk58BlLjULgIZAkIvbyeRXIEdY/RHgrmrS
LmPItw8GrbGwZ+bloOyN3yeQlGZ0l0lm4aoI1HIEwFjkQB0cgGzLnMUw1e2A/fMCdTJ5w35P6EGP
Vu8Rgh0iOWEqLi3qyXCBSFU6KKCJqmUJlmgRdadDgD57R4r3AuvdzB+8GBTaSUl1rM9PqZZCmRNm
u6ADR9ginKIKf+1PZ6RcpUsPPynniX91L5GLxl8iRfXdwXcvQeTI09POineAaSj00ICeUJ3iD0tk
jHPvZtROP0Xko/xhtZUNPgTzGEawQj4ggHLYKIug3uLjiTUuIeaX1+fGXyr3MRdOn59l1lzKU4L/
xbc1AisZVG0R+b2Adg2LgfH+VeVAW1L29JDvlikmMlTbpKzloHfBAwAPLRxo3SSNEBkjXxPQuK82
obozaqcdDDKlAHWvMeJIFLkgVjGWpCQHcblOOb8rAcSz+UG/G21JvNTq+Zp+C2t/NjqzhVXwHiGj
qfI5LrGjn5lBmWo0NCVkj4FPGpsJFQ/lg0bQFYcFvUsJ5W3sLFEpvqIx1KCv+iYFYVaRRRuW5UJS
/KobIYlXUEFI+aHkTLN/+DIqIgWfRwQPcOIRCGIPR4j6wO0+avhjzMRCkV0EYlDjdS3jmBYzeYWX
Yy0HyYXGI3pig7JTRwxCAgI21CRK05+lAnPNl7OrhGWTR9YvPjTzvQXVgvCInR8FVTw/TAJ8fuBv
ml+hENqEfFZP7q58FnC+V1GsIlUa33ytcGYtmSaJ8d1l+mZ3IFYpIVQB7Reu01zg4P54ryN/lZNu
jBwETiGoBK4jt+0HOTKWBrAUiwogLnBFX1hozGN850F7MRc/gtjH3jDn2pgTRLzTHLEkgyEEWEj4
hKMexV5GIY/cACiR5+txLL7JKf07EeL4KENLnBippnMYbvsQ0jg7PUXQhZjW0tGOROomyT3npniW
8vddPARUYreHfoUk0SvOtkLUbE4ELkmCgR145L69xec8eQRF9+/qvS7eu3yu4iDwTbtsJGmBIVI8
h6Em8CN9+ZOgr0nzpEINcsUeANRMEH+U2CSf/r38JAw8ASHwo92Bt2cHp/uHhF8RMcdTIv61oACK
DaYZFiaJOcXkM5WvP5qYhaA7+7wFEhPVAw6rt5WcJrI5g0qheTM4fZNzXFI9VWP1eIEAuYJltZVT
jwoosfl8KNOsPbme1VD4Q7Wh/kdhhJ5Sy4gROwHOGMxUo1YDBIR5yGakXh/LR3r/9cCJX1UFxw4N
WtSBhjWoQc5z4oAPjuMQ0fEwODEybk32hd9z7Qypk194368hgRL2plA5tK22wFjWkvc2774m070t
V2GOD278erdy/vi4huye1C/X7d26txhCspX+7VCz/isXRzNUYWr0J5s+lTHvx7yTnXU4hjcGlwUq
1FwzJS1uWIJpyW/LXgeTvgY1/WIMnP2CJXARXYeHMYno48ZuWgzb6S8hmGNkFkQQMoe23c7vT6So
hpChcyeXzHfGPU+0Ke8kgaH7rAXwPsACof5TiCgkKsYNlwGkhqFnQdzEqxOA9J52t/Ts+iQA0mpR
s1qhs3KznYsfAakTIKHwD35ZckaCTJ0Qz0mFcWB5FttfQaB1bK127FFgAFX+OKYa9ufaN7/KFFDE
iSFgX3Y9EyLr+2FUwysKzWS/pJszFjWMEeX7Ymv/bfperP754o8xu67Knwt6r0Li1M2ZnGYu6EDD
164/q8uUFGOsKVpAMX7tPiyOgpMXx8/W212HLXgzuB/b/h+wxpKRB/mToL7oRHUQv5UFWq5WxTT+
gPz3SkYDPhxenwfyrbhJuiOCytYFqgmu19zyRpsRydEbsPkYFlVZmKaqwBeK0dSt6i93piPcLTG5
FeQk1fmyJn4RacgJZ+7IeP5a9uzOmbhLy96cPSKUAAX6xcXmWgRrvrSiv2UTebJ9hB+w0L9SMUw0
7JbMlsBsOs/odnTH3OhOsD3r3zqSciD6g1F6B9rhi/f6G0/EQqBuCfM4CgXZ6b8hcl+2KveYzvg+
VOb8ar4ETgnc6S3VcKG1l3pfF5sPaCZLJbIRbZsLhrjuOBrgKe7eOdRn7hbux8bpYle3iGajzYt0
bidR9+WzGw4HOKrqznyAGqOE6IHWi8C2I1Pyekvk/Qyvg/CJ2XcE/+/Yb7kFlBhOlfQg9ZS63BzG
Jxe1Acnk7DpXRC01OH2NJgE/gPQuKrQskuW2BsmknQbFf/ReZ+TkwMNzumVk/Qy6D651yHbPom41
jip/K3xhQ4Y6Pn9/qVNNsUFSt9VLl4jipjLLuCqFcPYPBlDfAwdMjJGCXm4NER+k7qNMJs5hh9sB
K5+ORJTTWbhvx1oC+jpEej31zboXmbXoWcoCiiIvNRxg5+eV+dyL6JPFjkKF1KSX8LpGKA9sQLdk
hhfa9WpcgUF3uGv5Zb5Ex0r/NleOP6tOBFpVyUq9xE0L6Gih7f9hgTPmsE9DyglpPLLuPEs1dCyx
xUTk782nwuFCnpf9FOJAFyN9ohV+jwFa8rDEqzroSco2WPkLuYk8lV/xISagIR6bLh8R2sqG5SxZ
9ixx0Ks8iOLcA5mRtOlvMI1mpqPBvW76eEpLRl0NSkQvk2BRrTbDIlk4Qd2euN6dOrFDK0wt68db
c5MIHjIiLoCMN3IHolHnCMPjsyAET/Q8oP8knTfxUyrSzO/o8wJ6xhhUqKILy1FCvN2UTlEYSpJN
Y1OHJPjLxGnpkn7S5SgL4A6c2ye0BoVQ5QsmwQ6F8wI83hlIYmGkt7HWJk/81wBLeJ5Fcwx5g4FE
tcCShHEr5Xndz1rcg1wwZEPioXZsUvG7VpCWqpq9a8jU1xhC3G1vUgPQQluWxbxai483Z46kiWRP
DOB/pgUHU/18+CNbIT2WzEkl4AoVl/S6sThtiy69r9m2ILLuikvn8a7ngOL4JYCI1wxHNnsICJpZ
HlKPTZijuq75sUqu1K6lLZ+OEj5Y8V9GGmjhxkubKANvBh6V6GaOoasZ5joSOew+AX1Uo8X5G0pj
HlpmfWMOfZmuaD0K+gVm5bieR0pCxfOnUtp/WZ7IAvpcowEZhCYqMtpLUXkTnnY/VHLssjHa+wCC
k9Q3WVWdOaHRPN/BhcIFSdqPSH8F3kCFzntpuZ1cES36nWg/xHyj0DyTp4eh+piVh+XPSDu+exRx
+8RVzgaRtCM5jI7tLwvBP6bSO7UA9wgIwGL1M50SHv64FDuuxe/DI3UxljGOeexxYoCfv/z++9jy
8l6uHYXAtZnzv61OTZ6fJbQi5o8CxSD0hkkcwx4jZ+qHQ6ld2FQRDmGA5psyoRfZlrqCbeFXJ6Zg
WHoA+bx0j8zajJFBGStD4LYEZwI2n908jawUrUbkmQZs128bdrn8SR115VADNSK2YTSxEcyA0nsc
OWcNR2DRrkxWR3BwLIx7/uVyiD+RI6NyNxhtqRNZ5kx38qAizSH/livdNsBGun4t1n/PWN539X/G
o+dSyVG3Scqwfj2H2EHkf+doYys6xVz+twp7NXiwHZPblomvi2hNd6uSocWzsS1HMFc7AkO1H7HU
mw5ARQljilSEAgz5gwNq4v5QtDhQgf6ZeaAgRZXalRWlWbbdip61Kj70f77n0Hty5kRMlOZZ6LAp
ugK5CBf5gYnSWDVrrIfDCqm2+i6Vo90yAOsZonun9H5sPEwxMQ0Qghlu/eintftUUhoAdrY6t2Eg
TxmTEU/wBQsNn9iWkccYROpa0WaiV9IKPHnX/gqasVAtEl+IbmozehOMh4J+dv9eM96ATmfY4yJF
P2c6WeSgkVEVeaaCe7Vc9CDJdJuxhhRDMCTWlqJ8Q4ZVAlyVhzW366+SNqMe5W4DcZGgcJVJT7xJ
KJcI8md852CJr8wYjDd16h21VAVsQDcWZ2exXQZPgN04M0vNZA1DBzMQiaR0KEQNFgfHnG4Q65B3
m/9nMGjWXHpJsm0NWsb09gEH4Zn+J2URLuklJnlGPXKjWZdtm3tAyEyvUZWPwYyxKA/S+jqNHOR3
0wYaAB1fZsEEq6Fwl40lIpsFVDQs/NHHRDZyWrLrVe1X+TzafxVMCAWDGSNf7+opyAuonHk5WJ96
NNcNvrW7p7eGDLh80rqNsSb5Y8UI85LCYVGWokYHjRJBczrnaDT0xF3hQlTIgws3J8pDASTNDNRX
mcRu68Cz4FmM+nPux7AoLXUF/TWeb6ZxDB2zl+RZv2SV6T6ekSDWMuJWcwi+dtvK/6EAodq5/HgV
4cWcj1DO7xVBtkX94GZV29j2vEA7Ys97ardS83sV22C+P0sHZ0Q0WuW5Q+BYJGiBI2ST//7MblD+
POQZTpQ8tTUOoP5RY+9vOq6F4DW/pSwigfJ6KrcZjSIYwn8PG9nDbR4meJCEUSRM+fPKoUI2BMe8
qODnkAmqAGrgKAxxTjxqDd+mcdG2culQ2VaV0+iy62YhCB7RL18OU2+bHtiRQbuv6/Yc293WfP60
63VN1Sdfwz3qq8xZL3iHK57/DY36QGdco+a56AicA0P2FQwk2L8RCsASPEdN9N8TG/xFtKZfeWQB
XRI4vwSU41kH+jUIcQXOpQx0edKCYcr1a+Px3z5xrMXledfofpicb0y4YwesuuBNRE78358qONyi
G22yvpDakv9jLlTCAeJ20TqJl59zyp3AadzPbCoTNxyhQS+b8nfht+cAT/g1LOEJifECHSZ8coI3
S5KlS8je4W0T7PbafPBGdNyCAFdZgEd00Cful6PZLqqF+uWJgxtH3SN7Gw/kBsepd674pp5gcGoQ
nj4DfERBoA8FVHuUggWJKjy4U2GDX7fC4wK7MPwg4dnnnOxhoUSJ2Fg6MqFruAnrnChBB/8vMmD6
+SRnv0ZRzRtmWlQSEXysFTMG4DgnBjrXVMWoF6RpUUuMixuYCnrqafH30Q0tnWG4yttIFYICpueu
W4w4ymu1DfF2rZFAux7iMh4NWa3EJoMckLIEbTf9QoVVo9HsNFMjblNsYtjMWqngC8Hq41RqdSX0
9PozAcERxudx7TEJ2qUd7j8W96bbSqxPXRawCpfVS/P2AYWvSWTjGoxe3iM9W9kCNvH7CAiET4S4
shxyO4E3SWDKFKkWDqKDGe6wcM2fDaM7b85cA3nOpSKsqW+E4zuVUJr+ANtdasep4GZ96+jXI1dz
llNkCdkIlsBWcrM0Ns1rFIX8ENGzv4h6EDtuLFWctJ+WDhoDzYejPGMRp7yIj6DknNXcovGUBrk5
yPP4J+F16XNpySowkp6QM8Kre4eUvmv1hsFdww8K/UPscIz05Iv2HhVxqqgkQQdhv4xboyeKFiSS
cddFUsRg4QPStV/lii/tIMVp9zxje57qTFV8wqnFG0TbZHsVHaMJ1g722eoA2zHrgl6kYQM5VWUO
UoCIfao+jEvHEmW9TTLJRp3GdqLXz5HDZpkHdbOtnV842DaW8RBA6u0i3QpN407N1lPXWEltfKI5
MtyQooD0WPQ6V6iXfnJoJCme3VAWyyTlBkiLNJapAqbUQa5Cv7cil1MWpJeM9k+j+sc82LP4e667
HzsWjspfkswRxZZiNoUU1UolHCk+78iA0qgHAdXrxCWp/Gs1ZmgatYTPDXoKKs60uyy0VKKvWhWt
tOyI8T8UVMFayLeWhff3VBWPLiuaVF9RI7CFHvBDeteH+zljqRA6TKM4uvyyg34mOEAkwAw7nj/O
feAR1odj9A7vm7sH9ECg1fLHPD2yPQZhqsufvsuFgcIFIzVuczEJ4aIs4OLxVtfgRV8sCszvbLwU
yLIpTQMI2I6jurwRTUglLQj1m17bryglgL1/2Xf6wA/kBOXtJ7ePtetpBbyYqAkxjLBtikiBtJlw
E/9DLS81fE0AAEYqGlqRgK8esJXF4WwjI9rwM1TvVZf/Ip2H9GOsTWjCu4wy0L8+0r0RcE+FmaZ7
5fUhYrqswj1YEByUmIyJzeaE6I/+ZUuzi0/LZk5MyE0zVvxIVpdNCONkXnHEicYCpoohHunehw5H
F2Vb5wBnxzvTcz4R7Rf49r75ZQpj/4w3f34hxyXb/0Mh5AbXKylnDqlssZMoBlUKwLapLrlHjaxm
FKvcTqtffmbTs+RMxh7/DA1GEYTFUfE37mhxetVK6yw/IVkZh18p+ZlN9/AsnfZPtV+8HnEwDBtL
Ijtondm8iZ2HVMQZXXcx4eETWVljtBJIScTOUu6vHmSnePVEHCGJA+ZH6LgVmC/DdwS2CAshZKYt
dZ0LVH7qBN9TB+CAfXOzBTSXcy8orr26lWsuTzYLP+p35tLQLfdoVY+ceb5Q0iQ7+R9/YbKkDtrz
akf5zXzn9ROHr2cohHHakpCyLu1XtJLNYcxjlGuZ2bfJtzxFrfnieogs2vCa1nyj28rilRbCgfZp
WHL3IlLmYP8gOxUUQa8nsM3UdYrgBaGRboculOgYpLz5KE9hLurCqcW+t9VG7pagnsBZTXi1w6s2
Q03/o2L07TP0pMocDQ5TFgwLaHZMXSuhXTXQfLcrJgLBa7zMjG1QIHvZ0YAaiBJvB5D40JPkBXah
5e20XCbXx2uZ6e9KVhV8RbuTjn/Ha/f6F7aQzYzqX1AgnHURdg5J/Z5/x4eiFzKT/sOK4wS14hLW
2zKUD4/cnVUtGZHCdahkYX5/ehTc+LZFVHZb0t85RCcV8sLrukU7PGtaRaOCAYMVSs+Bps+t4U85
Jfg4v128uUyfQbNpW6Io3QJAYCPywjdMAHIGeeyCtOkSGF0e8gVHzz8ivFxUShVsnJK3vMBYEnVR
+8gD6A4P0FLzOL73rPgstCEZeuOuH9IYYWOqplXAYlHaoZxQUsK2RRL/ydD+XzaUbqYQFKNp56cL
2+RTZHxslRntQLDo2gi+uteQdXXaQ5EnXXCIdmsj1uaaFtg883DXfZW9vtrg7kTPl2LfFNL7DorS
/xdhGE3Q/iTJTp3yHa3DB0pZxnibmHI39jpBrOgiuuygxAXv/WP57Bt1w/DrWnLxWFB3H4Lp9yUM
UHrejrffyQUpT1tC0Fu3To4H0d3Tm+9ie1LAmuIn6R0ovZbaITwFzzKcZD9wD5s0+2swdYTGYxrb
19Q6g6+FUl7+NRVUXgcuaJfQRnJEFJwIwn+CFNJqyvCAl2FAPgw/YOfzTVGVDvgE5b1LyWDLB1SD
PoJPBugWm2eje3hXV6M0M8fh6Dc56sLphO1IsAEBtqxSwqwSwsswiSyZ3dk68cyykYdoGJR4v5ma
69M/4PiLIJ9vz+W6yM3K1qypWtjRyMTvHR/dYZUN3wm9V7DDpBjAB2VNuTYFUTpCqgBN4knmN6K2
UMhBoQpNFhYupd3TAR6KSUZW7kl1O9E+npiCx54WGxLmUqL8kcQ7j1Zx5pYuqS7jPSUcNc5A6Hty
anztXAWWyVXvq6s+B+4Pc1J/XNTeYZ++TiQgm64KhcFyC9aq9Jl5JSfjXNQrayyDubRhOKiKTPLJ
KAOwUXaiy4i9BoZbi0RG53n1yGIExRTA/IZtlQSA0YXB9jSJNWFMrPp7Vf3vLqG76SLjpQW8KYcN
TKDKzVagEhNscu62pCLRhYZMcEjuvAMFprqYLono/JJKw6xzXkW5sZOS987JCz1um9Kt+v2oR/5x
6DKKQmerAlEFleWuhpDZR3/xBJsrqwRXU4X9P6TRWhSTXi2pCIHZPzJNzqJweF7vGVXXisBuJQ/9
oxvKuKMajEJEKL8dBrKeAbT5OoZIRsiTBlCKFQkcMt9vMVzN1lNg0+D3nNiF9/Cyl4swjtuwbVjV
fOK6Fk4oaWHZ/py27g4mBBvxZ4roo9m6uMROfrci0YZ+aUsWT5r/8r2ASBN7zN/fRzjHE0ZTVKsY
ib2VoO+sw7P81AGV9KqSwo/mhrg+OoLxEJCEKDW17JVTaZZ44WIak6zKLYHPW8Zy0Z+b7/40gKkU
XD7ZHRhw/pKIyatDbs0KCfpLLaoVBj4g0xg8c8Edi6aO3mikqGxtnNCG5xTrjHXXODGe1A4WPVWE
eHiaw5ZmnrBHF3q8wLVFepVGzrrjxKIFT/xEnXgBwS5x0FqMTS3gN732aAr5Z+i51VmUBfRSR3kk
9SuRjlOD4U42VTxZFvz42lWZibVRoGdRUPxMBZtx6hUqmb1kWhR4C/Bf4OOfQ3dTjeLckYXtBRSZ
h4ZhJqW8b2c9av64ZGGpjWEiwqUlZPQbtaSjwbRhjHyp3BxySfK9z7RMaOlmZL9qW2Er/aAm6sxa
wgeHadjeIsgncN+L9uPPpA9Pri/4ABe5/jpxjQtRc9y/v0rKbWpRF/tbBJ+d//mLGAMz84kym7e+
wqu9seoPi1N1ZnZrSZCQ0Pl43Fgvm9t2pn4vqvlLCgZRE23RWSov48AOsNWVnUnYZ1Dc3eBliC/4
TNy/tBaGl/oQiPPmgTL+IUQnRLazWTdNHdX4cIFOgrwv0g/nFizQ9hBu3ee4xnCRAKJx0Z4fGyRk
ZOCR6o0G/qigdNFw5C5l6V8ioPL52AQt8/BpRA6tGJnJT5Mr2mZSDOjhUPODLE5b6RsparQsUdkv
3M/jZgLaOroSgKOTqlwTR/nyfagDtHaL7yq4pCXzLUcpBeG9EsyXQ1PTfdZwoyp/HI19IVb1i4FD
mB+Y9kRGCpw+sWc5HYjKKfDdYFB0nWzqN0WFrbE3mAD4szyX4bEAchiQFHz+XIvvwTcr5veOxCj2
OrFCnWyJ6VC6tNqSMLMkk2VhZmZnDhFRJJId5/zaRcG5naM592sHsSYHC2lPEBjYSv5Sk53io4h6
hQfd8F5nkpm9kHyVj3wGX3HV0JNR3LY4VP33TDT0GkspcKmP0vFtfB7OLNnBv9usXmHdZZIessVM
+Ve30vlYvV3/81Q4zE1sp7sqs5bH833FHaxcMoP/xSEA5/9Ky2ijyJ+4HgaiheSNsO9MXwbdwf3/
DTUszXE8d/7EmyjepeMaC5a2Gz8oZCWmfDbyvs3vlWMGuv6x8UYEIgftFhKckyFhE1Fulu3f8lY7
CkdlLeppmfw3N38j3Jd6R3qJadCo8QbmP6GMxWmifr10+aK60s1oj12y1vs+5k4udXGJdvAGAKZQ
yXkpyxCi7S/chEx2RxV8NMipHCmbvFuQs+jNWhU0j1yfTThxQ+TfNfsPD4N68ZQnd8CAFKLXaNsn
HeK2tPMgz1cfHR/wEoteXUMY2UL2SC5Z9sMSXpqx6J9O8g0ikG+CY22jLUncGcwL6LmjK+9oy1i7
hysBuqxJi8SfiTDc52LXZetrcDFJ3ZSk60B0d7oRaW/JppAVKvFNrn7VAmh01orKL06ly9/zF4TL
VcWNvJPCEghr+WKYI38bGQtcg+cFYfZp4tBzspWnXhg5uTqDtxYCZZIuiytgqcAf8ppK/ti1Suoz
Omk2LEkGgPB4UDDlzawCXXTwwGb3DZ7aML9nPpJeu/crRAaClYh1bJjE5KK3MI1duIWy2mtVF9Qy
RQHj96GC+0n3pAjmWChIRKauHrUwNLf68o2xezTXryCanAjhw2DKWbzdK5woVLoXhlTW7pPCNuch
w0okl5kHmDwM29xEmp3wgpdyXnfkeMxB514lXa3igjzwedOT8QxGqH5wOlyVDNNjLdww9EUr7Uoj
NFdnkBECWLFc/j18F2vvt/ES2zwNYvRbnTFmpdOIWiknRnWTC5q1hTDrBSra8PxOoXBYCP5pXoKz
BEPE+KNrRujaUpBe3Eak4miaFD0k6dBBx2+ITVS1FC/1KNBjiy74ZPgzEHQcgV6AAGyCW2Lxo29q
aWcQEhiG3SEEYGvoIhhbkqZvQviE+yNbVuH8SdioUaq/O2ZWcV1iQ+JZrlaZ595zFj0FfR3iDRSi
ob+RR9IAoqEgGNSEqxTlk6JPRoYpQPL/lZZohdV839peaJq5f4rQGKX16B5pUx8AcLa4TbynN3vs
i0Ra+fwHUHtbSnZRh/gQ5cWhTFrQULhCOyDItqGpMXczQsf4j49hEj0YAL3d+jYKHqxThIt/soPB
iBM95tht+VLaIiRNAeCOKSDVtxHJ57l00YkjJszJmsDvs9oz1uHLLkIMPT/rpi9RSXB35u/yybaU
hYOeHADdIZt2h5jsh6Z/X6lqIc/o0PtKVXYQghKsiNDpqBU6KxMMwfjfn5OIOlqcsGRzINq6wpEA
rv9U4/v98gfjW+/sMn8/4//GbBpzdQWwAIkKwCqUlijqANls3TmczT5rABr6k8YjhPRFGtP6owXw
noVup8kZmKFdWPsgRMyZ8DUUex6RsyXKVwW9eWQfGRcxWvpB6cDvq4yBBCTE4iuXkytjIv0BD1SF
UciSH9tStMxPhda4Vx8bcq72lbikeHbDW31TrkT7/GZ0G1QaD3YKQaMc1Wrb9OWbtHFFOuRDOASQ
W9tj8LV4b+f0Cl8cDBanijfgJilshRlL+LLBMXgvj/9gx8mXxaDk3SDcWVAAYkLFpHxicKa2w5Tn
qY5dx4zqNb2z99mCHTtGpqUgDkGeiJuZ3Z6/iKJ/LrK3hWAI0WTHr8EYKp44VxZYu7z7WLEb9J6Q
KUwjKncvC70vQJpRVt/n2nVwmopeft0/sJoHaZWppThd/7MgichvtgfswT9gSASxo+BMKuxowZEa
L7NrESgfUvMpOlQRQvPNTZwxsa2M4oTWZdhE66Gd8rRKZE77mSFxPtJOHd6ssCpPfGdLh0zfIbHt
afmgUVBNrSOLgFJj4ynUloosLdr6c9RyEaFF2LbS/hXYe34lkVmjz4+sLj+u++EFr8aOduyqkID4
9tydCdwDARIyAf17iNTfMywRVUdA4k0e/J3BlN/IB32x/x0yZYSziPP0uZtZVkw29Nd10bO4n2nL
gZMi0hHSfJmF+YKX4evPAHWl9j6rxFXAG5ZtJHLhwJO9IAIr6B17HCsnLrDqcp5S1KTm6EC4sHNQ
Iv+d1VBITAWRCGpEUZNHfJd1NZFsIKkRtbNOZTs3viJcv+05Q6b3k8VzNjBvgbZ7i3+GlEEOJpNt
QUr1vIZAwkYF8Jq6/50lVwnfaQJCDw1HWVE9Bp2MG/94cg2PJhKu+DH99+FOI1Jk9Bb1dwNu+cT+
mFpGWSymHrVF5m/ZhN2C/OfGmGklOXTOZDtRt5uoOf8At8VcVwvizqlpy052pR1ieSybjTsbcWxB
8PE/EPzamLMmRaK3yniPIkaKCNqKu+D5OiwWS2Nk1DJd6FNKlC6gCHR5AF0QA9iET2V6ZYqsJTdq
ZwAGioW7S6Uz7GYSH11slP8UMD/awMLqHajFDE5PuztObRybK65dFfINBbdYwgWAOSvLAJ3Jb291
wqNoVr9V7WfoHlhfUSYYH6friGc5JVGQ/0OTeepY6/HAas7TRfFggYP+5OUddVcNNgcyUyZT0QMe
oEJa5TZa3QyCtbFfADu4Hh+WHgjvCyA+qtKq0BXjznE+O3MnSnQOvw1Yu4ikV0FS/bIRvfY10VCP
p034KXJWF6jOU4XfeMs0kH2Io+Mut/tSB2uBETQ2HNaFaHpK48e5WIFiFLxwMzwA9MStANB0A2p9
CdK5BhLSSemqokF8OILxaWdw3MrwPSr7bmXtFPb+ufLVt9VFzsKM8pPZEY1z6Xq7LmAGjzB+0ZbO
hhVQkplarphUQ87nA2UX9rAfI7V9joLww64oq5EyyJJFUbryYVVrFNAM7ak+VF3TlN7cvjIQU5Jb
dBGomRUy1kLUXeoHfmaEExOo+cbl7foT/D1HIZUz0xWVxy5XzxSollxO5r65StTZXrALA+o8mDRY
zTfhRMdzOmgl78Ww+WDrQPK/9YvcqWMZ+e0Ex+i+vReTK1z5GfHQXIwAWljQ5aGXpoE+o8BOJuxS
8ptaDYrIQIJ0jwzDyACEXkI8JeDseWcORoTFXDK/wbmCdHxtp0xxoXJfTTv0Ht0oJc06F8AWtJLp
hOlZCOHhk6W0yKGU7jw3OY+EwLR5uAKfLr6LGI9nozWzzRpTsw7QZwdx/wrvNICNlduDO05C3kEp
xI7XErsXU7/o1r/29ffZZsVf5KptmTzfiQTpM2dE1rUSlmMOFvGCV071YHZyj7bOBDEog7kjXqZp
T0Jghuu4fhU8c3yxEY8TdzOVLqrfgZ+QgMtn7NQBfcM7uAIypg2DYV39b6MSo5ZCTjkFQEmIWea2
FS68N3WnLT5yK8GndKbdyCQtskoTEqr7RFaHg8uKAjS/CaWbYFCnX830SLhaaAFsf9BKC14vxrHH
nC3RqB1gv7n17J0ST6drU8mSHr3pkedwRrwKhE3pIBOfA96qTF8YmIl4RFnGQH1CjV52+5NWSSmq
qpRo2WNCF5PLgzfLEyNOaEGDWKhDGka0UIs1ZwaGIzPS7E/gkHezi91/S3wXFLnrN3vHLB4CPKUm
jyfUWO1o/MdE6t/Q81vdHAThrgc6rferZ+XXRGarOx67ueDpYow8vIg8ioiZkPZQtbZ2Rphwz7mt
5JxTCSNkEcyMU7y+ER4/QDsiUkm6vA/d/hlVJDK0pUIg9+/keBr15xeB/JgB71ZhOHVNbVUXGlu9
oL41Hg2BZ2JWKYGk0WyXBTLsD+VDOumFkomcLkipo8ASkde3T6VZvrYbvSudGkexNNXVgnEaEGTV
B/HFvkG8mrUdQ4ezSL0KY2PjHLsnXy37j8W2t4tTqMt1dwIsDhMmhwcZFSYz4VwGXDRtMUgN0uRF
/L8gUTGz0y5hRGa0DNPW+rxEkBRit+omQBWHS3H3T+620eqQ8LVZaadZDEPUButcA+iGhxmveHVI
zNZAhKL6GGBNXmRrVO6blDcEVJ/S2Dd1NOFtQORIVBQQYONUVZqkQzbmuRF7tJjwctj4fR6z1gxB
BP6rGBGoF6OrDHKs1I8dZC3mtFVoZR3X8gB48aRbPc7Nyl29U6hf3UAvump4967RyfbxCthA6oak
4vNqfCOxIo2P+7YaDew9kSI5i+TDFPKkXbaXAWgVRW/vnm4CdyUzVL5TBo4IFefJgrPtmi76RYL4
Snyzv5/tTtu6rwN3fGMtIUmB7Wz7ck3vgFYmNclNiNVNBGsc1HZqsy6SQ/M258dT2ifxdZIAQf8W
/D6zlYnLUBukDyhyERNNlJlwhMu3ppupPUK9tTRKnN7hc0h4irjFC3n8rBCaaCNNdBynyUtBBSQu
1soCjGFDnK5nA/SIjCd1IrvlaEJAnddVUFdsL4EyqQAjohghEoYFQNTkGCsSm0+dWJMGUhawYWGA
sCx+7BXMny1Xdb1+oJdH6OWL5aG+jAn4cXtnl41vX1PkKZFRgVoCWDKFP9j+TmwAm25QSoIA4xG7
8M08GzP1eR428HyVa6J6Zg5i0vrqSxEtP5IvxQ0WuxVlWQXfDUW5b5t3c8n1ZQB5Z7A+xqcGxJ6s
s8aAWs98xivOXRsLkPBhqukqURyxUgsalYvxbCc6qJLWPr0lbIZ5XRrSeCDYOr53qR9Y1MV9I+3E
i23z3O51vk4vTs43no+0WWUgj1CADhvJpwCMb+gHT28i9Kx9PivR3UkNBIff2gIodUbOqjDTfbf5
bpViNet4iW55IiNMDzKMpM/thvLhfSZ7e2vEYt7eUqZ4ejp0Nfc7zc1oMSEVdBnYH16maDsu4VHv
GCJLdjKfg+J9nyojoNMeaVhFP88DjfyODfn/o1Pc/diHLlH7xk6UZGRP3GzVB+8WoPezHMIjKh6k
rq7rtYx1dPaQJXvDQOrWaViRoFECEV6IJACQ1o6ILgovLQ1m8ZRs8D11CTZQQZBrYoBhlojaEIat
KvByl2TcgVHgUHrsHTsidDbZGw00s3/pAfP0eHbka5fmOfUIYOhfCKHhrVkPY72Dvfwwu3llBbUU
yJplZNRQ7z1RTK1bHwLGVY0rcZDB30GJokDNnCVPpfFhlJEan46w5v+yDsrvlWs2qD8CHsvH8sOz
mT1MvBkNn3IT/jShDMVWX8xRVlxQM/aIImLGcqHJ/oituqUrygAx0MhpVR3cLcArnFhHMb9YcLmc
yZViK9oh26Ksl9za5nNW7tnj9ndkrTFWwQOINvNtAIs2xLVVHKD7dvQ7eFvfkeOlaLTk5Ywpt2Ss
ULZcdYzIZc+mRNQuIq1t7Pw3QPHNAZUHJ9mzWq6NbRNuq9FD306szU1D5jBmdvqUqVjPnFDXgW01
UiBwLGkfqMpQPbPvRFYobHJTM0MNAg+IdCGX63qGWnlE16fDYKHfNX6yPIhdZuDYdAwxzongFw2Q
NyVle4hsP/hfhT14thCAnSiLmv+dBWOteBgxNg/VKODMLy0dV7OoBGygDLYv+eP5qqewu7IaFL+H
+clUUUij1YIlpTtwbuc99rwM1zkG+QAFyLrEMorb7sEjzZyZUs50gCQulANxb46JYBg6pxWdj7ce
1RPnHaUY7JECvmnZtqRjCNk4xudHzEj7PnTOebr2YWznS9enlF1a+yYNbLIu9253PeB3YdMCyifa
2ODGd6A8ZJW1qDtJJhCUr39Rq4AQuNxpemjERSdfKNwMnKij0UBMM+38V2ISBrJmN37G6Tj+QM8S
ctxjnpARfC7B2K/WxpMC+iYW2uanlpzyhymVkKZ7dBlZG7O9IcQ32T41Qu2OJ/oH6rnXuwLIALjd
zbv2WfXA5+LUGhha4H+DaTjPYt4BPGdC/yEjSlWwmHJyDsNwPqrdvjiYJOtWCi6IobapbHQx5+1R
B+cCitDPci1FuoJHXQhi6oE84SNLaOPDS3A1QEnJG2HplN+16IG3Owzj/fPpUIUvYguqcZ6JmflQ
Cf4RSk0hBGY7avYAJxsBtwWoSON58hpQ6YRsxErTn7cLql+pM8O+PUn/Voh2Sbrw+GK665ceZAcl
hVrSAnJxYvixvS038vdmvMTKF//hlHg45PnBgJ6pIWZbL5iPfg5VU8tPixMYHOwYb3dRUk404C7k
dFf67wIsDeybMzk4siUjIQZt/iIC88LdZ8M0+EN/EcG40gzzfWOF0n1xD+e8DFPsOoLsuUMLR0hI
rjPXJyXXcym09u/e/YAyKFDL4V8ntze3Cd/d0HujEoKNjpG2u9EjIanDoMz6hDzjoGDJyATYlOld
uAjAD1+fZ1U1C/KzI/sZitgKRVmvzBmXDMkOx+99Sdw3sQN5M2hIF5oY7ftIbwr5LJN12iZCL5KO
wAfJLHwMHDtrNgMn9r9usBAyNEPSD3RVfuKju35YaKD5zSUfw+sFINgzl7GI4FbtpuppSkWFxlCz
LT9Lky9R26tMdMu/8X2ZGL9sXe3bDcZP/VUxnZyTW0cFQm/ekY7FFEYYS/PiW6y5YcsiyEs5PrZ4
X+Do+SfLehF+1eCGLIimSca7EXlV8W64TQTTmtRSDO3dwlsl4LEhFeAfbtdiGr6Y0nKlk0++BiU0
W9t5p/Ud5efM4JRC3tPAMFCdwUhTAuHGrvz8UXiVewc22Wwdyuxh1Cct95qH/OcogvHpfCsDLIuJ
hpzvttHitCgkOFSr3SSHF/ERzYJQPsfmTsy3Kl5e29TzWx4bhtzROgrNmV1mXLvzHbsANfg9rpwU
ep7TJwFJ0gOEb8e1xfIKP3VEmYtYhUcbnpVgG7UoNw2rZ0w0uq47GB5NAkpjHEGL2vIcGHcg1lLz
yFtuCOvasibdf7/7kuZ31ePxlbZiOG1xl4HUN7xIFyWJuclviTMRRzhw6qQkOhI38Ceer4FhlrMu
GNmlnLqwhtef436V0Cx5QUeD2PZPmrWKP+i1+LrrK+ysIQFeqW68/yuHO/wj1VKbp8PAR8TQOBhH
C26f0bWchNBZD5sTz89JhPKufXaOqhPNnFDwddb53BTh4Il4mYBzsc/j1RJ7DKqvMbVnk9c9SKwD
nrl/FMdnf8DjSN75AyOkgA8C+Em/+8E1bybGYNPrW12Pr//xJnulICnYHOiji92KlBdWOFBKbrI3
jrJXsAB9A40xz04puhcHk7VX1dWRbHjthBtE7GbaoOcT05bzfsTvgOJJeQMSZSq4SS56MIc1Lubu
cZV1ATQMq7Vubddpen26v2XSMoR762UC5R9S70vZfsC6QPl6Pb43tJdld4ZZATFxJfbtFA8nV7yA
KTgIskgJY/7uvC8wiPEEtKi6zBOcAip8oPTQyuHcgWk0Ry62QpydqsU5uKV/cgywjy04Y7B3/doP
n4RRqfipZcopt3K4vA7fk5KLLs1L9HSOPQX26SIW10maVUyUF9K7NApi5NH9slqk3xfn/HvKff5u
aWZACTr06Drtn3ecvO16ibLs6FKbFp1aUg+mBNCT/4KrnrGiurTggg40UpmxFyXdqscIqBecZh9u
tRsXhLC0JJlrB4LCdIzgA0bThhfC7ld196I98UHgGBvOLrgV7KegEme5gm8+Gn+qOt7PPDIRSyEC
xknOhU8eygk8myH0b67/zPNVkY/l0GsfuwGjoS8JbwwuzT9YmZJqBA8Zh0yQOM4JLduA1aliy0Zl
1QHUcxKO4L8WTluWI1fVx58+Ud3NTfvARTGfKIKFxCUpyxfxuHmBWtko9u/1cCd+ZUUe9BDVEIr2
W6/XvR5Ef3P7h+1dBFBVIV34hka3DNcjcuKOmtI4EjFn8CSIS+C05yfvcXZSHticRGuQ5ijNvUBS
MgthqF5dLnbXhu+JGfi+f3VlT+sNU/JVvOsiOTkG+JviyBqiAOZoM+DtzsqKwVQ/QrE9lfyaFJjQ
3W6RrSTftrZR+hImJ6rR1bAKPgfM/jFWLJnGorMKWptAAHSYf7xg0m/NXRF9GRjyL7xZXqtug/4M
BbaDGoSLoaKebAlHQL2pOywI3DYdxjIJixhei/vxZg0IPKZpK1Qe9rTDUukw66lRIiM6GTnHpA8r
2FkjCW81kJAWsTIZpUIPxcVxX3hSuAazncsJaV5jwUPCkA1oz2UKNW7Ux/6HNmAcN6uxqYO1Bqfu
H3SvJM7jq+xZFBa1jSvEpA2aCVcB7ztv+PIQ07F2LGrZT6xKgLt9rQw5rjqMAENTHbV7/tVt5D0e
UOSU1wRKrJfiUvf3mX8loDNoEIvH0dpuoI87PXpSdf+386s0iYgvi1T7mShcxVOqFS8Qy/CHggtv
ZkojS3xWNixVzrQFk0Hm1tyHr51C7lDYdZNjl30iQ1zie+6NPlWCwgWehyMM1VLPbYhV/N8dlI65
3hS/onHKqTAsI4R7V2a2nvNZ8e8nwTraxKVgeBp2tPgYLo9IH3Av8ryDEU9VVgOqkUE9K1A2KL6i
KHiG/K/EXCWcjMKexwQWmWO8lz5lYfBA+IN8KeBz2zbSgFNzxr+y8n7PPOLmv9wg5sx+DUJ/MlTF
+ZwZ5L8h4bA25sVeKFnMM/PaduuXqCD0wi3lYrbelQe/khceXepTPZOe1nJafBckxVRfXns/xufr
Z9XVD8dyaQvvUlHnHDXTYNGCz/QgmIswpvsbRnCR+fiOl/MfyUtpc+aJ4jcBgP1TMqkc+lBr8uwu
hdhC9MG+Lznq4ipcYs/IXBZ4f0siYAzSqkCl13sK6SciKAUJaEBQT2tdVMgae0idFfY8lLDwZXXm
edNv9MmOrqv/jNBplk1iaBLmb7VkAIIqQLOfsIidP5u/toZvTb8V8gzdxCK5WEOVHLCJGJzcyMju
oBcnzXIGWXEl1/N11HIzNd53RriNlycAzrqq04mOtwVy7DVLszzRwC77L33KfoJWqYAIL3R2UBjY
i0MtUSb1DvKQa9QJr4BiTnMBGncMyXH5vE96kgVq2m6esTv3oOFSTSbtjxm68HLV40rpDiruI9eZ
+qn9qAvOznliFGCXIUy6s9HebsF53VFJupFC5/zn1Ko26FdQsHR/Qg23JnUZI5+2lRh48AbOWcxa
Xw08QV2XgFBH7oaNuoWtVXTWCeC5hPlbV26dRoELkYKShP4khjJULQMf9GEN8Cp/2HW7BMiQutV7
wcAXTcoKQygYfr6J1i4GICvLncmlhof3jT7cvkDIbLDZCs0I4qxzopQJS7EhZi4ky89om+8EZBpU
pFAFMjwrPE1zzxh4DYwbGrYCHFDqHm5dsai+U7NpjltjHD81//IJKODplfGwqoWhWOwVRF50BYF4
GtkvAIhRPUXktKR6H4AJsIdzF+1aEqeKfhJ68XYxdvM8Abi0RIu5WCDpMgj0/HoEPjXFI3a3Wps9
IMlOW+m3pnN4ngNsMEhzzk5/FRC0wm3qnGGtYVcuKafbsbhYFWKDXTp/BqjohOa95V8sKDMd5gcT
1/KzviUZP513PjgKMa8hcMBXc6FcH8MW0mqjjMFvmTbXtEr1e3F0KWzlqRUgJu7/IIYr/HKi02mh
PSU+CU07oyFO+JWTKPE4vZnRTjP2pp1tY1OMTS+v+EZxJ+BZmf2cqY2y5M5g/QoyAet92vlHC7np
yosQ83srMo2QOQsS4rJf1XeNYA+ixnCoBfPS8hXETKRuh2wq/hswdtGGheXBob59saYh0MZVlsAW
0UTeJEUXh66qadqRnCwdXdxOj3PT8nOOaTmCnHOt1BQ9Cy83TRl/8ZainoaBjK10elglCl8qPS3V
1adWsIO1dZYVbwiF2lH7OFC728Sg9A36OubUeQ7/0CgVoyzDOhPcTnJqoxJq4fhELcVlpUi1I6ny
t+0rloHN36pXhcFb66MDYBN71/U+mI8gKI32N2p6fPHe2sTRsU9h2X4UQLt41NePPGZIDKhG5HPe
/oPTLWZ9awW8UWgiR04Xp3ih++Tq6hURfhlJArKS+pVzz3s9uWY4aXtOI51i2kHumMLLweXnafq6
XFO8v5eCihMFANNJPnfHfIflmjrcrVKxAml9osn/MiQyPcifeDe78YykWTfqjgqczCwnYOYlG+s3
oDwRVndpIMKAPA7SZPdGNVVhxwTI8bat6ATNUu3wAxo28TlwNphd1Ql02C3vYLAm3GBD6oJMM3H8
JqP4T8Xr+MuLlG00HS6xpvx4tcj23TcRn40b5GFt+FreYQW1aaF1ss/Ik1DWRWgeFKaXeFjGwyLm
5wLfKQ+OLj8KQdQOggF8wFpuaNJREp5sjr3DTXumXmh+zLutB/OIYNqC12aE8HP+VXvy7kNh56u9
AQhjDYIOCCFIfjfaXyRNpQmDvBfYFZLDv+KG/cuqCaASCQSuWrA4m+UvfacR5xVrXHqPYBjpEL5j
e7DCqtysqgNhzdBG1mpMep7I5Sznn+BEBWw0UtO6g+uGnOveXxRdY3S6DIpCzbiY6umh9W9FTVAw
t00FcjrcOi0oVVNWSnjVV41SKEyTOetY8jC/oXwXusROtJYIU1f3qDFWfjYq48rDQwiJjeNH5EL5
aSYWDHeDmRepS9hbkm3JoCzgFqNjSNsRRAYK8Bn5gPyQe6Rok5G9DHnI/b+xon2gGsw128/BExYb
uDUntjV969Uc9U0oHpgDrCFPKPIRG/FKMPhppZ0CWQ8DiBL3H7CzlIFGqyWVJnJonnMTmq0zo/Wk
PwNSoU/jcQVFPZOb2UdHBYWmthFDNBJqlOsDj6yTfjzbmPrEUisoWHhcNjVzuqaB65S4Yq5a24u9
XF4tW26IUmBpACAkxW/o9AtoNiUTUmGBMAkzYVSVwmz9HJcgpwOocesSgZL2dOjSlDVvMH3iBQ47
V2FO83XEAPrBpUmlv6qM0fhY+3ByjPFLdpUpIUnY74ZQUf1h1jb//oiWpVvPUPDct7DU64SVlC7n
6bQSh3KGv0+fkyurtsPQH521lRwsx/srElSkIHyMvynFQmPRB9F2UKdp/rEaUeFOg8xh1zMZY/tt
T+lbF8btsQSbu6aD9LIShs7Btwbc/Cty0xXIZ7hHEZgcU4TCd4PFsYUpoyu7avXUCkoSfsFL/KaN
v0B4+/HoW6XQwDJVC8i7a63eKVg71+3zBvVmz5deptJp0DOXQW4nxSr+/tpXaGyue+965dZWA5ql
XhkY8dC9Gd5HnZ6/g4Z3mjnP69ER6QB7XxJf1guUNnyxs4q1fwzTf6oNz5/oL2xPBg/W73KKM6YM
QmD25slvVAFjox0gm/xTe/M/RekexL81Rx8fQM+Uf5OG1eSde+JLl3fkSIlLFLJ82uf+jheNm9ls
Ewyw3a51twDY+EZoG1uxOjFr8VQZkw5Slq3wsPxZloU4cYUR9bTv0NNK+s4lqXbfUzvUz9OlmezP
UoDK64Yi8jpMUSah7pxGxqHKE7VfQ2zRbeG3Ffdwalt99gAEDeKmRqKzqLCjOAyLEkXHF1yXiR5N
L4P00/RUyX7RnRDC2XekhpPSqOJ/moCKOesThePYzoSeB5gdVfv1EVGkhoh7px+emByE7wTFaZrf
7SyfeJfZLpqCC8hYwA+ChG464bkpdyVUySeO4tQObGRCNtdGc3hP5eH+2vDNmVU+AiBkxpRDSBDv
T4fS5BnrA82z04tM98246UoG6VD40JznqScgTykI3XM11ydI7tKxDl9YaofTKTsj9QR1Z9Loe+Mt
6bq1vN8K8LH2tlkrwBjSXA5QGzGP3QUk21twDUnWMDN1Tpx9Fh6H3kSwzyC4TVB+LSMrU7i0pg6i
KtcP7DmcFw5Y0wFLv0FSw3BxmXPrb7lO3TBKGf2C10K1KcR3EeVzQkP/9pQiD0qSiPaDZ6lOEHcS
WGKg2WbT7HZn7gtlicJlyelL2FoyNJi9hVTNgTtJh1skp1hi5DUMa4RB37bV62ZkPSWr5lkf1cZv
QCQGpp604DgXU+xEv8ra35mMXbldHNMjCTAyFBK/k/ZPJ8JwtQV0m5czmDfTTE6xiyLy40MQSpYe
6/CD1RJl3C/Zl5GVnVW6MffuEV2cH7mv9dPHiIxjaEwhhtNfAwJgI879byCx8I1yTOEzLwcrbjdp
D0At0YG11iIy9b/s6WRe/x/JNa+sVIrXQtoq1fkM4oNrrrObXyy0W7iBFtftNVy8Vk+nAFm8AiDP
LNahOBsblilV88+ODwkQyonwTgb7Mqj+uDM2y8K1QCB5+S9o/uQbez9+BtKeiyJr/7imNACo9Kch
/W4ZEnlmjVg6lOpOm16J8ZWiTudrNSwC8z9W8L2BhKtQfoS8Hr0oO2aU2tjS7nrloGQmFCeGd/M9
D+rDQ1Eru3NfI/hS6pz9KOrFp1NlcSZlLeEJw5USrkHj28qAd412GaAysSMcVRQWmH4IpgwsYacv
JBvPyehgNCTvqnIAbx0L7x4c3ApUPvk1giUIl45YjwEbzeF4L4wZPCzRd/hhTsSDdlmn82XFgwA/
u3wnONjrsTPlIoxXmOj7fs+sUZG9YC03K2zRXLzlhK3cisTSFBJ+89o0fvfF7a6O6OUJX/Vb44sZ
FEmQ8y5Hc9M+zDH08lf/5kSFkzhutL/r6VrwKerXNWXZn7y74KsINFM2YctKEaXGZqHkPwdYOLCY
TdtoAt0kdhAsE686t0+1PpJxoHnqoRwmVKLLB0BjRtyhP0eJ7KJyUJBQoUC8CmtdnqfKuj8ibcHZ
p1UxxyFex1afrc5E4oHnJL0PYhYdzRFtR2j7btNhHtY03wvZmNW5cR/BXBqJ6Y1req7jodCDBK+G
CigfCNok4d+1JAFXCYta/1wUImW/jEaE7pj2RGt/uGS7Ed9RE08UCXIxA2JPATirbhM6lopENpAB
/tZkHRAS9ttkbADaFxf3Lwp56YxhIru/XgoMB//p3uo4luLoIxPu5sbqgIBinxf6+beZvLbd0AaW
MlhSvnWD+SzyA47GtYLscaTTPZItaw11cwFKtBtdjfORe4pyb/FWRplynE3IV8xNzgkDig9RqPEO
BN+pyzgNMKTwLkcScJZ75XVy1CvKVnFDfebdx79ya1fEgEfN3oGvfPY0ULDYddu9hvTozUq7mASQ
0oIW8coydoqM7ChU+9ATmxNPcEmVObxbi7rXcJA1lIjp59k3Y4IAT6o+iNgW/y0MesD+pIOcB9v+
+9deOP2HR5jJ4ZnkN78YGp6v2XgAQr1YWjDZMrJcTTZ4XsQzh2fPETZMpxZ9QcS6ZjvnfBYQ6PR0
Y5FOgqYKjmLPclFgFYE/RVzBVVshH0pTFz2jraa9JtHsEbGFVHXXULZZJ7bPIpUvWi7W0d254Bmk
XWEf7bTl4+okGR2UZRrGnSjm34z7Qog76641ApU6v80jnvxJaHAdAvC6EjAHqRJWcNPdlIt+BQmp
8rjQzWRuBZRtG1w2kr8F4w2fKiEq1QxXGH7xdnBVK7XLiOaZs6Dt3oxfcJYu8CerwF0hISghaxjc
rSLbU6B5gHR/C6An5lpqLasAWYtSkwRUg+myo6Kccp0iDwLu/u4qrk5tC19Jn2SuNThaD0yKNO3n
QBMCLm5HtFaMYHrSxWiCxkPFVJBJvNp5VDtI2X3UkHpUo3+i+Yfm+EWdcSGt6Q8KjVgaeqsbbomu
9yw8uU5wyfv3IvtMAaRnQMYA8o0f1bjL0uOodK9rSbNbAN7he0yUr9yY5dQYNALpiGEmFf2aKhgf
3ZKxxqE9YH+acDll8l+3ZGscg2sQf6NOZXfck1crETbuRtZ1JxZyWVDDgB0b4+auQQRSvN5ZsykR
HvcLLTV+HwJiIlSOdkx/DSO+itm7fsxi/1dovFPM82aS6/E8n0i8sJ11jpQVynK4FBgzoq3QQArA
goKJ5pj8Gn3ar3sQ+eQL/iV77hjzBdHc/RlI8g0CLUk6F7+/CgB5HxJBu2zSlDMjxYlk4IrxN9+h
6OdKJgQ2yvrqpgJBF8cHnoDYaX51aXbzxV4dG/H4AWvRN1N2xSFz1USBIinqdP5yXOuCWseXnQ4k
vTrNSJv+aVFUACgl30M+zlsZsBB//4atTGN+pPXlaGEbHyDBsmoI57HyWcGqjfwO9GOPPpQFWk9F
XPCVD2u2/BOvsuJvGPQWB05qQ4qEV1wpGqnkpw8QJU6Rvp79OfQQLzGHTyvxpVyJ4fXcVm+iGI+6
FU23lb94Ze4b1J92eHvxaNLRbk4/KlJQBRE92S/doii4wj41PB2wnU476HCGErEWMuk0od9pmp0X
AZ5uRx7pRBtAPO0J3+sam6th5OtmfbZvJjSJ1dCxDOeiY4jS7hsCy2/LeStqj43Z406z1a8AJWU7
/vak2rsMyydl9BNcCCQtrTwB++gxQLWkUT++sgPQTmHSnYR+RIQvPPwo/eRdLdrGGKJz6qoY/K9l
Dji8V7ogTHy1x6HJnLdBUYtbzDyobEqorSUyw4iQAoAsHlvYX5WSI84nKxXatlxk6vJs+VI1xqMi
US3Uf4xAimuob1gUnUdS56WP6Yjqn/lE4rQeXo9WaJYz8kQEk641l7BZMrT8fSSzDgIQyUlhbv7f
DEnK99MBbzwWID03qghqcRQrD9okh8Qs7NY6DR6goecGAXR+UPSVIwdH6OX7/DXmUQJCi2LP9BE0
B8352Ej+gN2mSdjnR56S6RCrJ0MvIOEHmVGwTnl/8U2RXCaFyCZXEDnV+TIa9YuBQ+t67I3dBi9r
nsWgtqj3U8d2d6L+HBwaZPvOWZRLmSfsx6e/B5hoPiKZnCoHWnsAPNaFFivO0AeR3jIqYI7Top+5
vSyBpOlA9gj2MRg1FXFb+AC0DHHluRaZ21bMxeK7FmKIH/gXa7jUZu9gooOYOL11v8rR1m+bfki4
R+FKXBW8HfD1usD8NibuVXEP7hKolTzdkE3XtQVS6c0HgO3zmwj+jcA06rmoLUgTusCbjDEns+F4
8ZYUzjxZ1ewB+g17ZLzhmDRCvFA5LIQgX20cxTm/jZTEz+Mv/8GSGZDIYsEGf7LFtx/9y0H99Mnb
ZUoRedgrLxO7llKyYxB5Orzf/hMXZiSbtytuHB9F77HFsUuFEWdTsQxbYQKFCZLlEMz/MUi9C+HI
y05UUzeNZHlCZDRBJGunEdBVNCgkDx/zpD8DK5/VYtqVvTYBiBbFp18vdtTJ0VQ2UF6FXibpSPsI
+q8DXqerVuynB6kGqsCz0g+RR54EvkfNWEzwd1U4R9GDLaq6YmnSU42SM+Tjabrcm8RI7/RNGzLE
vWu650VdaIXMkuPxCSaDMOcRK77jYnOjigdP2jEBJN2zma41ie692Ks7AmAjVkYYhIVCEk7yw0hG
xS/w5g/Zj6MoEIWGzR4XyL2/fBw7OGLv3e9pEu8TyjEccbltTuHbWIDKyG2ztEX+VLrHVHKSMepN
HeMayUKcRaoe7YK6r99EqVGNyoF6BKiyUfm+dqk167MeRyq1NDwy15qTwpksEUmgq7T815SIYxQR
M1Fcj8GfeP0D7Wi93l8rMV6DDIvNsaBZXEBXTEkmmceQosbY8lB+Sze2ge50seV9jQSzPEVET5fB
ZphR0LPb0RXRQTI5FdkH1PZf9CKMGte80/w9DLDWNQQMBO5trBFV9UHmc8Zd5umZHPnTwuMHK9KL
v8MuA5fVD/iRsGxbs7OBH0OFODJD8z2OwOBRVd6w+67aCa1uKLOSTqymldqClUb2jY1rnH2bkkvy
kgNwsFLpesZW83KpJg5eK/7ySn5SczeJZ6e/tB71JzPvjrKKl/4RJ4jQXIJ5XYRJi2WOyIx+bnIA
tzZKFvVSc27jOeo/QnzFtDQsiLfQK+z6/YFW62u4m0VUpLMtcEY3qjPaO/msLYK00dYNl7bIzsKl
JBgTHxjC1T0OmjXD+L8Wg9lAuOtOg2KfHvvDsJyCD+KeaiIC5ffZwxu/Ozch7n98pxbwJJcK+6AE
f++ugqDhIjOhNbMasmqpiKq4Yr4iPRWowe4YILI9uPue0f4Uq/clAIVeM0e1vUtlUjIG87R+ka1F
UqqAncWO/JLg1KoEL4YEIK4lEgH7ABLjC0L2zoSytRH1lYfrhr6QmM2tALReShQo9EfTUBhn7Pv2
8IzhqjgB4mTHHB5nZhKD0lP7q6UfWniv0w0qPEXFntcFfcPv4hji4+m84R1FgB+NVm2kMuO9cVbu
TJhKV/qw9Om7qwtb65hBzcGQA2yfZX3Fa0sq9iOCA5x/qxMciIvS8pwlt8sNPtRH0RgEx24gSA07
HL1cWL9jOi38UHQxyxD40d2EsuX3HYwHUpF6EoRJGhEz3uvfWEAy/z+O7v/4v4apA969LSOBuGK6
sDvFvZZwd3/Hx8FPB7HUrpqyvPiJBCB7RKgcbDe2AZu4hVJ30TmqsGyBbgIGpXi4Ihx2hzhblPyR
n46R0jvf49J9NO497eIkKYqDcNbo/egGCnu0MRuUKZXPuikqDEuczNmVc0cy7WkSuTTcmnGPRlGV
6fn7N7TJU9YYqT/pRsAUgIxQIy1LhJSr7qlsd4TQA5gAAuF70Jxn7lAf1nCTnEwP0mP3c1uddgXM
vCOT9j2TepWOJoEwulcHyLmAiGCZwsGLhe0KG+eE9od1Q7SrTg5QUqW9+YSYIA/DXkD7FAaz4S1U
i34jF+oES1TAWvCkLcvNXm53XK2RPzJY1m1rz08UDrC0btBfs1dBbE8tRGRrdopypI4AS+zZYuy8
sPczqicIQQj2vQsCxa/MZIwIoPD02cynWEBAQQgvZsOC52aUWLzLhJdSVducweCgNgJDaBli/4lm
wp3nWIZcpBPhSEUKiMRxbCpWXxnD3c8jEndbS7LHKj2mWOOVH8Yt8Pq60A7loqKH2qmEvqW3Hg8F
uHhMxKUEwfZcBheG1kFHWAWxCePa+kwdBlwqEESbcGhqadT8/0EDI50a25vQ5hD/+5/lvyBBAqtR
GxjdsYGJJgFnzEHfugteTU3ULD6GnE6KoqccuNHLhnZTPNTLpLpugVU4OCAVopWAMzCXmR0qNfLG
iqSCRWbw8SqXqy7ucnjh+ikce/fWxpmmMM6M839Iz6btiftzRneQ6CbgvXnHxwpwRh+pzyS8NmSZ
WXJ5kmJaKAEFmG9dSZooWYoLfNlEPOIyypn7GCk+8BOnW8qfCfC2PycMyn+hlZRYstYAeIVk8Wn9
9uINKfGZiX7zIH7K92+64v5VuuuEybWiRfu6tZea9zuQqukv9vHaApe2TBe036eOUEheWW0FuR4Q
msW/zr0fNbe2NMkegHYzYLYGGhCdnxej10J4Qbbf2qmHQVbnJHC4C3fMcSUdcaxRnCBDcG0sYztM
iFsFnxHTmFMNkkucaLcKnzGlgUqnK3fVCsTyN7EOwpIRIqBY0HZ4I7ZVhdaXXeGmY2gKTyTcgeDL
a6Ykm8c2klfjX6nH+YtlzBzgsvGEBr3HIibgs3ehyD/LGnrjKDBiqtiqfTXFPeCPz9ZjPlcf5KqQ
9ql2uosuJp78be/JRZY3d6njC2MaEUEJ9EinQT4Qmr9H3OydpdQ2Vh5m7+XVa8OUmRRWNGlcWmPS
J1RlsGRhV7c2zO0qWHOglp3oAnLPIqrDX20iA4jtz9/DrJD1XaidRJNQrRtF6XbfPNcdLrNFDQnY
dyTp1elzQjPDeYWJsvU5Frf7Qe8uOC17XQfo5IW2NS8WLq2ae1nldIho5lBorCdS5Mqu9qSyK6Wd
Inxi6qZP9WdOGQlbfXNuMyhGYp21iNIeCQICR74XkqUmjhhDlOh5ZPUMztsdvI9umVUPA2NKR7jH
Zn7UQsMvIgM6qUbtvu6F6bGB/Oa/qXW+dmSFqbSNy9HMu7SHKvN7llYzlMLrA9n1sncT4kg3G2Ub
sLkA6EyJ1GoL7a243IFGwUZAiTmi8CfX42kUkGwqxsuohf8MTRv90pCGs+R2VFnrEI40Gj8fZRAI
H0ItIW3FpLMDyoW0uO2OWDvUx7F5BWmp8YRYMn12OMSaKG44IYRwh6Ts6G1sjb2QtlWgZhtgxlxZ
BDGJin8kn51KOSzCk+IigFdmczKt5qIt5CeuvTo6Aps2uSYcLTv3lkyAFeWWSpJFTCAf5BkzXVcn
nLbS4UjHU1nMZhTIgn3TjxjcapsAwEOv83/QuhAbF0YvJDLvTFlvLCYiXVPl4ugZAkBsx4EjnRFY
MiBOU8mMDjYJEHXdm3Zmi0Y/k3rdseCm/mSWE0hAgVFpH88ome1h0tL5tc+Nu/o+0ezZRxvtK/a0
dyVwpOwt4WzFZ52dyfzmgY0QcY8PqrjBlkcLzg2WFCSBKvW7hYPp35emOk3cGjdDLMhnw8YShpJh
bbv1RAnH2c05ztqv6x8rP4QDp14Jwstt8TEoymrute8+nLklrqfXygNtQRcL9d7ZQr6zrFcv+8p2
fudCCRmsRZpC2MD7+T3iYdkUgPuI35xsRzUWVbKWHCfFnfmZJIF8EaBt2NfB7KiF0cdV3MLCoVfe
Ui2uLpFH01FEbMzV7hx3gmF3rXB8HN8JANLAwmZ5VtlVlEMBwF5ngEICBObtOTy9/JPx6ZjmlZIS
/FUiNBDeriGRE1n5da6jTkpTUFMmfLJpzJ5dAQvjC4TOlbfeK/M6oSisVeMo/c/+O57Rt2J7aeer
G17F8gShJ7n4SN3pE9jjv3Ptv593m1WPpkjfGvB6ur+yOuNVqNcNuDxIcCtivH+DJll7JJNkqUA+
qRf+EXuLa+lCiRucAVvCak7seOrCuvPp6ZI2xj7B1LuxCWMTkxi6aW01yxWI2VM85eoc4IhRKDVh
mJxz0muWCGIzSSFOeSya4cbKqnS5day9P/EPjTA1VzmVrAYVyt6/bml0kZMrOgd8LXZyNbRygNFt
KeQbTZvykQZVZPjhftnjpGiZ+RUHjKJGikWyHHnIXhSBC6UtQPfFMeMykM3k2vL+Ly9aEIylkrz8
S1hq2HBG/6tbJtK9wNrBIMFFEBCEBpkAPifIEkv+rfW4isyFrD6SGf0NEJiGUGmSgNSgu0eNRqnE
fnXp1Zhp61cXOJ1Fp5YaDZf8cf0dmZbmmiFYqkDG0zSlLyFYUHZYnmrHjrG+4b/u3sEpEjLYklDe
OL3+uJ7McrSCixL6VBqboqWzB0+xXcFMBAyRGsVMGui7wu8zUvxMdbPCo3vNlIUyrQdLuxVJw1SG
jidHaVA2FApI2PIHzyTJdIZSj2R+pcBqgB/2lHdVjM59BxyCcLkcX3WmdAwY43FsGgtQ2nS1upNc
cj/f4AhucRWAZ9XsOKwLAo0UZ4pUvB9MAcxbBho3ft5SIqxTk8Tbc7yyhNAGFgOC/0VB5njenN/X
2g11IdCY0Lzso2OA1vzawtoFyXgWrotMHuB9RMfkNtLvTG0R7gWl3whbDLirZh5t6RZ+HOPH7KYo
OTTmn571LQzoEId7QK1S8LWaZgAmENECptQNHcIwhI2INLpHw7FUEjlbPpqudv2XiG48Yz2ldWtg
90pf7NT5xiSvurHQzaT4yra1eYVQTyZu8H4tQhWWGKEC5suetZAZLQmOquzATOu20Xqm1LCW1lvT
wKSsV4GQt6S2LROVQ8QQnrYTOOa+h+pudjZiwrbZ4XaPpTHCyV0WMo/psuD15DI7TiMZECGrsCxe
20Yb7N35wnbqV6p5OaNtw7GhgMSI5f176PkI3z7AG8x3w/XVf7v4W8iMDUe6JrUXpXA1OBfGUzz6
8yZnGkqM6CfbE8Bb83TfHQruvaWb6YZi4PEeO138SgfvD4wSeijAHD4gZrE1PCMy9xW52L6P+tQd
hex5/5FlU//hpnGsUv6rf3LmbxFxSf1rcPQxZWYsRW+nvwFiyBsvP59DHUKq+K4qXdqs1YFefQVW
mX6oX2iYmDgQkkk+b4k1JFjYP6XZGQ8NRRHjuauBnQVSa0eh2jtFUHdR3wx88mfUlXVfad4I0ecW
x/LaqUMJCqOLjlehmLZvUcY7U2OENsXdh97Ykiw2ICg63Yq7qVuCHGNAMbfaJBjFiELozJ2XXHI6
W6hv5QvXHPTpqBePB5rokW1qqPjJh+XBEAM+BNnwWzNr+qT5Tia8wNUtzklPvBw5IkIvTht0bwQE
tzii7+kz9jGl8L6sGC9suGx75cwQgHSkRG6bzQzzIk73xjIasfZ4oH/K3UoofVyT7UJYqBandOa+
rMco9OTSe6vV4wr6+o1e02NVXuZm6XG6BddTC/6JnJA1QityHQ57yjkFQE3aseprE0roLDEcDTHS
iMIXTyUFGzvMWVxHZZezT1p9rjnED5SGc3+AEfhyups/1+Dl5xIUtLLyOB9OqZLdEAzBosoADN9n
3a/x7WHEsYROHKzYMVQmoiOiqGwrer4e5n1h6fw2virEa8iOAwerY/w5QGmLdR5RVH3IPLDfkFlK
zuHBqeFTHMeQmURtN8ASItukXtJ4wCgLI6vNqS+cVsXra8qaQ9niTlyJyVSus2oPVCVIEgG7nHaG
47NtaiPU59jjyf6fNQlu6Mx7852/2ysmbdnctixt58tAU4P1jbclqsG7S5a5YAdUb4eqabaKhWir
81DzrBFhEhjihlsvLjTQEa7RpaXnKVo8jEuYoG7h44wuNP4KjS8Vr7084zsa4Y/z2nfaMGJ1zUW2
H7Pbu1hQpn5BvyktZCAaqHu88xYoBVihQkHGzF115dcBr4vUEAQot2Et1u8gjo4/Wd5ucSfctrkj
xvCFHAHh6fLH/XLnHHnxuK9zKhccImJFNpZytKdGfBDKvJnbsa0qICg7iUOVxf6uRpk+8NOFmL7K
42+7A+0Lut/ftlh3u+iwcPWzc+0beeOVfDOyI+mKJ618Pi9L6GqmfANIvzLTnYKp2iWC5S1hNPi8
+29okIUJLvCdKP4YFGgFiz6PdWJQ9pX4cvp1YaUGRTj/e4ZUfOR6/Fq7RfKGde7DyDPllIqv7hTg
+8AYpXEhnBHRAuMJKh7NQQLnxY5TCbDANsAoWqm3f4Pw4jM3PE6dY7x26XEBKJ7kKmPCkzCEXhlI
a4SpS8BDI+m+6T1NozRviJr5AcIsQxm8UwD/fW2BKMAowxBAJRg4S9S9FQ6QLfJsOJRipMsFlthe
goOIhWxr4ZmTDSm2APClt5R3dsGh1gzspgoe57NMt0+dxFJTgj4jqAvvQTC8NKOHarc9090GW/kv
q4feccPsQcVDAVBCq3WaZZydES3+ZZW1FJAmwB+BFqlC0R3jfSKdCtSE3q4gq1+LHHGBdqQkgRe7
dLnk7/5KfB/Wj1nDNB77LceG/ZtBkhHd0RgQL1AiCMNa4jcQM6KTlyj47NWt7vW5VRMvy3Lrcmdt
MTuV4QoC/7jUnLrKHEUzIU0emTFgmU2bxv7t5DJZfXemEpbm2R6wNzLFlvyWyu0viOKwJe2ABLu1
SIzj4BwbtUbbsLB4kELAC4V63PjYjELgBCiqmL9LiBo8LQJHM83e1SwlMOepyTJ2G+mBLLDYyQBk
5Wtd1NM2/Zeu5ngWKXdRAvUVS4c9SNjicxLNliZYmATc3jo4dtgynrlC0mYeJrgtck+MrpBwX/4J
pvfyx+cRHre36dYYDpekxsxYM9heWL15gmbd2bOLK7J27Ne17HpsXyZwQ2Bf/+mV7NMyqXnTwZot
FaR9sllXDySlCYhSM3cS6UNINOe9mjS5xo9mqXmG9Ac2Dwe9TTtZo8yLu+PkQYOLf1hVz3iZOJgC
rvOaaaWHOhwoza6orCamA/uRT9MjV2lNhw7DV8XvPGfb0pqQ9yU0o9IXyg1UdTQ6ao/WKFuqoHTo
i8yjnqEItET6Obi4egWX6x75llDeCJHX8Xz55fpaG3+8OI1QpGeFSfIXN2F+pXU2VO5PWvow+cwV
SDQeP4isn2GER71gfSiyO5cjmK16+zVuz/15diKSO5xkcrhmzB8raq+ct5eFKc/G61LnTP3wRR4h
EIeuCvJ41Bi+fa/KYnemBSjz36Vcm43WVMsZdJerQKOTkftpCnN5SXTA/sJlCpivUb5OKX4Ifmfk
gZo/3j289fl9HhGZ2bEYrW4tCQAHUaIFrQ8pTOGwu05fdy8u8wGP4ApQadf5HZi+pQanZpXsC89e
4Q3s72sT+LUx1cVZlzPQcxBMWZPJBuIlz3FT/ds0qUiG2CbYKXzlnqp0moSFdtgeLOGfndIfdRzT
2emgDWM4wUUbuA5JNDbnigmZciSM0c6iuaGwlM1j63RukQMkZ+8yIV/BN96E2ySjWBB277P1VvgN
UsNyKb2HjLgPEU1OgLNNO/zATuwUS2ybDuehdrFp8zZU1r6BaZT1Tppxn7hxIwa9RE0UgsxW8cBJ
hmqJ5gEEWbqcofwC8I2Ee58QsmDfm34DBXDFIW2JHbjVfwXqRvMok6zoVfZmHgEV6yroupINR2W+
phXcw6n9GmynUnNgF7e5yXn4I1XJDdmoCGlgCVV9LDuXfc2cpgLGew4GmV71DSbf48UmNklZVBbv
SNF2reeU3y/bIs/fI9wEwOFB+cVzn1yK0rdYR4KR++hqJQ1YnuMDZyAp84vpsYuTXKbL9+r+BUsc
WOVb0ByhSc0QWKvarA2tOpKiLqmh8+5Z6ahgUZ3TZDqo3r+jFPbUJr67nk4jmC7f5V6zbew9WC7F
4vCevOTK9yY2wSF4p4C1+V1nwZo6rXVGb+VrgY7LnWYqWvDlhejBzUZDkGjPD/jBxmenXZM7GPcO
3S8pT0aD7OFwIAN78BtJmiP/4LcNXTDsFYjyE+LNb/S0vU3GwCsSKM9x9n9Ynd3U5CMY4ormlKCf
mbaCmOJQbYvqcogMqr7mH4hRBvn7apql1qi98pKNp9SQaFFyn+Z845Rx5QqNTDEOCetc9Iqm3bhm
TqHj/c6rX9un0OmUxz3ru4Fjru1q33nuC50J6Lfht8grZLgpPdbH4Zr6gQnIbpl/O4OnilkLQx0u
IIfn+1TjtqDS/FANgy88JUul6g1wo50+WZT5dffq2HDYyPgGpSWxexxuglrUZ8GTj963InOQyMlI
GF28bhe7e4DT682eykYHkUqXtp6t2Bm7xtcgRf3R3aUT+tgdISoDKcAT1+VMJZBV0iSbD+xaLuo8
HxCLOzfVwuF4ZGNANSYPQINfqSaXSd6WSIkAQyKFGYcN0HAVJOifJWE6GxKnGm+4IJ8aIc1OKH3Z
8w7ZZ6FKjdfyxhmxk6xgQYJO9xaOMXgjzo280IShgSZm2n+YPeiTH/V6Mir+rXbSmPLDaWZg7YVY
ADhYOtnSlKruZhXHPRQ88dCqR4m4is/79d0nBwYwNhHCkmp00Y4I+6VAEWtziopVM2fPRjU1UzJK
wIJGCdUfYPyNEzJPHXumb7OMo03EuibxDnnScQSMKlsRLvRasdF2cdX55W4jw8zKRTzWv2PvZXK/
txpr4qf6by90BFZBPAUXUqBL7nCU2GLeqyXrFRX/Vam34pUqe5F3u2jpvmcwtf8TmAtEpOD+3OaB
Oc6amFx14KMszfSTxCmh4NwVqJUzptvO/YrOa9Az+/lL9+wer093xh2n8/ZFvn2X5XclCycpHpWY
MJtspsBJHR8uQSJnXYXwTKLq09wO9nSCaUQv4GqDxe2LaOrXFQDBPVS/d3T5iHZTjwgY+/R27stn
iQoYIbL66F3yQYdOAl5wludYU891F0S97RC3mi/21Tw+6AFfmNeSAhiRJxZhKC0sjiqSGd+hiVii
RKebcrTA2h+HlWpAKF1yO8O9yInFN1fQeyhXMeFQmPk/L5Atp77j0rNu7oGC7trDs6/tTtbZ7gvk
VRLwNnvfH9E0s2IaU5inagVy9HPZojiazNQWk5R+UIk0ClgZ20wK3toaODpAiE+FjLLdTDoKrgWE
ATX8QQlwzvM++PLUK6b1YJkxfKoq6YufOz0y7e2hkqU1VVcUwpzo/eJGToW8qLzsinuNa3+U03M1
hMBYvGckMtSuyqhdsBXI7vSIeusKWN5H2rhN/TWUzhxlmGKrSlh38IjXyb8xv8yuVKIiGFd4XxI8
Ml+AJmmQgHxVJtBlFAt9eXAO4aNJm4y7Vkb4r7VeeIwanT2Kzp1cdWOG4CsZYF569zgElpqUQ3Xd
JakVsTna/Lr4fp2DfZX4MszlCFFPOnvArmOHz2W2gy6J03YM8XSFCwtBwAcxAdx/JOxx9s9odSnX
iYk1gWr13z6AglXlAVHVPJ/7Q034OkwPz/1sYuIMHOP9Ox82eUMiQvhzxLdpOUDJm7PEsUmIobrQ
IvJg0T++ILUXasat7bkrr0ex0UNPzwk3GkwriC4aebKbqeQht2oU6eyr5nytuRiIlP4iRac8v3mv
+dTItj+sw0o4G1T/XwHa43oBb7SWWMKwoxniHtiO1VGWj57m2adC8neBi9+dxI37Q0gUZKM9/7jy
TNLEXWTisaLRirxCJmAgfgUErsAE8fFEE3zuYY93le25goWch8XV9dxLXZYxRxOpCINJs7Tgffcx
oUwDnBj/I8LbGIqJIb8VggIzm5jCt11nzT99F/MdNHr0ixQ7CW2sq37CXmwurgUI+Lvq9oZ98Nz8
8sc9d3kLH5PkjgJ1Y1Sv0F4uZ3wubOiswkJJmGmqrVg97MjHdc/2O7JqpGpjuH5VX94I1y08X6ur
iauqRdq2bkqpqRu8hYaj/ZSEjUW1/pcURuRq0Jj36Y5th2+YCV4ztRrNjiuBABgbYNH/mZhFYKSC
C9zie5S2uhPoeENHDQh+BgX0+E+P/M/CxumooOCQ5Wn/UPPGyHtOHtq4oU1DrsknSDQbbT8nWFfh
JGSZ+u4cYRoMHVYhLU7kVrBAMRklSw127x/UR4OL6pNeoNmSGZQ1Ji4In4RWgeCQLMj2kAGFDrHS
knteK4XruiqIpJRHScPPj7RLpAzVAtSmUoHerOzQMmXRRIBj//KsSH62sE+oaj/XJSuGbrIMv44p
pxYQD37X53VS/nxLwwbv1SmDzD6tWNxTyuN8oVwffnvfRaELw9c5yDqkW2XPQJnrluH+jPWAxKho
cUkJMKQ/IehOhnIrdPpYLmE+mtvmQoNkv9Kxtvggr9l6mDi1/zodzl92ZBZyYVipiRhDJII5oWd/
VtLgVCIZyVpff+qDaIt4+oztTFfBDwpm+IP6fcNi+wyH0xnoGsNfuCfoLFHrsltjNYEtYZpgB5dA
89S2XOVTYEoxQeFKJRURY99GqB2qVSylEFhgU8qY6Ju2DLI9PK/xTxu9oiAflgL7UkW+9iUMpmhF
eKHYQklx6KbyjraGn7v7dgy+AHpy8Vkdco+1NzvSdxM6YGMIXDfDl6cdARX8wDo30CqoATne0Bx9
HJCK+trsW+MA3vrRk2JjQytlf80rKJvTh/fJTFE5foue60NmaF19NCUPn13kcGtY4jPuAy0kmKrZ
wy+Za62B46IwTt7ob5V3cU/0VATds0VKDEw+aehmmlCqDuYnhi3fRLwA/Qgz7dRHSRuJZ7TDD/pn
rkR9q5GpILxWi24hc0depGHPso2/QP9gf3vFdfN8TO81cs+3zIRayzBugVTLBtC073wglsLxH5Up
74+txj2zAniI5/mcV/QySuFyKTLAXFxaXWhiTgxJwRzRWBtliuh7bWfDxixO8iBXZ1DfPaEhMI7D
GSkVOLFze27cls15PjE2eAozXSJkZY4XwPofc8xPYGr/Mvh05t/uLNvzyvxlgTJbN70cmkMJakvW
urngOGdOcQuT4XcA1E8ZTj8V7VXI+LDQZCKVZI8MIVxFKQGu5AgCffx7Iid21/Hk4orh1LyLeKSb
OQxMIlYEHWtuQiTimp502pFDw4PtpuN/rBDEzPSPEcC+cjfkTWjPT1jHRMUC15BarC8Y1b/PWOBE
ZyjOFYI9yVkHr61RGBkeE0VaD2DB7YP6uKRa7OidukT0XKK21HkKLkP++H4fCEg9Uv5LT8F7JYqT
KOlqSBry8YYHdS7u/KnAxfOVR3qiACcrRLhsLRJ+1YdaNwdPC3e2m7xyQgW1aaQwAa8PURvcekBe
ZZgoeMQs+z2VXQs2wHjZMQ6I9sjNytoChwLsNVJ4FbG1pL5tltkpOjMLXSu3T3A8GAM0Od+MVZyk
HlkGOoBDgX2e1xMRgfMquIcamddyu4wTkKw15wCIJhL7u+lwnfa01S9gBhhCBaX7WkA+I2F5LWYM
H4hj+64sstkSu6+HYXYuBDLWGcHaYXnRzyPxSb6onshsw6dgqpxbfmc5Q5lgiqQHi3fAGpY29Do8
bHch4Mvi/xdBbwZ79m5uKZVI1lMl7JmR9Y87UiRGiMmoUZTZPzeRRQdc8DgD9+4evtABnRdfPEGT
xQhGvS1YffuC5x0SyLDdcM5V//T23lFylIB2KIHN70BDc6r5ywwSRQIWXyL1PM6iYLQ0invb4s/N
3HMvHAoctNXqdz0G3UNGF91kVPQkvp2DgG2WJtBAAJyL4SfV3SqO9qR7KFa6hyX9Wy71QhF5kmFg
TsQ2hICdxuMRqaBEHyLc8GU2+0FDYmykk5fR4tFRm0b5edQCJ6au3szIKbOsZ8T4udJF32D79xTl
Xs1LLRvHPcd7vM4MYPxyvQgEYsNao3e0BBz4XesSU4m1nscMLJRYPamY+g6ddVoumVkPpqg6czym
eN8ytDGLzQv/4dfe8noIY6za2NKTPzH+0PwPCIfoTtBQ/EgAZkI3kAH7et4Iyd7bLpG1WWPecLup
DH81PQ64tRVjwfgL1txl86Os2biOJdb1zoj0J7DfjR9r+Ixq0S5gGsR8unLxaVynavtu/ghs4GZv
SH7uei/jpsAIrix9Qhy3akjd4I+8tXk6s/WZFUeeS43FMzTj79Yg2aRnklWTyCVQ+v1ZhuOQXcYh
O+OhD9f/21c9Po85OtQfX5vKHcWakdfH/1jLQ0LbycMHVISwsyxfT1aZcMkuAu6G1qcyIVQMuiUl
nGI0Yrn8hiAVEWuQE9cX+aIL+E8ecNWtPF7SwhF/4BprHAZlRmni/BKBeQ4fnxWn0sHdyo2k4UpK
aidR8F3sGdlAHhmvOBP0OPHctsZazTwZjkx5h7a7W422IGGiPZKvIpUrGuuy49PzmOWcarW68noZ
uBsobJMoaW4CFMLhjTaIVoLhXogVT6q4hoX9D1PQCKHtMgrmpB3Zn/BphKVmGIlPGHusTXv5UvJn
bAY8pgMfs8ohbcKn5bJCpWdQrzZcm2iOxJSOIjqiA+vrGeCYT+2+uMn8xyLlqGTOUShNdY3Yqwkx
r3NB2cH8Y2I1kHkI/B106BLX2YVIddjyPcLopvOHP802y8lqndoq1a9XhXjUOBypsdjAarb21Yxc
jANx4fFHuVEzUEfvHwyjuQVp5H20yJ0DMJqf6y38VKpXPllva2Kph/avoYSwXW0DCS/kNsfxr1vG
W++Ur176lZFv2/kgVrnTQL5ExiEuoWhlPfefmIenrUQz9CTXeanLTLBZAfO9whcNJDXp/oGw1GoS
KoEReNkiBvupTzmmbV1IunhHH9pt9xeZLlTwF+Kp2nZeZeD5sFRHG96tOBNIkwUZDOp/zgx9RojC
sbEIIgdugidE1Yh+6K9BMAel3U6T8CbWxKbVLjk6/Kjt3LmmWI2xIwrGFqkmPwYboenyO9FIIMTq
rb135DI6895Dw18yWatKOqZGq1VoMtRD45uFx3tWC0WAQyrMlUvOogCDkyjxPSgsTnHVEKhG2wZJ
MogYbqWIujKbt6Xziko7Vh8Ajh8BbcasTwii8XDBn+s1zQ2GUSxernBGB2enwrnNBlAYZ8cKYUTE
3ulI6a5YJoY1ae34AdIuZ/14b7apoD3OhsN0PSfBv1xx2FBmVIKxdlMf/yhOU8dchI7CojL1gqpd
o2A7CtnaBv5SGBdsLODN8nqQSL9CMrXpOVbRdx9pJi1dejHZ1dFC/1PI6Q5HPdMIIRz7WzmslLPG
nKdsdEn0G/1f/WejDJSn1Ib4/iYmFsjIweWYD3KP/Q+B6jok2ua/t/CmPtkQfC73mKKbt1m6h9Of
xc6RwNKO6L9sRx2BAvJXBlTZC5JbUS/y5lemugw/kAYmR1LFRN/AETbVknYn3dZlw5+gC+2axYem
3HyQatbddZ4nZhEpbPlTbnt9zciUMRYgwGFowoth8fTNG9girsB+UDUqa6xHUPXfb9X33cYWXIuB
9kxrUq+LA27dLSmyCiuJciIX9GHXcwomJ+7S3FGG0wr7C6BEUA/m2F61srtCCgZlsFEgLFHVBKcQ
dKTsiryfQIzFHCgiJX9HE8vfYVYdy34BiZ4Fm4ZwjP+jI4Q7cegQw2TfaoOgh88I2Mn3ssxI8D88
L5gEbAtqMz9QGbikNFetXo4hC4u7kAPgCSsSmdvQIpDClDr+7blzUhro3r6KmlBI3cBI+NCNRVEt
FDzGilWpV8B4fS+jpR8ZCb8IyB21Lap6YDJxDsHHGnf7ZE9++0ADJKHDqIhkW5MKg16Ay0HIOgMt
hWGModwphS00AgHKPxOxlkJANkCwKA+zVi3CSemH+b8uNEGpHkjFn/4mW6dT3UdS5RcgVDzkQ9d+
JJroxpKivPXYb7Tp3rsjqsK6UJKXsGDb205/asnrE85UqL4z7NCmroYnApXbXHnz3fSfwY0S9wtS
NuLUWiX6gbZsDb2KTmmaE2x4H1BW3SjJvKTl90iCXOjGAhWXTEESV/dKeKvvAj/LLNVKfnAiD6VH
7BdBXUA6q80bnVR9p4loWxVaJ5tCQSgCjL+Oxq+iUkcq+smrPlek7KWt9KA2Z/HahwEWWMB7wemK
bOPZCgJAc5DDDprAmBwtN1naNx7+00MgXr/H6aocLc7YFKv+x2LaNVd5CZAP/uIdqlaVyw5tO+IA
Pn61FZ8DEFUG7GAd8Ek6hUqK2MH5BhbXZYRvvG+Ri82BAjl7vChQdRBGKHsfAXVeuBpMHkgfGcL3
/J1OeGD1vxAGGnXj8SHJ2zoAIcdcK1k9bdVwxTfHm7PbP1RvWlJ2M8bqNkuUU/YA/RzyV+TvWmCG
bbyf8hCpXewiL0WYpyi/YiBtX+bL9LMEUN8on0G1CAKlol1UzMXox9g3BvNKGHzSP+YflQaX4Sy9
Culvwys1PMNAmmy9fqrciavyTMzBL0TemJmeRHJx3TIwQbQSsmBjNCgl/+I7HGxMkPHy1/tgUvPM
YitEpMmAzpveY8FgOtWxacEsHhXCsj60cx4d/qVgIC0P6kHLBOPPxi7h//cqtOPeXNMcs0tm0sGC
ojCrWduyVghX8cRkiIBBOr9jW5kbeHq17n1tiV+IBRrJ97BNupjrbRZabNQ8QzebQ4eGZby8x5Dq
T2kXSE0xLLBVDXtZLQgpo74sltQQRE+IVpyl3UFHoUls4v1qG+c/sMRUcpI1VNbi21IiMlyBV3Hj
elAnHedqMUK8gOyskmgWFiUoAwwK5t0idk5Xex5aRO6YnsOmPTZaYWvUjRr3javUmygvzRX/0aRG
+xx8Cqg4p1ahDIRcixHTP/3bD02OYWEXup/YYzGLYfHWhe/XPHbCOZDIS8BbvTJ2xjsjKqPiqHGz
IL6R8D/PPv/OzjmyTbXCP6EmTUw0xGG8WgQ6dfJ9qlLy7uOp7lIpsAJ4wAUhbEwgBnPwvT215YFc
DI6kx+Jb0D1N6Yx65JVUPaVNKo5rjTAk12aGaMDDGBzaPd+QHhXKKJ6+dLhvKGdtkvnMriOpinLR
EqJtiXPYA1VrwcNu2W5vGU6G8VVICzpy9zQIqZuJXOato8SPFIELRk5QB1hSWdwS7BvVb6lkGF9x
vUZ3il6roQkTnNJp68vtN0wfUGsYHJOFLH4zS3Mtpl7UGyarzEyUKuWDam4xXSWrdLmiWsetoQxe
Kv2wkkTXl41l3k6tfBoZbnzCM7myqTVQ2V+MsGLRf8B0DVM8Kb/hJgWuzcpyRwYsHYZyPlncRLFK
veZJ87cYHEapRzt+b9m8uewplkpVUkNwAaeSj6bXAntMIZXBV6UQ7X2UEi28RD595WQz73Eddbxq
rA/nVk9RG4Mi19dGY3k+QTMEqJBbBHjBFm+WmQ3GU5giayAalPesx6zZ3HipwKqyfign8+nZTuHH
IbzYvSPj2xzJ7mxBiUeXdB4KspQcs/5BC+RIWfoCwVeFKxdqhQwnxs5LWyXZ5BjsPHbnYoq1UX8U
if8ikgIyNg3PQlJGbou7kAnrCFZNMqhgMnwx2P+9XotwOGOPuAB9GNFivUXV7qq/0jJPrqSTqubv
w1Njb+tzlWsPlYPLuMdpVMmtytlgQbugzVMpVLfVtL6L2gVtOOU5JPxaV2d9ks9iDjJlSMMAB4ss
a2JEvLKBAnZESu1+Fna+gDobg0iX/xiYh5pIRujIltf2ZgpyCFg79Bqz7g+tl2R0J7F4fq/EYEMU
kYY0EEXbmTI3D42ghawMVRWdcWFKy6JRn/3bsIVOoEJOWExTZTrw3lQ/j4L8bO2BmZu5+LOwiEtc
JWUYSAFCy/H0uoFR3moRxeYe8kQQGLRotExljSaqzV3cO+KhIQT9rOrv8zVPnraBx/JwyzFbbud1
p3Xdko/tE4jKWQY008f4OIMzXJa3dzgJ5w1+8kI1b9Tq0N7P2UAllhDbDapUEXU6QDuWiSvEGhpE
LIi9iXOTmR6NnDwn3eJiZlSn9yQEd666/G49ovSXxamuR4kRvoKAbX6mhpFebHj9CHLn/fbuycKj
y/W1aaSLdGLsouPCBgO9QIelCimDoOdlKai7+fHuufQIrEp9tlRFbG9gJzHMGfaipNeBD47vqO5c
jFjqOBN+b7BW04nyzPNp00nIKcz4mZFAY7WeYIiRVSTmOlYnn0XrBvcH2/hkfHmMaMXiSDHlyb+V
gDp2DvccvGlLFv4HokxBBZYIz2NFn6oBINuwtjJ18uF+DhEHAbAK8aIqs0gfxh+L2KAlBTghMRWx
OFMVF38wBpCT9JTgp/gzul/2TyAlxmB54qO18xslicy9uPriGIQgGyiPXmlI4Q/VFjNHEZ+RF+TE
1bPE3FazunqIDFtl7yngc3TIhKhwUwAePATievOo8cXElBn1t9yLfdbM3ioneXd1Q216Cn8hisDw
CbKCXaeFU+vXssfb+9p0wR7L28YvH7y5DugSsdfiGqtnWdYgX2gUExIhCrf0EvYX3RYiMcLGKe7A
wuW0L9Pf7ZqGNOMZt7bASx2WrS47Nz1Dvtle2uMaAeCpPDNpDcCbWRSmC+mv8O4yav5j54oGcqjY
XXRl6bPwK4Zl/9vrnMZ3AE9BPcuKN4jRizX7oooZGDKFW8xPMep3EglfoA16zgnF24Kh4Fy1BHfZ
Ho/QJVB9rSmgHLr/EiMjHhHHuf6lGQ9xxTzyFGUQbTRUlcIAtKwZYYAiap7gwuomvPjYlBM8de7F
1qMK6XTPnTBL/rI0tUFOR4NIGJWx6bEcwSGP1xszjKvaeFlb6uoH6qOpgjDKgYl19jsve8aMayJm
N/1sVXiR+x5t/mEHUuiPk1AyD55jwrfo3INJ6Sj9DSlZZxzf7nS8NmLz1IGqIVrrk6rHxzxIBv5C
mV+r87YFnT8gv8559uJkX215DgVwDfO0ZFpjU4wccPo9/PtgNeQn3EGHe4X8Rk3kyie42eI/lVSg
0kT9r2l3Q5Kk0yGgnW2wRAH5FGxlAC0oAtpO6+OphP/snRHoXXc/ibvUIVv6HRYncbAG+1xFunpT
B6wRAs1PY6m701u7foTYZcd4Ug6GyExgEP52YTDCY39DwTGinNKlGECsxSJlPfQ1keSHLhXJSZVF
RVtckHN+0kJIYW0DenT11HU158C8sumg7VkTJUizBG+psa0PKkc/VEsRFTvgEoP+to5zHdgccdgb
NL7M8fN6PWG3pGugUoWtzAu+/CMh5CUguaRwEiNYDcPFT50BWfd3/v82B8eslvEoNqBJ/hEoAdMb
JxnLy+W+uJuCRtCS8wiKTcvgmnr6RKuQh5X+Xxw+ds72L0chayeCxB9pNiKiNwsMsfsY8mVP8vlt
fcw5xjazmov9MrxUZ0pxLuABZsMkXwOUmsRNgDnFeHzq9j422y/68sHvZ1evTSST24Dq1rgTIjsY
EuCneiVI++iVz5mBH8r2/PSE7CuAw2qQyXEn4FxVs71NAm+Vl7PxRiGT74fdujoOLXBUDEZ1gYys
Blu2pEgpUkiIByovS8ZH+6/gJhlJ2shPqoJxsq0x+NKNVLItXv9ev/ZNPu1XGHERRsNROxk/o3nA
K7ekrk0NX0LVADN/aRxL8xAM8OZPDBT2wdSs7+5B/UHkDRfXH0SHiSH+FPIfJLgWaiiJ8LPon4Gl
QOmzyOwQrQ1xbnPxOTAoy6uNZCstYBBMwJaSBXVjb6BbiXu3DSnSVEyD3MZCUJYD3Bv5QpKeKXde
yFAsC69TJvVywwOV1wqf1l1pAQLl8IdeZMcrNhnCMoexMGMWgCF3q3HiTFJCAi6UTHjRqnMosNfn
0yl/InjQVJLXwry0+VvpuVQ6KqZXya0rUDThYyuyvIPWv5Y+GBG1ShSXGxOegLZeCBlopecoqckv
72mdJoiMcv6ny7KskuMkZIOOLXbn8kIysjgRPnAJx3k16KmQC/UzJoc1Kwry1anbpvr/oV+5CCSx
PhQ0YXzkJ+QCLcKEKxSolDDl5kHdlAOjpzmm/VyCLo7xp2d5Y9TsoXjsyMl/vAEXNfDc/DUrVnSs
fv+6nXPR5PzBa4U8lO0UFNVM+Cypl8+3PpV0snS9YtdvjT1tMFx+ARQKlU3MeKsWDxLRwIXdPm6h
Aup++UghipdmOV5N6HGCuhqLK0uG6SCuvOOtJm1rEShWZ6cawjGrUbspBOMr86UpdLxhTi76cejy
gi70X5hYwDDyErmIGinHk5US9On4pjsI1BqK9UtaGeACZBBkHx9U1RdZshijBucmY+QVnN6iamus
/W11bZFlI+vxNMzvWwmfUGeu63L75G9tCF2cb9FlhmTmwak5DZNGdRMDBbG6ApHF8B0T4i6FeOKI
IMj43MQ03V+2oe7fDM3tlZEL9b1dfGn4H4sGySdqp0x63e4+ABWcdI+aGgeDtz30oGqGrm9rUa4F
40AllqHcMtsA/7zpWd89H98sfwKRgx8FYwR93zSXafwsJg3E86Rx3Vnc7LTntq0zyyk5QwtaO/vi
FHkedFFX+QnyJ8sRxl0b8vCMlIpBdfdt6yNkjaDRttgEsEk5g0V2q9c2YyogcXWpb+t/LOwSY1JT
gj856KNbVR8NZUpd8MZsXJMmP3lWIgSTVQOrBY0aCdATwX6wabuBfwUgP++e0oMzEEBDoXbyGkyc
28eiB9T+js3n3rxzYUCmoHpJiOU4eS3xQlM/HeFXRKqbCPMHKr9sukwxH9g9LQNi59FZbNCU6g7i
QQZ7XMNv5TvoTya86bLYQKE4+Y5q2qqhWzhEhq+lSLfYz6NRYDnfurd7WUfAYTdGdz75+S8JW1aJ
Sx6KW29zyiUjRPWQqSQgElt6B3T2uiuRL77AidhX3Jhpwo+cqZzZc09usCMIwwScP1F4zjJCvC4m
WaBe5i/vLcPiwi6gWLwjKJ8L+DqOk434eQ855RvDtPoLqiNQSQVeaqjV6QOJk/jDK8Em0SkvwE4C
KylCouTvptHZONyZjoHNhs6+CnHVow18T4tvPJMShtDP4kLuWm1d36pza6jLvNusEl6LgwSJe2q7
IPBdQfDK/pJahXknSus1N2uzExlKXJEQvfU59h0Do/pw3jWedOxlE36nGg7qHGpvTabE3BnGuFX4
rvFnRiUBUHMl9TbEiyvk1T1sLd5LqvvW8CrFwi+8z/jHg3jLj2vuXlOLAd/2MfC3CqxAlfpKeZMP
eNhTUtORTjWsbFHi1Mu4c7KkUBsLfQjAaOLNPMfsBqqaC6Ke1+qMMJ2l6Djuh7cXI9772wYDnPBR
tIJP15XURs0JyjKz318EDAqzL68b/MYo3bmvWS7OnS81PB+5M6XeAljJCc7G27lWaFnTRaW33aqG
TDnOk5x3jdwLbaozNShUUotxLsoihhQoAXjlriNRw00tsZzb1HbwO0CEEBE6coGeHAaSHmoaTncA
eUYwLf1kzzHv5FnU3bz91AzFULZoElrBACY8wZSuPF5J78zD7ZKFITm/Y7Y7NzInrfYjyv9E8r9M
GyZUASSN59oCSkt9xSIYdw0bdL6TzLmRMosknzXGWWPhSYTLdwhFGa2KLhx/wqC9zQiTCYepeArL
88Sk908Cq/E6HLV91JPCHgDs4Lkf0lJ+rNKJKLQJxAZB2UMmYFVQXGtKXYaMdmYYqr7KMIUZqLIO
K7DmAZ/k93nZO0bb6z9JVQzUDxAMJScwGUgufZCIxPDoUPBaQcP9GJLT0tMjzmqqHlAJpjDbbvze
ynM8ZCv9KF+nsEVEH5Gk5eUOXu+DKdK6AlPVNR4r/MbfYZ7AvUeiYN0Iuk2a70knQcEzW78OtQrJ
MUdKWBstFuFhoHc3ijT6zJLUqwdTPAyq7cEMvuvpOEXkNrvB00UsQVEufAPrLfNgHzLUrNEMiIEq
k06bU8FnYb40x7p2BEI8aGUpOOfbaH90IJ0VbswOiGGPBTbNyycHSMq29cWKbzjzh3OkxzEL5Z03
drSFTjeeEDYmJiS9xwaKvRMPrJCoMMYgaGgyHfW1Gx2Oywg9cXdQBD1sFc0WYd8A5zsKgzjw+QE7
zz37vWR+CUUzS0sHutuEJBIhXUc47So/6gknaLo5f0tfhLIyrjKvQuPpQZbyl/StnlGMvfP/JXlU
cpHv2Cj4F7BG6Qtew+TxjsmiaDMBAgYwcxzPv1PIxG5WE65H9H/itjVvPYiiROzUXmcVgz0iWlo0
l8pOZa7SE2gNxW44+4jX/c7VY1wmgDMV9goV0WW6s9dmRkErd70zvfDrVTrgILtOWCNp7sNrYkyr
jDdrsOXx3eiuvOc34skYJBurdM7xn2ryVCzl6t7RF91maHQNzdsiEEccWsZMVQ2MaMoxONAE2+eX
kAEPy/4X1v2YCBPFrAqJGscfz8gZvvATvyAHMOCM5G4j1M0YMRemZjHG1dArvMTaJ6EOb7KHzoMV
SaIR90h5Nw2HAKHv0LAoQTQHUSc73XUdWJLwsQ7bDwUYI9kUYaVIs9A0d+VZOBs6lX0huXD+HvKt
Wc9ipf+MeEpz1QmTM1vXeNO99fLNCsoYLXCEDmPoK94/bQ+0/fpfZVaCWdmYcY7QUVljlN6XKodY
FkmtHf8VcstuzrSq8o2744PfCKnMfbtDbosv8DjHmjnzwktiF8XA5h5SP7v8ktKuHMTQTEM/ESmZ
CvAMcHiMYMk3LNuxzPg2Iqpn0kvOyjnlO1BoV0bbwQwpq+bB8QH9Rb4XIGg+e1iyvfLtnEA5+Cct
ANEDAy7vCP6tQwdGMCDFiTCxi0jjuDXLSZZWo/A8p0mexzz9Eus8TU8XFU3DOcgeUG0yI4shP5uo
lcEiXoqN0BNhrzQeZxF04VXJr8QhmuWY65JQaq0bOO6EAhuTE192CvEITc57Ba4aZOAmBrUXI+oP
VDtzRurzYsTiSm+NjDX4Voei5irg+PSKfEOvGlyC2Y/fbHRxTyp789srWM08IOIY99ZzTXuNZFjr
qFU3+rngQhNlS93AzGQuREmeVGqqwo6YnRvxuzMqT+EHiGVo8OWiFxXdNWO5J28zSgjbL5yV/N7e
GxeEFT/rWdZIWT+kC7i2vpYTfUUeO2cCiuVGwAKg0ky4hvWbG8I1C/p32e/tWXLzpTqjH9ACtyvi
Y5oDbaZcElvEkV9ohuqqFeiAvQ/Y3VizdSJxRou3+qkelMiXPKnlS71BX4jGedr0pxTYigw/CH5Y
9QtgoB+P8SDJZJhFC98TzWdlgGoF2xrm71HNk4gniM+pa5ZYMP9PWgiw0i+fe59w/xlAZA18J1dq
z0FNBHq1CmL24DV9q8f4hcPXmI9RodngnW7L4N0hIFerUf3f3bLOaZILg0I1MIGCwv85g+e9OzTT
NQZKsRbQwV+jv6s1K1DdO4EdO5pYoCPydI4G1q/Mq/KVNeb7NWP8OFjBYIXgVDG/XNHE/QRzjsxM
MDMGK7vZxKvH9b4UixHsgs2ZBgfHtcZr8hO7SldOJqZQPDZGovngG+rxbgMkpsE7L73fZmHm8SFI
5Yw2zcl74FZvbC8uZgviIqVxHsGiJexS91qm2dxgf9V65UH3/H8hqi+PDYEcZL/5woG0thGR1TOa
e81V8g/CVEGvU2c4rUsOdW3eT1hd/+1qZnJYvEsnToWoxT4QoMEHAu/7FIedED0U7W/LAUXPcsFs
efqIiOA/Ext/Rs1L9orAkuV4uSrcfWMHlegidaSL+qek6QKO0LiMRCA+/spFEZ0iwz/4e9TDoTfR
BFdHybFqcrheA6dlH/U77CrEHyxlQhjSVVJan63TUnxQ0acAHqLXSavuJiqmO/c+VOOcOdCQd+kN
dw9mXgefkjQFYiVX6yD8AkOwELxqgUj3A3+orX+5n1m4Pj3nam1uPlOCWF6HUi1fom1LX7AVgpvA
3p7l+45gxzbmNb+1AwLQoJKs9hpTn4L0fh+IOdeHWUQbafGPOle/kzL4wyEMVzb4VpRKqV+9E1DS
LXX+du0RaKWMzCXYHoM6eEZeflvKfAs6rSJc3Y1Psh8OTTB3A6Pswbfaje+pa7mF/PhCevSlXGqW
4v8Y2d67IrQ43aGFR7pNgIIJ+1fPwDy/TE5MIiMnDtVuqfy78s1JMYSOdtPqZHJD46HjpdpmoWc0
72937AapL+ShdneJToAz1TKBKJI2YF4VLaTmlHarPGzRpjinwycqenSfllhZOIv63f+k6QIFnC7g
Z6sSAVS7RGzK0V7wJ5oNcwl9RTy0ipVMpbZ1MUzCI0b0/mhxj4e2Ib32bSukLyd0DPbTIyfuFYpd
ZiJHZKpvR6Y9Lmhcg87/11HNxu27+SNuCUDdyylG1H0u7rmxkmODu2fSy5bEJYPVQjVlOKeP2Jzc
X/mePf5/vD6UiP2GAVO+01asq98IevNOfcE+e/vSDT1z67iNVLj34lerH0tkz9ky4fw07F7Obb32
83RIoX+0Qc7L+nfNu8rM7mTnWY8OYB7AdPqr39OYUJxq/BBBXJalJfNCpbwrMSrwmX7zzrHSvwnH
G/hC7e/RxR2defSp2S6owIiZ3PaMlE6oN+jH9P6cR65ahD8jqhlWjmPgNg6DKQuY1oIF1cK9BYII
0oAKS6eCOU1HLurG9otPJ9Ub/iCy6f7mVNPRuh+XqhHw/6XhfXkV8vxu+ZMPJN+uKHCglvLfhfPC
BC3s2D/JTMQK6EpIXKY8yjMMaKPP4t1Zri1bybj+5NNIh3hMYxRo4KKORcYsz4fNz8LfOFpRUjKI
19+gehGU0H2xpxaqkufz1s4czTaoWZyeBo7XPsbmOFfrIyXGWnlf4TTDhBUT0OAeQSK6PWCZ5zD0
VlQPzDIXi26Zjm2V/BDHGBVoPnQo5FxuTLgQPTgKFO9lF2gp1cyuAQ42vv3Mqn6eRjrrxnOxHm3H
mnIh3x9dR/vxYqpicadiBWDzIPIVGyD/2TKHqH63wg92l0G1hQikqDlJvSoJ86hi2/et0IkEGfYg
RKn2hbm4RNjJC6zM7a/VbMGB53/OFRKYRYuUc+j0aJxC3RBnnphoZWi8zMyG5tJQ2PhticVKUn2P
8yU/Diszpk29/PHSLxBkpubPBchqVtEyHQjCqmQfCUeWoNEVD+kpm/yHwfRcQjdX4MMsMSNXtbo3
vrBvGDGp5m5vxX2XZtpUWYCx+KQjGrp0U6FRXmIvbl4fkdnDCzDVv6v52pi6dLtI68/IJOcnBO/x
xSwTnumTRA/YV/Q37joXOcBPEsqaW3aSqRPinydrbMx6/0hxeTh8hN+FlUpVP6Vm0kik5ODf9mC7
1nE7XIGmTD2lmxioVi8LGtT1ZejydRCLwRyHs8R4vnYCcpuLuuuAHFAr8NT8OkhEbF5Xk1XeKzhD
2NV1Of85Sz63yZdxqenHw1VrofdHWO2OIqBtICbPFIwpU7W6UV13FE3zl9P436S78yl4QFtqZKjT
7ei0mk1i/H9JrlGzLyt5+o3gwHhJuQh2vPquacYyZ5iGX9O4NEgzXsO3qTf8/D2npIXTvKlrorjV
+qEf4hGqluWRhN3NNZZP4y11DW/8qyd0FgUTHrOFxLAAzl9DlNkt4tzURmSD51Dz+e6cdp3hsunm
Ns9MSACoMCV4lK6JylYlUXuIifsjHJ00oESgBMfpmDfaWhCwlfPMOZey1ewvILU1VHShLTcdNhtX
tV40ht7lDMvCLCnCEOJrcUXZxGHLywAOqApLHW5f61AI1LS2HM/LpTIyR34Lhie6XVUSW8dBfp8p
FwUzFDEkJDT01lJLBPr5RChFGzmpwjnCXrvvvMc0AhbPK3+NVJpRdWhMCixmL7tngHEG6EOIdMEp
JEO/cHKb3w4DOCpKQzqT5NNvI0NXM34YIE8YmHfO0IjWg4GNshEfvvt0VAuqBesrgc0WxmcpVW4T
kLiZucvNY9DQmMKRMQoK4JrFDMeNH48iNfDgZSfbQ4zha21EP+amXZz6OnP/+Xgy2Ri2xONGGgja
j67j3/yp9kQ07JcnDCFgQMVjcYnaBtbPRJ0zqBW9WU3vsh9KbmCo6UCpM1bCjPwG2aDznwJwGI/R
vl14ncVasfJslPes0eqsbm0FGNeUC8qlR22WTCJnwYg+VNIug3KzwxmLZLhCqdpDL4/8G1jXMuqw
37mSVXf+c57oCoegNTBiS5IFq2QM+pkW08Y85lOmOsi+/gd4s4J95Mz+GsvAsRUgrVGYJqszOJYz
61LQG9+8sbV0JnOjHam2HSbi0o+2vh4r5Vna6kYHkpX7/da/cl5O07Tp+4ugQhSUWXpTonExfvss
+0lIR0HDALitXOgex21Fw3gfzfy55yERO1Ca+2tg5fc1q7yyTpqIF9T98jHJSX0xAB0VlvqS1yvK
DPvnztScSXK9juFVOabeKncVlXSWTzrUBPf5Feo7qY5Rik2gXXQN17wjL6d/B+4jr1jLi96xf4uj
v0A68S0XeEyLpD05x0g+2KpBUf7z7XqulLRFUQEUszdjf8+XbmJB6P6yvfcFIod1mYJjvpBc1uH+
oRiBPs1AQjlVP0abzwJNR0Zn1YtjjUob2mI3iu3NVfXYNAWxwDPzHN5OVplbZ7YqQxFmA2mRY/0x
ql/BOZdUCbLJbt2HhQ5VkR47OaAHxhOTRZ0eRTDLdkTiL8x1dF5rnNFJe5wcffQ4kt+l6EmoPaAj
vo6JwP+m7lpzVsM61cN3yPyychTKxe2TTiOj/GXoCHmuYzklWpAjYChBnhTueroGagfUlCGy43Gk
ZWnkG5ee3JJdNlt9rbYTzaoIcnKcLWuSc58tcYUQtbt6fxyWIR5IchH9NV81yWSIa6/PSSY6LKtz
5CSnLai//kzwW19AN1liolBlizBq2RWHGYWoSPXodhEUjRwjsPCkldtVYMv/pXu6y7HGX/6tkQnn
GcjcmTCrcsxsWcMQAnPF3eqk2Cw7OEl+dVhrenJg5x9Rgnbu58MhVhWdr9JEr1BUyPDSwIF/xQfT
HXk9Hsput/c/+Mj9vWnv2hF2GFrUZsFDLVSlWN7Te7Qt2KA/C36jZCF35jAdFDuW8Gv3UiY/zOCU
C4DGYZqPWN0YnwV2AxbGo8qJXCR53iUMuoIRs8AHRGHE8qeQt3Nwr6BOcYYt07qTWX8BRfE02KHN
eSvT4r5jZH8bd5CErvEQIdRwAQs1OW8RoJjNnxG9xmGNo8ksR5eUCCIJbu5E6UaQ8HVFSW4TLpG7
Mwevjiwp9C3HeEiO+11BEYXxPJ/ntsORXFoyUk01z5LEOtc1tMmZvpTb2iu3gavAy47GDESyT0wP
3birUj3/PGqfNZRGOzmN9btSeccMtdJRp5gKtTEqTBnD+UDpRUjhL2Esx5WItid3QRQNWNH2nuZl
4IroH0YUkbDa2XUtbjlSu9byDeU6+Pb8/5wYLAaudwTIeROxTdp79jtB2Kga521A7qoUQ5AgVbuP
YbbCE/FIwSfxzMRclt6L/ZgFPJ+SWaGEIGu9yV6Xh00ND5Q8O8aSS6s/8UZO+aG2MiAxzsxvXqrK
vqhTmjW8dLg3twVKE0Tz3s3NWiI/eem1CI+rmWB+numzcY53tSl/WNNI1ridylAVm8qWp/03rMun
0b5vX3XVD6P30RrpeFyk9tfWKjjyFdXsULKBzkZwX8h9EZj+kzvijFNZL4Gc+rlEFJ9iRRW4pZ4Y
dLH6aXEN2MQ1Hk9Q6wuQ3Pdu96zP94PcSGO2r6jx9OJ/4A4ElpwHBryNdClFKiUm2q8zmrPyyagD
7Cf/fXkgzpGvNG/wCwb+w/SWYijPvFaoewTtIK5yzgeuGcFOd40++P5hrGUoP1Ep4+ixK7A0Losj
3jAbi+mMxurVGgWj4DGsuJ4lP6CAXxJ/11z4h2RS2nx+nVTmOvFWx+02rmjxmSi4OTTVgtqg+AVG
A4TK+ZGNFRRpmJo3cXd09CWhvbdSeLACRJ5r8KRlvHlcIG9pRaXPVZcxZOyLor2FNnFK+EgbEt15
+K+xkcR1SDeNxPuwSHNw7Hp6L6Z9ihh8pRL3tJ9Ka22nIoz+jEwmPi4O/bwlgtZHciBktYSKREvL
dK0sn+loJ7SFUYqFpiEITDr4/EXH6uC4Vuq0jlOkzDcKX2dgkrbZAqjhPHf026v77Bab/a7Exp1G
6D3/S6JE0l369h9t2YnUMUEt/QH2CCuL5QUGntOXAl/PSj616ZX4xcpihKHcBo2hxjSbMXtm54le
fO5kbVU5Z17slgo6/jaftSx1Ju/HWtjATCBS+GOfdqei7QbZ5ly7P3kS17TKguUl6K+87zypbdCJ
aGIjDGCEHL+YYMsKsq+rn+kTZaj1UsUrzyB2KLXM0JhlNOA61YYeM1e1SOz90UFO5QoZOtp2107U
V/SNb1qtAP/oYSQmMAysmOwr/N61VO0bQ3V1pWssKvygdm2pNNp2ssRPg6uMApwgVtwk8jiTpAcE
L5b+R0bbvGqttZVhGzRLP+K3GQ02hAxhL+wgAc7CmHjnIoxD1V3o8A8ywpiUXswhLEqUdO2Pkn8X
y1RMUsd+IzbjmNbB7F7kg5dF+QcgaP6xor2aBZcUcyO3GWcLRGZzAcF/12sJEovm52O0RCC+IUkN
9mTbyszZDP+41acCVrA3Mz3M1fuxLQfzZlZzf0WxWnWZyRwtT+5thy1JSYkfdwU2Y8999Db/+8RR
HxanbXEmXael/Dsi20OPzXPN0KTPz/DNjsl7/5Dmy/iS+QQ9OxMedmJzXoo6vcan9bbYxhYlHBW1
8wQjKcKKQYR14DbUHE7Tv+VTfb2CCr+yEWC2PfBcdGuVud2TcnMxkNwQzg0/TWp6B18R4jturfBf
Q74kD0rYzMFa2O+U7EsKK0LIAo4JM1SHmJHieFGxS/PktjQ01X+q0OYX1m2kInNES/TB5ZsdtiBO
QoDHXcy9RG9LJC1goGoZcIlPaXTpr6SH0L6RUX1Vd/jBSOfWRS/aPA6ReEmqA02BYlovJeD4oJJB
uW3t7ZXFvZSOXIg/Wse60RpPKBf2ahapLRj6HbV+b5BCsgJyNtmnjLj06wr7YjW/43HVk6gHe3J2
DNwuRFLzlc/snk2a2bhQqs17B+QUJLLht15CRUy24Im1Aekp0M1llaYj1BfhVr+jnMThzyCzTzJS
YR3SBG06VaxoCYHltotzYVXlh6SqAIkVvYoq5Qm1bTVN+UQjvSXdhFkzHhKuD04Iv2U+ZYqPw3+7
vdoNQkiulTIJONNf+13t1IrwW1qYq5qPp2yI7Q/jcLd8FV4QXgIzYx0BpfwXVGom77n1Omx3GedM
AmqlQUteciiiMMBvY1rrn8rMKmQCWutpXCTc0q7JgpgIla39yUohBqc8vUf050OPktQVir4ympeA
LWozmdou609G85YDIH3sHOjD9HglwGB+R0tKyysgtQTpb8WQ7NVyUv9ftTa82UU5zvHax9K9Ye9x
JZI5q4+LhmhPwHkWLWYVCMOnPsJpsEh8hm68wJqdbqNgXFuxJekR9h25EReUT1yHKBZzgzanG+UH
h1lZ248d7/V6ykJNkrpRKRzJqjYSjmQAlIBPthj2TGm168On2npWOR1npGrSk0oguDTAgS0+Hz7n
jmJb8wjd/uw1u36K8yqL4WKZ55VlM7amc8+Z1/fL4uNNt3Li+zeEb50WMj5J3HGLPkBFGklERMyu
3+vF2nH7F451xijZ4zoeT0rjm5/rHqYMBojruat+TRRRgyEOcp+W9WmbuOhG+U/B0XQvJPdiqOc9
xwVSFgjkt3+6NGmMS4GARlhBVzg5kkZG2DFpWRfo6oG4+BYNs/gYK/aZTvaSaSf0+qhpkzs+h9Hg
q409MCTiLH2PxOIfkTZ9w2iSSrL6afW8y9faad+x7Q5zaqjAsdt7zCYq72zaTiOy/O9S+G4oN0R5
xkzgjgHV6Nhaca1LXzX3HHpa+UtNtTR1TmJbDTLdfoI1A+PuP0lZf9FjyRWS6odASM9QF1GwglnG
0HdHHueIgWIz/i/m6fds8aiD9b2BJnGadL6I8t30pxk87gFhaZw9bXAr6JR3ttFOXvMhlxuFvsGK
S1Clc6Uc10lH2MqJkNYWimhiEjCDXc9zwBtPpTttglQKhzH0AFYjM1PqlFpQ0pZ5UW9abke+Gwtr
NoZH2L143pM8hE6iDpbLEralvc8D978j55x1GDzDoYB3OSHrYFszWgDvqPEQi4vk0ry0F5FT3W1o
QJIjShZ3/lB3C6mlzt3/0IatfhbLUXQhkcRTjNAyvDnoCGyzlMbTtIuL4W6/khtM8mHxXTUOpWic
HgN7eTaobqdMqzfe5sIjKeOfJ7y+qHxPZ3JRmwfLrvdk5qOymmht7xIwxElc+w1mXW7G6qukNL/R
uDoSYuSMmocExb123mAkNkjSGo3K9Mf2DfsGJN2HNqwQCXTZlQRklegogOX4PYjCivd5Ffrgka9t
gUszAihtqiROPICpQ9U3EIT0FCq+04dGRPl1OFWpyLeUwix5EDyAyNQWgtbEDkAdlKu49MeSiaJy
mPA6HXYCZf//IcKDD1hDs/16fYZzwLg7r1F8cXoU14KmWcp7cn7IDbHZFbTXlZKJEtygxFLcNgIf
/bBmNzbP2nMCElqUngziJU4xMP6TNvbTwSUXjmtnOzUlwrqyTAZGcptCHMWq2CW/HbdUGfX6WLcN
cK/0qPH6D0HlBzBoG3OogHsORiBTO3AHSQXYIsZBsUOADYZEZFeuhjuY5Qr1LjePxvGAa/pAfxMQ
Z3IfVJifZOXgy71pmrkjh1Qo1V05wIQMnY9ebmgH9IB0wWbikWu5a8EgPlswhmqvoP47khyfECS8
lqbZABdHV6qKX/Jc2gFLTpT7vSdpNo4xHqRjDgIdHkJub5rzI/I0tafD6Fu+YyNCLwamGhEamE0l
esE6CQnAHqGVO8sjpP6stuN8roRQKiQny4Owlvs2pkfzKJa91EPMZkFKPz+78zXZ7W083gKppT1r
J0IunyC4gL6T/J1OfTUOjSymRUdKKmO9xrg+OeMfKmTje4s5rawLWIYFwsTwBi5UH/DwDFGsfrTV
7UX96Udt9BlTp8Kw8LvTgxhWTdcMEIMdfF3LT+F4jGG5+/xXX/Kf22W8aWg1QVhwem4md78Yiekw
67XHGYV2VMXzTLWoN1HKe6uZAZI1+AY7r+M2KynJ7UZE/ONu3+OtHLzbsyao92vY9Gw2NSnsZ+ml
QCknj1Z6p7Grk2QLdm709K+wDFrZAxW5L0s4PtIalenyv7VZ8nonwbEVj0f+2A5f8H0tGvP9qHTh
TIuMbZfPA8mTkDvDwjWSlAqU4ZxmKGovfn6lwqbyrK4aYwfJ//MFsmWi9HcIA+FwVxyy+EEzG0/C
M867zxrhHQntmwgJG1QgaMHgyU2FVhBo6WOYqRnrK2PeJKcosNi25AY41LsIZap6gLf43X5WvMtd
jLyh7n9C+bf3BxEN9KssdS2/cghzLVEKcBfzfzCqzgqOF7P8lDERgqL4EKFb3KKsC4Y6PxP845cO
PBiGVMVhC5ZMP3aafhiOYVM7nTSl3FCCWeijPTjEfnQ9U+XTfD0nmFW11A+AndGSS7Yj6lvChY2L
W+QCDgbzDw0/VMzDDkVooIPaDAFJ+FAfNRyo6DUlrQ33MNyR5NvsF+2boUMRYFTqFYD6fJTnaYVT
JKJ3IlOeuzDjdzp+voYOXMQ6VJAgSXM4M6IYDsz6i5SxkiYqc7cCutYoma5fK5GfCfxW3LbEI590
kqoMjuuA8XFs2G4EMiyvEXBTbxnQcmsGuAFc95iBznfUGambFu3oVLoxv69iTUUg/Y2mhLDg+cRi
2LGPg83Y4vML8LXazl+q8Zc2dBGVIJletLv51+tRsZlNtCz1q7YJqJXwbKJd+InHKadcWzAQXmGD
ceep8H8Ay6sWgyWlcIVHQztD4XN7a0tVKfC23dLFxSMjoZOKfZDbCsP31Rj26+bRhDiCr/LGJ4TE
Ti/so965kM9OHceGfvaOnYyqGZYdHv/A7PAQ4WpULAzFq5OkpKJNjMwPPlZjneKdbFkc0VPUPoFV
3JpxkXZ3f0TbbM1PehvrIGlr01SgWo6wX6Z8aPhRxZiohfjum+EN6kutQLubnpxcpf8zmlLr13dD
wHpFINkSrsnTawJfUQBmnaba/6+K17cpOL1kKI6KaxUWI1+w8cv0l3mecX706plFOiDntBN2A5f6
38yWj/NpZXPiA3rR6JJS9vSqrU7Jyo0wTU4+/WCs14Z9VKuMFLddL7gVNPNBmcr5n+H7RUCa+AJc
NQEfMGI7BBWvcpTzROjXlWh0nIRrpu2mIPZyV5vJ9ZE8nss7KHsaHEFsd2NSZJreRNs9Ap+bCKaw
S6srL0HyNpdEuzpjlVMxL1QyjqHLFMGew9+XTec465yB3WvY0GMbIdnDo7y/U15Dw4DmiGZmie0V
GM2LoXLm77yjW1HucB0TIYo0w1Oq218SgN5nStquxf6eJZvabv4lcad8y8Y7SJ0HkQY6hnf0yS4T
Msq4SKkxIuoOZWryJ6gqW7nnO1+w6DVmzyuKGSRJFWDDTcf3VWi+ATu3YN5Z8gk+ENIbMf4QWTz2
rCSG2+zdnpzmySPynsqtL0KucNHxaDVU+ZkQsE/VSkY60w9GfLvyKF6afTakc1LwsMt2fTCRIftk
BTyWdR2I9eqPMDW+ktETn97O8bqelQIcuf7wI89e3jbIqb1SKcm2RQlaN72lMTntfjV0gKo7L2Ri
Rfg933YNNZOkSaqvgIX/GHz07Sj5ST1f7GHf/IxPC36/ablxXGCBoANc4OXhC0EHasJ7A8+onJiJ
R6d7R8txWYl3rvUeV/o8AFID7mH4ENwf6H2XJhos19blhjptX3wA36Ma+mY7uby3WX0Ug7YciiaM
Ezkzt5nRHyRuDoTzIbuEjLl0q5BvRslnQtwNGUtbwQ5wDAx967angF0gPUzy5lFCy0DtiyGGy7Aj
z7Sv7Okd0sJ+z+jsQGcJjCxROe4kGItoP6dVneLj7soHUZaPl2xCZGPF4D4KdYUgu3qLxioljCcD
9d8EYM2QhXx2nnaitVDKVFUx48QBkZUq1j0MiZBNdIKvisXdJXcz07L5CczsZX4RlSYiVfnGbxzg
4ecPJZZsjzBygLjo1ZQBRcvHZ7W4tNVbwrNeQe2uDwdrPqzkg4ssKMwFXpL7TvTeOd4Ss62QFFoe
sSPRJ7G4BwZdxfCoADk6Bbe59J4bokUCRFJtf47v3WQWM3gHVU6wY/lkMLs33eqoy36HxRxKU5/b
JkTcH+wkv+TuqBnw2MlfZfb6dYhChYHy5lAU7JJFkDYINBUqdoh7GK44+vq0wpJ9LxjRNCbuFr3f
4UXOlHHQO5HQyYsj52XW6ZpV/Ncfy9xbd+3880lklBtXhb1yziryIZ9WyHvs6pxCsavZsTJkeYG1
wKaQH9737R9HfRdIO0GhjkBGvACnD9AWfLFKokwalQ63cBKzZy/Fc1h6+K4AzaeGN/5OPC8pfJGm
3FlFNxYxV+JDrjF/wqGNF4Jdm2ww4UKSV56LMFtOOyzJ48EcDWUiCt0VLsztyfwHZJVgzijYvY1V
8LdH/glxyIirIb5WvCdi0YrdmhaqMxaqIIyQ7NbDnIHamnKFT6XR/6Am2Bf8bZJHZjv0ABisMHZx
E59vbPLmhVqt9ALfJtkVYWfgimJXQKSDikHCPmakEHvspSWKzqpk4jLt20Lo6DUtZudyeBxzl4mr
NuWxVrJXa2kqazm8PAQDrAOBL/wOXW6vDXJK7wYovB+ED1kNIxyqpRyPQkVrJ72+8AaQYadh6Q+V
P+cfg5Qq5HMP1Ov+TbSTQ/jZLXmiQikHu0nKX0Cq7o8TOfjCYxIJHHeST/hxOKPFdlhOMDMK88TO
/QJ+h+bQRXPvHU3Gb1nJ/yagPilpx8YPbgn4U23axo1NVIigubk+Jxn+0DZVH43Cs19jr33Ek0F9
7Lv+sOY5etMs+ASemZMDEI03lqKA9X22XpS7abGOOtu9G/mDSwP48A0bQnDFA+2J/J3i+1GbCy55
ybnMrW0vwHeGCfNTwMf5VTe/BP2604Zs3XwM/n4vyJG1BtFMnna5nM/6rJCY/AKG5nkiWM2v0saV
MUvOzcSjzG6gp3/DA1VmXG95fIFBsefzkACzO1dSi3tZEz9j/GgdzfrlicgTybhrXeTtod7/5Oej
WI9imSgXTgI36R5jc0jMwTJDHkIr8ua8qn3JbuZIBOr9cNpnYNEUcZX2kloJ2OYslwQANuYd0xdY
x5PDpwFbqXS4qkYUc2qwTLtHlzKb6OBBZy9QBGXMNFnkfd39MT5QhcxGbY5P3emFaZevTOuGX9YH
kMdg0sm0i+ugOHZf0P9Hni49mT5CFQs7FeaJZYnNSRju3wwK1VRkO1cFbHfKdwtU3voT6amMWz0W
PjkYbjLb5vOIC5JeAjqXGQXoNab610a5R6aq7J8yOpoFOCucBNGAZ/0oLVTS2eFvytFV3u41cvNc
ufKKMfNtYAVANkSIdCts+ZQHu5ORtlQb9pXCWERT3LrUFEgHgqMuKckB1t2d2Vmz9wBI/GLMUQjy
5FMNlfHSqZRgf06YedQLy8EhECfPzY0jlHp6eaCyaQpjhASPYqjOKU8D+q11XUBq8uo61J6q6uD9
3L+U8CRPZvCUB2nhE+kZZoLoi+5AN+oQvARC9p3U1PWBWpyCS6kL+PEAelZmG88GN17LFAhMlZgl
bqQELrMkrJvyjmvcfjB7OZ6qAUYoLr6FggfyTY52vPO+RbEFI79mqmTF2LiB1LJ8V8QKzzi8x7Yf
UyoXifKGjiE87tsdDy93QuSKtO1Zzfu5LSiqQr8R2yKnjc9NId8yQr7hq757DF1ylwDU/XVgsrdm
yXifMFU7vAy+yXoG1Ed6c4gXhx2yF0p4MKOm1P/S8090XErZlTRYiYcuDpSIN/9FmjgRZQ55Dzw4
Yfj346Ia64chjst4lGonDTY+UxWGJMjwMw+YCu//Npy8D8eEN1fiFdK17YoRSiNSX4iUZyXtkJjS
ysKa6ZPPBeGV1m0GZURvRo46IAPU1ffcI1dwfqw7WpGYo5x72A4/otygEfRPzHMNdq03gkteyuRF
O3rNNnbkol3pdj7ESoh6O5xu0egFR4jU2w42VwpbwCsglwGgL0glq1ATsiHqAm7v6uJfLUsQcFm7
hxNRFYB0zxyNS4DDIAxxhibXVsKqV2WB0m52dpKIp2E5WicBCjBqhor0XYLcCzL0g3IX37D+1rzH
s7sQFAY0A+AUj5DFWMRLtxSnZe63kF6PDn4xjvM0u4xI2ey90erKVH6cc2I1WHTQCPfl/rlGlTmj
XLil7EC9JDAYm3c7hzdrR5ZRFdrFkt4B3oSE+7hN6KS4s/p8ER4arQ3uTEwCdqDsj3ueUjdXplSF
r6VnJc2oXlRfGetsGO+raAdqgK2GOQCch20NRgZcLF8E0DnYD6dsWZFp6lzlguvIVMv4wUOshNPT
FsOeeeOyBiu4lJuplI7P2MKxC+Sj8s5FJiA+IENvWdz6qed8NEbwqfrF99xA5iqmlZLJWaU9L7Ze
gTu8yDixsEqEDSEdXHkWteCEyqUmejG4pEjrDyRgWAiYeVpgi0XirUv63b+tjjAWHLUfbD/v04dw
t4Vt36DOHZM+TbpIBfXRKzd02/tRk+mU2Mcxva5y928UxhxblRjeXFxsT99nysrQYgO5w3o7NNe+
KMeoMK1IzsK6exBIU4oR/kj3hyph6CpzTIy3iwNuA7fUSiyZ+f//kZvcD07wFPcTaBlw/53u+Bi4
UvpyPuZ2MbMBvfx3o+E+nz6OhvzG4XgAmFxtDQT9bCONWwbqk4gtEuoKKLw8El4dYxmLBk3C2ZAP
2rHk/Ftrry4HiqFXe5FvzJR2/GBXanFpKcygPp8JhoxYf3Plj3lW7BHi/w5YwZvoARXnYu/TTc3b
kYA24R0duGoK5kHLsnGY67A/Z2VobI7+nlvoQErKPKGJpTE3PnutgJLTKEW1ZH4m9TqnrWv+AloC
A0yqC8bFTr234Ez1WUE3Ze2y60yAkpWSw8mS3oUry+AlkJH2LWEokX/DjVzCpHKPXAyav+KZVqce
7deUOnoPx4BiKaI3N5dKLZJlnm4HlhiTZKEwd2HUnN3EHLPL0NUEf3ivsD0e5SkUVy8BfM8Ogi/w
BcbYsSAI85X2zYSgPZOBnq4rWvQ+kIypQgd3A5aS6ks/mNJkIdRbcuaRXXJSQvsF+Kt3aO/IM2/e
nInsfDGxFFGRwEAMvYmi2+3Mey1m9Dq/nikYhy2cNufrdS7n9RBeIxS1cbCdB1CrK2DCF91neOdw
cmNtTQvsgs80j4atekF2LBOMvizCe5EvzJkTi8OBFwsXH+qVMXZV5kRqimNwcURjLXNIQoKWiJQM
vA8PtJAlDTx0tbL86a29VFqbNNgfMh93TKqHQaCv7wlMpOfBi/lr7zOrpEcAde6fktvU51wvhepD
uAUXuhBmMMM0Z5ffmlS3rrRqsPduNDd3WukamzbpEs9vxQo+9WlLheFgFKjVwKExUPn1o1p/pVCM
9VcjNyBFRPpRS/gkB2Tl/GXJzUsxXfmohrwX8Nf9RW2TGZd0W/vLrcg//4Saf2UFs+wKj5t2Knqi
lIbydgCBJSvi9kbn4bNqn5KfO15av9lZj28D4gAEVvb1qmDZ9p6BeKBj1W4+f6UbAqUqipNG84mR
uVDmy4aHBOmXMlExbsk8h/jm2Y+qYyiQGqTsZK6aydBeTX2l/BC0vmChKOMu9Oo1MeHJ5HjRlwms
QYCE3ZYz5ZwEv/2SqXVQgAmncr/MtZh93lyO7+j2TWz4dWq5vDSDSHQiKn5/WovqZmMjT4WbNx9y
y6pIQq+GjtIaneDnuShjXr08Sz5yufhz6Kt8DXMuR1hk2UWEe/Ze9m5dZ33JTZHPvG2girZ/LOHI
4nhI/Q7ES1pWsjgc345TBZAxRs9lwH7U5TGKkCkeEuC5y82mCra24Sz9p0NLFLr9emQzFsSUl5bc
T6PsB9itWjFZtBTnZ0vBEFomrn7b5tNh6HYalPYHo/Y+eJS3v+aXX5lqnalv9Xw6fwBIpNewu4yQ
jiUMJgkqIONUtW8eL53cjb1yb1ybUaKs/9kkJkwqA9CfQi0Ox8d83bWrCDLjvRgwJYkwnI5c3QOm
+3Yrk9urGbyQMFYvbferR5KFhAwGLRzRSCrI4igR3xGSRteHpv6KGvURCtSRRK2y+jaCZWA9LriC
MTeFJOjtk3KnhfCXHnaCdAW5gMUTVFRslRjBc8pApbK8hIDZ3y8+Fs3NQ4ckk9GPumardxYPKSRF
oEa0HaKd6wibFQnGbfIXsEkCVenrBDoQ63BxOFrsMbpYxJUD0o4tq00Wk5mzaadL/bBzNDQlNLG3
mRaewTUG+po6j78cLLePmP5/WCS+DBogtZuLpzdnx4MsxHHjvgeTdhuGBg4ptsUWwuz6rFjGzQue
sTGaC9RaQ+likLc1EVbU2Nkjo2S8T0PugUcbGm2vUFz7OCWVnCGpVvThrkVg7X4wWHQkzennenAN
BT269kt8fntMSoTt7scjUyvsxQeuRcQ32jbfsnX3csYUEWVXP9IrxmW7yhseBYqbVAgXEreeC12B
TkzTkxWWedCE5GKj7jCPaiZDIk6scbtuKl6tEqJsKSiANIiSwQGnzRicFBLJN5a4mwLijVfffkBm
w9eCFmhlOGsDZ1F9DFBgzX4oraa375BAa7GrZNdQhPqb874nGQ9TQ5zren0zhNZ2fToy/CQBTZMP
/HhvHkwH7MQw5/X8SRIt0oSA5R7qO2Ct4aCFTjPNCDXfONTtbSEc1cXRBZNmc5xKXlXeFSORoHrl
8BZykIOisinLLJhYR6fDTd+BR5TPbASRuv8veJGVgqlcNmoQc5H1TNhoThzOzMVMsjtIfHzgRzZf
K9HfFh5Pk3WiUezWbv61JOx46QpHCxXT/VHKzUygXuJFMNQ7NFE05W0j2HiB25OIiSGriqVzzQT7
KP6alHGHhzqC9XK0AV42H517wY7UssDYLilqbf5cmM61CoqnqSS/pEvXpndHxK/RS9PD+XGCVgIv
+mia8w4Oa2XdyIOwHlJ9aMGKs5Q65SnwomNs2Ark1LPd8DohBkT5Me55go3y7MKj0Y5cBsFBI2mf
/i/sHawy4/ISb17IyaQLk34gNFkAD7zQmDxBl/8sDHYV4vvz2mab+BYlp26RyQj/ndMwtE/3XLhT
NVnzZduVTlMdJ0vI//v7GaF5Kn0MxVzo7QjKVTLWGX1HxnVhXH2xcdTmjHX+LeuB+tLwiMiYO7KA
3f29TgyfaSrWFHvKOc822BqWVGRG7Zq1C/mYRDgEVorYjtSAjfkA6WMI5omm+2G4xGOSVr+4Jhl4
yO1Os+QqXrNto2meEe6CHVUzmGQSN6r2FD3oBqL2IWEHsNvSi8U2j2T/2KXxj/Ix9QiMkJA4DeCC
jQpbpuSfTU79rXqWFH7Ehqz9M0LkHXqcjH5kn6HSNF4J/p5J3dYGExcSoz6tjynnDPcnCYysOn7d
ev1ILo2BHQ2zNMBpHI7dmZ19oxGW3OFiENblQTDzWtQCpzXIoIEhhXp+mQ0ArJlest9o8fgp9Xiz
+baAzBCx4/WBdtBWszYh+l9BaAfscaDoGpzwvpUMbIklL1TQOzAIJpijG3Y4EmZea7riyuL62a2Q
Oar4wCGsmMQ2hUKrHVCPQVxGfv2MKvO1gJ6xErp6xBnxxpBdAUnOlmS61GohDuEuw4tY4et10qlL
gkWbplMA6rrLD8lCB3/5wyh1PkagzYrVP/3J2ksonvObkln/VtJh94hPfW8uTzW4FJVA/lxNBACt
b+7ff6lGaKOaph5IjeYB3x6DM4OiEY3aSaa/WISLIKeGCJh+0sror9H++9bATxq2IcjrrxeeJqIG
SMUbluYkDRuyGz1rPaMxsyXVk9Pz+rG14ZYGUwYdtyRomosIhEHpTiwwDtkUDqv5aqJHifVGKo0P
dLT5P6c+mH8ftjLu/0CnCAVEqKjCT9oodeDrhFDZnETVbXAhyXWXQZhGTN4AL8PCFc154jIYUynm
ZKAgBeQP4e5Um3vC8nhk1672/kZ5uN85MXxZP8vOuzZLRwjkJZ5/eeocDcFT0QWWLQ3P64c4ouRK
YoCHRseDBXkI5p+aanANFVd7P/S8QtR2YZPmYnlx9Fqc6ejfM5RkUo3rRXb2BINaDIelr8vXAUWs
NTch2mbbGgsfDnEfozyPpl+qZ805NBYC/zM6bdzbYjr4kAGEQwnyZOzPIiSEUuVzCmjd+uiPySPw
LN0USmr0vnMNY44ES6iNOQiIG3dDrAuwoy4nuSJCytw5nkISi24fzR6mLO7ysAwaxAFfIXGdvA1d
sXDzlzSle79d0STzooBEwhddT5b/OXirvdwLfdeGv9skHpAhTVisO0kkLiUAdKOivROF6nZsgBlJ
x2yc5qQWOAczckJRm8Ln7eXGMbpF/kgDgXgsRMj5FMoyMwhCIkLnXSh56JnhjRyxBSlccDiryDdZ
5EghaBNTiki/PDHX5q2eZiWcvQo8SwLTGj00A2zgLXT6/kmO06Lwtfz7JwINKsvC8NFs890HfvGf
lKDJv3LQqWkisJiTuX81YqrYOiI0i17sE6pNzFtcH8nqWtEgovxlckuJcqZl/hisoGTOgGxmvSF+
pPQ8F1S42bYGdAGZQqcywh36WN1cD5ddOxCXoFty9HD+xQx0d90+7LlTZDHvURdYDV1BNLGkdlty
WUDrdP7lnQmQvvSfSLlxj2rFlvNMdv+xW+WZFfZZ5l3UxQk89y2pfKhoYQYvPA7CoV+BL0fqJ/BI
5fdhfTGcKUGikScm2brC6niaDx41vKEYBi9iZIFgv5XfDmN+qW8JszqvrhobXbS42TZiRTEil5PH
Snpbm3Zw/63nW9mU35TqDLCq5wO+yeQx4ndclum+0kS3AwVCr+mUAHN/C6yUR0rt/+DSPWH2JMxQ
R3NV+29aRfEmWxO6lLpyuWg82cD9QETzlZ3AnfplZyzl92/P3i7StUjzemmYkgx3j45oSB3Bk3qE
KhzOc6nNdRC5Abm6wMlAar4ciXZVbzHao7bL6JnGbCbCRvx4+6Elm5aaZq8fhI8VyUNp8myD3R5X
BIbF52koEuPGgnzxn2Lk5rsEtix+d81mY2QUhwar4ZSVClEevcdznZiy55dai2EHDKT9wRs+uEWY
aqHKbKog0bXZA0LxpnAXqir33I3MF5VHNl8rT2yvJJNNK+B6ymMfUHartWjbnmOBSxYzvp56zuBu
+M3pKRMYhDAfGoBftM6sd3fvfTXkop4T+hwqjaUkesDaSptc6FjA0Jpfb/F6l00QZXwKdP0neoGw
EB8tJvfvm2Qrz6yq49M1a9wt0FYmy0Xs4pWlKNJAO9LUkGVr7pvfpuRhS5fZ/wDmqd3DmVzrD+5W
mTqZTFi8CON4lzXxoOa3EIykcYL8U8Bz9XvwB5XEQVjzG+teOaHnhoA4H0TQP8Mw0ajmqy+yvcqz
p/Xmh52vTLMUEFHuj21mPo5KRUzohUatasDol7L+NNICElhkbJRmSkuE4rP7tP9/Lr63qNU4LQ4L
0y7pqc3VurtxHWFcsKPEmCtJWvgsQ1DxoMFGhHGHsA+fRMTKnZ6JTEeG2Hh1/7jKtD8LPsCyNrjN
RDKRasdf022FpLknlm+51lrFOfZal4fHQogJvaxcMl+vKYB7AkBKALO2Ocplu1WPGyFyUxUSxcW5
PCTOr8ZPFd1qlAI+WVGELiJcgpPRQz9JMPrtO7WV9c1FTQDghpMfsI/VExQ1red3vfCddGkfF+NH
MCkxbiADh1NgAuQ4Q36AXend8sftRyW4AmrZFRtrQG3jEBtL6umnEDn92Up59NLgU+B4JRSLsC9y
TbnKFzzvBH+zyQaUTyS7VTLmb++zBbwqvPEO+tN2h2KSs/Oz7Y30lXS7yjWDt62JNQBjdbba7i0z
/zTNB3QEKBFi5IsTp27urAoZD4Z6W+//nPoMxcG1xnkkqjK8X7nlQgv8G1gW4ilfsiQp7palQlJ+
NMRxf51PpEByxqy5fyx2oqh/3USC63lFBXCHHqBJm+cCdUr72QoERK60PYw7LUonLfGCb8j8k95g
smswh0AwtZm8Aq1/KW05DpC0HSGdSYesCrBrHN6EKqzVMBWtUHcchyOLs/Y/4BPMFmh9DG4RayFf
Ln5xp+fEB6gHikeMzS5FBGmJo0qR3twm8amdH0CaTteB1q20G+iz79VPp0+OgL53meabszAyUfS4
vHMp+8P0doCWwcRYKtPvNvV9BuNETaLGrg/K7YHSOGJ7Swm3qGp6HYm2BHvIY2/0q4Vdke9iWXHw
wgD1liE0G9FPdYKYq53OPPXRumzZREkjNfxG0+7q9SSVyTioNIRHBIroc4kiYgM1/wXfCfq9n5KP
3ec2C5WYBhuW0P0IdfDAo6pbkQqCkKTigCIEMQiMCz6y7MOT0hGzgudHReqf+ahHlBQNeUezHloA
p5ARUOQJ/sEPNJShlX7tekUjndQfrtY/20gUHu0JsYNNWQrP9mNaeueBpOpyfnMOQC9L0JQP+k0s
7K4x9+CKiutbHWw3TwLqkwo1Fn8U3YB4LVyB84LwWVZB4oqqUWCXUs8cz+B3fXph6MIJ4kb/9bwj
b6mzj/MP89qK0VOKv6QYaOiIbvxYr/mlXKnv1PoOS+BGcPE1QclzZYD0cCVEZukWWqGZ8avskIfj
wFmC4PLWL95QwCWRYljZuYr8Dx308Pl/Fd2zJnSl7DQczDyVleB+F/scJFBvdVHcRPIq7AiDwJWs
N7B3GPYSw90YPbB+RueE7ULn7SpxTj/iRjIUNKuXMo5+0giYBk7nJri6Wz9YKrleNtgvV0QCKaVM
r7KBAOmubpx/Gonn/aEr5Hj2QbRBirUFny+66EVzzQHG5HGjsJVWk4VsNUDBqk8vTChK+AIvuvU0
igm9pckC8EkIEoRifUrbdY4VvNyW3gsVJqOndtK9XIjeYGG+Ok/TY8fYQPzbWqQ2McmoHf6xxwwY
mT+jMkGiP2cYVKkxrR9cEeR2DKIbeEGad1hwdfa/Vc9SzAvBmgumOWbAUualGnL1hhR/zXN68g5p
yDp8rmafNYDJ9o1iAfoIJIKxiN98yawOVb/0KkhiCwxjnpx2PG2FeEF0ER9WKFYpB5JVpw/b3B26
t8Tp3vS5x/Ek37/hKuyxlDe8j1IaCxNVH+LLVOhQJJnqK45NztYUWhwkejIISwUjIJN/0kOw34up
PO33KG08fzLhxl4y2mSsFuB+SUp8B2chsnRQk3kkhRWwXI3gCZpnPgv5buqqzopUD0iSgjcX5SfD
NlenhBN/U5qQNIeqLQYn3WjdsILaL2jBpgidNNJ7NJvLe9ui8vosTA5LWzjstvIhoE0a0rKaX1EC
YZlEqp1aVdEk9d9AdD5sNiSG91YjMV9WQHlES5uc4EuXdEMjwhs/JmBQ0jiP1Inp2+Z1ovJ6gMTR
KMjJOMQEUblH4YM/xrylI+Jbq+bRcdPb8x6kvMSH78HuAvDBDTAGiR2dAUDwpjm8YRTQnVhTujlG
BjSZ1YA1vnjfCMT4VmdDw8I80X8VEiXNJHc4gdjK1Ga4se9pklu185YNSHU/yVI/dmp6nw/i1Bjc
iqkEimcFj7LwdSam+TdHpzhrpgO2X+S00718iAcMyevhkakSxAYABRGCFT0BbUO/C4ZstrEtSK+J
9wjy7hMfvUp7yEuQy8I/4SgTyZOTth/IY8yaOuEng01qlnfF2WuXGJ14O1aqwUi6SrgK6tUf5fEQ
FqkLY1j7HPiXwtxOUJkNDEZyf7bkXi99BDEkf5zRKIz22iUBInZ6EY9BOphgYAxAMLwW9e0UuG/6
8F8q3jWPl8VeOx0Vs2PIQ2GSvJBotQ+ovKeXwZ0U+b8jkvq5qb9fnuElOJRNhffVIlEmPLRh/w2W
OCkXzNDW65T9BDs8hL/ZZz6OarL1bwL2yp+sz7hNXJQH7hiRAl8dIQdGR9RAojUm/wnQpsoZ8zpS
YsPSBuHvt28dg06bPF5KnTLPoAlMR71zvr1raFUPqYfJsrQGB8Qxm4x0tNLm88obrN20GMSWL9NN
qUYobGaQZPacLAJNj7Xx+G/HMo1jzYIlpF7nDs/geuDzaULucuILq1Fp3Ya8Chv659JtowbI0IEO
FTkea8huqvgEcSD2NQBB8WC7RmEsTgYCPfTtZSfNT6dTGdpwHQrTUtLOHgv9+dBVuSXW0c1GlTRs
CpgScmLGimJBkZ2uMgms+qsZkXdgkWNrJpIfqgzp8DhkeqN1gZHa/1bivU92/vPyCqIf5CW4IoPw
Vodew34xPm01vtL4H3eJdFGBOZHavvv38gtASgC9mv6YFL2FpzI43nWd7nbWISdREKRyNVr9bGCn
lNzKyppAVJrOwHhgm7V8yd1w+TFDsObhUZjCTBSM1u+RFZ2/bd4/I+zwOxijJn6aLRiM9Dd7cOHt
otutVjtM4fYo2Ttr9uj7uK3l9DfI7nLyAm2NsJwjiWAcwIDoJF2bdBLaqKkNN8iQ+eGaacipqvPv
yZfZVALHmc0w1jPS/umvJX11ThPMQguSmAOxbZ8lqBAyWaSZ8oQegY1YH3RmwFvgHFUv7LlLc9gq
RW4iO3voVKGhD+iWQQiHjUUAwjEX10qWKk7qi+qutWhIuf8KM5BfnozOekipomuhp9lO/ZduqX8a
KFTpjinlxGpvyJV0lWWGDhHamPsjMeofAo3Q1JUWvTyqORyudoMJF0+0R7x71ahzI/NeqV23DJoj
ATvb11xW6ikYnGF2oaEzEeJM1Bayjr8trBrozQ9pWjKl2FP7+ym2YDiDI5qF3864S0kfXtEyX9lf
RVbTEGBl/7roJNMxqXAv53xI55kfi1ALV9KmZkTpxQMnCF7w7T/1GPaC1a5mp9Cdf6LG8B9rsBn2
txI0/OtZfGLEAUEJ24FaC8TKfiF5XysjzvHB24vL1IGSiD3jHdapgB3zUUDn6h87VVZx5YMmaaVl
fk9HN/nTyZ6e0Ben2+KBRiltLLeD5GsWoz3ZIPw5cg3P4flrxWWnT8kcxKkfJy2opD/uj7j14FKR
rp8O+7ryPHI0XvxhgsjIjGuZVu1dT3BHifVk8dx8hRlQPq23QE5HOLIpG9xfWrbw+6IereGJJ1Lh
MivqdBPs4JNWgfV4vdw6navaaof0F6NqO2m4Hdi8O5/aB/9A+BoUZITHLiNX3X3tieFyLTEusyFL
T+82h5d/pRP50D9FdBlgTvzFN1vO8afTc5P/DgzYaiCozaYfwLf10uqjIpl2Kio2STnHukrWHYcH
4A6Jkmes3oZPVwkO0JIrg5UWf8eMhRcG7VnWnfeN2v58BnPvAF3gjdxHyFxRtHbSHIeRE21H+WtR
NuZhPS1/hfbxnoKbgPCJ3cKpxRCzXPvi7+sYPtVLcyZA22UDiN5Ykcj6G3IwKSM0iHesUD3ekYu6
vpUNBCxQ3sYBprOQXMpzqc75ot9n+TGylPaUhJp9/UpPrYkz/qjPX8hfAtxNOJawG+R1TEozK94H
uqrZ1vmu5iXeG6WcZZ9UkSkr43DiF88FnJ/AwZrofIwbwP6fsvLI02rtP9Vwgatn/OqPM3r4GamP
Zyj4njKOCErGZDQERDyvoYema7AS3XwajB92Oc3IXGF/QyNxHCZPxYse7+2UU/ZtjAjPsYQ5DqiQ
/Oeh9VyiRiu/1M1evZ/g4qvRJAat2IYpPhKyPoJEwB383UgW4VCxG4cjVhDRSRgliows2s4Y26yL
CsI2P0jUsFD2HLgSr/QiSCAodCyVE3xACNMnETGS54nWkbX3KY8OZhV4tmliB1E1M1qUjtUeYhSt
INbKux3XA8KuvgywA7dJAz/Lga0++o7m0FKGt+m6En66Q4xQ7mLldbJErnZKwJ+qc4t5gd6SGc34
EqkSEUta7i5Q3Oam0aZrDW9YtASbYVYLtOcsbC2CHoLBn/SATjivIA05F9ubaMbYqLO+Gb/zOdkr
xaIkz+fXcC2qTWeWE+IXg1WpxBsvsI9v8VtND4NojUgpiFuLtGQ0T/N0I2gIx+kF7WDAhUcZ0nAi
TA1fD3zb51STxveqxkkJpihpZ/8QmVEPiBJS8SRGT6McF9EIrqPGp3JUyIyKWOrG2Kz6HNCo+40V
6oKcnBZgho3FW2+yoZBLrCMgnZyVSuuU52AbToA3m+2ZlHuUjfRa/JXbg6SE3RuVgUlvmmHtLtmQ
VpG8RX3MPpIEQ6IrVuBTsq2NdciuhhXPhf5MsnJllEwJDf2J1HZVBeeqE9HX9Aa1HbvxsU2aEKZZ
/Xfd9oqq0NxtAtu0lysx0B2t2sSp91zx3/LyaG034O4Qb0iHUIMxoOEtEm1t8u/FmZ05qnXsDRqP
r0xG0lte6hbEqiFxzbuH1zVv1uRVxiRTYJSPVB1YULIiacOaatQrWQ6Hwy6OWSOkUIVlCTkv/q9m
plnlr7VqrE9A1s9G6g1fiRvPJLxAkDBP/2a93vi3yWXf7xMGnfZlMofqZ3dgQXb0kux3LlMr/+5e
khLtiSzTYghq5Vf5HOjmbfagyR2ONNdb00UBHh87TxfKAAk/DJPN6Y7YfrpNNGz1L4quNrSqUrWT
8vZAur+FHFR/elG9kGEbOmS4BbobLlDcrKC6RGaZ/otk2YtjUplkTtj9NgEQxHDwYhPbYlhhjHh6
f/jYxRzbDGc9+a9LHkr8iWhhaM9LNAaOgkS73bXvkLXENwgglv3SqQc5Tyw6P5KQvgal7IloM/CL
vQdVPuM0E5rysZSUTHS+Z4UW9gHK7azmEZiDPQbv/qXzZ21tkbvoSZULkdYfUa10uJJDVC0cdzBH
Shmwb2nbD/bjeE6M087Zcoyn+0v+or+GVGdP7apZxErjXBQXOpyOmm4bS3NcizUBuW/l7tAHYUxy
W5lZIYzOoqVb8RtbFT3OYjYyO1coRZdNGS22bvZcNIXqQSgKfmrjc9ICdQherVYsWqiwFJ2Rp6wM
7DLrk6CQcbanw2T3ApB20A2UBEKu4Xzqqix9ZWgC/D59dfP5EDFykhVBdpEPWphacALDEFcCmqB3
O6xhT1z/592LnHZChoEppVmRVfU0xI9vDjxO9qHqFCtrMbij9Q71+vr6ioSFRw0aZAUGm5/ifHQn
RUWLp9SqSyD6UaIZqTZLUT84vLq07s4aau0keIrEVwQAlrBOeKwrh9gYIqslorlHjOPOXVNTt9M5
/3mjiuEvli2re6A2tXF54kRfhtb0HeYOXTQ/H5MwyVM10a8rvpbIN2oBb1ATQibpSIU3alEJTMTu
/QayH/nu6yeHFKvsc+d4JmDbhTw/9avT7shGELmpiDW2SdpYrYv7V0+7ZeZ0DvWrbHarukGPCGDh
FcjTAXb4AyOOw4hMPDxWInMGOywDPxU8pNPNoSLMDFaD/+u+OEW6NhytaRvTHxUuPW2M92Dy6/fC
9FSNCnWqyede0yl+d82abXNw1/ipRSzBJoJxT9OzkT7FXHx+A9AXoYaP3bnSRdrdw4eBf3NiqG1l
wyqGy1rS4t6JflfuRh1U5X5coAIrLWk6OD28mF/92RtSw//IkxtDdg+d17GReE/Sr1vLjT1CUUSe
++Sx7HHzMI0cq4+pMbWwIn1/ljBjR5ZaPKUglnSQj1BBAf5qN6sjuvN3SW5dPemgKL/hYN75BTEm
J2HS4WB+4NsjqwXuRE/KVZDkvcZ061G9WfHY5w7gWxkDeXO5a8Nse2xQ/aRP+f0Ft7QNvvaZQCel
2QV43XdpDPN4PbxQ5vjaLYJbw7aSIIJK7aQDsfPl1K4+cA6ZdbG+fyTa3po7wNvgRAiZh0oz0Y09
3O+Ayy1sLp2ETNdDTrwM3ywAtU0eke0tM/v/b4PMiGx8AYqLsRy8el7/rr9ISeNMXlVgZCIXadXJ
OGi+wl4+S+EPvwGFhc9t8iQFFiFvXFMKlNSUnTwNPfyzq+1fLMASkI16JRHZgCiEbAf2wRqqDR1t
IOTOeU69jWToQTJsY/hTEW9rGZ9Yx9KkTQMauoDgLF0kBsppGhwaK4pNdEAfBlLLHXDLjZeFLTh2
PQ6D5frYkmu/mzk9s7JRTGRIQHLgblXvvfbjyyLWLk6vidXfOJnnA3hLRF2DLvW+t7X2qzn7TuI6
rH+xTVtkbTCVlVEjn/GCBFdFrfXB7FUyEOYAisj7tj38psL5/NKCA1U8yiEDBtBk9YwjKKuCbeIn
mvjy6hIhnQ5prLB9iuflcq83u3P09OKu2BtaAjEl4BnItbMWvQqj8CRgPLl9Yv2//iaF/aM/+waB
92i+R0ObLUsCjEsVJ/PE1uXi0naP680Ix/ur76lxQvQzqwiXu8+fV44M2QscoOUUYOvGHZdkCIVE
AFthYMaBtW6qvi9rjf5LIU8zkqqsvutmU0oT8dsV0awaSF4/e0dF9U9DzQqGXZD0EDSponOhIJ9c
hhmIjYp0TKUEjE8D6JSShqVkd8WVJgHmn4PptEfkiJoLbfwC+78m0DGWb2TerfafvjUNxexPm/Xf
H4Kmb7tvqwV4BfRgiVvu8yTJetqCIdGBVBvnh9X7Agu54+cANU71zbNLqftGq7UmWsDqR7VSSjRM
ja6gqZHvhv/U3iWBg/BOC4UJMlQhpsA35iTX+OR6VrXthmiUpWcpPc9Obk+R/+m0vnPz3ZXu/r3E
Cp8+Wdtn+scYZ7TA364HH0M5geOxTB/5mWDCn07+x1sPI81JnxdjI1buuKFXdWYslUxBYNBlzSdV
8Vo8cLHzAepsXFqoqWfsz/gpsauDL3qcpspnOgfjgGv5svAFNrsiTl9WByi4ldxkDKmYE0AiEL6W
+HldBOolbzq5Dvu9bHFY7OapNDaavXSadUwfX/B1b+vNrQGS38LRorb8AR489UtyTVnSYR4zCq0m
BwPBkkWmg8qjU9r+DWGZCp/b7zHayV3rpEBWwS8IyzJr0n/abVj99LbjwbAg39XzlzHgidj4Ye7q
La00fYpU5h5uqxuQwQ1ohNsB7ZoPRBEckV4eQAVVYTeS2epZNtp6kHfNMvWnD4jSA+fzfTxo+5s4
ZkQLrAi2/JRnhPBNU91Omm5B6zRlyu39oUWwh45juyHZhjmSTcsjPG9UBkj1raG0uBXUeFvJbi+J
1Tto0o3o4F3FEgTuYECTA7fZZvtVUke45cMbRCYgQ4hD2JqJQXsLGtEznLVqBtYvC0hkLfDpYrVr
HnCIClely+pt/jhCuPwzYXGRBZYzhQAdozWeScaRm2qlddtbAn/7UiY5kDqbuwZQBemxJ5Y/oAlh
mbgunQDR/MCPuUhXH4w1gI3sIdVP+HkWjzMC9n8vOaOf73PYyxnRWZCv4klJS/fAu8zRLyZqdzDb
wfLUEtPuTJ514m9V5qprcB3xNtu08iYBe4Vv2gqe5zPMFPw0xL4xs6CHnVTFUAquy+Iv20tfLx1v
QfXiwoH4p6MIp7Cqq35F62jfrrs/FXCj8tly4OHrWC1rnEBDQDnHFjd6ExsDR7Re4t3cjbuIa6CA
bzyn2YMeqCZea5fH1DxOFKI0li59GRTCxohVInAp1HUEq0CdADh2rz5b8ntQMHpTEuheblXnAN5Z
/daqL5bpAtJYvdyXVowrDBdnDnFZ1vAZs9CNY8tp1vNbIxUNa3Gm2e/o68C8BucZKp8Tg5IihqWJ
y/JUkwLaetj4r6wTBLBjVxkm93Q8muv7klXoTOmrUvTJMA5WfTMmz+pVG2SvPxbi3bAglXjLPLEe
98Qs9W3MKmysmlq+e8nWkUvPboyrSVEBE6yxC2aQ1SVLv/4WC0h5VmavVIfMNJdl7n3JZgVr3BBH
Nt88H5tyq44i1klb7lk7q9mUFFcnl9C9xwhdarUj9cU3M3sRd5JOIr48T66cPJl/OEK4vpInnTwM
jHq1/58inqOxkxZb5/G436EOTN/jcG4ENy4ul4RagW9ZLb6V/Zn4n18nq2TeTC+fcaNbwyQ1Ebi9
csWm5YxU9Zcfunzi4a6S48suMAggNQQBgMUPSH6aow4w0NZ9xMBTRUAcIOi9ab4P35VW7R7cE53X
0J8Iee6MOP/akueJ5pr3Pl8kA5M00VPdmQIjn/C8TO2QkXjsKMEZLSAy1VjsTFLGfSSq0kJyjF1Q
h7gZ6coW+0OlxtwZ65IXDFB0Cq0Tw/aZGo6ec3EP2GWHT36lcL0hRS+5HaWvAgTKxWkkAYQjSkMu
CxqnHFnM69xxV7ERumNPPAyOxdTqDYfC9MrkjSzSZtPaFWy/Q4Um+q08tZNdNVkErc5v/HEt6Jeu
LFMs3y7Q8rmNKaiY/oo1K4NXuXGVuRAhfnRiEUNATHoeovtkfKGjuUIzB0Gv4K/GXdvU2WsioZ7L
SPMNQOj/W+nSYsNMTdeCXayfD/1ocUoiKUUTnCTp2bgIHGmT3xcT95RzxqATRzhYYiOFE/8IfbV5
TI9Jzrqo5e93wZU9I2AZOfZOu6UNj30Spoh5lHOPtLgs3BIEFiwPbDxE+JBuF+2U48y/bh0wMOrI
cN0d66JdYv8uQdnBgcFP0CPBqTJg4+XJkh6h6CJ3sDsk2u0XjHS43WCwFN41p0oqBPv4gK8ALx37
YPZ18nK4xxrn7eHPeWeuGwboJ9AADGz5BKhqahjuaHOYSQkP8YcqmN7kvSB9Q9feXY6h2pSpiGJn
ceJCP+7kh+nhkDnhBlDZb0LZr9hlg08dfOgZ0SCNQnbF3pPsFy59mB+YSxQZekHSn7m0mABPNIYi
rsLpWeaDxRdgI/mESdbvp8pECw6bMz08u4+8wr4KVOLImnSbO4scSHt9b7/ZMp2bL74Yc8wT9XYM
jq3azsnLp0aajEi95meglcqB4rLejaq9dRX4aGb+JZFgpBmJVpW+Iv9H1+Z4h1kXyoKBOa2s1iaa
48BrwlB8/GOzTp3Qhs3iTI75riD4e6fnJ7GkllrTpdYujSrWY8jYizeACA8VbHjHNrs7jvOiaXsb
AV2rdx/RameqOphaYPl6e9dk6IJb3AiinCqoh7aQahFx0nyL4PoE6TT5n67UihFr4AYkM5EIq6ZB
9Xvv+eRDmIC4z8EDHDYKNSa2hOHHaMU4ZJgQgrq6vxAOVgfeMtOSscUiFRELrS8bKwcgSxAXNroi
j8VxD3NwaeE7DRdP0itrmCOBM2gb2BrzloiBjyX79N8ME7FKQYk7U6Kacx3slfx0xuhwmUsgD2nB
XACRGhPpHZ+9CuZkXYGMuRYzGuL6pNMjG3MCSlrhIZOyK3QA8wJx0xf2X66zW55hExgq2tevWX/Q
e0TKvojURZlf4l9sy4QfLUEWDBJFRFMbWudmTha/1c+c+vkP+tc3qyzJPEdTDkyxpUcNTSMxfdcJ
RKaU6xTBnWpCg9l2CAcTczsGIMwU6I6n7SEKCjceiyE0/tSQA7/I9wAax4+jp+Fo/s4xCF5A38Hm
gkYKLF+TjnX3ub2emlQ+zwP2GD4yiBNL5HLWBhKJ7kLYyaVb/l4UPM4qSNuC7ntGP9btg3mJkMOl
YeGUBgTVghoXsMD32qao7waqXUHH/CBveA1jxP9sVnuaZASzMt/VVTLIZoMWkIP75ErL+W/sh7tZ
uguJJd7nswdtGwn9BLO+QECzmbQusASZRy3YzdyuhqxqOkLz/V7FE77CRXoDQt2jRyoT9armevXL
cNb+Wn9S75u8BZHi01+hpR69hYvRQBw1+PCLqL+FQcFX0q1Nh3oTIOsOZXx4NpSsGpIRb/9BAqEW
QuIMApVrMzsLT/2c1C3RMvqN/2CkbFOnUHPATCGCrgQGTA+FNxFMRiksvPaaKeTWdfp45goW98bN
6lwyIWdS0vv9GIPp8iEraJSIcfG+kzKkXLQouWhc75bd2J/eLLsynuc1NkG+IVEe5RhBjyiP+zlw
OQmjAq8SuKB/pgNiFEly6FYSrqTldq1uzbCCt/bcTzRcYKz9p8PdlpHFtaHh4hvCIwfDivC4OyG4
Td/dUIIoVQv93CVHOprr78HJEW+w27Yf5in/6SOMSCgbXnNiGj8Y8twpfZxsVut/qaW2R1d/SkJB
lNFNofleYNYfRg1Dmtwl9yNwq24u4qHGDQfxcE8N9b03RQGs/ZuUbumHOJZW+P7YlKR6P6ebKX08
hsxt7HuJRchejuyOUBbGN6vHGOKVi65Gpn4MTq5EycCOFr9h8B3oyhTbkfWzS+3LEohRATqtLlDy
V5IeRO2H/TObDs3MaSFZ/iY9bf2y0fMwExrpLC+DwC9kGfAT2iIo6WMjQUCvjvxgHtSg8+r5VxYs
3BhDoKyo5bNjESwncxOBm8JDhZRyNrOSMV9qtJQ8qj+bWIWq8CQZFvUQS5UI9ESnupPKbzhWHy1V
6Cqppi3B7ip0KRRyktNop/ik2EBz+PMaf7IPdFJ8luJOeewmlhf9++FRcgL5EjQ5ojgXiHA6i1Gj
sLqiJIH3S7EZ5CBwkAvIDTJWAUXAu4mbZN4XjyEXB/BF3gjWCzeYu7ouHPNweLEwFagXrLDMiMZq
wEHpVGZqDU7VKGXkzkWpynGRF2rPcpqxJMszls3tyZ759WkAvIf3Mn4rZdPib7zZe2e3BkP9qdFk
98mkpuHI8i6aq8kwQF+0oKL4DQvY+tKG5M6wFDcRPzKjHfcyOLNRu7zMU5SK7VoA108TktalYsup
mDYOZ5tmoNtcaeTJM85hexvBISQCfEmN3T0ZYeZ64Gc1iD8xuaToiWB8Cxzxhu0D/I+9mLzTR/l/
qxkgu6tEw+0QjWk/wZwNocv3oWF/JcRO6di1jrLruo6ulm5SVaIecCoUP/AGHzGrttGPpv4Zf7k+
oUDRjiKiRWpzj5d7u8+au2H7DCc8ffIctXnZ6eezoGCrnhGEMPuBi/IQq/vP5aEmH9dSevpWIhMn
g7TGQEK8anGQ2ITilPoyTiSbXiFhA2bZnng0MC8rwF+y8z3ryskrMBomjE9v6X/XvmeOsSxYRAHH
h7itw/kdtXyYfPCT+vPS4vWt+nwmYeoY5BXyxJsGIcjoGUdCLuVoimqyWhJZiqZedOAzEOBKpAXk
qTLHJna3H40a7lHac30RMiSedbm8n7oN1iafH7xTlPd1ggv/posaYcozI/InYk2sAlE5DiJjUhll
0QnBtNtnqmrZ2YXt0r8DZN17DR7jERCNvQxScpBAMHIvdKSTbo5yjS/+sGmy2xV4MzSkzdzB2lCH
G+z3aAYsrY4HWnd2VqRPU3t56wVCLSniBdal5N7YnA/CMfvEMRDkaAEHLc2HijMnDAehxXRTruAY
doyANhy2FqHVP83j0nyE1jIxFoS1fShOoeGAmO7csRX73bTUfRO/88b3DlYWoyqtsOuaxzcSIcBJ
XyDr65xa6oxS/FP5Iu1F+ljV+ZECNlYu2Zf+twEoqQsTzRrC7n6xVs/t0+nO+VU+OFn0GmabMXce
qIgUM+ha/m1XGrMC3Jgyic2mbe1SLWb4Wc5gTInvlIRC7Ec+LEyW/03+FyUV7pVGqlBywAwa7W2Z
h5CBskT+nBr8C2SWiX/LiQroBlfjmLB5l6s8GbDM0FaK0dQDv38cA5A7h3jeRbMFJfFj80/hPIMw
zyvRHk2nBkbK3tdrHgdWbQ6rLogx/6gi4PgSUN5WdlcjhxO6+ItXqMtviaF090sjJRTbEnsVyT8P
ON0cBpuRIjcdP3/IVJ7qTjm0YM8/TwQra0IaX3lPmTAPlUeCG831XJd3pcd+s0XOkPC8oupW/Di+
aI0BQRHJYDRUS0qJOx0zXHupaXvJkMurg9GTSjb+msh5wd19CR561/zIoSoh0CsoxU0ZpOQuBMgM
xHgWQ45skJHsZ481DiwwhHUel9M+nJlnZjyQ/eVYIg763HhBnXt3R9YtHYNlzNTyl/UXA5OXVuXv
vSc0ckYD5u3NRZ6eo2N8ZH+0TzwOos3yTEpt8mL9ay/7lmONfnd364nfrqfhxW2LPEXxv7RkFmtx
x+0NIy9cuT7cW1zb+bvqGSl60E2feAkMOaCzTPwhItcbnydF3LQcdirT2LXwGhhKoyHII3ggJXbq
KxmddQ0Ud4mqCjYfrAS0wvqcjtjqLcP9moGG8RDWPp1YX91Gt0oJ1ScESHjN5GPlwl1BFsL7sITj
yMe/KKlrGCHLNMv70UmxQn2HIvKjW/huxJdS1XiDSqTP6zxwLu5CRB5zAaxySLohClu4jSIa9gJj
9QKL/yPxgXHZSrql/4uV4PHvwsFLEEOgmZIQCw/IKqbAtBMhNR7KiJ9sQH7Gwtdj/N0sugSTUXDE
pKsM1NZu0kQy41ZdUDI23ZYQ4/hylgDqRxlj+ai+rV4fgR3uTxGFH/V3RTiSohvXPBEJT9pLd9Vq
FE7+z8uCmoXolrxGrgdHtJTtsd1nmNrt/TnRKkKLXP9FJuWG0S0xbQkL/zpowHMDqR2xzOzSJxoh
6f9qVh7g8YKtAToBFHg7XNqjBsnSvxCnokbhio120d68xcR57rBJntjYR/PWcNCuZ5e1+P6JEp13
KQmc4fl1NFeUTinmfa7YzNV9xjyv/BTdYgup5ofXGGqYrxUheW5dxpPzuuF9N/XHIPrqx1Wmfkub
uryG2AhLVUGkejCwh2Qkrq+GLvEPRD25qPirrMqxUtz34dt5/vW8AJ8GQrfkVk864rCWS6dnLHPO
9maC15PPbuyYbHYaKUEBZ0gapbJkRxFW//2vDvhMcEMnn99llpY8xFFHTNRSjlj90nly70oNs7PU
pWy4vP1jhkgJnD5s0IA4NsGlHMLfn2HwROGlvV1yNmooaHvpPkQhqtXLNFaFwbPtG+SHB6cF1J1u
YoYJB1Q15T4YBCEGh1hyNgQRTpOpmWVeUcaBxkhXbplnOsEBPSol1qUW/7Xf3cmanbGnj3NV9ZH9
RSLKM8raKx0hW7VZ0epBjVVXukev/9Sc7QeEKHgKvVFqqr1xYyyaz7QlpeMvlmCwAFNiD393YZma
6U7rrQwzntR5OfoX8Zot/PT2O53spYquE1AItVs0Qr1GT6qLQgcQYL/4iWHqlyW7NmONo/SjLTIH
W4a4hVdwYKHU3UtiYs6s2tkPWjd+sprQGvSFqRxFnjaHvxsmKbiWKlWsDurIJYe+BXqLZZLXUzoZ
DTrkOLVNH5TilGoRT4flVM02GbEO9g8zV+KEFOMZA2lWtPVsR3UyszmAVL34OUyOGvpv9/6hFd1p
HaFA53IJNT+SIrJQojhYVQtx6EYpXFeFOHcVmVptzQm2dk5xvF8uOQkqNGyTOLNeF9zgHZCkLg+M
Gj7VVNGNGXY/aND5x5CNZ9BSIev7IFgT7ecNfgFDeXxfb4lWdw+Bx9mA3BhAeu3yOWNodVCiT5LM
NsvutcwIpOFPSGVtMsWmcgXlOi5z3iRZAleU850zT/AYA3dvelCho1meoxpgSCpgGKu3b3Yex5xd
WBr2Kld6dAjZ54mopSum1uS9W9EW/kaiWoHtxIaQzNzYbuXBy1x1aVEjz4EDNZXuohGJ3OvQs57r
ZCa4CxmR54E+XHpr6w+tj/Z1rKJRiUkCXgwHATbCSYtjcVlbRy/KFKvHVk4S+JkzDhsUJCJtRxS3
bNbOltPR4cQBszW+DGI8aZJnJ4liHKUJlVVGRz8LjnmJtzr3ZSXPE5mRaVP9/CSZ3Z9BJIOcmbZ4
ZgFbj2A1BI5tGge0h/CNXVl1PyKbdTXaf1xpCJ8fZhIBDCuuybdNZRKl8lJi4FZc4JwZsVzUWY2F
Y12QST3sB0tmpfrt2D10btHuJSGcbxgPO351zkGb/ZfzpS0RrK+UkanM2bpEtUZP+PcrGTtvDKPX
KzdNNMw0OXdgUGGN/em3AIzQn0CEVF1MJdBVtkycBUb7C+r1WU7InEax/JZOItjFBqm1jdTxvHkz
xb1P1ZEwSVfxrpG7RYmxaIXDY1j8Fpv182Y9r+PDE6ZV8C2wGQodyEHxM3M9BQNib+VPKBw3tbwy
YsF/qrWuNUbC61HZsP4+u+1wgR9oOPtHHSK5fBbtROhS5J9dPI+40KwEDXaopeG8V4zHa6goGrIv
2+//eNLhlEHVw3MaBV8VjULr231BoBA2SsaZsvf36eUWSyyqLEZ7ndbu+SofO5QKfrNN7teezl51
X7WxUVt6wGqFYVWg50vdTlTNG/IitgaBa9BCwId8NbSP0UWGu3wIKQIZv7AtmvUH31TGreflmOeB
V3OyQpnUS4GyW/FVUlMvk+8Fq9o9rfjNOoDsuZG9CknrS+tpkG8Vj5VRa5keAs/ZWYajsXDtqtIT
6mHB2jz+ctCl1soH10mqAsGx69IxFq5QTwV36fAdi+cO3oDtVzXfUyatm/WEltIg0KOTi3SOOvyy
j+qrz+R53MeL2MVmAweqS/Ljx80Ilmu6ySekemCgxNZa0Js50arUTPo/Bm5E8pX32ZFTYXcyaw7B
jIOiR8XiNgrcBcmwXb96aqqJkYWrZltU5cw1GlfI0Lan7ZUJ2uzL7nUFeUv036yyuw1i2YL/hs//
4QVPC4nZC9h+qXEv8Ruz5R/F8aOx/RVet9XWhycp9k69R+DstdkhUnYaCPYFbaZj/soeuRqeJoQ2
fsjV7h4r0KyPMd7ORMBkzdr4ifnv4Ocf0XrmoUAkDzqA58uMz7NCFb+ukQVpchlS3gxRtHKwT++0
KMO8XLzgc793UcUkmZ61bZZP4wgy+znEJdOGi1sDugaCfSYcUKcBw2OmaFx9wWAVb2K9etELEqOg
ILV8qPXLgTyMuoalXQP08xkAeUEkfjn9Bz87575vhY1gsdc+gg2uHo7g8F+I/aYAMdG6G1Ms8rj4
3aPbRUNSX469q/LmNtwXlhXfm/sdYvUWvBzBSI9OpDJ17oy0waOMRwOck5JYRpQSXmLQc+kEmjl7
htqxjMR5c7ttKD2QJA7Kt80oII5Z+BkLFTmYbCsZLigw6rxgmhEPN6ZBz83/SoHi7/AFidYs9mVo
M2jA837Xxb0Pw1hHgBTMpc4WHxCLgZj3dMNzYLMhpTIR5rFWnA2CwOKkQlFP30n0yxixAgtip4uz
icBz+S8fGNByXaNJ1A4y+zjTbBQcxrpN5K8DWzZihRDeBvO18GPMQYDixSo6dXslRMlFJO2TeX1Q
9g5V4hcr8i9rkTFhxcHj27K3YUXaQyIQpq4pkjzF0QSu0IxbG0j4oKpgBokxqaw3KjNK2NZure0E
+ztQYly54dzw2phqRy6muDNRqT6TJeAdGRtuO3isjfcn3tpdXOpWPCRuoal7PCeR78wpwWwp8Fd8
nvXht5C/1iuvYIazjOjnTejQ44KE6UK5L29fbHQb3rJ3mM4wu8UFtT33SpXhng0SPNB/ilz6ElLt
tMY+khobTLYPxjnGZ6CxGwIbCl8owI1KpQ6gIJRd1iVEK6Z8VFXNBSTxHomq59Lb/dbFBaqyp/x4
SZCtkU2Ow6vDjag/6HufXTtZtxapWW6GHIsFO5T8QQIubWIsSequYcAIXTLhSTFS8c6BgLTuvNuU
MUBaaEQ96kMHwnvWet4SeUjkBwpnPSyeyLAras2edkqdAZ6Ga7sEh+rJV975KUgvuYsK36kR7npE
PuxTwakv0TRM4a6RmuiXA6cghfQ0GtkT5gE7C2OE3V38cnb6+WFo3+TVNZGEEzzTh7hUjw7SQiHo
hk8DVVUHMA5l+sh2hgs1H2nkYKox9//Nr+vH4LKjoXOblGnUZULDZhHgjewf1SBsDYpOYuUYTN2G
EMAZFFx+okJM3EJt2kzjBSo+3Hi36eUyBpz5lLF5Tl3nZWNJ60Fe18ariru9UzzfN/ibHWXty2rx
fQfh5SOzCrLwb7PkN1E3z6qWxIF/2ixnEjCsDOfFGJ015qNnPq1TGoR2ipQT7Q1Kd8qRm2kRb4k5
ItjpRQguywU0aNZVI9TUM/asZhAP/2xj/+Id2LPqlIYt4RdrkdTle+r3GqJGuVqoC1eR+bIHLDvU
sxKFiVOTERe6exWylSI/LBqwUQj1/rw1/Rmpv2JSeVOJxLK08qeCBMmbkkDj3Wppoqrd0Ia5PA6S
Pm1zzzHXhC/K6WsxmICdoyRZeTSd9hPHqFTope84SmAoECpypoCTisu1QnVF+n0iABY/RqKaRjGg
0/nYxsLvRHVANCLowl8cG7rKTYZuQ9NFIte3nWHB3/iZxgXdKSOBXIRw+OG7tSYIWC5a2Qe9ffgx
jvH49ah23tAeufMxXMMmCwHoBzsWXhPoBpUI1bF5ZeIc8JfzyLy5yctq4MTLKDHiIeBoQXGtjCcy
OYIkrhdgInaGCaPeS2dg/5ajR5tWs7Yf/oC0FPH7MbzdXAaOJv9NINgzlCVrimeTUHMPJXLsKgGm
yyld03iD2ICi+dOXHuCkldpx21Jazuj5W8BL9qmldR5cVKgAoFGSNs/IE2cfMxDe146U645NOt/z
9bx7EDmghlR4Rxovt5SwNRhZR9IgOAbP8g+caAVW2QmJ8oc4I1Tng4Q4gPaSoDsL/6LSzKmDcnU9
CWiz8Kai2W5EVLLmFK1SI0E+6RFG1eaHtCFsxg+vaCwUV5xA1zn3WZgbGOBZf96won8lxYG3EBmS
+tnhMya5PctBsnZyzXG+IfVcNIIfLheKGXCfCV+tUfLwhPx0pFZrjesaUtM8JgLDlziCMM0LR9FJ
Z/tuTkFB7v+qVbGJr9OCs16w9ev1r2bebJBtuweybDJDM3yvP5Nu+Y27oPeb3bKrq6EMiyZHjTCS
TFvdJLggms4vA/AlPuUaOHDJWsWNjoQAgaUCAwMrBag7KvlrTGJHhAjygKg+RolWCuysScuFR/gK
iCp+Zy33/WvuCmVkBTo9lCC1ybhTqBMlE4jtOnjXXoDWJjwjolOsuCMin5WEphAuiFk8+RLMmnMD
Oz7hQblD8BlQBP48VSTHWp7TihW/bBj7/b7spQmejy+W5TiTFZyY+TNxSLO3wLLw9tBC2QBoHi5U
zOiBJfyq3/zdBofAq9pgv5qhmCUC3ZgrQstlPr8dZZzMNmB5gWk3MZpVMtkf/5RO5nkoYUwi2ytL
pQQDrou/vGNlzwSW2lj5S19zt1UxndlF4utbVZngfOgWp1IenTrUcGv5rjqoHAJhm0pNkA4W/ZPF
t0zdatBIMmA9cYPWyvm+vS5JSYbKItxowmHF4Xs3qZJS5rJ+/jYct61Mvi5o7J9t+qeOS3WBTOfx
rg8ZNKy7GkEFx+96NcZZHPPMtA1sdhS5z1Oy9Wx+wV8KchZCBpShOl9iilnWc3E5lODrfOD0Y0Es
CVKmV5aOP3mj638ejYib4PbMt4Jpht27Zw1hcX9O+ZeiI6FVcpumU63U7WY04RlZ0O7pOdgR/09H
X1wT1mgjIB4EBWGtEluFtUFkpntp6eGGOdSSIEDyFth65Cq1b56YwRfcGB4wrzK5Wei+Df4O4L1N
LXEzFK/E9Z64/unihT6uRpXcvL7ndhs5HFQUaS4PL79aPu8GFd69e9VQETF1DkcJova+cJFCH0hL
RvM56s4UR3v279epY62G36j8aL3SGFzns8b9KKNCDSDPJnQUZXrfjPmRTM4xsHDWSjrfzqyj5Clr
FE2XO+MvweFUEnQC8m83UwAzSMneUPZF0DwBG4yWgtkUbF3t85n4HQN5+CFI86vSzxUS1gPpaP6+
Z0QAh1/9roXsC0GLLSrXlQS1eMGNyvpholrj7vL75Ps/s9GsYxXRzsMewg652C4rjo9/jAQYXW9S
REL3zRUqqnNjqLgZMydl77nkidjpIwHZVpXA7D24jiu7daZnqF/3BKIgrOH9Bv4wS/RaTkhMlqiv
545+98pbxDtzwdS8D0+dk2wpgFNuo3gehdndqTrkxOrsiP7ZC14xjBOe+jFFlbZeGrzmFzSmbj7r
B9HnGzPricrh8+FRO/V7GxIuc2W/BprOjP/a6JlgRr1wHCWc9u9o0GXlkiWffaPDyUis3l29H9wE
Npr7BkOuneoe+DJUuW0unRkW7qOl3MpTSj211+hi3CxZNUivp2MLNAvt/RuwBmsylH6PWcyQveLs
u9mPhlFeJKuO1ZCIPMek3zZ/KrXEpAdgOn1DLDhoyK5i/YmlEB6NlvSH666CnEr2KAP3xVOvaL77
LpW7pCmiYLWO0t1nHv3i+fFknDcZbxUpxW1lCbz4E2Uqw07s/hohpXSlSViE8qR8iUzIWJhOsSkW
mLNQgejy4pdoyy0JqIPZG6I4DAnyJm1IhZDnpDjg4XIcjPXoGYXkvFzbQHgg8cBl00QrR+PEcRKs
ka7newJvO+AMgZOzpZ7Sv9q/bICSpZHesl89q1dJSt+bPW1mqkZw6XdTNxUcnRG2iuQTWtiaM4yT
zQZjoWuduxFRDNi9T2I7ORnLCNQs4y5xBowZMCc3L86/FtL4HwKfYaP7vYBW19JzGiTGljnOg2y2
Cci+Ks96uO3i262uap/5UJCJitelrCFcVnRecd6hl+JG35BQZgaJ0rFbuLEawjKuHL/2G7Q6ZGrn
X6kM97XLmNpXV20nO3lIc+ydLK61b/I5qz5v2B5GCEk+Ryo+4BWPdASEVTomG5FQGOCQ+1Djucsa
dZCM7BQQEroK+Y8F53SfZo7LdIWRMiZI4UBBBhMX3pQsHm4i100ODAE6vL8lZWLCPAe+I87B7zj4
QNAG9PkVzYY/rC2JLEA/kN09gsOfbyxQ55ZaQP4awYHGC+YCUmdLypu7zu3GC7RqIdZB55HZsyZY
uvHG7Dyyfy3DWWXb+/ShMq1vR9aXwSJdlzVXUOCbKNus9/hhqhjVHfZhWd4BSZ4RU9Ti6ZZt05eK
SgLD//alCAoK1YBIY3nRa8oYw4WlJ4Azz+MmbpMLVU3fpzYjeR719OU3CBXfRW+sDJfJSV7kuFjf
Rxo/F2zyFI9oJRAvK/tCor5GE6OFr/eoNwcNnvODvz8DRLWCR+9c6za2ZKFeoN0Ut/f2J+5iV9pt
2zlZvy8rtjqNYxfSlYBvvBTw7D+5kyRRiFCzJUHEXo40qthnkp2wfg2AbUBIKTGuP4W+UcTcp4/V
dpdHfhTRbum6wDUxiRJhBee/8XTQqX5Akite4M9wAFRp6sDFbynvQcwvU9J8VKrdb5bZqeD9RNfW
k1qM+h1j6aSFWlbWVuCtuBc7VqIarvXY6DwldP0fE6ajGUIOL2MJbyvlzg1Wsxz4bE2jP5As0HOH
LBKy/498zxXGWed8AhhERuayqsSYl25XV7tGsByINyrJrzHCcHUu2iScX1BfYnfZhnOcIQ86lGn9
m5YQPJ0UGMwt66yfGJaRIZspcZpxNjCuN+K3GTgnydU9fKgetirojemqv9R42q4VLgctv3xDkvDP
blucf4Np/vj1tqbQsgaANCJ46SI9n3iqyNXNQQ6B5wnsYV9+/Wcy4eCy1iaHN8py7hoAGOetfbhO
RSAAOSlpdfUp+s5Wo7K3e5xz8gaEXsV4fCLqr1JjaR8DMdng2Lnl4qR1vv6k+vvmCS95nWC2ALVs
KB3kTb2pdVRg9RJxXWYyGXhh8m34nXid7RdR4po0FTn4fppeC2e3URtTPflbGaGF0hVLJVvjZJLE
hGBz5LqIWxiMErA2XvgfvXy9WOHLR9zvtCyJnp7kf/FMJ1RoPRjxjt7Ho3BCIVNLRNU0k1nPRGZN
nteq84EyOD2HrtuFaa3M6q9JECHBbOsNSMxsRt0Qf5tpuLXefV+hs7HrhLb5pPJ1RdRYEyAiNPrs
8kL26l8nU5gjuMEHGXtizmwEEA8sQUpD/cpsll5A/klwDIcq+qn4tn9tqpBlZGFHk+5O5NRWYhio
a8QJ1mvUE9j4OZpm53yAmdRqoProJUnyq9NrmBlkv8nFWlDIQdyZDdHgp9VRsTS1rJNVoOq9wzjP
QSxtfflQUo+ELgH2S3bL21arHg6HClp/kyKGRYauvj+tjz/jF7dJSy9IXcm0yD0wPYsbxtu7rW5w
lheEjOT88+TibSfhPgz30WQB2uyOrJ5dSEHUcGTVjd5dDtR/CZivcyyPU0Zf/KThtNt4QMszkPD5
8YyU/j4yOUg0vA/wvvCSLt9UyGDa8MRVS2Gwm2/Jemh7+7ebcZbqhn0EwL626qdqoEMK6Nxl6c5M
ZsyMZYNZCkjcKaEMMYuwouVSTE+a9bRDIRJ859IeulMeimDGIrPaU3aAPNCqbepDpo8MQ5TUz0rb
9BxIhVVzfEtUh6ge/m443tuUP7hQwdueQkvrOMhfwW0JuSdeG27ooJFmNITlAby+Df2GJTPQxFCZ
eD9RAro8PfAr8rHTAwGLdb///lLoafJSDyUooXc7ogUygeRhdQbkaIYk8bsYkjZ2J77c6M/0x7/o
dWKKMU64BM1fin6kQHvzgGB3GO6pGaBWfg+d/szCyL+yCkMOh4lQ0RtqM0N5PWHweLUCtW0abdHb
U6lPGjasYp0jvTdF9VzjkuffggBmxnvAkhimfwnYTBbQRHnV61Qci0w3BHLkXCLKSWvUfyWNUaF2
ZH3Hz1R6Y7aGNbmB0bRkGolVoYl9OPe2YHKiBZAs679FI/E7jUXkHOnbh1k7PYMUioFrSCioPwWk
V0Hjozh5NdkX070A6CpLyLCb9TmEZPPHCGY2YQr1n9B6WHsZNSggvHwNrGN4BW1f00QMFPKAA9U7
59ZgLC8Qud0mgmHTuqPxSvMRwT63sS2EPWXVHjpxAR46c10fB9FUFv3NJeO1WzaVDTVFyL7i+npA
woI9pDIazewYK/gLgzHKUaeCgcZDSVAovUF6LgpZkC89P6xYsC7HFZqsIsQvFGubd7NK1AMXnOQg
AA8UMlxC+JjfgJPVy+EzfNVVnwS6JTgpXYoAyVCe9p22NXepP2gYNCXWKwmrv/CmNVkBvwdXtjaF
eHKh0m6FJvAIigSb7f/Hyb2qyal4gZPBnLttdHnhQ/WAK/JU4KhvgLqylCeC1l1vyYfGFTqxwb10
sc9adVtG+i/WujfkyjCcAxgjxKjCoqAn+mwRbIFzvVO5VlHr2x5osN4aOQQB+chFxdIcHTUWWgWO
oM3nhDWvKKjcj5Hemlm0l0h8sN3TWyIMC+M5n16agam2SmQEzyCkRXml8I9im9K6Y8u//mLl8cvI
q3aqu6uWI207UqkK2B3l1OP/P21eE6eHooG0K9LkCL+a6jseuqSZ4yyQhKDnW8Ee1H+Mly80uVTX
MypKjimLyC72RicaeC5Aw4rRX2r8gBXu6wezNkaLeEOOWX0JOdxAAwsPLUKUSWu6hFIIHABTjBeu
5VBvHarXtHp4ufeISYTwpDmlBJ5RJqwOt3b+gIEkg24GkOUZf4r607/lyEBZm9X5jRs/CP6deRv3
cD2UIRQbVCu9QcHB9Ziy4s4J4LqvKMuKtIrUsU3/87Za7kWhLG3sTvxmzrKEgQ9u8+exD7Gd967F
QmLE/oEefWvi+UjBtCERLgnBX/EibtTrKzQEznRUEAQM0pxSPG2K0iKGrfTfemeIdh5pwkG58ikk
6IX6lntUTK/bgCwqxv+5l3zAG0awwAluGwp7p/k8SIbjTIcdFhX2YPcSMmGQixiEbiZzV3GpOwvf
A2TdMYseHG9IXoQHwAq9rhMcQ/gK+un2W2Vnu8VJe88DIckc+ZnMn8puoujF11BC+lVAXtq21m4G
9fc2zut0/v2oyLvm2Bor9XhMEXKh4fjzCJP2nRlBBOPZ3P6BlnrzG6H0suOSoRjj0q/RX1ofBXiv
QpQU4u+ajejU0XGFAjDfcz1etMGvL9aS9vYEm0kvw3BSkqabVXhbQfBG1aZd7v8gKQosrSfLXQ8T
dc9iEC34K7KtetCqv4VUvZoybWW1BKlrYI5nYlmhO4PL2xOMdYMtx+HuGhUdovQ4zwqYo97A5bXp
l3f3Kev84Cl9fVCmDzEb5/xhwEqRvMvp6Q8y7GO9tEYEZZJtUTL7POad/mj44D5GlYks4gRsLwqk
XpeV7fhA/MOvqmdnEUKM2gb7/ht4cefW12qsmrwGRraWultwqVPAim8/85qzJDzvCksP8Qf2niDK
lpWcH2jZQ2JY64IrRU8lkXpWsphq8y1o8qYg2sIaIINrEujcFy2hp6MIpldP67iVy4ryGMhm0Owg
k24VjWSS+bTyOpAYFtn5iZx91Vl5IsL+sCiWDUOpv0LaMvOuffqDDqv2Lwd1zRywFUpIBYOI0EG2
3fCer3deMdRgTyTC0WpSHhfpOSrxl9Yq0N36ocjZCM+mhrw4swasegbpY1KQlT0weQU3DJX63uKb
fWeMKRHwjzwpep4Tho4yjAAzEQaF8R7tzJXT6mfxTfcBHjbzclmsXmU5oz+TxX3RZt8gHn+qPYkA
/sRKnb682LVmeuyQxT+nC9EZ1PnJtBbwhQGoIEocDbriMfpxaD8kRLbI0TrBvqSluZ0C0F7Gqyq6
YsOrGocTFghTgaVjCslF1KpWJrJMrCM4WwZSAJUqWoXY+TBR4Dw8RN/RSoW/x5XfMsIxTHkuppJ4
dftC6ZZWbIxJtd+ZkhkXhZLgwAfTbOSRyKu6Z4PQVuq/8TsdcbkmhD/4XG6RXDVhc3eFZ1/4zyla
QIiel9Z9sapcyBk9e6fzv04AEzDHkpj9GGWHh/rAle0rAVLTi46oP5/n2U/QA3XckiwlzPKRJO3u
NG/FgajCU/3itqX3qNxw51tPfzXsNG0Yu6xLLyn3D/LRWEK8tcT63Bb1rXBoUBfAfJZLk6Rl5myt
b4u2VPR7h1anspx9IMQL5LPNhGcD2bpz+pWHQxwehbQN13V7p9lR53Rnt+wzsKb5toOTUNsDTTlA
xvf7N46c4A7DGZgrk0g7gxlrYii5AF5P4gTM7w0GC3T1/HglYxMWpbh2b0F29oJhwB8mEZpNaABe
tSwQLTiLtusQXUg+Tq31DuiEDRaZwgznIXEZ00+wI5+SYfKAuzppHVGP2GbytGOr19WXVb9T+6aI
vvtQqp770U9yPDnI+uv0CxJJoq3rZQ5mWxnfqXhFum7XqAE6h31lzU+6q8n2kDFyvSjbXZoqwuat
+t8Chal44Wog+T+CPjuSHlof4aUlfZKCFPfk3QHufaraI6vyglj7ft6HbgKXWhLswTFegH60gwm2
N5aCHl29BkkDb1mwbPWqT3KD7F26GL0TgXqdrezHqWh5xtfF8G7/Rf2n7dSiYL5tq5dyDFxbC1ja
htUFP2e02eFvQaFTao7sezhyxMntdc289KowD84JPs6tikzFCiH36VddK9O3chUBUzb8W9U8o4+H
5IMj+Z8IMKbnX1Sl9jqS0wglJ2Iuyh/LVYFy8r/Rmj0zsp/VgjvKN+Bb76Oanax/NKrcBUuKHhI5
IrE3PnmoRFNzOohFMzVvP36vHXIos3KXEIFc6BF0BDwBEW2Yie59Ak85yYYrcv29T/6cwCC1Cgdg
lkz0paoAdzdWU18r/wtU8kdCwo5wyICC+z/W7W2nOWN4P0EP0spoz8YGDIBONjIgsLaITvKLvVF+
TdCSYmamuNyiFZGY7LcFBtEXtZkWcl80C2DDkXajWrzSFDj4bhk991tWENSonpJd5FsSOsds1oAR
msxRLNuMii2SEcliBnbzXJusIxudHilQ1mvUNWVdH5EBxlLMXp0iKtm6UBwnekXj7gK2+AJvjfxm
68K/lgM67UqKzgB0R8RrttXI4Vl/x8DSGiy6k1fkJHR3WnSH52C7OuLUvaZSqbWqJnd1wbPN+1C4
MbC5twEJFjJcLOKRT/jTUuceP26HGo/A8sen0kQ/2cBY1+J2DSsJ2VoXoXAmrmYWDcGjMfm9TphO
o0eNeHDhZA+T2ffNDMfGtvvTwUpyFESkqBAQEBpD8AkLWstbFYMR93obbgMV5ISGuNKiKogyUDb6
SWIGKyDOhpsfQwlTC3mmJew/FSu5JT9OLVcP/LSBXiJTxzlkKqqWLZLfwzT055SZmVIVQkmVHS6V
itzRowirF19mwOBjjZgxxSaVSXbhiTmwaGrA+5FA23z1gQK88/QizCgWsluJW4uhSmpkrxLJR4Et
uFYG7ZsHQISmCp0Iq4LnwWlvj7Pa4V8wpmaF16uL388neAhIotkSm6noOXE8Wji+hXDvzyLYorAE
EXBkIKIJwGSHq68O27co4t91ahqmrVtzgUMAFTZWQaB5MIMMCIbY8azx22RU7Z6+gq86wHIXxskm
do36ynJKUsmlu9WfurIs8ARCyabvJZqhNwtLvGJcpZPxZ5Xi/53ON+fZsMLXvL6toB8Mtsp4+L4e
DhJcMBrPerXY7paxE4aDLwlSVtBw+RPi1FxxMQ0bxDcCn6hOL2eP3yrwyWF1qCLFUt4d6l/Ax3ju
6y+RiktmgblAfS52wvYdrXLPHYWbbMGW+w5jX7107oMaOandlC7+vYHSgDI0NzwdGQ8Vlq+d78ee
NbXZp6z6OwxiFBZiSeqQj+8hGCYzqOhGAh7Ky4qlO0t7r6JN5Uv0MmgxrpUf0PZfRJKo9gIyZJpD
Gqaftcg4bRPB/AElWvCbVIaqaabiney3bo4IAcsKxD9zo9Nc4vyWQ8E7gpmD2vt0nAxGsbjsFz4b
NLLMJR7hL6QP9YEdOXbVQY+o/NyysZyDwi3cqVwbu0j9xzInnJK1pmIGwkG1PaP6e12K+nfS2kHN
RvPBnBErLDqstzMWvQgMFuqyqMnLyykmvkShm0gPQB6Jmfw+rgGlMZSgzfBjqpGETEfr8kfEBcSo
alNkaZR+qFVSPKLuDM7TUUz/BHqu0qfjW9naqEgeK182HhvsUDWb6zGNBX0HqTagv8zU3zfw8SY/
ufT593bkI6qJrVFq95Q9qmPNOidYZRW2VL68NN7x8ZGMIhDONqyZgkg+OvvFjPANAFiH7lPyKwEg
5G70qaXV/k4FMgEkvQD0H0MPUtdP/d3T+tdsfurQ5P8Yc6KrZsx27yXbyB0lVZzycz/rpR5kNrLk
tD9b6OL0MCihzUZ2aDWUT2MEpu4MVDjR7MovYufaEWfPkOr+Ta0VHzy3D+9Ux4m7TP+NkRF8Rh2G
j8Xjr/bRh/lNMzMkhUKCdplrPZVdZ0YxTzkMHOfLiSbmVaiDPTks1QofjyKrbG8fpyBoDUnPvl14
9qpKwXuncN9PytcJVWvOt9xmYKBRIv1nClJlpKKtuhb7I52meB1TlAWqBW+Om+MoZf6lPf0SlUoL
qlC1Ca3QMHY+uFmlVhDNJPk8zIrJ9syPfuBF+AiXmxX6Eax6dBth98WkqOFgVLu27DyN6ZQfPL8U
ZiSEJXsTyStXIePNVzl44r1dlDFPNHzQuBLLmOKB9ondLv8xo4R/fXp7P5bceLo62ffPwR28Ki/9
TPeVCx4h3NcU2aVFh1pPX5oFrmFsc4D7Ykk6nIG79nyGYB9fnSQI7MX2+Na7PlJ3csSeB7NZIUkX
bXhOyrdgdItS8FtGc3lAJ0TNITz3mf/febAV2x+cmoIuhXuvUG9Wy5nHQwzrKMzlFuNwy8K5cCCu
98313YRo5qSD2uyakRwZs2w1Jrydyy2Q3QwoXqmvPVjV37W/LHCTIRbV/zmOXqkvzfa2EzaiZrVz
CxxzR72mURzkaYX5CPbSA7id2CLVI1GN2BWpSq0BqBhcP7qrESFJtzqo9c/PDMTA86YAMccDy7tP
diXGYBVGdYSfJYLPOdkYx0cPr/p9pAy2i7a9aSIqDiSY8kko2ZltMvIEm1VrZQ7dX/Y0Yn+80qFj
vCQ8QrG2+jd2IBlntrV+2hgf3AuY+Q1fX7jYHJAq2mujgNWadAeyIRFXa9JM8FZOHvUq9mH3aKg5
3MsMP8lFAydKxfGIPDDQ8LYoCpB0nN73TdQ8NE//4nndicnN509S1tKZNQ5Z8CTSyc9gaRm2Qg0j
bYmWHRj+qDG8VS7DLFzTVLq6s9LTcdM09d01FnliLW4IdeHlzIWmAe3s/zhZgfD3NO0roaxyyY3t
mMu/HoQlCOIxFYCzoNNThFQpT1o39AGjlxshERvV3ueYr7nZ0G+LjHmUEVFK3kZENGpA96x45/NP
x1Q9gi+lzlvBC2z+zwEctkDh+G7DHrHRLGHxO7uhBkkVNhODY+Jvx8CvLXjvhqCFV6bf8BuJ3LfK
yWWCgGcVqrZFUYI32k0IFk62zjJXfPT7m9FdSJyEEJ1lBey9PhlK246uAbDNm8STMML4+2IjUTnz
ab/LDBkufgzPNNaBPhDQoDfgrFbX3BB775zMfwAEzBgQ/Co5ap8dgzfLlw+Z+wy2tY5qXaQk6txh
3wlP7MKTxjYeCIs50ept1wZ2ApUeLT72j2LzX/cV2NbbPv/yZEc4hE9w7TfYoVjuqF3qLHUpOppC
4m6hXYGb2BL4ACUg6BQ/ngLZDA9fDbeRG/9bbJfeijIeqUzLfN490BQYV4494jEimCqeuXOf7b9w
jUV0hr/4WDHmez8WqXPu7I4pgPSCtup2EalPmCP2nf/YgNfLUGvYHBENXIYBqO+Z0wpDxU3wRyO6
IX2wL79MYps1rt9vK0J9Eiy8bgw2JEA5B1RnBFTbnr63qSmmG2ZmF5xBBYtqEj27Cjt76J5rwt4q
tz+IgbJNYfROS9kkdRjmL0CTD7VwutRlA3R9YRoGJ1AliR4lHGkMF7lG0Vv8a7X/5Wfpu9SMhyZD
7xOCq5I0xd2Oek6aZn1/XwxowPnIhT0o81K1EnH3ba3KiXtZuyp+GgQ8NZdN8siA+7ksOScFLiMU
BAfiWcs8Nrg5isPiXCOsmjeSuwGirNgtW3+bwr+SGeyoRvmyO4u277RSUAZqL0a/Np6HkMrT8oon
guNZ+t5wcsHPrEN6Y7KR3gTpOJ5T2z8f529cgf9lUu2GrEyIlhsFX0Q4qO3f0mmfIYXC36lj9rwC
iATpmgH48ZvUKqygW3hFqfmtR7EyVs+jZtR+CnGzYNQ/OrOLNBiJOtmqGmY3PomOmzdzLgxx16MK
Th/Bo1Bsdiy6ps/SU6gX/z4If5C8SkkLqO0WwQKUBq49GCyqCUoN1aSmesoLNQ4rmVRA0AZngEwi
NFNOAulEFey3+SWXn9FlJRL7amUKZlkI2TmJ4b4QS59ed7zPUnH51nquDcA+j95jkYKlPA3owDti
A2cY/f+R0NDyef148N0JPZU7kB/msbze04ulha+VSvkmkYsBBhUipXPp9bf6YVwZTVKLpAEAICaU
8MVq9chs2P6hCr/jqCAPQR6RRIdTylI0ndzUK0dljikzB8k4zOLGmaA2Rscshyu4tqOP1VGoS3Q7
pTI5W/YpEKA3DuyN6I21REo6DhqADbZ1WdPgLbk/L2EsVu419nj548KdvkqZBtM3VKKTxIwLYx2z
SSmvrdZHgLhkTYjl486+eY7aFnfD6LmkfuHDZdD9F4C/KaA37NP3cjGEFKWVz2rjEGIJCmIbZaTH
EE8/ANAxLHp0v7rTCMze7+X0kYERxJVAqbhwBsF3SNrfaZ2IhKOc7VDjCemtgKxafyPTer54ufSm
Iuk4GeKWxv6cf3xjgcC6NOQDBXjJYm9f07RBsE8AQYx1KM+NN1htLatzbrGuIsO6K/7LCwtOX2fb
eZcQUE1mlzq9utBEyqUmopgFMCLMCqWSv+9FR90Ph4hTVjcsWG8y6Yl7HZXYXv0aHY9k10RbZSRr
zPURknfWsheAE7qTK8BD3xGrSSjpUeZ+ZrAdqHJyHsG6JLt0TuDAQACHnwMXknFdB/9FMnWSVr6g
f7W6a4WcaHCTJRJP3LClNFuuQ7dIRrZ8rFRzAEDKDsUryl+wJqyTHKKRv4hbRaj0coyJlFUtiUhD
8KlMGHRS1uqcNlwJKRxUce5arVlBocmfUDfB80M/LP3KnLogM3jnyLfs1YK6GcVV1K0oyyvzxH6q
hAhZZed84GlS8foohI7/8QjneK0irsJYqPGSVaGX5higWWuQ59q3ks5zUpelvnCLNFXgbig7kszM
AlPwg8AZ1h4YKXhZF8MXFfs6WiIIGq65HdJTwnWKXDlOcNugofFBsJ6ga3D7Jo8SligTzIu7azpg
hFBUrOpWkYZJfa5n1xkfNIfK7b7MmIRXnL6S6X13OfmWe94VH7XmwF6hWt8rOECHB8KzLNFtVqck
wesZLwSYkfASuig7iKPxwhEdB3drGTHAXURyjp/EIGhrdQVxSci9EEBDQt4IdnnjVRh4eX4/Rm3+
8mAXt0rl3QKFCgPoVVAbY2OZoBIqk7ghK4VS5gU+c8uPAlXvGgsfABPSiVZxmaT9OB6onuE0ESU+
JJkilsHPqnjWgfSTzQXiqD8PSK/eu/G4HFXrnMoX/9uoKWyL1ZHurJqLkP3AbkCx8rW/fq/5ApQe
sXHPCp2Uq4uNpF0CqWjuVp23thrsuhmiTwWfu+9oksiQ+WqzyMG9nFBilIhmcyOpwRrfR0AEFlJ0
UdG+vg9pT2HFvegYHj6lMGkb8exk9NaGyIwlbQiFIhuZ4VmvznLq1Zo8Q2Tmg6x++z7ZcuSFK3d2
gVIwSgeFjdkX5rI0O6M/QVcuay5hr3aPyv2/D0K6y9xgLZVhdQoQ/dWRcG7mZbA1YEbOi2Gl3Syg
/L43afMOF6hPah9sJ3Jxuc5xyIXpZ+0tnpYRO2rKBKUhaNfwH6v/TTvPnaXd1VLD2gQMgIArMheP
veC7XpcjOWLYBIDhUmvB4yGkCksB8CPdIr7XDg5nsRC4ZSWG8B7NII0ShpzsWRKM9rB0HLnol0r/
schayQmCxkxvxuxnGyXXFfAmV5QyocR+zNCqd7TV4oWBuflh9XLfLDh6mgGT0yvbF5vYdo/7C8Y5
T5xEn/T7rc6OBWvgsvkyVMG+ZDDGGf8N3LklVj/l4fJTGsB3I0DWYs+Plkk5CUS2V2pbar1B7+0G
97MR/bxtOYjKoKDCB8a2GhhtxgGnf+E8o0a5XP3i07fcTSVPVxTedE/0PvoO+tGhAjSipiPk+R8G
P0cIRR5zT1c8HoKiKr0nq0EBybuYBBPJrqMJ2suA2saMRRLmgq03dWq37oUKZARElJK0vj5V5XTr
YNBywzVJQ/bP5dn73EternidxrRaqgLdS6UztS0JpPIxyLytfrliDTqBOuAiGLcD7kKD/jSxIv9V
WabfHWaD1oyMEQg0X4jM3HidzEO4TCX5ZKnCP1aw/yLmc9OJzbkULKIJSHPReNAR1OKAGrqEmZhY
+CVgCOMiMsJpc38Undmc28/nBXYrsPaaMVbsB7f3cZm1ARd+SPHRkUVBaYSjzfVTKyM3uYJ1iYI3
pBsfdWpxDPN7vo6g8Ixbpb3GdCsEyLSiASKcfl/2OT6b42WVczsC5BiFrnVgyTA07MmcPz8BglG6
PRP7BHWqESBinTF8ABvvGCWN4cb951yN1rERGEirX5YqxpZP9wFBahSJ3XLXll/S6txVVIOWKFHt
8sMSiUWsc5yYcPc67uqWGO5yWzJlc3aqQf4mQZNWe59WRSOg0R3uZ0Ms4jGhvEji/RzDnHde3Slx
1ji/yY3Wm5c6tEIUvT1E1Rkt6JnnBgIP6YgF03AKm9XO8nPXzM3uqUlCTrov24BOLhR4Kt5vbrVg
pGQ9ODHb3pQ1QYTBw0Wl8GnEW8eKYpWHgUEB6/AKD46BzsXnHKGEg64CpSq6mAwuHk9J0bo7hwjF
EgssdM3OIiZyKpAFBWWmZzmnBanCvhjlq/P6wAtrzHlcanH0rVeVP2ZP/F6jBQrPvgmc/j2SJrHv
GTO/iJtDmczS5nibyoa/XB602IWl1+7szILJKSBvFMzd4333oYynXDH0cX53d36nGqcxeIH5B6KI
dHilomek5MCP/3HGEk0hGADC1QA6W/7av5kG2FHvkepSrkA6zFRNVyOWJQe5rn0wP1hFbFweMjLm
OlaOV9uwXT8qSG43Tgerx2lnkSEY3OFPRM/T9nbFSxQJ6dgQAzyY6+kgX4KrO2S0mp9ddFNFrC64
ePVQsgGqVS/D+cUm+q2R7ArGuSQM5pgnbqGIkOO5E13A3j6sgDFQayhX/49vbmoI5pCviXQtazC8
Wt3C1TiCmxmIeskyudmP8Ci5XC/6MTHiisUgQ8LoP0T/O+Ho8KbNHnPXkP7VqiSgQoGvP5SfgGwS
hxLxBzTNmcQKu1f4wKEzuF8apA8h8AUq9afHqr+H08EMGoQcmvtyfwGYv3QyCFB0mJT3KlxssjMC
ZGnbvzDHcB36wm5lCTScDaiZNze33CQAnULx7dnAyx4Kl3G3dIEYSi2DvWCzILLlAHQ6oTzjN2DE
GeXW4mCYGOwEyj4yLrdd5h0xD2zxrPHyJQVq4ares9xIxpVdtwqb+YqEiMjqTlOG7ZeJj/MS5sb4
mBKaZcn+0b7bcv5NsBGL//5NuGtj+rhz25KbjaSSCYTUurVhQIxY7U0X/nrAAN6S+sZ+9ZrUg6vw
RrpVHbvALrlfeOqRreLKbktmm5uXLn6osSoBGqcgEGighYZ18fHMB3VfVv5+qBqJm1j9+FGdPrFG
B4canmII2Hz8JXvSj3pc4R4ALaxfxxxj+H7jNfbWX+YbIP5R1eLZOkYp7wpUTAHsB+kJjC+4nnmC
jW9soQGHDgRDAg0sD1YPv7gtVU691g6DKoNb6HswUr9r6xNFwzlE9x6CDSqjU4rqt8GGiAlXjNTF
xax9xalLoD1TAqkptbn0NHPptF9Zh7+FSCFaepbT2VLvjKCNg9rklGygzro+oqC308cGxLHw2Mx9
KPAq8uWzaK5/j8lAGuTeNhhWu73yQiPQi5rEvOwmH7prY5jTAIcfhsv61b2Rz6SGcPdRIQahS9vt
dY/1v7BR5CS9GGKdUXpkww2FGDgA/mTHEozGUkeXauMDxWHHpjMQsL7Uad8/WZKdTHE5x35qq7T2
wz4M2YDboEdrtn2TD5mt3WFerFXzkSV/dUsx59ZuNSVgiloTLQaxcTzCiJFBhaFDNhU4WEkWI7eG
z+oBNAlxOAfoDa+fbW9PKO4stg9ftH+1gqN15bBfsi9Vz0/RyGOr+8Xa8n+OhHAmnv7dOevzMJ3z
5ZnspnuaNEaRcPcvbDapzjAu660oJ/hAo9xf5e1wYU9Z6wpwbJnV+n9W7H7adxNcS/rFsr48nou4
m5f17tU8jBDDTgYLGt11XPyyuBQNLZEQVjzOJb+sRMa5qyF4wyFkzkKFUseH2oi3Im3SjXgHZnUl
o7jPZZU9xBAQxXgxzoQu5cjfXxNxc+bfnoNHrVMPRJH0vqz3rWixr3/PyPpy/z2bmjJ+F/IoHmZA
SkzZL7CKdMGv3NE/eShgJV3WAMnzeOMmqaSGlQVXOLi2uuSuk78noRpQvUTqUMOgOf2bxSzahuaH
a14SG9pepgNf/vwUqwJz8hys1QeR+jh8SKf2h47Fj32QbOpmdm4WAVuZRz6G8+BHz2lGVzAjEl3O
jazuklsY5oZh6b4WtOqxn8pFUKw2X/WNcZTc/2sUpg9M11Lru+qC3TuP326mI/4jC0nZT5CX2xX+
Pa2TYNqxG6Nb3rHEQuKsymx3bc/L9k6aksSJmk7dLUqmIpWD+GtvF+E/Ibt1GZXGgRdJA/jZsZC9
XRrtNFjB24pEhCQ2pOpX35P/VeTN9yXbzV+0HGICU31Wxp+nSvZ6VhICakeWzBEY4yt4zzLY2z55
5NCVYROn9bqoeG1M7x7L6aSPd3fHHjMXUr+lwrCzvECXItuwP9hruoElsvg+cMjc+m3xbBzk6BCW
qmrbqZP1C/NYdu9oR3Kmi0HOaHZRMYLfxepp6lsE3Lv6AeeKGqoXIHQ4+ynwMQDiRPIrHJTKrPaq
QtGlmTObLnyoz8FEFM6FCPVMsV7NP7shoYkRW8V64uFe6n526nUECVR+i0Z1dpYFrxPCe1K04cp7
VspG7tgRBM06XKg1+oG2Z9Sa7Mh4829RlNsVreCROMa30BH/Ay3b5pXNwP1Vh+ue1YBccBt6Z9MV
Wl2Qq4tSEajmMnaxVBkZ/ui7WoOBud0yIYUF6lJ/4PT/wBOHkLKsznYSAduLtvTlKOAvE9fDBi3l
mVUpy/iKKKp7qYYZfC4N985ocUP3RLO0VowmVwIqdyhoAhe56Lyahlzo0442kdOvaqWSvo8HDitL
rTikQimDJIeJBfBkd4pyZqwM/V8mgbkRBS/1avt7XnzOosTJ72CuxAUIKakNy6X21tL9yCTEwfzW
yof+8vJsqhfEd/SRCVwqCo99QOVM896g+4LlEQIJYzlOh3/vPh5hRbdApNapMQAo7ijdRjynvMlI
MBlf4tuivPg+eS/1JwID2wr76ZfHKzlTHj5C3rtQ18+KYlDLHNqp9M9UXZJqEDQ3O/X0/0WEJPRi
6LA/GFnJKJ5elRCUZacyCc/wAv+5v0jSP8N46BibQZjd+wzW6pAQtfCTDRI+WrOYUfgUtOVfyMwI
7BiIh/eAZVZW7Ml8c4Z6bdqw88OD4YjE/J28QyarJm1YSLAS1rGlorv++8ShYhjWtQcaq6a7YMHu
NEuxB5M4xaMYr1QELvdofu0tXgklA6KashzZlNikzr7Z9l1+hOxrPhlZKNMJZ7Ljadqot4LLRow+
V0VW0KuW4FzL0WyspyCUnCFm/vGjjgmlWgGsTUDEGBEz2UpOFJn0otsYQVdZ5BR0jvFwIxgczYaC
ja1uQ05k8W0/KUv+yLocvYyspxxasBIMvaCZHEug7GME6usT7mHOth5a2gzyQHpEIoaej3Lu7u18
nAUkEbDorNc8YsBxQSnZ72gMgVyYA+RMU42ZZ90MK76VMrzLevSUBmBhrvK3b1xGqVKN9Qb58c5E
5/MkP0emMoJSJH7TkTXYPoQ2LJaFtScyEn6DazTUEFu7/t78KQwyP416X6BBPWbPXegiB87Tyj8H
lkdn+KUu4OFJpi1vEwmF/aWEZ5/AzMFEV5v60EoF5DK3zM2K/4cWYv0LszuvBQ04MRzSEFA1JNw0
EyHwzSqmWAgge9UMgjinhciwqCnxk97yOPrm5InNUXNl1YnGzQJOSOA8dRWL57iU3lwY7B3BBc1l
cFaNF2TiZu+zXlRFq8IpOrX/RBke83np6LJVEhf9oq6mam5mygAypLRkMQ+QczRWShBrmnIqr4D2
MpirnLv4CrpDKGxjtmgvnyX4qxrYRLeR2Py2cQAcYRVqcs5Z3KeO4fkDgJFNH82eDR28VIm4Z3cc
xVpc4PS0CgPNhfNqCcP9qmbx0T/MkI5frC5I9VjBaisArLciqYqpJOt6UpX428AQJtzkC/9dgtDG
IT55Vekl+yQ+M220Xtu9oZc366WKsMQjY2Blrq0AhWlSComNgX6Kwkh7y1AqUa/b5mWH2YyJ5lfm
kazl7xejZ0vnAvPJAvqh4Kt3/vDAClgPQSgykV585tFsZ9YtsSp/lyMxAaHHQA72JBuyzmGgsWS3
jdh2STcv9qY8M0FHVCXdAym4xUQYD00xRUtPogn91kFLrhPTSTzhAgrK6quSiMyCyFaLuJb9YNjr
QL26CvYxXnZMcBoCE82WYpb5XsRB8Infjn4G1QwPLVK/wToBmcv7KLIZqMmDs6Lo8j5xoYfsuJSE
o9ByFPrLCwo/xiqNd59TcDAf/mxZVpLpKyOiO0ih1e40vIPk1rbVGoFramGoogoqPMC6GEyR9TEu
fq0hwrrEikqCedS6INPzdDUXgQWK/enLGe3FtHbx3IhtmTgcqnWUkaOJMSneZS1Tvj15lsaAHDS9
17fck1EyTGXdBITDKgWOzDeiIbuuh2JRvpxrjvNs8Ellll8EJtYbjhMBrcrftGLgNrM0C81qEih/
aCwLN4W3TCQMu0hwHPdZ6guYHpVHyJi5alWlVM3Si+XxmjPe9jAC5DDyVQKMsgYwFaMjOmuh/DSc
X2EWhxyjZonFMpkqsoL+ufVoI+y5bGRsD9omgRPRwvRXvxDEQABQD5uWHA03tteh8o4bd3uXcc8J
2KAAui9AUrw0xwmf0FLxfDRZ2ftmA9NmQWyjzk/hmT3g8JlKDgiD8jtxY5+EiFFdancdLyx+rBWR
ote1U0ZrQ5rm7NH94kSHKbLxUA/9Cvjsc8hA+RX6ueqRR5frFwXDEE+rio3LhT+tkfRp5oUtfZmi
aDfHif+EEC06Xu4XwlvPjT0llnqnkbXWnLddMkdO0qxP8ZIERGHMkqjwmFh2Ucgm9reXHjWktr+f
tDCs7r03NP2QlY9Yfx09/JJd4P+blURi53c96jN1jB2n8g1SV9xL0euqmZPNnupYMjP4fpy1ZoAS
mrNRMrDHXbvkKilYumn/O4xtoTDDPX/oooGFOrCb9IA7+69PoOWX3HbkSmYkl/Ejo+WfNb0a2eRi
Vrp90IfNNEyTKydrB/Pn/InMLx5DeAYzq3cVOUEBrY0uBtdb/YRnDfgit9sRca/HT3NEXMZ33UB0
IbjHswQGrmGenZPWr0v6d/baqrDcKBUYLgo20B0bDeo31L/nwqv5SOZVhL2+4o5kGis26ta8L4uP
9ysbRP650vQWKirwcvxY2oowm0Ec8gUNZ0zwgPWCTAflIAYylblMsAM210xWLQ0IEYm/ZyW+/Mky
YyVKV0TOblcUQc7YSyESNVhIfkAWzzMblm/+7E31x0xBOHfUFRzQUKtldov747L82KXx+6x+ZV39
9I7NeT/bFpkrtS8n4sGJrWRWLhbLlp2KBd0JkxtytA/AXp15sF+usWjrv3RNAuoRSMegxka3U2tN
lR8PQXLUMN2N3oTeUJEB/u9CdK1zOcq+iWGb0pkfmQyEn++pPGw+G9Xw3re38YgtgzIpU+Hjz7Cj
EN8e4u8dT3lZszYsEheXI92mr2G3HFLW4ifkJBKrnHHYuRBhjV4MueVqoe6o/XnnZJmK3B85EyNz
8uzH+bMeeuPDiIieAj+3n3HFVTiv27Pevs+8qBNai2Cj7IZjUgrySU7+HFN7BMkNoj0atarKN9ve
BxKhsHrs4vSYROMVRmXlT3XogP61Qw3X5jgksEsvzZEklDTYHF951LiCvhURAYyV/9WxC1qvprwX
QoZboBeSbG4v86xGaQH3jkWVxmVfNDsxoOudUSuD5tRju1YidDVvOFceXPHrt5sE3Z2J5ADVOyVx
CxOUrjqZMC+k7Lg0zIH0SL9yDeC9T8Glk82y3y9QsrOiUq/9f0e0XONIlqAaNyqQvPaNGhsXTTyR
oAt0tLiant/sB4z2nZIwINHQelzYOWjpXVuu8AHwe891eCs8dcH7EweGJPj1h6TmJKIMSqFNtBrh
jh0iYH1PfJITI6x2zEkN2ckh3mZ0n51xLSjdgZDvlh8sDsaIvm90a4Z5KKwYwlA/XdcBz8uA1pir
7iAWBZC0AW3NE7rQcQFW67vryg6ssTLCeXJcHcijlD+LrGXp1X+Lh4PFPGr9h572RWr5gJrv/vs/
nUDO8tvHY5qU7DKXVGdUx4CySNb1v6wwdW1A4uNXmUH/uTAKqm56S98HqidAS2v3kQhcHsN+OvKP
oTFWEthfyl14CQJOoTNDD4eU2R9a6asyT6s5NLChGKhn5VqM6obXkrYj3o3Qm6Y3YColLEZEM2oF
OLwFDhCbbYEiGj0P2x+NHDdPwlvDpOANPHctoVCHFLcK+fUDCFJCMOzU1tTmB3jK7DAVw8wxofDV
PtIRSL9LdjqLyD3XkF3XccDfylWeI9sxJVrEV7ekjy91+FSjRrxQnpXVh2Ba+40C/WhTUYltwHNq
+9UakIBjscVRkDYixv+3AOdVFuyu7t4JYh/m22l6n8C9tt6Ag7X/OCiVUEnViQZDYyITerdZKzHq
/FPYAvaviYvlCT7/BwB/IDV4Tkm+TuhswLPR3Gxb7fo4JVaOL9vtphu3YAOQuX+MLIDuvq4GHchp
eO+OwXlJ5T+zUqLS/3R7aYp5KA7yg6Mq2wz+1fV0g9PIOfhwvJtJiWari2NDx6CNyTY2iIeUazLY
/AFTXpZNnlsQKBtGfUJw1jNftKFhku6IaxAlR89p2Z5SwY7FkMD5B+cdrwj9i8pt8EpZNs1YcaFz
0kJKtLgcTmoW9oVdDieDf4HmtroNhOYaYXwRYbc5TuyAIEMOfQoim82CdoqnEBAI3x4hBcC//2Pc
+QmyMGP+D+mROMJQNvD7vPiIsSEdgrBSYUllK3UqpIz9QT5Q1MBQt6nvWU0k8YTngVTs4+sYFFwF
/UxBxsPzo+HotjBFPNPLJ7qSwp9bEgMVfrPAO+xjn6CyOXKYAHzH8VM3y9Z3HW8GUXT1PgDKkqR5
U11pvOLrdk8tSSsO1HF3JCKc09bSY3reIRsXtutVPSL7cC4fdTnLnqRu/oF9463Z8MlyPfqzSyDH
ZO5wG+Z86hlqSP1sYrjRxH6fAadeYzwf3kfu8aH7fKv+8ke1sRN5DGr+bq8qRwn06tMTRmQt86KR
en3BUd5hhR9wM2zuV/QbUhxhw1kDHGmsNfTXLd/3HGxdcLT3mO2zJtDUNSScnlhtGlqE68OzheBI
iiiqDFFARbaJn/9hYxZPFoXWTZc0TbaIdsPOefjxc/XTEO5ox8zxmtkKasGHu2hK81rpl9PgnR9X
4t4EkK6iereUISnwBd2polLZmp/7bdq8VZLF3mgMTs2Zbww7DxtIp/LqjV+a5tkginvOkGaeZsbc
UzANjyna9jTbJm5Q2AL3Wo6GiNFCmbHqYZ4pSWsixIz+wF9QjnvGCp+wswz1DBzhmb+3ocQtEnkM
hyOLZpesPTCz2PI0O/7JvnGnrfrUSiae2hsSjtm4vvoc6KtK2vCPtA54C89sTbBs0A/hOf+9Bp+E
vh8GLV+uoCG+vsNVFQBm+wxERM3bSnORXRTQtF3bJeRaFwU+9y8Ez6zYg0GeBEuT2DkMNHZiup72
ot1alt5Zc3XB8Zw0WRQyfWQQ9eSWV9wDpRy18zP3YX2wQBtHdTnG2iZX74LKqZ/qL/6JLY6TFE/D
SJBcJZ0+dhM+Z4wCgcEQfFKExoolHBg0hDIY32uan6Xb+V0LFtkNYKgWwveor/TteA4BQhrjE7bp
KG2vu5eXyrXwa0hVlJyyaTHit66UJ+bF99OqXk0cUZMvGnhzyof6BTWHJzv+TTKXEfTm3UERxSQN
imtvPtEkk6DdtoMTX693Ct7zu3bpL6NQ6Fp8bXY6DA9/8T40xyKV6wn7m2Bsm75fxTFmd1pUgxfw
xUBh/d/qcgrrvRLHrFOsIixqPjQNkzfuFGz7j3r1x3PoA/CAYSgy2owy6wucNPXIxag6d8zlSc5x
dAxa/Ghz/PaDzJ9xXYnNur80r6N3glXLnqouhTTlf1Rns9i3JYEx2cOlU0sN/+ZnfM/luPjKALai
EaNRBKTAg9owm918Yi1abGCORoFMV5nA8roJHjt2CF2+g7CyNNcsw76X5m1+7zf0f32VqMM/+Aho
B7n1BwvwsGllupNoHHjL3npo+J+uSig2ov3pbAWzf+zpo+7c3/t7OfJFhfzeYUwa1sgmqsTvS/35
FckbaZwDgGvJhwhFD7Ud7VdebEd2ZZhjJ87wVHdd/asIuS/nrpU1zBpR0Z3P4SdiNpv27GdB4aH8
iCwzVjr0hbxKHqFYQTrICUoDBu3l/+rL6MkQu6OgY1c3gRLljTiim5I5YM2SkI6VJCMGJrZeLoxD
kBXCbgFj5WQXTfBP6WfZqtx9hmKaftAkfrJvhN9mohIO05IW59a46pgpwYjWlyB7gZO+aQiYkmuN
na5xWQl8qYITL7RUpFxeaXGF+xh2AjcZ19fX8MbH7Pb8d55VA9BoIpSPSbl+EE6oaODCiLSfz11T
Rj8683W8PaTf+rqbDLFgUqmjYlqtYNzfciuvbeFekABTxAQISox6iYjEYzP3acbLdPrkEFQ1MXhQ
iMvtFWxR/tpphzFb9kYYTMbqw09j59bgAbQhLzV/3MOwZVPqS/6ujQoCSIYYrYqaMKcFROaMM46H
LtMME1xgy9pXU4rrEW94DBo1OAxWKf/sLGfY+3++ktJq2eyuI7AAgTMzD/jVwbhk9Vo7X2Kdc2wc
/lB7QMW5EWcL8EztNOtBMrCLcHAE2TLBx2MAtB6scRXwz8peLyrkRA/0ck70kc+jpXXNVrGs0780
Sixqss1bZrb6fbbdNPm5glEkIVu6xgm/5ksqU5jDPJhHde8u4GS9a2PlTK8dxiL84g5JX3KS+6R6
OaawGb+03ARjN+YwVBemtABVI8cU1YB2qvzT+kxq4D6Tku8CoUXXWXb+6eCdLijiXr1le/ADuv3E
JDYQEawEHFzj8QgRx2MwY8OUaT6unlHFZSBMHGKCzLS9noXjJeqGPBa3HNOrZlNbuRPTwMIkzmwu
t2FNMU54/co6Ymp55okRz050ioYETvLpWQKaBQ4gHZm9Pwi19YfL3E+xzi7MC6WmDG4FQ/NQAF6h
iTSqyMBz1sP4Pw66OpCM45l6SFPtdunLYRFWQU2sDJVfjvf2Wo15WNiDZ346HjzzgPUaplSi4NSa
U2ORqqG9LviYZL1yIpMduvUNj6luPsgW3/Tz26+K22B2YcGDc4sxGpuqHehCUtGfwo7Jbbe+DTEQ
oUdfn/vHWxapl9HwgEzAvO3HhbzwKI1yQzdRm/niVf5d0+wyQkj3Cg8uTYXhyXNFlzSscXD/YWkD
JVqR/TuCDQHipxMIgwTwNs0sWpFVuU4C3Dqyen+WkPtkBQ4kn+ucOnJqowd4tOSpzf4RBLI6Bycj
qHKqkx59UsD3fg/95pi39lVwSy8KXglMIoVH6lJFKJ9PmS675SLX8uhU98vxp+OWMiOl2l4qvHCv
xpWdse6KiE2spAQiJp4UJviroORwfixppR+bxDRLbXizML8dCKZZK88j9SskqHqrMJgvtbCz50LT
5seDpCGp0WNX0KFHvBEtyErtyQrDfNEzRyfmaJhZOUrrYIs3gGKu+C6Q6eZ3yHN+3zpFNYJ8tDSg
GVQfwqLkyD6AtSAxF2MAjQxkfrt5M2gByyJtxickWWuxYCN2QJBTQnl/TXZRNprGqburUeLgyLHy
AUcVpj0d6LxlIRVZOpZI2lfM0fPGKlrn2XbmHixSwKwkG8oHu7ZmADrRgLxoGtYu5KMFm3v7C9Fl
jXYSHeXjt3e29TIwM0ZsgoXlYe5QYMD0dSh/kWL/VGJe+mQGAomO7jk4xDU7FyD+yAFxQ+VEHm88
TIOCI23jwJRwdHwo+EsM+VQ+j54be+wnfOXBgSUNAJSmFlQ79tbJdKVwrBmonNlDVZwkHuQN7Sqz
SxxLP9BMMpdfKn0JaiogbwkLIiAt+Bq0pXSiNQlk9IATJquMSYB9hD5A3QN0Pk+75RpRAihm9rdN
S2kDynrwYz3WbJfXQHFPsKZliBfaBh5A2Oj96vastyy+rmjwWBpvoVJc83cJcurY41r6Z6rnGheD
eYopo3nfC3tk9D8Lm2qVXvicFh7Q6cOG0AtpDYFVSGrSdXrZaxOC5xHRjQxVILirc/8TCGOkMSwb
mMGC8cOwmC3x/hmdu9zQ8ppdAgeKLFJZSOxY/9bQx2LuBwKEcJ4ut1JzrXbmi0dzi19meSrBKo+o
0j6+5WCXXQaOGINxCV8QmkVndxBujzN2iTcxFdtioIn+iEPGYa96TKaPPoVQuqQ33+776WmieLfD
/NHyi4EPIEB6wwn077ZMEhpO04aKiGYX/Tb+S2El5TNuPm07KWeToUQrnOQmha1Td0v8W3JZrlK2
SMbZj4p57Dv14N7pPX7iSF9Rt4XsevQ59OjsBfiRsTQvAZsspr1GzcPBMdWC98yTdP75tgvMfk5O
CAzkIYPVBmP8NoCYZMunj221O3Ie0kugOzooCewNB315jaw7STSCOGPI6sVpxlXIS5ujjCIbwGE+
vTjWiniaXxUAykYF1f9yNpNgbF3ZL8TNEcDGaiwzAwFqnpYAKOr4CvNtWfEryQ72aoLXBOVr4eax
/RCq4ZcoIHwgEF/Mv1YYJTrPXXEL5hxbR83nUjLZDzjNF28kxLFw6MFmBub3IM3PtklDowKsymR2
nXg9s6DZCjs6CWb16pFUyJJ+0Jv4KSipxatiJ0hmsS3pa3AE7ZnFGVJsd7fO963u51xScJHqKxP3
Z4q/cYnJWyuWlOY41vTn3CX4QQjiSIbfF/+FWhq2aiArZZycsrzUgm+UI8nVDMjZJesi/lqILLDZ
44KX2SORQ0tggzblUHpcgiWT6qnPs7bS9XkZyUza2YeqmAnNF8+hAID17Ug0g2rxaR9ej4UO1N2d
Pzu/Zvu46n63xuViPI1y61MgFScRbwnsAok290yW/W33gw+sXgKAo+84yD3QOP9HKRW4KvLwOS2+
bbtbE1+iqQcdsKOejgYiplljSkPkG4tBcEhJNc0D2ONJOVZuU/KfOULBMrzVnlQLKu8ClKhYoag6
1YiQinRcnU7nO6rz42AHZVUX4sokdotHc+FDc1MwCuqXDnWqBzutPRlG+Dn+LxMW2BsULK+1Ta9x
/wgYc15KYu1rmOzPgCxTpwAcbRUElA7xYs7Q5S08l/xZBbIJ09tu/XvmcoEc8ny/PQBVnQyVZ8Sw
HdgtpinrjjevC8YIrcyrneSkf7HG8KHS9t1jp1RhaWGwpiNGQNvcj4EbnsBiyl/96jA13GouU7Ti
xFbFX3LlVlNVsyPbwrahN62MlFOjaNeyaLX6q/+9COcFCXrrIGIDvGJ2Gt6x0nKnN1+uWe2nTK+Z
hWYaL1gI2jStLF6V1edk02znMwUacKYGZk864xBhuRG7L0R2CS9QlUg8hJ2F5cu1Auyv4hQAskN2
uBJVTKaUgPfDITT6nyHn62LOlPmTry76Cdon0ujDjWK9TKvE0byYLWFADLEBKxQbEnvL/G6nf+49
JBsJnWvPBlpmATkYu74DRwkp+Jm1tqq4tnKToAAbnE2/ohUjxi6oB46CuGmL68qKsabYQZIitz1/
BGE/JyrthE9E6KXsBFOQu5sZ/8Ou8q1vF17+HxMY4Wb8IKzWd1Dl2n4bKNhiBag4blvs1BuURRXx
OEPZGAQCnKwfE6MnQe72JV1CMkcYufCifHycCLTqwC/pG7fmLpVJ+1k7s8tpnTVboViSruokJNQs
IIs7ObZxgyivfcumL1varyfV025O8i+CjW+V4q6o4n6xt6dVw8mrkpkwfxn5ULNxGqHsHY7nmKrW
DALHRoZ2cEAhvzGv2nNguS3ZXN9yca05UxK9s5mm+Q2Qzfcg3Q/2CZSWdxTvylj5VbGyWwwyG1ko
FWvNQgoYmGeqyX7E44bZPjTV4x0GjQIeOJG1undNRoahEVBebpWbkfU22pzvNg94QQ9XYH2v4XNt
mG4+eG2JaqlI+mnt1eTnKCZEeTljNjgcyD7r3MqTirrpNf0zLK0z3ZNNE7ADKrJ702dDdNI9ydhj
ZqgPA2LO5WMsNJ4cSNyF8B6WQGBhLs0srHuF4BGHbd/IBS47bFZJp/Thv5EZ8pnw75L/xtowSTJ5
yN/jTRO3AxCxjJvzqvpoR21vXOpk7tncjHf3FPqHOABpWOH7gc/kLMV4/xC4qExEWV1SnlItQOgh
3PAt9cCyxWEABMs7Rr3yly5O9m8EK7WEdm4eouX3MNN7KawtxBpzZSq2jL/jBWXBvntTvCs0mYGp
ZsKex3MSSIDurZ9EmJcdrW9z1SRYpOk+aNUoLjnTvTZLCDkGy+gwOXRzb+juy+c4yvz7NsjpIprW
wMkn5UGy52B16Et68dYCBllA+l2t35TevFRhxRKmHue5iWxzAC1TIMXUBTssXK75t1Ip+fcKoBWU
Vhjdg4N49I0ElJDsHiihX5QkxVSZ94ngAwfHz92maDJyB+ftICK+VuKJzKptIXkiNpyZRmKEjmgj
NCfy1o4nbYz5H0zDC/JEdQqUnsKkkjTXBH+6pcr0q57rnM2PkiyRZI1DIOHv9eSDa7IU/Eb3nYtM
CjXobnJj45kImPbLbWrQtTGPvDr8sD7RRrFGTaDsG6Ed2ekt+TwXT7PDBCUP2yCHT2BInZ/MP34h
VpE+koTJu37n1aZZAsJo6IKosCcjTPBxfKoteVyN0lH2TCkQZqWRljz/WuULu1GVHeZ7zYXMAdbh
/CEvbIktPx2sP+8+drZxwtmXGr0aCWms1Pb29MjH50BA5lLaYORsK1h6c65o08hHNSRSzlBE15AA
vgHR0FcesdjlF+WVNWATFZmYfubQQldkTznBjgldECeKxcAqe8R6OY2JFlQRFzvl1IJjWihY3f40
svVwUbUrkrIU6aynLYEAnc5F5AAbCHDF+cOLOMiJmQ346pM0f7A0KjkpBfrezsb40qkAxrQU+p6z
XvCVWcF8j2pylsVz6StwaLs5lpmLROwZlB92yatKGcxU6J5sJz3SI7acGjjz6etAipCbPIc+F1fc
tjXpulZbSUmsVSFNJmCmkW97xBO3rKW17TA6ONqWzRgs0bWIUqsTgJ4CIST1b9WeP6SErJtDg9qy
X1paztaSFd2SUwCimSgFITMcqfuLII3OC8/oHtB09foGqtnscPpr4zRI+e1MPKcXdc/5svuTL6J/
oODlR7RG2P3TWuYtzAkhzT7Zl2O3RJPiJYZDaBfYa6Ys/q45/r49EGbt7xyDmsRcWIIi7i1uiDDs
/DnfED0wimskN47/9Be/mMVfEnZecm6iSZA24XCa3x8GFN1rwSJJekVMfsffDX5Z9OATIjiyDmUa
kIRNLj3izbssYpispwpCH0vjmxSjxBMpflLbGhWhul/fwj0edA9G3SqWE4HoUh1qpVA18Vdyuva0
3p+lpoHzo7+FdAiMMX+7GBpD0cDiYjoVAKBSNc1Si4oHh5CeJy+CQwdRKyYUtCUlyMhUsCunwxbl
09zopAcPauAXLaAmBrgQJIc72b8sSf+fbrbhiOM5rwszOtuTHhPBBKBIOA9c4EDlvOPJc1Ys7SKH
KObrEmO8T7T9L2PXej+W1BolxQjLsEKmkQ1wQH/QY2TNxP9vvogfVGwUh5hM7vI/zYnjnl3nXkKJ
728Jnv7GWDZehXzNhhib5ocVi19iArdksmxAXU/obwYvYVtKBG+dla0Z+A8OJKUCpf7s02eFOQSv
nWlEb3koNW72XGo7H2vzguw+CmhOpNrb42QSvoSb841W75agDYeYdHIsQ8flWoFGq37W/yTojvJp
4J+lKxRb1HDJR1kCMZ9lTqu4Mh5YEYxEEJfSTMMP5jOEFwtJQFM6hUa1aZ5PdxivC2G6uObo+Bqf
jWqrPuFV60d44pafCpy1uU4dd9TWuokTcD+4gaCeVi9E2EwkonXm/lSQ9CI2WwA3OjuN+wTjFQkr
+W6hxYyunBcHK/EN+1XpBMF+CJux2VGg5/cqYg43oK3K4nHXrO9m/N+7mhzlr3x5BJ6XUWzh2cbE
rmiBK5SY9hSVzovzuE3gAyzKG+MV6MqAiZ+yUO0Vc+tOr45L8j+2UGfNvYaSDPl2n0oyaOBeg2aL
U03TaGsDs9kbb7vFnejz4gXsIFChtAOWiySmpF9at9MvSiaXUxMMjagPDPaEqFGmDfoturlONwEU
0GZQQiHyvI5+WjAiWIj2YBwShb7LS6q/BBvdPudxJ9jEPslDrtUknto1hIGV81d+kTMDB181eTIq
0Ttmrdcajpk16uKNoWUgU6/+QSpXHjgVbpir91g1qAPuMfg2xmF+hM4OBxSOXiX6cNBsxPC40clW
JoqXT0uz9LzaZVPciW46uQzH7GmV5iAavGdZhRQBohkBr9rCfU71IKyydQ3/ndtqyYTIS8PCgiLL
6Omm4vSP+t2rXyrcDfwnwq46bGeqaBixWZiIrr3Y4PlPuSoEyEy1Hs3Y1IjPRO0TO4GxtoySF0zB
hkTGY0NaOiwi/KFRszOLgRDGvMSr4fDw/6tngGRJe6j77riFh6d/qeXCaZKbitETgGQBnOoK8hPq
Y10Pf++CyqJO3B43bExd2AsMlFoVFxcHXlj4+YxPq8z6WjAAg+V4mTKW2tvJSve6T7Q7R25k9nf+
sAxCm1K82fsr7azh4Ff01jne0jzOkmAqAgGM96ZKdaDc69SJK52b7PtujxersWErXEZPESn6ikWu
tO53qtHGyv59i3xV/ciZPnwWjbFFupgiKCPWylF7Pf2QWVeMzcG7PRfwNDmH3tVYdHUONyH26yEv
sBd9Mv6EOYPbcW61Cxq7lwzkKt4x56wX3AXhYtVhVJcxUJfaBdK7mE7pJkualSp14KsswLyeOwkA
KAVnttHi8QPq5zq+6l8Q5K+uXykq2hWGzhfHwPVkFctaN18HLQ0L2T+B6lo4r3IObtWJbTGsow1m
ChDsM4GBBxDhoAIp0mmLRgRylLj0FbxgSfgjwDLdd9VneE/76no/gHQAHh1VK9pDuS8y9vWt7sD3
hOhl2qzaVMhO87Iwi9PkBOAgHGxcDY1kaYKDcA1V+BUf6mYyyY2/9l9frD94BTfbP437JqQhcnIV
JscM2vhnF6C9SGBztBeVp+PDiSTsn8PhBf1IVTD93n802JnSrwq01vXqaAlQ51GsRqhFLdMZhypH
UGyvF90cC6EqtEm32r84+/zqc1dq6qH6ks8X1dVNvuEb3bO17VPWP3Z7Quv72UPTGLKs2PFALlWK
ZeixmauNJEc8QK4uG91MnChdVWk6mYj9BiQBXwKCc2knvi9NDLEjTXwU3SqIM7s0WwzlUHzmUS+s
JY1ffM92VMDAX+ennXrHtahrj6KiH4PtmyzFMJpvLmyOA93koAR2OTNl+8UOWNTUVQqr+H1LPO7s
d4DdflfkJrjbfO7bT2l3ZIKPsUdatvjmM2J6Ct3iMEnToCHoKN/dOCMT+82kiWI3WRueeN1CzPGs
BMed2mPssmOU/Q/uo4Y3WIDZ1Xtn/zbBNnFCuGHAdg4p6FuQdgj4dwdzrzBmlDSjMASo42OJEh5+
Dih/bdh4ZzEOR0pyXCBu8cLtsDJYABbLSl+0fqFWB45ttzzbH34iOAMezXXhq9cGQbFv3/AaKUw5
/9Tlpv/B9OkubPGjd2bogjG87ceOu8H81loPA6/vPufQ9BAmKfEJV1qpuxw57ouuPiAXc5hNXNrv
GtfPVGERGWDWl39LRG5rrrX44pcTfDGkp5casJSO/MTS/uFPQd2XyeNiSgWCqMywym4oYwtFNPS8
SLjgDXqTobvtiRgCLhWkIDZNKlk9Oie/1VgtbfqakADcjgrr3kq+9InUWJ+E9IC5MbXlsB3SKfK/
QT/h8qrF6G7uRv57We5gzdexOM9kd9jUEnjt6knC2M2zBf+OXaTvjTn3B4cZ9gy0R5J35dlY6ccD
Ko3Fxxrd1HH+eZN2gptgfa8tyKqlJj8JM4pqHNE53GZqNPLrT14q3nG/ag5uSlBHPzGWAUY1qSQw
5y0DzFeMkB6kbjxGYYgJOU3RogZHRAnGBa9+YaPz91BAjZIZwxaWBT/zdFtO7dIVuCS7lxKQPoZZ
r+tfm7w/aq1zf+5Gn4UMjPGiu4jVNHpq3Lv+Cc2rUFCX5T/KholHaQbDdj0nBIrOKLuWeu5WMmOg
QDFRhAXYhflYMWNZKQY9P/lW+hWJgYmR8ELAOI4t6TrAnE/bUWsh8yvB2cjL82eotVpZTbs52kd7
BzZfgqcZX3oMo28PD8/s7XgXKRgqPDpke6H72TAHupAM+dvps3hLbiEqSbfhKnYvoo9OCvviYmrJ
y1GHckTGbHvG22CgKOye0STXCBuWx4Dk18t2H1T0//b7Nm3Ih6OLZ/kVnbJ/ppNHMufJ5VBM5QdR
muD6z6sNjUQs8dH95X4VVrqjWXlO2/I04aTfcpblPxUuB+D7RA7pVVAeLu0JTSnVMIfsx1JDEFhm
sQN97qylhruplgXtK4tkYmGqAHwZjwcUOT94dI1EEVgz3KyDyPUwAH9LU8IhvJgfCIEgAAtHYYlt
rGAqgbGoAfRclS3SOuIk37D484N9ZVcgxN6NpUXuUlSMdJkTylpHebVexUcHuGfs8VvUCqPQNZbR
Vjm6VA/+EIXYFjCUftKU3IhAPt2z9SbNLYvisY2dJH9akJaScKrkt60v+2HA/N11zpaZLwd2NIQu
070R2uvNcy624LoFtgzu5zKowSvwB0sriDExWhSUY+75vUEkxd7VUoOG/5iFuhtnG6NXsLxr36YW
7b60XLUxTtMxXZn8zGRBeZf+71O6G1+SNCAWW+4rZayZVvJE9GPudBgSkjUswpEBB4FtOdoR07DO
UJU+XJPmOX/CctlqGfRykl7r/3ZdFYnumaoLl4rScX2/m8Fiv2fEqtg6veF4ywQ3NZDXA+m6BtvN
gBC++p1nwU07zZ+zqI18vVo7OWByVg2J47tvHNF+wj+shsk4o148jKYG2weixZSvFGjz5iekbr1M
1KQ/fe8iZAIf3ooFTfyELLi74lh6iH8HdvUoIAr6UvnXZzzTRFdBacn6u6ZIe9/K9z4vRI0O0K16
4rRKR9z8qLpU98ws2z6rrQHxE4bJM+liug+xRlnV+eJkOv7tP009SmCV4CxZ9owSwFRbSciTaDPe
bvMLFmhPA7+PoWlZ2EutEwGtAMa9yYPhbeX7EN+CdBEzAJKjNUkMy/zil/2i4wkNGFsj5Ye4flnU
xMiOOc83RjA5cjMBdBT5DQ7AV/xU7U7Upcru+OLAj3Tu5Dnk/Jw0xUUr11MGl9Ju6GLWpKqzpkw1
GoMXwCQagyS/tUgtJykWpkw1Tk8cY3uNEP64xC/lkNn/WwybKu0PNzQWkdxyuv1qxp/vPw1z5V7u
3PADN7BlRxbYCc6esiZ0w1A9abDUSBOcCX2KeDLr6suRUdm9EkAF/aFcBGO4kqC0PVxe9onsAUz7
vhMm25xqbzxBzlC/IiyVq3Po5AEz9HZkSjS1hJxxQ6khUXmdVwWfLhWHu4kAxknjUHePvd21UFuk
nYXdcXz4feLHOBEkkvL1dDrUAxH33C33C59aCiDUwyMlCgAoCg2NOm5EiyQtNyTUWAEpjbP8mp0h
07dwnW2b9CCwK1iMKXbPhsHXGkW6Bcv8QRobAlFbqSDrwo7czRLF4zJ21uK0qplxojuxSfEQFkaH
trhj+tVl6vmSVRrG6KMUAYyrkNVkCy/5mMtDy18Zbz7GDnebThh84OSE4jtp36EaehJhv+I1IyqI
Au6g2XD97sVq9SL2QDx7XZZXBg/7sbp6Y6aOthoiLKFLzgLpzzBUnP+aM/C8GO6aq+fuRw0R1zPU
kgALBPxa3lhvDMdq0dgzZomfJE5H6Iczj21dsy3G1AbiBCrpKJ0fScksWMxSo2rUtdIBv0plXHU8
GYn72TuFDFN3huUaxOf7knikNMc9orwKoFgZhq94GOFnMkq3/fzsa42bYTMOAR6szsdfXEnlnXRV
0Ve52qLKRCpIuqP1j1vKzJ1ljRnYmSEmh55/YtF4ubblDQ4saVN788SOb13LkQw8tiRJCA8LKzYL
sfUjbM+C/nK1Hn2CpFy9sdQAQV3mdvrlJiV3EkLxke0TRajz31tvZfsc0Ov13LlvdNtyaVNzVPqS
DEtSyGbR828TeSZ/6bMa4Fy076UTjJ06wf9rCehaAR/EFr6JG0iQHxviWuouD8RmP9A2T9+oTKv7
d+XkAYKPXdJqKUlAJj3t0VrBpOBni0JzqkDJKP9GUP0RV2jazaFRqGFVfcYMeUwBJN9ViNKHxMGq
ZzVw/w2wdbr8KsxxbXlwfrO5ixZvldPxA3bH2qJczXOQT+spf0UCxD0FZ28d+D63bpcz6nt1bReK
HQf/YDP5wjyCTjgGj4BozFqFOb3YiFciC3Gh/kUZ6O0kJFBlvve84kG3PLmOGubNo8blRUotteT/
qOUJBp26Af9dDhEVH1sqc3E0S0MZL17FiEbcxVQoYg6W1ad4mH0bpVxp0MAWe9f3T31UTmw9diga
qCIRZjBLr03AGZSAmZPD5sXDiXigTx69gHSTsQrWjEeIQ9jZRckFcnStNEs3fUl5bE2PSfSWrk5c
JMV04GZq1AvphaRAhB7RlpxbJFSiizTbwRgzqgz5U/a8iNTdE9/BXEdK0hOUX4nYLmkF156i4UHK
Vj1Vj7Y8kTYOLGv74F7H5ZgpP5WEyo3jjYNLJzujM3g5paZ5zmiM01ISdy2eUj+H94/CZ2e3Rlyc
iCWvZ4Mtfgp0wakP9+DH01kkW+TWfPbFG6z3n+O9fqA9Y/XWNmK48mYOZN34CZw5aOZaWxrkci6s
tJPxjn/u7PXzO/3Ov0zCKB6GSxiofBb08hZsFr9FIzW83Xk9ntXk/CLb+hlAF6283lRsGh7SFLnc
Exb7/PhxMYojYVYx0sJJry88aJfAkA3N1Lk3YvWmKFtgNx2Z5KW2wfNPy+YczwQdeY0fsdq2u1sO
CXHutGhE1J37BoA0VUXLomKHjv7QUON9fcPMZ5J6KXfw9t2w0rd+69bMGA65jafLx1rniTKFtYld
F/131o4o9c2oV7wowt2s49u07ywRiVtrq/ZKDMac4KdBthejqsTpuJnB4Z91mi7GdzjnLDjXSPZH
m2ITexUNr+fPSVQJSLK6WKW8byie9LORbgS8z2fwC0RFjlRle9uxXkuKvn5Aj3FTf3mrPggXiHL6
tUrnGlBnk2NZp9xw0Ls2yylUSzBRImkT3EKqskk1QrPp8KPiA8P0FmNAJtn8imh3sRVTncr90yHZ
4pTnsqh4oJvwQ+cplfcSu95ykBveOZ8bjserZljrnXPzl2YqTdgIzq9Ftuo21hdmYVmPlpFpcGlj
T3SOTxPwV48wEZetNxPg3/chYG8TLCKCKK3k6PuGzOtJTkoe/7boazc7H6tXgRQFMOrnwkVaQdDS
o4FYL1Wni4zlttN8duhaT2MIEXd5Yl9ENcr6SzLcHm1yT7rCK0b5aQr3q6dDHl2B35pDbapILWTd
EwtmZQgGGOMRWHSVo5zFpXMCdLkBV8Fgrupc3YJn24/XsqqQhsuHuV3hqAc+CtiL5QTJGF+TuzH8
98PurgsLD20hNIAyurqwuB8x+4JDMSU5gR1IrnXWvJ9pX9hlZevE/ok1+1jno+Dw0UlW2iN9pFgo
o1K6v2VqvaBcZP72r5w175i6eaSZzCnRl8W+7XaM+50kIlo6cDxG5bNhKBxVkOVFcI8cj3J8l1vr
A5pxvFXqDXXsIpi/qpVBXW/1jymZpx8ggPZzz1ji04Z+6XcBqjCUKpo+XPo6qOrdt8rcIhl3l8+/
sp//f/IlCC5yrw+wZPQB3sv1iPscOs0ZU06W87wB1YUfbehP+h+pRcmRYGcfv2w3gTMo7R6oeULQ
cDMw2FBBY4JreLlQ6uQ8hvwQiChsh3kGl1C9+ZNMsOy6A0D7JjBDmg9tLlTrGxW76o51mn6CGs4e
uSwSYArNVo6dZKAZkLH4Nb/5cK2Dw2e1ruaw0WF8LvOcS+771McNyRlFEnvem5zClL16CLbIjiEW
jjzpn+VMkK52VrbhzzBzsZXrwkxQ5AUfrXhab3GZBGTqzESncpAUTE8yHjOXN5jbD3WGS/36y8eK
o0/BnQiX4Yh9SwTrgVVErtt2eTN0SvIuFaYzq0BxzraY46l88+SXZuk0tgFUxsu1q8X0IzUzovGZ
qIVpG+A8HHlSSo0qOnYfBwUukHimN4QW/pY++sKe9yQF+dbmL3PmYzOgXJrekjwxQGhKEXXnu7Fs
e9AFNOr5o41TywQP+8ErDdTBuu7z1bJJJTy/U39/rKEsRoidB5LKJYzk49mW5cgqmlCARe4NMLJ2
l2fjy8Q870sBbKOIwOCLAIZ1ziZuWYp2YCy/6mCFKClawq04UDCG4JgF9JU7fM7wGlqo00Jlgqqo
6IG7T7U0qekBcxg4rMFkQ/UkGkaFA18j0rIZ4qvEOLlMMTp2oa86I0XfvMkgJWr4Q6xz/OQftT4z
lwlCnS1uexhTHPQpVh+DmWwXMk4c6WgvslBiATIWCsqHR0acc5+SniQaf/JjaUIlLR9KtC/Bnx/9
8E3HhELg2U1/GOt5PQWw8SIo+8uSyjSaS9X9SAjnHCcNQjQmlCP+lLJ8QPvvfzQoV9PpES13yDij
W0GQeG67k89HTQ7cIFRBWYRo6kdc1tzt5qD9BHhrvrHby4IVGzJYHkBIzF13nLvd86rEiNYciVuB
T1JLrO5LN3yEy22wExazceVpqyr6r9tw1yUBVp8ZNR24tNGBl4ymTQSq8dYxQ3ly70ueYmoUIa9g
fo06lUn4K6vxlKFeR7vxPYqE1H9db1zr7c7YlBDsB8xH6ej9wa1mnNh17AA74SckMpiFOO+GTl9l
uk5CHn9uMNZXfcIKXfRTI0F84kOrmYkxtnKN1fYal+PwGUUI0DYTsJENRMxaU3CLY5I2yFJmAVg7
XibU+4Wc1JN0sM84xHrZtzkl2nSio5wC8RCWdjZp4eFJSDhPnQ8QrvI54k4WX8yr3uL69OzLnEOw
+9d0B2V3I8hgCvTs8F5tyyDALQoKSV8PsPBjCJmXBMdzyZDwIaZyYdqbIJdGN32HIZHs4n77oP9k
80zjzpqfCtAkAoBQAZcHdnfy6kbOw2zI4Dq8+VOCLwYtAPKbZtki0Dn/3glxyMMgFsABWamF7YLZ
VMAbgtsKvSCAaT3U9enbJDKxLWfdoTWpb8JYObCVKDL/RQ/E4oOs2sd5f0x+Fb6KOPppBKmR8I8f
w8hTA+G5TtUcuq5x5Gobhu36/0Y2sMuh8MKdCXmtjjHXl0cGzL7qBwdzK9kEJG2CHHq4iJAo6xse
CfUyYW3KMIiaKNjRML+waa02LKWJlufDBw76wRaBEPBc1wwjaowcKHUCgX64KX8oFYlV/PkrItFj
puIAvHhJr5bLFIJAJvCou8Y7zuJniuPSeTRyH9Q5tpbY8M0ITOLeX2Hj+EkMi1lwRRdXPlE5Tsiz
TIoKbUTqVIRXk69ndJ5NybyXX2S2RlSHHVlof9wXZDVECOTVkhbOXRLM9HMDrXUz/c8wvWilX4Qc
E4MTRsYKXgXoTIdGAEqfrN6wSCBIC0hlDbkpICdnKWJXW72w9KPfbNstWyA74pC6n7Eh3R369vgb
G1vt+eK/0FahXaIobYFI9Jd/9C+OL0zvqTQuUa+OOx4j7izPUJ3LOSCnx9bcSi3ii2lHRO/6jh9V
hbnScyzfQowDKRt0SuW5NTSPJ1ksQ+j3RRKr8IKoh0/tpdBT6xqk69dHmGwMO1GIsJHm5C0ZtlwC
FGhCeTLlbrgJrD6O+8ZwelIaEEn5uwQbwa2S7WBxS0q0hs+UzUgGXY+HCKQM5/kTbMRKSYWE6vnK
kt1oY/ZtrFKuYDCj1w8kHBu2zjKVsklWBP6iqWF78R208fruk8lyVHkhulS/VboEFLrQEYW0K2HM
qWDJ+6oj3c4chAXJMxgC4o9Rm5AWqwxVaqSetYN1i5C2c4dUTiGB+HPGHHvKTJptkT43phr9F/g1
+l02y8alRiZLZo9xS6LrpeuTtzvFkJETqno/tcG9fDPPHV+l8JTbacW/OkeI/oDy37k0MUaUBjXd
fJiwWqV8KJzFBXgqeUHDcPF5aL0oWQgzJhUGOE5DXNvadCfUzjsgeNinqOEbN2JrcUriN9BG9ZkO
rUALdQQgeWFfTb6ZjOsx3HJrc+CGMS7UcMuYMurZ+1URS3go2yj1EnpSYgMA9tFhv8Z0FJusPs5z
H9kNrPqOwHzfbnctKoQFY0Zb9aJR+WIJMF0/+eLay3UnqlBH2FVN0kcCPRDRH0uEVVTq69azRwJp
AFZEstUI553wfdMTn8qovCKOIftedQEtb6p3nwuY23eGln2P5Zn5PWDyag9dtrOyXHqVgzn07ayR
3zhAMDTuX2OWpZsX1GU6pa8Q/TLelNzyTl698bFl73p+wUXGxuSZ1z+s0sDTTqG0+fGfkQ2gKkGQ
cQKr4uuiZhhi9oDHa3mi1IQxfUqK41EQynxtm58VIJngbI1bQALwZpT/avG+66lGtiRWL9ZVPo2W
0H3lMUxQZYXay4XQBmVOEotE8RBPYYDkNp8ruUMYfiaPT8aPI5jgOVwm4ND5Desp+3ewAsDISG6J
SMH7yB6zTOLseMofU6n7FSxF9O43dRLGmL0DUC7HC5OC7dmWT1bNTbSDNpasRJfC2RiLeQ0OzGuo
J8PeNx1gKsg7W6lnXOu0Iid2V/6xkBIZQYCy9iRDoYI7/3BiOIdDuKuW/ckVPt/IPM/8IMq71Sux
kY4ZK/uekzukLEYrB8t6lQLgct0FqpcZsrpwbR9CXeFJmBJy+YEQfdspUx+sGdFgg42fDoyWlkKQ
LA+PyklNoJ7hILqRhZXF5QilGoO4goZRG1KGypjJ6zUDGHUz5feL2GqtmrTG5F2427cfTJs+5rm4
5tEI55nSYhJYOpbXQHA+3KDM+lkCqzI2+KS472nDnrYPwsyiXzVZNSu+or7D2R1sP3LRbhFgB1r9
8ID9H+86u5gu3J0bUf1Uey/IUlspGGN8XlR7u+J2IV5KmOQ7l0ii3adLL+WwDBjKB5/bwFwTCj0E
V0sGCOCQgQOMHXyXnLcLlhJalJ5mjdaU3jFkPTrSDzqMFpVD5sPc9rQuRh1iywiaiNkDWRsQt4ps
NB0FIjNDv/dTaClYd2gSMz0NXG462V2r1FxMZsylKlWeK6ms1zSaLLrYuLNS+Wruw4vItibYlSfk
v49Z7v+lHV81uuqWu0oHdIoR4RMpI5se/a/DpVfdmSzRp5mp0SjrFek3fK5Pn73ATWBVIfnFw2l4
4aXE9C8zYKyyVNogLjZcIELt/kA9A+nEXLzJf5ORoyfRpx3Hme92iUdDcAxe3NPslNzVYWfy0AV6
Yth+lnpBH3ehSnZmZD5ovlEaQAQZrGHc7ZWbSQIm+r0JarGT5X3IGeA4XDIiRBM23oUC/sFWQnPn
GYk13QIwFv4FEeFBiIgPUYNrOSFCmThEoA6Ps5QDAcBo7Q6iKKL7SWPycl+LfKg1DTzZurfR/Gsy
Yld2PY8pfRd4Epx2oVo0kVrL58UQag4R1raQa2tSVyXX7/HwzOw9VEsPwy5PDGSrvSJsySBEaZI3
BXG+QjVrhGogboUKknusZbKAjXCqRC/xPtsz0wFdNIku7Eyp6+8O57yx9oxmYVmMi5U1kdf3o01d
eTOyGipMDWg6TrsTG+KVh5EC+Y8PY30EkPVn/2FoK2mmjiPL9aoGP1ukeLVbyyaUfhUqYcBAUGvU
ZSG+eahVIgyWhgwLEl/EWf9q3CVL2Ev20ryiBOlI1jEzxDfgtAwIoWEjYSH+k2W1VZIl5arbCc7+
x/oFca9rQKQD4hWjkVgI+RrS7q5UB5W3Q1HJR4WQ/bdXqzi5mqPm7UeFf2pBZznzX28KAv6u702o
ZOLgb7W7V3zI53A+Hzhm3maXnIwuS81JxucBXf+zoNpW8ot+ozaCwD068kAcYh3nt1ZG5+fIkTAg
Em01T3XlygvnXrXzGzH9v8Wf8dP87SjSScDxU5GRwhlUv5SAoeQjytY2TrjUG9LJ44SmdDa1QAa5
uesAj1dGUrmyuI2MaYDFlQsw+RQ9T4bj07d9EyjFUOM1m8cxtc6nP22DFTvRz14Be5/gipkVXTsj
M1K643GHNfX1RlVS+MNyMjsqCeiWQDZvnaoaMseKI/Kbkoz74KxToKrQrRxQbhDVsNoKzk4wrB7O
Cl8zzFST8+SPFNOAkzetJ/kgXRaEBpTBcti1zDaK/+gOzBp0tavEH39FvVmwpxovvSV37/EgrlBb
+BOxW8U0WKOARbzLn5853UhmKGcBmnrp2AH+vUwpBxPT0jYdWt+eiVHv3kG8LU2hkDcAOf4zh05l
NRseaxlxKmrB6yFhj8hPviNCm+dzGb6zBbxfrvD0LCPDO8BQ//nrzuzFIIZ70oJdl4I5v3wyUDaG
m9EjPQZIDesHJQ82ILnlPzVKOZgHgaHksXCmEpEC4kPvA+nEc0rmjCWAN3ko10jCtA8ef0mMi0rJ
ZpAAMmSn9g1wtoXzDIdcVxGAkpIaWTvLdtjxbCtGh6r0lNf3LfTsZNTTGVtqhlCuULcmMXgxqZDG
QlncQrc9xI+AzGPgW7vl3StCv7MyQX9xY0oDvAdQTh8nnTySLlBGa7moYHJoIUQgJHC8tTg+U5Pq
lIMXRUDt7g1NUCsVYHUKeRyCK7rl1OKG12Z4N0LDMMPc/RiiYKepDzftRMr+6wGaVnsvIxtMQN3R
ET8z177nMgc3t305zTOujqSyJ48aiRKLfh2PUbOZS6VpiBI0c0q6kDZ8HT4dZxUOEI3QNOfaEIFa
9Cc012Vjl+iyt0/EjJApyb3ur5l/l0Ru6dXIK1NgANZc7Q7UV8x1A+IJVhrxmOIABqDVtKEYXCKm
mA2jqskQPVRJSA1B2XOncRQi7i/JHX63DU3WgYA7XChSsKHjYrr2OeJEZCk+e8q8tFf0exA0XASX
chaP17QNmALnXi13x65ErkXFq8sK2ur/nfU13guNQC1h4vpruZNS3BFRZDHFtMnze5Ddovq8xSht
MrE4xN0e0D/7V696hx5FLHPrjGz9igEc+X3PJbs9RWfoRFxl2MtZugbFJUwqXxIc3M5LMDS1JyN1
yD+TVjUYOA95Nj7wfohKr7Q0T14EEYXh6yqohITuxkq8SZgkrjOJAla7fzRCF5yd5iqxuAbJSBlq
uJyp20tYJcGl7EXWqhAaRfaoGcLx2mkwGydNBHSHxwN1p1IJTH9oj3u5fBTpb0H5wcOjjX39F5pg
GMla6FK3RWzghj5x75aQvkIcRgyBWAkEyHr2KN8i2EmIUi4TsBkWrGM8xVrP5g+QN5uiWHoEn3bd
TIk7269BqCztNyemWZFMUBA5iNPbk+/kTL0f4+Ar+86J9Rvw46gutrrH2bpui+httr9XrS0SqKio
jU9HIsAmGP8ze7IehAMIXdFJxeYXXqNuPOTRgfGHOQEKmUYgfNjqK+hcZuUlLVcTmMjw8n039INs
UgY9x7WSkJbUiQhZOV/e7hCyb2Udo4/lTLOMW7mrKmb6YCP3WzDObBvzSbwNox9onti/tT6ma8gI
taGAkIEwVtTO/1VL9qDAsrgOUqp7Pkxw/fScYaFJb1qV2wlMUTo7aMLDY4pPH7eaoqnSy+o698F1
gnw/d+Sp/zod3QjbHnO2ImskvYKEol7auqTbOpJ/6ikNckf+WW6Y7l4mFNkpYva2vTdNl24/qUCl
wprhmZ1bnCaQBEB3QqlNmE6IIwOCBg+F6XtOasotYgU4W+x5vLzltqLYPhIk9PhbdzhNA8FJl6pC
Dq1t04fR+00/ntDMkv19qoV5e2hzJkhx/PWo0R+HlB4kdf53FS/jW8ODP7tZIKIPUkfnHjqAHiE+
/osU4V6pe6YrNYer0omrraXXA8U8zSqQDNKiWPRjbahuraW3a5jkoo18DJHMQ82zor3SuE1f/XH6
xU41TcZKd1M2/6WI4YUqy4nsUcMD16y4sz57L2noRSxD9hSO9DeRz2iKd2jRjeUhI98PZwbBRFWF
WhbO1POgOmPjqeQq1O/rtDTyaZUZshgGQLEc2DTKewEX6fvuvmPFCDRphhK0q3Bq6ZyHgzVMriAn
ar4CA0oeVgOwVsr6WlYCdBt6B4cLszmznn+vJ8Lmq38HawhwOZSMx6P3o+kcg/9wLyi/UQPsru3v
Qy7MCcjMMDpfAheWsV2yAvXhUY71pmrJMd3LhAIkzJCGhSmLsuKbjtjQTZsIcfOcaPXZ3hjr/pTz
AXG+cAqGhhh6Io2D6GL/VG7rysiquUaNmxcVCUJXv5nD7+PUBDv9IcQjm/og9vkLmB+2IlXIom6L
j2WjTcWm2lBAcD0fC2TQi+OCKn1tXldlnSoq9fO//43qzOamQWWq4MDdUI9WwfAkza55RNItSHb+
9YikhqxRGVUNf69+Ra7P2mBzvKIrEI0EwGeCAmsfAXkWLT9gkpE6qpMtPgcsoEfq9vwjoh0RfdS9
M2WV68ePKreHt2plweokL4J9JSoab254uPmP10mBWymEG/d767pzOJ+XgkUIhdaiwuUqCfFOv/Xf
DlFpu6VyJfHYzj+8x1AlRts0lsKRos+YEDWzuB6STLm+6cYNcJVfMzbbs5vLY9XOjR0gLW5s+/tU
zSJzlLNcvr8m9CiHyHr9m13X5OgJXBrnTpMbosCMZruDzPkn08QT4iGeWaVw6A+f68XvaFLVpxV+
8eDKL02gE2DWNVLVRyv9Su1JFFwuQAftXKq0+hzvB+FgZdE8iTh5AKHRWhXltczOC7gE3puz6uHq
gFWFNiP9PmLgJnE/l1M0RyrxD0/3rNXORVwzuQ+fFilwwRYcGgL7vKxVoXJDHpoIB2HNs3Uh1mou
BMONM8Qy1iysqu6m8Ub0MTqZCMB7B5SfdDCknvLW7AaBM/HRksuJsoT7GW5Cz/tf3wbEMjNDWBVh
xXVyfFuUERH4SWPEIErxb/wwaxBn5rpCxcgCi8Hy7pwldsIe+0zuu7M86Qc+VpHfvaEe3koJ+jSK
YZaBcwl4Ebc7zWXFpjmsfSCGH/aEv1HGGtGJIq6To/+Nb+v7ubHwhzOK5n6YTrnnOAjz6dZc/bpl
ZGFD+cq4HLQ7PRESO51Xk88831s7f4zMtYM4YAR7Xfgsut+Cg4ZUXlIurNtyE0Vy7MiMgbbRkOvr
+lfc/y0vxIWiZaMdfo9KpTNoXtfQpvZm6NXChO5WOmjgmMqgavHfwkeSwl3iN9QNRZj5JtxcFl/k
p9qDk5f0nQqMJFZ22HgUhNbxhEL7EA4DEhomHcYbz1UZ8Qe5GEZuKdsEcNimFUbzFMGulHonEhB1
/sSod7FFJcWAoWjkAqJ7oJikvgxdDhhHS5bqtTgFwEPN7yEQhIoFM1LaIRIAcVBEk192XW9sYiPs
qNegn0pwqFBVuW/Wtd0JXYs/eU9EIPHC2K5dOvAayi9AQAsAE5EkgOlcBiJuRGWDQGkzkmg20VWm
72yZcveS13pZVZ0BV9eJ8XfZ3oJ8M+95CSp8XooThcg5gIc/5ny7X8u6pFlzjpk32hj2EHJ56uzw
Rq+ebUvqIUHf05zGuOM6q9akE5ryXY3LpCap4aOMYyVJ2arsvHRqF2eGlP/MDJF1goXpxrm0KXUJ
AUfHwlRzRugqvhHpHSbz1PnfqisgoJyBuE6ByVzTwA3kHJMvRAd+FiiB2m9ug42iRnRNaB4a8ULW
NjoSH7Q35NXOn4oVmNAYg7pegSDqqtHQpinJHoM0Jk+wK6ygMpzJISUd2Xz1N8Iw+Ki5M3CsIBdy
whV7+ln/KkdQFC2BR+pKBN2j7oyY5mhz4ne5FceKjqRHSd8+fLEjtMaObmuXCiBwvB53PwSG02e2
ZXGRlj4J6YpxRgHa/LrTJyKDLykWndbeUgnumr8FrthIGYfmPo8/pUVKIYfyh0aZ5EB2dZSlDuqF
BSKdMG/ifQWmnstNcf7rlk0+hLiX9nPTEdNsWL6wmJ6QGC6slitWOflTULqR2WeEHl3dkCfoNl5F
sQkipdsX5TwSV06UheUxoRoWp4Gp715R1HJ1N4+rey93Bb3Uro+AzHjPGh0zHXdMXk/n2OjIADI0
2laNlbXmPFY18cOggpycdGDfqq6kmaR7Ksl7hWHdnUGXJxMJPfvPQ/qOP1kjqkXRavDBbBMtiNjm
Bm9GPwE370/vHlSCd01bYeAvWwSMUtZ7mBz++61dDhGYwPqt6XQc977NZIowgSW+mvMaM/JEfC5k
Y7fy1XoX6thx/q/luK2uC8ZfMBfYpcWsXAXG2chCccSHRTM6LruJdwfZHupVOGJQHVQD1y5nopKQ
1KfcJPmTVmWJBC9tpnOB6NXDqatiHnWwum3eqEFMQoKGY323umXt59pL2dz0MDo96paiSpmGM9We
cO22G4Y++cdmJyxpLIcHS/VqdiMFhMwdjqBYxJGrurmfM3/a8UbJYZ/FOF9StqPlHHHaK9hPJ/be
A6s7sCbfHVo9Er9lzR4DFJJAJcPWKdYwoeVyOXvJslawseMmfiFgxAr6djrYiOZlIt0hMumo8M48
OhieMe7q+amhqkB4/G//eh64aWF7ajPLOvum4A513/Wlnj/S1qDY8wVaXyMhyhhK2KSejsFo2/CB
uw/cvYVaZbq2xGBITyINdDISy6vYXK0vnLSP0DJTYt/pLNSfLAwJafX4a+DfGGpgS40ZTm9ogSaf
DDTjPldPnG40HBroc+BS14x4dCQDFhFVS2zjnfcNVRtH44kn/PYOkM/V9RafrJj9pE6RAk/mnNZw
aE6T5TmQK1xUTuN7b275KL66UoNWEjZYU7+iCn8h/An6K3zigGtsu9FYkLcSOhPZFVnFWoqbRtI6
PghkPc+UykapviYQdIYbN2sD3E76RpYQsYEnG4S+27JS9CUS/uKCWXuwelFD7r7ZV8iDOraYiEo1
oFidPREYbsmtsVjW0n/y6t+jxyjL8T8M+xSPIFKirZLkAPGcvydHSS4EdJvsYscntFQXycn3Fqio
geFP+/XYEwlO0XYG3zs1QwclFNIAFkff/fwh46KMWfeTaMcdebj/BMwJlzDSuMJRKDdZgBr2OomI
VU7V7ZWlfAskaM1KfSEx+c8cAxIfrCkOGgVh6WBZdRDioZt9qFsZ7SGMY6JsD+jJe1M0AzOZ+m0Y
zIMowAQ6iHWWj9zwRXaWnjiQWFC1Y41CDKTm4i3Mf7/MmkrWwLVpX67kXq6q7quqRNRb+J4q8d5q
2AlFR+VceEccVB8dRxjLzKF0zCQjeZ4as2lQ4/HeSHixxHKhO1GLPFzOmqPVbWiQ6h2A2Av5sJPp
0hB8uSHK/NpqErPO2gPw7eZRsdT+KGws6rVygTcEvt7Ghk1bzlNvK6p8Ky+N9tFCplVNtOs5QD4n
Awn7ebyNjotZFBgFRSsGDMkgb/A5UFWp8fg7hs1gQHz3RAypX9WHgPmqv9XN1gjf0haHOB17aaNB
yp3lco2VD8ceTvu2lqd9V3I9GlgDT016onGlS9MlSFrY3yNx8f9r/1CZVTpa5Nku/x1FYFOhvZ7Y
H1B3NM7tKyXKWaJmG70IgNEk7HK7Y1Iq5ljnVJfBUEB+X/NsL6ub4pzeSgAgqt2GRsiFTM8wlyiA
B78mnuQuBDVZoO74jeobP+HZQm4NjWhcLxo/4U1FZD7v0QMeZ4rwxnQexbIvz00kT2WJ38K869ZS
O9fHfc+OH8IQcv29+dFeGKe1yFK/ZSIArUSvWeW3P1qYhPUsxZayJSnCSj2oIFupFUIR2Gs8EOpr
UlaxND1wCLZnktdRedA7WRfdYHO68w3/JYXpuXimDIrH8LHEOOwJOLjpcK3U0hm6Ol3DCCPk2SFX
ndYNNYJnXjForSWYKeacQjoLj3FINi9dKcZXgBBDL3ztL28J5M+5f6o7i+HpEaqO4hsi+magai98
pRltdXE4k2uaopTTzO4RKRcSR6VtLBjP75o8gbqP1SobXRnwGDEllW5UPOvF0cwmKR+WhpzjHLI3
ghmNjV34C/dLaK+DKas1lMDFnNjxAujfyIv6xj4iLEVspnXmZEpOJVDw9xvtX9CTJOOF2oJGwzmb
I01Gjd0m9/exBreEAtzn6xRubSrkwuXTB57iKnVSXPFr6Y+ZIettHirnKN+NzuwIL5NeBv43a+uP
Awwct9DKoh2b8bQO/ahdAo+D7NLeXGpswhReOoG7ORcERiHJTwqjMbpAVYwocEQLVZoPRbsUD+mY
pWJ87BWbFsnapI7kgdCmx1kx5/znj5TOa1pzBIz47CCqKYIZmVuG9ms0Qi7ps5FEp2a+XubxP6cc
dEQJoZt6tfMJ1ELTDvI+l26Zyc02BEeiqHT3pF0arkQgeImi9bissNJlMGYKAzGd1ZIIQ2JaupA8
9qAjsi0iEVVDJZsixjxTHUTeCnc6gaTJ+NqLz9BgPSV9nc3sA0Wp825Gs2oqsM1QoDiBkcHtVEtZ
+4elWcOimvRv7M2Ov05gwwpqNqp1HzfRugu1CClS8AurkC1ehG2uvPePoT0YTg80VwdQf+TpT0Mm
qodHU4unfrbWbyOsgA2oHR0cgJh16uZj1Tg4/Xllau/ENbjyGpx8HmevhtCO8sl3ANZspPUHJpqw
qB20m7GoQ7wwoIovaMm+FXzz193TppdxcZ/hNdcH7Cu1sApN9sTK+uhyqq+EO5I6ZSOCCDJriUHb
I3f1GbZKJxhB5Lk6R5u995Es/OJhenyTU02yEhy8POwiPGlyXk9Yv11+mLM98rFXPyknRrnRWiSj
Z0L4lalz5SBWON7wUYkHmdzGDTPzX2iVBUegf/gGDESpCKUbPauTxip8gFq5OuwCXOwkUzCa3mwz
5ZKi3zYXONvwnQcjb+c7uDNgAbPs7/EzxoyqTicjFMPuDub7xhgInJHaVM1r/7R1r/Bd7ghh35Z8
yHSGB7dZB8xSLq96Se7vzYsbQZKZoZcYZKB3HLK71xXZY+253XGp2SLH1pehzHkHqgEd4S9irX9I
8CLmdrwyVA+Kf0OLfvly1m0vOFiJbw6qXvzDg7ySwMe+K192Ss3mdrXKpm0wPhCShuc5Vc1sCWrW
voP+NOYKjD+XC0W5VCsrRQ/l7vO7jaA6+3dzQvmjs3MDxRvGtzV2op1H7xJAh4qeTnT7B6xcxbKR
uT96corvUKTEBJ9dpjRk8FN88D3RuUTWc+FtH9oqWzaoJQKYJsw2eitF0BbP2I2KVQd2nOSrHUlw
kK9N6x6nS2CmIzDma10iEbvpHobDF1fu5XbaN564uQkVy7XfNx3fCpKqPNHL2/U8V+wXxEONLtTH
bYR2Hd+N5UbBgVufe7gVBf9+QC2kz59kQRVw8Z/6WK1MuJFyCmNIOnEombiMeQ928tR4b29qrmxU
70FKxiAgY/6+lpUQ268ihysgYvBl4q8Lg6rKhjL7+WXo3qUf+VAhukQdffGd4c401pgVYIGpuHd7
6WjZywVJXk0xFZqp7jOxNDRXlOrP0yhIXf3t7K6UwSrqFmtGOk0XIlZntAM/ZCWKWENovuINnU/M
p0liDp0oJXnV12ZJVH9fCnqMbQk2J6YZVGdt/+l8wv90I5/Sxr3fJtNqYBVUyfaxWv/yndDXMofQ
1DOF7Mxdd5WnBAFErvMTebzXdS/qwdoGxmM+T93A2ti8GAhaY7uK9ZMXmJwdaE0x5MNJKhDdeZ7t
d9UE0+v2EM66WoF47fhRnLjC05o6TUK7eMHFNAJ4ONo009lm2KwamFei/47vasN03CTnjehnVe1y
jZ8jAdndvCTNZtcSV7hCZtNPLBz8uPmnV5/EK8GdhlU+tS19a1oGQ3kMtH9FLmWJfLPCQzG5Q9my
FImm4ToZ9Z1fiLxJRXc49x7o2mRNeh05iBYLZNm+2td6um087cLSHhlFVp2TVyqxYV5Ok02/4JjX
0zE+NDEwjhIDXZHhiQVDof/vc7kl8bSu+iC0H7nkkXLMGdg6bGG7WtAlpY/TFBuvW6qLxR+OZUch
O+/VuVc0+1HX8Fuz+xXjcnJ8Q9ds2/Z/BxfwK+XNp7rFmSrdyjwUxzWX7gLj39+/3GLSPpCc7MZM
X/i4SAU9cnNEFC4yQtWZUNEMiItQHedYHx/HbjRN20Itc2iaOpqeweo+x4M5qgiGZVM9DgOx5aXT
yGOXAtXY9MyP09tJuKPrdMYwt5Px1T/hqFQpHWZVetUK/WNeDsmngKwiUrWE5PXavqUTk8DPyaZE
iT9n2dT0xn89PRyf6zVPoMBMOKdqiSJPDTNsICWSXAKOqGAkveXWfWh6oj6rBGJAWIpYn8ngxRGA
a1WG/J+nLwvDvR/4a7oE7kzePIu3GLTkFjlOuJpo0dh42akjo4hyjlFqa9yr+n+7Wz5YSoPz5Hid
pR+vCHlfk5OC6/XXyxLcwVTwpRFHIezKaqvVhOeofBNg8dVRMQRBw4VnYevqVTXWdrTkZzwbO0y3
uHQSlH6kt757qtR5SUyb5fTBPeC3GI7PtYqWetr5S7MyBz9m+2H4v7SZ9QJ1jjENH6UYvQf3v12h
Z2oB/XJJjRUHWtlAjpTzACP9IW5qKUt/0EwJY/3QL4FMSBWASpvYK9yXMZczpYwYkifY0MT5bkBT
Y1c5L4BYgmK7HkaasA0sO17CiebYvFJFtKpr3E0Z8S7UFaAjOKVrLwhZBTyw6YwNjGIe268aWZhE
MofJwVk9d9+SsjPAwnWmgLBncFeOZpq9RqgzZpl9aGQfgrRa8Pat0m09LrUqXIXeMjpk7gAw0vh2
2hokNLxwDbve5A4Ak2noD99dKCkLZ1CGY/ZTqmEVFbUbAaQW6FxWXVdpckSNHPhNJyOR2nbX7FDV
aj/WsoQUb34HwJ+DaEXmAzpI9vjjafyaFRw4W8ePX5/SiZHCZZdJU9raA2OQmJJhy7alhKKUtq97
vk8LW57g6dSff13h03Ta7vtDJ9sDCsJJ0yfZDONdUqSv4405bVyPcGX1R1escsW8b+1uw4Np3X1l
ESGZ7kR0H8K50bneujDUZYMp8ybFEJFDZcRDPDpHL23v8PSzisIFkqdLZcmHXtZtx0h1HuRMPXw6
wGvSytGezip36ppefI43KV5Le3hGO56GaVycL+jiRruXxf0czehxavFGh9Ltu8oNP/u6dBgX1XId
KGvoNBYCngWEHSmv4bIpqZhIo2XVnnSWLknG7JPBxcAa1jq+l1iRDw5p0DjCWUJgs1sK3ZA68Ugd
d6sNV8MWvpKbjYSlPZh7IDn8TF7eeXBaatArQFEilr2/pJE9BsiQh2cnLONUCYD711mJ1wN5spZt
mKQJKXaPkUMTUEYWWtLqsgLss/A8EhYWHSpKNCP9rPocfXmlOZUu9BDf4vqgtBM5kyXCGuZSkgNO
7FTjbRjLszeBuLpa2smpduN3hzNc7kR7gEHSZ7VFc65Y8oCGsCPg7ytqEf8OaBnZQGFrPndzXA00
2LuWxTR9+I8s9QQr7fdrRSTzdxa4Gn9iBDnKlai4p+m23xPpiYRrNt7/wdV0LTwuDimI0cNzwAYn
BP97G+gEoSwj5ERcusd0QEhDnXfYOn7TDKjw7Me4GB9wnBTCIYLratg4j+7i+ylbrpoQbo9cfH42
UZBrfeg8r/tkf7bBpHiEFw1iNRzLFzxHiKkTps46bM/1v5nm2HnoKZmLBusaThGlVJ4CKgCP5L7Z
AiRWAgiJ+YNFzC0KZw++8ugEDeA6sYUS2DNHJFxdV16eWdetxwn6iGWMvQvWXEyL3XdsvbiDC6Mo
U4W8GEKA5w+Hynxg75Wd1RzIKNzsA5b4HRFAdzq8NZY6TeMxzKlj6NqwV9sBKUKe8010sWic+lPI
e6Cil/n/DD7SUN6XG2aGf++qF5/GgxwQo2HqEr7tfBd2yLACLhSVveF5PUHnSCcO92rBhtA5Xy7V
iEXnvvRqFeEOBs1GaSt5/9RKLrbAfT4ZTIalBxdSLmlBIgqZKMDbw/Aqz9nVbZlasDfVvXqZZnYE
wdzhjKSISK1ho6WRuK14HUoVYXQUNui2cAQd880tjrvKSjV/NJGMFH4EmwaE/GrE9kjHYvXpoqbS
6Es37cbFMWNxiG52wTNeQAHVE5020tWQ4ueGS5x28XzWUMQXAl3NODNkuL4h2SOyWvp2xesCVk9A
saI3o3zK6s3ZxSUvfPY8n6ayy+L4JTJUh8xiRaHHjhwK9mdrpMss+8JZgVefeltLFfKwmiN7NaPK
oOaoRway1DOvE3oOtJj2yyMEK873FLx2nG0wNHYxT4BNphfefFB7S5aS0wGnFFPCcQ9x0HFczxVP
ErY6s+m70+mdaiCb2UsaSMVNA2R3ZZ958jVGU5ZkRYzqAjlFUwgjLwLUwPkqrmF0WBcsFpfMItcp
Zy95EQCdwmfT3zqS27dxUvgf8oiBFRab03O0OIEIpkT925enA/6w+8HE7dsz4pWpMi9j1SHnjg/Q
X1CS0pVu1db+vUG99OYzYxvnszt6zHDFwp49bXGCc8W4Lt6JA7fYYKprLXy2wEYaDF/v+QBcu5p/
iTsNQUYu7ktlWhTDjpK0iWCIamlHHSkHN+eknYwGdgV3VA7Ak22tMaVA0tzv2NA4+PMiizBmtaem
neA8yxjrY+xNY7mFMc+WvkaJhwYuEBSe4PvX9iLROFGlV4eJR1do4nD+Q4B6kmo0XtOkOfEIwc4S
svHPzEPMdniDI0yRKivt11zYRN51PG8iCzOZpof7Fh5QBi1VfslURNBoyYQU9qixcSZV/LmMYFJ0
ClN4IPKYZefMD1EL3L1jxd5yNv+o9bXo45ctmEh6abAFRQ9t2RDUVtu3iaC5d7ZLSQeW0c3wk3li
V2Fbu5E5uEV18lCUQ+5NEe9waO9ow+MDseLCC4h5QtbMELXZx0FvBtETf/CztEUo89zvmveKW6Pf
SHaXMjEUPWJvo68NZKRhZ67N0eGBz90xXb3fL8z1aGRV+2Oh/KTOvKlEEbp/mmMbzSZdIiczRR8K
0U8FZBDZiaYy1XpnqQ219l6KvX5lbD9ghcaUbIJvam0jZEtuoC8lamcfBfTUnpLPNBqVmS+o0HB7
s/EyhiTRZj+pg3EGDe61APDjeHntbCDCvgIYHhymaA6UHVh6M33l2aRxBkKO/nkG6PrGBgsLGjB7
IU1pZP54b8l5g0MFu6kvSKrEfxFugsd/up1SAKu2OlmCDVuXBYR5u1kvJU7kkWGUOxIiQNzY5pZY
l9YBSM4Id3PgfTBWKR6m4F/zkEK0RvFunahC6ojbo/mxLQVYYV21/zHYCFbm1A1JtL0ONznXLl0L
/EjrZ0vn2z0mllOzN1QM9InFvBe07V0ceKkbh+4KGCUPIJtE4PmzDnOynCP7R+ehROO/jYKgx2wv
smI482n9bXByJ9hQgrfrfkGb5+4ztuZhYSjOCibnpUA/XETelylJ6TGJAAVKlZxnZyazfPEAz0wj
vsLAm2D/OEMIu8ctHS4X+VxrG4Te9H2u8cLRcMGdhiZFB/SX5DYGkdN/WrlJ4QJGssmDpRBC+ZfK
fcQgxTUjaJzUpFLrT+6NaRoTzP+sP9bkdjEuWJ17iT7Rzg9oVeMKPTCx1jsoaEGN+mK1OSHL0p2c
E9sEntYW1CCTTFBSg2g2x1uG2R1vyhVjT8wIOa1tLNMW8nPUuLFdydmZKuPzsN6UfAUzr1D9ovJp
8G3JZmYkpcsbw2CWAm8q5LdRvQjcXVwrWwDWm4WToJu2+/8BjMKl8qi71RftiZvdn9KkvDKt8qXe
raL0QJlZ47RAsqb7l0o3X1sGVb0Wp255V2ovYoBE+uIJMRtkU4yBtghjJm9BRTgtOfrDWYWfWnGc
2V3Dp6yYpZ3ZXLNYrCtDo2uY2QvqenZst9dtRqA4fsv4XasT14zoPWlhJiYbaYqG9mLKKlbv/uMh
bK1xENFvLr3xDlpyYRekE77UYFu3tMPneL05jSSyas+lmHHCW3OlMZ2bA0je6DY6BfevcNQHp7GM
VWNV3EXUNSTkWgI7ooYNu+nJCE/oDsa637WmSZ/CsPeyX6/We3v0GDCcVlfmqixsewJsFPox95i7
J6JIL9HYUcI1KiyN5bmZz9EKRaHSJNCZi6Ilh2tiP1E+D3qjMzcBPSVvRlCN127eqoc6/DWt3ehh
4Gid9ec9VoCZkeDWBUrdxsL/IiPtAqyqh94+DfoDO+ZRxgmdJ0ktY3GBL6fxuAD0ViJ2RyJbTK+A
L0PFg3O4jvi0OfILfiXApG3RWRjn2x35SeHwGqC5lENTeNGZeZCRXTn2qY0YiqtxtOtBGAZigOtG
+MQrKtzdiuYkNaCrvLy4utl3S40ySIg1Eg2OuRFLdM/53I7dPkU91G0U+ktarZAAx/Hew+rOrsFv
O4jMZFbwJ0laS84D1dHXLiGZngTsyrV45g2ssELX+7qmub2fyH/s1nCg/Cid1NhUAQrURjNf2akD
9CH+2hinNKThDbsJzOZIqx2sXK87SPg75G3X2EsCA1uIkGtqj0n16lbXoLUUS+zIIsot9GYYV8oA
/vcLmj+DXOl4wqEMhB+07rwq+iqWOcAcQ01Qr1f8bQbVe7yF/JMhfKHsRNUytsHwpAeuK3jqHvrx
9cEQA9TI/RtWeamQVTn5Sqq0SGfYDsSZ+nXTh3I7nNHKlqvYuTMTwA6jAjtDrVSOd7oom9l4Y8co
7ZLcloeLFlpPXqYT+NjUAJBDzh62NT3MMOBiwHVnc6buTvcCfFPd0P3xmhpQ8yhv5oeCmaqoFcSu
9kcWYdcZcp2j3YopKDVzuDjZSvj+1hV04PpfoE0lcQYJI93/VRMFnn7c+PPSLKMLZIvlFGx4ZDMV
gAtZYD5dVoJkvWK8xqZMlYgAMEum3zUGPku53FyPBGf5zaa9d+xTSIZHv6z2iqIh9JcogckV5cHt
L9WSQI555exwRQslm3otRlTitjDbeN5E5Wn1tqkos7AdYOwFxOzmgNGuiC/siIPnRsj95VuEXYX2
BEnGYEJ7wc8ThSG15slPOYqhnNavgA14QEUSFeKHQHKfcfFhMp6qFErwG9Eg8+yhqPJJb9c2o775
p+EBbyYXk6LaBc+v43cNFUmoBZl60JsJUYHKk2m+LdKV6FUne6Mf9rBIvvuJIzpYOUrYhV1T+ByD
plczFRdGe5qFuNVgQjV7fR503qw/d12v8HKcUO0KYW+3e5PR+pL4HhOlA13ma6gr6rukTdeO2t7F
Njz5PRGLIDezsBNdTzifA1Oi3eMCu247zfesTjRiZAMUYryX5qa8s9evl9cs7dKvFIpouQPt+1w+
fOvyNG7wbp73TTT6cScozmtS/Tl15yMpF8PWBNA+bK//CSdnA/poTPbUBM8ZHx23nlJXxO0wO+RW
4iDvu7uSgygtxFH3J7xVup+mDWJLNOaDZFG21XQIaGsb/tKUgHLF+1QWfS18DPAIkNjncn61OceL
n+hdqrjMI+QQL2vG9ng8PmUobIJOt3SIcOKoFLYo8d9H7YlOlTKGqpGQwIS3xZIpIGvKnUtrtpXD
a/jBUtCrOfoeLUb3DhcZUIcrCNwKjOcr1nlV5nuiiDYVUqLMzo9VFS4fJRVE7JkKRUV7fLjrb185
C30lS/ivobS/ah/xLiwylUJY0CpMu0RzkS1S08gRxj8H51ihKGLWh2E+W09P3o27tb1CyxJwJ+ye
BfH4YMdlS7hzSoX21+wkGvzepBEAzjKMmMDjEEBVKHEkIP3pneghUwFUl5kb5Ac/4/vU9JAEbTA0
d2iK3OTBg0KZoB7tFinyQlFEWW7Ay2lSVrrlTFxp/AVwg5hZRqKstFvjaWdP7AZrvwr5/hjjLwOy
awHnj33YK5ycqhpYr0EooN3EfyIqy9+k+ytHJxIZN0pPvh2smjBsD/yiTKB3LLq7wBZtid7LbhR6
ZS7DteLGLZ0GIFfAKQTWEG68ky1Yzq4fgcefxqNp/V0hEn/ldTJMiwrnu5uQEYRo9WyB0Fg75iYd
uBjJbSfzBPaz91Q7gLKGqQCs2uSJbjPGQ3GoT2PHkZtnZZt91uD1ZCuye4fqYfsPAzIXLdPtOj0d
OMmbmqIjbz05P+mCnxHwSOEPks+6Xv5sldiJHk9MGqlZndZbvsQerqNKGl3/cn5VAP+PZr9Bovgs
0m1LFt0ljSXcjzB/6Ctjo+ugK/KbYHxVjqFhRNScyG5FjII/0jmOL9Ikrf25jOq1MgoDoa+d7oPF
ypdP7lgvzwrAUoKsnTaCECGPtUdq0KrMPJiRInSuDFpwRjtVcqDBPlqCNzVD4AFZPR0Ld4yedkRL
kPsQ984ktEoLstWHPjtWhxomqaXLIQH2cV2nfOYZX4VMHAcDfmjdXkxrSZZayQj1RxD+a1JBSvQE
JHXgwSWZDs7e5zUtBRxdZ6GmDITDWJslp7ywft/PABsjzSxkQ5VTguzI0wab8R/4XIAtxP3xFLaz
cugasLU1mQS2p8CPNEfmNoW/uE5QtQMwrhVVJXmmNGv5VRg88lnC/N3ZMgLXjtA0UjOeDYa3wQQS
1mh0Mjc//h7vKVMigzMYEfL4Oi7EHjTpUO9JsIR+yzxSSZYr8CSULN1YIk+KEmpDqpLN4y4/iPZc
1b7u4jKEzhqJNObBzOJ9QHVm08FwMojP6l0YHnCsH7zSBaypALh/E2X/O/hzRbSUglyklQ4Rtit/
WOg4wbfRAtaco7FRl5F7Iraw3S3BXVTCgWyBbg16fuvqnjj/yRV0MB4lAh30YUvIor31RRPPS2US
9wmNoEQTNu+fxW9VN54rl4mWQ9UQIvUvSIkiUcXkTx9xgWvHhjROMwvjuS/dRg930sCm7r2zPmot
4oKEvcWoH39DEZVyK54YAvyTEfk7EFYCHBbX/ozSEXCAocfvMOdV1tWL+giTPqyZI9gSu9bs4ZKU
WiUSu1omJVPNWlPU4tdQmRtdMyPPulDB5uMGdvFlkZf4+1qRGliEq4O24+e7bgtQgtpp99pPK8jH
krMGI9frN+LsZmBX7+Du4l8iegSiL9zOvyCwoxg2b6cCtJsWe3qPgIV+1WZ4Xs3AHgl8MoqfwyGe
Id78s/6fFCaQ2GS2tpaWy28ennMJhodBIY5D0Bge/eMsbgacssFF95hxVgfW1EYmlxmW1zMnEXBm
c+h1RnkjcnLy/QWCV3etaTg7NMd5Ukk47BkBz45x4Cw5Ss8kudc9JLRUMSfzm7xtWplMJmlblP82
ziymn6kMQLOgiQrkSCbSRqAOv0P/LE1fwGXhRsnCj9ZYECjqkMyVL7JF3lbxserrGT96nnBGI1E+
5MUHe/UrWY7LCmYKcJR1pF0HEwCEcsLRSIaCe92qU3MlucVA/WP2nlsHdkByAS2cc8OX8G/1Bn2g
41pO/PVwgL77HHZzG64rufZMB/cAFcFg6m0oilXO8Lw1jMsUOWVbZg6sQB7awPCL42BZ/kHZ5TDx
pN/eGXM8GVL7NFvtd6rtcwzMbb7Bou8UrWgfwwg0gHdZXyu6Ot4vTasERHjdVIGSOnAoyq8OSDay
f8M87AokKEXLIug1JmUT9WGOmKjCq2jLih4WLgNJ7/Bd4prD0vnmTQSiVJw8edmZzwUiiLMpT+Bp
ze6bQbgTJ4OAgcqLTffyN3TwbX2i8A1119DFhiSDUyM1kkbhJby6f+uHuZ7TQLoB2h5L2ND3iQY3
Tqfedi9dS4y7Ur4jqf63JzquYqVHpRN/9WPavH74au3FE+xvEUuJfgINf/Mb5j05dYfwIu/UZ8CX
lxA6o5ZcEF67eD4BP5p5FUFqwUmjoHuFwCu3oYd7aduPoLPrOSyMF3elbwowdIkTStyx/D/BfU+E
QlMypClHc8X+j2fqDLvgXuQVur9JrCLiw5Z1hFnuS3pYiZjFJGiQu2Mwip2JrLolqD+stAIGtnRk
lohFPM7fWhIM7HhnesbrlUW2Fj7by1xzz9wxG0OLrzjZr7319T3DlBripB/78tViL7hpRzZc3BIm
NytciiIsAXx2+CfSOY9UQFNncaBuXc7MLqr4vNOav1aqlSDcU0KHIA5obdtBslHKsPMxYsSRNx5W
6YUU+4bLFOjn8icIyuCWyXfHSRAeEQfqNgygrR5jWRzOm8ft8kwISQuipTSPMO/5gXZQqp6FhRYy
vRVeg7yXIwV0s8cuPAsftHkVhlDFssEEGgAXzhsf/4dy/cpxPdGncVymAzlfdLXWZxud+hZjshhN
gj4ZgtWJo+SimQN9ehZJSHjXFsdPLtrQEz3L6r2bCVQGpTGjTr11AwK5dS9VBYLrpf8j5x2+kjny
C4sjw3bd1Df9pmEuW7qjpJVVYCuIzULTL4NXmVWAsBcqaNxD4EUjD9vMSlzA9LMy6wFMuqwv+oZE
SkB505I4m+7R5WAQGjHltG8QlEgs0bC3kfstQ3NeJkUAVBDHfMIA2f1uSbO0SNzJTr5hws9P+pzT
VVMv8Stryg2lZ+sOxnthz1uyOXF8dPQrrFmJd4m6pc3Bge9EMKVlveeIEFyGn9g1fGCJxsFZYzEp
bkR8ruJ/rd+IoPSdF9yI/fqqC0e3w2FM9fhVUC/HXFIJYg4OUEKY2Vc+wXo4pHRXq7XfacXzl2jp
ztPeRxcvAy+9fXKriHM7Q1kBMpdbbXvJoojPjrZ7A5frReqNvFs0bblazoQ82Q4a8ntj0ZfRNUOs
DRunMphP5b/MAMWHznapPtZSyuj2UizJVvv0aa4E4RVGJspkv1bYoSknz5ZTLrf0avLRIb7q6LDD
gdFzQybIPOeJWSNigtbie4DDkOv6L5irwL0Y0vjw8se+Djc18WWJQgym4OvLFt9KvQ86QKuyyMWN
zWXXxf1vx/7qD/aYe8RRDi82G0XynIaJx7VcPouBBzmZc3t+iWUNqYULaoSSUrI+IFrZBMlZG877
Rj6KYpdy3Qm0+d4JDb4MlskwCWLd32XNhwKroB2XydEHYfRHd/80i2/dpzkvY8LT//LP5/gff1+R
3O0M1CBGDXir0tYIm997oRtAM/+zLs+6kQyc/Wr6mZ4mdlSYNoV2/eqtwRC7HrsVZKDaaCF9cQv8
SH2E4nPq1IVTNhAi8CvRfxeKoIACyaa17W+f+yNvmL3JwMuO8ZsBvljzGpMB0KuysAhgX9WOZLXn
27ThN91veP4pcwcisGNn+sXRufzoJbiXkz6BfY1g3gCkqkVMgipZV8t/88/TshT9gbtC4wUZ2FQ9
hsp5586FxcJ/nfz8DjN5hNppuOOlrWbPrN2vGKb/i7fWBU2MDLppIQZZvolZNr7sgrLqxw2t8mSl
9d7yMV65S1S3HYuRp908DBnI8PIJMetDv1djnIiYXT7tQ+0sV+mqZ/TOPhjKcwfZTcFYngA0o4QQ
+r71dPI6cBZKE5VIInaf5E7FrJFy3EX0IKTrfs3Ve2OGR1LJkAyJQp54IHCoLljl4iQfW190EAyP
6SENk55fREsTCkfbOr61xTmoT9B6SAoV4VqaURrZynKA0iUH6IKt/VuB+km1yagQLEbFD4MaNemF
eO0jWmskVjS3uXP3ZBuYX2JTjjc2oT6DbqxuIV3Ol499+tmwqNuERreGMQziefW3slalD01nrN1p
atu3HhbrUrPj+/a5p4j44Cssr+a7T+3NE9d7UjZJb9tPltLlp2Nac2FHEWiLcZu+utCjGwKMVPx2
lw1oQPuXzyI+mmuEHGFIS0kQbHcbuzGRlsmVhZlVk9HopfQBD+ZJf42O28n91Kmmjuoa4XK/jEQI
y6/L1pp+PpPk/RsWUiOluciFVT9Wolpdgo49F+YqjREhmMjmhRdN2Lri4JC/g8nxwW+PQMc2Lz5/
dsC1JuUAywRP3PUm6jwVN/BUrT7AK9uZCDkJPPwFtHuk7OxAjlWhlb5pTs8E4U6Yi2r1Ciebe+D2
Gpg6689gjK4fkHDYKP55j2HzIN6D2Kjb6p6nENwROA3x4pSRXGh2PnZLo8NwQXQqOQPCEMHdutJh
EDtrqCOi/BoV5J75g1bMMENLsS5Gc66J2kmWxR+XHNpf743yIaEllmNBnAcsEJt/MFOX/k7xnWWP
/5N4/pQBGgb3GedBb+s+OKqUS2DWlhpopUtea7PWkYsBsecgPuWLYff6pWvMJ4v78Y6TifBFJf4p
QHo5uDfq8VK9fBRmDL1ywcNYfYs404ercjpEoHKFqu6U6BFmUx/3F4aMiUZnsBmV+a6yULFEm7Hw
Whek0NVRF+Fcn0jvz+ec+6cwa4i1ZUnlXZiebVlw7Y5CK9hFxTcFX/RBlIyNPdEpcLi2KHWfsBhq
2lC8/ghdrgX557gzg9rgCBXPreQVpAkPzCXcZFU7vCW5/ZrO0xU0TejvpPgUHCBBInUDRC5APxHM
3Ymjs6eiNuQxvvCPVRd/oq5LX9f1/LSba+IX1czx9TRZghHEV6WflNLfCbWaU4i6EA4O4rORXiiJ
Q/N3Hrtk9pdu5DOAXMvR7FGYAPb6pWba17rh04bzObKMdH6O9vdQnASwekg4+PknAP5Blaow1KbL
gk+rCOlvHijsZqlO9DD7rC+G6xsnLddMiJsvobUgMVxMlWks2Dnp/CYAOjQ6Fa1XQFLHitKWgJvG
E/5yhe29BlCvpvh45cHqAVZlFkpn4v9KN0oqauISwk5OO0Nl81aFk+JT+AZWzCxX4o+h8u5b95iY
6iWI7aHjwK4sK7jqzThzeQ6IJ0V7cW4307O9gcLTxUzA72FmtJ5fcc9oRE0smZRff8yQOb3FFpfb
c6AfKHRl4aZ6uCT/gmtRbxmw63/+i3BGCk13sD7XDOxmUrYlcDMaDCH8o5pWA+AaFX8ge5T0ZeF8
wMjZkgl/qeEtzFjwkwcJqcIJMPUmTyNQmtyqRmHDJzVo/POKtyJcHt9FkOeMRDpgeOOpZQ6BFkuy
GgNcwB1PHzdhE4oZFg0rvRxFLRrSOMPF6Z0tV9qzZB0/TvtPPXRqdxlbnnK7ZWk2aMxDRQfUd4oA
AUsVVeZ02E1+PWPpLtJKmQblN4H68AnL8CGmvexkhV9+rrPF8BiWUT01OhBxe7yw9pgd2OEBWpXU
VrzJz/jjpNnVklf1eHJOTuFF2W/cU5ABTC/X76MDfqbyexYyMyFeRvZkyXBGKYLU4Cic1iRaVt+n
no+c1NpbsBkZEyntTSXhPZxDH08wcnAG1PdBRgVk/gTx5sAii28UNsg6X70/PKWBSzPcB7hsbK0k
rsVs2ubd/e9Cyayf3/EWeaJkxlYqn+vzVAWq1TZfaHstO3NtBST9FatusUtQtFQ6XNYWe9oH9oCA
OUA1Mkc4wNztsAKavOUVFM9o/QsNG3uWP10jtdYS8oK76rvfIxDDMIuT9RsAzN3BlksO7UZkHaU8
CyxJSKkuBFQCk1Y7mkRi4EFHdwhdVK7LAdEHpAobUAHVz+BDydb8lHfAZRUff9YajhNkPr5rAatE
ZDBFxNn6jg6ZpxQESWrA7US/BUCI2A9r/isgkEMZzHnbPQSoB0TvlydASSczMTVPaG247NnNfhYw
IuoHHW3pZGGHC+5C835bnGvaciKoaQAIN+k/I5BTZFKL5bbLI0BdezJlzl6fnJrHh/rZJ/kbOcfr
6k94NXqPp3/osyn7ZFQH+OxUeCBgc0sckGh6RZXhf8ixA2lye/3YeeJCUmz23OM5z5IvIEZ97RDT
5ki6g2spUskZ2M4XmxxjeVQ/Cq9X2ukirD5IR3Rc60yjtQme2NR/eQjy30dAZ+9TsjUbvgn8RY9z
+39bohMBo4ppzo1cyMNM24Pb7y37tPxWMXPFaYRaL4u65prar6ALkqH95PdoE/qV8lKSEJ/V7w42
aHhqTYEULJt60jANE/V6DyeQu9ByF0cOkdcyVf7Rr1bjfJa3P4zGA2DRrMjp/osGdaIlngLSRVlV
u23XiESA0ZfmNtYfolkmqkoprNP/1QQxakJ9fqhxylejMB/tMWSRE84fsePWJicG0d3+iKooCrWY
3VAfdVsdMBuaOHwTbTQ0tTFbltzv/ktCTw4q43oTpuvXuITwHsB2OJd9yKPe8iO8SOwvvhl4G6sR
GPXGeYhWzLoajJheUx+t0EQ4jsxU5ovAPm1IqJk5pMnbIAM2NvumMajLzldCav669n/rzez8zHVY
AqyY5nmYsHxZijT+sp4m3aDi9cWCgCIQkImbvTALRcbYgCZKIbyDkDbkhiKx/HR2ZMZyxXr/4uS9
XHd1N10CdLwYEAZjp+D7IIHx3byQkwNlYWLpsrpen67R14blyhCSGemI6BnvOO6fZJ7ipRMJ/WfP
qMFs1v9oy/JUukzEdvbOXxRItX7KdgBcwcDPedepZ+z/gv19ZBe9XQTBLf3Mkk/rKawVMHcm38Si
qq7BceKIXEqEjUoLSTVrbTTwMvde9icKSJ0LjbsHZPUq67rxtk1O9PUxdUWM+Oqjr+bbOPQJIKdV
wNzqIADHNFUV2ikiw4qUddMQ6ZS+ANf2QUqI9vOl7qJetHBWACTPH587b5UmYbL2MajITUQNZrlr
BU9BfYxK1fgxiVFRZGGv64Pw+qIXQk8EW0NHBBKrL/xBIerrKpht6Yo6WTMaxkifLUhkqxrmqyHq
AwEdQLvvG0mRUhZz6KVDLqogBejcdasTLAbs3BtxcD3H5ToJf4Z1iB0pC+gbRCjseISxcGjV4/OQ
F7/qPAa2lGYv4FTohrgsRdEwGceaNRGYu6bS67pPgATIHGx/QKxu80rQA46bznCWdaqYO9wjEB5m
saTMtyEuh7Ftkb8jB6tVfvCWmObnF8h9ayGxaGsgFON8ps8pehULyQFb9VlmSlO8iYQlggzaFPqo
gQYhrqsDGcp3T1Qtj0+gvPcOrp7U7Jb0extJE+iJIpavOBGzh3yMbAmSYc9RXZXttV7xxRB8EvSx
JL7PCRdbqeSzjlffaHMuH0HPAm9MuR6WUfmi3fMdz71F1s7OFyjlNLMecAjg4mGu5qJU0w9rlO6T
XOhhcNmNM+TCWkSoQNd0g845cD2ZcgEmgaTA2Xo2DmbKgzET57hIsJkSHq8M2s3EZvpX2HTRgP7W
Si4B6dFoFiIjQutXYJ/lB/kFK0U0bjj27Mx4Zj9O87jMk4zDtEg3FFx7qeZzjFxIGDiKR72B6rA0
mk4BM4PApYm7h59+dF8idXAZ2GIBvP2risOAabm3shdzHXZWUwBD/sVkGS3PVQhUiQyOUGccOhPi
E9/VdUvtaS+6ovilDyUVxMbZWoGxrVPse19mnT/9kqzrNBQUlPis0JnuBPbeMJ0DSFftZ/OSQ4/m
RsljeSdZhuVFkGj6It2DyoNHS8x6yEuT0fUe8knF27rSmFwLMd9nwjpAXojbc16vtDZb7k6L59YN
0ERfyfWF4yZxYfeG0d22PRB3g/yunU3R4j7pf0nHelsbNV88YbcdQvoE9aSOrMPULozTNg2n0tt3
viCcBnmKTuZE/dDMFbALoVUiMC27U8zNvw+VuZKKO+s8iCEeQQpG4bAv9JhEjJQpnL4jN7jwlRwg
aCUZvDRXLhnG03SqmWQcesxJ1zU852NUlVXG1ezkRfuS6m+lhJsEpcC6sDg00CpsVUlKgtbz4Y85
hWIEVoNHL72y3P2vsPiEwDx3yTs9en4MZDwJbqShg06nqHKDPjX5F6RcHjHw/yVjJWTWDdXQH1zi
0ATdWb42f7fPPcOw7GH5vS61QnF7RgCtW5lIefQukMJFB+Bu4XEGqCbYFDcH0U6ToOpM6b009gxV
xYIL0X8wdynMSdgG+9gyNsqf1+uM1qE7Dkg7DqtP1QqO5sXgCl/Q0FduLdlp1ZcRHNk/TzBVMcYF
nFQqQ97Dlobxb7MykIwH5ocd641IDFg0ONM05pFJK0LU0jdj2byAzhHXFPPVmmUuH2oj+blINDLw
w6rmiueXFKGE2iV+DTmVR6zCx2rr6zuoKEr7U3fygsMcpYkHsay8CatJvGu23ecPK4/jks2Rp2Ui
8ssQoVToYn1GEqza6zhbaWImyjKk17Go7d0tJg+Tox9k2TewrxAK3fM+NdIotRjJRhmCjaHol9+Y
5UuQ09ZB5juhnqG4YhItfcYpVT89+Jap6IUVMFkrWaY28urnp8C2xmhjzvuXcNIsrlC3dA7p/qNQ
+0v89SftjseIcHLeZPkc8Jl3N6VbCUwaj3p+sL4ZGDqJGLnYflHJkVNKtXruAsgZhgC0b9xMulDY
lVzSgVtdFVRwo/qHcNtB8k58Jrw3VNXXDYsnits52WowtuMtLspPu/Shf10mPePKyVqfcELc5qnO
oTQAao9Xc1Yc1VwX9NLTQds6cvVJ1hpqN0AXH4dMCsREb33yk66+D2BAtgwFX6Wi5V8C22bYG1Wk
/2V8NAbWvBoJGcRmFq+7mwcUuC3g+gKOQsdt0ho79ykJlUXF2A/FNJvZKjULGDbwEjeIn5AtsnBN
z3jBY7pzMI1ZxiMkmnNo3giGVqE2k8D8QyW2oxMz0nzuSO7nhvCMk95ED+UgSgRW0BQCRE1vT45U
k+IBtsfvN4kS8reiRoqySJpj+Dy26VYrPwdq/EWgGfu43eHyvALG0+FILqjNhUYg+47gFO/nGEgN
vFS5QpANIBgV0k1z3aHEyi6oCIur/3H9bj8E5/aN++G579DB5ibbNK2WsCa/okkLzEY2RFNvDCHk
/d7e+7cH6Ax/nlwGX6ujTXviG+KSxhtHrdxTNKM97dTB5ofTDlGaKbxCAhUDqwrMTk1fdhRcgnQ4
3AwPGYYBe6ptZVKeNtpxLv55TAK0QhVdkQNtblnXu9WgRxJCmwFPgaqrV6MyIj8YWJ8/1qS6pR9j
UA7uk1l3bt46wMgm+rybtn2kckGLS9xz3U0UmtGhJiOi9V6ProkNtTbKX/zt34WEC7uX3S+Rew7P
ijhwwHi02JOPMCKfjE6j85UyLioU4j9igxVr6Wj/WtsDQGtD+Qteej6a/gziI5VXUNF86AIZLkJG
dMlrQbrBwfkWY0o9GJnB29D8uszx/+iGkw6/UGZCkDDTcF4CBvWJ7/0fse1TZYGelICub168Xl/h
h96w69gSASAbiLhbpe7FHKEWXGpzOtN8fJd+SWO5SY3Tq3oN+XfcM9iswk5OsPruuiM/yYb/dlKN
+JDbsDPsLXA7EbyJ4X+m37zZbNmu3SMtdlZMYNFo3NhIiGba0IHtNEd09t2cshA+qFZue+AcvYJF
Z69/uJhJFu4iuu82X6t719Mz0jh3T03GHapYAbtKZkkYdpgzUeCKHFPWCiqZd8NlF6loE6tDUfNg
naZ89DZs8duE6ABEMRhK1GOaNmQxURRx4fV/bw+UhbZEfkhHLd9buIv7EU3XbKX2S8UjD1EYfSG+
cLgjVN7orh70DthN0nZ0FXPpTOBC9h10jp3txx58/kAxdksvOBTfjeLzs4KrpX5eQnUCkJMafabY
jiWF1rR0dt1roGT9X+hehzJFjZ85ZyEscve7Bkad411ympTQz1JvO/IB+hokdmhFnqqX9TDZoAic
Q2u8CMFWY2GomK2fSkxMKmWBWkcDg5XnrPVVzTQ6YY4a2n8wtemGrK4HQRURlaZbvAPEKYVtzF38
fOQvFfTRW9EbhimTmBXXM8h1onuPqJeV+tbkzePb2bkR9weASU/r7Ae500zvNNWTD3ofUy/g1TCZ
LaZP7yb9xCS48MacYmf5mD+8lkhZnBc+hjyQtAlSRsos+JPED/lE75+TdO55p/Jm7UHJzf/mDl88
vLFdg3b+f9kDYVYwbegpIu7x71dpf4Emu0NNYqVXagn32+cIeGnasofvBy4wC7XeeZu4bh5alXCm
/EhZKxlyiEY0eNN4vRZtoU/SjoU7LabcMVQ7Gzmq6uQTK33pZUBOj9YEY83uTMf/JmxSDFOM1I3z
YYQS0XHvyQoML9QZLyqwxWCFlTkv6pUvfa/sHogauqHbHAAbvCDUH4fDjhOVjGZo9aB59wGGp4uJ
Yf+4sbEj6B4dt6jKr2DZLWjQ0JI2uXUrdl1jXwjWhG2MBalntU2A/W9pYVb4AXx5AUja0nWjpnmo
zT2rYRG6fzgIH/IBLFuj8vL9VVqhdfWJsZSmlsP7csm+eBVfT6LV18eI569KjyACyi+zOq5cHWVQ
HnRfQ22WPvx3cQxI7dAkDF24/+gon76jupMY4u/9bROzFHoHicnZRA1GLFOaumKeNYj78NkJSMkz
xB8RT0O9UdRSBaA8S4YvMIMXXjgjGzjovN9jrMQajSQRhyu6d/7i/ZVOZb+obKf88ZNzdeSDJXhL
6gAdpTtMuQDyJI0LuzMi+azcrjVuSvcFCRFbdTPSl8qTnC7vPAtFptSF7AVlstOMgUq1XIkTXf0D
ct4P3U/wzi3Khn+AQCT4NUZli2dn/7cz7bVG4wRj8jeIRQk8OVFsxG+r+Hjg95cJS4vCn7+vay06
ccuHV3yR0Rq5gYDdmLerK1x/Xzz0u5qIeTd/KCaQ2JbykTNWJEkTeGyDY50la8XJNRTRqsgbjf7x
dAaa8bOLg9U0K1DG+DEvP5ovbug47Qpz7dRDB9O1gl54y+/qqRpfVUX0SObbVmOoZCq8pB2EkyxA
0JYGSB4BOmDHaG8wzyV22SW9wMKlsx32Hg710RyEoI2Wk6Qwbe6b5cD7ZM+3ElsJrOwtY1tFWNRR
Orjnxt8ZB/SJxDpDNX4ln1+kf3Qff6nET5oR1qc2+PZsV5Js2QUqJtNBt5VD9iYYXkCeyz+e1VrA
Cf3mP4JPxEyjrHCiJVb4KbhyaL/S5RRy2a+6PWzTWIDfR9KwYkDLK7qBkyUZqGCRII/e8XsoqxIc
mO1s+OBEpXwwa9Tjj4x0AAMwD75KlK5Rv8nFejLg0WjjHzKTPOdbDJGGnkCx9t5MQjImpuuAjhXj
CiiLdkH/7qBD+h2UKOG0GAl6OB0ABlyh6ViXaLL0fcy37bsv0ctC8yhPdFAMOEJ6F7uWczJ4USsM
AjFhlcT2WRTqmx+b3y1poyJcoyAiPjfNMfJJlp3uzrmO8XgNHq9wihTrqHDB4NlPCI2EY+TX3Ho4
e2m77J62zz6IFcUUa6+4Ze1EkP9ZaOES/ZO6Z/Cys9LbXsCpcyqUTCW8yQpPqzK8PLhjq6xuCcxF
fQKgHtPEhOhIc+ZbSj0iQwGBMo8KbMOi8wlUSbXxgTu7Jd+xXV6bBZhm8eT+r3Rp/6PE28NYnP6b
iKT5uXho6G7SwOCqZ91BPR+KSVsY9TY1u1mRihzenTMiHzWuuX9ukod35wSbzll/ILXDCtKPzUT+
cJ2ogFtLCW+Dm5tjCk7MPrdPJOf2Ez16LN21aNp2iOF1WGLWnVsOAoYv5NeFItum2uRCtM1Y2C+H
kDwfizCIGDEMB5Vc4OxRx14qtRRxAygswSa9cGnCFa9WaUtZ6Yi6jaOKN8ncCjKgyT3bVTfz2Os8
ooQHG42Mj0wnWRPqo0KqEQ9LBnGAfgV5ImC67p3UORH2aVTLoGLFfX2mtT2oc/POhJmgBADFkOi/
I5Y8uspfCVMwVSihX5z4PYl+Fkvykbpw3S7tmAssoGW15qVKHHf+oPBncwuZWfmM2CBArPiKkNFJ
/bfQKdKxJ7TmLam12RLIorGR3AlXcTZdPX5fhM0ls2tYEeUotafeAW1Dw185eHWVGf3XLll3/O+5
YNvX1I/y3nifIuxWTC4IWEWDvRH4Oi4bXHQEEbnmKKlPBAEr2O51fqYOXXo9BAtiudOq5ZBBgVk7
y+kuQdE8zOaG3kqAh5zmYPgXHIiA2/VpCZ7qbb9qEU3cP5AuPBV9uf/IdKK/HpQ1SZWtbZzS++Qg
Ktz+YUvGfJWAfcehAkMFspAKceaCyBH8TmBGqXKi7J8AuryrTeVIB5GDWaBi3qky9c8fnTmGvmAX
JX1A4I5g9COG3y5NZbA0Zr531bP5oTOfYhxariwKXOA2FDFP43tzrsfcPSIdOsvhWKMsMixxKQjV
YpqAoXCVAjGRCHLS3sckV14FGYjUF0vqAluO0exVjySkdPfbl+A26U1wv6fAYLvblWc6F5cvILjg
DErESChtN7qmRyJgzUU+yBGvgqlQZS+ZL7V6vZjCNx2I/VEokyR5sEv+zZShQHRL9Zgtg43/yJ+y
PvsmKRKpKQvqT0mCvFLxZVtFbT8Oxy54pUpgXhaGAqQ2w+pBFW6m/BPclw3b57bofOMW8V37XRsY
uzHoy+iV7gU1CIZU6G6RxUaIZlLzvWWP2C1ZTFsmH3Uqq1n6+ubMsSXbcKyJf6IC6ugm4WbtcibL
rHIkoFNVAc+L++NYwGyBALgmqEOy8QqATFBMfNSbQYq247SN1iSQbR3WzqRTmrN6hQAwwSOk6k1i
yc1H3IuqPhXtt0j75Gb1h7xYtgLFY3/a+685lPE7KdQbL6zOM1Ais2heslY+pn0X+G6td/+yHpYQ
Jk1hB1US+IUVOEhoXKFaHQ/LeWbDEKrbGPe2uJdjWc4orLdcQo1pvVWTPH4Ip6lMxncUDshXjRqw
ejGdB3l7FJmF6Fx7qC2lXIT4TBrdJpezbI96sukJcOhXAKxiYvitv9gOypCa/jXfv15HKWXGBerq
eIJinu4mbCeAC5z/Dlp/IwnFZvRHC4WO/Ebecp3dWPkJ7XruMMcdZlBcIlbJamvtHuvDImFXYIDb
KrM7vfdnnlXrnrp6W7x4vdJw/2cR6NZzgLdgFlNa5oTPYk5Jsjkn6UUzxxnWDJGaBAfPiISxM3tB
xA4e+tAGyZhc5ab7yutnZqclgQjQPI3rHG3qD6ALpwr9MS9lQxMyJqk92bSFeWiE5cIgknpuPphO
ff8AWHYAxHtzpZIYFpNWwUnuridZnbDnivkmhpL2+BrDfiivMYDd3EWv/H68PrfxNcTtI3gyHh9A
6hwarDXs8b2xW9Rwh/Ry3wlSVXBOWM1qz7cwc8CMcQy37v/eamAKn4rJ5mtnyg6BL5av/sLSSlZD
JfWkYCjZe5J3Ag3d1v0Awtckw6ixVtgTU1afrD3qpw6t66K2T5R9WXgzR62d1oWV+GQt5HVBqySk
sqxzTFygSN/lpOipFq7J3vPv5A1PP7sbyFbhNU3POiYQOFhMF4w9bBSca/MRM4h+hjsF/A0W8yHB
GukR+99myZmFwleWFfdbZSmBGxMG5RBBFnKFE6OUdDfG8wimYfUThBWXzmASyZO2zcmEb0s++2qZ
goPtsnKO5Obdiw0Rv8JyqzQ96vK4Th15FROlKQRIBVBCKbV7n2xkgdXtVYX7YidX3Ie0Mm4MWoey
JkIIJgQGxz5W1psAb8bnsaC6l2NXvkuyNDbVClegabZ92yQX2eia22vn/xYYGpaH8Y4cK98D5mCB
3P8lWleTgngkQJP0fIqSRw8KXGoLUhcuP5YAiulEIB4rTuMMIREA4LfJj7qLMabnEWUBoalGRcXR
UOaZK/TsjDS/pL4TJ4a/WekqojARzQ0KSbX9ANay3q7On9Sw6oa391YP5N9pTzZ/D2k/OAt5QiQb
ji41JOxcjL77Uj/a7Abwg5EXJygHUME8OFvF36IpHyK9IsCwDNFK+au62Q+s6Is17hyzc3w8WR6l
8prIrMLyhFWeIrp7K4hMz9z17SgV392kXvb8cPvZudMzOsGm8OVb52cIzSJAhhRWGqaddhQujMsz
+ieDhD5wjuBOg38qj4/4+a5513/Umy50HlqjlitHFg0QPbFUwR90furJ0uzVp4OA2F81es7LchIN
vX2egJSPkRl60+zldxxSAlCQlozGTVM95rMO+1UETzSNyNWCECAZUf8nH7iVjPQqVqvMJ8zS0/pa
+C0roL+BjS9XKusLDANWa5WpocZ61JMRXXX1YZUVOlvZonC73Nx5q+olk1Sn7/DLZW1E+4Ekms9R
E0SHvED/s8mwK3FHMXIFiZlkjU3sPDAmuD/rEH4zM32jEQr6xz7s4HOaefD3O3j6BoO9r3guKAcu
Hds01XaH0YkrJN22NjEome+3WBzHxU4ACCURUkDeV3nD4LM46GOkKb9CUUMpWIMI77MmxkicyVZ0
WJONepr22Xnv98rH/mBd/FjvmbYjUg1I3c/zderG7GGnXad1d8o3Xe8f92IyZ82fR7gY/A63U3G8
EBVoZm86r5/FSYArpm1sGiAbRS/lgRoiujSOrCWoO270c2gLcpq73XshFcz87On4TzaKsP4rKIlt
LBc1yLghwZw7Sd7keO9A4Tf8kBsWFx2LKSuYrzFOeebByAhSiN5VTP5CBHL+ovGcqtY9V9P/uYxp
sKIZz74C+lB7E79Yk5qmV3EPlw7mzH0/d/uUj78p2sZH2FkMHmqSKDtz/p71hmLg9zP/T6VL8jM8
SXL1kcgdfA60kmR5wBSCRSeu0TMjpHwxjvgPyUKaTO+ECiDbyq4s61OfhUS0wBx62tG6yQlpSw4X
v2zvqHVgbSjSSPQmuPM+TifhJ8Y0c0XULKHf8xbkXg4/96X+C5itc7/Csw3uAQu+fitnRPfUvalV
y210qCgy/NNkwyr41DrDZ/NWeQybNgcE6a3AxqKA+kFBZN/uMAj1Hq7a/imuaI691vxsWccF3ZqD
qocAdnBuFd8UvHd3VnNHQ0KpEGvKJLn6jm9FxVr9I/wR4YpPHfET4pnR6/UD2mRqWQyPVA3GKqXZ
QeY+RMjsAI7btOMk0G0tUGL090pB8lp2gCbdAAnW48wHF2Azqhccdw420Tjmcln3WlBk9KkR7uIm
U1E+C1iQsidWx9kO2v7vxwQnTkPPHUIeJoks3U2lzvp3XnMgNhW9CkrJIm0P8NRl44SmR01es3r+
L9/wGGODCSp5hzP6c2qzB5qiDwiE6L+VMfVnV44dc8qAvl7PqOuWOddIcrmZfIFgXmq38XE3Qctn
b7gwjJ4EU9Hhzd+KKGSlhSsESMlF9PGTf7cLT0OrOGCDmMZ0L/EmQ4+ZjrMWMH7oVa+d3YLQjKF3
P9Pcch7fc6/P4kbKdJm9rv/HpcLnXU9OK4DGXBKsRhD936YioLZR3+c+U+9SzyVjE8lCQ99At6fy
cG4sSvdOfka3Yyxj5To25iY7MqQlaWwj2hiIOBKjUZ3V1h0vxjOGG3iof1TMo9M11s4P21pVd12/
F2PmYidylRUUhR3frMW0h3kTEpNhAC5nx4SX67OLNeJw04F/lLVHoArrqmFwyee4DMdx4olrKenh
gNxTgoWdOeMQJBoMDXoYCcgdYIxws8rRDdctOfgrRRJ8MTFbk2cOqt01QTTSBkBw64jd6o6bVQiC
e5P/6FGat9VuTmDleRfoAjAH2TA2MlmQD+v3SdaAu62nGo2glLAMyCO4Mg5UzCRuOCSlHBFmk7CL
ufB6xiHG+0VNe8AqkU/6x1DZF1R4oJ1b4ltWQFfeZF05qvS3YN//0bE4QVYpuRQKAbiWLkmYPjtx
VBcCT72x30QHro2ndVCfyOd0oysqpCQKigcII5mCIkQ5K8b75Bbqg8LYaPAezaNLCdpLYq5Uzlg8
Hw0mwEbouOJzPQ9ZjK0pb8xJ+qCgNJnpYdtLbMswaRcdtnZ8Ap83aWUiA+h/N8q5e7tqW/mEjRf9
GD8Y0DT6MCho6DAeYGKMX19M+xlR781p8kenF2e9JxIt6hpAN6qhMN9IzZJIyXxqneMbkdhqLiRB
81NVgtMIyIwnafHrMqRaFdQw6Jyjwfrm35FhtlW/NSrJ2yCSc8o9DKR90Nz0PPkgTtgAmboanaCm
D1oHeQWKXuFQMEyDECYI42vvo5HI0qGZgZvD8533Wjj4ea6fV4cKWSIX29141e5VbDWFwgPTYlEB
ObJ/6Peu/XE4RJZ7n9pk3S8UHSQUXHB6c/x+PiJnKimzmXWATPM6Ijab2wvA2zjbXkM8+TWgHs6+
/uP3rrsMrI55/1DWrsBM8gGnrWCHQTkko6MYJXpLbMUh5XkphcuLl02QoMVBOBJJAiMnLUIY5vK3
iJHhJBAl/IrdxZpOx0LWqSJESbrfmXjG65tE9iPRMpFYodB7Um/qYsuMvCJlXYrqsQiUTV7lYDpx
NlG4lssITESJ1jowQyJDtDBkoe2nLlFkU0VWn9Wh4AoWGkw7u22ygRgGi/rJWX4W/DmJI2/oeAyn
/f8GNblDhSULFGxTUbRn90VJyuMd0U9oZuEVE9lHcv8O+9i0jN7U8J4fJ+MG9nJk/w3bt5IlBgIP
VmdoIDfBwz9mRCcHRO2OPXfjVAX4BNE8kvgSw4UP8alMQkg7qKdYwmGe7sUzKCqHmrsfPuKG5t48
meQOT8fAPfJHnkvbJE+xuDs1szDV2x3HBEw5W2R4TDps6gjFriMS/792z2Opm1lhxZHTL09ajoIT
7QjVUav9x3HSsKA6Ygux8cgENfh2B0WYt/IWneitCRVlpVjDN9O2NSAiDlhUNRdgyg50JM9affCP
p4TREn6iC5zTpROIAkKBXYGseIvRBkz3ASD38FJ7MN4X4ComwyV1OAeOaCt9wpPaI5S0zNT398pq
dWjr6iE/0CVsZftjyifJ1i23JsNPS+efcmdh67z2/1iQPrkGSabSIgxJ8xl0KT+eQA8gcoQnj00Z
XGGiW+1sS9fHQwFcPgjWO3f38Xxhu/O6cgWBx5DOv+XdOoQVN5PNmd22P5uwGG/PDl+zpuOkEIIQ
TnWC8qLeCHFQliGy99DE3he5ikUPTXgYQpNfJ7kyYoYZuPOGhF4k0GNyPH6mHn9mk/tSo6UP248J
LK/vYP17jgdjbSUmd2Sf2w4Vt4SiYLVu3BwPD/gasc5yrKc1BhPciV9V9AVd5HSgwLcotZiv/cbj
kmpMxGK0jNMcRvh5Os4AoH6tNSUlpQ1efiSj0DnKaVFxis2chOks/LxDciNs+HTumaX2fC+AX09f
ERKBuswaeYopn5IBY/rzJ0GkpGXfC2/E2/LvTsAzNzRD7kXs2wjUQhL8oJLq+Gyl5M5Os5LJmUGj
rAGRC5WRPx66FdB5GgwvKaDQbTF7vMRyGGGM0pilXWu9SvToudGumnEGtr0iWUN4svc8f+mpt4OB
B2L5YaDgSRsEzGk3F7x1dSG1PfqyeHNecPTBQFdGGcBmf34YVnsHmqZi5J8q9xLMwg5Jv1egQP7a
BSYlLG7mX2QJNX8mC4ylt3uzMYoinzL5A8aYF8xI07RRhnEZfQ/eLighQOR7tUtZsd2PdGCxghi8
Q/C/NQsAiGFeGXYgj6uOWMmyTsU4/NxQAvEmCdirv40NxagzdT/otpISEldQN16nNjK0wQF7a0zN
uY+QLWDDQoeK2LAwwrdNF4ZhVyOAz8cRbUmkm9QsonzCo1dHWCT19XBPDunKcVLmjufSnmCqdmSt
OnunhyWrguGdVUm5T0NW0s2JkxTqodRk5lsmka++9SU7AMh2I4LPp1Y+SzabwVtxHeWGFvVts8Vc
uB9aNVPyX460uwy7PP4LbL0i/0lRw9IpF0p5bOfPnjV6aQ3JC6dzTRyuyq0Cu+n04/BYhcPRhweT
p+hz5tgcndF0laaZHp3Q3kS5DZhQ9K2+aXeSh5QiySHSe0MrEtk4FdviLiv4fTT4otSU2E8zkqvv
EjptGLvBp491GS8h+vJtfsc2GypeXpLBH4wygv8F7SiMiw4PQxSSfJG7WNvrj7OjJM5hSNdNXawe
RA/L3FJz1DIP+Q3qOW7h5nkeeUK3w10TLj3s00bkWp6cpOd4H48PRR0tSS+TLsneDD3Z8Ef59dxA
U0++BrlegEFCAaVSoJf2B7OnArctrHUAErrUztiGP68jIh2HwFg7hPGsYvbi1exQHohq96o1kqoQ
BMMbTMdYwEGTffsT2tslchX5xAZPJegQjN4po+V8c2ThkSXGV7G/1e4V+3bV6Vp621DLNRoq+U4g
rd5/Q235n8ealf/GiQWlTXFpkmYYgQaK9GPs51pq2DJM41zMeT9m2YkaSxeeMxRqpa+tyMIUjj58
keQZrmKXmoxoTprc70AAW4MPl34JbXeZo1snzKEZb09fpuAKYTfZZrphQyYG+LROVW86Goi4oxGf
Pu/tsOeKdlS14rbLeF2TE7A0MQSLyx7anX1IDfyeg3qY/YBy6ObmpTt4UFvcb4TPN1f6MFFOto0+
prNtY7+tq0NfRWSKKyWT0qEETNMVDVPBEcGSU9ApMFbRvkP8DqHTFCk1fDnWYjrXQV2+ixhL/Hhq
d1b6yTVRKROdK9jxrb02UWxTV98Y11Q3UMNoDfiO6Z9g6bajUZ7fydRUSAUHWkozvMudHNzkhv/G
a5NGWQiUZSv2itqbEzDMm/MHzz22CwKS4aayIoyAaOURd2XMaMRM7is4jnIJYf+Olur2RySzhTcy
MZ6Cc3SKIbl7SSOEnwHPH/yIodkGNJ1/5+rwOoj6dJQsEQtrn7CDZ6IhnW10sB/nCY4LrENJYvN2
kB0Y6mPB/UAjuq+QT0s2eD0ZzEIJZyZ07obLhaEO34O6I1RdlFH8yYeYiAOO6ZM30vW0AInHjrNG
5DaSladyX1YSLMqqu9fXmJCJNOdqpSKL7IRIIeFhbWCOZXgYF9VZsf3PR35B6RndoAgutvrCrnKa
16PmTNRcwK/faeXTsGnDXXnV1xgTHA8O3xkouB3fJp7POZNTF4akMsQSV3Xa0LpFCgBOZvT5qxge
6oS5dsWw2sFwiIt3NtPYMTtA9Bf66IYULmG2eDC/hFKLbVbNP75rCyJpITb5EvgC4Ym8aWbz7/RI
azHNT/6u1ikj2CNgbzKSjVBjduT/LorG/N0GBVH0Cg9xKxzWrR5DGoBiphu2DMu9+iqDj+iqVZwb
OZZUkn66iBCi6SA1EgQ+DZBU+Pcqe3og6sBe1ojUHTLUVyD8YOHhC9KeFQXwLkDiMr8OvPz7EpQA
OQ7Ug8kapheMTUFmVpoh3amBw5dP6Ch/z9ZNqtB9c2IqRvIBHczsG0TlMJxZnMA2aKgVj7dGjr5H
c1RKppFgXurqilvObImEry/dutNy9yewzLIeWcExyG6bM1h9AoDSuYzGSZ1MI4yznuzCy/dBv/Sp
4hvtORrXCJkowGuDLNM668lr6ehA2YbZazyfVFhhM/Qia91MEX/wbQlJ16KqRCeEw4ar8Ki6vA4Z
jnq7w3aKqL4C8uj9sSOvZxwkWSdY4Y0h8hUXbjgtPWlulMcEPAo9bRBywVuIi0WR/1fKGpLX+2ed
ZSe1KIgmKcQYZPUuND3cJ3Rsdi7zvU/tZ+mJflmNecB8mGSTmhfaWkWKLxqg7TQ1h0iVnMr7aZCD
b8cQ3d2ycmkOXbMNhPTrwIefB9mnec2ZVPu+LtCh/hfOz3RK1gy43JrFWIl53orCGo8U44H3+Slm
anj/EFdheT9joygFiOU0ZICsycgeF8Up1VZhwTPAa9kGeuP+uDQVbVUt0BOiCtxxFjyxax0XTefO
8SPmntNOt+jmrUm6E36ALqD5DaSXLJYm05npzCjaEl42NEt+kBRoRSJDZC1yS4R9caRyLCikGj92
Cz29i3dw7C6AbwyOr7/pyTXjYV/sQBXirfqyoHuKxVLEnbei5PQRt8dQTZahqoRb5GvT/6w0G0FR
gV0osdyxbk2R4T7uLi1OsbIhppHAcwd9pqquTbwbfBRMJE7MNJ/Q9LGQdWyQAilCIZdvWLtR8Y4C
HQh68eB6Hv/BvjkdWjFlmCjh6SZ2ndUDKxs3rIqU8zu5e1HUCdY1Fc91JgiC5Gy39HwTK0Ekkf4e
U7nJi+3rW2nIDieM1pBf9VLsPFCEip4KqQx5uveT4fzeuKL+sVe9oUgPwCE0isbxo475JtIkT8Y9
6mh3UyTWLHk/QDWKdw5jRucSXc4/TV1jOp2dFDj/5CI2rREV/Uv1lI3Pz1obmbUV370A69W+E6eo
GlqUPcpwle3Gb4UXMuHWipv/+Q9lDrTAruUntoVxR42KVOlnMDmaRbDsWLrvPd/+dx9ZV2RCKb/S
QaAXXKauWKvGcHz4KH8Krr9667LtbGIX7j2Ixv1Gmg303+siodV/cBzkAmXX/w+qquyYboeVVd01
yyuf1SmRqWRY5S1sE9PpjnONdSXhYdhEdmzAWZmNRGZrI2jo2WlNSLSY/91XDGVj13KN1dD8/nYM
Xkq7S8nU7NuTgKi/3RfZFEs1JZ96gk/ofyZlRPuwahMWSOLLvbaGF69e3PJMzg2wFQbdNNcA5wT+
vQKNfv5oyEiHLRAs48K/aOIgbqRQaym6dBJs2Ibujte3jQrG9g2Sv8YBg4lHKbjYi9rQ0RZqskYK
2oV01huVbeP7P7PRH24vuL5c/znIzZ4/FxvPp+VRqqjOTDcsSHFsnTje/MKSmeWIg46JsITNQx31
FLDs97FPBkn5d1LMNEHtMJjl/W64pDNHy6pZdryARWpHksmQNZ0cKno/cu1LQ2L3t3sEdHdiR8VJ
pMLofU1KRSS+r9qom5LmobZ8/CQAKoQtC23202lI93RDJhJdHAQZfXOx0lqA1eYPZJQmSSmx3PEm
jGuZGhHdM26MjM8fgWyOqt82+ZXPqwUqp3Mf7A4lv+tmYU5FZgsjVxcUuSKscy7NvflgQhJYt4oH
/fbfvFFC0qXj4Kt6rWhpzsjDzkPykM0DPgJYoNMwYTlbcqgLX8e8P+hpCRVc3aDcJ9o8HC44sFYL
/N4YOqJ1hyB0xGdzgajbG0G3iYhNAWCBvYvDZHSQB3YAv3T9QPJ980+ZXvNJpcEJFalqPhi2pVzK
cc+BXgCCCOFApRfZPef7F5DbdjR+pZGdg2ubhUHN6ApEtQaP0brRFc9kqgLe6Jz7Njr9Yh7Idep+
oeRlaf7lsDu/Y7HwFgvNzF+igUE6FDsMt5XGDWUSjIZV0BlfYV/P89z7oiEAOy2Khl5XPdZk5s0p
ak4TZ2JcRELbWwmz75zr6EY60+tmRFroSDLosB2Jpnu0slPJa5qXTfz9Zx0eMBmASS3QTPv6Or/N
TredoNjhLD3P9wQ+ljsE2DDs0TTffauyY7CDoTn6O6Bqil45bkrYfRyh3oXFfx8Ez7DWBBwKdmRj
UZtJ2/wP0b3tneQ9nLsv/RQHztw8EMWlWkxAeVdR/uLy9JAdz8j7ZFwjoPdPMB8wNmqZ9wCBYbcw
tU8J1sXOkTLh3OoaTqFHXBHujpfFUzaqa4ejXrSx7r/WQOw/Zenuzax1Loks3Q3IFl2MD+SwDcmD
hTrYjzHlCC1b0HDiKkD7qpL42pGJ3LbFn6uX7wSifK9neeBR3vl8hJGRd+kMb3KSdXYTFVnMzojU
pPf8iAm6bwXDyy9x2I7e6g/Yswd5B6rZQELqy0y/WP4gd7oicrVfITD1gGXBrIr2r/PruQl0Dl4S
BHfuU9eZPtygRKbCSZ9B6+X5VSRlYrQFtpVvrB/OYRTuaLAyx2m5rH16CbqIGVR5HXbfUFXTBKHt
OYLWjZ4AEkpk3MEILgJ00SSMp3sKAekFdWjlUjVU++GnAGahEkv+MERbf6Q12FGhWKxwCEdUJxSW
byT+sLstgLfdgGugCtQ2lzexl3GsGCnr7jhI2pUEZUM5yNEG657/aJJe5cD707c75WVqS07xWihc
K8VMxsdnfXBznWO0rUGjySA3toL035vdAHfHN7u0cLrNxM4nmTZYBXkpvwfl/4HKi/P6y7shXEvf
IYPd3YmpzfoHB7H6YyVCucDaJW3XxUAPnssAfCYXzEGcQh1hinZtS+nJwglq3FcIsPy11sAGxTW4
+XRQpnMBqqkmrquFo5CZXV4FeuUf7oU895ky0O/6RE3LHuSixpGjD4MbOhFFrv9WQC1brNZqADqy
YfguFpIJ9F7cFSWnSA5szdikfCRaBob20vs/i0B7pJS8GwI+TaYh70yXCQN+N/K6sXMYJwUZMlt9
QpO0DLPR/eT+vQq6gqRlfE0S0ja79SS302R0SaxhI09VLIYHxRt7t6dAx2lAmVia4vcfcwVb9HL2
GVJ462kreCf3jFamUPIQoRVq1akGuFVAGugjj3E7wznvsQSf8MazuTOsmsKjIyrEAsGZ0g3kLZd3
fHXcuVfbwqqiu9Bh9ZuFnu9M42xwZVPbePHN+no6ePvF7nVUHX0KoFusBAAo/Ag9S0U0M42L1FHd
OUK73cCQhQ6p1jHqt6Mz3aD3QFy7JY/MyX73mXu30jSzwDjFzwxBe972sq2BTHnrCgjoWnasvQ9n
CF+AhjbBTdhJI6zoPO/7TDKp6GEs5tN7inzhWVBGCF8m0PTrvAwaxIvapljIG8GqItg7Zy+hiWjo
fhJUpXJ0iavK13eDqaX6K9dbWuyiTlfEtL9SnCi0Z3e04A5wNjiLOwiwBh9V6vddTSDpbQ2F/0SZ
I0WZ5U7LeCW5c8ed8KKN66x/uTj8QbXcOBViu78IvYLna8khXWZv4NvZ0Uk3NCY2WdlKGAwmFnYW
43C6VrNwec0rz+xnsurvD2t6kjdFo4TEvPVjyM341JKgtjDS/h9l2z6AYb1TkX97WedxluzzAIP7
l3tBR5sQ94YdBrvGN5BiBIntCcolWzgYiBhWA2myv/C/RLfhabwzhNJv6GxFFmUq5ACGLVI4sP94
dKjtvhE+aC9dt5D488wAXyeGCe+tySPTyi1TDBXNBim1Buw/0VXCVD2pN4RAj81KSZ/0+5fwkr9w
fMWKHr9ydMmeZUWkF9g3y/dXyMGVBq177eCvd/0YPk/Ovti5Dkto3r1RrSIzVwdyPhtWhq7GjoOj
HsM1AhwwIGl4aQGqooekv0fK8ydVEy+mf0to7HpChZIFSL+Cm2mhdL968ybR5fTqMKFI3JikVv/M
s38ofwZEuKSRuTZTBckcAbocIl/LvLun0L0yEgGdIMm08X/pvti8YgsyUYh2EeklWp1pj6ae81Qn
NjlLP6sbnMZ0xR4LHKxVICI/fbfvMP78h2PE9gwYaZGzFUEpwJsCIVpdIbK+8RHnEqZbX0X6Wyr9
7glDvHwAv+oJMzlGKa6jr+Xcdu6tHA0xMRDldE2LGXh4FpVUfSmDj0EY9Pif4iV1mHkByoSjunUY
K3zomQF9rHY+C8vAdoEkDKpP1Dp/yGPf9+ozJZTosWxiLG5TSsjAa6NnBgI4TPi3g4TDvM98Jk0i
4X974520kSa/SFVD0y9sauH2bhECGLFdkdk8nFKaP76B3B/HUv5Kjip/0ZT+Rx6XXM05uuXmH6bW
3sJblEn3Vxtm7PGou8GMhy0K+LoqZhPqBSMmVb55kTATyXgH6Nx/bIVLwwvkwlLvAMQc1Fcc+/7f
NbYd5OXmoZy5yL6UWQ==
`protect end_protected
