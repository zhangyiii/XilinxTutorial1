`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAC8BA+RJzsxIB/XPsWvwRe6IaRZ7YciaN+XdlX2GshrZrqzFW0XlcSYU
2rQIu2iv72F8+NhvISgO8SfAakaGjf9nNzNptiJjxJ8byEW94MTciuzcYlWn88lqJ6lE97ioMNcT
xsj4rWhHtSwLQ4WedJvucaPKTkbe2q4nNXy38N0lAyApMzlFBBiyzfBbB6o4ZtgGFyXjDWfuyvCW
y30gLaQM7BDLCpHF2z2rwGcXF6Q+Eiinf0wOMftNC9VPosgajqTKA/3SQTaZzAt3K312ysScwByw
OJnqzYO5oB8RlhhoGUctmtscdG/kmEQI8MekFcH0HM+0noqZ/ZfdKBZ7Z68jYyqZTzdV7IpdeDCi
yRRlvDrX1qo7o17o4EFx7itx+pWXo2X/TA0dhf1UdbEVOr4giWDzHbwWfymLjFtuWgJ5D9Ebdtgo
+RKEcPyzgU7lPgOfMTempxb51U2FJRVghjE4iIkkS0C/ovsBehtH5d+hrcOBJQ8D4PXaqUS6iiiP
OisDrkqZnAgN722bBISI26LoX76WGS3kqY6yYXuzsXhNAHvqzFvlU5CXSGsj7NQWTNSMBVOhzYqg
DrRrTRzc/ajrERQTzaUHCQ8vA3kVIrRoaPg2IOiH8wiWErAH5YMzS38enL+pE9/sfxXErOeuZbyO
YmUX3fzfQu0a4k+VGRu5kQgqn995HpweCesY2fSQrEM+uxrjdkqK2EQ5lm1KWPWI3ArzKESA85o9
yGlTIATGgL2U65uvbqOa8dDW/tXivMLqAM6nSdgVUvijg7GV4bWK+Fk3Py6kESCjpxq72JOjajHI
2zA6ud0OKyU6AcB9CTBPAHNfcBq5MwB/36E5RI+La/qvyU2f8XtDbkVRvUTXBuxlUS4Zk/6Q2TiM
mF7LXTDrL0rtV4oadBENXpRoABk+BtTPfyCYy3RrS22JtdxFPaFoJ8fA8G4Op/5hKmG0gB4pGxLx
L+u/UELm7JkUoZcuHSHBzIDsVbGuWZ+dgZ30WNfG947Lrd94UZbfR6Zy/a1dw32QRJeyV4FwSKqg
5eNmeQDUkO6vrnG9XVHiCtFcB+IobReGiVGeIgvrB76lfn4fVVvkFwgeZPCziRF2NNhQWjeAqB5I
7TlPVwyWSep6e4R3eX2XYfJL3pFi0DX4j+x0Xi/NOgv9FL+M28OStLYyN1ska5yPqn/Kgy99UmCt
E4B1czQcbnPWcJKsaVVUjp32ANnzixYP86ENhpDih7P8DHpW7SXbx7MEzr2w5sTjpDMFiRxHh8cn
z6n0cM9MTLq4lMZIhC6XZNrUrIgVKGtgJ0zA+3fNhcIZeZvDv6JYyNqkg3IfgI3/070UwUl4AJjG
XlbdNY4zKk+PS/LE+G2tJaviWgg7/AwrIahUqJA/j+swA+JE2b5n6YtFmZQceUovijsABHNY1RtS
5mTaGgcygk1kxsxcyrKG1fSc9gk49uLMGnYHfzznukidx0gQXS0pcvjWPZlWeBIxWLJ1khd/nLC8
l7wqUwFDjeEWCfbHLdBmPNgUln77Zn2i60RHLxtImOT15opLSzVp2gCt21nV1OTf+xGV8f81H9L8
HdzwGNVgvvJBhYQzidI16VMF3pUBMbRYzr8fUEEbxH24h2zYz9ips1eSyzgJDPZQFNt9q4JXVUPl
PBfK2k+yKfE/Oz/RX61UR8H3yCGqSh/cMa75WX/1s7NFjIFvLQPJne7535fAsZKQ2mYyye36DNrC
UlcSPaVWvl/8Vp5VYoGrijM+RFd8fwLNSkKiXHqeIYYO9UimOZKej53Lm9DLj3mNRYRAvEcvG4FT
pjpSIq3vGIYECynvu48DCKdq2YqkteKhAT8Ws7qj2Fs0EN4F/c0qGY098y/j+RaoGhZVHvtQMlwa
YIZE8A02a5tmBr+4+rw5FSG9a0kpqyieUXRVliLTZ3YFj4iotNZh/8DJFl69ucQNCrBrOTnEVEot
NYn81XNgVbsdVcrM9dGEN+BZqUClEqpOATVISxW+51We+zRugyQJ94f1jV18MxE08AFG1FhL6KFe
jq3apooW8AVWcG0FGcmri+90DubEoCJ28rtTITtHIHdS+NPNKLXFF2Nu0D217CBcvhDBCZ5rPMmu
HC9BMSdkrdyvd2/w1YV7KPE7Bo5rzaa1tTxRpfhzHQmSXKUepeO/LJMpBiNZGcjjpEG24z71JyQl
cnKAAyRDG8eRVDkDgEJUQatisUnjajI7AydDVmZdRHLXV5xGTGNPh7ZG23UBLh0MbljUhKOINu4t
Oj88+SJCa1a9rUCvB9BofQSsuipPg11GSUJFCIFLTi/Tmhv0uZBEswvZ9Y33OmdF5ccUuEbsc1sH
PVLk5PXcT7uL6sXFhKyqV6btCEJ4r9SjOmbVx+zkdPPZnyZ/Cg0o2YcmkxBJNXbkuNPgknSuUk0j
IRCmQEhxiRMXQ73SIbOImUxHcruac9Iq86jrCkvj5PNG8NNpd9KBDQHoVwV/yaHfldIvKL+N/Y43
sqPSuqHQ+ZmA5osezEi8YXd0RFbE7Pis1huoTuJGg6QuLA5ZepnhSgtDengfr5h3nd8ne6ORL9MA
AJUOa0qyuLOs5byuUHyWE8xKY4OZ+pDJBaXIRn6mfyTowAWomZ5cO0y+tXSs76fDP8RVu4Ku7Cdm
wPSG4qQUAzRCYOFYv4SufERIDclHDXJZzJl7lwCfOUXKjldLKqdVjoLP3Teurl+T1V2WZxeohGYM
bpfvaZuC8qNrzKSkyYrVLwf/JBlr8q+8yk2t8TiK7Yj/wQ9JgUNVvStnpCPI8V8f4kc78h32TRgq
AliRzavkqviEm6p4Y7IggWjH3XhvHUjHbqLs2jMqPqNUOSc+IJBXPSh6mbSuTSXmJRD8zgfxLKfe
EwXbaQBpvuQ/gZariC+XRsL3tTbSaDyZo3RWzHEsn0eKrYGjRLJTM2YQ1pzwg2NXpjg32ZarSuWh
HODxxxxue0wSRpYgda44BMN8b9SR2HHXucWe2TbKISOEvGqdQ0V/JvFvWIJg8KiFVZT2i1HRgxH1
1O/hb0nXPXJGTtyOCyQJMQovC2lxkJw2bnnwDRGRbycsoCpQg4HwVkrQoPFlSm7tQP3442evoXDp
2RwPfM/L6aZ2ADgPnE5qbirJ8IxSv4a1WVRlsdo5VAMud1PA0Bf1mHvcW1sMcCcr8YAPbp1UWyLE
vN3jNY87dpXHDkA2QsZyx89ba5LoQOTFkgBZ+3OrtIz4TvlniVBILNFS2UQsv3o5gax7i2xHVyP+
Ej85sMCFFtF3vZj/2vnMReToQMQEAu7LNbobe4AcYAOhceV44kM7w31Wx16hiYIp1NHZcHwF0Em0
LMtWEKK1LfobybZm+m8XgS+0M/4xpeYIqys+rSAqvhGecQA9HCiDkwg49gBUwoOioI6lq+QY+TVt
gN7CwQsOfbz9hjDsdEjysNb6XOlcXBS2qOi0l0hhm7oxkz1km79BN5I8QOXPyo5efaX3JAw+GGIh
YKfgj+F6+vrw0DAXWpCL8C6kTjLCO05CEv1Txl7Bmj+cIe1jbWET3apR/hx5luuQUOojeUuOdY4i
o/BpkIDAfxOlME1BW3PoPhrzc/iT5c3mby+xANXU7QxzrUw/D8lPwZiS1IkIQGezQFHbBWZctEML
cjEOCnYicM0w9Z3MNPi4NgOtfSuYivQufjBhMxzoej+tbLM+2rW8PRIMzWHXPgnM47jRdJbxXOfA
mjuihOAgQiZ5+cZMJBwj3cpwnCYCPnpo7+wwofNghNtQ7EyDfg6vyUrKRZuLTtbxmgcCa0PM4Y8B
ymvfz290MRpkYiQx9c37kD8vl2Tnpoiue3EYZZ1hWPrjqcfUycE3OPmB5fxbsdJJGI7eWAl5Ok5a
KM5OVsyzDRQMBLu786KE7+IkLAWQiwn3XEQYQpGBYibH90qiHMAmJAXrHZzI6vowwccPAA5E/1IZ
xqf8q2AdUl2t9OLf8skIUldQhdSgTq2AumcPB6/mqYayVVp6xp5k3nF8np5qdUnVDmiAlyaz1tlL
pNymAjzEotEgu9W9a8bwhAcFvj/+qWKowsqTIytQmnqlinMB5kJdGlPMqHWM8nHUfCbOvEyET0D2
LfVuQK+Sw84gp6VamRPDxXk12Bdh3U8w+k+p/ExmyRNGvoa4FcV5aUcX6qU/YxMfbYwfoWRLUW++
WTF3zHDd0dUQCF2a21f1UOT4yAgvSy+KdPImS7bhkSWcVKIi8A19y0w280X13cOmxf/Plc3vHxLn
fxM8pwxeGqC1HZ9r+S7gaLJR6qYqNXjqdBEBFddDncA/yDr0SPnqhrJIscqZKgE1otO7iXrh+YeB
KBFQTg/1vCAnTSu+IReP1Y996rShkAgFKyq6eb3/0CY37gsamlPIXdZCIzGIwkBVv5Y6XhUf772E
8nxfNFJess0fWrBJjjtSWfffTq6WwhRXYeWxJFRnDXUxt64RvyV7gZp3HfIYEpX0a7zVEkHR8lyU
30Uvbdqbl5NI+P4Ub+mU8xOoJTTka9pHww3X1xMpuKH/vuoI9IA+acOEfFJ+SBmX/d3AlhPh3pjw
+2aWiCsa4OUTKQcQSOW9xRkew5bdq65QR7XJWBN++1D5igseJ2sjr7mxkjJLMQVWIQ8NhK15BVE7
/hUYcV2O6sMa+i2pVpI0iZJl+QgBEeSUxX49Z6NoEpaX8qe/Wifk6u9IhjQbaKHk6VbAud3/HLcG
F3NC9KxbFlqvAvDQgIpeJyzAuqrtbdob8/1XZb+37o+vwmh29Yq4kvBSmUtOQGBdSpzHKX29EOhz
zeZGbyfICa4OdLxPUpRor/dVCwaa+GM+HN4cKS6OB0/Zj9zrKfr6wjlyDSjekVH6pylrXLDhHHnX
hrqX6bS7gYl1LXLF/uvbqHozgdrf9TLfMBD/vhiAkObQXS/I+hnFZodMjC255V5YOimEgxqG6vYi
+KG89X4uSZZ7Gg46EC8az8S+r05/iTzKYgl4qsw0VgEwG4OuTh05nIEOyaz2a6SS8jkUR722aq7v
tlNYLhcQ/6jsZk9mxeTY7QR/+4daHZzrJOnxyQeHzHwUWMP3aVQudHa8qAGedMNfdx5LJOjW+qz6
wyNoYGAyGpXIT+uptBRkaeTYAjYwMIr47lyPx4Cv107LN6VChZKkaTQwDHQJ6eUgEiAnNtRhs51A
ubv4uNjekfc/z5sFXfWLhsZYs4gIJMMml3jXr279QMrNsJ3zPdIdhKCD6ZqTFGDp5CluVPKUkUyt
2Ht3pI+qo12YTr9Ab0T5gR+lsOsQKna4VyiSeJXVnee8/Wkt61Kkfmyh5xIERCbTsrpGB/QloURE
1p5DRG8zWcExaGR++B5VRG93FQO7t1dTBMTxXzTulG2bKscVSK4AbpRgL/ZUd0/V0Z3GLZl/pIvM
hwOApDTen7csWNhXwdsWjYqTeTUWe8CMYBX1J91ItKqME3JCmu4WivlOjtRnebld8cvnbwT7dJ3j
2R+udj9EcTFIrhCwUV9/tAg5rYWEbrd0Vc6mbmJ4LHdDwCrP7loXCGF+1RkMX9wKM2JLW0mGkxRp
Ph9CDb63dIs/5qxSb1up/G6C84FjYh41StYmR5tYdIn29clWY+mzT77eACehN+IB/kd4k/MmZI4d
oY7O/Re7KN5KZLwyZ7d+DSOHit2PRxznAhhgAHw5+Ha4Js9ndP6EVSMrM867OhveOlkPrpXHr4s8
BRwXhTcMrOjGMfAVaIR8Q0HwGafSlh+lZD9AW269TCfnbvyCSqyfOToCIFNk7wTCcw4OMIX2hWb4
daQYnUwxu9vgQlAQBKz6WRCQnSIa9gwptW1w8cfvz4J/N2a6Na0rM/R7UP5TkW7m5clFXRnWtiEQ
ntaI2umBRB437+5Y2LOgxhRr8bOgR66oLW+UIkpauQStbB2PuG9Og2QGNmUvK89whP2uFLs/DUzg
7XF3u5XD5/259l2/06xSv3wfjE1aHG120y6jl0B75I5j7b1y7K5atsY1jvscghUNb5/1UUz8ylWD
2GI+6oyu0Q15vqUd51rfDa2HjTfgqVsJjzuX83RyL2h8Eq9VWkosJu8BOWCahejjqR+Qb0zzLzHE
VwS7cJ8WaeCKSuy+EfwFJSn2rKeNYthY4Wc1G3bfeEy4XWwbLKfVOjdt+m0E3a90pKWUkZw9MtQi
nLpAS345VViVnHXrcQuMdmogpvm8TFGvpj64IxPsESXDDQys3ay/eMJaYtlRtlPYE3N7+KljNs2W
o6z9lpO7+fF+1dKYtqQqmMfy4ybuamnuGSc5p+DhpxdQ2xbv2MVen5igsSz9Tam9eLMxtx5pO9y4
mtZa+FMX2aIqIlLbognx0rnkfqtekDg6Q40O98iOVuV3DDf6f8MFElUkQFS1segwvWae7HHKa+6V
sRljStYUtesJ2N4gAfE7quI8DqX0DDToV2cB41wUchANiumk7Fy+kQPGYhOFCUN24IcgixXbY+Cz
2ocNML3ycDkRulyk6R/x/4ZOldf9WboRa4mcY4c3v7rqp1FVp9ODFaHEqAffK2mFKIF6A4UppoH2
zBB30hb/d5NPBksvIO4P1R6MqjBWoCgDE3Tzb+A6jAv+k1Qrq7H9/Z22Lwne442vF7NawfGuMspL
VQFQkjYJed1vNqaBUqb3f4MCR0ls58WNoWJmRf3mjDoEvuCCZ16zl/1qHaEPSni77FqHIVPCq4Ul
G9VVPo8GoUr9QLpQF7raysGmVdcDT1G2W7HCHwnyHd09+jh+paNLGxPTQxAjXO6Sz2oWZFM0oeQM
cea6r5wKB69TO0qhF5/5CMew/H69RdrmSROLawkRDrA0uE81uXtsAVw+zA9QVev4tWgMe4EuXs/2
fMcK+v1UxJNEnFrp6CrQOXNfHEzA9b4itb9g4xcGbmUocQXh2t96fJVp/VNU889ODpxu2QoVYZVN
quTbW3dOwdR21KnSvwXVxMPIY65RH1iZI2yfzJQRTh5JJxYYjcFLY485E2oIPQkB733U3ymWyA7I
mRi77D/z8JhzdU9P4KZK4vGklKBOA+Iq+TPTcXkc42u9ZMoj1qDniB/tMTJNsAYc8Av+NqkYDEbF
gRZL+3CuR9vD0ec=
`protect end_protected
