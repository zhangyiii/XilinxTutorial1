`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
d5VJXu82JfSwswDjhvbEU9He9tQ5/1Rw+4/2nB84LUuT0wfekcnbAADJNd0/JtXdeaCUlOw7Zwks
Bp1VvQeB3w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T1a12gH9+o/WCd/uq6lAozrIbwFwnflilDyEA/rZKRAxvRmKOSqBXtjVpxVSoEgX9El2BLPK+36k
Vd8y/iFx5HcwlteYeuYuGTvgQerRA9ycH4Qwt9s5DC83MaSGod9ecMMI8PPrmdJ+hCOX8sXwEsN9
IHAKBa7h08XDRsgW0os=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZE3CBd8eugZohbo93EvXvQkUxCnosHfYT2eG0uuvFgW4E1aUdxFin2hcHpeAodvxBTyPhYz4Lsqw
3nsUxnz9hTb8Lhj5XnlqKx2mVFP8Z35n8lJk21C09QHBGoSukklDPI8dbQUv/KxN+k1qsLBHfCBA
FWz2UAwKlgCaoOPe87s5MUwwDM1/P/D4+XgEQCRDz/7JDN7p8ZFVtltMEx51xjJOCvfGoEeTzG2k
908lkYgt+B4pvwsuFOHwC28xicC9lqwuIR+OiqTI+hvqIl3tijnK9dhEHXmlIo9PqdVp3p9K5niF
C0wKwI1gK4zk+Z+Qv31AV2g5KDXjXxSpUgHlpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1K/c2Exmx3hO4tktdfNX/hsUCqBDw6bH/vDRPja11f/SX2mhefMgy+yYp/XXIVeJlyTPI7AwLQ+m
jPsm9qUsxInkPzY00BDkxz+XjPmDvPZhWK1LaTfp3S2KuDInJ2AYP1AwgClVQtpRFpipBFYqQeNS
QrfV5V8iPYsCh6rtCZ0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z2R2Fz5uoP9gCKKJ4H8ByaZdL0II83JUVbmmEiqboGhJOssYqqghHZS4Xla1DO6PE/W7lUbFZBMN
taobe7WZ5vLL3z9KT5znQ5u/8vqZfQZBnNTCM9ij+NRl3PRmkUPrtcd6xURukGspBspXFvJDNTq6
HoC8rJF2dAK3E2hXtQ2qzFXYx2JspRBZw2ARE4ENjzYZSYK5AhF3nV89pEvyjDlChnkSNr7Ec2sz
zSK49rQXLtbokqxvvzCHRCEs+NoMqKlklN93OyjJFAIzYffS6GiGtNeycU755Cv+/fAQynybNWn5
4vdHnb+JcudvHzAJFK7/azTzKOJrOSm9uJYTZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15232)
`protect data_block
mvi3i3MBI7n8zvuunOT1BL4eDGhQlMnzDOzVrYI8XHOS3ZoKFTTDP4UmKkCCDyXvukS63/BOGJv3
NoJdfMFYhDx7pjz50AatTRm5dOIAKktHZJVnSGt5h4GNaEO2RZrMb78Xxh3U1zVrxlZ3qI2EnDLt
tzneGFiBIXRoOP+GoM2W06jBPrrgnMLIYYcuoKXoUGoy0Tu6kRojjd+rMZQgJ/YTCFAFQ782Og4/
vTA57reBXbFiXcNw846W22hW6Wh2b/k3ES0Bv8jWE5mlls8Eg2bW8lDyRrbFvs2qtuj5B8/dwBWm
MEtP72sPcxiTduS9XBPqnMKn3K0sAVvrEoENUcZLfkCWr0G+r2JynFIGKwV0zPqeo8Ixf+NstxBT
JGIxg52SOXcZ8Kepa/HsjgHFZ+JwNdT+dx6JRDR8yKPBYPBub9Pf9bmPBq07syUjwwMnGp/2pUde
wvlC6k7B9pHq+/215GUQ3dXpc5xlKT4CRR4/4O3j2tnz+lkuSBqhuKNMEkGhT6pCsaWavsXlA+Mt
2ut5F1Eqwz3V4cpmSnhlRrv4c7qbcoSek9mpUp1aMMoBFdLckn/r6qcDOe71/1KsqonhHDelycBr
bkMhOAsUuOrVTt3RpH4Ysfg0AOXj54diS+XD3OsfxKWkWi8XvChQjOBp/6rsyGrEncxl/OwglwyA
kbD/R5CtuTnuV1vfka7kCxZwyAZbRjiR//no7IhZ36v/qeCm69gqtf8nByIdBGstNslFDHKv/yno
O2a/Ecd3kC4LO/FdruoL+WcWJRmmNx1UYGWbQyfeCVdoA5ieZ2mwv9PTch6ZerarpYiWX3Mn2E+7
8K70hzw4nKvyrxjr4IFZXtJfDM6SJrdlFeKhB3yapSkMf5W7gSjDHPpyfZASF/6D98lRwHTIynKz
8tHJPBNjObYETnc4um+aes/Y9sKMH4AVdx3F9Aolz0DWGGMqPddQazZ+XkmAxrB+ydGyQL9XmQK+
DSF9YbWxWWzMGQRKBiRq+pKSbL2d8OTboDDxIFHHwH0bWBuZUGY8shH7ZTzgAKT6UbojCUl82kVM
RvzNcHmNa+za66fu1Ztfeu0d/R1MIrkhj44EekCDEMUejShLRuH+noVMiXpcgF9dQuWVWhG0xZkW
HKfrY+ki3tJ2CLv9BEXkD5fJ/oTryqkXlqxBlNWeHa1lFxa3AvUizy8LA8c8dtVGHbRYpPblnJ4f
1S7PKasFTL7+lPhbjCbRskXF7KNEqgkJWVdvW8ktbV3XoK0uyr12ln5P/k2IZ/h003M1SbFkvJ3F
olU/71sLRLUnoZD7JLz0JEMQD8GLH4enhvnQCI+LUgLDFcp6utYZoYUqh9PIXZBji9pS5ebdMyxi
UIvgEL62MtRekto1d/db/NZieedcHqr2VfXfr9ukgBX9W0M2kPXK5Auqwz6vYljoSEu9uFRTivaz
QEE1LpBrZ1ng4pWvKHBihJiohBKSV4I5uhRzqyPCBFs/j1Xtra4t0bqpWgm5qlYoX3B/lzHB4PPF
g7FT7vYrPb2ejUvREE9ey3ep2oau/t9qKN0q2NhB4bHJOFwXk62N9U6Suvgl0IrZ61hnx9VRpnvY
u48HiWBj2Tf6oIam6TYounmWrsEfI9/rJsQW2BW0kO/GxWWZHZoAsFDnU5VUrq2o8ym89k/MlnZZ
8HKVRbElEOrXXNBx+dXNYu5JibyNowL7YkQcnr3jgSSzR8oVszZ3Mo8Usv10bWShGCI+M1mt/KBq
MkeGlcJjoh0NNjHRmG/GK2oVvekIO582nRT6qAc4Csyoo7Bnr7vSAQ7xdFP48wGKUjSMRhXQGiTo
vF0fa83/D8fEw3SMftTKtkCvils4trW9J/v4TDR8PytvlYvDKwgImiTrkl9RJ3N42gd18uZJdEOU
bvBhK/kU1PdZwxbwsrk15q9qf1l369555IwSxvKVxPdSXfrQDt5GNxDx/90sbDy2d8ses+rtlGDQ
j8mMCOeHXTw0jzse1CltbkjGIzt6VjpbGOrsStAuV9Ggj54HL531J75eWHXeEKQkaQpRxjcwTAB+
BHEjhIuArnzEc5tyPdANuckN+SakOco6FGwXZmCwDc3zvYl7Hh2tXz1ibpRBl2m3HBGYLuKuCDvo
dayWWM6ZJGTZQks5Cn2KbEo0sWopGnHMXaVUZhGbRVpUxzpkfrpDmQOY8ZFnf6n5o9Kt4i896TQ0
GoHsnY3u5rL4BlWaIXicOpa6jDBJTspewjGcn4YRE8mSB48f79efn3O/OCYtePCES63t8g2yLG/d
tPfF9kVn8qzWYDyXm/907qcZ6/xp20Szz3v3881QkKs6dUCjKra2DPI4yw0VqxGsy1m1AmZBxHkO
9hPG/nhYNAfn6IM380svQGuYuEomyH3i3yfwmbYXlCxZTNKkYN17gdOdm6oX1RSI8LFYo5Izg6GQ
5UnIyIqwekWPKGHEAo4N0cIjRpW/3gbeyujvMj2V9sI6ATtmIgKHfABJgDW3weMPaPu3X3QXTRJ7
TK//3GHKDZBbNpeXa4NH+J/ZKKjVQuJG4xShFijZiw2UGVhZwH+50BFHONXoxDQueHlp6NzpltZO
RajqU8FPd3YgMgGlyvo9pZRW3N2mOfPvhJ9UsOaVUjnVpXCpxD2VrkIavWqf4vAHYlGteDXxNgry
b1nfHZ/SCoj8PHADVI0SR2Lunsn6dXNOM61H6pj2hHknwBp/7EzP9qwxNnqlYQAc5haYVSGOXugv
IPbzlXVMm3CFefARQS8HoDgA5um8Mn6xNK6uDQBQpKI1KjdOHR/43Og0M2LMS4WU7y/23zMNyFCw
URXTPofBouuJV4WS14uF5BBIUNzygSlP2DCLHePU2qaZT2eztOHTtjbjjfC2V+yxAnApFkw/36tY
3+KKKbiCZ8p9xfq2muaRaVyWtlidGpPDQaoHkcBtZ41tAHMDFWJe9amvgiheFMO31nHwIu4S4JCC
HTgi0cKAvGY63cWf2T2Jhz+j+0lTuIcfSomkKvSxMCDaAvOH+iufnULEV+vBHMSQtAHzuYAew/U1
PDQtmrkxkE9cSS5ZzzYp2M7ERPbIbbKM1mdMlxGYoUaSPZnefWdXcNwRc0vCa/QBnsCwoZoL2Y+b
FRWZJCAeGKWBEFePxG2JsVqGacAmlTx9EgFG5WPYqv+JAl6YqbGtHC7fhUiXkKohqqu+1Elp3D7J
Uo0FJDtZr5ZSXWmWnxEzfdfaYOlta3t6B+NXu1yaE4vB58zOavFnK7zPKFu8gR9eJ0gGxh61C1ol
iER8GDbmdVAnZu6Mtt892PPj+IC0v7F0P6zms/CT3rVuNs7FEl8/kH2kJJ/QK2Q5TTHCg5BU4Fn6
P10kgYM/dlQoQiM9JHeUkGsNrX2gez/cOFrjbLIk6tFOQkagTscMyYbL8+nDCOcuV1bLJpP3CDPo
GKpZwNXMACWzXHLMy+5h+jpUYLP1/SilCyhNrpui9vivh5AUbmyZCvf3NpVZaatDb6kWznSsCiiA
aNcdKhNz8IbeG/p/aWTbGW2R8v7Vh8INyxbxK3LsagiXdNJGvjyUEeRE5TBS2sSZr7mfle7UmLU0
4JC9s0/TaNNDnYmWOESVnKRZGL97TqcBUUTzgVO7MAmQBRium+ea1CRreyzHH9GBy9wK/fUJ0jQS
sLVT1G3ardq38xeAz+fef6cSpbNoo4CJ57hrJLOZdEvN4QIXdeK7KHSY2qvhoNTn6TdZLVVGTe0Q
cYApj+vQQurkp7GDGji5pdo7fmVbad2MxLISpfB+x9wzOARMhOJTicXF9kghQLiTiN1p4u+cDu/U
iJaUyFWTbdfzTrn+OPjnrnfkEy6snC0KOK6cDlvDg+JD4Y9cAv0Jdhm+Fx2KjAGTgrA/JJdYGMTG
+P5u+xfLO0GbcjEMiUTIhEA/061DeRB/RroVrt0k5Lcwl+nfIlo6Av/1Q/JkPICRoLS1cONooSbP
jjLvVIQpK56QlWjCOIFime3GLxfn7H9JQk9B6mL8CkVl697bIA7HEoin3xu0LuUHOg3zXSkBEu/t
C9KFLLmFn/RuhVjZVckl0ZVdlBQP9s0QTVIsnJJux2XYS++px7hKGGeiv6ziwZ2Pd6bB538iVJca
L0mHbo3ot2D387jidLPeFeyz3SZ6tEQm/AmzzOcryaLfNrHHOtp0d89bfpY1Lfbl1WTGKSucdfGP
EAAgdpkYHZJd3V01XkdLE2Yf2P5x2luuRgOrKkKjCJvZYzxWC0AEhiUwtfWB7oArrrk5AZlCBEuy
XtQgX1pMEoJAy2eO9YyldpaN8CWMvz0TkZG5dB6Zga0OaIVYkBn8zIiWVRL+01XTZmhZSTjbQPva
u30qUxWEQPDvvUD8zMvNUJjl64RVLiaxs07eKsBe13oFVCDaAqeXtmcTAuSSA73IZd4JukPyQCgA
BOJ0YUqTDZFlik2Od0wfSq+Ltm9YzO3zaPBnH9CmGIgUhrr4qE1hPTXxgDU7EKIqN/XQ3pedrooK
PD982Ph4OlqP8lXyWigPfXEapVl7aaFqE9ZTEOzr49kYMglzKdAdqa3LfC+4hDczBlrBhgk+QYlj
IvD9Psz5G6BxbFKFXTGPbM/83GTN3JBNCVNl1MCMDc3GiT9q2LbJrDo5v8/009P8xfcuGEget0kv
biUV2q2sz1e0MbGBE3h3+wtH4LXbul1WwjOJ/3oe5ConXvX8HxSVqButvD1YBRVV1EYoqyWEzYPb
SxpSkWA2dzPyFljuqeMBikCOGbDswU12WPm8pFff722cSAlf+OeZqC1i8CYGK86axC6x9fB7erK+
fQyQ8Zo2vgWIPhtVQt4uc9UrZxD61wL1Onwa9ivKcTQyySZj8V9VYeLxPrkw7yDs6pzYEbV3oTfR
r99rPOhaT38rERYOPy2hLoXJWR1ersxDYC02dH19mNlQAy+ogToQI7qpk2wiiiaWbq+k5e0cmjV+
h2DpjtuaeOkkiweft/U6+B8JA6nxMCjPJ42fqaq4js/4JhPRxIlY+jqpaL2KniRWNb1ksruZYXzm
NicpSrfYyHtJ/gGnpgxDHS0yQeOgUvVpII3BTiLeS1mVISWhozKB6+u8VpURNHckUR6036r1UEIv
+CHEzXdtwN028meAAakzFeQ0AHWcas1bKdC/cPSB6yXU+u3liWbxeuiSIGWqsbEVIPb80Rm6BOdP
vspevoYyjhE+O7/VHiUZlp3sINYxL3aBjGMdUYW2NjQtWBdprlztszcm1Xnhi2w4Uxj2QiN1SD3J
Pim5eI6ZUwaLK2ULgVhJ9CrEvOVwE6NS0cSMFyVb6IiHF1PGeO4aIBp8b97q73bxiSTlQkdu7sij
RMp0HBqWBv7MHWSr53hTWA6SOlzaEN89hFME2UKr3MHUD2C6j+Y6sDCRAKu+0U+VuBu6Ay5AE2mU
iAqrX/QY7YqJnKZKIFcy/JiETH6ZMlicn+n5stLS7Z8U5jC4mk/HlMZ6XjTr4G0W7dBruDtAvVt1
g0w+O/IDxDNolsavE0qO+HEQ04U6DoO3O1MymEo/b/gDCO51jyra80ZwTfwMMHRwiyvvubkBIXN8
Z9wJjXBvo9iWsOZ4H472FVwctmFTPoTaL8eGyB/gmg7miWJwN6vGIgmdEucMXn+KEmUzZ4Ciu7hY
rbWgGgOXoa9dAxaLtnf9dHyyd7xrqpy+AjYLTQbDkIjVurODih+l6ZrMLnGmo9clcSkQZhR/SSPJ
1rdSrhNZpsXeCiOsUveqaM75k34txN3E80O1prcHHdrZse92APcgybqUeRJNVPDAoBg2HzOk9E6I
+eRh7Nnz4UkcBvswMh1Hm4bbCktJmbNfhELncbXfrkdJB5gRAVRCsmVET5QQ+IAgdn0TJ13P3mSo
47IMQQAkmPWZgHVIlxg3DNZo5m1uci88vS1AdFmaDmc5vAsmsJqYdceK1TiKVCSthjIXTEEeLlfG
xzuIizBB4kmRFg1iJopwgV+pfZr12DSIrc6onZEGSUVOI40CKcRBn0HMGQUGVj/FYHxcCu0cDqV9
k4VboOw9mTdHV7yjdFmIDkzTuZNA8P2zHq0gRCu0QncRVnON2T3ekGBHotul4blnRvx6YvqJUgad
Bo9OROtfK8U1CEX2DztZ7EyJ2uGOghlKNA7rRDuXZIsbrYqCPEV/sfQLGpW36TlE8+6RUmUa5P0z
E+O641xXd9q7Q/KeX2ckNMWxdH0hEVT7znudoVnxB9wIT2K3m7a/T1YUEcmIs7ZRFFbVQ9kTsY0m
JHXW40vBy93qra/ggQHgZeQkxMs4mCaxKHXb+Eos7jFkHsY9GuAl61eAHmib9K5vPj5kvvNiVj2c
PbPJm7ejKhU4il5dgSNmmqY8IAUIvZU1Td3vxDv6Y+OrKWRjpZEOQBxY2Cjs441h+0oEpbwkpPMV
vw4bNGbtPaLiitYpTkc41cbSND/gk7EGVc2bqrXl0/FkWMqzWt4KD4Qo94zlcHMzmw/raiB9uWVJ
1rC3B3cq6qlP5JW+4MfGFJgeX0Psn54aOcWv36YC5jdnXBShXMGMgamJrY/uqrkS6P8Y2NeblXW1
gK41vPQhVrCfHj7lGy73cDF9mMc1/Ao1Vi/dXgeuO3uAUf0uhV74H2bXGZLpNe7ZKhH5k2N4Q2kV
eqOC0Mh2pE2vJWspK6HU4PjtsAg9o9zteKcxkRo2+K3qjx6V9j6yJ/3xj2VW7dwXUg/rwWWezH71
S0mW/zwxu3e+nzA9AgIO40n1kOGxEAQzVUdBAys4uA7rLY6e9vtC0hugHOuigwuu58tvq04XlmVA
NnastekFHwhFMvAQBm6tSdFY85JqjPBkIQzy1tgdfQeTobuHGOnCYCqQ5eC6Dgmd9Y+o4rK2RXbW
tqlFQIBIAl11WEqDwQbmXAY+01XCvQpD8fxD0xe+twRbHq1VhiCBIdYCGY8Z4/m2EIuyRzl47aMD
RxLzw8ud6hDZblZgmJo+cjErBpaMMVeLidFbRxNcTWNPZ9fQVawxqHDK+AD46M/T69MwkRrG+tvu
OpnL/1WHDhSMbKKkEiZykzhuyKmjbDXRyXYMh7P7niSpgFJyLtD8lUMZpf0Py8R0QL24WKgvQ5aO
/2/oVGg3mALaan6skvvILsFNWRtZBly3YLMcGdedYZg6CfKKerqe+zG7Pxaiy2WPsGiH8d8RFKV4
epXwmHmIhkni+GkruiyhA3UccUYzw6AY8cybPEJ7EIZZ4RSdoEbnwcy+PETbxIBFjFFhcAiCDhwm
pLkJSzJ6SyE4ENrmfRmcJrIy1X8+fpRjb/Ajt3Wv+fp37tRJdqROxFou+GBEYiG1kzSUtTw4a83X
9Hx64jISve4UYr0Gk2lTxaAKlt9C6JHa4XxpXbicmuNcEq5Kvy5g7+qvMYpuzlfcye4Ew1ephK74
tTQV1lafEvBM7LaCDJPDBsm8mJvcKg+X2GNUrZuRkcZGYQtlukTPJzmypM18M5vjNPZ43tginKFh
g+6LtjQImcabN+AkwnOUSwxGlk7b+c7IDK9D0ZJ3vftrpXnqYkoubputQwlFGNzx6EWRf7AWyc3L
y88j0zKEE4TfnMJ+NQaKnOiwX9aqd5wii6/oWYNu0tEYmJ3g6BDP2+ylArJQnta4l7ntvSGuO1xI
zjiP8FCvScPfzKhpwjmyaVRW+LARt//4osoQ0O5DVdcqnPt2mvqVK+nFfIXuup92tVBBcMAmYzn9
hLLV/Ljgt1jmBKfixGr/P3lBcj230Wc5k5Xxx8jdn+W6liI68T6zMB8fLugywEQ1vguup8vtgmPU
BUqzn4ihaxFWPJlkSb3A0UJbQEVZAw7nlDxW+BPC6PtE0i4JgfRcTTcvhr5rKNU5j3Npcl4aws4C
Zl7BKmBRvbOsE36JnxcICqGvjjcfRSFEqGi8njmL/SF2jds05L8EWCYBDu7kcYrMTCedjxxguUGL
42++FjaNMh2wJHC8N1VD7hp9Qkcx7PlWBL1+L/bhCyKJjc+SSvIWxGQp0Fq5nNFE7MJDBhVD34W6
h5xONnsH4JZuhT0pi8iMEDzfTreFoP91KoaZSB2g+LiunV63UhK32sGgQfYYCo3mhSDQx7eI+SUi
Mk2B70Zf8prRoM9M0aIq/xbAm+2Ii/M9cTD7jF9STG+LlFmxu6zMiYk8CCOQ7AbFU1bTI/ZHMJfQ
Q7y4ifC288Tteekki+U/yWpdg3XeUfZ8NGJ+adzkVFv5/zB6ForVBE+mC+iBkPNSfOb+vyL+YN75
Ee8nB2bz7ZTltXZP9u73CB29f/6Bf9EfDzspRd7qKNd2A0npmznCdfdR8iw/MTTtORAZr9aVUq+h
HohZSGdDL9MUOeGB8ZmKf7NvQiHufvk44MWoUhhsEWnLMkxwrQjvQZddMOnGLrLiG/jg6CkBPd16
zoZEfMc/xnz4ZWFKXdofOCLcv8P6GvGMmlNsy6Fi2sQWEyOh+ZHUiH74aBqlAxgu0LtKr6m7WUdA
vjErPkAfsZryBYJQKqdx8PgZkCfelQax0FFIMvblGLJDCExrFAVQTQ/GyY2ShCEEXQv5hmSJhLA/
YjgSdou706XqaQHeDpnr5DC2cCXgAKoy1PcIy6jjt85rIEUJZsWz49/iNpxgkce9FfN86uL5L3bA
++hpXXOyoyo/z8oY4HlhR2uNXfCT9dxoEpFi4OFwLL2/Ek5qPYG+nd3SAMBqzGurUfPEqbsCYLVm
KDpSnjDPQO+fxFrqwOQR6F6l5b/AooBUyvs6N/IjzWgCoQifc20K+5gksvDWblJktJ9JUhwf+F8D
1f+JJRGzDp8zJDFra+ogXMbCe7JU09Bf19WaJGCdZucY4LocLDP2vr1iNGrekq/tbkztJFpCvxBB
OgJS5x8rVH04nZJaeIVDWFZ5HG0tubJlOB8Trm82I9YADLo30/gX0UlUA23hzaoLeNFqhq8CBdh2
pOGMDXuWIvkgenzoBI0v4htOLCpohZU2hD99SHF4678S/CarevrmJOHvy0i96gKaH5nx6PKRa6DA
0grnKglBWSPTVKbU+prS2uakJbof0fFOry/AhmhemQ4/JX0Bzf6tM2/EPWDgZykXmhWxQ1WpNG47
1uEOebI4jicJB3hOXr6JB8sh8EHrAanbq6A4ZlbJmzvxwFLr1l95YQGMHYHAiYzz1PhI/zxZ8SZj
N/ioz8uA+/+rCGjb/tOPD5tliTOFFToO5foBhrS1NGBg+W+i2aMdhDgBiQ4M7BgzY4d3c9om4D4x
4u/BR7Xssh37gycAPP8xsrTSLmhloxpjCQWKTOBV6AvMd+fteU+oBbf6J5cfwVyAxk6HDVbVG7C0
aHvV/Lj54FUbCrWi6l+mhFYSPlY0sd4db/OnpRQwMcd+XvxP3Q+/cJ6b39VCXUCD1twt96q38Tyn
7zST7p5jR+jAqdp4LjEOecdb+u5xo+w94YMz/KWLgqj/koAf1WL0bDwjJxoKB1WqRjzg4OaT4EAZ
Qz5G1L0ojAfUhxE/EOwHwnzF/P3ePoDC5ZZPQ/3UeTVRD0f2wrrekJZfWWjmC+l3zw+iRxoXOmo5
g5/iiyY6JQPtnfudReTLFA9qHo0LrAwEJ9W697OCUYoSrHFUE0uW0ce3aPtj6dUM/n/tTgLcFXug
2Bcc29ASFWDnTQRiAsYGvjsRcpXgK9pigXUuu0EWxloO3wZFtLvTAX26bSk6cHbwQJmf8IL2DDu4
6E20jILFf4xyF2rOwh2rZqbVylTXhZdkrOdJUjT2kQMSTT5NpQlg2eIcEL8PLP0jN4+6/dVY4i4A
nqfuBVzo05dQlxJEnTUxw8TGyA2I7nlcYkIVWacqvbgeyxQ6sa+4TRNQQ0ssO6LXnT+sqz0Etebu
6F0DogFEqY1xYY3CMxeQ6eZziturqdstP2b/fwc0ZKa3Is1pICn2xQHuG2sH0w7jnxcSIbXB/993
jja+7hpbTYe3hwD4nJZER66Pvcl31hbr6Y4LjmTJpBVwfjolvJrQ2ENkNl3HqLvOFeLI9NHUR5uC
fuHS84AArXmwKkHxEmAdegRsZR5329QQwn5ok3e+rZqSdrqlzS9ADl7ymWQsGHZe1RjsoxiENkNn
MyOXLEk97vH7W8QTyPppFw7FitnqciAwUbPRl9j4Hz5tX8orcN/Trxgz7FJJnpsu3JEilUX5e7tW
w828O90i8EZL3FAECLNxJ81BF7TbvW74NcMbni6rusDPIObYhJiuFNScGAWG8WcHGM5yd9Prlvl+
a1SRxSpxdRL45PCdLeSWEX5yfkKVmO4+7aWQPQkDNo9QCcAcLwNZ7mXDXeLkjDhsMZWVUJcQyKPD
TG6DNN5OOYGRxh2qECWVFXHuKFY6j97Xhu2pNV7pM8bt9asL4Yd9RZCWUP/ZuklUzJQlrD+2M9k8
ac1VIk9wnmMWaUiIvcNNkcsr4a1uXv3WyM9djM4a9JDh1dYsjvJmW1RHQqxIyquVHbWxYHvTk4+h
dtSoYHruqNvBS1Yh8YFnY76IFCo69V3P5e+PjaXsAJWxSk8yUdrRuxQwWzFnz/GcILJbL2voBbeo
NDfJ4PEBO2kNuLWtsZINC2iQ9hucCUgBJtB+KMfsShFwZF+PXy5Y3BWIod/fD/BehN9xOU7Buwrx
1dh4yLi5nT95T8K+Z5rWjeylG1n9vGh9BEhjiIpRsZ+7yujHNzgQTvqsFJAMRBjxjuC9WRFUaBGv
SyXdRQV7YofhEBLg3CbTSFG9yNLbx2CNgqyXLTnN8X7RXHhFHmMAn3qYn3+bkqCT8zsWcmkooaY2
qDhqIn5oi1zQNsnTJtJ2ozo7iHqFey4kDTY1o6jb8cIqT+1yEcpmmFCVJq4IPh4YESpWZluu0+Do
abhcF/cqPFZp18zzdVosH8ydYQUct8qEoC6PyaIXW0ioRcjgiN6ii70C1ROpOXwE4AhK7olvsGdp
52MuOiyI8wuL9bbQVS6tZ1M49VPA7SWyinvbDV88CzuSS/wPugwEpPU5EF7ilX63VWaREsIibOKH
tJWXRk5I5kgSbYB9VGjtbTHL3zIJZKk4KmiILFzxPeIl13KrMbAV9QH6GofPnxDj+dF5+q0SqSoL
QSw2jUVhZXsqzyaA271tO48TyYNSjSxJO09w399xMoabWnGxnWlagPozixcnNR0k2LVr7kVPEK2u
MVr35LFt8KacFzrfGIHUApU3Y8LZbJpSdDU0nAY4J5mWe8O9eo9FhaZ2SqzzBjZYQ+dr578gq8/c
h2GsbUVCUOGx83uEgJblSO2pn6+tWnRNzriZIw/XTLZ4lv9kNYoyun8IcGbDgobipY9GjItRWCh4
j0ifa0GcovviBzb5aGFyDp4nHMJRab6d2UGPOyzw9YEk0bnywl4IrIPstY4iRMedB6Gf9gWUYplC
5CMzzRw3cL1ZiewLbJpF/T/p34GehnMJNqGzG4v0wVNwWNHAG4G8V6BXOUQp3uynZkbtjQ33W100
PPl15gZBz4sTtWFPWHQ3aAO6uA/Q4LQHCh5ER2XfUubrxG84AIKF4fNBclrrXJvZXlbBlaD1SViA
XS/vwtKu+DbpYpFQ/mAbnb5jPzEjkZ+/5NwxZjn/g43oB/fynozzjWsDJ3P6ZvNJKqeRBg3ak7Uq
XahWmD16GmTI2vg1hx9WfjVXFSXoBBSxj9fzZpQ4hczCFIwVcjRrijiy1xjULDlmCKa7yw13djRo
BDC7916ShugVEr3i58Ys7bYQITlljC3vor+9DsuXCcpRkYIZI6kuKhIUHKlOMiP8uqMSUa+wSh8X
tHjILIczhkMGswA4nNouU5rNCI+WAQNpGWIaH9v17CPSmRtdy1r253vaWYF6I0cNkQxIja4kf5At
0gVl1HPBu/ApmdKcG+WQy4yL4UO/dSu2P8L+tZK/GJ4n/Ro4aRqK0eiTn82Uj/RUN+LYBCXaNRcF
Y9BN9UUgSpmbcRLXIxRQ+w0U1Sd6SgEQTgBfmXRqA3hgsRaqx5OAsAaBRlHll6rPQ5WevT5Kx2dZ
xYYZxG4ZwJh2c+hLR9IvkKjkwl7VsuwqM/3L9L6YEu39pIlRR9UAUyftGORzHFYvEmLG4pUbAaQj
YdZ1xohg6w7Jy5OooBlDDZqCbQvl2UGFNKgioc7PJewMB46Q8KWZ/M28x/SEjmtmYOXpSmnsw3qF
O/U0FW4LDSzcH+YMPoDyy4a9b1vh+hfY1MI/Oep1TCgRXSnPOzNj/ckpmK6OT4oPrTKuAFRUdD8X
PVomp3gIw377UPhLEZTs6ZSX6EtMHYH7nR0m5FSbMxksrF0ZbQNKVaxKhZUo4jycl/n/xLf4um1s
JIGQLUrAshAtC8gcK7lxkpC/YbJZQ/c1EuNyKR9dqR1W2y2n9zu1bkJ2RcheNUZMqQ0NnoIcY381
mi1gDyAtF8JEXxHGCaUUJBEs0MfrBzuILCgh2jhtqGgpCk/i04vH865dSv8AvOrueJlDmyutkISJ
UfN8plGO9w2/dGhnyixmD9EC22f7kvv9fW03LJR3SAS8ra1jVbZa/CLBsGEuVz5EOX4F6j6YqRF8
SIoED/DTDLTCV/14C62iEVGmI+a7FJQlHb8KJzG+LrLpFuEU6KK/9TN8S3x53rmMYL6lM4QiaV4i
pj2a+udlK6Ny7irciHITY9L4HqDdc/1BYWk7llEzb8BIHLc2RrI4ubuoECfKVJZGGpCcp183dRmZ
JHKIgyp/GeBv93aF5MVVWedA5ahmFWduX0DChFbYZhoqVyGBpL6Orj5qNd//4VQKV7esTy9ag6m0
kP5gVwYpR8T6afRFI7WQ2/1gSLxYFctvn6ZJkH121BM2up3GDKy5kGunXqPN54jHxtDPPckm1QIW
y2/39PvEW5XTey7KuMau5gpC9nM2YtWU6webdoNkOXIPgGSPj7fRFpYFIO52UgQZwY844LG/yp1r
izLrcLy4o6YKkaTF0AMtIUr7aWEeeQHTyetz1skl0VuZYAn7E/4LGn+ZRs+jDOG+u7PW0/o23uLN
Fc+8jyu4iL+cS+5xZC3pRSh+dxEb92YI+lCl1zb/K7O7TgxWY/cu0nfZ53UYlnbkc2RgENRhIUBG
OtJ2CS1Hmz+100lmmP09kD8WKugeuIELSdrXcKn3Ea3UXQNYlWhI0FQaTk5XLb0x1qLfyK+4ALuH
/vJXppyU+zGA3rrq9ia4COsL/qGP6DVrrCdnkoK377TSw2rHYUKMVFPMHtwO0zUHsQDtfQYiY62A
1P11H5g6p1WFkoLdVfYW4EAsp1rdQ01G7OShP/71SiAHaWLgrI5q2AvGwekTSRz4s7FVf8GONn7u
nSYR4ABSRE+g+ZUZRisJtmTqAYoTmjjfZzmSaa8ehIFAdYe9+J5Xhf1yzrNz0D1u4Ckywo5F5yvr
eI0xmz6HnJEtX5mkwRDYogquRGPpg1wnqiLPy5WbAuON5OrYeGd0aEjaic4cZbuZpR5heU5sZ4Ze
y5hwe9eo9Tu4/Pr3Zdkb6z4tfM69bn2V7zxhbXsbd79ZmsiTPjrSAmpU4KecWlgt/B/c/WJFaeOm
re72EK8Qttq+Ls5QbANK2WdhS3Qa/TOXJXw817sEi6R5+CzgHx2yKnKJzqNDHh7jiZ3UCMO8xt++
AcvIjkD5g0HJsKenbBXH+Iib3mlPnNQa5bfgg1ZvlzRh258eulrzyYNh/qWlb48eCuCU8ulMcuab
6bUPdCroXJpRo/hvYoooRAmkcYRnBzafRCNITRwUpRLdsCFYnBY6v6ek8nTGqKaK5GWcK/ryUTjF
ttCivK1xFpkD3Qe160sjvDkRJeD+dMc5U9AL1o+GHv2FIQoVD1/a65MNBgpqigV2N2NqY6MXKp/a
brcnwfjpY8Lz7kSpiwd6Ci1+xpoI9ZPtfyaMfLUT5OEf0AmH3oC+e90oXh/OlaQmhLNY4pMTP1Um
UuXUc11wfj2RFhpAmKk/hJWf43y1AqBMU4Naw2+0cNw1pmE7kALqKHuSbyRy0NLUbOe3pGO5tkuU
E6WDQrcRicRzyZjzYggNQRxtoSwI9ndLXrjqEI4l0ddyF2jgiNl9RZwl7u3/YgYhhwrg7X1iTUDm
K0sCDLlCkjP6o8yaDDsHN8t0N46J5HjNDMSfaRRP9tz1x9m5Yhdarr7tq0CDMKYHlz2nCvTnsmAw
bzQoZucZecHqqfZiSeJ/+IGk0fwV1YfwJ/oHNJhluDDGKq5/AukCXj0AhBUgAIF87oIwsDK6BY+G
u+zUuqYhIYGebRC/dDMvV4AjGwZ78k4fYRbqt3f3jFTbQ27qK0PNeEwAtOaCDWn5xZDdx328xEpy
neTDeAhsF1EnEFmAw1EzJsuU7186Z4zfAUFrNDsn7oRZwOHS6ZtVAND8GHdtw4J8sU7oZx475tlq
pc9+DToIqLHCk+L8t2AVUbGZESPC4dEvlM993Re2u8B5UYXwA7+ckgJIdaBKTkXG+lNDh68qy0K/
1BMD7cofYqpQrfhdULyEVUXYfeB2E1iMWpj95aqMXQDq5GyYjbzV8l696mJEQw6T3wTOX6U7oWaY
iMdraN9mqrkUbJiF7GEMmuEMdw/d/axaTf6yCp+pAr8ToY7SxTCkwRjXLHLXhCP7hg4kN2f7tDV7
cNmbuRc+mw9Z2c7E4Z03771AjXI8Lyd1BfOAAsHyO4CxJJTydaaRxcAl+JPxdGa9NhAwHBKfS35m
5llU9K1IZaEouxFBpJfN2dXHfN6TJCdTm6CaQINYOCc/WBZV1enJ4WllG2D2IVw/b4IGxtCEyEIt
2ni7mRvBiJmVvOIEZX8xd4176jUg49AfJGo26Q4EQ6goGIxpgCKnhCjGLpmYXxcPUuTfqbxZvAup
vJs0Y37BU2J9mcjV5vZtXdldnNCBJ6Suwd62D5uKGMucMXEqfSDPPntlHnbilyYP4FPuEE4SPeCD
ZgjcPxKUUqEC71Nfcau5ftSoBt/oTjwOvLUpa5GlhiBSF/CwXZghosPi5AD5aUrWl1dy5BX9cXML
RQBsyll14HvWHaDYxqmrEGQQNjxYn3TqeSMa/+aGxa/DIWtlBQn54iGNthnUJtv+pHiryynt4XeS
Jl9z/NMjFe+6rpTHUan43m5zwxRqHJr19h1d2//otHZMdmHxNCt2ZYk2BlQnu/I/fabYKl0jF7DC
Tibb9O7ylRX8smfN35sxiw14eKEqYaDv+P6rIMBSHLVKRdQ5SliSrHjizF1gSQ4J8HREAQPdSaus
9B+XwMnICT/OjPIBWCnPBBA3jQjXHMmvuhOlcSCvLea3qhk3VPKewtfc8KlC7Xang+MfbJDJjNTP
IBy7/wiq09crnEXIldArUqJRTYjOiPISS9uGJaKSHZk4UimXA6B2wxN0Ui4Yt6hMpmTDJ4VqwOEF
QahPu/BKEw4ccCOXIYLEVIYCIpopDKijeZBk43sfZcqsdtDahCFq/drl0wbLINsaIEhgxlvSOUvq
xYGy0CHv2mdHNyN8ZvlBbPsuf1WsFEEnUQpACIMDfQr5vzzBYgGa+ao/igJ/ul1up/v6+6yEcD1O
Y5PD04eR79sMLTff36hAGoexToDPiUUtDCD64HRo2ul+4K3/0fx6nyHrVZSgeC6/ccUXTT9iNgHm
tKP+7HytiufL/OhKPhTTp0rDWZSUT3Tx/93aiLhAULn8T4oK2WjD3ECDmt7vEcsDv016tZQLyZYM
pfUnlbfD/BbjXpzRceWFfN9FxVoqMOXTEypU5svDLL57iu3vYE1f/RH0k8FPQDAP96kKSGEYc0Dn
z8m9A5aP749IPPuiNdJ5Vr5WMi8cAEKCiB9QWkM6Nj1hF7/3cs2CQ1uhneCvq3nkk0zJ0u1LjLAj
zqGlRLeIxicdnMy5RRrwn5hItM72PaloJ8A+SBYFCN1RlQ63b2LaRVQIGy5K3DstE4mukERveR9K
MNeAONKReQJt/DHoA6f1/0RKFPiEsysfCq8X+hY9q2D/lSAjDXu9hzyQHpgXUyjzyHKWZrJcTtV4
FJb0tPoDDihRvSZ4mpPMWLfAUmhGWziN0iWbr6Yvi1NbRuzd/JVZXbdlzSQ1/QBUB7ng80EVsRCf
lPVGpo4YErgstQl5AVO0ncag2ygVZwRKhdNgHx3icUgcZ+bL6ipAQqVNAximXXzYVIWHTffyiowA
o6bQKQR26YBj7KOzpLAsuTFcCySe3OFUnfelPfkcUXl6aihpOa3MO2Fe2S0zR1sBAA+l8Pe14CSg
VOfM+YM3Q9Bi6PaeewcThlnQFROwpgfvH1STZuxwMBPAke6K+batP+LcV1caPeXkt4sHzclJxKhD
z5vjMAmd0k/g3oP8WGwnXFCl5qTQgQGBDrXSSskBVsNb1S0pwoxmD6+x3sR1ZGWhSVbzF1Chk+tS
bHgHAU7PcDWzYJU1lMyiZ5XC7HrB8IHazfpjdA+PHX8/JdA4d7jBsBd/HurWwyaDWGptyTZdKLF6
5pzD+QyaiX4STM1aINHCENIux3QLrMFGGQmYKCw0criRedahESUYaE/VJ6lMVPUSDPalAIAQ1RNd
PBCv1qnCh+FL8cB1stoLfP6kAK8pvZsanswed5W8CxburaPLYf8U4popvwR7ykhUHCzi6TFZ8xU0
LmKfCr7NVCtjhVVPePDlKvYQUSgrYFRytMCpnLpyGeaDZOl2ndSqdPoCcaLDIOea6SkAjqFdejOU
JRqSBOxSuI2VTL921PuIjApzN1G3grNqJLsu4/+31kSlVyVw51QyNTia/Re6deeXGJpfW4Uy1NuF
u3wBZZUqDVjSFHrzvDoJYnrT4cZe01pOUgPqNIZ8ZIIn23uIoZmUbx65Y8P8zVof0+0SHFBd6UEG
lEonSgukAvkdpwN4qVgzbY8kH7EWhetUuHIf7gxPoktU/wNi147ccLwEA4/luLrlagg//kgDYowF
uMu2ZvEbweG9AdOhHT4+NDopBCeAN73O6F1AQccek7PBM2LdMDgarlJT/ZPH3WJOPt/hAF/S11/N
Z3EwiRt9RnwajPm0F8LYbLS23LIsbXmg9Ow8GMpjm3RX2rj6FRpsbnurFvyv5xpJSh4e68yJbqte
7NZgIRAbatWjVQdEkmjFTE9cbcyFiYGnWUx6DlBuJ9OSEqFGG9nLu5eHkpC/68bWEiL+IFzWvmag
vcgGhFMVVvbWhiyDQrP/yoq/7XeWyXHDWcEKRCvxgAKoOkm6O7W0qdvW/MCZfE8I9tjBEoYltbso
2L5DvzrTHhSuUVFNZgtiyuvvH1xhGxzT/AqbX7z+gGHj/Oyw280/9dF6pRmiqy7UBabymW/coDWy
b4IvEX6JfUI8SMRgHAGUVpx6shfLEq2L3fXOGy5pS2dKQyjsLGzDudDb/4xLeE1/pCN4Z/Mmszhe
qrKMKSS45aH7zMy5J9KdQwONEiVUaF38cOlE5UZi1G+T0/mS+fsX0mbGVpFAjSCVNPxQrYVP708T
2bO/f7KX76iW0eA/eiOZSTOC8AfsEaLJ2iSj07o6ln3Zez+aMSoPnpVtmsbcvPd5QGOJ3wHwa7Xt
oaUJnmZMxVPxfUaVRbvhff9o89TVEkKNr8yhcRcqoYx/OIkw4+UyabQSjlmQg6GScQg4W18Ha73Z
GSf5SKoOkiLl/3qxRLOYzzt6maWHn3oUAR7BOD93uvD589WjNClYStAw/pbownmJ59UzOh3n6Yqg
fYwyazbynbvu5iX+29PVpo0bQnfrIKSDya847DYtBx6Yhbbq9yCCYU3kskbuiWk7wJdjDcFgkj3K
UEr/GmbOIr8kNI9/AT5LEyQNGgKoGI0obP8dlaCgMy1WT+yuyYteFSy+kNspivbr4fBTqOpcZ91+
tNxECypz6oeEdPLZTXn4X1CQhq+zsi3R67ixyGtkp8kQldo1YlVdEdzP/G9qNRpiDRXYWjOaDUoN
e2PEU72mPZkoIlDOX6vvpluNJuKN1bGMmwZb+nmy3hqYE4cvwTZYhxdayRkft7ZSOetJSZ2DValn
EGOhHqjCVGPlYWL2hw6r0/V5HTLo22NP7HvQYe9PSAJSrcQ0nH2kJzDPoifOOQHWdJ1wkqM4Hhfb
MsD8G/+AErheHcqnB7DbjZA+4G2vLwuzkJ4POKA2hzQim0CoHZqW4HUgq1F+rkg2R3PaCfYATlJp
y9XCpmhCunCwF8TeiFDcwa1PEuOS9fzXS508Uhv22Qp/g15/rrkdpHgiHrL/G5NpSmrdaqmWRKWY
9SAJb3dVFVWfQVdLxiopH/ruyuRkbXXCF3GEkrzWE1WcCMIphVp/2/SW/l2cTPM5Q/k+mnCgtUF/
+ycBxuN/xdqTfuVmjwpOfQH+2o5eX8z6FwFDa4tbQuJ5sB6EIMeubyU5w+0eKK327yscAllfi1qS
8hFXRPoyIO0lUt6OwVqeFMhUFlVbw3YpYVewugiIMVBWfrsrFLcXagu5B23OvOveXnWRfNAfib8R
9tiFwNEcVQCUseDuXV7ZIk8N/t3Idc0/rT+phvtCnF3mji/y53g9dwrphJ/dEjFRQ++2dtb0GSCq
tl9yrnH2wE6emBvLWj6vNqD2Mm9NNEhAd2kuEIsAhgoQH0aUonVny55v2qWfsrFjh0A9XHfs5kVR
BsZbERRzUFv6fHh1uXlnbbt+QucGB2LueVwH+9C9L8hhFalcsJz57osq+r9ErAkXSCX5DSikZ5qO
XqI/J/Vl7/Y0AOyHaP3RYBRdD6sbpJh7bZNWrngjkcWrsviq65S5eyu4t5pofTAs3irZmL6pmzwg
Ovi7cH9JznykU9m4UKUfJstT+nnYU0Yp/q+1lo7F6OzfJDD4ky1srNoxi+T/LDTUhDjnqvZlKT2E
T04OPStIrxE7jbk7h6u0Dva2itKkPyUqSTmEkzYA0dgq8dH71m3eFadM7OW3nFLvxpZipw1WROJV
uPTGcPCS8DeCAp/eBzap2teOEsf3h4B1kNWWjqkehMiNLWnPAsoBDmD/HXGWvPhKHbxKfn0V0qn1
87rp+jKZS8xRfuvE05e5dtVJRbmof8Ml1h2gB9fjLNnqpHkHoqq2nirW8expPjCzF5Oh9QQ4GiiX
2ShCzHVK/sZ65tiWJJvG046qg/1S607LEqUKMTm88mRlFrlFj1n4flBkOHtB2bv3XfCoZfy5Jde6
fvYXMZV1onExdK5j4QA5p2fN496iEeQhMh/TWNVwXfMSACjNZQ0n/F/b6I6BFnNMlenlKMX3VKWg
803TplzAhLFgfGjisl6kBAmb/SMuXmxgWd0c4jWCVDmfBUySX+zb1hsMFNN/U0rn6iFDv6+TN0hx
NcqSo8vpfShz9PSsoSIVMsSgPfooSFbOEUgPh+73hJBBtp636XQ2HiWVrJwVmZxGMiuLRa/AIVRD
xuwn1jzZJFESENWO5EDJPuil2T6z+5QFN0CDi8DQz0WBYaiQP6RfsHjGu0fBNzPw1uDp/SxsNDjm
FxujvByYvwADB7CRxVAlerxrzsKlGLjSGptzUEJAFoaqD/lVSDTY7d9gi/c1r3/Ggdt1aGOmfFaI
dqftBCRhoST/64DrfX4aN/QoscciniY7nOOBhhSoN2KRa1mx/soab2uKx4ZskfsBngDm3cLBMVa0
mbGue1TUwrLhhE4RT7EooouLm9s4TTIRFQr0JQJR2yBdQnW2kGAX9FQ7t2bFc1gkLXdq8P/72JOV
FQSIzqFPhTF0jCdndGNIZTfmze5h+xA9h4wB15KQqk5QJpamSnyB5Gwc17r9GvTp1a45YbtvcwsC
jA8CNxR1Q6ipjnS5BNvnppC2j7Sbg7AcPI/VZh9MH5DY2i6fZpc2DmmWKS6a9vruDKQTM9eNtYLL
ZlALugrup2TazVnIlzIMFfhsklcVX/BtvH+jmvd4wb3arRAE/yHbxmkGRMfvcnTEQkG9QEDUVewD
lLpMxmdYTcKg64WQjMwqhxrDNfl4H+dhM8TR5hcUaKBKGO8WbIOOfjxthjW/lIrYVp0dmn5MyShp
YfByhPYhZXB5CgUP4pFPTE26JdLQ38NWR7cktrgbIao3U/UpV6AMhk0e2OEVZclovtZuMzAMcQUi
HJ9zG3LCT+I/Gsbt/OEeepx5GBGlaXWTd3RUsvZ3fdmUzMmvuD9F49A1LemVudN2ra7SH9e3KTpI
GWtEOB6UPTPbFFqFT/maftzH5JHYxMKHM3xipEUHCYfsNjYgovkjl7Y4hIgWM368IY3BJiZO3Mj7
IzC5P7q8piojDwa2hoRkpAC//Y4nXDTtE+7uaj6lEVFAxFdIVhqrxNoKepJIMbBt+9clHdKLqhSg
9kbzgBEkVry75YPXtrccC6mjr7iQgliMAIm+8+g4OIGtOhMXQrPnoBAm2hF25gEwYPwmbxFkNemW
X4abihMAst6qZwvkRyyh1adGQlTL/C+vb3P3HwGjhC7kOHzFIZZjXxwPNokZ07kL7+S/1GlBIINO
wclkYIFYgvKNT74/7A==
`protect end_protected
