`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7168)
`protect data_block
hTX64IeLyHzfa3tJyS5DfurTWusqKnbnCjGoVcYRbJgBxbC/0237+CrXUZAYHFyk2Su1fOLuEcws
22zl4nSwcaa14XvZbs7wW5oaZw22FirZbRRg95fFd8zd0TBYbmFPpC0GjBWlEI4RkcHZ1xAQaR6w
5IPSDmsrzAPJ+3ESj/KiQ9wHIgIFH4BQod8s0sQViAXLXWsTiD7EdiJmWJc/s/dAFLoUxWjSPAV8
2q6qB2lqEUXbaDtCWL3ta7volhHRnewc9C/etfWePdCxCGHuEQPZddqVbp5hRJtGUCNBQSHYGFe0
RNE0eaRa9fxG9roMK6bw6CghFVtFVMcmwvLTnLhZPTFh8CyIsRDrjKopsW7Y/EYJHNrgpRKkpIH2
vjHz7d13bNSJIJc2CXfuV03GkjIpmRyWin/7hcoGKU89B3cposAXc1ztJ9ZrI7yKA48SSnawha7k
eCnwPNUqaO7vNwrNSoOCi8oPbFf+dkeF8huxEr36w7GQqqFwpS+WrjIvBqWjt/5mCEtKpH1HhHmo
+Bps+Y16LkhCDALFCArM3KG/17FlSx/e9R+qeDZWocenxByhbTCRF9qod4h0/dMYQryInhLNcNyC
7quRACcLwyg4aTQ0vzfMp9LSwQSA9WdBfGMP180aK743Jqza38q+3FeCcCcU3+D7ydVf1IUm/gLI
6YOhqkkI3m/MBsEqJsjAtP37eSn0x4lwl5hsISZ6SoKa8lYi3sRtxyIqkovUZ4lCQk1pVn1LaEDU
kxkpYbnqacfvJi+enybSCiSGt9UeZtpL0XkGXHLlfdxC3qtlMezcO7J4aUlAGBXkCc46iE3+iHmA
fKlf1OUJAPAZADF2nxc1iGHapAbgvC6NJErqMt8ZDsxnsDRqh+FiH586X1tI50XJ+auABVybdxM2
DTVjd89mTMskG/J61VAMseeyB+/tUeXA1wsWqkzMeyb3x0Zg9N0xq+uMIsrp3Xvfz4bpPPpCOHjw
yNotqDZZuOyk40EVj4cwa3Gz6DPqJh40s5N7Al6PObjypqdXjbFRk+H1hG2bF7sf41i5LgBV8GG1
e2uaIkwZAOitwvi8DVB5JI0TMX+OttfNeYXnTdt+rg4jTakNV230FlihfvHgRJNnL+L2KoKG2Llx
RSVrFejGFTA/2slEQlV6OJhsZD3b16YeZjNgqYWsRRdDJ+xSQup/b9GudFavNBB8vnEo2FSSla+Q
5xrKOyFJxgU6Sb0VpKeNqE6RCZIs9wn/UgTtU67/7lxIDBuzDJP4BEGlFTa62LYJ6CQXoxYZEOKJ
bgtTm8+/z4kIl+dUbChjlz8MT287ov+bPz5fb04uXUtzn5Yodobw8IOr5nA77xqkNnGSCeSGbK7b
xp51OkBz1SJhcrCLzo+mmizI/e6huegRQUWQMNpJxara1T3XvofnW0Co7MqruZH599Duxft4EJ39
VX43+Yu5A0Lvotl6iBc7tFooCn3qT+6ZEeeVI74AsHuSwL7zYI83z4Veo/1SxSaOSv3mJv7KyXxB
oPWeWgBtwLBrPkJuJVguTh3xdkXcu/LgFXZhzwcld0QDw3BY1qzYq8r4BRZ6pDAKOohTDVGJM+Sl
BJAmjECqQIIAFIFDjNa/Mer2rCbISLz50+Wq4J7XV6v2u5KIdJGKi2YLeF6mzSEEavLfkTgqpBTZ
X3kIZjyOk4DAK5wide6fRF12tdM5hgat4K6nhhDnrb0EMQO3f/XGabeybOtSpPQKel+nJQWl71be
KaJLLfM2SbGGEmhK4aWnlsiLiZKgfCWJhHk8YF/DsuhCQuBcxpB9RnJs3oGeaet9OqMcNffrkZfe
5tsTt/eZiRJy9K+3DwyzhLomKqNoXsWhBTT09CiQExm27IVVb/3o6r5vk2icVpgh4a4mPhbbQ/x4
E40dyxtlOjg/i9H5l+IMq3aXxSvtn9WaUxTAArT9YpfKB69DUSX28SPdIPeJW9VPbLbCBctP6MqK
JrGYIS3/MEC0978wSnADBUZatF4pny86lr0WRD8bnekC0CX92r18r5U/jCgHVWxpLmEhPP1KfJwG
BtiwNCu5V6RdPeHEP3VsrXDYMvVfFr8ZrJt/uUIBsoIS/dzJNI/qc2dpam/HNiMXwMNNbm/z5ckT
7bPTXcVqzNe3DTwz0MyM3CYajJ5Ok+1aDP3zrcHowUPoFTIFY34zv+a7YzEX1la+WLNewwTUb+Ch
YLq7W/uj42MAzYJXBLn5QDDO9enu4CQrF8LK8SfG15Yel1GyLf5MdOMRwokrgyEfwlYIWscnzF1w
QuDAPOYfNPWU60ve7YY45HKL+z8Sz3AzWbKkUG5ZzjPr5sQo3YjPqtYYntOS6OM+qs/678W9DlT3
Qwx/jnlV0QuJYFwiEiBfV3bbENSCT4dvCDvBXVvv74mqgYH6/RxTV9Ilnr/qHrtJQ52w7sFkkJcb
omQEb5T0OLY3m42ViIJg+9REWq+hIPu4S56WnD4GQ3sGMqcbYv/NFucoDWrG17FPSO7MqY6YR8Zk
TLzi26Zz2YbR3nnVXsTevP41chZusa15f/3cz3QQs17xKfd/ZC9LsD/pvhHrmYin8+lnUPBfP2S0
4isIhZtm3I1t4PgHZRDNjvYniBxyiR7rzloTE2RsY8zfef302yt4gYj/rEqU/ZvTQURHOANbPLas
0DnXnuZ5odWKThrDaOWMp1zlWeti4vDRy5WmjZS+v74Fb+Cunc+Oh8v8Nl4tqKYkcl9N4Ili2v4g
LxUTmICDABJNsj12uxlBSRtT9o7vcOzNzK5bbs5W+K2pNEQbnq590ZFyhBRRjeMFmY5yASRyK2Qx
hT+Bzg9qkLwTxsddgPUP+Qyp5nbTunLFDulMSmzr+CCv6SlYmVuyvXQTdxwpW61zGZnwUkDaKhLf
hlzlQSSze3l+sxwoxsSvHAFthVSdUea4YYO7d6ro4vBshU1ikx/FMEQBvd6CXSI63f8PKyLC+PzL
N4SSE7wdy1Zdv1dEeoUHrdCpM0+WWIdIEp0Hch3ivQ18ChbFGu2BjpZKaZan3em5A2RxXTNguupF
l8O/KWIeFpA0KkOlpKt1pGa41HuR0EhLZaK2gEUix3g/hAm647Ah4tm9OzBSjlCWDCqOqNH2Xi0t
Kb6v4v4IfmlbsAw8lQyMXwygWPCzWOqWIkFfcd1A/ubpA+FldsamA5peJuJaHzYfDZkE2dgaqhOG
NJnojdKoAvuq9oxgp8KT+cS4lZ8xezUS1P88hZQ9dRb5wwsowpX2HVn4RA72zrrq572xMLNnrMzc
+XQangwo1fkLB+tWYsy1FtjsqDNbFL2kjgym8MW3Yv3rdDI12NzWUCXoKoJfgDZ911dxaGno7WSB
rP/cv1otofWPUWyVNGGkdKwRu2o6SdTIh5Kq9w4a90iY9sf2nw7VxmteBJzgJNBn/DIQJz1KWMFp
dXfFPMf9Tjt/YOeyMymVp6CnT8cHx70odJ2wa79CeY1DLj7bmwyopP4HnHHiGKzhFWjESZggPrCY
FPzMJViEwtcIAw+2ALNjoG8Sd4f2dXOJv9HHupARM+hOe9xEMgmMnsp8d6IiRVYlWNNoYGkcxx56
a9vmxSkA68A304KghHzyD2lWgZhzGqx8D8JtIw1yx3GhpALBmmUBR/SC4fLisi6eJy9zbxNRLId/
KMXrl9ylOmKQgLhc0CkE5cI+cyeMZMsnokw96TgxjmoMLfc7Nn5ka77B6+xUYS6m/NP30Pye4A+K
qCMwK6K+5MLH8Blw/vPWu67maLkPYAWO+n7rbPTprTIwv7UfdeB2kGHL9vagPEQl6B5D28gpZn/Z
iCP9fNiXs0niZS7w7WAsxXs4HR51Uc5SGuyc9NRhrqYiq15P7R138oxa3RUo7s9EhYSMNFokaarc
4KsJAuoaCrhAF+haPlyzRZPekTXwcyKRvXhs0ywLAQ+n6QQV62UDSWluaDveikZAq2sHWQaUq8zp
pEUGN5kYI5Jxw8douxdDuFajL/vKEj+TDviPksA+8l+fwL6qbbEDYhaQdx6jjFGf/InMFuzZ8SCR
FE04/JrifFadZciqrfz7FGBFhPunslm1kaK+bYYaKkSorEhe4h8AxOGKDOCgJTXHgHC3ZyS7aVZN
E+Lbrtg52qAkp7sRRD7Yx/Rcm8hews5+b7NQCS3HMqWE/CO2XohDC//qWMYkie7fDY/l9vjZh9pI
Qcf8D7FMjm4QApYMNOQO7XpyHDKWNn/adddp7tybc7HncEc2nC3fa2hREA7nS+8kHoONQvr2awzF
Y7dRREuIizvvT2Ar4+ZZ1F3auI5UB/xOvpwzBUl2DB4KELKOmygvdKcB5mrg3VUR8/il1HR7Phvz
3SPVDUFhZqu1uO/j/ojKlPP1wycDLvJAekZqOaR5HJv4nzndSB52z+S+cLQDDD9n/s79w+9sTBuP
0HDv0NHsQh0R9OTcI4jvML0OXMiUe7K3gFlrjfFURi/0M948lgRg25s0av1rDSQvlukyhaHSpPN8
mhwW1Ibrsdy0xjCmQ1xPOmzFhJtKxETNY9O29ADQCbw/K6HYq/6IjrnuESjJZBr1V1RlWcr2MrfE
fDgh2U/vOGoeAK9bhIYuh5+aFhUtVyDbNyoWY3hopWV1BYU+FBUmhccocZ7+2mJ1SQGUcOu5sZCX
iIJGodhdPYGOh5WIP8OzX4z/6B+lQRCzVK4KA3oY2rSqN6cji0CGMnYju/1deOB0WDuM3EwyDpyA
+nXfo27Fr6DXnJ3qqVaMyQRJ/61LyXC29s0C35VdwPm7cN7ZbTSIAfPa8Leqc5nAvbHaZKenQPM6
wq497RJj1SdPtp23BPUdgFrpNyqVfcB9xJJf5NGMXm+qCKGrF++RTJt+ykgZO0OOE8GVSJN4m/+D
umXfy/tYh+iNsc4bzwVWZdNuiG4wR0AfBhTwcBQ9H/SlAItfREZkQ38785DxLOVnoH65cdBpnzUl
ideeAuKkHMjh2IVHkhRJ0cbATIK9Cj1ilqH9y/Dl9YzoO37Bd6d61V5/yWr9guww3J5h6ywqO85R
U60pfYBL8V6vrgsRMhCNr2VmELOS8ezjuuTWjYunyeH6Oeu3yuiIl3TNVYBMYM/WMrePLDpHINfx
JKJIsEPfojmaVgNO698AlSTia6Nkk1PFujEQQ+ddXfK0/PPoW8TcE/w+t4yXbSwOWxeuNIsELmAN
owdV9nVCe0TdBwFrvDd5a+5g4XShkj/9pa+lld2sRBq/RlRLI2qIT2LEoJmwzLsuuWeLSRCFV9UK
44a9HE3smDcl2lqfzD/gMiE++NJGjgOkKA15Xv6HDm9UQi5tXsZXf485Xt43SXtb5pZtd2JXFz9m
e+EOqRCclaPRcBdSr8oz1rZ3RX0o6E4zgFoYBwhyA7fMvpgHDT0QNoRIHvK0N4RPBt70S6nPKvhS
pSIzKJBPX6JN54/HUCrwWtutQhQT6wPOILP40YorpbnaNmkIf5miKC/1CzTkWtfmMoUTz1VdPWLg
gP5OGeLg4NBsKKCJWq14zDTS/TIkg7LHiEd+hR77aWJfPUtHr1oyy6BNlxpCzcPf+bN3qkCIBMi4
CIIY125mqCqrpfr9Qh4tZI4sn56BVkeV5a1lPUqBkNOFpZvWVDicgMXAGwN1NbDXBKvTYZ+oYpn5
0cZwIAtKmSgFRwGh6GmhCAIjDtxc73wlG9/X3wjeGRCSPROs3DWl5gOiSbuvXxWtJ56Fe63xIYa0
2RdrWVkSDXhViJL5Qx8/5L/yuCiEnUaIQFrSD+Pt/DFsTyniRY65Gn8F29+lT0uAoFyTMSq2epHj
i1zkk2oPvPTNrsYZZapwWLtRm8dMW9Osr0xW0YGLlTCZimmKP5dOyyiHicU7y1Q077wkJ9PaiuQi
uriI3C94/BdWeickLen3/LAEfJm0fjvfUELZTixwT28G4hOiHtH6siBqIkUOpZilYZ2ZE7E0CXYL
dIh1VpXU47GRJUrnDdNz0lhXmIK1aQHX4dMFU6VIFbZ+udSfRRRR5OEDAm9hN3jwLLqPP4BJyWEu
duEIO6AelFqlOFmsvBcS4Ejdtu5rwOUA7J2KQ35m3DpJJjCZ2u8B00Ua329ylRq9VlQyvvgabDuE
rDerQI2koMzwxDT56kBFHvrqpR15fl5rfx+E1PJpY1b4Ft/OtLCId7/v5pX18yq3wTvDUwYVNxhE
o5wExDGVEJPSjqODOfmtcoS8Q6BfNpgrDbPnOdSP639GKHxMRD1q6wjEvFB8hsLB6mMUfVfJJnGy
vr6K6hja7oS66xCYPFx1awZH2NuofFSu15FvaIc1tNFenpYFfj80I17dph/0ecRsLU56VgImpQsq
cB82stSVLOVKaEPYqqqEWhnZqGU9kTJNhfPuF0AhmF0rw/GXNtCAfVB6RTxIO2JDps/Xwhmpr8ZF
/4JF50jnAKT8sruDw/Cn3yQljR8BBaockD+p65AIT6VYTa9VRzBfSk1njjp2IR8J+SBeSNESY0Ee
6ipBeO96pbBK0O+8H6z8WVSHwUnsZeokWemDRSHJmBbhPAsR0JDyqIRpxSLDLktAmVr7+pTQHT/d
8ouH7hSJTBNKQUHloJHQKhiU1aeJEVzwxsW0KGNLwrWjA1HkDyn7EqVZ0y/qsdpTmECfMeQXmW9F
vZ2H0vSX9Qj2Il4JJBw4lvbJSAahmnH8p0nflQuAO5zf3l6kDv+go5C9iXuMOD9n7j+24sYW+Pih
BSdcwiTKsYDJy8N1AiQAzXJXjQ9jAh3vhBtaOTRWSEUdnOf7N9KSiBT5dSoGO+ZZNnj2etBZMea1
whTtthno6OTW+fCUVJylUbAjHniRQtKP++ZgDWR+10TcHgdqeOr7Hh8YqN5PVmxiG88KxwatiZBE
BW2j2JKE82vTeaIUSlw0fJdNnybmtyQzCUXBkrFT2BrpRfhpUkwGSP71jZ96NP13g30Yk8QvvZFL
bwuiJuUXtPT69esJ2oYSbDvPEdW13XaMqsqZSL+1MT3j9KV2x33FL1+g24UrMzMDX42x6OC6k7hU
cuqBl+diHGhPLN1Wbxeb9cH6LyheL4oUM8kM3nOinNT65G8oYmiHBNwJdTkwgQ3yMYzgevoaz84q
DSmChE95nwssjYPaDAmxB52GCb0ZrKGUxNRVHQHMXEbiQxa4Ini6VZ/WjT0btS2e9NUAZWZ19PnE
t0OAaYnS8bT+IIp8cWtPdeXra1dnpi/YVUYbSNtqrtCQjc42zSvbLvbOv72gAIVxKZJE59C8ANZE
10t3sKu9SNCH7E4SGO1Txg+Z0jZDd2pg8u1QIw6JujMiARfDRM6zN8Bx5lXNM8rCuNwbJr8S8l5c
OpFuA66q0UaymppildNXo/WWo9XNWKWWBeKc9mNbwzWVOucuaGnOlm1LJy6F+KJPrLB7CqEfupEl
efIDQux7mNQlP0bVn2CeWIZL6ZIutad4vr5io6tEFi/XBXze8ZrNJdqBsMtumccKE3quAuf/KZo4
NPQ+RTB+b6bYhZKBqldsm4XnShXHfCLhtTjeY4kN3fzqv+UCTfoSaFGxzmX8b39LB81bQjP3RESM
cmjioZ0wqf+5sOHh05hXK5b+TocJe6WBrcyAWZ7BflJMjCvq3q3TZ95OlaicRsFm7b87elP8g91A
Pyyky3hY+TfIUCw40ty8z9vDjZkPTDBEVZ85Cr8lWecbws25CBsljQMS7kI474A+KsYMIVsVjL9Q
c1ie+Mzlk73kJkStzALupJbeC3LvBYHLdZ8yI1olrv/y2uVu7ezoUXTGMQHpf8gC9gVJw6V9jLqF
VEE6BCKftpQWmh+jYyWjs5qs5nQU6MkFOSyDgl7d5L7vCAfCmGIwR3eZDNuRk16LD13NxNWV37QH
OXMzau81iIHwqBJ4btfk/d1njzv3Ub0augC+Zfp3vqSDvv0swyqOqjIvt3XCmp49TZpnL1vQJbQ9
wUZSnWO++Z7ii4caf2fBHaWY3JqSqHQYFO2edGdYCWsvKZt/XFTYDbK2L4SgRnY6QhAsn/IbLOXy
fVSMvKdsZrmaQqvs2pR3sx9rRS36352ZKq3tcQ59h9zxJfDUvTlBfYC30WFX9UK/tpFnWKXhM9In
x8e3jY6ZX76uoyaiXjLQ9g4VCgP4yjVEsIe+ps9Qdn4AdVe2QZ0/ExCHWmsZ9WY4rb4mHuyKK0s8
K919lr/zwgwnhghW3p9WO83Mketcb5cvt60I/CJhYMvMJaakOnFMWVo0mk5ZsFJc0S/1IHPVr2b5
NJd6anp+yhhSmlEwMMzg7wjjKmMQ2OsDIrYn6tffauOkyA87QYOvWNPG0lKk/6Ce4ftRRrhU1ApC
xjUlGNP3ZAx7ivp/NVZ2Xjt3cJuX2K9kZ0It5XZKAx5CZjCszGy8q4bcWRRAKESSb6OwC/Y3RTQ2
8OCxCDaPAFx/3zfAp0kZK6uGbXgicvY4p/5IBXOjjI2U7Zbj/0yy5CxbkPVvKyKjUip5xF5h4KmK
YdpRXm26BPK6DRnilnZAd6k+iaGqvY0L9QOC8D8b5oWRP/zTi1GE+8/HvcaLVNrkaO8n0RWUGNgj
I06IA26l4Tx5+So+HdP5Xod08GSNhTmpTsMUctdkuW67n2vwalmR/og0DNZr8O5hGef8v7POLleM
CQpbFCPA7g6ltPDWyTA/k9ofkqT9uY8w81vZzOm3udT3vh7u/Hbz55MiJUYFpQfBasRPydsYRnEE
qcIOk9kgA0iEEJ9DIARYBoDc0Xn+OfHkhKORJmHDNW6WfZE6+mR3iOVcGOfgYqi2lWDuiKPrV3iv
9+aTH3tM0E4c3b7STF0aFd0nQXJ5HSoaLVKBAo4rcnZEH1ux+tqQgpXsFDPLe5CxNdfN+TQzxE3n
JLfvsWgEKrIm6TenvZdHy1M8o9QblxV6kqVJSZCBGtDEZYM+s6ny98P3EItVaxm7nCiPJwXoXrvm
WyqqFwPvIwNO2M2W3AUWCxIJ3Zabndy0bwcyoUSzCxF25MVkrAQO61fmzOm9HBUWAk9Dm4m/84KR
1euRcoKuxyqj8VY7l5l++rJXYx9+ItNaVcTZIl/bLjo/VfcMlyPU7aN0HwltCO3vv0qRl0QjI4yT
P0aX0WpFzKPHezemQnX9a+7s3Gmv6ok/uR08b7/gIaRKOBeJ3FKFFWoUkbhtKiXFO5W1tFvddPYr
BpVrV73N9NHv2AXcBxjww6Ulxh039yOzLY3ewsJxxwBDJTw0PFrlvgzkKtRO11HxUU1/hwAz7Sid
TrwR3BZoZ2QFEnbCA2wlK4b0CtUai6/dYobDtxo1ogGyu0mx2vN3Q8YzjaAHWtk/b9hHZUEUZ4Qw
epYUa73biXU0mP68WS0wI+NftXRqz7EYX8nfyTrWSLuJVlELACfJnrTpgm9XkTjCnU8xdH3TuIyQ
OOfZnMqwrA7h3qacbTApLx+j5AkGvPXrVgweplJsop3cQ2T6J4K2q0KsccM5asqtkRsbt/UgZiJs
HCFqFJ80dgCDn7CwKRRglqiwDxUqG7cd7p1s4bFK5E+6Vg6vtBFOwPFl3bO0qxLjdVOSNB0DfabQ
6tP06dYuVTC+Pa3eHAuWfM9Yox9zhvGGqIvtXJq37AxC+KFevE8aqT6AHQ==
`protect end_protected
