`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56560)
`protect data_block
hTX64IeLyHzfa3tJyS5DfnCGfI2VwUPJSF+Bc54ckFyvAd2I90/gLhJIdZrX1uTC3SnHPiWm4BsE
evblv8AbeXGsZICdONQK7qvk25eOmgP858uyTTAJe4j2e/73aoj6J1krcMM/abb5UucHsrMTgVxU
UvdLBUcTtwx0Ya9Tb3sTZ5+iQvuU1fcKMycKaF8GR1CMo6+hJC6xvDxSJRYnzcUaz4vEYPgtCZKx
rvZb1Qo2wvQbGCal4c5US+EdGr+J0q67fCxEGcTsXO3HzZRXX3S0xSoZVnSR/hgiSqWxyXLolCyK
YArTdeBEnHE9xmxRJJjxcMpw5RG1WOaIJkEsP313CS6XoPKj4I14A0PFTK+hWV53djzkFbvN10PI
jEJ+esd/N/09Y0yWICLiPStPh/JdcVW1bVfZr0lcUsMmEVvSR64Jv6Lb0M336DNAhw/b0/W5t4Kf
pmNToJbvd6GDPTMhGVo77JpUxKH870sk6RJx89Z/gkChDqu7t6oC4mpLQd9w1sL6AQz1pFUN5p54
S7+Hawq2bH4HS8MVQiS39Xg1pkvqjh3u0p4tWsrO64PL3Xmr5nnSoQk5Ms0vkETFgdOhDmzuHTFY
i7o+W2SdpqxVJHpRnCqPcBqlasa8aVKU9++vSIN/wZbhxQl5Bwq79mi9OJbJKKtuepSqFvqYusS/
Z1kEjGjxmDdfMKRHXlKxjYxB/DzUckUZPfYMxgZ4gVKqMbcyiaMZ1GVfXwcw+XWdLfGz9NXOu+HZ
hDzbWWnFqS38HdH1j8xnm3lwA4j7dVN6tTpzUXAUwNTqAkHp5RfxIAwbRYttcTMkN3kLPPab0/w7
Wd6JHV4c6lfl4zMp/BM6AG6jLwBNKZZA3huk8+T2uuOYcLMWwA9613q3albp+P8bM5iSwDu5Rcol
FYJ77b+7KWCkM/FmU4zfiL8qc0kwk6uIRkfy9ZFC6SriB0lMfC7HpqWBtwMiGJrQw3zzhjYbfwfl
c9pf+vr+hIQP+qEzbm5dTjb6PuXgdl1DfEFVXdRXpKZ4UeDl/lZpecMvEV7NoFNIE/on7teGuQ4l
Ak16rw9MmYeU5W4LmJyn7rcpJmiPVLGuBHKBWhfntj2F6CMCQl6/7KHKj27yLDdJPdHFpxW60jhV
aiAme+HiaVNenwNU8mEo+7GqhMtXBVGp6pvUGgLTCYldMH3hIMSxgcgukyEJ5LjrpKYfZEstngfi
kaAHR2IbOpw2URWNZy6mBoHdFudIwHPT5GjBsNd7h1LRhPgtIBkTqsMnVCUfTemA6e9i/d1h87+0
PuhHpfQ3KZtwh62S6JqNE+VHb/AtNDtejsBgTe3KV6Mdc6XUJAIPFEoX3xEf6OsSa5STbAesr3GF
xJPrQ0kEAjVEmmc5s3j6+hIoMmJDAa9ex1dWkRkNdCuxgLy/ua/+YJwNGDgftb1XOr59eHdfqqnV
Ce445m99IeX5F4daXIdjbNcIA1iWVR2382FLakjy0+ZokbBx/acDLv1KCr44hrgCMO78fhJVni7W
usqTdgf+zQ8XNvKXSqWxicVN8thK7K9s+od7gT3pX3MWyUbCO7zSRnMNgZlmWfgPLntvcwVi++5S
Ux2LL3bK+uCIFLNb4p58UWRjj+D7M75Bt2dMdD/e2cqGkCUzbULqa6X1/8Ha5yrhmS6gEReT+kJV
/K0vjVZHE0mqfxIs24SwwBBu+U7s6TVD7kpbY6mvpQZtpqxIl9sasT3bVpzC0KFw+z6Iz26WxuFP
rt/gh9OohdpEYehNe7TCtVKrhZ37sdRwiJ9oJkRIVFu4hWs0SnWRYhWaqoGtH6Lc4j8SI98Teitn
HIfdDDhUsfaR7UBBKm1gVD9cDjMgbXiCN6itktn90KA7NW1jOEXOsvRnkbUQSfInMMcsNDsQ6UPW
EFASL6WmGlCqP5mLO1CYXCluGre5IsnntvvXHO6kwvD3gmgK/vUpnHIdfPkF+nrCIUuntvFrm/iq
eQtYymLKpDhHJdqb9iiwsSo66H5oI9qLi68aXn2BKDTKd/Rp0AyIc5AizKdQG/ms9j89YKoxVkW0
B/6Sj3f7Da82ivVgzOtRPgM+dEQgJAYMYtR89QR03KruVvWbj4MgNfwS4EFurfG0LjhoiW6r43T2
BBPuFdwS7D2GZDG92QpRAPaGh/hbjqG5N6VdDzZHRNVoolYZXOkAcpu0spg+SPCTJMIHsVLxW6Cs
28gOY0nL02k8kiK9eUovkLjF4/mA6cccCb64XGoMyc+Rdr3gTmVXq3xXS0Rnpl/rtwIDXGUh1CSy
W3UYON9MUMkhs+rIfKXHGvKFX41vVXLNSK+mzECjzVEEWKElTl3B1234+Zfl6sfrsN+t4N9Lvhd+
AJGtNRNPNuwgGRElDCRyCK0Vt1i/JAtTCfji5mFjgClNbh32zMCRf5Str6dqODEZ4htLmXm0+6qW
lJzTPVAlRyEtY8FiYFWKgKZX9kdMDMe1JwBHWV2TgVqf7T7e163PPot0AQqRMGxcro+8B2wrKEbJ
NGYRmKQoypLFfzyAyTfR+qDEz0sjCApnLJ0IJTCQidotUphwY4cnvCNZzeD8kvt7TxwGa0KBBMZM
062fI0yPjbk3EZHNhMZD+dTckAP9aSRQxdZQKFrVgdX0FD9e/BD5eGkoqJBXoY1DCTZyHtx2k25g
zknc6oLGpv1vz/RVG9FGLgXypf1M07yOJUtkxO2oTphNCXH2hcPH0jZtyfvHF1fyrGuHyoGUkKWU
syPdkiKWOtjbvC2dP6AIS8NM2feHdZ3AMiWbcIVskaIu7VxkKyigBkFFY0rtF0WOE06So6pPZugK
N3s+tw2bFndUHLS0Pzu1bShGb1sjoGlTFcM18GM+EbLuROvr7ncigp4GxOzPpe9imWtTMKVCESua
OwB4Fd/EZedrQ+uOM02vQaXLK7Jloa0GgGf4gm3w/ldJBxoj1/9YSnXvYWeAVRIm6vsF3evZZjLe
wiLaZgRFKi5sqEmDrFJOnq5hFSOR7ZQnuyt+rYL58laY7dRiNQxpnW+nRhAGqTufXm0x+Jzfxlmg
NgMWzz7QxRLTG4L9O5IzvAX17hWb16+keusl6fxTixfdzBSiGrclR/2EXpKr9kQX7bxRWHx79F8m
9r1AqKvLg9fLzowBRa7gIZrD8m4HLt1mx+nEga0w+QKE5rCeEMjD2eNI2oZDrtQQrFMEIz7q9wmM
zcGHGrlwpE7WFomiFqUlMzSRaznO3kxSaeRE4gQNKhfECYqlQzzLdVyZ0sk5EpI0SQfsFZAl40YX
rgia7COEUfjd66Ldoly0CDzAOdFyR8UbdPS045Dx+QKp3ES/NX+xkDMSRM69/iFvoo44NvUX3+vN
H16As0E5KFAnyIPtybKGwmJUpm0CQl6unHL/8DOZGk2a9dBRYV/5h82gTRXfWKop4c0p7sQgJx0E
n1WqY1jl05aFE//jeNXAA/vovuVoKwdS0PK5F9zKzQAqgD4iUWytL3Eh0s561fzWlIG3JhPJy46t
i4iHw8Q991eJKn9ToexqKKBNVfnmHB4ZcZ0YkFSrLpej3hjMKOhRCb5lkBjQNBL8QfA7kzxKe1dU
K3TpxmXNsWNRZ6a+CAmT7nxKjvp1it8k03bDf9N5wBitP5y/WC8tslXWLqs98EeapMA6HOAH9vRx
4bOWxjXFiMKT7QblouXas3I+ObHvBtpV1CyZixTTAU3x8MeNHOgaBVlx8sMo65ZFK6qc8avOm1sm
meVdrUO22Q1j6X54mm5lkeGluSYG/Xgu2H891zvokxXSvUDl18AYiwCcq8HEk4jpZubxQwmNv+24
HToclnYSfjmSeUgmZU0jfUnRdT8Fs6hItK8E3mtphszARqV0nMUdfRGrTh0J1JpkhyNO4VzhpNOO
/uJZOr+P3Pmf138JjXoOGG6WuRVJzIatE8d/FhrcWjZy98G0mTAkxgwkk/fneYvPy6pmnYocLnS1
UXwYfOQnShQYGI4ikjlYxDYXftk6WNxc4ttrSZXIzWiy79CbgQ4R20mnc369dmXV1dYZ4/nWFcql
dfC842F4lnyrsLdAp7iwmnxxsTiKyoSQQbqPKe4S6EowK2Ee+YlacScHFp6voXL9vXcmus9Bi7Xj
SOdjZU61etAwNDWDt/EaMXqUqx1+Vwl0Bez+0cof+D2oGkErUlEOpNchLa7JsqwGzBQWB9rK2BLp
gFJRGLyWpfPICDxiUA6PzrGFZM/L/vOTv10+f0skuReK6Kod0RITWNVq9o/425dK3tB6FmS1KvNa
QU+yOsKplRbPnLlQTcUAM8D7u7GLATSkUDDHaKKv8vdKeHSBkcMPNSJ6m0wMZpMgTz5zYxNPwkYs
Lz94NrsRzlDpHk2a0TbVXJ/DPaMaqrbyUv91aWs7vp/+t006Y2w/PhS+Eo1WN0rOxJGjkh2GoLcb
yMjCc4rDwj+S6fyzZ99602ZMiAe+z8KQQoPKYntB95SQMtfML8rXevPtF2I3hx5XbSuNlBJxmEa3
3beSH0rD1HLZDxlAcXdSA7XN0g3hA7ySnP9xBEBSr+PTFmzyMTLtOgkHpp6xzZxV9mLp8KVWPuGP
DCSm5duzGyii3vIfTiHFgGbGgcPICawXJZQOT180Ub3GYvIQdv4AzDuCSRr6jHniFD/NfqDoOvnV
LQbltL3hZDvm2b/5rSaLmTU0VbA90b6uRDtF7S5g8YIeBGnma5N/nkkKdHwxhbmsGMX5EhScyHQ1
GmGSEBMfdlkzmgih/YJs3HfpqQVs6FX1bEpnUX8dXt2fwdc+uI3uE2j5obZWmElvcxF0u99Yd5kO
U8WRef55fmaRq1WQ+frTh8B/i8m+hkCiI33I/gRIquowXLi5QXG3m2c+72Vm+pF2liIkzaRVxvuH
4yRlZp/SGTLTLCF6U6qctlTzAh0HbFVZqjwUcgmOtc6357Dmg9RvmlmXTgF+7kQJfaoI5SFElv/O
rWJBcqYah62qhEsAjkeE/L6wAsevFdjh8lsKiezHhlm3fatZY9NRWG6mJPtZD9WpWcZ9/421DN9B
EENtu3WAg9FmBEwc6jNmgbNweEhmaj1C8/jbi+Tg9nktdQSdQ03V70afjGXf6DMxV5JpZRRTCmAG
k7Q/pU28aKGOf22ykeZXH4qun743fswr76erwlU33NvXGjUw+zXY6w1IRC/nxMibfeBqWZUeU1ys
Vcxgqi/+et5RFec7pxcix7MxS3gZbjaGSHgIpPHaKcqw+UjVOm8vMx7MCpE6M6OARign/vMcvsdY
C0b5STeOV4jgwXrslVIfNqpIK94oD0+s24Ikaad1ne/s1zcZlM9kWdSoOFmh1bFizap96snic/t0
ze7uZaHIDBKc8LL/vSnQabQEvKq0fkYthoOigCdW8BdIhKltQEyVJEmIZGiEdGUyojg9DyVKjPoQ
yn8++SEU/S6+uv9FJHzwemdGKCH3DzK2PCwOWs+7/WSFUjwzuBDOmFIffzwO7M23e491p/YAvWFw
yVaArl7PYDo2xdFuDsFMM41J3yIXdSCw9EYCfOSxV0bdNWKLfhJfEi2+NNJQsLxi4JNWl2uSnk/T
ZEIAcSGGXYW26PHlHGviAFgg1oQeyrKoiTg/9r90mG9H75prXLL6zWutOF1KEXwVP2ZNn2Zmdaef
queABUm9fpgmgGDFO7VsZzgEhlAhwQt8PHBGhzfuxQwgD/et4u7KJoKmBZnQwH4TSWC0kLp0Zla7
Y0qb3Jhh6VLmeQJhpRCZnuHWMw08ReXwsppB14UDPuLD29m3Ow5zvbiOI8pjoA8Vk86mp5SmX4bv
FFTaDhCLLH8UV4ph+wmuu7g00+UqXYTn9LaSbFNYjLcktndId0zuDg1XDiOUs/jtdB+QCEAp/zbV
VkZW/b5Bu/al6enxgGdrs7wXQt+Mwj61uGXo9ceP1Cg7kdkbyXY9cuYXi1U70L+5ehqfnpm6w/8w
TBDPMA7E2cQbSlWq30EH7lZJVj7Oj8vmtbTmM0QEB9HQmvF9Ojcd0XMWRFWYg9N4HdmxNWHH87WB
rBkqS/3JDLEi4i9Y6yn07jemA2mzXvDECTcD5+VpHsWgCPWGhz3jkNm4xzlzEKhf2vOQcrbdKprW
BWLARM2Rr8d79m3XCrqOJ8rF/OeExmwBqMTExqZvQDeyJir2fAFIqxmBncci6JgJy4axYQammmYB
fu1jWW+r9GI60j1YJw4HR1rKzrHhvNEOve3+PzBeECWiVWfcasXLB6xN9NFyr0dmaCOFn8KCGtwE
FzrS7u4CyQApb0mKPNzthcPsc30f2A3zESO5qycVHIUiCmQPbTWMmWOMetdlfpNC+tGbO5g+1QwO
4P9HFAN524VSkiGXXot4xGaF9SOXXouYnQJmsBVN6+gmgesgijzp4KOTcdxTuHpoTOCKOUJdzC5B
oKPw9ml9Q2+jMIVizpXHX06K+lKLp3jrw5f31F/Vukfla49xguaZRSY92FrhNq4LdKJ3toXtkjCV
+/7HJXE0I90kTKBOuQzLbvPHcq9McscsACpTfE5l2XoKe86ImlAqAmgeo/+oSD2nOxo0tsuoig+h
DS1ZKMc6qX9yb3MPh/+FuRpKpV62K9bs82Z2pomYJomtI8znyEs1toyuV2pJRf0eEg1xSxCARV50
TvqZobsfXrVV5r0dfUgUGWg9tWVFb1N6w32Vc9Dwy6GYBKkXgO2L98RwkcQySvX4IDs6yM6/2Ly5
8oGIOROqVYpZmT4J/vne+6ls3aIYotQixqs+dD36WDYuOrrjXeIWidoMek8v36aoB4vgIhb540X5
r2apJ1S4oDHBZ0ToFfLulA75fvC5yJ5qrcde2i42tbhyEARCIxV6LA9k99tcC1MB9WEV+ZdKDr4A
Aw13DoK5en3amcjKMXX7qUCZY1ECpltWNEVighIhSn0VgNgD9lhELCJLhWNupxAzbhgNuO7AKxFe
jcIfV7KCFnnA6C6kg8bEzU8oS7vpKt2PkqLPTtYeYJFAXoCBLgwmpuy5kO2fv1z9iOh2JzmiVL/r
9Qq0xK9MbueJggChX11OYVtSgNVQi/L/i0Gg0R4VHnlZvodgeSBdj4C5nTTnvc5wZPqzcCTYk8JR
fK5c2LFAY+bDTwLXnNYLJS40NGRe6/kTKrP2xwXrs4AFe5vvj8WLbLrB1fXuf4XDElv3am9xi5Sp
4vBlQ8R/Tu1LSQoTfD2d2v0M6ikqFYy8EjFHvxS4nGn5IHIqAiKglhu8mDvAfYztvcddhMW09WJv
vdvhl8FlriyG/rQVgYAYggT39YnFw2x6dHkVn7QfCQC9i1thSoD5HgglZdAF1mM2zSLjkB0NmH+v
lT8B0J63U/eMMcYJ4BQEHd4jvoCFtzfLlwlGktFNzUKh+st0ortkuPhwWsqZCTl7tuwgma6PTt/H
QeEiddAjt6fg1C0HFZej+1K4YrE4CFkj5txQGenaX0mLKiSlQ0k6KKXQCyxWMZF83EPt6WuEolWT
G64f9+uxouVVYqfIH38E/o6t/35wl1wtcx3cKt+/Did4aYA+WN2Pvk9imKGQnZRYVVbamBnyK8lj
tV4/QT/VOpwUZYkwTOjOuubaCgu22+Q+xOzW/5XxMhVugyx38czMvFxcfUGDh+wLMtMHmSivjIQo
vBiQCx0JoB4ZFcqj/rfbZOccTZKsbJvSfRD8VaJQwO9evlsPTyVUmpWoAMhCj19xWKb8bbLWtELz
9lOKs/ZSg1k3ANqkZF/AkPfoG7uXw/OZFKB0w+6imgCkJMkjcK+QYVxd33yB0a5/OiM3UD/Bv88E
+BsQpRizlqPgxPg6q50Ye4AdMTGGBO4g9I7Q97uAHTaY7+THjIRd7waXBVaB1ojF6RxCwxk5tXKk
mqmU0/GIGz6FDAYPe1d9wuxkYHsqD743yosZ4DPE2g9ozaFC60gInurgyMzr5KQ9qmRsF7gmB+u2
+4NI7BwpQf9RxlJY/OvEBPjoRmo0NTk1nJ/Nl2gHkuIHWNFzTnw/c3vM1gnohpVR55+LGMRrsIo/
OPBXaoa7NnRq2HPbv5nTh/SwYMwXYZmxvENQpwLqdmIA34D6Eo71Qs09OJCTf7hewHwU7607czmm
N2ETNs5uUc/+ZEscxq/zRFhuACwj5KIQuTlarn2Ium4vtbGgosb+JSOw0s/6fer07e6KFaXi1Iee
+HTbStTwNjgyUc/Frvlvr4XqGAthbg5IFZjZivdXK2jyvqhMTyC1CRXnOh3cc5NzVAyXKr1OSISj
R1QyftltJpjmUWIo9u80yLs256UIutLI0+TIZzzlOzfFU9uI+7MhLsT+SVEo+Y74tQ743SHfctGq
iVRg4PcMZRIoKDpuEEYPKG7hITHqof+a6h2GWFU7WwoDfLGDVX9jSCcnRq3ihheRJ37wrq1qb/G3
YadOutl0jBnBQS66Z1TYggGM+hAtFs2VAqAwzkULomnR8CVfCNcyrkWQPFkNq1c4tkEfDeir5IYU
8L2Bxh/9Ngd+5M7CrWLKAnohVHc9XrkO6nHp2hRbYNI9Xd3yHG9NDix0CquC5FCXJCGS/b4U8OH+
h7zQ0nEk8Nxq4R3FcBZyETMWFVC7kFe3fbJR+rDMzBxxHRYdBjnZd2hZys+X5sUotN/fcRa5oHSC
aVgQObTU9HB85kX9RFQOaIwyyL9UGrao5ZIobQyZHLHWM/HxN8eBX2FYriDMnDtERhOhmOM0D0aP
TY5fIHNIqpITalFbrApive90rZB2Z4v43xdN21G0qGRADbBSHZ5tvdFa/f3dSMpFit2OeGJGDhOJ
lbKcORI1qQHkw/jvXS7H9/dtcW8kX/vETMhhJFnusQbECyycLRG+vXmwbpG9Zt6j9joJqOAmcU5Q
GzMjVaNEB6TUZT9VN+2KIo9RnEvry06E0A2MaHqrRJ9RX7ZbDbbeBVSeCu4iSdKOsBCUrvEGz1dY
YUdZUiYR8tg1eQQTRABkczblaAe31H+0gD5A/Pikfov8ka1nmhDyM6aS67PNEEyPUG5kPkN6HjCi
sm1xrYIebF8qFy59dTt3ZXslbbabuOGyH+jJgMou9V8IrU14z8hWLY16I1mNr9V8s6jRF5MG+QOP
TaQw3mB8XfqnZy/MuD/5YD3z6Xmu30SO0kKLMKACMGPGIizwgl/CGJLrWHHuQCdPbAodid1SmfmV
XjfLbdJsPAQlPHJc0ijKuhdB6etT3Y5A/hYoytkPFx5OEdHf+oyTPsaQv/nFstpuUZLm/vCzCCP6
nVGWTGnqEIWazNddgQttLw874BKFdHs4/hKEZ1EUJxRVWxedfjXV5j02BasZVa33EFkoTjBcWyS7
dh79QrXr7kKU/B6LswL3iUv0Lr15hJmjPGh3CE4E5B6B3MIHn6FFpnpK1wohdqvsPWsRfUVj/Cut
6VFgdsAL8IJwK2Ar8WUrLAUA6FZDLjw7ien67yLSlsbxumLEtv4tpoB7NmE6dpp7cmZhPT2fafUT
1gLock37I5rS862ux5yNwWGOk8OFyxkEelJ22wU4Tp3VMazWbwpOleRRL2VgrtzCdsQcKhlVl8dC
btobNDpDZAtkK8PSE4Oh/BRG7DcOpOuIU47OTGzMp87DVBkr8qW03GjcDhAuY67T8dOwPPlbTKEI
VqYF26HeGEK+Ui32+6zBUK7LfhACbGFRUroElHc7bkqrTEYQlRurpiNfITEwKY2li3q6f4+DV9ul
IQYQvjgaKOBu6CTa62kWkiQygM6P836GxbL3K0NiyVk4L10rLkI27tuuisAn9PeNn1pSaYteVv8U
Z7Ram3Bs2uvFLXQ1xv2c1wuuq3wh7TO1o3J/EEUyMzwcBjj1qHuvHauFXFx5H6dql99c+NVbhAcf
955PS9CDdwTn36q6xoEIdljaR3CoO1VR8XeCW5h0lmbg8bXYZXFmjSrEjw2XiqyWnJliDrvrYSf8
eRV00BdQNh+sIo79Efv2AKZVG/p3NJWWzAIFnErscno+OWUMBFc36/VdII9RYlsUD5JONvQ0uo+4
jeOR8Fn2lQjocc41o03fgxbHgvyjssQwO+SdHvNbtdRXyS7XJmOzizMS7ZBd5Su9/ezW2Lm01JD3
7jmnpHrrqxVJ25oAJZMKCkRlM4UEO9HQ+sGBxQQVsPd416PG6tNcRVNMV0fUT4VdOjmIAX2dmwDl
8MVsGh5uBeOPWLC3NZS1klPogDCZk10hv4A/aUGT+eraLyTotf2CLB4/g2aKVsoHj8bsywdCQ066
u2M0Jwfq6qH1wTD39DkZBnL/q3+CzceRCfIirC01gOMtlITBocA89mF/QcsxBem+WJ91S135e6AW
7OKyg/SuWFAnwFkNmV+/HRNwwseGZZZHlHg4yN+2QrQclq0fLdHlf+r83MoDu2fnHK8iIkCvOOyy
GhdjhH54lI3zZdps+MXpFw07tj55D+PNFFHlHMDv5K3YJZLIJ4cSRvLy34jrWQPlshlrXxLq46zo
CxrtiidGHyLMgTc1WNPIBpPhW6uPIBBLpbaQjYto0ZxjPKl8nGT5uccqVPa3Uys50rpRAPWsb85K
RbjFNNBCI18AKLTh6ht+i5mVp0EhDNHUBD5FQPjVNdvL8QjOcWrqGPOOi/NpVzAI4nVLqeMT2qQ0
CYR8aIYUc66HsCxNY58w/Ou9xdHWD5ZmhE++3sLbZ/kcHW5lOYxVgo34SEjNWSdsRqBur/oPPWY4
gmw+5k+vHGHl2e5nX/yJZY4crhomo/Sut/bOs0AxXHCZO3tKmZirxA4io4BhOJ7DGI3ZdalC3nCc
Kfzr8nxAwYuv7bDfjCDvTuBWwjBXRoj2znu7HFZTTbQs1Yrzeoau/vew/G/Mp4rQ7NIanVIEvBFN
64Ro/qyF+Y9YX08wlrv0RZ2tyjRBDghqiCcaq16UCjAXjKQ8JSRgSf/eQyoPXCJDD2cHVeYl8wkp
I6sCs/PtipTdIDtyMahVOQi2GITtlskulkE+v75rPAZls+QsRusKmbK1fPnXTs//RYvu1VnvgIpK
8e+zCQqNKDISF0Q5LBUH2s6Q7r0dBSo0Yp9ZNo0swN8ocH6Uq9OJ/itUxZ1KwUXGn9P5QEX4m/TH
wnDjVoKilWuiNwTYqyDy7ZZM9tTtXVtigy3HpTf6QYNPJtW2Uj08iLnWW4rR4L6qVLNO/qxHpDjE
7qcj/LBPjfUD8pZqAVyx5HaV0hszNqbZcNDDKDc/KBnXNkFtZkNLummldn12xBAsNTsRseNyWjS+
n+AB/TDYu9YVbGzYW0x99xNY+1sKduHiUTrmdrMglc7tb4yRVC3MxKp+vxvJPm/uTFNYWGl8mZeY
e/3lRbKLqQnDez52ziymDTpKvMhpmrGURNAum/HKsmKD/DdQdqK8xuqHefzLPs2wkZS/7LXG7bfV
/Yzp817Z5lrC8RK4YbCDBNb8gxeql3prVPBwQ3xpFePFYCpdOEL+HWPFDjxv/RLU4ZLk6Ert0RJR
ueZZQaUvzeXt31jsUoPXwIOfdw92zzEU9YL/DO4ZYYyJJp7uJjmq13h+ycUSbY2eXeuOGdKt/xJi
kx/NZv7rxblorQC80MynqmD2HlXvH2BnB3kED0z8KNNkkiEglf4FUmUjWYKMvT0bMrMHuwsQ+LRs
oUBtuv/Gvkgd2tWC05VCGkQPeux2h/rr+YQQNSayYKoG280KHSoPTHqU49+rxIeTOFSfUqUrSYJZ
4kAXFYf6MvsJsLD7p7dhzf0xyy3H9cjBHCxFDEMO50jXT8X6vCHX3b9/N15GzvFG5d8OookJj5ei
EIQ78EiJfOa+yKsOafexzX2RZsSyk5a9RxAxM1S18lb1BZYD9L35ngSlQ+cW557iI/0AiyOIt6LT
A0CYkXb+Q7dxOqCWp0ol4JsD0fx7cVxTazQSJJB61QUg4SFPuFB3rpB0y9FZEEfxW9CnJfG3vL8c
R40bw4wle73zy5e+YAoR3fw+fCKrWF4Gm4Avy4Q+4fG+yMdgFt8nrc5jJd2X5htkSi+hcIXIeaqf
ctGxJe+V1XbgAiyTMZXwlrCt2wONCZZcQpYrZOc9zon/Svc2y6+4YWT6A4dvAuH9AWJwqvoqAhTP
V0WXZka/78wPoGsYCDhfmQIgPilDhX6z/yZiHT3YlXAL9t5XKw/7P7++u/Ek7vyCV6R4v9A13i9C
S7fZv5W3tH8SgHf8BWyWdJwIyHWaQSasTNfLHi6IhBaE08VcheKgI9sEAZLuNgW+JKEb6W+ZcKso
syecN4t9okkkuuk25wG2uZG5QsF+cfpy0Y16awgd7/3Fug00P8FK8z92Mh73/Ff04FG87isqyUrQ
gJhS9jRHx0jHDCHvmuVpGWVe5a8Y3PQpGhiVDPUDw3w50xd7GCDJ6HtoMyF0lDHmoW0fk0e3WoEL
lQJ2qqvmtXYjDp5nF/euhnulens7Rol4JI+DNZQ8X+M8NRNw5MG/BSReE10bkbhjA6AOkfTKFKik
MF2RsSkswjMuxuOTDhcoHM3ZOuak0lJOYTq/cb+BeC9B1ufbT5jKeGQSvUtpoHTcVknCYX92mXlS
QAJ735nwlyoqLQxh74X3F6TOSGLgChqEVUOwhWtD9rxBRruQiMw3+T/TyhfMnf6NgFfjaDNAaEhX
Q9dK3MU24In5fIW+E5BBbOAMGom/gv+FU0Nj9vwtIVgS+NDlOfC39iz4jnMMFx/SgnEpic4IvXh3
Rk5ZcP+TbCaXyOyNZFXJ7N++bIBBD1gtCfOyI8UzvybVpk+KG+3MzrGfVfdH868IfiAixjLhiJt3
WYWCxtLiB4UEuCXvNDAPRShViRfeFsmKdplCdaSTkHAiLafCi9YP5nw12YeSEcUIA26cYL6xi2h6
25McTM10hOaOyh4UKeGvkDmICV5+vQXT6USXmC6XSBH6fgQBIDT6e21irA4EkP+59gQno2doZeoQ
NB2ZfvuU92ezKsGwDDF6TnU3zhE6bzNI6BklIftW0CXIlo5uCLGuHDyeROMddz9I/6bxu49ea5gh
Gtw3VECeeLY9Jdrkv7/09TUVRpYyFms3FR3aeix4JBAIwKsi7TmdWEtgSUosfvT2OQ6EM2Ks91L0
s4ITopHjpn/BV8yZtaqcWxjk0tu+br6HmaDUILayDnnMIwr8JYUItSuPstabf+WuJ3n0urXsDt5k
37686g/jpxStfZprXPg7ExUylJKBX+FbZN2bUhONleQMj0+rWq2tN5uvQwjzPHkJcvXByZA7bllS
Xg8StLE4nB8+YoeA1F9YqD5M/NdSq3M2dPK+neO78ApCmuVld1YLOwXXVsYk6afaDwsoc/oWd54B
B/T8AWgit+5aDW54ahPhEC4qia7rRxOUXyjRHHcn/6hoFMjTwP+iUjZonqhloQcuas1B9i5ohzWz
C9JLxZqPjjoqm9xSP0ENelxBOIOE6xPA13t7PJ1pAENfIPvhkxHgu3qeAlsz7FSIwyD3VDMbPlSp
EBT7AjcXCMEFJaCQg8o5+vu46aGui//lD1vGIRfbgGgkmzAfUiRbSdVvhWo10YH7k89382NxBjld
gs3E8B+kKCQhtxga3h7i+setk0DXfs66I+xF34FdKz7FbhCKVkz9xEnhTF//hsk9Rq8AbzuqGn4Q
Ov3jNub/8StN7KzyhlriSbsfC8rSLAXWs7QhMFMMB6CvvU6bo7O/Sf0mprbi56KTufx84mQ+dbD2
tXzoogrhYlw69C6eIn7eQBkuJb5bazoCXnZ+/PyvaIn80hoOImYFS/S9oq3YD+9LmytyeQ8w7E10
c+Q85hnkkwg8ZhUrKCpT5d/FuXUiyf89YzedMP4YF1d2WN4eM9P/qJ7uLspl/Fbz2UwWqiLrMvpE
E1lGvNd79+Le4Qqqw44oR4J8mhZQu/UnkXFrNJxL50cFGFpYtnmHKcMYDavKJBB4IyevepoYXROi
Lp4lzdnHYqUHJS4eStCjcXdlJshzqEUOFsM7vJFRcrH4olXESecqrn5YuxOCUpKUdFZZNOyYJFuf
Ny2IvXD55jp2E8M3pMOU6J31Cic2KdnmBy3317ktI+sCWrrbsKyxisSCd5Ko4cBzEpLde6OuDw16
gtzS3XxXCO7wYOJ0mNWjNw6g+0kyautvNgkjDAa+jXkcRm7eYSAI8sTFZGcZx+ow6o58rbPpRB1I
W79OOAdXm0AlUSXypQtH+T7KnL6KAEIphq0bvJysTiVtMXKZdOOMoFRd8c7rbjztDs0lMybsER+m
SvyNixv4sBQQsVvHMXfQEhQVCPS2Cduqq+NETwCOecVUg0oi5RYOsupcwgaM2RAYJfi0c5pAgCUT
WjN6reTvtCvvPApBCd+Rarw1n44klVGmLUT8snYA5opKZNrxUba4zgSUxIVrQYGWn2GKSIGUy6j7
xKvLH7yG2LndspkBuhLb+MjrmzV4zAc4ogfIzBQ8xlH+TacbKv8MAn7oJ/eTR8xnqExg6h9M42BA
cP6Yn4mhKTLPzwkvPNRxHCvEqGbxKGllgdFtBfkopsInAEKw03iMWZuNWH4lFmNfEeEQDurbwzLn
SuK7xZQGiTU8wHzjqvBMY/CwOm/4WAHzeh73kPY2QcLt3KX+PNotSRMs4zkk2gQb1RI6vN5v53v9
delGjPwJZpgjMjWIcY1mk7jzdyHQpiPG1QeZh/gd1bkAe5ky8bxWxa8GM/CMnZbEzecTuUQp1maB
3HtwI/nLdsgyE0B7gWtbsfq0EswsmnMy4u4tMvm++w7u8Hb9TZmuUNjJNoGtY0TXIs0GTofpJe+g
4UOLK4FSFjd92gkoUYA79YMMC3XUrrkLuNqiMsodk3gorhmsC+NXrn/+wCoGlnkezDLUpL0taCsW
riTxsy+5fTDbLGyVQ21BTFOnUyMEBXxamWxJEGxKSdeWA99oXzWTQdVU6K7zUZuaIQJb0b+J5phc
77ZyKFTRj8X9mIHaG7PWmP9ir90Br6WAZFNElbz8b8jKNxwXhAp5Y+Z4S62ba0myoaSNezi4QR92
341/f7hvX8ZM0rfhVYNSdeTOvlccP1PoL2Ih2lv3I/vVws2zEnNl4yz6RdkCol8TSjMhIy+S5IXR
IC7XBOwxWphjz0oj3qhSU0mqy2KhudVrAz56av/oFDsXqLciKLPTfmGLNsOFB7L3t5HmXLYu/iO0
jQOrPM6WhFYf2iMkGdzVOkzKKdET+5WWQQ9UHW8KxTwaJfwmKTnoLfixcSrBzVKHl7KQkV5r+fo0
p3r9BrgW23LUTlWjvqNZZpe/VioPizsf5mpw0LjSVLRKHnvbYiC2oX/KpvyDcirtCEmcTeiw43iQ
hyLyW67vXoEGMdFikyq08YRe7lNJLsEcVOR0Y5wCgl8o/GuXC9eMOC5K+TqpRyc9qjv1wMfQ1jmb
6SsQ/egcOVo9hMsmz9X5sH8sMYf2Pi6oDjCLefixv+0nXJ2myobkR2s9s6takk0pelJUit4tFA2z
N8m4+STht9KzbVpU37aiVPzNLnbRvusHdQyheJSRIeUAjLEB4fFe98YihBUgrbXxO1iIa8X7zzbq
SCzpOikKQmhmu8ZWV0TJPC/H24r5IdMPKoFOhukuvz562aO4TeysHnkAKED+ARvnTJl6flmGZW6P
Cf4X0ZRVrdCGhRC7PLV8us+89jltVRVvJoWjCFfNsW4ypINKZ4GrhUrshiBFLFS0V/71zeGjRXaM
vY1dM3U1K69WvgqJO0a/7ptnwSnhK3M7/NHqtYaWBIEwJurNtnrELC0IcIxeMQlPUd40vI5pEgDA
evxGXxSAnfSzyzqGXE8u9+pumlQ15cDXEctmsFjCRRqgvGJdrKKItsmUOOiBDAFDzmMiO9D9IMw0
4jVFy98U8UR83XlUHe5oSYY7Vikc3WoIdsvtN+JEknL467t0jqtdWmV+ZzmyUkWChMq4ZXASsY1O
aDkniSlTIkug33nvtR/yG+0BD+wowuFRpMT1L3z4l0RVei8w1suo0Zep0lVvFsPwPceywW5y99Ng
ZYIPHsTKvAU1XM34WVJs+H3wktZ055a+zWZsbrwdb88vtWmcjiOZEHi6QNwNXHb16BzwFqdO8X7s
DiY57nJVzNGqxlMgsv1iRpITWrfx6WMrIPz9o8p7zz0yA5whFr50nYBFqpYSFgAmn2EM72YfDxOY
6wya81hJJD4ZnjX0b3pK3IwK7hnndAeKA6nN7FGA/l08FyTVdB4kZNW3f6rEq3Zn+KKCJwDX3OVY
Wf5L4CcbIJwH6jcoipg2nKIdco0bj8VNX39JuKYjuHsXDUoJmYlDcBOQlPSoqSxMkxKrx7OsFUfh
TZCbGAKavdZhtkudTmu/Pk83Ggxljk9dtn7u156f0FWs9dLXHG49wKjVjdhnHAuA7XO/f+KkyLWk
Dpp2xh54EiaNhFvAec0JxalAz6wK7Zm4xULPnZLlulM8SdEAMJF8uNBujDSa2Se5yF2pmQRV1JCT
DSDl4lDm71YkcXO/TiseulWJog4ad7ThyGk7SqnSAenMZUB3MONNSqw+CFZdMP92KN1vEG16cm5+
M19J48X8KuWqEhFqeqbh9AbkeCVIpBJAHJ5ihEcAFOWr3aGfjReal9vaWSh9KsZsCVYrCjBH56E6
3cYfKZM+BpDEPilyNrTp306M4xO4mt3mtT54loSXBKsE0ibctJ8KO2NcnbaybDuDX44cBUhAgO1A
3edaFzNkG1zUIPljJGw+nlBCRefGgunFiUGkGG9c2KbmcnepDB5vDSS93KcJ8IXFuL/AAowSmomc
t385MJCx7EabIc5qJ0HHfOLFv4KfqGvdyJmjILJTm9VFbB2iG5jgjUz/ngYdxEdY4nUETWn1/Rwj
+yuVr3t4Iw0kcoBvtYrCM+vKvZacBw2MUD4VU2lxqPMsFlkZOkTNC/zxI0ofl0MaOyOEPVxKlaT9
rPDbnB6xa0Kq5q6OLxNlZSLC7BUmBcRC00iDgm6UprqYJ+ZG6sEzagSLlh/BUXVELR2c/qdajoHR
dJWEE2gX/W0KC9C9QFkWIHmU/nLg8Y9AnjXlcnfRwdhbuQlBTCbIiqMvVwD/HSaxXhzlsxG7/YOs
zTKs3UCnGBf4xPiomwpGQ6Ey6b1MwM0yNGxbWEujdMH9p1lc8yZ0v+0oRi0FlGcctwitGPePKGdy
1Of2JL4NGahDOAcbL28IhgEmS81bogBTe2+j1SxehWAEME6lIff3hPuaBP3NbtJ+2kLIHAzNhINT
0GfQuCNixxsBh7hwoEpzv+FAsRWEWMFGP8gggG43TBmc3lvq8S9Sl5aZYQPJhe8YwEjVtw92Npuh
476R4MXWv7QYeoLTz0R3wxXhmD5DJoskBfJ/FAy6HqeCHlGAkzgS024iUwzrYcfBy27zWv7jQKPL
4UyGNlhBURlqFROyPOH0OVj8Voc7gDKOURhHYs+WVhU+HeBtPhM06irPitYsHjdo9WMQqblMmLbi
pOQQ9UMHiy7oMtNLNEQSB6rAFUbbfLrwRXmN9YJP+vktidjgfhhPd48zrlCvcxjzqPq0TUD7ZYBU
TxMw4IAVHPDzJ1PpUerVH/6RBsvzXQJeIt0dESjKu8OMUDN9o60oK1P1OmMualsxCeQ/AVqOTpev
8eCMe4YL6I63nW4P0Fif2/vHFPlfRihCHcv9pwzUw+3Y7ZXGRTwathXhVarVxj4IkZXGzwWIPuS8
0DqxbWwBBKnkJHDgRvvuzm7VKu3Ui2JTsHgMS+jsBzXSLhM8dCpIZpzPGPgfubma2mfJMofl6V83
5oI4Py4gLrJO8Bz7miHQnuJG/KsUoWuDPEb/+MXMIs38LAdDDB9GavQr7abFq5qKqkqzLa9XQDXR
b/z1OTmw0O78THKF74C48OYSg7lIx3ctemXoyedKD8B6AHZxbseUcInHMQOPz+WnRainhOClVGwf
dv7vJEZIzwNHgAo9zX7erLKRmzWj3qCyr1oZcCmtQLNQUJNmjir1cuKsXX18YiNnO2dKliyHnlFl
804umi1JUuZvlhbPWYzMkY4am/oetV3IRFWo7NgllYZQFf5/wtji/F6NEAuJpzgjxKxAmuhMO0dt
EBJmPompXhLdV8+gd+zJ6QVjScqrJFO1ta2GfYXYp2UMkmbdIfT+5YUc2lZD4ZDvcRCVHIOhq14h
/8Ur4NCnLHLoz4B8AYaQfGci7OPwP5MIndD+0UfK6wxs9kGY+FeL4rrYxNB+QoANrVzefZA1olio
BlnAoVdPepCaKIkYRs7HYr6mlBljtr1DtWYaNBVVyRdxO5qpjOJ2k2/rJPwckPapUdNml8/gSmta
8KPeOv0rx04TNc4rUx+Fm783dfWTo+E/G4isJk1P53BWkdEBfv95sGA+LSSGe/+jdVTOnotCxtuH
U/UsdxcWca/dh9ogCZMlpZP7Rcut3ekF2PwUzlZwv7TWni5DkFd/ofv+sqAcC6fJsUSMZs0hZGvH
kBnOYjiljralcgrFz40TOh2ZGufAMF8CHQhh7D9vKB7P5LwQXkkdEGonhiYeBXhVRHGApeq6hhB4
/VeehAC09hIZLVG2/0cuUQ8fc3N0A1AIcvP5CnlHF8z0gfoAnQSZkdFQHQTvfJiTgAs6h0AaU2o4
PyUxtw+8MoDGBO8g2Lwc9TWLod/9ztKxSGL+0g7SrN2gv3na6ndTcMRQ2g9uvBWZAfSoKb9Dog/i
7VfkCejj0xyMaN9V9rVJ3wicNAYzC+ukduQGQ6EOvl+dC4wm2tBoA3MXz/+utTFx9o3mA4685IRt
tcwRDCyJhDkb8mT4B3dgVj6TbbLwR6i71qcDaf/cYcyvh6ayKS5K6ssr08x4D4oZUwb1MujIG7f/
1jZxPKLCwt6W47WX2RlhtbLNEPj2ExbX9+bS4UemwWHkag55ZtfzzNA4Hno/9Q0E9Dt1OE++tqlV
/4O4Do8xw1aSJXzMDM22omleyAXupfIsUr+WavS0wB016YC1KYCfquwIZjW4TIHo0dLuZR97m9Z6
MAm6N6sT+lMVIpf36SZ5ClQH2hdndpJXqHXr5hch9ALMxEGMovJz+mMpZN0rS6SCR6t6KkWtZkgV
nTCgvN4KZ+jO6r8Yx7Azw3msIJsDoDYcZRl0w0B99U2qJiHijs4GvhXh8xaqGJvrXoypxZKmjCpi
P2HRuUdStOVIeUI2/CAGgk3QNieQXpmCv29Yx1cRCzVzIpGuOQAK88Ll6s1WZzuArwCRs1Pp56JT
C78UykNUj/hgDp40ZIOa+H0Fdiw8aeQGmsav0yXrZTN8pvxLoOYyShmu0LC1bTalLZJ91e80cmOe
5YQnKfFSMbI9pgzBHwlRO1zb7CWhs14ev718yKZ2Zotb6I6kbtUfd8ZM1WwWQ/4EDqWPrpfIf30G
euqp3ltANm3pxXqullpwAmSugE0hItTN7mzbnd8T32yO6rx5IVL5OpHjB3F4pZAeXsJt3sTcXKtF
sbHvKO0ZUU9CYQvVU9anAKJdPIaAYQQtRjQPi+D3b4UI2UHf9x28xkScGYGTB6XyaHrjtTIWflKU
F/O+BeSPIV+WOlTZcePRbRHmmI4aDoxXAhkMHJ5XXfe5Tdzf7qTVdhwU4Mlw629aWMQU3JLt4yyu
fCGasZ2ksPRwbxYd6K81IYVZxwTcC3gOA3Bgkg5VDLxZYJO6z+WLoEEufCRcP1c8wxZHlg0+ZGOy
Bt98A7OBoXAgnZGUFVDgzhPnkIPFbtyzGXaVP14CoQbTYebJv9Bk/8gtgWdBa/dcwWwLM3y2i01A
fbeuHvMCK2E+Ff3QwlxULw9ZljBsyxIwf9VyGDKW+ywCbLkXv7SyvfnCbqw3FbvlgQk33yOsKHmp
tMWeUgpTDBoIlzqvAnRCOG9pH4vk9pJ3PVBEFCuP31Zd/55xF9wWXiLALNh6ElHQsYGrq9/jZYPV
dOhTZSINvKUylqE7ydpZ9DqgWwmgthuxNCffr1/qF7sXJc8sgPPVvubSuz339FYwVJA2swBKPwst
EmL2OrKHQZPFpbd3VdsLxoOGGpDHWRUFcITpxf2BRaEe8kvWMP1NnvMiiyIvR5vDyjUzRd7xhFsn
/aRFQ3y/kZhT5AdI4fl56HgmhxwYT6SxVafZnqBCvOmElLZvEII0fYt7P0hNprcyUEdtd4KIZSfJ
7ItNGv3FuDfaPpu94SHOAKYtbkjNrNWsbDlh1oqPC4av+ZHHRCVlXUjqL9u86/sESF+5ODbKtxQC
gI8/heDtm8yE/h5XOan/dC130uadDlRvwfG8EUvcQcxixworXdal4nLvU/JsxPs7jBYyePFI66dQ
7TnuowrATPm+bdl3RrfAnLIUfBQUzBgFmOEHTHv3pe3Zl1Ew/ZYB/vRKqoZJGuBrMyVSopoP4EVq
DxBgBLT58LFbgcseOtMo+lZIykAizXtINuAUTbGGUTltcikzaNvx6uRFlZ/ZP0ymsAVkXIdRPcyZ
nlDSeOm6tcXfRpobJ+MyCHO9o5cAeHgL93gHCW7COodyS8ljXd3zw33lREbCg0NCkxcDkDWnhph/
kI+gKlbGdhIqCp39R1sLDbj9J0tg0vmfECdbvtMssAdIUYJXhGJP7WZUls+vCcBVgeO2+ToLvh0o
rvkghQ3m2eG86mpo+OcbhvU4c935PLXX+0lUA9elPf7vwQQcknTYDnhKGajXTIqW3OXet3Xo+DiE
HlscSXlQLlECJh8tUXhC8ReueDIN7C61vX2wecO8ycwS6kJIGXbRQCY0F5RfI4ZQwmD3ceQGlwp3
YO1l7O6kpD1YIEdEkqg8t0tOw6os23IiAWwpXMcCpZNtYsXa3gYvWj95HysopSh6/0E1hZbBEc08
znGdbN0uiGe/UYJ0qlHPnbsnK8xIeQZ2Kb0/ZhZc+rj3FvyydwzG2DEzdTwMtLFKiH+IT7l//dn+
98v4HXMJtbaLDzLkHNk189qtk8fHAUvI6a4NbsFz/ObEICnfkqL3GsSIonNssJ3zsgft6im5gsVL
UbYQN2S+6+wHwA7GfFts26YAmPUkBy+G/Xx1ZvmWVmMMNrsEu52Grryi09yojRwrjl+BOudiqnXU
O5b913XJX7m4FbVjLGmYdD3q3SpeDGmKnBCrxcuCXnnPOMP9i+uZf2nbpBYZIgCb1V8Ebdk97x8W
nHnIMvTHD+CDxhBLJGo5XZFTv2StgnKhf3uxVFjerFEsTLrJdHpD/Smq2pThug1rBDT0n/KHaFpa
3xiXZDvWIjRf3nbnBlJSBbT05cBStV0eIa2qJM90VXP8C/gS0VpK+fdKydCsna6OJkjnx0HOg1T/
pwbQ8Ag0jIgtNWTnUmcNl58Oktjx/XQ0R/dV99fyOWaQ6fVpwxmKZa4+GC1n5QfW3U2D8SYUJN2h
W0GG2HINGyrR7EZjHRfkJS4PmqrHpU82F1rpYvjYOID6WecZ3Nd+LaqKFc7R4V3daJA0AzDY0p/b
sKXTNXJKwOPqHiE2R+yn+yzM4zNkY7Mg0hYWAPpjhypDEST3BvsIGBTI6CibidCyWNsWhYs2rhd5
2Snybkx3WXGO0jrXfwHyGtrFKMMvgzJHjPQE5zB5Xw4YvAd59jNVjAOpGhpt/pEMbOeUibgc/NDt
/nJhk0QHgBA4sPF82m2IZL2kSUm+tDxfiwQWqV4F788cp8odoFw1sHs4iSsuWLYFHCQOlR0bi8k3
V8gaEBGqEhCwnQIXKyil/VEzEtQ28+PZD/klnd7a62XmhgJ5sRuufjiEu6rr2cmIvp8ObOngjwxI
abl2K+Yo73zE716Jop37pQ9mPMpnW1RA27bkrt/jZCb7aMcIXNGByxtMA5CGu1xqoiS0eErfMWUf
v7J4+caKA5heVu7n72SS5Ipo178XCLTMsvCJgzlmTmsmxPrwF7xv8X6RjNzNEkaz/oPzeaISWDdS
muLQ2VkGOjkSjW9OvvQK30bIE8LkXMPy/SsGSud2xcdA+dBok+F1MkS6sDMgpRn90PRwaZaEGDn7
YODop52Frl7Suo0rcHUfJwbfi7Gk0FfoKpyC3lY8Ii9Nfh9cij3fLdPBtscpgdrv33Wis7dEyylz
ThSagQQ8BC2hpCEob1QWld9SKrwFVRTMnpxC8WQrV2Wt0NwyorYMON/8ngSFQ0ZFc2+T8SXzXB8W
GqWxRLiXLO1S/fvFBQm7s3Q5L8hu8wNA/iVVzyCg365tQ9n3bjQGaAy/9acJUkEjxUq7L/DE60UE
MZJktXeZAgWYwIyJ+E34z62pW6+9MOQc9A6gNAn/Oist5O4DlMcYXd6O2ODBSDdb2aMAG7ytE3vL
PNTbF1uqJvLZnOK8DprYum4QoJ8SGREzlAu1umTMvgbDyqVZ/MSA+Xqv0U1nWLvrtsytW4hs6QnE
EKZ0B2etF9Z6BSCR5TCdakVm0kGEhdHxDjjciHAOt33E6bKzYaAsHJ8yVHMlEpwOcWFeOwdDHcYt
xMDpSrTwo7FZTFNgM8oNgI9q+WI9gUImM29bQCR2b57PFrVpOpnrviv+n1pAtn1tMiljFjIfdafl
n1uL2MIJKXPJeuzDvVJYfF/PxoJM+2y9I5ladCtlNiSvYtTWJH/jpU6dFN660sP3CsMjJB5zQo5O
qbHtqVQ7BhtYwhEFIGVlmZwXL+tYoDFRxnaqpaYfF3WTtsmBsO5QeTK4hMXAGLqd/zFSwPtwzqJ7
ciEyHzBmHp/tIhijdb/qcZatTvWF++cFroWDk6z26jgdmqJJfKalWxmwUVlAlkQvF2EuMErCJt1k
CKgrmo5P4GVtwqO4AlNwbpSHWaGzjtmQ08HPbeJgRZpnSXLEPnB1YSe/icPal8oYGaVk1i+hvGIc
Z6++obVHgL4pouyPn0Ko9DDvWUQrlN2o7ODvZdlqew4EP/jguQ2GGXlVWzFWoO1fX9/wKjF6YvCe
JMcK5lz7mqcJZH63DBaAlnivgO1jLOFeeivQk+vEwJBWkqmaiXOA6X4TVIoIg5NdCBV3UOnia7uE
jrVjSNsqKZAZFDNVLcb1B/Gv8pdmCL9xlI4/Ku0GavfNvMMf/swy6oTJ148UGgYZqVtfZsRKkEWT
DN92Xray6glHDYyDDwxLLq+lYRfuM5D50YH4dqbWsy0zwpvYBo6ProFXOfzXs6QUiCIAvhgRyK9v
93LSmnUNuglN8jhUGsW20lMiLzqjYFdE1uQXbgQfy9YMbAmKp9myaLgxt6xpbmau/yxDXScWPAH1
60n5hzvz5WpDsQ0LPYLLn/UPlhnsKdyCyqWWL1ZbaUiDKvbHx08Nx03/S82t+fVnFqBnSt2XEi0f
c+84+PWuRIwdpvykq0LsdQhDfm9NbVyg1CKxEqA9+FoDn3SN9HE3TitpbQ1IFObU5NFFYi4xwHSB
RR4a/jy46Kdqm/TdMRHFpVYLmNo/dS4ZItZd6TPAlRN/uaazDlm3V9IHoQlWI/1NIvOPuhDojfbD
PKRhZv8zCu+xbleZjU5y+gCS7DwNrKGK4uz7ZoXN4EawV/Kl0X7WHXVnghLD/onCaqtHlp+svPOg
Kkpm/YQ4dOgzZQLLsaMPkqA4Oy+62WZ4Slyeb5hpOSa0DvpX/CxMt65YFz1AE4BReCeBdw+Zz3hZ
NbHChbADB3/2IyQfQifregujBrHWKbstSktCfqGg+VSIWn0csbVo++G2CJ+VgoVsSoIWvGvZcOVl
dFV1Kjbcnb5LyYhISBm0bogi6KMK2R3ETIW2WUjmd/HGvY1wbwm7602gPzOZrSJKVTiU9zfLcYWH
Elv0Zd27RsqerArfT+81ZVi32wEy6SH9gWJZklsIfNxm/K+ntrznB07gvkz+4/e8mmmY7F9UYSSy
WmPwOnczqy5BNapyNa7PzrlRokrD1MeL0O1a0R85SgVJijgRMdPCZdUweobLVJWpi2qrIAUmHXRh
gyW5Bm3uSdehKfzm+iDBlmzVc1F9brxabIJVfcXHjJZJbbs52HpH06qUI6AnppCM80MAVE8JT1LX
ZL0pTs/ttAyUmupLHcxnKz0fsp4xp+/X6rCr2ILAyVm6YpLcaj35r3dTq1HDGKPop2AXS3Wzh2WH
q9/k7rE3iPqobstAByFTO5pP2eJlDXH48POaDk2EB72ma02TDXOYaHQgwzCpp4PcmjFA2kcDXRF5
Iq2L3Vg2ijcSY50Bel6MGpkK7SwKEklV3+W3iGQWXfs4ZMXoOTrbEDkkOGf363ka7hEyy4VGdH6A
gR2zFdzyh+6h9Qg6REUgtE+tTLk11ayrpMovfu9crL9vy+D0a7u1UxVjsFUOeGHMxsKSXKkPCSlC
NxoQSpRg09d/r7TiqxKi3HUvJPfS2nxGpWVDwdFgpUCYeA0h+cLHxuDQ5596JSkgNT0R7IB748wn
QSexFINVaaMAqvqOnPhruux9tCkeJItnFqzRyZWD44ULGzKmc5gybscphCfoRSmJ3DggDUFlMNbb
3pA69QwM5zmLrs49CpN1DU49D8jaDiBVh4uAy8o92GqVnAVxm1O60Mlp4jwueWWRLQONxWyXtZ6f
Yb8Sc5WXP0dVqmRdSLYXbNdPgqzJXK/o+d1F0J0UaZHHz4ej2ctL1mJwtwmqxE+I+eTmeL1DHOan
9QkZT3S+mxTNCPKBhmmutSUU4YSiqkTy18xqJ4GngrEsWZinYSJ5Qj0BGkv5pqTCJqx/XZeQGkvQ
ZHveJFjZJ+Z5juCjo+PmNFQQU7omdaPUsCU4rlpE9vIRqricVfptvxcQM1uUQyWD+gCtyDJKjH9b
thkw4cgNmYEqDNcR/vsUCbyo1qhvWQwmbQ5zui7k4eGdGKqCw/CKRpnzUMd0jVemn6podBH6yoXg
HKFcFt+9uJey9cqpMHDRwezA3X1aCkHaOuGd8u7GBCpVIgPXBxPtxsCNacpotU9SUedN8Y9AT4Gj
n5Myh4bE+boq15TcXD134ppdly4JBCZk7vp3vZKr4sT5JFYc3HViO/w9KdMJwYEdKC22WlHvby3U
3XpECWrqYzPRmBAgY6ex6saxJEil9HImeBFJEtq5GJIJxvOOvZkHNj0QqE/zNGwNeZFDnfNI/QHP
c1QiLLY+BC175EwN7Zm3WjH8iZssg7ME3s8TCd3Z9bRcRaIBD6CSox+g+IYvEiz4xfLJIPNcc40L
Rk0RfuKj/yyCUBANBXnZLmFQqJYWIkT47M8o1jtxFg8sgUz1SnlEYj2edATzztJtgFm5qEwEreu9
DHtpYew6FzzuQHLw0zgemMZD4tRlrD9ihNSxJYkADlZNtArPPu3jdN2NWQwPkoQ3QjRC3bOTmlhh
aCBs7Dyrl3LolWr8gTHZW8uJfxa6EaMaYElCP15dQm5eKBgL617QkTSPpcPpnTiZ2CjJdKP1Ikh7
mUfXbTKXLl1eiRQHVSaJn3RbwGnhvfFL8jn5gXoV63CKgPf3fxhs3z2CPO7DrW2Y9KIdj7x0RaaA
kEQJnSdzzFFaeWZpWCUIBeoXBC5lEbbynDgKHasqV3IjT9YBW69Ey+368TvUUGDeSoRqRut98vtR
lLof9LW91pJV92WmLS18dyazFhrkOUCyBTsdRL077pfqNx5U15Ljn03ZIxnoVOIBtD9oZzPSlf/C
GHkWYqMdo/GT+wMT15cRwrWcBFaxiwvXQHqvfLK8wDpfA6OzqOq0m9icLp5bs0rGliduzdtoIuXu
LHpyyBoSJGVWphMcvBUbIpNThDp9PSRwUIyzKYi6ysLOCnZeEoQs+eBQq6u05zsbEdc/E2kowSdP
ewcUOFM4hs38Fmeb+FiVLHrb6GbcDgafzaQA5oid5IeoY3Ujy5A6TWCzyQGzcNWwZiEwNTo6GeMV
7pmQOvWvNYpfuRZJHd7L/Kco0O8+HduiKxpnxffayYmNP3XXLtbPZAeJoA/IAHKvg0RJ2s3+PKSg
PcrBBmT3EKfOOYiE7JEMDM3ttX7AQ5jqlty100AJK7xbVc1V3fHE3rwk/KWa1Sxw7YD1gMVRYBWY
Fxjxe8mPrfebCPPNSLGcmY/JHijkZMpan/IRbHyvi7gWHHIlQp9H4KSXvmifuR+4MF/Px/pLu0dZ
TMuUyF+UMl4/Nmo9T4cdrPiijip2G1sQBIqfHdVEdLZ31gIKpXtwZNv4s8LmOMMMyCHS4PITBt1T
pV8k6ofedJWLEj7ZZelFmr4hudMiEtWQs8d1a7HdZFTnsBQPr4JWPFh9kc4D6awJR7UdieHYozjT
0xuVWt+lT3VLXRtZ/jbuSk9YkBvrMXg37E+ijsZVRBoUBQk4WucnZg6N1ETZmdZG/odVe+YAfJP+
pAtLk+8O5y8WW8Da8+JrSGPl8x9eziIyUrZyo18PdaXa0aOgZchLsF4C9EH1AcbamRgnXaPaIj5V
waGh+KPH6WlryjGaswtX5C60RGlaLH6jUnlErrE4ZfOWLksheRAkrqMfS8GKYviEk0wYI6UV8ney
a5XTCCivwNZVUvlPCYI7ehpAImJ5ZtBK0zeK1kJe6oHU1US+Ah3KVnDVmBBvcygKPpl7HfYpOQaf
1lJriwf2YXgsg0c/KU9Q2XyqYez3GHo/kKG/72A7v8gtXmAOewz2lFjGBEnTF6dB+BO1AWxUEjZc
REKfUSgn+7rH2FjfTzEonuq7XhCDuzjEe2Fsm6LvE6CEbjkoU6BbuK1h80NXC+AcMIk0zmXbDkos
i1Nr+6TGouoaOTt8/K5ZD5puI1NkPYJvH2w48wQs0dUpXBvwmvKcdmbWIV4C6SYTQGzRyuUMjoLU
rsKtLPUt2+T6aTyJHKscXfYQx2EpwP8+w1S+M/Fmq702EAsRkKvAEKceQVLWeyNT9KuEKlgP/hDp
ung9kyG5Sb02MmvbU2cuxOdY2SB2o3qtZGvGHZ/jd3bkgKAvYffPkA3s9x1b4qULGH+X3s07MDIX
7X0LV4ui3sa8sVuZ9LvtSvjySOkYHnpRHHu36yFZTVusr5zGMuwBD5k1pjZAfsN+edut6oJG0hzA
QuCFfxyzWfqOGtFYC5Ii+VInXwqp17DdPzSX2InI1qN+S9wlkbM8hABfcLOc5LI/3Gq96ju97hI7
lqDaN393DWiQQm8zI4rEGUX8F+ypjhBt/a9vqhbIBFLgwnVJDonfzYEkBodRfnlmHLjjyCHSIJwB
gsvAb71b+wjfWzwwsfUfckZjwdBLBmx5tB1F2jY+AFrckY4m4oEu2UftqGtiveYc2N2IiWyQ/8E2
/s426wLInGrZYH/O6Iep86wL+4CGKyrGmQzBVagoYHKbU+LJRtvX1mmdPJYAOtnpmcCMVZ3vBqM+
e2ZqjslHqtkGVYtiC9vRS++voCuqtA6WwtDAZYjMTOc3TBUQ2tX3N7cG5oRQUZrocLHx8/0YvOTg
3Him+Nj9ic5A+BJZg2KJBatS8GA7r3a/VBkUlMj58cqu7iD5MLFLeka0FIidUKhpqjHINYHAWuJl
O9u2aghInjAzQH/9n2SzExlC25XPAKU5EqljvOQmkrypMYS8F/p+uVH96NpEOgAIta+/1DMnJcuA
i+eNGP0djg+kAHDwjBz4jRiU2YNGNQtp5Gwp9R0XUpIbWrxhvcbeuhDRQySkQpoUmuzykmAlhpC/
fGIrM3K1l5Rw00wlsQWvYiGuPKxruhof7NJ0zKNBnltSxerp8jbv+2KHGUh/Nu36Ne0AShfpfCvI
bbAoDC0FFaJKXRhXZcRjs0K0+2WecRfINXg9wJCVK48KG63I27Gac2DxM5pKXPLEw2AOatmT87Mu
lrITkjkptCmVztTUAyeAgAAqlH9imU6GCn88R/C9zNDxBwqTyaJ9J8jC5T2fsdBpqSUW8pWGh5DR
KfQjo6KIRYpozPYYPiNxG3TqXafl6vdxaAaeMoncIfQVcP/j9qaqeOmd66mC0fDWj9O3/qgC41aL
QqfoFjnPlpIeOBxbvfQ8gCVy5W3gtkDDSmy5iXXJCpchKaw50Z8TuBk0QqZ8/Tu2eIs8aX+g2YTl
mZlSd6gUtTCbbvOyc3L6jRh5PnVc0JzmCFVBkUVNgpRuFe0nxfYzgVoaV6dmrcprGMPNhQNUvGXP
dwJr+1LqGO3IJpa3jvW3LzySq98fOIoSJIed+EcBbIQQmC4nGkHYNCCL63BPyEZnT1E88+ens4nn
m3n7egpI65vINePfzN2P7KA73oFGOd6CWc+i4QvOMIMzEnv0M/dHhYdvWKNBff4O/MV9/JWR0PvP
7/UIMxypTwrkfKuX9l5UpCC6C4B/rLif4TiCZFJvN1TNXZCQRl45GYAtTlUiGt7iIRstLccwajUh
Kw3BDLcMG8BRnaCX0rjHmqz/rogDC8JRxUu8JQvtMx95Wa9swh9sqUbvYaHQu46qcZagibc+gTWa
pGAcSB63cScZ6aS14/P86LCRceZ9TzcDhnh6qQLJLgjLHEXY+oIJEML6DEwEalkOYEH7JFrO75pn
9Rw+KYUrt2fvW8oft8vA5fGhrKqHQW5nRZkEH3ufX5nglaHBKBVoU3t95o3KBSiIrTDTl8H+8pg2
11GDrA88h6T5yNZ2qcU2UpXGmg/TP9rZ2+4vXXn/15cIJxhyIhcusQhPN6qCS3bfpIOES3gpmzO0
zvRIdnw1q7b6oi6naVa1LZGH5vfzuHYQvUwIFpyK7xQYnBy9zl6PaSuKcBISSjLv2tlZOpBsCdHy
7TBVY4f6RgRbzyBxxZuSIbL0tNkvo1M/Do7xy7lvMEeaxstZV+5bhAdP8Y2GuUgS1OTi7j4CQ1AE
3MHE2mDgcqinsb1hTFcbVoKWbsNB88c6HNQpIKzINPlnN4iC96Jj2fcKAI3lHS+Ciz6uJ7kPgYGd
bKJCIp4NfmKdlcc4ikPmqd+Wf0k49dDjVnOipXMS21X0SH+BriXPaxtL9fPozRe+fgGQcuv8Z0Hj
F/TMcudygN4mA/k4Hf2TcGrLQ+htEt39BFfZzGuor498HC7rpFQIv48qRt8oHK4uwfzo3ggvIxGH
WtHWHlSTOW5+Ay6gF3foIjoeQrEHfb8LCNnZbTS8PVOXOzv2y+cGwTngmjf6DmbvjjnrSh0z5/ox
BBl3OyjxI/MZcHIeDk6kRHuonF/Pj0cj9IQTrl5WDUFoLHT6nw7hzjaR6C0yjoQj0DEZA6pzQMEP
SN9GPARk7RrB9kHBeV5eMT+D6WHIXnf3dwcIo2omxmRVW3GdVKc0WBaTqGMfhnGiGmD6Yo1RhuTA
2LrjVIjHgmgJMNV0lNUpByiYcQqc0p+hW5AhkCSeCL/oFoKAExUmLIjOn3OJODnR/g/ZiJqvKt47
yxxsBoVfvX/81vTSXbJwEnM+HcneItUnuYbGNMA1ObLpPJBVSldce94MF/csN5nbyZ+exF6FgD44
WuTU5TgFsGorPnAs7CqdSxEkCvrMktaDX4kEkj9seYHxuvyLQ48NOWctwOjUQ/LosUfz2QQKXDKU
aZ7iNvNdCiCaxVlp4roOqVX+ea0CBQUoEdJwGuXvvfel+H/KYlI1W0TxDLvKkJO0KQVHq9rX4CK3
fWfFenHwCvOlrLr/mUMtsmNpdOR86G233iZMpI33eSkJQvrt0mYsmE7pI654tiGwauSB7e1qAz17
JghNiK3ZM+TJQ4WZSaqSV/i/zhY61nR49SH3d+zggtwhOPlMIBmaaytMoGlTZl3Z5ZKeFjPFBIB+
M2bL/r2khAOmBFoXTBXY0jtE1RCb1mnTyJb3zLOw+M5PizMq/UeAYZSc4Rn4XMdG0Q9GMfeSsJ83
YcrydsGxjPHpepvDh0o9Wo7Wx5O3G4PWhdE/sKlfpjutUbK40+hyafBrnZvVDAa0+TTZGeM1sgvF
xhqXn2d2lq49qS4Fc0L9QIm6Mt6+ABIHbZRWM6yjZoDTmVzauwz0B3sl6nwL58mFzchG1J9xvT9m
ykaJBlfa7Eo41CZmtwkJJpOPdvLULDbWYGanhwnul8n9xFurUlsLhgbCIqD7Y7NSnXLiQjpJ3qJU
zkjJoiniQqHHDEhXeP+boqaN/GxBM4zYj/byKC13MzfSMHxgvdgfqXsu7oq+BMgW5lXgqdR4T8Vs
lQW1BfsGGwv26Fs0Q1GMwh3vy+/hJaoBQE28+mpbRd4aTLVfH9K4B4nLr/ODFiRh1gdAb+R6hOFR
c+gsKnfS6L0m0I2Rr50IOov5ZLLAGKKpVpxBDwE3kKpZrf97i7uQv1LGAK5MXMoH7Rx3/rTGVcXp
7A+84UPoKIMRVO9SEcw0dYNrveoVC5YBQKLRw8/r+0rvM9FRtJQCvELC/DtZ2b4l8Vln6sBjjJ5Q
M0U9BASp7oHTptsX4L0em0aEcdfkUfc8+cAnOrIBPWraThCj2pVgzYkhNvp0dvlSf3jvG/LMEJ7B
RN/ri3+3+HYRMsffETxQmFqivlCj5u0Qq5uwqG6AmxmmBWhiUKya9w2oMCqZ9g1+gnlZrYZvUu4G
h17IaPh1iu7EAzUySUUE2Qxg7rgzNRuEvOjd4xSSNXBbXN6I7hCSoOVaD7rtQcvHYi6Wut+Vlgun
+EdsJmlV2OARoAcpydOjhR2+mS7VbuRvQhIBVbn8fo1JFAQ4QjxUOHMrH34jBNfbKcafSj5GfKYe
BDexPpjQniBkF59W4Lyo1aWSH0+0ARNc6ckQ3Gk+eG/uk3l+8/RL1d55bZbx3xG94mj808DvrB2j
ACy9WYRUpEGfTfywgQbuYOnx5rNaa/4up8VgNbAIdLjzvOg02ottQsiZLl3Vm0bQwHJn9syfAAMi
rBgM0SAcygLtSMj8nrc/+NtkNs7sLWw9VNn/UzDppDhQeIFnqIcb9J4CS9ZcyFu78hRJdG4T1296
lnzs4vX8f8h6ciKEjfMH7rTXC/gGWK6x1c4fXWvFLtjeuMz4z+77v33315wAttBNpzzVwGK1XCOY
ycx7ZWdlueLWFaQU3tXooIWVcmFOa4OC5UT3Hll4TARfFh1j4X5DKQ/B0VRWRfY+8mgENhZzseHA
73Vyng04KEARkfRuTdKHzrcVMw4gPydKVInj6onabcHHUv5/u20Ja6SbklUBHGW/gBDHx7wB+VP9
eSm7/6IUVWEr8xAXOVKCmdCSYs3raVsiIsf5pZbabFZCsh/sCYFkoaBS+6v6PV3pa0/qI7RGsj67
UDgF34F5Bzhbpurcku+UU6MofN/a2XpN9dFdf3VRZfu249nvpM1Fn7Vp//zREIT5/7wjXGFfXeXJ
w3GQMS/WMSmYzA0ytg8SZy2DWO1567tI5DfXKvUnbRhQtOT6IQ0WHnRgKSWx2fbFLa5HHyKeOg4Y
+0iIpn3VKWgQxtncRK1wx/BUUbxaEJSbN8Hg1l7EmKZvroQwTgQVvW/pBxyG+t/J9SLsjlqWkeFr
7f0w58lt84gjxWKlNiSw4ZTbU47BQkj5m0rtvTlR20u70vUSKh0H82JwLjh+dupHCPU9MMtRCwBZ
S2PHkV6jKtFPmzzA+0iohrsG47DSheeYny1i0lYHYQzWXs4s1WTyjKIFqevGgoyh+V/wE+9ysan1
VEHDThag9A1XR3PWzhv2o0k14HcsVN46FDb8CIw1f1rEy7tj9ucUZ+zesLWy/UYUQF+UpchMfPOJ
yzEikm8e8BRtM6kmHDDvAnzSMPN10/q/QeR/++oCcrUnmx9dniBIHJ6bILXP6OEsNP4mtYe4K1XL
IVn3lT6PNyVae62PBkppDxl743riQwa9vf1x1slXm3crFkD2Paaw0Zahg7FOZs9JKb93NILx53Xb
Be1GmcrgJnVHWU495sVjM5aghW5XNcpogtMJOZedqJ3qLWR+QyGLLv49oJpvbdc6aNQ0DD2stK8n
2HXBFKJT55Aufc/p2L1rlxdIuthw4eY3bkx+se32GzAyQFT0P0dLi56h7vhsP0GNE26J9sLNK7an
E9vpSc7VvK/kmrxXnF+xTWr8irRKgqR5vQWd5Liy8CX9xM3KJoOXY5cn57Z0QD+S955LVBwkjAUD
wPoK6U/AthYnAeIr+Kq80G2UxW5vaFA1ZB/v9BX/LT9e9RmhZa1G8uCfhN8zOXlwztNLmmWcXUs7
Dzo6nR2moeTmzVVxB8oXXjbPemN9vRWgyozX+N52rWxMovJXXrdwYSqOv7ciJfzxARz6QYsCUkNt
mpa/fwsKFw/CxAsT4dl7trrnuKTxacPAjvqw6idewb7r9TKkHeJg2vdF0XD0s56xYpzAQyRdaySO
2jQxv6fd/Mb/mqDpa0sP4Ns2k/DUMCeHRFpszziu32IkZTafWsNVEv5S+MOlQTiOmwsENI6x2ZaH
NPRSegLMtjswT9DKIveCiQysS5kH9z1yxPqCcddhHMh/EHsW8SB2pOGP3drBvPGLY9ChXd9sRXVR
a6zPCI2p+WEpwsJ015n+44eDyYOCVrmcVLNh94qjr8kAO6e08aDq41Jk+dImbfgQiPq24dXVBww4
ETRE08Vr7WiBImob6gSlLg/7xFrEEZ0tJ9s7abBIR4iAbtW9T1VhrUHNuVqUteGOAPNIeH4vkAqw
YO7gPVsb/jntUmr0iaxeoolAq12Qqsms4d+wdyK8skzQlZl6UijPuh8RYMf+nzVfWLhE5R+Fg5yI
ecuoY6DDPLRNrg/iVkcZ1Ur5PH1DsqUTkOlQjzp18DNhBGLlF5RC4N2O+qapf5xHuXJjzTSdKQMP
dZa4UmhF2rQoFjXH2ZoIXfcDGpkfmHHK+5PxzneuprEEwNT9xT9KekmbCwDWJ7UqBpmjV1krDTyt
NNftDq8Pa/04DDyi28pKeCGAlP6o7SFZAYQ05DavinLpgxw7dRrg9FlUKvMBVl/bdMqMpnLWphlR
Sz0Y7cwo9WdqMTDbz7coWeI6auvowv0goCtXasqcKue2UbLyTQTd3IQXES8wbaZopxdgcw+xQ73Z
lpD+ktglPiZd2Lx2EwdsHLa64kZebxEXhK6z96a9lm797ALwDv9CJL/IlMogZUQ33iA+wIrn/dBd
CB1XN5McMevkZJXb2Gq0UnfbZPvWH09tX8GGRu8g+l52KovdtCY6H94fp9n1Ook8jJs2ilPuPO3h
XE+nl+SOhZGaEyhAijAeTRbN6+p5cZzEuUUKdhFDhd7m0N4Wgs16l0CtJkPGJKNo5xSkt8VjvUYa
LpA0Y49PcqR3FgNGHIM6vhBEhXIYcNATwrrA935G1MEqHqCHWtCSN5RP6c4avcUcyayDDrEPe+T+
LF050cABeeUt/GfiQt3mUG9JvQiLPwzDBUuTt6jYkH58+ZHMl6+OazGOB4bT30L0s7Nyt+QO5IZf
F/PwSPODVBIIOJSrZNbdDaYx8mTJqxrt2nhcroFBeMnNeGGZFes0m7PJTsK7v2KciepICyvThGSP
XOA0UVV3Weg33pndZcQyjupicoeq6XIYVPorrORpjwHMWSdOE2nPNvKHde3j2tBXWqSwNxgmyebN
a6Go18+Nc6VAuWdQoYCYoMqgRA+iSm4cWyjxuj/2BAT1ONqacOMKL4098UCxBTby7Hbs9d3XMIdo
tm14zwrQm1/AlqD/OPFtq2Ww5dkJERGK834WfEJyQj3nrC2a4XtBmUhehSMayb4R1L9UULczICib
W+6TFtJhWJPfCEs8kgNyZk0RRbQzoBPFYArFju3teY5e3W0QNEj4JVDF3x6omZs2oe4lg7FvOePi
XVQ5yhvSqMDQTe92pGATfE2fHinwkNX1ljJa0crtnooCFZ7U9j6B6v8EH1LQRszqLCwaLaiw244Z
4b6QvorpIYGUj+k9xgWX4SSyra9icBFND0kW8efAecBtG0sMb0tVF7FXpzC0h4iQSL58RNV77P8e
Tyw+FYppVsf4d+dEfaaCBnM3LjRd7rkRK3YWPxF2b18DSTnCTtUUP5F8ZTNdcijYgzqCtltH3Wpa
jBan/nbOGZON2M5xwGhtG3B2gb6zqR7iYR6L/n6EsyBYrFCrPdwjj60DAk4z2o0S9q7WlUeUlJWo
AI9mpPnxj7VrtpflOFKMVt/SePyZMDHkVeDcW00NAlaY3+k572LM0usFzlCf5heSMJ9TpHoGUmVn
aErmm54ZcLz0wN/hO4P+FKgqKRUKHTQCnhvKy/lyAxFpkwqOWT03kF9Bmm05qgGTe8cve8l6K9ES
x8u1oyzQl7g4qjwGo2mt95SbOR3WR9bh5Briad+tfMILsEnREoz724bpjZ7LZtIdC/7UvRANdffP
5lkcqaiwQzSzrxqRazX+g4MuzHryLZ+0c63gwZf7VY6wkbLV1twW1wDoK74M2H4/bEB60SIftygS
MEha8IRgBPlkIBiK5Ncr1x9nyqNX48YjPCGeoi32FFV/ExtT/aemhT7wz0DQTxCyB7uCpzQstezY
/LDmQsc0rL6SMKMOJ+hp1XkmFRKxuTqv7xJB7Rp7NTaGJfA3yd/9LdYxOVDo0yr5/DL1S5lJsSnH
4n5b5wxG+h7EbkLTu5VFkptDovixfmer85eFGCIDryXze9vmW3rc/7TAaUgCMIOseln7cmsOHFgC
byDtWNGi7a1ppuHrHFTLFg6vXJaN4s+QpMcqyIbB+9NQjaVuKXmRd1XQ5Du6yAK7p6CIVcHDpZgR
O2MjG+Rh/LaPjUUcXfXOmIuPv9QGAXhZ4qHcDtTo/oSa8s5qB0p9YzuR7xysm5QvrPV87zHZwkaI
PjeJXLDjB+Tbj/kSqRDOOqX3hQ/HfpNlQuFJUijAJ7zusbsmkqjXkrKfW2OXvChQpBpaJt9dR496
+CNprtJoEl0djWo8G2L9OKEASKwvgJ4i2OWH5YmSGxvqGGAjbCg6wRkm6tA+JnA7OUKAyKYBBC+m
gexprWtf7FvN/mytoMomrLWkNSs9Ic44CMYfit7/FFVG7fqvu8FjcfD4rX36JhM/PKyP56S+rhp4
u3YbTYc5Sh1KyVzkMz128bZoZMUbNWyjldWs8pNbLjLq1sJAlcuoh8chKLko74A7mpSjlh2kQ9ge
73rPtQ5oaOXRRMd3kT1PIB0Xz9/C2EvnUNjsCsa2d/ZEYP10Dpu1DshStXm8eyvhDKmNLoFJNG3J
ZHstvi40ynnYEQYhvJQCsUwPssKBmaEB1vOJRXUznjMsSx4wRFfhJlgxj2sSiQgETRExy5g0YJT1
xAuCi5ezXRCcPGUEfYsLi83Obw+Ha8sdJuwFKzqiVY6u/bi+dfUovVFMn4GA1NXYsTf/LQlKuW55
95Yeb5cmZ97U/56XvMQxUlWgDVXIXg06zMKKYzusrxMjYyWrEjX7/Mtp1bAGGWtzas6rv9pgWPP9
mOX04lF10jojl9ez4a40cl63pHj8lfz/TEoytnpEGqW6MLDA02h6EDoeKrBUMXocZyJ0Z4qI6OyY
XzTrx3RbEemREHmZw89poq/CwxXhLKXFVHC1aAEQt+RUizy2pijxoM30VytHzxjHTySnY7W1Tho9
cejUYY3Qxky2SKZ9gHi2GuDmAqcSCv2E+tHycYlcXOCXQjiFvJY5Ka4/k1Nu3HDpq7alg3+QBBcX
PcGDjGyKKyRJS5j4A4GOhpriBeiNyPTLKN1Im3PNz+XI5wiHARGbZD/JitvD1ho8XpgzREyLQ1zK
dDZp4sWwF29iSAjgwVQ/C26GBf7lZJkYkJ3EnrLU1O7Kq1OFp/jf/ggTk8tuFzKBh4PJKvJAh+fQ
w/5uAA++ugk/wAEQxzBBlUQl2gKfZmTt8atmFCKpGxjilB/vx7/jBpMw72olsT/EMPnz6sJSDrff
s6H03Cf7/hFLyksC+iQNZNMQS5QKx+LB7TX4tcxwB6dUec7q7SqNF5qvIiTyUSzHL4+kaOK8FDvR
GpENOZvkIZiHVWeBkyVQcjKN9NQ3YEQpIHeyK3JY+HWGa9d4gsBtUR8EP9FTPyPIWc0NyMSrZWJ5
MdLEaVR7i2uJHwSIpLqqTyMusakiRuu0zeaObousMR0asKA30aVrnhAypoDj9nnypmEqPhTLlUzW
ZrOxK81lOHmYamHzM6STD4LrmmCcYe16myWUsvj9GCYp+DE2JOfsAuO8wMWjCyB4qNUFUJpC0t47
lbhRrtn+kp1k87TZPPOUk8U3fq8Kspu2Q41MZ2ZKeKT52UgmIqP6zjdMnthjX6AhzYYe79/sBqEZ
QGdt4TGZk3UHfu2qUSPEm00fYG/bnNpwdGTmnp4ryHkt0zFuAazLdr8AQ3gW2lsAGGN0AB2NSDWx
8QP1S7HiCZR8UEu6oLjES/T1SkDZ7lHLGRC5aNdMwQDYCqgQ8juHFWwFyr3c2D/BSrl9EuVQ7e6O
fjhAIhLOBVg/3K3Zor4FsyNqn8JLVXscr0YTXoUdDRbTPNtKy63xaQJqeYZRxLmOUVpzy7hGdKCP
LYH7ncIT2r2Z5/2lo3VTy2LGYf18ZBiz7q2zA8Mo+fy5VtT6rrA9wb1XZZh0lnWjUQUk9OIiN5jn
4jh6abQLklhTiF/9LFFSiLP1IEhY/wMoLqD0PQryjhx15W8QTORVBCXeAudZZt/ms+3IyNarkIyL
Q0cV4FTXGRLOzqpnAJKKmOAE2t8V5KAECDy+58UeRjuHzuP5vl3V8+aB4oF8jhbGGT2hZVbo7X/C
ZJKDXvQylFlDw5/w9QXHPBAekP1VOYVXGnhklwutLdNsxzhAP+kmgpT4D9QJs0aQ3//EayVqHbOY
Vz+ObrXJi2wAFHzuwcBwjfNfeRWorCKB77fsUb+Ptw+1DJu6GWzF/BQ0OvaRHXLatfsTHw9vbFKR
nLAh/KFZa1MmMw37SATZffMdjGtqNFGrW1yOWPckmy8lqcRoFVlY8Xk6sv02X5z4UE1A95msGEv9
BKEO72Pq86JXQQ4lE4oPekifY7lKOblcSW6Pt6u/sPcPxJhrn78pU/ZVcBclcjPd1DBOI96fwN/J
BA80/sUpEVHZK9gH/rJzk5vS4b7fjaDMZk4JaUit+Hr7NUUXl9SJew8LVnZC5rCE7EQ2KBzbMR+4
/3Puo7NX8PgMvju5SkVUT17roknp/2A2aA7weEEzuwylYhcE6GRAzyTLRajsiGZr8MGxO1Ux4rC0
HsxLn39GU8/ndL198f4JjKt52J7a2HvYM6EW2U12Vk+rtrEG50EpzuNkCAoonPn2ZUvuQRGPc6fm
zxwhrrV0pHgF1EtxamPRyw3Kk30n3HIOpurW7cd6ZJ28vDX0lh0YBvFDIOx12FC85Pj3kw++7VD5
NMjbHDXPCDFZYeNUfr5Wd0yFgqWgWFVxQ9svl56P8TBvo5JoMten5wsLZ6mp+EbSIUPtajjKP/S6
WcbEQh70rXwuef3bnqzCAEfPZWUJhBVQPMnAKXuq9eDv8FsO3bJTiKyiK6n7+mXW2sMyxOEnfcdO
MOorXg06vbAs9JC5izQDpJD0jn0HDelczZjiZKq8VgAOPyUm3ZsxaDb4r1jsR3u90PeSTwbNvLSF
TjntGl5t7m0ig7juv82pwR/Y0XNwBvCmfSSD+gYqGk7WZJP9MRyYflv20/MuN+GvkkGpQubEOzYD
2I3qVY7JlOUca/ty1tNAGqWjfSpo5kfJkWFSpQySfY7pOb6erE1HKcoFBQtC1B/8HVm4OHPF72VB
BCnZyf6qTOZxyuvyfn9rFzcFaijz5sWs/wdq6RtlXqhTFZFCtdw/tvJCYnr52JFW9Kcu1/OKs2nA
IKSc6SxHIIq7GzUgpldTdcJxtwp+fp5hz0Rui/3IGN9WkDWWcDUtIq6dlTz3cAp6oDhXrHLoRhxF
mKVl+MTohMUZineBHR63yJ3lMVDomPGSqveQCmGsw4ONVAmYxNM7byZbwVkhYqOdIxa5XV5kgc31
cbYMdTw3p7XmC07F/TTZ+gzUfHhYRmqVzXVBZ44b59qV+9mcPdAg2rcWoxVlRGRZpHw8oiiGcUfX
MxUy8/SRltHbuZ/7lG3OIO/XTm7Q/KCMBWQeOFsAD62HTEh5lrpfGakBVERfNpz8KXf8Gb4FrUAk
74Fqd98a/jSm/AWPWY7swo5Aq+1B0fIbz179IUFxMyBh2ASsqNANAxR6dPvAWJXG+BQsKF/Ob2z7
b0QyCDhXgyRxB5ydzoNtbvaa/7sBMySpeQ+wOsQUAAMzkRE+gvhLlhJPd8spEOpbzpaKIwRAm52f
yId+i1gXpaW0DSGxvHmkekVimkQzWBpWeDdXHQ0kmow0RYlkdMoi1JnlYhdGCX2VNOoJgKbQFUOK
VORw4o+v1zDX6C+te/bkJnd0f/9dZWB7OYv2rfCVdrSg9Q8eXEdseQP0d1LDKW8ejisMa/AWum8I
SV+iHfj+rSQMhrGdsQIdy3+6J0IiDvmY3j/yZ/xj/NfOO6E3y/fDl8samRanaEKRBAa7MZwEstV1
CAoPpcvtnEClnd69noW6wt1nbrtvstjwZVQKOJIin5N+OEt58ncGszb7oyVTR5RylCys7F5y7rop
R15a7WFpZyCKQus3sLrCY5QTUP5VvlF2Igu+JFG4q2HcsgWEFFu/SkPSVCU7YpyNQcYK60tEs5w4
J8EMpB1VR4wdnhzv6Gq5pnDPGYWeTZTCsAT54sKrB9gdXH3MJVHbAziUwzHyWCKHSca0RBBTYzlJ
2UxjBI37eSlwLddxaKzSef7BKV0Fpn8dYu/ElSqQNvy0bdyMcgzTzslyvkAv8/TVLej5T9ttGMTd
3ZJ3GOmO3MgCg9l4mnDGPRFqSUB9SMnkvNCy9cUCF0Rt0jgv0uMIhc5Pgviga47jCElt5NcMMBRI
KxPprz8iXCNPJREL0IelEegmLg7uwQFRGhW/HYhe4CiqEy4xCD0sxvtiUNnRAH3anQtw3ub4XTjS
ucHHAiM5InfBO9/HTbunci8/3QC2EGuZ9OfUIu2sCE7t/8Wa3hrMJpaZ1JpO0wEs8I587TNO0qNW
GEiJrpM/XWaynYD9l3wx4CEP9ihZCnsfz/fObiTIPqaZ7SUZmdk0KkRtK+W27h8T0tAE3DCt8qRQ
S/UX55IcwqG5PzrLAIwi01h0F5zp1fMcUVzhjz+LlW1YTDR8TRVaqiyDdfoVNGW7jn1QpzNMWTYZ
flzKqniiQspl9jzi3+dQoiRS8sfXFcqFPnGz4gLt0KxsQjqyZMN//7ACuqBHwkC9rtqsqipjyPpR
dFOS1KbvM7LP75RI3u4+e5l2uH4TUggp/cdl4R5TKVXPcoaUYjviASjggngsk+Km5RCEhTRNVvR4
jDAwFhdRermh3//FIFLDPWBC2jL/rgjqfyGFJqMQcL4lL55PH3RwYYcdHhsttHYgepP618O//7QZ
2ikZSvm7K5Re1DxvwR/emEAWwYjLNKby5IB0CpF8QVApIAdroX9oIt5JD6haWJC37s2/xQmuiMHf
CR5a5Xcaqou46sdvKIlv4aj6UtQv7h+3u6Z3yB4N24pyq7Qz6pnzfWptZ9GqaE2dAGjc8/cqSNxn
zIXMmhUs7NTXqdKN/qH9Dm+tAetN3EQEjK3xWdp3OQ5P+beBQdBU7BKEgQKvGmr/AH8IoWYdViNw
/jRRugqH5B56gkwolNyALaC6w+82DPSRc1NkM96eENKVLjRZriHNidoJflhXRvsPWKMehqVYIIVb
wmTD3WTndROL63xnZmUjcn9eodZac9IU6Wqf9HE2kFDOoXr7/EOGukwHNb+CE5fBqEVQGzpH50zB
eZJlL+m8EeGkE5w9Ka9MMoB0pYe7WipwIIOfeRIEYi+UX1jCKpX9U+vEcxVK7Fdow4k6UU4PJRY2
dPQG3w6/nFAM63xnOPsFv0KxbSTalFdRacCq46gfNrH+AJwIAfgnoUtYFbPxecg1+XBVpFKUK7pE
T8QRXKHuHvHFahLL+Bo7Dzz3So5k5vpr3knLHZma7LaVDwihpA6Q8zHm5IGCB5V54xWMHVU9NmR/
F53ZbR+qrypTBBBYKf3N2p5VOrbgP20bXG6z5nAB4kWZfngPTI3toK9Br5jMwRgOl/l7lLbZQZmF
bh+y5YlgSN7nyq5aFa2qn8VlMN9JHobAvMcyzUG9AAvyrO0BR7ttk8qnl0bS7sxPo0a4vBxcUMOi
chF31dwit8BWMFX+bDvssWnU5/oCKB4KX9hnTKcu8h4IonhVtMSc8J2V7/g/NOUVPJmiaHACAwxV
rEwLxhHexNiTfAKM7kPo1Da0ecxDKRzgf5GB24LO85liRFtXbpB2LPaz91SRpfg/wUELW0qQyNF6
ajomXaEMexXj9lMlCnMQm9PNxI+zS334MlQYt5aIobpT6uR8EiDmMEu2QWhH5fd4h9X42QY8X/Ul
E0Djt7IZLsEs8PtQvUnVqvLBhrnQh2Gnhr3lP8NknysBvm3FwSAKgOD0ULaKzpHDzKl21FsxSEHN
OQjo3wnF+3xuptJoiOUBDSEos/C+BzMrPqn7sqNAoTPdnw+4p/FqzOiyqnHWLjFE5vABt22ERG7t
uRfkdIOgX8wNhUhXMHfqwoK0wVWqybomCWXChh6TNNFNEGDgFKuIz3Ae4vMAEeqYMWjqJjmR7M3U
6vS8vVwgshl6hfGrJ2u+HJj3SRdptaPOYWc+4uJfPzq9NdqvQk/nWFLzmNesdfbVJCYiTSGnBEI3
MzcuAYtlj17gbgMOuwITAKcPZrGre1yrckOzTqROCJZF0f3LpgwsRAJqox0Grqby4qd2RzYyX9Pf
2kLWipxaDBrFDJZSC/+g/J5DkHhOJKSOiBzTeI0ulEO358oNKoFCXo7Y5M6kKoBsaeV+NLlf8ObE
5DQXLppanWcHYAKnJKLfjZ9I/xDEwU0uRgqHYlTMHrXBkYLdpv0/mxsx/Kn8QFF64sYBeoC3vM0v
3Qyu9COpk9RjmTcDfIuwb/ao+d2QMziBb/fvu2QHm+mCWKiMhxg0GlWNk/qY0K/31wmf/tVSMuDy
OJ5f4kAiIGqeeRS+XpJBIpwVJSFlql8QDCDLRkTDvkmKzA6PMeBgDb8DUvKCzVa7gIbTmOpI4xzg
7Ik7HEO9IFdFBHjMLr0OfTJcp970NiwML/djYaQzHO2zAzQRaDt+Uk+3VI5SWjctaFqmJLgn9UHd
+GqCnVPqAvhPK7cafLZLtcjvE8CiTD/P8LDpoyPJHfNGcoY4RU2xMPd1UnNYzJ6ST9F0/KHWkFOu
iJvCeR3leC8+IUBx8hsgdmuZKEF6Q8Jb27lNw0l3fs0fON8X1VGHLfcBt7maluOz+8xi69myWmzp
PTbUq2Zh6Eal5SIxEgGGfhkOo6nEYhSkHqYOWzHseOeB4aq9r6BFXa2C0jnuW47xqGoKIrT6ojPn
NDcFcdgtpArMHWMijCzi3gQRjulyUiVZHY+f2lGaWyGt7pk61VJS4N3xAbF5tNE9q3M3P7j0Q4T8
kPJLinjEf6oIDew2fsgEIxeYLK5nbn+yf3YWCOeSdhrfNKJq1xvd5EJtkCgVweWgOtD+NQpv9EkN
R9sIixkQ0z2GfyKUkpIqkNmCPqzVqRoU3xwAv3EEgWuW+cyCjXR/4rW5VtPnBG17EpYgaAFWXCta
h5D2zBGjwbLuRMqVDmdeigXq971dYqgxIGLWb9QZF1GSADbdWjcK6qjnbaRNbjTtlDMJpfrhE7yn
nOZDajCd/iprVJpBqIa++A2S7K30NqHjlvMuLvQiGJRDI7Jm+YIIHexxaxePajAnaMWO5UMyHFxA
txrDuXTj90HsYpI55Jn42ABd6EZLQ86CgIF/sPFP8+LUiCAW9hjQxTRosuUzOGnqygPtH/Vx1x/J
vWZc6oJ5HSLa88g3MsXc+c0/2SRKYCqBhMgZLgyQjcoZxgk+2i5IvERrAxjjE8zZ+gJDuVrIQQOS
aClQUnBEc7RegEBefXFnrPkNIl9anmgOR93zsr8EFccATKYmRsiInGVbNOWT8BjzvVVCYDAUknTd
UIXjXfUUY49ZedfhQLSqshrt16sFMjqv85r0oeBcct6FTrvoIwNd2b9RlIjV1qUXmUo11ZA2BKY2
z/FiBgpdGh4EyWUCBFWtxJdcja7nnamCKEwVm8mM0bFtNg4QHiMwUx9vc+vBis1ENKIU0P8lASO/
NwC1XbggbmsN+t9fJbUFmow8MuHQaa8QlRH5lczpv7k0KEKXkMIfJnnS0g1IMQjlQuguu6PWrgsm
0ZJD+KpYeIzQsHvr823J4w8ukzSSEMuMx3NtdZNnvYCZ6bxtFbHssOHrnq/ctrpAjDXYXc6TykPE
AFa6u5GMSIFhuweFI2DvFsouRSYi++cd4SEOpPNcXinPjVsXHyQOLvKNkhNfZXaJzX4MGQJBPsqj
ZKh7sRPcLS7Lcg8Jsd/U26nJt4Gl84BIFqTpXJZqKOZI+DQbEW8JpRaxC2RleWIoZdahOQhhnYtX
pYKw+66RugRDj3U4z0Wwg21h/VNXhf5twGVPXAIbApihyAblzbD1A/+reQD026puwhaeKHzR3/dS
aRJRIAFFJvQlnv2CNvXtosvcq1j3QUAVEv7jHcFH6mnku3LHlZFLXhNQi386HCYUOof52deieuiX
h+Faqn1Q75LmcA+aPwN7iFt0at9Dli9oiayMaUBxVtG0RAhBSpoRiM5m6Zbu9TnfxIx7ocWyqObj
Jn6HLtTSAiLaQDL/wczR9IeTzwIKzrpS01+7fbKEVyNQV1xHMcCPUZoiK5kC15fnN7gk9wbm8oM3
/xTl6RrpSOiPHedR4cTm/tUkoIrq9AATeNPxvs1SIHKCDljZF89iZWZVH7QkjPqZwrQRYgJ+frjx
WbFltnCgN9yvRim6E8BV1+it+M3lBzUtEsF1hMrfphDdfunevj8OtigCPXZDJ6Lx2JiGEUWPFUGf
5bamrwzcaOocTlqcvPQ0CGJCJAn9SGOFt7U+atXeCSmqkdxGYcxel/WTISWUScdi8UJwsShepP7F
nzj0HChncP9ciIUsu8gjzm2g9ZDUlCW8RqzlsyBMTbEzLqRFzi4BeCpUIDVCxOohzBThnC2VDsbc
mRlxfgDdFmo0wDjzuA/gsnQ/tkbjeA4wo1/QZ5WnhubT06x6p6hWhH/FUAe2ps2hTI9uJCjlFF9h
cHqfzUnhL3YTqD3vnXYfnnxr3BMx2W1SZDjijgpLU1mdKIKALaOhuV5vceHStD/5tLzlyFytqdg+
d4N6ELiKxFluBiZK+H67TtAQLEHsK0BaJjnOL1b5gKHAuBR8eXC/TZWd9T7sRxS1lAxQsi3ch9yH
66Y1R+2cEvVGS7KQQ8OJGrK0DxeDl1gAiHz91SoEv4oMIpT6vc+YfNXbobK36OLqovBmyIKPXqYo
/NL1U9vWEJ6cYn+T48n4Mbhu26A+LUq5eF7zBOlpJ+Gu8gagot7XwSYLXrAhaGyJXcyFSV0wRN2B
6IapojMOM7S3romjNSXL58H1WCKnlJDxUqxnkfkr8bl411KvX4PCeIa1uQimlW7Sq00GZeGQ6Thm
SMDt9KcTm7JMM2uRjC8IzaqncwWyrIp36WlRAYvC97n7iwLMZ4atl7VI2zVVEJT0RJMGfmmk1PH/
o2IOJiKygNwuhtYD/HDhQKnnsUbjUqx7OwkQ+Dy0a2H8rEF4irdFI2bqDtKuYgSgEqgS91BfwKQO
rC8NvzxWKqAZZbjCEDiqxrhnZPy2rjs4KIKOMpOTWQxraT8yOD+PqbpTjSYgMPwC+F8RrSElhcmG
XirPgbA2r/yKUx591+gOMtmHxcGKdxJD2Qq2LSKl72OJbCskwdYdB7OWYoTAzDkBxmo1/SEaKz08
KSzA7Bfy+5J8k2rtI1yi0SgQqyCYmN/rQciUqCFVbIlkQl/gXbkovnXFP7RsTjWjzcOqYdh+P3Ls
AJzDiajcCS/BjDpHqnc1G8euXd7JAC2P6N9Q85ZbCyQNm0zai2/2jPP88igkVT0yYOi2tdRqWLHG
nYvGqPTubgvzkhRlfTB1f1V0dof5DNQJZHVo0qoXLxSscRrzgH6WJN/HT4dMSi6S7/Iv2XWNpdw7
Mrv37f8e73U0HbGG83+nnOGWahXNedbEYXfOahl+9Z6AGRF4FKla8zq/FD67xJ8hlJzUV0pLe6gR
jGf3ksOFQwx80q2LGAFQB/Qk+28JEfWDbWrLO5AQc3tm1OzKqRSbw7sPjAGjwPfMeMnGmc5z4RHa
BVVEqy8FPJSXzctqCSe/4g+aGFJJoKOn6H5/B1YOgji5zDwT89dGotigIeDjatFTVvM/MOEFEJqH
AnAReJmgzNWqOCIR5DelSLv8zF3VZ7JV7LJWm3EJNVdoTAKZCTJBWe48dTKh7mM5mPjJ/VXdVMSp
+8uJQpvwTZ8VXGZZEwnVFfj2ky2Su3OaQ0gNMdYPeHlUvX+Qf1s0WgSyaPEAymob/9UYwypd7OsN
t79WCXmEbIgRr3EohgxymtbH5gKHadHueEr8CNHNH5xtlL20AhGQdTLMWa7CFESwEq8NO+dobdBo
12xWkEp4romnbss1DRVZ4d1JedmBhUT0zRZ6piTmzAqteHH4JBOT0co554Pz3Xp2t9l8k46AWjXi
yqMMlaVF9mxAfLXlinx/J97bAp2aNzCehM07gvA+9r/C9sqHaYLq2weFqi+Fd8wsLI6zP0W+Ydcw
Q8j2v/sm449XfscKgg29adGBAmEgoccg48crLrP/wVD06ciqWVRK96HTOil30su0Kh4Tez0OGh/s
g4Fa7jD1/ZK9/ZJsYJB5cGJc2+Vy86orWN+znjIJjCFTxynkD1PPeFpBJ5hz6kjExwuRpUylq1hx
t9aeex/XcwKkfXfMAKitVN6fu8pxNjVDtogJjNFA3sPwJURk2ubQARoV7jHY70OgReBwH8PC4Y+0
YA+H7I3O6lFfAYAqFHKXf2AO4yQ7BPXYS+UEDDg0Btx3JqgkR1DrJdZfTy00Mfr7DuvzA7KmlW34
3HQM8t0IQQvXsonKhjP5XXabkLguOrlGL54nu36+O0uhT3b7brfAj5LLkxIa0YAUKHHmQscxWkad
PggMD0Z6mVOztAUeGL9cK2t+A7HG4nBLAlPvH2vgEzg+GOJbz8wM+8BWTK/CVt2qzPSVb+2iBVNI
aGiMnqy23i3hTrrItqfdaVNvsBhx/Jovr6hIcxiFjmn7bxPxFBCRlI4phIphbKXBrdFs03+pxO8l
9Az37K72Twt98qI/IZuqyFw4sK2Oq0G7OkYIyNXznaDodxiId+t5iFNcRN+uJpl1FF1+O065w4HR
sETgPecifsZkGIalOQqQ7G1mWXi7g6a47+N4+FC5Mtrq0IQWHOMazycjbpWDkdfCzSdGpj/dd6Tc
ivagbfGfRqlwjIfGOovn0hnpoFEnutQv4rjWs4O+IDprHKtl1a/waTEEXHBtTYo3VORepbDmdXuy
VjOiykW36TtImmBOEiAg1MOJP8+P9l2cEvP8GjC1PtJF0Qamq9/EdnzWf9f9L9EqRMUD8HF9HLwJ
nnX71ta/hhPASUa6MnEQaQouggvcDJi5V7G9pLg3f+AcDFqCHe0HETX1Sgrpx2HM+Ugu0T9uWeWv
datDugGaEGIOx0pJkCDt4cqkpVOhxeDyfvZqg1WtT17081sS7BQT4q6fGdpPZ6uCzmXBHsKa2l5v
JmkK6nyaE1pCtKDo84VixpkliIX6TmJYU62DyemrFQWRJbcjxNMFIBFdScWQNUp7+XbkbQly9jTv
5gyXuDp/vnf6UULL4pzKWpnC+U6XpXeNYcqDbb0t6sj8AVXHl/r0LiAY/gCxoCCEAlWgMGIpiI+2
T0rnOkxJyO98+GSu/kiwkEyRmyiARXm554xZZo0gZBGNrfKVfnclAbcie5+q1A5JBeIOecvbzSle
vCgjdihRAmflNS64qn/yWouGl21v5QHWwCpEvujduvPLZkwe7OjJbyXIoExqSMy/q98TJfZx4qpS
WR5094JV4qN0m68yQfdHqGNu9N1REUCfT8JPdQPWSCbPKgrwf8UcAQPu0w+fMRQrtHFsXsGIjO33
l3mkMJa7E+CENhU4DYYHq0WWI8M1NWdZILBQm3r21z0j+a9Y1yF5/jYROH715wXUX12DSrq+ObHP
3E9H+EzwaZRiv+cp5iMvxo1hRqsQmqisY+lIHaPvXak61QOQxTUqZ9J3GsWSBSPEthipDZbMxcAv
4274Oqgk4PU/dMhYgwmoNUh+IW07E8YahKBm1UotepHhdH6vn90EayP4P4B1YbLinHo0S9a8f5h9
l73NU3XDSoBSv+CqqVRdW2SkIhAu4BhCyh6wTG1UAYYbyvPYLowau+7oaWqU5Ih3HIdXh2t46bti
GyOB1yRC5JD2C7PkFPxHkyEKbpCawAgvvcwO+zRyfwkudjKQFHbegcvUT/1JE6kzWUgW6Dur1LTv
McUbHS8pUnS0XvDNa+FR7VgMxPy6b97RBB41dJqSIpc84RhOedBfbODU6PvbsV4lz0+G87aHkh/u
CdvUjvlDHOrDi/EHXC6MyhqA3achlJd/nRWfWHVcxFDCHymZhdcFrJ0bAYGevFyIzaPgMI3CSeLC
xZhrSjkc7pt0funDSMx0nZd0Ry8EsCSqdnHHWD99UOc0obirkoqQuoh5/2IG+/FaHIQuIlAhPH3S
JE98hxRas15oCrl8Rl5ub5kL9NYFU4ZkPe7xY5gcjW8eH3oZ+v7hngcIApUasLNUe3fBMJnxYhfC
aB1CkjlhNFs7YqNBZ7p92d2TUJwjD01yKxzKG3dctMWSkkXbX1HNT9nhswPcGjUeFmc9v9c9+LmD
9qAdni0FqPbLsxaod12Ad6yOy6pa6j4Dm/tQJii1yDGt1K5WPIvG22aZhRaj7/+i3lGPtTzb+2fO
ljO1Q+d2YJjdcuYTSFxtvrTySpcb/pTYHvpW2jtvFzxEI3SVRuZDO64cocXlZGKkbFz4WbO4iCuP
u1CgbnbnSBKexlazfdZFIp46n1C0xU1hcfosGEzaY7MZEROMQVyyk/TdFD32+uT5d5oUHA0m8KEK
EcxUw6GFOTJcc2GEew/Knnu3VehIHy/HAAncd7pYhA6Xt+5uLpiORMMS6UMFC21vH61RbYBCMT40
M8a59mRKunyOUtA1AMUHjGwO+XS15wXtbWPguvWpOPNTcDAwTgLR0NlexIv56dz7gBWc7b9jqI8v
aj4M+Sdp9Wjak/4wDII0ux4Seueum+iHspB2/ij9XzDff82hfmTHfPG1/jo3gSi4atfnaYv4SXYJ
3BisJF4D0UnQFq5JX05fLiZ00x/DMVaGZEYZmvGasQ7c70niPKH2oceQuuPVhEXOmClkRO+z9qqV
2CF0Jbrx4brKng5+AJ1uZs1gSQzWqXeR2PamtTZwsFz1+zlg8ctbs+l63l6NF/vRTWnda4wqTVen
5jGTccxXTw9qKvkzP1HnAMnCijIlfjvni7jAYokGx2Ud2YXyeHxyQ0nqXfurEIvU1BbT9ZFYut4G
RJfTxuTdi+/cuh57tHOCnsTwbP7v2tsD7KO3usfSqCt6ruYEdW9F+CYkZFTykKJGg2dpnWGGMHnb
DCToYBi3lPLCHqIuPBDLU+BjE0yhRQm/aVWOsvUZeriSsEFp0TkBMxp0GF7zkQKL+UQ25Y/J04B5
qty0/xdOl13VAgcEgRgurNHNUVV/mvOB4rLJAIgfJRn1aS/aee+9bAlf9tYOBiZTB0CPa1lmgTIL
oTLx+9b2MIqKtHvOa0lkhhc5TyhwWhGBGGjHlDBOD1lJijpctLZ3Hcu3RMDoS9UzGHBlMki0M5Ek
PUa4Xlfuc9wJ+covE2P/3lrqFJgCIFbrDQkAuNduLSLslLK+MlWERiMWBPAwrplAe3Tiu2367Upk
w7BdDVe7juOibc+vHjuP+p+o7w4+1EkUiOjPUI0KQ8L42appN0wxjFP2LK2H7LBvltxEDTBdd/+n
nBXAQOLl27MGKsQ6BFQhENuakgKAqUW+aO6bZHZP6CJOY3qt0z7Yv5kT/SJNszEdRfT7Q0IFjSoG
WRUTemYMRGu6V2j6KCOyD9Fz6KUG6H/KWhCU8BCPKwRyVtFHdH9RW0hxNRjeHsvbiQ/1VpR2bDF4
GI2Tq5+dGPgnL6D2+sG2neWNQuZCiyJhVm39ouzcgUgsmOfmydf1k+HW/60wVkns9qqHGR3TOgE7
JamRNlME8yPjxjiGksQkKZtY82iXRgiin78WksN1P/dR6/2jTtAlfauNx93H097aLaUeI0TT28TT
EtPeNdRc/HFw+qJPL+6cJqMuM4KrCTfNek/s+KcWiQx1QJ4L81qub+Hja6kqo/cOqBtBZO1xj2AD
yoLCt7/0BVaxJYvGa4tXO6u7OI4zh9m0oLgXl5XtEmYmQHNi2P/Zi3Gw8rrWsXUOOQLL1avxrLcZ
30xIQC0GA47tdgXkk0YAUzNJZsu8bTD0nBmJ3F5zWRm6QQfoLcOjBD5uQThwqBa6oNLCE7hZmOj2
X54BGgBUvNfJjYd4dLgeNTu1kVzfZ8DhL4cwRNfuK0uaY2MDIZwz9uhs+oZPbWFq1q/A1Wy9IfaP
ivOogfqSvTsi4LlwOGsAveNvGyCfDUWir/0hlNPslAM7MEWezMIZ66FvKCaanSoIgTnYZR6BY78K
pjOXHLXY4q0gDWe0ehZNv6b20FAazUzwDB3wZiGqYlTruM7FPUGfwvOrNv4q9lPwcBc3/FPTPJQq
/BDxWkOzGkFKEJcZHEKDTObIFXLzdC2c2InPb13wGKeStmewV52aeTqD5Xt7QxbuPoMlpdg9QaVt
paAqAmMcJZ9IUJJeyyLBZOWeQyIDPXwb+bsajLn2+v9L/9vx/rPxoIRWZ+En00QfPR4lBeqq4s7v
aV1EFeB1mfYIo6cEa/V1Fzy6hvJ0B8FCvaADL36PkBsWIXHDRQcSm0+D1fkCIIt8UvgHClF+lON8
elPXKrPW9QF10MLfOJ/UUIsgpDYhUpVTnkeF3SBi1c3pjQFiSXDd9Yec2RXdNkQkWKmGN/M5acvF
NQeRHfbtwOOcTbzKCKQ+akMEPTqA9VJYYfW++ixZzfW91KJuPFMYDUqudsV0zfg/OaplsqAvC3+P
a2AY+XNZO66ZrC0apvN2Z+i/UwHN7v9bWA6A5qDRsVVqOF6TCQE4OnKeCPq5BnIQ81xwTzEKRcmr
SEC6k1DsuEdS3pwpXB7ArgKP1jwwsii16AvpTD9PHsxMwnCVZhyqu0T5A99f2e1d/Uz67aPL380p
hA4y27nbbhVdBefzRWrOW2KhahVslPtlGuwToQtDpWEGr2nqLP6xldNtSmJd+SoFmQib7+aJKHyH
ez7llMwqv0chbAwUzGl4RUT2EbWFp9U/2XiOuZDs73CxM1U3ODtj5iEUoovv0i2G8zT6iCk1JZX+
gtrC5wiZdOAnp0Ymw8sf5Zck1Fy+AjWTWBMtKf7OmQOwoFlkY1RTRE1xax9rZXsP7cApgdVxcjBT
BgD5i2OD+YPw+Op8S/Dv6Kgfl9pu71xQcV4tbiRCWiyfX/TLDMaCeZmeT9yWQ7b2fpvN1KQAtIL/
SPl3H3a0yi3e4VrbMgZq4O8HPkq/aOcSA2KrSwXPnLJQosi6WYl8hsKxz6QGiEtOHzY8chhFSs8g
IGouqIBgq0R8OZkGw5V2rkNDQX5Kb9VWiNUOcz/SbdQ/J0wBadzi4QBwNhgrtxaOhJSpbHKofr3g
cqwBEjVGEtwKVsPbXqbyRUYokJg3FgnF950o9xED5dn+NYj0aVJ31g12CqICRMfYzwhMjtBAlujV
iLSaNxxlyenqXnsOrj0gLLMelMfuSrSy5IJzKyTpvZ9v/2tZ/4xkov1IrE4WqdrGG18GMScesxO7
CshHgrskGtDZmwM1v/YraUHQPWhdQlVl24nOKxzfP5jndClUZwPLUu9VepdB+mt6EHbABpPEzjvx
+v8Nvj8jHX81ehUIl9OzFcK021tvRuimMNpIt84Lo4h81ggCcirdHR/CVgGvPEvK4j1dmGhWKiXO
OF4XCY44u7bGHuFmfX/vBxo7FoI8bSHmDt6+h0EfQY/70MI5yV2CKvDkXDylsMx/EGva7BGBBmMO
kN60m0FpPAT8K1VUWHsU0ESHJw24sSA45uN/7PoaZ6/ugNFuyiESE4lBnh6rTEsicGEevquTBbbe
1gLsXaE+2lzrNOHIAnPDJ+PFPi8Ox8iPWDetsFbWqMe1/xRSkM7ZC4ml0boH/xXE9RfZAoATEhav
RT11+SeglHmt07MbJWYx+fOGMvcg9WG23mdOHzv9WBjQ52LehUz28ItGFEWX1yWuXyA/Av+K+k8O
rQEkYhr+8JdyditYQW91u7UHkraKGxZXJBNuyLxl31c1TPteKD3AUQcrHlPhJ6XqWtYttIAMH2Bj
3rUHytbC8aOQhhyukCZ2fmowR2ENRZogjp5m1ffMj8dGCCdalCBoxZWnjSa+2W33f0eoMGW2Qw+3
nw9PnwZ4ujTtP35f6C31XiONHtojdv5rAmjzCMGk9Gg1BeuB02BPy6Go2odTzLLIRpaXSn0VMiiZ
/yyMizlyOl+lT9ALKR2M+lcreOsuZmvumgXPs/nlIF6aBIdYA05IvGmvUaG/yepZM5FpugCm6Wzm
TNz0sL3kgZqPVGycTeZPCsYAuYEA+8EKr9ex22/69JqhK0KTQznCrvYbeGQaIU1/K3M4yz/PZyEs
6guVTF0EIWGIadWnVKlAftWERiuC3evY0FrabZqxhjGUGDZd3k4anmYWZsk+DWwtt9KfFM4a2AaZ
92Oi/5JgllTMIwTnaQNra+A8QAZnnUT7ObHY91xdwYjYpQHKNmap2Y4gmrpQDEUX1NF70itp2UzO
nexNioqm3TZ+vVi2sN+YqscmSSadMmNSLnIxBsZjlmq0aCUu5E5Ik014Lz0FbJl0uLruz1mz4HMI
BlBGOnumWU7UpHo35c1yCcPa7FXfL7YpYh4+LOUAW/FS1rsgD9S2geWFA/CkAyOH7qwTzmI/A8ix
oYLtLuGkavashTN0lUQgMWNbcElMCEyvENGUhm2C6/Y/9Qq54LIr7WXrpOxgpaSw6mzbgtRHmx4y
CMXDXKpXSeTJtksN0sTbDKTx7rlg/3/6uz+RHJ775KmFRUvIS1vxTxbtWFvOLt1VqtiDrqxkAP6b
h8kKlwxwj+5fleRop8W0N9hndf1bllG5m8K92z23cojKjDERUr9u8FE0QllkJIAa/YsYS19fRtGC
Qhit+SjlSVOgP5vQdtGDHOZeLDgbP9NVzzqjQwbFdWxVk1S0ygk3//tl5Z3FuHXoUuPbYjOMSdqA
ylWTZFd9LMMRb5M3olNHg2fY7BiyThjoezKzxuiAPYGRWUqUEVa03kegxax04cy004l+zrJrtMPg
46++uh4NZSMu1GQYA+JwPjoNgvZPofU/tBBqV/A3YehqxgF55yUOQCCq2TWzSlCUnn6cMJHwJoVo
8J3/JdPVcWrIjSf89+5sHW0V8kWc7nMkjN3zU+tLjXYBauHOKPTBYn2oryc+0ysUZKExNMzR9Ubm
yK8zIOtw5iky8FtFSjKB020uqfSi+gcddAgHdY1p3QOzbYJjaouzlF3H41mz5ebW9TSAn4ji8X0l
4Bz/3m5NKktfkTEEwhzwtSUulzTELvFoxD4QFBQZ46yXstHY0Je+N5oWtb52RXy6m0cQEyhhGxyo
WpRep0HhqKNLjmcNGOi/0km/r7J2f52/Dz/I/Y2npUnHSQmKSgyBa29wQGF5dWupdREbi+Douvwb
J2+jY/LBNYHv6ps/fHVVP/V5ZYoRU/V9b7/rqGpL5UcurxFCUNdB1iXT6Xu2P7ljSYI//cThTKjl
QqapwNcPXPrqnB+Ma+t2cdTJ+0xSYyqhXIiRN2kNJ+K9d9rPOCP43bO2jLZNtm4bNg3Fhq/PBFcs
TtWXAdlFv5t6527Ha5bdMYna8Zj9HHVByR202i8R2AseQq2dNu+2OQpJ0anFaLq0+6yqPBR7kEGS
3U5Rd4EOtbnCbPPocB+wWNi0SYEQgTZJpNIOMnbD6nAU2TIRnt29K4hQApWTC5LEoowAQbw4t2Zl
RnkShcz9xrR1biruGdo7H4kYLI+4wtchxkfWF4QGy/wRqb55KklPbHmb3zjQuKLzkjZyz/eH3jvU
1Op8XaO7/C60KYa264DFyNGF3GKhAkqlRLV/EZgkLJSMrNiTsOJmHwTBDd/X7VhfcyV6e6V027t3
W6w8DrTy8esKnyFRTlApEqJ8GKuCDOwkYA9vAcd7Q3b9reG+tXba+tKd7SlJdyKmB5Od2pfWHH9X
kDndDbZOQglUVm/fMhKdLAN+vKuDSS+NCQLHSW1r8TubxvwJfYa7ZOAra7E3pgqW/PdHNEj9DwmP
4J+RRjwSlAkXowYQYwq4+5w9NsHeZ+IVif23uAS76nDDR8NLBWvXqEQgDBBsTuWJ6lkozd6K1xuT
FlWy9XhngTYWnCc139WJbHZD/xY1BvPLDOxylwCpZ16NbYwcGIgaBSra5RJszxR9+ddftF41rS0W
bpNV2M9y/si4x+GG9panMp27VfAHA3VkulDbwEbalrOla4aBHrYL9R+nV/Jjjqd0Jx+sN1zeWicm
W4foWlBp9NarAkZZHWYFAPlLSZfHeU2r4OUuhE+XqkYhCdGLWibelGZqa7dQk1rNVcpzKeFpK2ff
x33jn9xuHTAk1C2TsEH9fZ/NaGER0SsY7ip2LblCmjrL0qJ3zD7skODNXEXzMFGl+s9vjQZMInxT
XAHTv6HixZEKjkYPJIm9CV+oT2XQTL343u4YWzzrfvgl+BsZ0z5OHxilnw+TVOn1WvAdFKunREj2
Jpo2Rqrk+e34+WM9pviN/tmNLi+6tqGg+KvliIrO6+qrAFu3ri1mDCr05V2JofahpKTUAaPXoU+A
mefEKk8uWLESCgXet4oMUETIHSfXzUhbM4pOzcy57RwbQQK19umpobT4lXwqd1XlkJ3hbE0deCmx
xc5n+GZzQ2hOQHEacNtnjDrcqS48QXSfJBP/qvbeplmuTYdjZVHXFvgpbAjKl9GWdaGNBFOz1dyc
xm90tnIxYrF2mF2KBrIhhvrdfywJPyM6UnFDAwvI6Lus0ebEE+LI6tKiMcifR0zTH0PRIHDAN9sf
dbch1gGArRMYwZaVo4Sr3F+49r55BWFWDdB8N9Gabk6+OrCW/OSOzlEc82FXySApHUyDe7xk+YTr
zDMJnQQPv6lDpjjyKxjdYBaWG08zvi3tU/1mP2D2dBimV2kKs3AbjFRZrQJ+wgCeXIPIsnjRfvWd
QEG0/NBFHswtnKvSJdRDYGDz4C7E30DQ7pmntBt1jnZySNsLQpBVSzxSzFdEXPuf3yeizjoEOUwb
KKPoWMfV5xBIfzXeCs7orYUXDj5FEJ+vG6RPJQoZ6hkqtH/NZc5dxs1WG/WgMd0nKlpKL0RIk1uZ
ZKmQ7JqkR+FK6MltFWFCPAMM8GxTG+zNnEli9fQCReH87xZh1NdwPbBSAxIW60pUwi1+SKpdT1hB
9nAzNdKOny4H40jCNZP2AV9jrLr+ftl7qIQGJWnz4HqP79QP3HKsrkK9ogQaXzYigbtcDtP6P4DT
g0E5k/oLdRgNPNimqbI9rZu6yrdakWmK1otH/t7y7VSjTqAyHJS0h41AVkXVNuq1V7KHNwMXqmtc
5wxDWKitchOZwtpCDCa1xGIu4Qhw9okC8gsa+n6/7PrPj6XRngCYBJWcwsJDwE5boXfGd1D8J3Nd
zEVf6gA38mQIJh5LSRHP6mozN6cDAhHBaz0vAfcP5vh0uX+g4seTIqg2JAQqg9zQWcm0BIkhr1ee
fu67ibcPSNCzOFzLSEghTWzFD6BIpIGVtFGGeipsHeD87Cz6+eLwW6Q1okud70vp1UoSlbrjgUAp
ewZl4HoPYi7KNjjwpDXtUsYqsYsybEKjCs9UkKT4PMFlwsVTnT47XewVUrXw1/Pmnhk4qTvVHLy9
3rzdS9B2xFRSIJVdZXja8YfIjsC5StxIrF+L/r5eUG1vyT1D2Vm6DYR1RR1Rm5wqSaTcxzRtwJI2
lMULBWTdfnbYNJfN2Uznnhn+u3uN2dtS9S1nD4dm68TmPqlS4nl22AqGCCnwRm6YbVIfKOPW/eV/
87ogtljmdM6Rahg9RRU57Y5BeWBRVT1cmTOhrTi0D3tSgu1Ue1rE5tK/dYTiHKy3CMhqu/DY+KyS
vZnuqHIhjYiE3E3BonPavjRrO394hJb5AnbRcfxojbo9r3wOHxe7XBH7/rDFXQVB8fMK1d8W0waJ
XTXT5N0KtGlNX+T6XJCkuGQkdCuyGWownkM5CcuxkmFfOwo5GuOi9kvakiBob7z/QX+/HqfxVOrN
xSns2A10pIaXVzJnQx+lhhklXnt2m025nWvOl2gM4Q/leKYfT4FKDEOyNfC2Y6o4ZxlhHutUYjW5
csV1HXBsmwzGz52NZlSj8Ba0fN/iZmfA0l7zKlmTXxIhRXfme7gFC10xzfKRwmfPoKKlqpOqKcdS
lW/4iz+vcK0pKstgniLS86jxgSYxspmn5Mdbwo+HqXYOY7db1/x3zycwEFuzr2ix71LFfOSyDxTA
iHwrxVKR0Zcdm9yrfjWxmNBkdwOU7ADcEj1fP+v//L70VS6yD+psVKFzyfX/mNK20gq/6MaqMZ7J
m7+KQlpIaU7WEIdBnFAjXxi0cW2KzGM0RWuCxruOnlqlqwgn9RciGM7x61diJHj7Y8CVjLw+YnRN
JDiwoBCyG4wgy82cILocc55JzPOkJuS6q1bzc65F3TM90PO+Pn4z3ghi1ZXgjebEmEIV/ZaY9byl
pK1cX+fOWQDI0m3o7QmydOESOND+O3pxg4NzEP0zYapC1eiq75TiOPTWsnpwvvar/00iA8rDYpG/
svLxfQBoQsJEQd+2cJpdgTVyXmBrmJDp876dPjBzUv1GQ200qU31e00HKlEJdHRsg+jaJOWJ5t2m
i7LntrGe521/yuyMyi3+skPRapZipEooqaZc3EsVAZOkgOCEvxvrdwERHfS71sWz+aejmXe7vXqv
ELy2wyF1nIgaSm1M4g1vZ8IJtxw4alJ0y0YGgjjcmSxzYIV5jJICuBiW0+LX4Y7Z71616Zujtv7/
4bW1cYeuxYoQq33RUgP56Zr/TXJhWajDneSw7/QlpEhEoLpyjEHmb5vMb/wcHiEKvSxDw7aHTYY/
XJciigmExKpf2HCimbJcjWqnFCSa801Rf2u4Rs43KhD/DIlldyOPOR4mK1ROJ2pyhif0dZa7e9/o
kNDheBYSZNMcJ4i0uqsxT84c07HukjGFwnfbN/6TscZImVX1i8NNBZz49MFYMvnbDwdiKk982meO
xSxsnxKo/a6IEzHNhgixseHjgvvnY+JzSrPydruY5N6LjDZRoilyRSCq2csAdYq/gSbgWUTHn+5u
5RZ86Sp4ctP8sTSkKtSNqpq/YDmrmM1UuL0i4kE3foC4f5tMgsc03vBOvfLWPVKzSddjpfT/bfGF
YptxiQRkT7B81pB7Eu69nhQvzXRpdkhJxu34ygZSGzSK7ZsImooXKjpSwbNJ0hxxNjzJIjbSoh4K
tk2PFOot4rBexTpWm58DeU/vLq2CzjrB/MaOPBdW9fUMVlp9CP2HQzd/BQ9COQvHwY55H0/P8oKr
C/IJU6wFqANoWL8/jl/hLs9DSiqfSYwOS1llJPAWEH7qqOH7/085keoSJWemQXcEjJC8JozFI3C1
o+1sdnXFM28c1NcWKY31V/arTcKxBKoHPPBJD8FA3LyHnCe5yEsuSkpVVUh2XUufo7Tg1j2ulfX8
seyqWMyVWz1QgnI3ENiPluIygm1zwm5hBKGGDbn2tEuWGGodsg7vaX/oG2vMKduzf8pLR7Lnhn/T
qOhphCtAK6oJ1eYd3I9hOKfpol0LdXWRiE5j7Ok9yiFq9Kvh12NA5IHyEf73QOOhCm/T7rO2/DTP
gWbo9520rkrhJ3sHWMo9wO/JfXWxKNMPD7KrzHU8/A0678s/w7mdp7wiZ+EfgXut09UVjH2I6FuV
g/6LkbrcbigYaw1RD9ydGtUm7dTshDXvx2+ebNz2RZ1f8HraaEt1l1UwNmz9Q7z5uLf1Ow3tAxK5
tWkz8p1VTk+mZC+5ScPEwBbl3IgFuH1putbby0avTnGVSEwfS4z5BrpO4uk/oyFHhD9qh5kzQ1bl
zBGc7wkzWxYWtcRXzrX7KKaKj1UqupSlUAYBpCvyZgPjvPJCMlknaBrgf20rtxqpPaQ2m39aZmTK
Fafme4M4orZtN8jbl0AftNjpwHdg2CKciaLqWnrSkXWgDo1lXJxt3jC6Z4xbk0u6GoQWHnD9lD4W
IJk/q7N3np7wLjhRxF/i0LSlkAFifbY3yP4TOX4oBq8l2/mXwri/1oULHC9MUEM6C43SOVABLS6q
wU8VyhOcXtKzqspWGj5LyV4nmSAJ94xZls4f7AVH1DTPi+ezM+gArick1ouG7H8U/GjZtrAZJsm7
FTxbuUHUcESbMUrSCUhVH1c2JTK0ryl9IqOm+azL53hdM4Pgl0xpZ/mORxc4ep6zU2cZiDugl7Mu
JoJnlJiePf4XcB0RAB4dtvspVnrZ8p6glXaq393qBjrSX4W8VnJ46sRQFlQr87hsPtQtkbufeeA7
M73LgbovXls5mFBWPZABgFHtGyLmp2j8ms8hX+Yv5cEsf8G3ev+n+7KQ4hg75zJRgYuyNFWG9Lp9
3aMY494K0ZRW/wcnd7KT0i8sxClULWAFuwe5UT87NcPEm14pm3Ye1n96LTQKZM2vV1wZdonCxvw4
Y2A+24zXKamFbF/P+PqSixtcTXFlHMTINIfV4CrhQ1ebQliZPucxvfoFqsZQ+DEjy55sihixY51x
mFy/S1eh8574d2RLKTpoaPE5WfBTlA/8eBBM76ZqdBEqCNx0bIj7vrn0CZ8sszUDBsXONpfc4FqB
ij72FozcPHg5l6J51p9ABoMqCNJoS2qncBgYQN4V02ly64hDEq1hhA2IfNHYrmCocJstzGWBUqvO
/odbcCJpfK+jI9OYXeEHkbIif6jqCXtdE/d+4RNielwMy/0T0ezg8EpVrrdI9o4SEz2TaiBHJt8i
2v+GXTLaRo+J4HfleCvT7YTWShUGFaOe3CQgMA7ZxJA3Uq8vf+993NgbsxPuCcQlGFSIF7f0QDZ/
o02vmVJLVdamze0dVKy9IdQ/ycuMmuUgzeb8rrbJH1C2CzhZvx7hOvbhPnKgF9LF5YedS7sZOJ0A
t1hfzkgTvIxAuAEsOlG6/gyF3GAJIKSlGITznN22S5ZnuNTNBLl7oWW+msGh0yeibCl1omkYeydh
WuR1GdMq/zgkxjOU6jiEgl2ifEpAu6RkfAX8TOVAd5hDyldt29P+bRM/xAqwPO+Vt9AvGDLomtFi
HLeJr8X9+YisHG6myylYxh5fHPqMe+oJmBXqoDagbzf0RgDm8HSWAJ3R+pjBll1a25hQDsKd+Fz/
LCPTwg0oydMUWex7EWLlQFZCj112zgjAEu5Ijsx5tEC4coNtT1O4ny8EXGBLI60hKLn/so0pNrJK
lrfCrSIebbbrGD47+JMJyfJ0YJk09zK1/5L3OoOTlp4V04xQs/B5VDtLBHG8s4/FssRrrz/Xd2n5
VCzpHg8Sg8IE3QOm6n+Ky/wp/9yAZ20NvrrnbLPCK051m0Rs0D1gVp9mE2b9eSJ8gTsFtIOgXwO7
whGOkzJWKfgYfCfw+QNTIJW4YA5Cro3GBN0rNfgYl8ZDah5pwJxsaiP8FBV009DV7ZhyclAe26hx
gDsM7YXqDY/3WwJbib7shyi/0vHSz5J1n7rjiWN0cI6jqmsXshe81+AU4NoB8Gk0eMk9yZz3oy53
54CnkKchLizZR4JKG2e6i/DIKO6Ahg6Uee/Gl7z/qJ5IsusgExsAYwVitDN+8IEyg5Y4bRAvtM+Q
2tL1tEKbG9KsxSR63QEeRBQE/lvfnWuQlZ3Dd5J7w4NlB1W2zPj+TelXlHIbRcq70ulh4GBZl2CQ
1/kYtvtNmAvOa5y/K9QqLK9zMG4+r7X/jnw8CDhWm/jmqAq5akrNnDREa3PFwnP1G0f7qcZFJiqV
WfLsafpVKYKASu/P0fkiM3Zq0tgLau3aubdpBCdUeRmiPi5R1KAge50dGioPESBtWJcnsFj8oxCu
gI0ZpZb8twMSgM71PlJ9XpprPrPMP93MKpIl2yY6TaVIP1SDeYLsB8/HkLuwpZQsKvrVDWpttuRo
hm0YsikD51wWXES3JVPA7ZFrzwXowyoDW6wW8dPqZo/09LMDVkCJs/2a0qme3E8xuaG49AJGVaTH
AMIbI72ghh6YuguVnuktoeheAXQxFgA8P4PKO0WgMZ2S0p5C4YsJ68H6ofhuIhxYizEOuGfCE4xQ
V4py/Wy386ZNfcOyiK1l3vD0YY6x8AufMQmQDeWdnZruAbU0OXTK3MjvMxLGz1e24EYqCNV0J+EY
SSHHW5uGGWTVWLS5sKsjoB5jSX3w6pBdCqkbLqkM66/Ir7OpYVDmHlmiCpv/yGcQu4C9Y/sScgI4
FbgMKAbqTJxuDEFlfvOw4PmlGKvJOJYatO0iPV4Q0nkDDAZb/hFzlgYmx4+8rotmmPDldvBYqRCg
LOUmkXURkIgsqa/G/w5plpqJzyAp67Q+b7tsP+9x9hUUyjtMCGw8tFhUvi8rsKyc/IqZXBKNqnYF
a3mUsD0h/Ofs229olk9d0mjzRyoOeEl3xIe27mHYjvXMsAY39+8DmwdbmlePQlYSlZ9xvTcYfCv4
LAUfxe+CjKAF1q/KDZPLAtUG2qhpAmFjDaFV8XIni2cINkWRQPTBS4BQZkQ176hgVwdGiDKf3WnJ
u2z/gjP9fvCmmSDPuwG5MwYNSFP20bTcN9YO3O71DyGHU8eCqt+eWMAnzkvPCrurvhmNalniM7En
if/RvkkeS1RuotsYmg1ju86vxeGKVPJ2LuPLJKFjZhzJ/DDf+Mo9cj8M+QSdYoojpFB2juIW8vIE
ypBST+mszWmyNsF8WEWsrAbo2EXsWiCxo/KYp68PDtbGaOejVaAJU80vxEXb5f29FM+A5SIxDZ8D
ybx9JZzXnKT+51Cd7beoJIgrMuEYcaM4w+gOjLs/hikYJnHnCiB38ZChUOqiO0sT+w0WMXg7C5A1
y0LVH7fcvK4vJ0wrOgLxuu4ReuYAO5u1Zzp+emFLR0Zx1CBAws+BX7i5xZWzQI38+0mg9s308qG3
J8yuhO720G0Yu9ScJ2Cep6Wwj3qvNCrsCnEK8cm9ATa/vzueF3k0ntayR/Grp5FLMNhw79qCVuAO
nixITzjQoJruOSQbmiV3AL/Z9nadCwnccg3DupmRXiM7Gj+vw0NlkQB8YbW+ylpb51FCk4lOFYYw
lMS2szmJhhcSG97HAoShulpkTjqoiOkpcoYxOKHs8B9jUSwCoNN3lY+mLxxInckFJhNn5UbUhwcS
ph8AAFfKVtPtt5fUtCgsds04Vzl322ii4aHDolIEVs+wZjpw2N/JVpti7CWRsXHx9RIlyspRhMYZ
tl3T1IsTHFPRqNt/vvqYX2cBEP1Uv7e6eJ81fk3eJt9fse0HwDmSB4qbi/pYOCaZYcz/W5a5PrCe
821rzXLr/gluV3UWj2Wty6e7+9nDE5ozR6Qx1ZTAzw9BcU4OsimY4+IdJ4OExo0t5nt1bpqjFYlu
UN9M9zbGFALitQX+hF12BmzABcsY8FZwpSOH90G/XMDkJh0+HaFzTmzS4YDgZuUGDZRCPelcajTd
rmFpIEWjuRt4KF+H9fHx7BtfVSx+FSgmJbVN+1DZbiuPUa+Gsg1jeMHium+Z+ISgWLm0ZoC9H3Mj
1dv6ENztV+SlpMWMZ54mhizHMSOJ+DB+l8JPb1tlXzz283TzivWUticFHtUspg51Czq5xSGB8DN5
xVBtKBQPi84VRjzkUl4ENAMUfOjwvw790FZ7gDaLs0o1XDBD2uSaC+TH/0aeR4IGv1Hc4W3cJZCY
HS4MiS48lWfVJaTW97NYm+UNE+4zJacZt4+ldPJuIx8d+qSKA+fuRn6+JLfESlL7+ytlqOjA53kZ
m0moaitvE+7p9624QKZsnqbhugB16yOMi9GzBB8Fo/fpmr5wVcF240w+j3ZQFmAdLBFDahiW9EgF
it/4R34eDqYXph97BgzoAwkLQJhnJb2U7hhcKLwWN1hzls2dOuVxBh2PG6NhmQ0KPUFWG9XYgzJx
k2hDqMHXHQNKq9kjeSh3hpsahfOj0n9Bcmw7ql7G/TLgcL8CqY7l54yZ6wE2VO7sBxF5tvuc162F
5CYa+d2Ml+3fAh7J3MHRiVWFzDmb/WLTrgtSGEpS5+79jMeXiQCYkCp5Xnmlp86epcBGhhj/DwQK
r6xJ7jNheRWYiprCBGEzfii2IQKQvop3atu5zFgCSmqZqSPv4h60VD43Ru+dKRhXZS+sC5szCeHG
7rfg6uLU5l4+NKOPztGEsSm3gVK68b64ZkT3szKesvWrSixoFvMK1JQJ+diZKddinRcM1TaaZpP7
YG3ZT4CR5NTezYmHAZZnP7Ck1RMidT6lROdOS9Yu5BoyfOBTlL+st2p7kzaLfcToJPwq6jup2ZWp
SwkRADTyZIvsJcSbFcN5Z66A9riHmF70huHZErj9Wpr1TGdUbvEiFUOO+BDatHSjbhKpbEeHUm0b
DnQylcGONuAF/AM9uxdTNe3XUCrTmyZNGXm/ybMm1OZkec7BXelDZhnYJyCoTabMVjpYU5zxtsw8
v18+LEkwl846b2+LNVNB9EzGbZaz/2N1Pu9iOpNeUPMQBNb67JNb9W6AFYBR1gVZ0TAjjTmVHtlA
5fwR34raoekN48sLo0mJrqZx5pSLmFtjq6zJjrtUjFxkTRiRbKRSFU5KY0ykS/f5JqITQueO5mKn
ZBDksSrK+wKtOLTRWQwFukOVo6R0hfDI5dkBqHSCtZIw8HDH1nDDDGrjZWAksmzkam+l/yKcnz0G
HUAykOOvAp9/ClHXK+t8SiPOTeChy2lkR27uBrejB/fBjRtPcdPBJofZxHxbNeA6fnlaDSH+RulA
92daRuFo0d5I0Vqy9BM3HEVxgVjbv4SQ7bPDPWt4y9p8wzzwtq8mp2W2TEmB6Zyv+Q5xjTvKNf3r
lnX1sNelWgYc+OgC3o1BSdQCOsad9VFv2hk+50sq681bgQsIJenS7ST7PtOrtBcG5MmsLcFErh2z
8iR4tXPomNnDMLdfiGK4BiOf1/Lsk1Nlq4x5qOmP5saVfP5KTae0xZxg4PGTNFf8G+WIGvGmUbhm
Wj5GgcobpMvoImC7Y4XBX8b1ZziGY/eSI3paXcc6WCXCNolmDcOPdvqx+IXot79MRJU1DvuV27mx
NQr0wKzSuLPRYvKBNRkwFFG4eipNyL6pyf9q4CmL9Jw4JKFTmNCoByUqEshHOAKNVO1ULNimm87D
LD3bDL9FwM3xjl+BuWAsHxc/tIelgfvx0dd3y+CW7mxXPqMYON88aR/ZQgmBL+J6n+ugxDH3XwpL
ltxmchYZbJa/mOiG/vz0F1zA8IYlIyhYR9gPG3ETAUBz+Vx839urpl1Tc4xqrSx6hw+qyphri0rr
GiNHoZHk7dm39ObzxzaiA38EGHegtv9DZcIjgV5hqqeophEocluaFyy/4RSTE10xgk9rxUoPMdoK
SczObthfjpgHEP6m5etCcxqWnJCaNB1KZ7LWcdJozqazlMjmE+dEKaH3XPZDrKmAkCMjJJvNqR8J
3MZkI2vnvbIA6cN4FiUKBP4U9xJ1HaKbTzAsEzyWMvNdhBKxBEz4iS9QFi6Wk2fh/tGm0NMcML7V
acYSNbV3Nb0jzvvNkMdAEMlMDeV5DiJYNYxZiFk2GvF7lic/AXToOOtaOOLvd99NSmNu38m1joeX
ukQLlsCjcMOiUvFnh8kw2Kx9kc53wB4NmpCxE519IA3yU5PZlDQFhgZK+BwB+MKwebTqgHdUPe24
DX8h7C3uUaxC76mtz+w2etEn/DGy7QZAPQs+a8bGtR2OY6yW9Zte+oOtCOoiVM0u+ADOsvGAlHAR
gJeBIF2FbuMgw9MvLaXqIDQIatKoZa+CavEktioknC8DfHeXdABtH7ke8sC4YB+DSTgZeUzY6POh
3p8kirP2crFQaGD4tZ85q9cTLeslePRzIoGTgFWeU/rH1Th5Sox+EalOPEVKxEDmYlpDe//7Htrj
0hP6xUBNMZuWEpYoItlanRYkfscWZDfo0cjvdU8wbDoPzPJWXa2hnvx/VUiYleAwLmoaeC8p6eg1
iW+7qrYzMvG4O0tc3MCxPnEI3CT30zje+i3kZ4bTCu3+QvhL7UBwl6dbmAQxZjtrgFgN5u80SOUD
rrR04nA6bzdMiuyWhew8OyHmToCrufT20LaNMHJodJ6SXAzyp5Xj0/wguOtgLm9Ira6zDOudw5I5
AVPZRmpM0WxJ4kQwSvHQwmJiIgC+MppN3UAKNpRtJvJI/k8zklJWqNjhc6Sussfew2j2y5P0Q77V
E8XulQNqTWj7ftDfw6xVLVJ00IvBfXXjldoBCqjYjHxifOtzQ0cQU554zNLmYuo7uOWXeaKSue+h
v7JopcIYYBgOO+/35lUZxh5uPgEIr92QxKP/JJdoaGkggM6dKDRaKXAYc9+2/0FU7oQdyJy7/duI
gwfnG4d2ha0/PdBDLFS489oREx8EoIkyM4rn+bSCtScBftD9J76raCp4fqOsYY4WLK1arvXSDJES
ANypD8pwh12dqSOR0FWje+cq8femejKI3d+xvHilooOQP5GCLrDWNeOU/gsofPk5vOpgB6gGmzM1
UrFKQ/Q1yZbRcfcJxs6xjjNtO2YN2N/Aqz57/wxAy1ZN1Bx6TD9b3X54fi0/TLTIfPO64+c/jy9J
0Wugs9EDgaqIOEUFMd54yZeCddZuAp6CjLwikFohR9I4LbvKTDPdAm5ST3P/sUoihGKxumE3yRX6
ap8btWkQnIOi+crIswMDM7MdgNDwOcanFmjlfCu27HaR5RbkVcCF2oL0p2wiKq85iMbD3Lc4Sr5U
p7qtGSD5tyqTOR/N4fhTU7a3uAihLFiAJuOIuJv+opmmfRXVY8rgvB9Ay6kL1e5cPylaYhSABWtA
Irjk3BRbzU6USootrcxLw5Lzi4s9oN8DmK1d9stOMjr3J2WxyRB62j3tkpMS7Iv/Y+N8p9F2DK8O
He9N8m+vKfbpbWTQH6R4pANf0ZCkLH29y+5QRsErmzktGWogA0oHrF1IlNn5TX0oRvwWJ76hoz7+
PEMsdiMdBPMh3uTqVWky6ws06AbBKDVCAVF5ZTQ9aww/ozWwQW4Ws/Rj7gDjZWlqrZ1RnePotJRt
053tYgMTpIY1noZPy1cuFUjuxnb5PSmKGVAAWHz2B2mdkVavuVzOuNempLIRFo39jve+FrYFkOd2
DYwFy67SAxKc+YuwltDyNq+xF0S8PbAx+H8Hk0q6L2CKqY0WuK/moTOO4tVzxx1BXYRd9JG/KWBG
28nrBuXXWRPcgaCc8E+wfYQEiAB+AdSW2EhIu9Wy2vmwa4ziKdXpd3M2lsAKvccPeoVAxJ2+O17M
Wv2RxcMLkQ4jsVVN15Uu9ormlQQAnPnre8QY+HvwutFNU+ZQhOAW5WCZMQYo1oXmyf4CHQb332xp
KhdNF9nUokBZ3CwWufTVNVrIppFAz/JMgSAPEr1aSZmPIh2PYejaBvXDbnLroaNsjVTngmDHuZaf
j0dtTQpwWaH2KrUV5o5j60u6YRQ7TYnhWayt6v8hD7N9rRbBUM6JQjD163F7idA7Bdwjw5GoNzqf
AdM8KhNbvVWswnUMHUaZcv5Pz1hk//fJY0fYFS5Zyc7wgoclDXXIek0arRe1ZVHkeOvUbk8sZliG
uieIxTOGhUUDk8M3i64rDRkiMQSk43nYxJkKIYxKEYchXm/rSWV4goVSifbRUOibM+GE3+kMhlQh
w4fHq1YTHfcBoxw3JmVs5G5d0qOpEQ1+8nBMw3lBej3IgVvsdBh8SGkg/x5v1398tA+WpVZeSPQP
xLK/hf7tdhJEaAc20/0vYQwTi3oGwrn3xk65aCRPluSt2iiZYVqYIhJ4gVqMkJbAszKoEvXHvoBN
2jo/bhKT1a1NYNKfzoAKaWcvzqg71zk/xMbp946Qy7OgQzEHILjUP2Ld9U9y+WgoPe+wjGN3202F
eQsTA3fmj5XL2UDAEXnjl4LVKzkc7j0qi/Wo3Xev50nu2nF1qEkxlKnyfiYVnxpYggrZUjGjmOJi
NsR0+viZrcTKIy6/MbB89aLRkLrBhsRt1eWuYNK0k/Ib0CifONaGiX3nz0llp5dTlBT5wYyAKN8H
WmCSMax3Yl9k1o4PdiDbUmlUWapKmrI1wyKrqNFqBX0Jp0k1X5iBhweyLlzW4SKo/c/rIBNAKELr
ZZV0ifeHzsjtHGehk6d1ZbFDZd5WHBKGU6BYB/HQe6tK60eqyWCD+iJsLBM0DXsBt24GLlnfQV5w
8G/g6XWWQvgDwoQRFwDJd+8QithdC8AdHPO0cE9QTBZNTg5oUSaDqLqjq7x8M5kizRBYfBbjY9nJ
t2n6TeRo2VLmsE6TyAVq1+2JQUJ1Z1H8oukgz6kGshrCz/KWYLU9+JjcQAka9u+fVA3ROIR1Q1GE
SfroKVC65q2sYlyDTnzsGDw4wdlrZlvTWWsEohO04t6hPOx+FYXwNASdf0d4Wyrsyy1yDj/2dOKC
t/EL7yKsH2oUqOZqW5ljtgrYVaL4xZxFhrWQFRqbrLcpcJu8r5no5c7089KWkJR82nf8hQfWZMIq
ZeTMDONp1WnA/M/vSJmCLh9B2ZyxSEGgsPBljHBYp83lOeBViQ24u8SwTLVrOb51g88taq36wGxq
LN/xWb9qv5ta5pcAEA4j1K3KzvCnTwX29VdMZ8gavGdOdLIdNnapd68egpnBMv4cLc2xy9C0VLfu
6cxFM5yVoQBTq6MZtcm3lOQ9OQPp7gH3N15uGzkm2iTfaydCIwVS6UPRq7U9j+NOYxx89rR/qbdk
9HFOQoaD5dk/vqTalm/ZVYXRuWLqrHcMl0jnY0da/AI6hVEvHsFf2m9xpShN3bSH+ByS5kGpsnyC
xrF+PTqaZtYukQCt5x4Hs4sB6u5RAS1/JH0NwEs3RhO29wT0//zxGzhBhqiKr2WrCa3L5b8FZBjA
Yqsq5Sq1VVN9G4qZgtSfkgEvj8l+f5Q+eCu/1JOYAZOtZLwPUJrMK0OXLsyHXur76uKzODzkgznm
T4q7Eiv+0xCQphUyTQROn4jKkbWR3hwdT2UZdUf0EUSgu6x+U/qDPEMtey1MX8M2u/DM5wKdeb/G
KCgRLY51RNwgS2Dcv7BRRomVq2lXkfPkJa72p9t9cRnA3A2hsJ43tSldF6D5pDRIxL41UitT8ok3
zNxmS9J/SqwaprTb12zGxyY6pVMCFQc725mNB48BrJaf9EecNf5/U4Ne0FDH7g9FZMA0PjguohHF
yfXsw+neMQZYZS6LRmrGpNUtDp0ik8kz8O+FoL9d4X6qElF+/SsnPY2W6V5NNiCSV8nReMyXguQt
Z4uprAADS5bDFRPlz/e0P4xb9AFGkQGjBPZpoX23Fg1thsEw0/LsbMj57875d8XrJyobpEEDlqtp
5kJvvKXOzFOnUbUR1LDV1CsvN6fgsuM9GHCV6Uo0/uX0xNgzsjJzvob6l4GY/XZpT6L/sMFNPLqn
1qkhyXVUR8y6gcplDGqv3F7vHKYw+v1XXVZHkfXcZJxdB53HKpFBqnpGMIUXODYUuvuBniR9Xq1W
tPYydCc23avvSgZdK5kLM8ppFeyalVswKHzbgz2amRVo9E34OhV9OGuTlHzQRQnHVFugG1KYLXtf
kdkVL371jnLoZ0tR114sKu77gONrRupvVZtOSPrii8e66Pxc8XTpWCRb90S7ME/3n73UdQeTWbzG
wjsrRTCebNz+qeF639LaWC6+pnum+rWywm6JdUzfkxAPmNxxTKubOfFSJzcWyUru7hzwlO/EQ+Om
n4XWcSsWD561Kdu9vufQN+EvPjKB/Wdp5iyl0FVg5FeVy1o1+mK8pLj/CYucuK4q+y/4w/Zfrj2g
1tondzQZGxR69B32LujfXHhqP5saqp7y/hxcHVFXp3VTaTS4asYH/yCN+3pgqPfUy8B2Kz5k1uOR
6R17ELHDHzKxx0q3+fq/Jkd/3H2pTLlmTeU2kOv4mEUllSSlFt6WftVD7AJlwnIEhwW3RsRE7aoB
rstHjtIWVeN/vRRjEPWW16CIhkMc1Z1YCAAegFo8hdPq8yMPDVjSX2czQc0IgZuOCFQcZeDxD5sX
IXudD8zEdMq46gvsyXZWnRx6v8y+zz9W4vnsn0IxoKNK25LMjUOEwGTcbvmql2xYfmXg036qs2XK
jiRCqdxO2dJJmay7QJvjY/e48YPZv504FRgOjkB1xZ0GTtiCKlzubqkq70KGevOlw/OvKV4axuwR
wZ7TrQdNlpStbQFJHDkiq/A4zbf3BwoMbm/TV2DrNA6QM4gffsGojiCaEwX6ygB+qiswgW8NqVSo
AdyPbWfCSY2fi7Z8KJt+vbvxEpf5VHQdipXfNolmlyRuCUndCqRRanFoCQjPTTFhSLST/jkbIQvP
LG28f7ngIKyPy/xzsQwpGftjsKz/qYK/SB5QgjFMf2Zro6HN3xNVtpqaDJuw0ww6DDEFHgygaRxE
NA0sPCExCm+GDENZySdWPS+gWiXwMNNFnj3tMVfjZPgpxV+S29ZHOdK3qik5ps4BW1fqXZF2srnv
3f7nb5EHIPA3s4eCl22rtM/F2oAZJYmLfbuhKjW3/BZgpqZ/KoPni92DR5THLU0k/hbPmfc8SeU5
uSoQPlf5PhDnP29nhiNOIfbLiiF6wksKUGHkWos/JFKs+R+dEWef3qo0rJJ9FpTJvMuPPVtNBt9D
kUFG5wn5aXoeEAaYMZgwMBnPvPeMbilei3+ALSzbtGaXkwaoSHn9SfYvpYdZrLc9XNbC2L2srFD3
qeEiGETBpYwgwuruTVYXFv/C8HuYhjUKm0rgdKyAsaQPnroMKFanQexNRFwIWbO12+49XC8ISOQd
tMazsAwDLB+xbZyJ5cBRS8xaLAvWW395YOeyD0VP/S3doc71jXseYfgM6s/dmxZU93f4W3jzj911
THGIgtR1QDB8JXsxX5+dRiyy0gJiKVq2j2gC5+wfPB5zlJLwLAjrYt0K9QeNQPjX3207pWFbJcn2
cx/9CiGTSzDQzNdMPdy7lEkrFtsTgKP5Hx301Sw+d4I/2M7cdSvn43adKo22JP8fV//hl4RZCJzW
p9Wshq9mpwYOiuOwe1x/YiHTLVNwDAHog8YsK7SXcclhLG7ADsq0erzXVzkerY4WF49HvwjAr6zr
odUS24bkyc8J/ISRcoUPFNJ/0jW54OfYODqN9QNSZSBkgBHv6dcG7plCx3Xse+o7ZjjxMDOtvtmP
m4QCR16qDh9zL0IGN885VVIV83w97Dw9vAYUA8TVSUx5xUQz99vZfM0ece78G3lCntnGe7rspJ+C
wnFMRZIlYswtbYswaTqBzG6BrjN4aZxG5wRvu2t2Ohbrcf1LNG14VXN/nqQImliUkvV2R+UuodfK
89eoUaFAYnv9uwjoUukmhqYbBCBMLindBxrJBjQpsa6/uNES/D7psa8nOonG/rapH9mDUehqmmCH
RnSSMhAFem4yZsEhUA0eEKHbFhIUOGFHy9Pp3gNXuth0UrfBfix+iroXEwEzugCAq4BHsMRO125F
OFOyT3GPLBiGsIGnrKJYgGrYi5rJQGwilxRENoRLH1JKgfCIU+O8OenR49CmeaasQuuGASGmTuLa
Yr39Qm4OYpGE5xRuW/m9HROODiFWd2iuHuZcppQYpCVBuFrkdxGySVodLwCBNGKBg+eRNZJMnIra
SiQzrk4YComk9jfXekI9pP1kpGOLdLPv8nQkCEsWTwy/T19fe6HUPJKPHuDS/iXgRS9fPH2eNFQr
zzBgbyIgsrXrMTeXePIa4Tot6r42sOiR79mL4rl/mQmUR2+lB5AkoeuZHgHngaot+BLgh9pwa3aY
ApDLa5zsqbLW3SjFF+pJqD4T7yjhMQusU0lT/8MfQO52vLS9X3ukSUZ7XqrwSXxs1DvrfUbieSUW
hq34h2R15/Ub33nFlnm4c9afkMc5sHm1oRViVMA3fhUGFCgWPnOnNcvn/ZrWX5zilqKO1vjp93g9
zhO9Cri+XKNICwwUOnW5WEqlB3jl7j3R1JEsbCWIxb71owAeo9R+zHRwIo0hxLSnId76yO7mKlp0
opFOBXocLSJna1FkFAFd1jhvdccCkGGnDGs7IMxKLazwA9W3OE+KJLB/v2S8quF7llXaPXcqbBfN
Zrlcns0HOUu/2Lz/15CPbhaTVfzuRL561cIn1qGN5x1KCKlmHtqMaoIXsH489V1kGA5y31CMabjI
J9pJVov36fOosX8D2/s9bIJk8pe9iNDiWfGxQPXH2GG3Do9i1Cszs5gT5hGTb42QaI1mWtGe2FOZ
1DX75TrvUJt7yE90VOjrwot4X4EWc5oxSjCFDLrAQeaCgfOs5/8lHkS3N0i2L8B7GEFQC4WOafkx
QktCAO5J161XWUDNgoCJxfNhDr+9FHIECVxSH2gp00iYUSbNgL8QXohg7W5vbEtNK08WZsIUv7BO
SzeBUeuh7hXAENi3xxjavIjx8uHmTbn5bRzmiApRfPgFFVgSm4O1rZktrqgbtMT9VPGF+L92reLp
jNf1KaOkGwrU5qaRS5LtWwbopkzjqq/3Hr/QHaAiR4+9YBY+rSubC/7xAB6tWG+m/5bOYYyreDUZ
K583778wHdyfR3KquMlkzuqsj5hRl3Lt1oq4JO7Gz/YCeO0jhBu84J4/OhCDxAqdLTo0tvaaLkvM
ZJgW5BrcqGmWVC/geSGSkd5+Z4JbLDZ1VjuyIE0qv9SoUgEGhbnOs0Y5jk2/g9M7CWGqtY2GWR+X
Yp+LEyjxxslgDW01O74ldOR8/Q0XjUrAqxwiyDdnd53NP66O+mWgOxK0xeFdzhqqJl3KCjbV0GBg
TmjTWbcv+uSAcggzObPHJ85/zUacz/4zGWr0/4OLeRkAGHf0zvhLRUI2S+8C9/K9tm1UDoPa4/sM
rOlr+FVSCZYXWdfzOoxmWgIgb3dewbDhXSmkFszePB9bNE2B7sHFCW0KvUK91wYHia3gKXt12CmN
Oo4dFTYM7wtj6ExBT/RbrD6BEzgdpQUPJN0BFcCURKO9l302XINt1KmL4n5TtkLLMqxG0z5lEflk
9w/UfDkq7vtrA+EtLIideEVZgDfnE3ZI79x3p/3KprtuVlZZJb/y5m0lwUqa/EHpAcpTUcoFChZf
ydyCZNb8MrRYt+ou3JAVN7S0qmUR9O/YERUqSXMjFy6/7CC2an6naAtqzTmiXiVtZUW9VUHGd3QJ
aARpPYDfsN9Xoyvw83PSRvRu6SM3BW2lhu9dUgUqMaZodc3iTufoCxJWHZuAa/VXc+3daaiAhr80
BibPSOt52eSH8uWeY2JtTfZ/7zXv8OEJpQ5gPdTZgCUkT2XV8G0TeZAHdgxqFcSWVWI/e/T3upe0
JRVcT1E65Wzhuk9N89zAGQjcDScQasGlSzVhhOaRTKP7rWGPR0q1ddo959QZa7/G7cyi5rjykzeD
pRCSu6wUnM6hyQBLwhN/qXqdprLsU8Toi6SbTyoXU9Xm0uLrggO+3e7calM8qIblXCZrC00Kw4do
OJJV3+3piLH+wSaQaRBGERxaH5VeFWb8vASKj0xOpBELcu6knNnSdqOPLxomdSnvXrH1QQw+BNAa
Z4Adi4Z9EC8POfirT3C3tDYlVxwkCZDDw/DkVBcKQTlEBgJFUozfwaNIW0uIT80Y8EohBVYZl0ud
MyG8m6bT+yU13dP+9xAO06id3kMVuUp1Fpk9MG+kI11MQAK4BycvM8sGcXOWVV0Iun+W2mcv0RvD
horUXy+znAx0Pot5gW1x8XckYDBpXph017vgVzL2wEe9UcCunhrf1oiEBvnRlXalv0Cjk4sFbFKu
6R+B+goQul7J30OL9bCNw4eQsyKOzeueN8LaQDK+Zm3Gvsd3k4YlBBGv84l3a7LtqCOuq5RnuTEI
OQh6IqP9f0xU/l+tVSLGKHvxzkOrh5UqAPrDlFaBUF5ncXow1SRGMf3OLzy/6sXgWb+8tPSoouHV
MzfEEA0mH/S8WinPQTs8rMq9h+CPvLGBJlqe9ypTw5McrAFXePu0wSH9ZTIiRHgXHI2WxORYystr
8Cng1YL8SdeATq5cwyO6ekB/ErGQkiGEsxQRWSB90wAeiuwi9j1+OHXC+K1hRY/nYuas0jvsS9A7
fPOcLF15m0HsuXYxMooPeIwXnJLQZK008XHYa9oGoj8uQhLMgMxNiR6C04mh2iPqxCptBuikJ9MK
WT+o4jfuA1dVuPhHTZyLR4imGYuJ0Z0ejVzC00EK981gvaWt2g00lbByrre42qe+ZBcruKvUg916
jq0+fmhrBqvJTe02/7Pn9xqr/rsfBiJ03pL9EtK2mbFh+IrAKl6COJ/iw8N1+ROEQFJyH7fcsZT1
fdcfCrh0acdciUTluzQjnke8wl7USCxnuzXeVOIjy00iskW21DabN3axqMTpHw5aY4DQ3EUGKwGQ
PD4/AbIGA0K//+0TdQJQuW5PTGcFotXds0RseVpxzt0T2mwopY2jKmIHqV6Rrt1Q+QqOocNvwkRC
brMzs0IvBpQLPG5iHM3nGi0ujqtFbt1gwxCLwAZmV50FX7VoU0vRUqpj+7al73XzWZSE4ReVLX9f
VPe0d4H0wl6CXnbTGrfbyzpRn6sB9a8K+z8gfr0FNczy2rPsFzKHUvOlMtqT8/EBfUxm9JMpJVXk
4JvgprdynLbwmyfj7faQvzHPLxKX+VxecXcvBZ6nyHWxxXxvEol3rrYOVE8UvOsiDs0C7kKV7ZvM
LbPIoDVA1yIx5Qrpj3h83sldRjKYsn9SewnAjZLzuzxfpGS/s4pi6bAz2T0nn6slAwoF+2RPC91I
dWkqCpNZfHWuyvjGMKFGUcw4uurOQRvwl1x0IvP5pABn3BHaryjGa9c5zQJFHK3rTjAydaOPoOHm
eDwhq39xcU2Tg043yPDbbKen2VQvF5CG0ir76ADcbF15QlRLK/BxGwosRobEd0hlqXxgn0yeDYTg
SwYFCtIrBtGDMNFIy264VbeNTva33W3YGJhzsQDB6PnENO30cbBogCp7nH/wt64M7EJkKzxWSmft
5qFgWrUwQkCnV6z6xmoZdK9+oionQcxW1w9mLdNkin5HlmLsW0COvAAEudNEUfSxSd2sOQBkLTOr
kbp5I/fP8U07pbqbh9ryFvwZHNuHu6GKsIilCIyjFQvj8PLWcs8KXyPjB+22MreL/hi/ShExbTMX
ju7FexNlbMz/s6PJgHxCLZfKtDNVKoC0ATS62d2X/NGCMsc+BudG7WGxnAn76nRJ9/iCDHUBTavB
NkGocOeGbHy0u3DUFRgUYtFuz5FpkuP7Bczc9iIWItmHyRBUDpNyU/pUDbRwUPDPVmz7Rhpw9dzu
ibjYIUFQ4+OB5j9eP+6WteT4zAIGqrkaO0AF2e3tySjiSuoIEnQwX9g2sgNOssVZ1JKebOfT6wBG
y3XS/Y1ESlcgpo0+TyW5D4So/C/68nfJQWbGvnndXu/wERtTHg2b/iU0fygaphJv7Sn6gbhmRMqs
McipraLFEWW22UjZqqa42+QPvL3MEz65eZclYk+O3xUkJl4IilS2gnLu0mszt9Wqkx0DaZJNYRAA
3p3TjPVl8ZLk4V+GyLVYZZjU9KOMWbB48fbHQgzi4TRj3dJLsve7EN1H54AHWXfgo7bjCI04FLFh
jAIl7OU7YoGBU74VAUstZjrJrPdmRwYbNOIOz4CB1psBSTSK6NEWxjzyPqqlSQKT8K7lKq90qMEG
qvYpYp6sMxwNhDVp1Jix+W5MmwAKqqriv8YHmYcZxtaEKoJ7Vn4OCzG/VttzgMvwJPBs/jMNX0L3
e/rCqzojm8wAp6XP1kWzIX0O/6OnH2k6DK32dYPuElMypKt2nNPZrCDkXjlwVDuS6iMMUCMcHqp8
UNwF0xQKM90TPC3+gmZB15Qek5o8S37obfEusG3B5ZuzU6Ewz4rFwVXwS51IbbSMqkiP4fugGuNA
XjPgSuPaZCqk9KXlRjaObVNRmDTdAQWyNMYk02IVn1KL6QUI4yhF5nN7/rpJDnE0FlTwy74GM6JU
UsfXKNeEhCRzbpzlijWKY5wgrTV7sQjLUnykFpGotAbaIZobNm2rPosbGOIosFk3lgyFKFrOIFug
VFhIf+WrCF1q5vz+1W/yhemA/CeLrWj3bsrGFaKIdG93yCe5vv3K0mk0fNgVZdUwb9EJtX3VWqA7
Mav6OPNj47gbOQr3Fjbq6eQaav35F0fWG+1/TMJ27V1pH5Fd4TyeqYvkVq90201UyvrWu5VE2rbN
uY2VBfR2ovXUFt3LJeWaNwqppw+IZmpzOj+ZYoA2dzCn0vl2NLly/uzpvzU0J7ljdUQ9aSKgt2AL
8DbMyiq/BPt+QWOrYYhJKk2AzY7Q2M0D8fc4mfRj0SVkYUsZYK2oXR20JsetX7rLc7h3131P+7t+
BkBcO9ZNcdYfzHdg2WU4BPwoNvZXe9cV/jYS6TiBs+NF2stjqav8L4Gx+iBourPOcEtpMB28Wry7
YllwTJ0Bv0HFmi1p80+Vhc7MpGH7LQpenJIhZ/KSOkn1WzbvAn52zpkKFUXEYwrToVSDnyXxisuo
00wDsL0LoOaJ5cvvg+g2YSozlhYmnyFoDXGQikdvhJRxjSKGZX2RviAPCNnsS6J494m414DLs9iK
51oUK1JkSYv0VGX5YAUsMOPEYjnnlLvD+Kt5VP0m7xYQ3baPWSiX4/824ajzppeOQdDlVfvzlaVo
QjTXa65L/OBey7hxDFMLK+btbQb5DcdImKS/switG+/gh88NTX0qu/97+RCxyqc8uruXGG03tlfm
VciRJxtLkPy9XN+ULcwmAci1UZiyGei/nErmjhkyeFxzXL65CZ7KAR2lk9uVZ7UzWyOq3zHOpUgR
ZkTZu7cEtlLIP1zKy3pAmFpoQogfH45uKC8GKDuro3E+RTwSRATtLqo0rClQCeaJCDRom1zxRsQx
ahnxN1sqltabXmIHq7VzqKTz1Do6Iaf/zZNXTDjjNkqnBwr53wT/YXg/HxiT1pJMGBVAFynbePrw
ojYaDL/Zu59NcbhaQOSZ52dfy4sm5tCvI+AyfSNBtJYts1lGtvkfAFUuiHrCvSwAuS8+yExVSCww
dHjwY99njBO4WQNf6jhUAcBRv/OS8EYy2QBqDh+kiSHXvOG6i713/4XyQL71S955Aq8u7vDUjL0J
0Ls6eOnduzHElGuHEUTr+wsOQty2GEgLkjPzgK1kK1L771/iFRC4PiFWMCRKFXehb9Ok0DEH6msC
8AyYz9w3qOru5saSJI2AjdfFF7aTxuC/FrPFX/hPCGTfLdSx9TymLViqzawrMRn86AXhjZuQ+da7
cwI6m6mvahf6B97VG+X0/WG3oqGXo7dMPwfgvGRdygJsrWX7Rzltj3jCjmewuIUxHKUrL9XRGqF7
cjCvBsCZKpofWbDdN02YtesxUZTzbHa4IAPCXz1eQcp2z4Ot6oBurQqsIGqdHmwSzfyI09Pu4lBg
cgEF+31wLLPgmQ7R0YV/k6LrVPzsJku1Qw5XJHOdwzQicAKeR58eEW94d2iPj+jxfeDAuraE9a3G
0loFcLwoSZCsvPhn0si9PUnoUO5iOhAtO0fCDGizTF+Q3QqMFOgQveLjtTg4U4ZeEniaUPaPx8Q/
ACifuIExh0WS0ai3wnGXoL7MGWS3RWLLib/fLxEhq5FOLFLSnsYuuxo6VCxZH42YX0+j6U2nNS9R
JMop6jmuXuTDN4FhntW3Ht18oBGGz/d43oQXFF7YWrbp19GNbCVN8CrIwicJ8M78hZiQ754c5JiU
eR4rBLt6KPwuzO1ThHlH6OwUka7NDv/hWatoW0cfHONHTX2lIlrjtYMfmYEka7NjVH4ScfBdqT3z
gOnlhl+kCQnATqd9h2pUTttM4SeeD8KUpnBYuAgXZjggAFFfLKHpQMUF/N4YoG47dgGM72RjpSPg
Npw5fSLtsETQslCXzYx+Rr9MGgp1uWUUMblI1Yrr4269tkinSBi86xIHy6bdehzQrwzG2Qav5diC
8Bp8NDg9b7mplxphUFmwrNem7E9kjyB8M7jB00X0JU934ig1eu1bPXfqSrmrW0Lo90Z2V86MgIVy
UOR+rvkA0TJRFCyWyQTGCuUQkRy0u5Y2Lx2sHFurc+grQudVUAgViKFcxNK5CI7G/VMI2a3DWhof
lxgFwHcj0h05BR40B+WkGHaTvAlASugZCmXOxi/Y5gM8psCcC9obv74grd7UieALNNDx4L8kEEQd
MmEuXPV+/LiRwG/FqSNUh2KVoRpbWE3e91aTPioLrRv3me9EmHuIU4SRuHb6ZV0C0Kifib+1/uwH
cCQHYYO3EKqQW/JkDd5GvSjyJVI96sLc5o+Z4JvbA1UMr7TfMLA6ymTl2NtdjWXawC4ya2WCYMgj
m4ECD8uMHTrAJ8cGks0DyxZaTXnsMmDvcuIFm8e6lvRXRJqqYbmS8QgLHTeivLQlR297ZCDPAkuL
TeagK5GhXKN43iCqEHuDuW2hGUahDfTtnxcB2aH0Y7t9WWMcOWELC65PG6ud/haOt/Fcek1Y+JBX
ahdvonxT7sHyl15vm3VMg6cFYeFWK8DPhy0COPQd+Z2GkSXL9imDNF23rtAfKwlNN4NcC1PrRxOB
Mhe1wYzX/ITYDTbOJPz8RIWGiMnl7028VvBJqDQlCNPpkzH4a5NMKjoAosFH7Qyc41apeyScSt75
b5Vu4H2FtL8RzGjQRdMl7CaQuX+rC+0dS8rSLgJQf3jgaC26R/m6C2GtglfyLY30aINXgD78Nkcy
R5VfEGNSvQVjqAv5MahlGFm+ANBMNm98hS50YAGI28xkIPpV0BahzEP+1j9CxiOhEXQ8z+0I2tid
YXxVPYNSFebBx6Y0BKDmSfSKty8I3u0Xye3Q0EFP11kKoIy1/oGtC8g5OJxUM3jR7iiUX7xJXT6k
fMlaHwpdOm8+vdYbj9SLOwWchRnUHTlQclibIBlR1mHS0twDEEnykewzM4wWX2QE/eNkefXm8u8c
XOKevi0qXhTRpgGTOZfKVlnzHOEV/ElGPV8yy1VTQlaj5lUkjAqxfnCOR/DwUTpHeQwivu7vV6pD
BP99tJjSvDt+bthCUW8bJsPDjcNTWAnyz3S8eMQ0ZsAcpd5XrG7R2rYcm0CXIH+cfAyYWSvHUEBa
6Zd8iw0VxcR4JrLNC2U2Yb64FYs05cC3G48cXHzYdBla/5FA+4ELuJ1nQEb3d/u+GvIuWu9P3q5m
NMhST/P0Syk9CB+ZqVgAyOokykAAQULgcuHtXJiOFAg7dwL11+nG2FSoCvQGjm1TSencbZfQdolN
sskpVJXNJwoSV9nHJbXfg915CFPB5sKRwn0KCJAQm4LDprJo89gI6K1mx5oGl0ItF31PSd02yEif
EFjtJagp+GBQCrf4x/iAKwYkVEIaykv2FlES5aMgUSxbGf6vVHCslBJfyBwX0/tB/D2Ten2vimcD
9UeaoQJ0tPcA7U02LdxnAkjEUy5EQyI4tlmeZqAExiwSnOlVneQwgKbDkFEWKJ+3mpmcCSJMpb9N
A64lIATdPeuprirTvrdEcNAdzr8beHrv0DoFztTnVxElTLj7a7fEncL2ILQfIKBn/Jp63eKrqD29
PzD4FX2TyxsvSIow6JVt/qOZExIKIVI/9qnZ8EZa7LdD2LG3EC+h712EWfXyCkfg+v7NxQOrtxnE
H483l+otz13Sf22uytrgZohLcMgGVxeUtQ4zIqS2e7lWls9Nu4SFU6esWHJpCRmjYlpiHSpwpQYR
4LvKpWqkdvoiJ443Q6cgFw==
`protect end_protected
