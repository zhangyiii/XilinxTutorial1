`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
l9rLb8eyF3AgALThasPiNG8/4BBm1wwJaB24bneaCtyp/I0xi7SHB/t0Ctv1xqonweX1MzV/pVKs
tQdRNspPIw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X5KWlL148JabgR5weT9wBUkHFWddJA7h4OZFLd8bdBf8Kop7kg1WdkOhUDgmpNTHeXS4I+xH4Y4Q
HjFAExnYrGUC1wm7p5WVL3DFzD5WTILYoEImzLFNcK9/mSAIwCGj+Wtr+9xrMpQDaly5jC8Sj+rc
Nr34z/YYnZpZdFjSjFA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XOX+x3GXJVQTrGGT75+NpApkQTW6W42cmWaYkzqsNsDYv4er+FitAoIemlb3od3AsSf9WRWhCQnT
6iXQilkemT2DzV4Xsw5A/7I/FZ1E441abMpjv/w5Z3kwpJvNtJvcGvjcX812mAAPcXsPvrB5LXuC
3JiNsCaNzfl0IQulHvHCqzDHmgFxZRkHPXNoL3EbdAxxa3qQNIHMXziT6TfG6V4ioLwZkfmj+nFw
X+PAA+oZbdjyO4IF/qvCl2mnZ/REv5vdMZsnEZ7xmZVfOO9rMWwJcGnuuXesJxcZqnyEOewdy0X4
g5x7ACzMTBvW4JyAsNl6ipSaUUNJcxvmP1Z95w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
umhSCUCmm4WZMMJVCjLiDlzFgH/9KhaxQqdvYM2gFaFK/BSZmXwKtVD0oGzsfgEnaEnfAZpnMH9p
W4FaTz2HfMA8FyEQD6bKpLwcrFDP6FLYTus4W9auRkdWk6MByslYcfESnbPd9BplDCjnq5X9FeJm
J+EfUISXG1WULY3BqQc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NcJ7q/waCn8/m5wYTzYlcTzCH0J7XhsrCXDcbP801wBgwPzwk6W1YaeEGpz6w5sg9/BVkYMZPdHy
s116tGvxEU4yIAoLSq1V4khC1G0CICk3cYOL6Am8EnS97sHVRnu2owQQ8/o01YRhaorvw4ApXGQo
FWXh1RTAkyoxms7xpWs910xGCq+5ztWRsH4I8eissSMkhuy7owGmA0f/OPnBvz/16ynnHSqeTcgH
5zrPaJOgTZH9aMea2bstTOpguVDKDnDoAXUHV93yikhxVZbDx6GaPXUh5fshHVEaMG3kP839Gx+j
prw3SfsWydM2YztaOjt4rwHOeUOZ19sYd2Gsaw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4944)
`protect data_block
GMQYRLdIBu3cBPESIImpy/E5KG52tElpRDp8X7vzNtDA3AK57qF0gJYr8K8ckEqqOqGzGbcmYpy8
TOOsLR/OmOuuy+ynRB2tioxFaomvNhI7IGjwAZUEF+aPkfibPW5iwagbVZ5pPArrjpOks5lOMRwm
bSB3oX6QnyKgHSehE2jRDTJV9qzGOfvw7TjiBoGfdVLSH+RbDlYT37n4nYysE+9NufZVFQOxq4sm
nEexuoy01fngvMCi3y2NdV8ttq2WXVfvFsY+T/V8yd4smbUiLdXgoe5s7LKSQwZo6IzWYjyq1Jxb
NDcEw1+Yu3daFYS06SZeVKP2rKTgd7b/ooX71Dg+2gSvXUOB88pjtighJSipVOwrRUrelft3mUV2
/m6ZthIrunQ+VjL3DHMOJ/y3K4A/nVgmh4mrn+Zd5G7hIaL+G9LUAGZNobzPch0Rmw47Y4+OSHCJ
c1h8uOFt9rkxe6YUac36hxaQ1SYRIWAdBg5717UVFynf7M0r7DDzhxcnhh3z3g5kxrRejmXM7yz+
nEWTMLHcgBcSrHVN1PUzpUxEcYkG2z6M3jW+CFqjuBRGYQSgeCY5jBjgvQf/D2RC9G0Amp0GxA0r
yJmlycGKS3dWOWhpvlb1RehnGyNbwUoiSHd8s5uuVGpQSCdwk/9Ux6uHm2Yr22mQaDQ2PHsur8og
tfryMA3S7T5Ak7saSp0tOr2Rs5fn7FvLOC4WN9BBiVhA11wy5XB/y50WpKZEYBgRT6GReCh+AjlC
5Fh6ozBWfP9B+2Ct35vvJQq1ybqHAgDND6cw6VthmbLfA1zvrISC3Hgqs3ay6RFBUcwNqm8IiXxu
hUDlyaOXnlQoa0rVxzmwh2pRNF6N/Kloo3KkxU6v34fsqLNKUxDdMsKNyk2xKD3AM3KJ5OKuSoqH
VzeYqZ/KUanVLXni9g/oSmlyOMejfe+pRLs9EmLuCxY9YULJyzIhTAwrMtT6zsW9Y5vz/sTNzePj
67rdDUclnZQeDK1+ZDiepLXqlUqchzpihDEwcax9XlpppZQK8RVUrMwZfG0YU7lqGcQRuLrLwep/
w8fOOs3tQWjDQOBJnWJ702+k1gM9FXT4IzoUplwjgUJTvz4gYocJ/n2XwM1wfSd5kR1NvkQDEXqP
Z7S2s1BkpyK/c/W9Hxd6RGtoTDvKaGI6G5XfvTJvRHLJiBHmFKlENZnJOh+tDNy1rP7LeiuiNYZH
8Q0kkR9UKJmSeZsRE2xDYmL0LJXl1p2DMeIA+ocKf2gq3H9GXPNiMzLqMR8T7x/DdhXzDhKU6U/y
lhDcUSQWZrVq0ZB7w72kYE3ebBJssLvLwG/2tI8Aoy/wpmJUDmBSHAhw8CYQ62ZPPv3TrVenatyT
GuQZV0yKwfq4nU/THEVLEeHLTkS/RtE0Q+mme29hBy54GLkJvyK1dshu4XdrBmXSOwrEBrS/MVp1
AZph22VktXgHmXFMERjzGmCc1VmXLYiltoexVe/9H0c3balGjT/zmNJ9bRB8XOQwVCpLTLSuHo/v
HqdV9NchiZEt74GfrqW5n3IxMljbDvt4RWYwbDdyd2qherYk56uyiI2zONcfMy6yRbBFs6AWoXzq
eEe5BxI2+Ti1j2ukLsQOAk2JMV05lGLaFg7I+AuHBZ3Xfmkq7I3X/CWnVpiOQmoSwe1vluvhjpNk
oRXsrvWdmNXCiRpR2Mju6EQ7qlsKL6mTSLhkm3boTG1G/TGOIXQQ4UpbxPdGeBthV4FOL156yL/z
+P1s1xfmiLcCj74fRkO26Dw0Czq7axlOxIZN8W6Q9Dt2jGBe5clfw/stU47A9OCexC1BQKLAAlST
e/CTxT9sx0YGJjP7n6L9N69SfH+wcizyJfj4SCHeoYAlcVeOivbmi6xGk8yjMU7LMxSNIkmS7ezp
XoQVjGV4BQMoGWugYwgjS2MsPvPaqDvPyJZY0hLNhHavBXV/tdhjfoRds77gqi+VZiUx8BzJ+P6R
McZGfwKoWUfwFaeHp6lmcFW5atCayD0mpKvGPX8SCEAH9HtxaEn1Gz/QXln5PMJ757XSOURMYRi+
qm8ahrCNUHsr3xycfuj6LZe3DvzpEluMonszRQv1rex/bGYK8E/53fzLizWVR+Z64zS9ec8MjMxi
nhbgEe4fgLhv5nG7ymjySOKViS/Dew5F8vZK6QalcepwdAp/3KhdwUJVDSQ7VED9ls+943maEaCF
ZPk7Ep/DoZ9O3NN52ZC8XRJBJciZUjBkqjKmBfpexG92DIoaVBgwuam+qXn/7qdap46acvx2T2wg
ruazuibBcfLL5dPCHj5zgGJg8alpiKtGL+TbwB6iakKBCDLv2kDY4Dic4gAp+urrTZENvRMaJIrl
ia9PSkRnZ01YJQCJ7XmKYjYyddIB9aCUPHRwq2+bPS1Vq4HNYrpkFzk7eHhzYDBbGC/bJOkZjUbn
ITsdAILF2RHO2wh9rIrwYKapju4Fw5xoiCJYJI+yU+W7VRin4TdfPz2bc9pqhTiGRS0hUJGpWYLz
xqxFP9nrWXEoKHCsv+a+wsd2dZ1L+VrDlugQq13jzWiv/+MGpuc5EEpPaW1uJP2bgG5vijYKbhh9
i79eyHIQUlzdxLRREgTNdNCRJeSH0LFyvutoZafLqGjRwnLaO2pKk6o+kauPSTx4JJOi4s9XhxCv
vbEfLGsjBBIpRESnQ9Hixkv05i0mkVOvRMXIhGq4dukuPtxMYu7y58F4FdJumrZIhqwUSMupEMY/
Lwg7dK+SmPk0pAwrILnYdiG3dDTTslEttOxHGWKZJjRjYHeL/FSeyABm2znEhhs+dPDUTqvBYTaF
7u4NWux3G9dCMZlpp+Txf1pumBHHXuAz42lerxAknN1qQnk6Ui74IytAnxD1532pJOYtwf+n14hk
aejd/ra8pExkg2hmTKlg8P/MxxTvuI9p0dsWJjbbSKIgGOZxoeXhQvpqJphk7WWXBRwQg1rIvb/c
PCYJlPszezX5nM5s2DVmq6c7u+8t53NR1aCZ+wSfXWedlx3jVroRtPb7AOcGs91utdBB4QGBFwZ0
CegDJzK3LOylS+sjy+rkcnMA2Ux+SxaWLBihYrXl7mYSwLOcL91zge6DfTM/aQ/ezz9nW1MtNXrU
hcqNNT9MyFI4fwJwNCdcBj/GpvKKUCm4nuQm479StrxtJCQeRXQynxRCBVCa/f9RgDcA7Ea3c8EJ
HdTPtrvwSF5YPKtK8pgl+lI3niDVEX+rjJCibUNPfzLr2ic5p6B/T6viIovqfAn8ECaHs1eEGPIf
Cx3Rn/CgO1OieCCSF+xKnXeYUR1dbNAAvqI7ZaBkhUwbQa0hAE5ljRnkbw6jwkd1fe+Eo3mdkqWY
6clhzOsFeUDzzGkEzwNpjRnFg+iu23aW8xHvauKYv8nrlKcsWOtntuZzu4/kiJUTPMIB2wzrwH/3
7gZpPCZiC3sucq4pt9hwJxyXxZ+MeUCS+uzH5BgUHaIm8cuXtmGgcSz3OibcaLQgDrxqc4Lv5NUS
XITdyNPL+udLkP7lPlleWrLLOu7lr13I2vvPo3Q1UdEsqdKzkPacwbYlPPO7OU43xj4QisK2xr/G
EWLUQQ08KcR6wCfo6frL9ek3xMm+GvonmI8x+iwKK4k5oimDHLx+Os75GxjVUgzc95xgpJ3vTmTr
t0aw3mXxcJs5OEkBHRPTCKORZG+6jBxieMG5CwdVk0rYdIJZ5xa5EK9cWOfzuIzLQRPNLRznly8J
/yJ5UhRDEX2tsoaDBJRbrPDTKDGj5cDOF17LiWuE/Khq0iCo4/01zXoTZB5FGTEzi0u3iVvBNct8
istjI2WzTG4eVqc2yqglXZf0+dL6CiNIgsZzCj9Pa1WGqzZtiNb/0Dbnb1xknuCXIlIMBpnl1vz8
/tYu9XpMUIBcK8SMlexjtpHRzTBKG5gWrSZZ2kgnUVhjle+lPfLd7P3onYcrmTe2OeXFBVjrkDOi
1a0X+Bv+JhUkqzDBVsQ3f7Sw2lEsoebNOOEfmoELWQTqM6NAeQBbKM9foN/hWEJlHNwZUSWU2dLY
CJwhRrDwTThiaPdA5X+huM9dRjseT9gAeh9KFh7vFoXAz+9i26dsTr0s2yKhA1oO4kmdPnAbpjtr
2+yv/Iw3K/eD+l/U/nkdpgK49vb8xmiD8hXIy1AEXkuJ0KRPFlZ4GY2Us/iXGRx+hBmnNP3/b+Zr
NvFYtlBDsiOSpHrhpihVlf8wr/scWuDbWBhkmR2i/UeiofR4G9zw1REyjZXPESGyNmMLvFw2pNRi
l4X/MZtm0MK7qzEoMHsrSJ8Bw5pEa4+QGDQUmUKG0Ea6R7bJJHq9CqgoELDkqt+2zCL2mDkRUhFo
EmTxvva3yS1WBeN3isBbYBGrozeErS8aMuTmLPzclAN56wLB5GRDgD0mEQXEgldwnuKxOR7Ow5dd
HATHsWDXDJA/qvtmrV+3Y8u7B5NicV8sYijlnebyWdj3+FW0F59qvTLruS4za7kKcnH/8M+7UE89
SjY3201LNa1nHmbhKgPNpcxR+LqKISiR6ytrSIkvXPJVwK4wgxy8VV4XoCMKgMZStagnpX5k3qY8
hpwefeRBD5sh65rBeAGPW4bdWcSdWZFdYPEuCubH/Ua9YoEbd5Dhsq8haa/yBaoEGQczxA3tU/8W
rz2slSWptrNQABBDjfvEb/gYPQEpx9eBHvMKcIqjMTNk4QvB6Y5+1Z2sVNoWR9NhUZpw8eMlvc4F
/1SnWGdqlrmRSi9UWz14rC9g+pvLwIosCBZudzqIm9HDZbKLNl4qPAqrGp0Ss2pmvUF9hJFo+lpr
QGk9a2X2MHehPlc2037iX8YCT2pyuay3Ytqj/rxzTmQQxXYTKdJSJP6tvOGc5KhnLyAyB1xTwWbz
uBcI5b6lBTUbkEZJmyqzGFYmzaxV8ag3yBR0BU/SzIJ+zQbsaUrx6pLwNRw4F34H+kxnBOldoKub
x8rl3oYn/88PVMpJYtDqVJKm1R2Kc22AehJVw50unY5HVLRoYxHtWhLvhIhxG11ZdOChcuJNcNaJ
78o+6+JqmaHXOkUqkI5D0vfweKMJpTlqpTkGecAkW8+uH2nzvWn9EbFXMODncR9EnEToHqTCb2Vt
KQ/SeHnCu/68OsLJoZ8+MQGPyst4eJycbEXhSZtzdw7Af2YOriJek5NG3xKH8ZxP6W3gZoWl0qUM
nEeflSbHYfs6cjb3E4smxhAw+hoUONYgXTKGayk28Np8dg+DS0CxkvTho52nNv3TJUM9Y3dZHKGL
16naacwpF9Y6raVDbaZrFh/EMOqsVx8dSbjbAEfmCjGZnEH3CGASFjhAC4lRXXfpYgi5Uj/949ep
QIEoLBjILQZAXDnjXdL6ZooM0V47jUu5czq1jKPuNDvTT8aDIwI3iV7LjsrHIZfgaE1BPZiiUtTB
7n2GhDUgu2REcUk9qHCD+E0jgox/tKZTNLI9AKarZtxjWFXeYpJ23xz9DKWJ9fW21e9dTtSUbXaD
NdY2lXSNXO4S1GC+fPSQE0nmlhv8IMa3YaOtrCaZyib58W9kRMAyugN2JsAJPDVxDNib5/e00fvh
bT9KgEhzc3fD+jsV2Y/N8GShhe0sjhWWyIzAgOocUJVNy1yUI4hfco5Idw0aDHhL7Dqpyjo4uWQK
bwBQ6dcpLoMidwaBJrc4nOgzm8yhIATuh9UghYJI6NoWttsGgE3RjVU9BPur7QMqS+wQAapRDDK7
TO317Vqu8wfWMIaHw0W3U9+zUWYxbuoIRWD0Jlh1ToU2f3FPGjkGqToiwHKylvjXh19nYWhVFBKe
E9Rqy32MvrP3Bm8EieXjKoFn7LBbgZd0t8oyPn5n+EqDVrPW5nk5pBYjMHjE9FoxQ4Ms6Cp70pTW
BX9sFt0nAgY6/Poqm0bFoM+8l+48o6It+CFmGvjWyquWExGNccat0wuDy2ERsbOtlcWt9e/ecTq6
lV+ztzcBPCaFug3YNpeo78hqBe5zeKB8Kmwlm0MgpQmTRip02JcbQMCc3bwzQojCa8tjIWIloOaO
gySYhjIYZnknWC8ALmAStJFOP/olRUJHWI8epkHyHXYA+7fC1zcBydUlu85PaWR5wxnCg5MDGfB0
w9j6W80GDE4MfzD3ecrfv+MZI4yr6jB1uoi6Mrm1BokNs7bhswjxYm6x3S10hmZqALotnaGxgVPI
OU76SGHQ+/dEYxrolxM9wOU4vb5JXHn5lUyDooxIyastLDE5mdIDCi7/IPAOvE5lPP0n7XiTQ1HT
I9O+lSfrQTKdX6PX3FfpM2Rckkv/QjPH/Dtn2LE63DdFdQLmsPiIUHf8pUsbRd4G9RdO99ePPKdn
qgxxs9EGtIRuWKulbFbNvU5LjOg/TFT6DY0/FrfXT43jM6/wRzdIjDrF8hIVjXsylA53slT/N0d2
ZjUBxtk27H2pTszadTDUp2nZWYVuctwQ7zBxXVGtrH0lVFJWTiUmB3+xBScY4w1nB2uxOnTfJbMY
wTjpQYCRorcHxnbR0rOKLrqts7SYRebn05nOUklaKvZrvfsszmDSSYOqrwum/KTBAvBYxOsPwV9K
4vhW6dQFbh80RJbUS34lkz/F2ibtHkQD3vU4wcrJRjDoy1yog22L08Cs
`protect end_protected
