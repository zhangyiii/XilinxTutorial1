`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14368)
`protect data_block
wrovcHZ5qwQL2M/nAAAAADeCTRrTnvnNgJT+JPGsdI4nsAyG7n1TzmeUsYWeQNNUs0Cc3gcKgNV/
KPhTo6rwSM/jRKiQrhDAytWjs7xX+K4+YlRtqwMUiTg2arQiSxlnRB5xGnt475/+y0N10gAJ6Atz
J8qDnJkTpYJeKmF12RYyKSSIEIuDYrDlgk5BDr3gPcSh8RfUrxfmYPXibaj1bXkVKVsyj8mwsl0X
59QIQALLPd4xRw3eD8DxeQRHIJKZLS3IoX3PsAoxMGV69gsTrrB8vvsQC2e7zgyAFXEzyYIzCF4o
tB+azSG/5D2UcTYBJLcWHS6mMbLhKmuvIwSkpbioQ1AvxzFRCYB3SQbRmr/z0sG97yRZfCXZWMqk
aUV+Paw3aBMBc8cVDLGv0BeUJsSN4M+THBB1bQjPAS25vJQOpl4vnqw6CpuBPYSwAQBFck78pOkm
h8LiW5tOLydO1Sz2ROFeerhFg1k8Ta5RCGokXSo3VHRfc5aNDDDECcAu49NN1ijPVq9zuP962gXy
SUjP++I+gywLYwd1AVBGXJoG70w2MX7LCsUJ/S9ea1dDfJzaVdIxVSJC0YOtEIS864AASy1jf9mb
64apbAbuFXHPe1ogf/5vU93vHJnkRfuQQET/W+oDIGK7UU4t+pBWTOM8Cbg1cphBnQqckCYCFOIr
0etz2lA7l4mAC2wD4LxHFpumMLG863XumtPox8gnPWJNAn5XLMpuJ3nC7PyzrcE2HRBxX9ugU5/w
3UQilEscHIkKSAr8ozQTXbGhofYFdFZLKujpI6VUEGpGKYDld9HccSDYc9QTOynsKRRsSdJGg/Ot
v7c/pJC+p6vm8vioW4OZmMs8xrkheIMTZV3LD3Py2KFYu/kHT37BKtJ2c5Vi3pe6oGm4mfonsqtT
l9JI4+GEOkn4zkLocjlpUguWc66NmcSzJVV5czmNp5My0hL6zF1Grk8h/Vq+y925h39XZSiGfeX0
zr/ae+KiOS+OE6J5j6y3ZU/2yTskYD+BzqqB/8GrE3gi+EZV+AHea/0GVjatl87yNpqlzjpDndYT
dPv7RtHW2X3Z/bT2gJIx0ivzyrQWeKMoIOK4ZPCcL0r9oEHw3+iCtplrAi1g7ZjVlXti0YxnrgMF
xEM9GsE9pGpVVpg9L2FD+taeSs++6GM/a6pnnYTB58VY8DqKTLXWj3qa7MtsX+HQ96VSy85mtaa1
Sbl2UJ9OV6qHRuoHU5oYNMeK2StACjVKKk4fJmTOjagjMHyTF7XWpdfdH0kkwWTmZk9rjjZeL6fn
46PEkvoipWUZRVMM4lrlavjASqFMgsDrtmqQImM5bghFbtqvTN6u44CrWDDMSXKJi0RnkEoKF61L
MN5Anw1a7jkR4DlzuKK1BjjT79y9a4UT/eyjlCWGB0kITVFmx+lpTbzR4c7soHDJwPulnWyA65Km
v/RYwgl/wT53QwEJtGtan6HcDAGdyXpZABiorXcATmjYliXVuN2njkPXtma4XhYkGMGJwCYVmye2
8v+dhrtEbyuCPrRzzqDpfajMhLqa8+CGEz+BVG5uQpfTIcMSCeLCiM/uxzKV5GpLrckghg8E2b9E
0zTqc8BK2S7eLulZrdqsTGGAI2DFogyZb/VDAhK8gadC0c7NJIf2Ruz/aPPYZU1+pRa9Ei9K1QMy
suvDZvwrFPsghs1lvNU2w7v5RxoB9Bu5li8P5Q9m0676lGBFpX8U24D7JYkvc0eT0jw/h3XZ0jA7
eHj3th+fqEijp5YKhefatoZb6G6w/9ZCog1iwnc8FI44wQNgllzkEck3sPjlblaFkucVC8LBemKr
rNVnOTce+KFREiqE09o45xll+0+b35pFCP60eMMKHfJpX6wJorkS59QokGiCc48rdqjUqqXwPLwx
KH7VNyhgCY2/NB9eUvZ3EsGsvLMGY2eQF/T72D15rGsAhl83uory3zk3wToyrHtaaPmAeUQm7LQI
RW+lpmOddF27w3utNAnGo8G67Yq+OKgXnpcdz2JjOwLGWOAO+PxkIjUWuuLYZiKYO6kOFFfYciqc
dvefCvlptQeITgRKV+b5L4+z8WZlhq/nTJLMOd8Zf4aabhbrrJYF9WCvo2mtwcnuc0/Wils/bYIo
WhrFoSyx1dr06EWz6U06WE1fp3qjR43AhKkrX28JCPWeBj/c1lHqKGsf/mptFI2rkuijShfw84pt
P56nvpAoyNi+g/hTsJcd0HLkuD0baOKgfOOTP8qYs6UZly5q+WJmb8tmvlYij+Q5RRqpkV5iz3DU
pvy10QUw+spYebsJi1umgxofZqCZVKIcW4A2gKSQBnISX61d7rAApJ3qbeaYhasB1r8N1zTitE9R
TsL13Qhp5LfTlWN0/TdzYhHuRVEepOu5WJEDySm3oknym88HoOPf6aAaE0VnhxnbYhmmWvwDrrV5
0mPhbKWSQrNmUQWoHY3IhbtYTA9Vd5UL2i/amSiFIb07WP8D8yuCuQs4gGMWf4ycGnlwsuFaiaVW
1oHgFOvqAX2sSyGzn4HWrFBAhYAIwBzgz7Gu3hVF+XX+Y+By03et7BM9D3LLZLlrjC+/MqzS/oBk
QQycBclfKrVWe9LoxL0pBf92BezL++ohq36Ppo2t4soekJvtgyI8sA93lZvyiWGrvjDRtVbndDXd
9RLl7ESUNuzeLecwbS0L+/VKqejGeOTjOgiv4JL5pmBu7pjJ3lZQLdoIwVvSvX8V7nvTZ/SE9z/Z
jf/4jYhlf5rLuvIl5WvGr5BQ/uCzCtqh2f4s1kkgKs2BCu1uSE90wEUPhDiq3Uy7meOtFwe8Qfee
y6ELhy1CE/+CIUM3mfGy/D4b89Pe/dERR/NmUUp5LfBEthpzqKxXK3xBb3hHhNL6D/jpQLaOLZZ+
XgtXnpDH0FovrdrKS/w9O3T6mvEzZ3wHTJ6nm+5RK5gvFzEklK3bGHy11gkztE5viybKPiC17Ljm
VX9cJsxJOfSK/eBSDU/DJjh8C0/1qer75R6Yl8Ocv1bpj6DCxVf3ETlc2VEoRZm75Q1FmgX13hSY
cwxGZ7njewoMBF/unewTYGMlqAXjVTWyVM4Hlr9n1xNQHXyMd819dYG1hhuxVaVnaPvXgCzQcYG0
nHCR00J93JfWQjrHMXpdmTxuhLbH4Ge+WoIN3LXqmOngobZDcWdx2aBufWPQC9W7trK4xORy5PBO
8vBEHmdV7+ZZUc62I1q7B67JeD1yPQRU0CfhqcA8nYiGS4FpmAR0NKFC5XtHgzTfL/PLcF0Hr8af
A5eMEVVUgKtQto1XJCkvDEWBtUAyFf5G3W1vjxmgvv7IorfHFx9FBMFY6/RPjDV7yMp9f3URGFvR
2AUM68QfkqTNz2np/Ygfu9QsOjgdScbmSYObX3faTraqwhqwz02FRF1FeHW9wk7V7Cfj/h+8iY5E
uwHVNSBsRQhAkWokvGRkC1JKahFVqyPKcZ6ANdC3BsQuJ1L15JOqVgZY4xqEfpK3Q+x+24H483eL
/Dizk8yCRwUrypfEZf5Ps//ldmVeNd3AXncp9emzVf+JlQgKY1dv7haTfDOOvcgCZI2EKm+XoW6m
Z6jwYFjMcyq1r1quxn4SLkU3aom55/zkWrs1b+kuQ7WEVK8SLAyM+E4EcWhA4ia8hsTozi3z7Psx
Ab4dKA1AD2c8/+AHC+Kqv7PPUjVK8rOKrU9HzmYc6soxdJqnyG9LJPnswqvAqId3PehbhuUiTrLL
h0SJatV20l9XQlZUP3o2w9+uXHnXRu4JyWRmO04EJPFx3ob261A/vFjE3a4IB7Vl4y7IA928qJeN
UZcRJ7RFGEgJf5kaJXNxFyY1kR6h4GQzGjNQ0k6vjgJs6KieAhIqlV77MgY5jRxEMxmYFMctTl10
8wiiwY5uP5mzRoBrfTldrJQOGta3zF7n4Il5vbx1hWXstdlk/MGZn4HCc/USdiu0tYefSIycmHNx
gh7yAL+lsx/DJdPFa4Yn47bWoz5tyJZR4IbQHpFwU91D2WcupByNpGUXlBbUzHxvufMxcJBmXd3g
Im9NEQF2mTmuLWlqZ6DbeWyT9ie05Rgu6IeF+QhyFBr3rRkLnUzKmchi04O8HRhTxjTb4JLhzTBi
V4KtXhpOIgFVJM8lQUVKoxgjTpcXhqXZFh+GYtD9r4DFtaK6Ezj4gNvW3LXpiB8pl0nqyZOYmfUA
yaUWI2wvyC54BzP97gfR1rHozHdO21doAT/g445r4cbSONs4pbGl2XypnVdN7p0Vpf1WPN8Eb4Zk
SE7CAs92XiRdd0jVn88NMOaDBRKdVLoxuagHkbbam0gNObmYahERxEx8QCvvKHBR9/lX7lHqoz9q
bhu+R6waBVtAgK/4dFSQxWqkyB71Vdl1JAA9fi+/FETO28juecSSh53LilqCeqZ3T+STkNb8765C
yjMerIbzMrNN8OPd3svmIwu4csooTogMHFpYHhcFYsyQTSdV/hlEJmq7QGhCjOZFATYujB7h9EbB
FMQbhibLtJACgtDScK+JTnjJMzd5oXqXSAyqoWHpPuaN4ztRR1SIRPO5Boqf9qpYisBUYkobXt+/
18NK9oV5Jc+xyg4TZavnDX7VVuOzJyl3SshIS7kecSEoXK2dghA+9NaOJIG/frT6m60z1a03tiuP
IGaOKTnuVeopeVO8Vj1S4JjXe9GHjoap8hns/FL2InVhRdzIa8nh4ySwvx8mT+1HGyc83Vx5ibit
J3WTcq1nV98NaSC/Ievi6HS3HcSs7lrXCZslxPDqaVR/t1Oxr7ynZCZpnIl9JP/UmciNQx4pkiNy
wSwr5nqo7jMqhMpCHLYVivTeDZnABKFPs+ggXcmDaKpTUL0RNPViuwUFX9xAd98Rk9eMqu9S1R7d
cKD58FdXGq4NA9iH0kOZEGSqCnVB4D0ZcJ9xkyobL6ByRR/laO5vlWdLvcKHXxQ9Iv3cPrKyndR/
mZMQU8hVFwdIutQeBCaUQO/4MvyBOOJLuGjLQLQnTgIDhSKMX8rKJfLgQdrROXdaip+BWPsLJmFw
+qqN8z2SbiWcgp0vzrDbAFEGbfldSFITxx+k0QILtO+hFJ5Vgj74N5i+DW3UZn0JWITGQTkv14hI
Jp+kF5dpRUlBlzvplgD3HRIwAeJojTFKsa77pHmuhA8cT8x6yXCKf5Rh+khsLPIKKuQsKNunjEmy
4D9TdxFPVHpSuFxd+FxJLucdJCBmPLcw5pHQXFSeKI2y5tKj/vVQ8KWFl5/02RtSTP8BO355wbJP
edjmaEEBWvOSMylnc8hebVHFNh3hHX2X70mJwMn2qvMsdn0DM9SPhKk7wdRD67Wzb90mw3E+yN5R
k60aroty09wH9Rfq41cTLtzadBVitZprBlpuIMnP5nOcCdEKpPUzT9J1Cq/JBz7Q4TdudFN/4Ltf
DTlpbju5XihfSkMmu24yNTzg8QpXC70t3OQLleDkQOHYWyevrk/hte7aY97m/Z5PllCuA+aowdn6
AkymQeoI/QizH1cxrUwBNaUNCcwAPRbm+vfiw1HFgbP7Ukbmh2Jrze0pRykOlKxar8Pu1oXozZpK
F5/WuDrhhUAzKTiJYZkMXmpKwQj2AE+C14OFbauHL7wVteYHcLe54sJHgitTdRdQVzWvIXnuxq3w
JcHZXmn0vZmm/2ZYzuczkwrrQYh8SUaf9GrTP7nOergg2cPGZC3mbm3YbIhgDjdlbiaNKFvXWxeu
9sw7DMbqZp5NyNZA95j+H6XigSYhDeBSueU1dC2QXmGvXkfK3/yAE1k9qFgm9XzNC90EtMK/hYFM
Y19N6EhCIlyFLGXXkOnn9s4se4SBHID61oA6dCPpXalHHYUdt+UfO8Fk3k5EH3yyttHGIky224vX
SRD2CJ1El29QBAhBgAWX3rG9CWKpgmNqO/VpEhUi9A0W+BJE14pe7VsmW21UY+MsC+04YUAgOohj
4PtDhdMzwnbFZAcWWLm3u+D//JnrlwEYJvff2YEJFNfWVlSHYoGrCG9z+/9LU6ySqyAKzDGU1sql
B/W6t/SGMTSVU0JoMl0RJO1FvzdBsi44foEBgiyddp2y+/kQ3qRyons5CAFurpa74opMUtzzPyKJ
Bw1vfnL9fT54XRneiCBRGLCijSFFK/jvKIMUyXWq4cv2NWtksEOiXSOMxMEGTPD9ZHudKTYI2tUE
1X1mEkNgf5I2R0F5ckuARryTdXup29QFbQ+ZtJhzsoGfuZiw5btHoS8B1ayjMEyuz9+bkFN3eYtX
rqqDn6c3YoCwUv/+DcpB8TIlEpAJCIO2MZHoR0uwWUOMvayA3RxLGwn0HIRg1U6bXn2F7CCeN3Lt
lXwJH/I2POAITePZ+9jlYRUv613T66gM8bPehzxvl2xJay1WgQ7+pHUwNEB2cNyHiCyfLU5FUT46
knBimtfp1b/sHi/84UwGWhgi7OrtXGHmqPRG1UxrTAifiRS2GELoD5GJzSc12TNSVOmcV6OgpNGr
GO5rwwJYwi4JAJPUbPVF+s4SagW8FeiggCOG0O4vTfloEqozKnHeCpnZOf32+63m6ABOT4vpJg+8
EVvxx82/r51lr4RtXZzk/Dk8IdJn6TWnwNAix8YzkqPhhxPQO60aJCrenpdE3rOPt3fvlH9KeBBV
HaS3gVRUYZ9Wk7oh/PJ21MphJKSWyt968pLV7Wvan8tezPgsnwTZ0ti5jZacWFVvq6VIWtJr2bu7
tx+3tFmWHCTPswMQLiEprwHq30jjrts9BzhQTQmiQeeqqAm8/88kuR5XbnTkDnamkQpqEFSrRYLy
Nj77h3GvPyyQN9MRJlLgOiuC4ze2poU9np9w6Xg7PExzf+k6X/P75cfbE31rcQFPthOExZsguqly
g0ObatO/jhZK0yVyxPe3MxABKgd9C9b6clFo+/VhLXDPyD/s+zQ3ay94GPc58hs2uqRpC+yFDKc6
M+bKTAS08rWqe4d2F+Cg6lSAWBaOzNkdO1VU4OjQ6VV2wOOXcAUInJfW1uD+J70CM8C4HsCxVV32
f5qO7ahN2vBTEh78MO0CcPA8Pr+eRuKO6ZG8OBxnx5aaecUABQEl7YTeQ6KmA6MxnbwC2ybBbm5d
J4Wg+jUVQiZWH8R1ziTFnN9Q247s15xDEEfJm9oVwibnoNuZ2zxxIYeB3HOhGpYkBUSna/XVWn+g
ZbdEKzGa1nSzsWF/gyhyAaC2rs+//KlQXJpOd73sub64LxMnNlDyvQ3wGlScnYbPT1VpPF0AID+q
RxvUE8cxKnZqwa+fZZWw/qsMNkrkVJXEA+uQTsbPcnlkBbJJv/vE23IXpPZEK3BjH7dgqcMehtGE
ewxiDr9irbA1y4leJGbTgbZwTVTSqNFa/slh8dauhZaMj7Vu60tNhOwNMaDf1M3Ix7LuoO1Y54nG
6r+F1gwbhrdkIu3xwGC8yEqzeEl+c4RlrT9Y2d8M1MHa+N6n2VDbs5bfHEfwYPvz9lXfJdaHZtPB
H+z1NxOu+n9qKv1qbEnYigHKHvAN26U6bmMp+dwY3A/B6Tj7AO1S38oE21qNoh+NMuEDtQ8cpvhg
uA8hS9e7ULOBBIjO4GjRWk2R4JImD7MaqeYa0UAkRnBtN1rPxv4UmqUda0BJPb0Fivw+CBMRnXHZ
8mx5ARIjJa/5bvzNBwS9ARp+BAr7io90K0yN2OE+vDCHUpzRPGxbMGaB0nKMpNEcANfZ36DAmuLL
o8kuwJ2XgyEvzV5fsdWH4uBo719NlDeprIzPRn+B46Ka5NlQu9hqq48vu/qz2rWy1DA/ZPuja+s9
FyviuGRyb14fdlVq3DbkQeHNW564TC+6qgKtu0klckBDN5FleCkB8iYt8r9TGENrpfchT97U7LgG
8pvnrudTxXoh1rni0rcIUoVUOEaCCy0z/WxNEHQL5UhS84LeycRLyEG06w8RHzBV7rfHhYIWMxPZ
6H0nczjMkiw0nhMVECXm3rplOvHgEfOG1QylVVUlExsfWAzLZUfoiBFSKnvlucYtqFEG9MSoRBM9
tkdLjHzj99i4C5S+s1oSg7Z6hKMlrFAPaH1qlTcO2vslk3655tjH9SWXsbtjqaP0dTDT0pNfAGvC
jIPlirPFAfOJmstnwbAIDqKZ/jf6AyXKb+q/yZ93qGHGP74nfFieeQWrTJDA3U+3GVFe0qom0dM8
OjBmp9oXu1r0PX3BahiEY4P1NWnfujNkFAwdi7+dbxCzmHDvU9jqwA1RnwKrKg9fYMMV00g9G9l4
CueSe5KApJtpbfb5pOGaCoAFZ9S35ni2xmJ/hGxllXlFqopeuRVolZ+PJYMR+5D74MU7gDrRoEcz
p3A96yHVQmIluUGX6PF3bW66mULkqsecMhAGRU8laKMQrENcgb75CJ9njRlvwuo/OzIpdnPxck0C
MUb85A8qGXxAgiLvRSGrGfPflBHdDtQ/hzrNZ3kF8RsokPI+qea6R+e6tAm8XzNfxYAvzT+QOSag
4nRKziCU3XkT87pilQZZtSeGylpmylOS5BccWwARx4XVxcnH66Y3omvIA6wP+NZxqSKYFBy3OHar
imAKt1t+ELlV+LAB3Mqu5+p4fCUTHlmoW56yre4xxHvtbVb1rZsEHc0vcp6L1yu1b70LAZLIrZDG
eSX/l/StJLPFDRI4IeOWcGgaNDsa2VukS2ckj+maHzMQcbgUcTW8vO9Da42aUBKFMM6w12oJahgR
bAi8+Cj7OgfZPvUvDYC2nzubxEiaX8pSurgZbBdJDeKhLID0+0vGl3HUngdNQ6JkV2zaseMu65/N
bnBlkm6PnECkXf3Ff5HL577ipFy0VWBoo5XloCX5pUM5ITdBKAQVEnsbcQ7SvHm5lSFmYgn9h0DI
GYuP/iIDglkfw17Q5oe5LmnFklnzilZFj68w1xKw62M4R45Z+Z6FbTw1gV6YNs9Pv8j2Od3h3RPo
N6Kr3XNACKnnEvbHe14q0GAKW6TCZgfjZOy44hyV3BGegWHKH52TrKfn+Rb6cEhs1LL02ck77o7J
WTy85+3g2/ZPlGAH4y6yLEjKmsdAZsMxdEFskBDoAvOsT+oehxYJCozNDxhvZKWm6BcWW+AOqvls
I1wZbsKqqt3evisH5F0opG/IUFe0YFc5d7yFDEYMOVnfuO+O0W9YXSEdqHtkMxnNpSmVutog7GXJ
iFEaM2oBu4c1/QS4nZVVVvyt/D9ln2seksTjHgI4SbdS53SpsWnHByQJ/pXVwl1FtAgwsFGyUJmH
CxocGxfG+ZYGMjk/91CUTzis8Y6FtyzM/nI4Qu8d2vuzjjyCAmJrUj8koBFz4+zupw5QWKxqyQcl
H7+bYx1c9qJTcCxv66nkW7oswDhVtLA4pbGiBjif4Ea2p5WXbj+z1FrALTHFAYQcpijFnXwEA/hn
0G4vDQ2qP/3zSSZgAUzS/qHPY+bANdrbtg0fRu+3q0i3uXQuD8qJUHy1td1URBbeok2t0NH0Sn5x
OdC3U7tkMs5p9VGXJ1+sLyX67SkyLHBQ4adopuIrCDkgEZnlNkykzAISeljoW6qq/5WPTVbf/8g/
N1NRrPJyKS/kQD74JTnTKMtZQM9U1uC3XqzAHv00nS6jA/Ca3Mxo/5/0azBTHBUSa98c1I+rcaR2
/WYS9cSrtd3Dg246PzV6BN2Qz/bj41Fo1gciYeggD/+lCVEKIulp6pkBfiUKJlvtSp9wCgU7IMAf
TYd6RTedsWXdDHUTFyI7gPD4fnw12IL4nMcnhgXIIdlfI0lVozJzHAhSdaQRrrCw4u1vmi26HKuk
/Ntd4VE+vp06r6a05nzceFRCghjc+6daIPvtRdD9ukNefMfKzBu1gSPMMW0tiV0SjE2bOfODP500
26av/NkxjHeAkTl3GGMR37tsdpUqE5TNrEwULuLKfC7leQapbOGwpKlIn/NvL+y5XKFremO2hV9q
G6KsTTF3yYtTLrbH2VMAxqxteh+Vw6EKxxC4ngIJzLd07QKo/HsgW0JQ3JcF4dUALnR2jBBRWC9J
lgGZR7ScIvxx7FUlqLOdxR7GOqzozURm7VH8Jp/EbntKwaBDRtRcngBUqKuA/WwL3ANT58PXv7Vx
IBPfqKLztumFCaKcCXx1+UVplmQed9orhmYNQYI+miq21FGKQTwv0QKKp1VchK93rnRLFLhTQIo7
eFLeS2J6DCVew4TCBkHMQuY3qXxRQZIwSKeqBovNpG9DEOCSSeIvlRH6S+MMCQNrPYfTGR1JTSbt
/lkTM2rUvrOXhMHXH7ANxPIzHzXM7xaJ92SLc6Lk4buzUr/dtOvKX4wAgjWV9O2UGEvPlJNiHN+3
sDF7grc+/Cy5lAroicEyhnh0GnjrFhPfswcLaNGqL8ZIrwRoMymhDu9/DE1NPfshAsAtzaV1OZAn
m0cG2bdpsq4XQD53LoMdN+jaS8acBfmVUojJlksJJliRmpCBFYYbV81ud+fOniXkuwXsKv6cOfe3
ioenLK4LHYzUk/iEMBj59LBorUquK0RS+zxpl3TOtqsnwK2EbcvFQdFpM7zvTL2dIR5HEbvI/Xej
s4XKo+wvtnUqjW8+OKNg2wXtiUhOYbaKUw4syumYNnpNbNgpT/SYeImObmx1rBfRdoUP9NxfAQTP
QmX1ALXFaZFbIC+8IIBZrw1iHHSz/QHplYtT9U5euhUHOcsBfMHh2JxpDQioS7L+340LsS8eXgDF
8gxdoMN3RVsZbZZ5IxA2j4D0VdBefIby7teR0YCU7TSiiuwdqsZcw45qIKT9roGftummRILSvjf1
0Pnhp3qFfcYRYiMIRvzU9X5lNqkrwLLKBY9V2xaaj6J/DTCvqwu/a0HACHAPk3qTjqAmCl5Lbdz4
Rfh1fEu+e5iNLtYSY4uguqvvRABAbm5BCjU9ZfO3uzclSmvBtx7SRpO/c+6KU6Iu54yEUkvbDXYA
w3nQK5ZHLv+/ybO/M/PpZe97+bZMxhN8y1VzvdB3yNpN5J3lBbshbZl+oIQqTMjQ5p06JQFSaljo
bogNGlE/6DeSHr3eCqoYGs/uzo2DwHb5QG3BqBicOS4TPGuMjKl9nc/srbNmkoiJV6jrXJi1rbW0
79/gvGcze+PmTYpH4Ce7CwDyCLvFJvQyKuMNclwEmqYoo7SPuPb5UU8IbgV+cIr3AOlbrqrjuBgO
aWt702/sGAn8f2X4sBa9xTAt76QvTcQBrBwMEJCAfYh1EZ3WIy6txBgQPvtSnPgQ2YtEgPjW7lXU
OJh4JDIXKgprOcHh9XKuV9eQaMpUhyT1aAcWfPTgqsKSvdUexIMfM4iBjB+fGjJ1UqjqDiolghYy
OYOmxXWqA4GPS1HTQ/8MnMsPgPn+NNbW0xyAHUfgOZvWJ2q6lpnhWedAuX2TKP7PbeVzD2N4G8Dj
xKq36pKkL/cd9VeSP+XpzpTuuVDxjXElNVzG7KY1h+LZ15z6Rst3YRv2tG7oy8I+BnG207DvnBtG
sVKegtvF1CZ5xGczYPL2FKCa10iXDvvRcKv6hf3ED2V5aR0SCCzvwLYCMKtntXt5zOPYDVIHbn09
4qMkjm/XmtyirQqYORwR69Edk6aYw9Enek1knd9tmaOKOfBJRl2BPgN99hfYQCPQ88l8+qJdRwSK
jNDkwjQC01LeL9NlepP2WvHK/WF5JwUjK86R4SJKbEImMoYUQMb+SkmkzHxYIRlZ+9DG6D0VVnZ0
zaCjp1tuPqHmDmD5neIGviMix/1hkrlZLvkfttCb7jeGOogSPVvvoR71+MJguMdSemtqLSaehU4z
JZ/U98ZDQpVtSUH5t++UqNKBPilVtK9vG1JNNsSXdWI+ELuad0bRjTyVUgcCj/oCtxJhclopW9Ao
FoIYCqPfv7qIyHfexlsjuz5d2Ts1y6C17ecikSV1bIdOCzbNdFR7jAgjXMK858DsrCrXH4i1UDhi
mGISlQJFsS39Gs6TM3lOueZfMckEqAs6TGCHrrxvaHq8N2UrhwGNl4edkEiVjcXHuC2QUM/5y4iK
P1cYgxjkO4EB04AoeUDz+YPS7UHXlfPhk1Ywgi4H8BeRX7y3NJikluBiDL7nYQGgUMKxggaEOhDv
0SXne/yf8JVIlOWbYO0wDpweOsGlICMa9M1NYOb8YR4YXHBptYnnA0PzCtgqzpTUywU4Yfxol41D
lb5i3N45HM4M692Ki4d1wYE4tDxJ/SLk4HJpr9DvtZdfFR0i9Vl/OoDHUj+ugsF3BpIPUKL5ypgi
qd5tClnASZ54yVYH38hHMycGVoqErKKpykkJsEBJotDjUQsNDaaPy6D8jf6LM/7qjopKQpPU3O2h
0j04Jm5pBOLHXHHUEAB8wmQkSPWwOXbf2qXX/BXXwv4g8HfLIn961YUGkMx+gbIzmHzhn/mw0sXr
dNVfxhWXQB8lNCoq/eSIzX2OAAovlFz0iarTds/t0u3AnULj+cCbwTbHIp1Ns7PfN9Njepat3HLR
rSf9ThS+ng7pAxQ297/JEh4zJ1P3Lc7lsC4ZHtVbA0h7yWd7xbWzJSaQooKGFKDIbRaAmnsA1PA8
lLTUFaVINeEfsrd6fcrYrfvaG9kiQIkm6kb/dTZnSMQGzZcXH99YHf48xBtVruzFQAOikqmG6Ydz
uXGA9AZj2o6rHdilNmaHt9p4AuFoxVxVM+okwxN3AwBQYYXRrGjGwNMsUSHqmduEIte5uV961L6V
B4s4ZK1wZGWwFAxjkJWHQdUxJQlhTkW0kpezWTHsjej7B/D6jhvZkvnzeZIGkRgUEhiYF1lyLoZT
CtVS/yG1dT7mnWQ7hDgeBtwuKB7ExMKQLn8cRCUg29z+OUkOfmwb92sBqnzvzu6TMqrKGtcso74Z
YyAOLaoz2uX72SAqQ1CEA4il9nkzPc7xy4pYyoJsHqfDImWDx4yCHUBbMwNqSQQRDd5Aj/uDnQsd
2ABzKP4IZrMiQ3w/+VMRSyKyEI+yeT3gIQuegQqEj5fcd2Yh79M8gFsRitSPWMDAQTLOR9UWKmAE
cM5i3DFx4irfSjyRdgiKF0xlkDU2Nn9ykHVOkNnVo+GGKhJyKErViCMAApTTBxHJ7Pc9dxP/nXtk
ms7ta58tJ778bLHAR4DzeeVmwbAc85sG4qRys3hycCi/pQdafwV17jfdyNns9eWWso9YKi1quKgS
gQfvhg5liQyj4BwGt43hVcAw6DRGlwV1vwx91V5xB30BCR0GhByBTOOZWgS5P4kDZdsN/yRYuUZA
FFKBSZWI0Xs+01Ly8K22cPnUNtoIdp/uvyzTylKaDC964P3S0raTqPaWi9DQ1qx4cfrcaUiaR7Sl
wNijqtUGjNVVCUkQUnGKf1j8lMF9R0R6r0NkDihVxf9vleE+piRv1D4/ueWLv86syREPYMG0rtdv
Nl2P2N43ykOvL41WzHDHkI2mlTD28Y5w7+r1g4pcK9uSwGkoZVjueXYwtTU2LQi/zdysRg7LsqwH
/mG0/2tJKxbmHQAxudkukctvnPfbdN/QH/kYl9R/BIGcHW6uHkRzfTqBzTuXNrA5XwEYjT8yCIOb
yuXKfYRa4EKmrtv6IsNa+bhCtAhfyAFpYzJAFqEQUGPJf+iL5am+vYZSVLsRw6UqT8kQTcEXEkO1
LvALY83mNI33D8nj4D+8Y+qJpZh6X//OzLoRzj/mzIaguVdwLVGqJ5TLhreBe/A8oHjn5ixFfAaH
tZhC8zHJ0a5u/G+l9i6MImF3HluLRWCiNiqyuwIsQKeVzkcnV1pxYEHwB75oG21K0ArUcTpdL/BJ
1Z/mgCjaq/BqzdnkytbHIon7ImBKAlM+h+3YYnZDeIKYNUNEI/IX0p3q6vJGhqBrUvbkoHCFdgQA
wCd/96k3s2qGXkvnkszJ2lV1yFAjdrgAt+fV5eJlxZdPKRl2T4BBCzKk9g0q0EYDkYQrVneq93Q3
4Nwtg/DkZyYSYXQG0Yu5KhHLvJJfrh91ZrsUWmFYie5SETMqxDMGiAqROwNA0ua9HWbEjY/h2C8+
JLhfr8OWCASi6vR6gaZBgk0kehsvwLpdPiVHVg0/ai+EpGUuSSyOi/4A6YX3+MAU/FBG0jf3ROMl
zCjO+7Bpy1Zom+r7bii9OdaeOxZGVnenXKDCNCBWHRru49QhP8mcsOhmihs5AQRbWTtgnikUQ6tZ
pf4UZPxQR5e6nc3d08/p6a1vSvHSwb9YuRkAM93Oi05ElmXfdbmilAFDovP6RJRlTvriIH1/AmZM
DNyIQNWZWZoxUNKmNtNMkfBrKO05sSWO/IhRqrkjqkFVXndWWtvtIARyB2paK5aqLagVonXcMGdg
R2TnLNo58CPd2BzlauzDgbImoVKoJm5JiWo+v/pWupKmIxiaOS5/eH8rKXadackPV3PN7LT4gGbe
YrOamwtBrzVsjOHAbvEIkwW4B+yuPgN8/XIcIigUqu1R3uhfA897NrKRJuBNe/3r00uOB/GOFCwM
OVvih/GdIWAUedecjPr2z+Bak770SA3V99XkvpN6NIfY2N/YO1BhhzwJ2ljbTjYaxo2nmWRsjwKM
F2rLu6ZfI4r/0Y12dZ1Z2Kaq5CnUjK/3RA334VmvmsBZZeFdlYGqRzVBkeM2WzLDyW/oT5TW0A4R
qykLsOkXRgCwRYfxlWx4N8lTh6hWEX8PUyAEiBoLdRlLvU22xCwcFiyMdaN93yLL5tvWTTS46I9S
vicG+KNuobefH5XRbczOqP/4UdNKA/VLQccyNF14GsyP4OB2lalLU+ybmgABgStA35Ed2Gzz36hb
I7qO83Ft31GA9ce5gJSso1a6S0wlsFSUWkKuvfPVcTHlvXvhBTh8WCqlVBdyxOTG6K69t4o4LXUk
zU27+ZxTl5J1hQwp9XjPKb/aDrSI16uq1HBKWKjYJK2CTnHMz3sFdG8FP0M9xNRqkFvyNbBKJNeB
1mk9q9lm1A0gZB35MkPfNFxJWWrWWHEpYKZUqzFbuiprQSl5T4iAGCwi0m1zhWasVeck6o57N2+G
AA4OtN8y/WfZvY1UnrrsdNs/38t3ufCFVYI0LB55rBRtaU9hb1FnUnZemKbLQ6LQ3QIX3RsBkvVj
2TT1M8XN2h5+wcNDsWW8KsX/L5PJPyOdToYhKeqO6emcVyJGW3NaDz6sO3hcG5r2y3vNts7k6m7J
GNSex63uofNaLnSuPFHzjnzEhYSZoG/4V7RMo0kWwvRmDvvONzqYmJtkAZB/wXcoSFwt90wSFkkl
vMBSI84+x63/uj7J4StsVyW0VzgQQNrSRY70rXr7N3Mf20oq2gxeojuMs6cdV+5f0f4n+lJts53Y
z0VyGEKowoD6Rk6cBLylZyapgiBtafvXCGOKePf/plvAlyKPaQ7CKPN+6Mx64J65CRROMFQlNFY2
qVTVzQyHtiSi/0PV5fNiS/InsK/ZfVXZkEoA6YQ3NCLuwDh6zd65ChYlxY8+S7dpXV+NzHkRkuxk
Wku1rDSfClrzJEmoIx6m73zItqE8rovzm0LqtBjS54lO2HGpRIWaU4FjzQ9qJF1jdUlst5kY2A1c
LvANhgwkE4Z16nnvUmqE6qxYGrHTYMv8vW8IeJwoGEU8G+k6TZ9BG2ICegTKzw5LYlQjNGbyg1XG
P6kSRWthapBL1drCI1qxTt2PmcKjTAR+UvqcDpyf9EiP4kbUhjhOStVjZrE1b3c35akXHMfapwla
D1pZwtAZ74V0g+La7y+2D95mo7R83Y8irxjPTo1XY9M/20VJtvxBj1YUwPXEgEKucBRQ2ETFGADZ
1IZmVMeNfZ4Oq5dfTtBIk7nSEw/arkquGEaddmvLVkow/vBYMM6MNKZZRfp2tw5g9SUW7gqaj61t
E826jyJXpuV5gdv9ZGTSsiEK7AhvD5VWd5d2pC21GkAtaXVBsnTx9lNGs2cISrD6T+gVBl5JyN+k
QW0DPDqs7k/0kZfKbFlZkl5JGYg3S1JfK/OJ8ptMgcVxZUXKADS+cf09kDw8EVZvH/LFRIxoXV8f
eFL48dIjINCiOMRctN2q+GVjsRx77dB+wzbF07WiUzDRY1vUzizNuKNorYyl8TaBR6yXrBlGmdlh
OgROGpnKY+vwIwx3aqrqB7F2wc4Xc5CZ4cG+A56LWgrTubKZy/qtBQs5quFo29ekA8pli533GB5F
IqvSWPSJtMo0sr4cd4rWtWTKK4asajBFn+qMHTog+1nf+4CWB0Nr6CHCS3S7z1KSBGjppvdbZVcU
geclvxg1c5LJOD0u8YU8sgm1q05dCIvYWMfcsKTNTOBODYTznIwejnBODZ/hprApPkhz9OPPug4m
zEDukWowKZNUecrgSM16k/fXUzQ9zGSlcSmg7rBqc4rUFBenXx/BkpxdpcfyJDu0Zgm74HCCm4Sr
u4JIfQWWnKGEQVZ3Xn2+YYQcr2YXP7wojx17vlXFeZKIvQWbB1xSqic4l02IclhqgA+uFsiQTeKJ
XrFRK+jwXwJ/s9fWKnXJ4ZEniYqCt2/TdRgN+usEOCsYfOlB/yY777C9ZMSgIYQZN25dJ8muQLtL
4bUFP3tMoVcJbgzbvG9tuSsdd1j8f+z8oyAQsmpDrKyBqutplATwcZXs/LsiWZM3VXGfN0aoVIWd
nLl+jCn3ArFYWHwqO5mCMFMtRJn63C3pra+BCaF5odvYzVVmUYJjULg8DjNeLiu9aKlF0TKKgU0A
MSV9p0e7+7ZMtw2MeTMWjYvd3dPRjXqw984OgEl51HfMF88hQYnCtqecbLPn/hSZODYRsvQmEixO
gwvCfzTlJhR8XC2PwRBrdLC9Uajkc1V7V8gcJA1aUupa3z9A9yyjAOhJbjwjvxcAlvJ/HzyJetMX
nM+rM3hIc2MY9FB1BBCvtMNzztV4FCs+GN/ZvF/p4ijeYLLB60n9hnh55EH2wuMTaqbkl/q0Drpb
yvIulolu+zhaPC8Xrk9a4j494l5PsH5UrX8mfsZiyuc38GjmfnuP+/FB8zR+dL3aLO4y88zFyLHU
n0FiZy+UekHO8B6vdkfqbARi5OwSm9kN6QjMaAEBtS3qwWoaJjdD9l2yT4bJJ/+EuPv72I4sqBXe
XscrVhOjcZWypqqOaS5IAuFDe78W/eitXq8c98xNxCk3nCepwFsbKJoZ7eB6m4OW229vdUTy61tF
Z9ZgMH4x0+oLfz8Ei1lOUXpkxEYOlgPWZTHBjWHBmqnE3H0N0GI95YxOhA9aL3Lb1fL5O0k1PnlL
5ycA3VopRK9XXpOF5pR+TCkKsakyTE7zsNceZuL4hSa9SQYR1R2wvX8xcGCTfxCw3DvSt0OSdNS9
BOrVkMM/is0AxtXltMn9zgMCFgk5J4niEe482lNF37ls+ZEEWtcda9JUuJn4QAzAPJDiUCpzFjj4
rgkVgXwYicEpcp/1CGISv268Cc4ZYJH+xriDXccVJtFhQM591+ktDYhMqrQ7Hq1QT/8rr1mO40aB
jT7hxi2dWE1dPcMex5lYuTYDxOHFyf2ujBQ7r9mhSOjTitrT3QTYTO1AJhMw/Ov5rmbRj15221JJ
SkG5NiHKltDU/E9v1Pf1SxfMovkTLrXIiNl32/4kfUXXo3aATlosboZdqp8yzbQM58Eo2Znnw+YM
mnVy3kGoKhly4VIrwSWaPXULOHSBlZ/gk1wWoLRDrClHfCGCIprTC+o5uSZLMu9mrOduRaF7eQVk
DVq4SfX+hePGCIMwjaB54B/f76ugxOKh6uv/4vwzkVbuaRBsg9y8QJju5wTej+kf7KnHMJTM6+Nx
WdCkBjNMOsZ42qeR5BCuOzPrQpfMXhk0sYq8Dmp00VOjoE7WJcFKoGdNW78EVzHNtQgt4ZNPnm7q
/6FFtrNq9ZC2oSRf7juSFPNVTMrWuRelCldgqNBChwzEUTswdAXgOrp5/+X0xxSuO+IyYzlsInPC
3oIZbg7VOHrWP6pR/tUUtFXZ0ejrMTFY6kO5A+LPDGXA+L6/ToOalu0glqCHnRxK1ONYCw3jKSWt
P53mx06t9ldKqKlx4UPxodbvePE1+OZgaqrsdme27UEb6DiM+y+MrodFbJy+686ggtgpWrFnS0t5
3iCdcjCq9OMBkjv5dS7KkUdZVITiTaag2J0o7iss8+KWY3VKJqCSdtkWEt7moHefJ51ON3toDtUz
4C1KHBBSwD6IaYw2MDoubYVRtbfln9nRIf1adlyFDuqiTa0VpBkXlh5aslFC/AZJ/FyF+EQibeIL
pZK6lBN8YG9PyG0T4FzSTOdB617PbzmmaE+RGygtMdaTfE/H+7e75afMCumF751aTcgVp2F3jC2B
JiapRgGC3Avip1e9SmhaMBPeT7GZ/4hvleocvy6R4kh2ve69T1AoIO9weezLeNFQjSCDaz1rs/te
bco84tbA/zNW9nl/sumXG9gRN6cyufk/AW2u242h/964XWDnZSp+fU5kdw4VazW43jxlrP9gJnU+
cCcDYWZir6izc61dYTLQmpUOZh3anRn9mqofkk5gBkJw9N8OBjzXLkT5WwLzyf+Md38reyonQD3d
siXt6EzNF6EN2WCePfX3hlOZBxjzz9xv3jPlfK8yActYqXnueqMJ1lslTKAMZnSY9mWavd3QO30Y
xpYpN+qdldaXx6IZaGN87yb8wXplFLDXaDcNvZikSdo+3r0aCWso+kICt7nCHy4TZsvQa3rIyYKU
cXR0dOe6flb4fYcFbi2y8CZFVoCZFXPV4P8gQUZGcv3N9/ORDMG47lKLM0jERAPGIOyxMum9JtJV
ShloRAJ/4cjEmUkZwR8jYk/mJQh2O/GBMb1DUMFg6JX4bX2QvwJ4OCqP1v6ITwzbwCbtP4mgOdkW
XnDS+pb21bBDaOYltUuFWb7nAASB9Ko39b7Em/HdeeLuadbhfXSbhAwi6xktDCNp807LQ+b1Ea4m
4yzYZOOmOwjexqikDUexHqQ4SMKrDgyF7krjBaIiGOLyMHA0WDXOxcCEBdFmgBg76gAUuGrYhAiF
0NVo6/feSMXcOfIi9C5fzav3QHDW+bWnE4zncGoXmlkqqj+9eG0syMw+jXG0QPr7T4SsqJyDRYVv
7GBIqUXkMC2i5ULPMnKkHUBdp6r9E3JUEsRYE7oyBVFMp++ZZdIn3UcKelS8TU/8TcdqL7UwL6wL
jGlSYQEo3UrwI4iF080htRMCv2YmpOJL95p1K6mUqqLyrAjAiLAqBP1Kcwl/2rRrdSyFIQuuvW7P
l8IEJuSUdzM148YHaG7FVT+4/6PGJE05qB6gAwidwRkiDiAW0CuYm0prE+PN+JYrdn8olnBDNefo
qjNU5Q==
`protect end_protected
