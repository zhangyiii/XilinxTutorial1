`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15344)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/Y3
LeD+qw2K3LM++tksXDWlRgF/znF+Jw9c2JQAPXKM9TKRvOl/czmCOhE3aNSoCh1FUwlKG7QK7XW5
1i+Y/6fuS/CW01hotPrez34/+2hYr87se6GBDorysLqVAXMsLY/YV9B7HhDUSw8jyNyknIEmI3U7
WudHo8vhLWlCkMQkDcMf+Ivoy8TEGZRjbwDtOXoE24Tpyh0y7Szqp8vQqEDariMqKoVn6oTmJYLq
2DpWhIEswln6tRI/+zBSleCqwfAdmXyYA/Icw782kOJqC1rm3rVrW/fPVK8K9QJVLjxlLtCOUsdW
MXHfW8zBcf+OJ6M5Ps5WfxcGaSo9F93JhZJwtp16qQc943Z5uL5S7F6uhx2/2/JNEiZKR4nwO6YF
9lApKneiqiV4lMknv2GfPf3Z0yt/epCJ1D6rwzHUxOS1WE+QGHCe4rtK8iJJPU8gdqWBAV0E38zX
DrRSC8OcTDpaHRsM4h45UtUZ7QHuncOnjyjfle45UXlGJHuJmqtQtKoBHlkWLaWs8IxPTRJdashu
kUk0S37b7qinz8QPzVNDizIo7tt1mrqBCLYTAlFjqwSpg+Q2GoQNpEbhhjJSmvYKPuGddRJZO7Wl
OSphxyLgZzVvmxDSH/t87kHgGHsFgjp9dviohojl/U/zWNmgRey6ALjcz02ZkQE6vzh/zBsU36oI
1XLzZdPOsmsFTW+hi0YtW4QXrws+XJn0lDvqAm7a/4zSUan/YXPqgWJAp0UJnu6AAEQbDjLTTbka
rmLtzTc+KBM7Qh/MrR0nLXOt+vB6+4vpyFW6VF57FxmXcsdwTMv34b7IGNAHXV19xTd61xcwO0FS
hYiDkPuuZYyI4HEIp4JXLUgW5zvyHVNvmOFASRRNUBRiTkDYHnHp7Z/O4tBKX1n17fF6v/fg3mwS
2JeiK4If3PXvktkxXJaPGyiZmPmt5A4Bthy7HLbet//JHNLV38xyJ74gKq7QU9oEASiPXGEAhbM/
x9I7SkQ7MIJFc8uqyxac3MnFNurIiDEeYdHyaMERPao3PN6xhb/2oFOdOfTFP1ukLGNEUsk0hPd1
LgkUtfW5A20Gbm2UqEhuCsZlhhN713pRuj/0GuH8RmIBQvAjd/LXyOWfuP01wImCTKOjz7332xEc
vYTB2ZLyx0dZNiESt3YthzquQ30BRv2JZ/yMS2L3RICN8EY6volLZIQ9J/ZWNZnto43SN9PZ1A4d
KcVhHcitoNxEjWlorIlUHZeWcgjrKzRKTms/5Qvq+XK9VFq4xnGh7Oac9iup4UOYCOq/mhqKA4j2
JlpoYNdiV2q/qk1GYiR9lF2o5Ecimhm4F6Qr/f/9tQ8wUUD6qfkiHSEpOGq0Z+43W/6hQ3pmdtRH
CP6CKYahbYpyAC5P664kR3KSyU3BSn/mcTnKBa/6NWGyfV/dwudwQZYVTSGWPphViyNhg4NXBZdW
VpNjfiNyjHV/WD/NL12VW2Cc1vUJznM7Ohc7WOPoxL3rTVqMbdkgPi1PL7rVXfy3t8gZU9LEOkRW
PzJtI3ekd0GtH6hpTLnCd4KmXpUwUPsqehrqFsbkKH7YNuki4EFBpsExEHrPqDWOzpH/kcA6Kdrc
YH3a3yqe7rPGOTbbq8kMXtkWN+YItZVlgy9BxRaEYkXkPwPE5k9IeceOrVP1c98Iv+echFZLGGt9
j0QBJm/V8zqFl/WSHqF+eE2suXsp689eqNMH9JYhg2llYDoxhhS7WHFNPfDyoEWMj1/FlOG8ECsl
8hbPn81Rxh9ZGPDmnWU1rLYxp70uYzLoDW9knjjlU7YCZd0swAJvYRhXsXf3VpO1kz3iv6W+nZMX
Brg1+/LfOSXBphl/YIzzMLzLBGrPVYuVX6U60QduJlfeyJj/jsupLa0YCq10Y7+A2WSQXESFHfnp
Oo1bNau5NhQE2DlB0tGBKT9+EPIslfIrUiX61m6Dkfx7lrqNHGsqror8LWJv4D6YsANdMsKop3y8
ywyUOABWxCDeC4c0Mvj7ZXbQ7mSXzmcBcrunwbWP74A7PloqWvI7iteJV7lKc7ctjR9u2w96DihV
W/DwvdUVHlOVlxCx01PJRop9W1LKbTZpY/0ZzTe7UocPsy/89bc9AcwM4aV8BP8oa3Tq0MJrZOMO
mP8yNtdJbBItrltMSYPKOFrGF8h5Z9v2p0WPw/sstYnkE2z48Rw+6hSemnVMd0wzek9T/E1AS1oE
ZrA3f8QL4jIonmJyBqQNSc2KVR9ezwV6djyk6MGEmqbDiHCADFai9EZ365ggEep82nSHyOwH7e7k
WAk5TUhv+Z/kHNdp52dLfVakxOtEHSbneCdm8hkeGJ7HytHDkfG0EsgZqwM5A1W/2scrmPjhfeMq
Z5gZil+FLHuqDgpnlqk6GwlHJoOLR6TnOa32UQ4VybJP9TMmBagp/su2C8/eaMBKHBuRVk39v7FX
8dhO0ZLg26Y43Dp/r3gPiA1p/bUv+HokNtQflnLHrnfgcNwAFuo4ChGQr1suF+/6MEZ39+YYcLQX
aZIHry63MB6k2POVKN1jUp6i5HvsZkxmE+SYqfeSDdTzqzoy3kdlF3NsS9UON2EiPWysa2Qu1opo
tMApEFghS37Yp1yaPg80jFeZRC2laiYChE9ZVjVUsteBxyUf277ypkGtcghPr72TPqQ1zQtbODEV
01nBZ4KzeBhaYwC0n8+Xh271Ug+NcvgaVLmitcZexDBHRfooei8SXKptlrX0Oj+5f74mAi29Jmga
Yl+J4Ze7y68N+bzIJgr5GmTFfbhcQWOQtM+BOeiDagj3eW0qeSPaLziyW5Otu/hbEIob2UQETk1p
onrFt1MwZK1hw3fcZGOjClWT219Jhfuyy3lsb9z/1Y0t7kkhyoXH0NKDKRuDurkJ0bKhY+0GCyGQ
H38L1GYASu7gN5ku/Zk7VkFeHIldz1l6oisOIKm7UGg0hicb5B93f2Pf12QemWqxMQgJ63mSrLMV
boU5NveNGoLsYDtDnaV2YNF+CNcyA/sJMBZrLAgN/9Y9uAUXs3U4HPLd5x0+voXUhAbX4JvYJBIt
lCVF1LiQZRVoZ0CoPFcTPy0oqZf5t/B0waoz6o3QOXzVHLjS+SJmInj4IqzXOmBxM6t77U7imk18
bLYCgkajPq5Q2BsG42RmIsu+QPpn0N4hg+BdsyTRZhPEP6EAVaqRoVBNIdfJ8gn+tTTv+OCdZ0fP
wJmNdiPolTNcs6vK9TbANpZeWuI7a6qtgKNBsOCOdc0zhjb/RF52S1BKEBqc42VuGhh6X5yU2mGb
ruL1Fd0poo8hfojdBetT9uzutJqvFkx+1xuUUrZIfuYOY3VMlY5n6iS6tCuK8VerRYRMRQ1w3ZNW
TjZmBq0MOs3B64bLdjcA+Cb5wKYCtVDrfS1jPXCYnY11vEYxa0lbOLvnd2vLtQkTwluYDygDt8eR
Vy7ZGhDBf2KaHmfrIu3ziboSQ5DFEaJ/98YCNZiiNFKkMhf7LI4MzhlYsZmfTO1rnyW2+tHTEJNb
Vm1wWgpcmdwKzr0Rhxk2U5n2bMUnlklQo7Rd0A751/vrh4wBWM72FBav0E1vSc/Uk7q1Rxt4CkNw
3cc+TXM4ba0WI9RUR20D3i+E5uc8RgK4mdiG3Xdej9xXm3EEVLc1/7WkFLICH/3coj1VjGG92Vj2
XccRw2DDMcGnzd+kziVpmJ0nh2Eo0HDQ4xp80/oPecR3NSVNrGXFqVRnBSu/f2Pnf5Y634shqAvt
Hr6aF3CPOBpbbi8pcV+eJv/kX+fqiaCbpA0MiJtk6FY+IhtEYOC7uSf07TBBlpQuCRfHbt/spQ8s
bhkxVveVpam1mckRxkk2SHbRznUfebNmDRoIT+4Y6plhdlsYMF+zTcGKIr8sdaEMJnjF1WzfCyUA
KDg1QWyzgSPTSTuzaiszYgYdNhnqC1+kYZzR/M3YiZalajrP/05oE8Fy77KeGpzLTx1ifD9HtfX6
lYwRXFkD8U5iurWvuPACHmb9YtWHXHpc+8ISlo4pBG8SqO9axtSXtja1RzfrRkHe2m0+cB3nz44k
/mzpz+D423Ex+LY4KqJqTWWjsgK16vDfRaA+RkW/mhXoTFriZUGubMtkeS5FLF9/9rk0F4ovlf2O
Vl7MFbPiC+yJ9+HYfAkaI7yMSDvQs+Iji0e82ZYgHmhV9FoZkOchgAQI+dq8duqeV+AIxztHhj2r
JAXNtsUPSmIefLqmbGmxlNLylHaj1ZvfTEAk8mEiDpMqZu1nmZefBwHu8p9PMrfe39FbXCIJuWO0
4gpozT6UVAd2Mf0WX1d1tj2+IJ3ZPyh3IwJVDnbO/hxuafQa1lR2WgPEaaK1w1wHMDqxdgrRenlH
+tsLxWhy7mVqfOvTADV1hPlQePraOLm9qld93viMxfukItIswbwk2cubLOL3dVcgtuffL8c8bLCV
elJT2VE6teRQri8NfZLuP1UJJRuJba7SqVdMXCzPwAXgFBt+hWEPbvi/oPDmnckECh2daTACCTwi
FKnf0jS1zZwwd3S6Pj+ep40L7x2/9J3RX8muaNFITrSEx+U3ZOkpM5W3EESHeNpkgHi/UWd/aLON
/3S8tzK4SnYqts2lE0xQ3h0wQTQqB7TItL9nY9p8g3INfD338voL76qxWSjEkXbbOkClooy0fU8I
11RTx8YB4V3D2cn/dyfNrUb2uwGXEjKHlSCeJRqAoSz9OQNQumj3LB91/+9tYZbpoZMvOMA77/TY
fIWOU/BFDjxYpGgbVXEZKF2OFa6NFsx3giSwPbtrM2oUeUNqqi8ENOxHSa9VlRZoLTJeEGCCp5SI
zt2REBcaexc204qJNcbWYe2lXVcJj3QVMq7hGqe6DYV1DuZOxvBgSZrXOU7wYetTwoxKbB8QSv4W
uSiZ10Fqd6rPcMwRGnnzaVD971CnqpTvAiORMwGc+NA5CyhAO7evhUXz8kUpa1nvwHc3Rxi72R6t
7ge45Msv9FONFF7cL6wL6vaqCf8rCGC6CKx/PGG9wM8+pZHHAkyMJiCIu/TmeT3KOFgp90QZ2JvF
bc92y0z5cUY8qIMvgTwzPHAKh8zSXvhP8Pgef3lioPxS2tpI1Od+VG6P73p3iSrpFIymH3mM8Lf3
ZLgnsHkRTEVHtd8i4QDLNxQIyEsXZQcfsS8vndLzkuDX6GZ8kLyxN5cv9y5YSxVdvTui9TGSTs6c
KR8xGq4Lhk+oppJG3hx27DW4Hy407z8s5+tcfNfHVGLhrQ6bEVw1VrolNDGnPU+sd0kREKRPZp7G
5ynWT/GokjMXLeLrkv3451gFxcjIi88tb+rlkAgQjEkctA8/X8N1eVKP8hk+Ha1iu9UBKXGV/efj
LrLzRJtSrULLhxAP1XM9stxNdLFYMyhFcmc5lZaQ7laYJE0TU3Zi0YdA84/BD5vMKT6rrhKqMtC0
0qMbfFd8/aaf5tGpdD2Rgq3SaQQcrm/n6eSY8d6vQ0AjNJrPnmg+BX/tuYCi0n8kjjQMcaYGUpVx
AqFKdhL8FYdEn/bpgWpwCNfsLP5sfnp93GSfZO6bTps8kbM4EOtk1LEsmmCQ/S9k/s3u/gfIi8qG
9cMo3Zf5CE+gb4DUFQhA3vZ1lZZ5KHuLAJqMhtt9RZ4Q09C8xrjgvVXW5SxgC+JxM2pqdrkQgS99
9CY+ITJ6/ryggXK5VL64rReYk5AUGgg6fFY/Q/D4VtiNz5KUHNoD0GnFxOmXSHNXll3IwQYx3aw9
yEqAlHU69sfJrYvxrsMMo0Xj6w7sJpTSws3J2SXN1jk/2pnm+uSsVePahuWd+KkZVkmR/7nroBE+
2nSAtQZuYh1jMkwzYu9RHx95J9hpoZytzYkQjkgF61xnE1Hh3mWOxF5uJPG1qLlFUCYhw8MCDD6s
2uZoJSktLtJaEgWeasyc8+GSzto4HNZJK2R3mWht4IgGxuXvxf2ttv4k6JALHANSCuFMUrcTwas9
7cg4QqMHSD9ofpUhc8KcRoV1ferdxw+OgobOHIbmutrMrSVU4F3jPLi6yYAOXKCAhaKRz34YMz2X
Q81VgPLMkPafdakysPkZc4HdfGXOukqBzzestrjujvdjgJXtuCmCGcgB+3GtuL/J0lLpf/VFvf8W
oWDSqLDRnSde5EHBdP3EIv7P2HOEwuWiH/dbGzA6jsM6YMCnruOFs0SIDtpIsAjuOhUWfIKYQ5FJ
EVYgd/vroTC4t7nL+czkJnVn5Td2gybwxb39wWYgNLMQOxKGUBDWXti+EbKWN7z/lBFvnxxn8tf+
jUUsHUf+7cS26RZofgzV68tEIAFZvKj2qPv0hegC7lJBaWvvskLwql23gtNGMh1qFTAIBZU+/uY2
9LIrlmX/yYbu8VKBgUqGH0VjnZj3QkWnR0PyUGFptSqF9GZmxixEw2WdBU3R7NPXJ7vg5A+DChoN
1U13BK2fjgpo/crFTsPYNLEwDzoIdm1gfixHhLlZzhK3M0Ydf4kU+JH4hz1+xBoJ9eg9MvGWItsC
MC8oFIZrDLwGD5kMRT+rpuqd4v3CDagzrIdV7wrEFIr0QLbXG9KQVTKzHC3JT0hKlhEYZ8+CAZ0I
XthkWUP1iKRXWnaer6KbLX/g/BnLAQCvdP2I0PnY1gjSh2LXMy6TETzFdgiijgmceWJEwSHbuI5d
SgAtJy6PVZf1FYn75H1PR8cvsTmHxUj5mUvw0FxfBIuD9iWYznpAxx4q3xI6Xq4p6r3yF3MPIxkg
PVio+pP9ymMpmH9tSSQIQirAAN1TbVQgEuaKdw7MSxMmFYwzIO5LzsvjMUm0jYnhlPMS7Tjx7mHv
nsl2KkVNjgp5VLasSGmgS8q4emPMZ2cv19jGajATyoOPZXqwEvDYUxSpFJd9mld+gMUPsrCIwI4w
tkw4yOeWqC0hsfIcjuf42wumBBfTEJGt3rgSEu7Jg7t+J0frbZ8gCVMKATAdJYsEP1k9c+9BYbOK
ifT6xeNxuoEBOAKHCe/UsNOrgBlkryYNvVhLZnlTVfxA8VowQ9j1D6xg3xWadTHKFj86MXM38BE9
RxDDIIKXfC46zdxdVAeG5vacYqEPJ7hk8B0cw9VIxGKNi+jeSb3ZmYT+TTa/9SpNZJGH5EZr0tXR
u7cyza5aKjWAX36N1Q4pCH4m4pUCT6p11r3MkJfcxJgn6tZXF+rEPiDLlkMM4A+EyiAbhqTrFRij
muntFgI6MCk7Up/vi+PcPM+PkU5j1BED8rsfZbs08OWQlu1Bx8vHpQHCxkvO0cRO5vEl1RQIrac0
yvBCrO5nh8c7M/52Zptj6au156g8tuU2GuTm1/GOMZ/Fbs1ohKx+5m2iWmz3cRWcxisBj2PYlfoM
zL7EOkhHxMCH2UjZ6q+q9CFRxg8a3ELv0LtqPEq3GPBB125OjTYOghHXzU5GHEMTTaSAQN4ggVSB
S8UxEToQ/y/iVE7g+jTmqjuOHExgl7ttz/EWglt1q3b94xCvWgAlxDHzEp8dHazHcCiL0ka61v9F
kXYvEUccrS1+aqmQ2ATfehgHlRQfrV9+9vcN3o6q/IP8K0VduNroTjMaEHCloLcyitHT/C8BDYZl
E1eijRjwd/lmDwFJCXOn1LBMPL6JA6UQ68nz8CtMk4k5+HBQnpURexECzKLgXAY/BOe4dLGwpo96
N43saGdsXfruepS56CA5wYO9E4axR9cqlQ/HhNXR7bNPz1eqe/XHb8U9PJJQCVBT7OawNagWRkHU
rTcyJEBok6KMC+mGdDg1mAS9lJ8cmwlcmsL8hq/errPBBmjTW7epAyja0BhvcWS+zBGxJYcfFwYn
+EGiqYmAm/XKTbG7D4h3GyPtGrE6iPB7N3++olBK1wzIvKx8yGJvPK5BOhIOmzI3jr/rcs3+kQwG
UcHa17278i9F3XGo+p7GPK6fue+TRiY1rM8mQLUJgPjgOqHw+x8+thri+nuN4fCKJe3f6SvOeRC+
eIvFgNp5+LjRP92MCZX747pFPsJ0dBYtRM7Z08q7ru9coMTUqWc4d6tmSjtqG9dINmqBAPiviK6i
m+Lr8EBHcSCovB4NPm7VYodlB2fBYkzxDqR5N2vMbJywfpPzldVrAgdXA3et170vgpZHe9p7oXEm
1m0+nqnpRUycO4kGqhQirArYtpj86Woj1Dx5whQgeBA8HyXrZSACIuSGLg9qLz2BhUe7p9ntS1ln
fjdzTIx8TT/emdIPk/SZ3R9eqTNbZDhHOuc7J39qPNYU3Ey+R9Dn0aQM9eLLMRfZIDqdTzS/rVAA
QKEZayL9UUpGSZj8Ma08q7v+8xTK1JAluNqYdUicraI/MWyMubndd+cw3Ksh2SRx4g+i6OyOxRI8
rET0xFD1uv9pEd4ME5dgh/R4OQxnN0bD+onieJcsUG7CFm4km/YVFxpjlQNlY2xQuxi9AH5eF42z
o5LRoqLYJXoijUH6YsXKATDDhA7fk87KCtemK5gXGQgObs04JDh/bukCXtUhOVxh0uAToIQJKy1G
sNX2eZsc0HhHPh4FWbRrlrKbgbO5UriyBGk7YCst5yDxqsfiHe1puCUzNCFFTg04vzYZcydLRDrl
F9JAYMbsyP/UhY8ErZmDFGqIIyFp6dSYQbotHlIxuS9FedbEzuGuGDhF2jAV3LxwUrR4uF2wO47H
SdUIAP7N45uBI4awqoL2J08lCRHfieaitW9GSW/4UIn1OBXkq1FYqHQm77pTAgH2Q0o7grrmgsyd
GZThtbcmmnbDnp57bFYP/94PexWvgot/FEdCKvOZMDJy4GitLM4K17aGb/LveU3XqZUzLo2HDoNA
OO4giamRiw/GZGW0EH3fLc/w6MP4YiGsX6zb11v67qRO5iWUyp9iYbxedaJwRzSAFckqpccZkJ3o
FD1l+TAd67huEGWI3H+t5Ju0jvz3RE+FUfluYZgWVQIDe7RqD4v+jErLwB6+uBMPghii2heuhwYe
BaKWdxagNEWklkIpT5Zg/qKROjp39mtAZRl+K/FWILRKvmvcJtnw5F+ZdItJRxFRYWZdGCEX+cWQ
HaPsEhV+EOF4rc4j5ImuvAJVKmwvkaRRQOTrJZIExu+2ZhU3hOoQfE/dTSOebQClOzY9ySw/tFJM
/dBcz7Zk7u8yKUOjsEZpd5B4Wk/WfdL6U583HLN+Vr4scow2G1ZmoKhxSjpDUjdyiFgqC0uI0K+p
P6EzUEi4nn6elHlARgH44NP3dBNEjNrrZfu7E7rJ/ei3N86KoDcgWt1an+b9uH2t2bCkKGX1/ATP
s+nIOQ31yFjMQfdkshTssGJXzDoOTvxZa9KXMpvRX7bYSsndkCqngcPDqH89IlK002cN3rb1Thn2
A+vvXPgJzM1oT7+E3gFgJThJf34SnxGGqMaAj8/Bw4wdvAnjC3ojnjtS6x48Zjmt1evmNotQ2Z8n
1zKCNzRHKehDB0RqTcQ7GSr3rTpYbdgk/u+8Y7aOM3U1eYiVKe1WPBKaMNYUx/rU/IV/fIibQCAP
aPnA9xdTalJVFmJkH7KtqUD66IiVDpDAgZ1hFNPLQw3KlM9TUjyJ6Fm+sXISM+/Mg5Dy4Y30ipVH
1XP0Bo1kum3MmZbLFxfOt6rw6UfJNOQr2psuhFeNXtHAHl/I2hdQwi6zr+x40mLXSnRffIfaae4z
MrrRQgXD6fz7c47KdTJFfvyMRLAQwjDMDjp4EHcfCan6iVbuoLB3PsgyJb7KL4XmzH6A2PerqFu1
HJ7oCmPpTmDLif8Y+laIrZ2DQ1wDo703ru96IhYGj0HZEytNZtMgnFLjSaYxquOVat0aOywhw8n5
S8NqQoGGW7EkBh99QrLh2uha/kDfDIEah6+TDDOkN7fJcBzvWTgH1CXa2ahmZkMiJvZTKrb/4cBQ
KVCLKvNm96caTIjANA0yJW6oG88WIn08XQA425fgyuSOmrYf8Jmsc67ziL9Y6nMFaUkVHpXNus0S
R23HeTAfIF+pB5rz58mCmPXfbiYyA/5L7TB+1rtf3/2A9Iyie0zRvjCfCjnOCfksFhlfriF6YXe3
TgXLtSaPEYGPghe0IQkSIjYVZTGEmUguFwIslwjlalttG4m5YCjiP9W5ZMigE7B9lollBGYqq8aN
gfA+qZfUnFRooRqhtt1xGe+IogUam7mL9VzNzlboqsuy1r2izkDpiieWpps8g2na3CSrEem/QoXf
TAl2WqVL+EQ4C366Rrfxwktm1OpijpMKNSOQCqFpr1GVRjdIAZjyQln6ZBStQ9nwcHbaDo1qOvY4
7s6Iajz7hd79oDhd1pnwAOljcW26Eg4zlTWFzXMjefsA8kbykgIs5bJhmNn+uD7vqAYy2p05i0Sz
RKcabk9/bxME90CbLI6HOyrnIswfU5dQt4I0S1AmlqDeeHLzfzEEh6GN4Zum1f295h2A69iKvLc+
bh/zI8T7AESdpE9Zm40VxH53bG4mC9vmvbIuHQfVjf4Bodb3p3PkhaQceq4Nis98715BA8dCoo6+
YsJBF12EU42RkIIBmipNYKZf5TYiTlnwyazByzNZJPo/FZ+QmBUoU4LmJjSAcahE4c7e4eQkWDpf
poinYYhToVlFYLUjHA9pQWjKBnWGGF5+3WACkBdyxedpsRRtcmtlzRyjI6HX4+YSg5nNWU79v08h
N9IQ2+/RlB93o0D7sF21Suizon5NC+x30hI45EvhYR+8HQ/hjpoO7oRvRAHQNfBmCEldtaFs86Tl
qT1cfvBkNSijRBHxS4Df5Kcw7sWTfI81/4Zdct8CfFnBqyD6Tq5zhSboXRpZ3ALsv5tDYU+kyC9K
RpeOtMoBzEll/e/Iv2lmggjzaJcxso/iI88En4FsqecN6ECVuKElfcboxQYPPkctPugiCKVVMTRq
Cvib+R9UPKK0AcWn6PZXYORkXcluRSKzc7wdU6gwRfI5IUUtw8k3axW1mhNXSkPH/RUAdTyXiYF4
9yVhAA9uGhrIewAUlOTftBnVm3lICo3SIN6tnrdFh6FFNVACDrbGPNSUXV+KrjX4IEyOfFOHodgV
yAT+80TKomRlEqJstFdgRuZnqbj1TAWxDpSHMv6Fogj/euz3617IJxTUsmqquqeS3l+COhPBL8+X
BLZoXcKQTbO3pH0TDl03bK+w3kmdhtisvPzld+K2Vcny7Z+crVyTMTee4hyUcnf7v7ffNMpfa5tu
oGFoUEz8FUSuNxxdLc1cyxP3CJeqddPyiolfdg8C3FK3Ya8WhwIi3J0INaGT6IROfccbSlHwRTUL
vEiyxAh/y9ONdxx8WWpbUrw8cx8S8bgfwrOB/KJyH3psqgF2FDMEuIkhvlr+9609NMLd2r8UZTh5
l6JJcjRTK81MAB3zNYAH19wynATbpSq/H5BSKcITu75YjYIoXZ59TYKgaHEh8YT5BlkW63hvUhwo
yzHTWHdvisw54QBYOErhZQJJ8dkUgzkRFEDIAxbVYT4vzd6F2obFzm5m5nRIhmK9k0FAoJlr8G84
KipHD3Bhp0fawN04tecCr5JvtbRgBJUqrRevgGIySFrslcVD6Q9QpHDLQg+LtuCgA9tS6SrYNtWQ
xi7gmiwpoDKmhIcFxT+qji4RYCA9WjtazgGlapBTFq1iUqhjD5Un6/vHm9PEXSMyivudb17PZOel
9rZ+XqgmRRFRxwNTnwSJ941WfMGIMSEJoXXK3lf6/91TH0ZhlbBTkIQ127UW+oqAnF7TU69OumA/
+Kuc5GmJXCD+qP11NMlxmLbinSXEaKqg20ia6A1juFkRvyd3KJiu2H4IRmi+wCidUL6RBNjKu00E
hIIAZmzD2pS9tY6RU/f1Xf/KKhlRndDzTckr4q6bqErO7Wno4YpZ9h5xbtYW776C/SapheA8jvSU
xHChKiOc/L3DUEEIZM8vHMUwTi2e6uUvJn8n3CzzUo9lnCRc51rWxwwMsTmx1iVyuMWISFA1/CQv
UQwpdl+GKlpMYOolJGefScgdw+5r9SgjLLe8blybXKWzAxm/UXbD7crHzVNapWcqWz5Xwe/tmCt4
cYuuIevAFp6baXmq06fMwx/vgAAQlhIKjAV7vjyRaPvBipnTu8sFQIX1T9W25Ft4X9wwpIjzbm+3
4JR3A0fALAJjvOioOf8PksH5Op/5uqp9S1dElCixBICv5pcKbONGF9BIcEYGfNZ+MuaRuVstpxjH
K1jiH9lKnaWfUkFliJ/nmJH2d9zDWjOm/EnUBQqb0ZOldanhBzmVbbaEeD6Nq3RTUyKxCXcjwffZ
SZQrTN4imgY0orjPcCkrfp+oaVtH8q0eg2mYD+ML+Fjgm5Sg1ycX1IuEm/WGa3OZWNDuZlYP+IKe
n95h7+Szb0TQiKtGLDIw6kL/flA5LP9JxkLEvRH/5FeGm98U4p0rKFUZSI98p4yWGwBl8yvvz1W+
/mball3b4OCe02e6qccc06ZsttgN904BjXm03K458iqnbudrssErB8D0LDUpfWxF+zl6QG+sNhVj
jdWU0RIsceyiiX/3NELZCA7WLa5nK/q/4OQGbQfNwymgo8dBfZoeOiVZqC6vieeAQbNodeXJhVW1
enkZHXHQ7FOixNvF8zDYqatGe78gvdwOQkqfg9zp74voaYqHYLRMMCnmMXgPxuipFDca8KlEvNiC
NSQzmeoQWwJw9qibSrK+8DsykIWUJUugEzjf26Mz3dtL6qNl+8V3ZKsaIPqR+qSIQzF5mMec951+
D2ixwGbtRLV/dhkXqlfdB6gfrRllxxuEUOorg0Xs/wOHeMh0HF5VwBGSQkKuFJ/j820FftYEI7/A
aoxZmW4ja/TaJ4N7VpYk1akCsaEyaQI3NrdS+rA5LuD/cWyQDmAN7dog/49Z3weB9EniCMZtjp4+
GvkFHo/XCmk7FUl9/Cqzd5ZLng/fp4BAeDxAbDl0uQQUUd0zWucHtqVujMLs6+f9Je1CvZZXzL6r
1jGz80rkPS2xN2tL2BCHg+okTY7zxYGapSVZYZ+L8Ptanf2Y+VOG95IzB+p8ZPR/RzzrcaFlWqsB
fnzuKTNqiRWEcyKM2nDfpfhYWl1N0PkU5JkezgIAdadH0OCna1XHf1gs/FhkQMxswMgodxvblThW
Mwz9YKGB+uTiJQ/NSsdRK0Gbp6fYRHIdHABjZNKx3BhgYcsxiDG7Erp8mk5gvcF6gefWYXkuYNJX
VHVkzYiC9P24q3t8OlIM1ByiWxGsrE6GrGFHrzHll2WmD2uCaH1Xh90Gc1eCkkziQdkjWAs3tvlk
fYttPNO/2xu25/3llMg+Ur47TYX/iUdA26v4e5vfMNJDi8NJn0J+y36XihHhGofNKXI54XtuEwEZ
FN0kfaBcnFD6c8u6iIiTuKTmkPrXWMD90aUJ16XJZYQAJ2wsUVciSCGckYtxdTqjCQwqdrkb+jjQ
JkMfsg17a68DbC9xPw8o/rd0+SF3NnTwsV731e/1gRV40Vb2pbd8G8L9Kqd04vo8x4MvkUJSpHlU
sWXOaj+4bUp3v64nEGtXqMbHgTs5dUui+LmOtBNDZP1CAMgKr2BVkY0/iQ6HK2d3yQbEx2vd+moF
OGw+qbLALYwW7mM1gxjcjELbx3wLmPBgqvA01BONvOhQgp5l/l648d/T4kxj/8nfQJQ/qWx5zqSO
5Jr7zTXfGU0Au1rQFYgv9wAIKiZDYvCrGSGlDhFEskPlN3XugbHmFxhK+eaI2UN10i0wRNFjdZpY
JEISC0L741xdWZm2etaEwepSiaimaqkYktpQyLaNKThe7zLVrt3iM+SRaEvMfr5w4RuO8rI7dkIO
Pm6C0wEms0U9mbeDYrZTlf3VR11bwO2CdfRZhFpJzB1g1D3OUnp9uatUnFpeQtaSN/K+az1bilw1
4TZ+THPKe515hhxDotCLP7uamMW0tjVFL+IyLtQ14nNB6oB063gReigy/C/nAZRi+tophNx9AVxR
IZEppCYgd7TObPGM27O3ZP9pcY55mUkm4IH7RJ4HRuelmmsrXJtPp+Fqu2y7nJtsUZMqKvXz7wKD
Ceat0wKuzPGK/k0kFqH7YqWbWL43xCKRhb0vIG9juu8eFBrPFCZGmBXFFcdTLwwzaBObX9225Q/D
rWRRIlHj9783ATXw9H7TAqyqnXBMb4rrEDnXcQHsLGAz8TjJ4swx8xoLQ7zjKmM32wK5XIguYDCP
MTG4g2gjnWrEq55sRiwhtusffZq+ODRPDswX7vLrmbm8mhOMCX4xY9DV/vyjtQgdSB4mQmovHx48
IbnPXi30du5U6InMhJ854Gde4zMwFME/bo7GMPkLxmpTHAM4r5q43c0BzTdNVykZwr/GFCLdMz+N
V7uDXDiEGWQggM2Zj3/MFLDMobSpTx3sfkkxfhh9isf2ykFRJ2edbWabzLTV6jg6XX+lBfkK4VGs
DC/7Q090gBcxUnoBYgd6B77IId+1RoN7bga0a4k2JkHnvsMChhNnn2tMlnfBg9Oq42ar4oSPOiSF
VQnozhEjNrzVan7nk0WZ9XzZ3cMbmi0p6h5EL9I1lN/cbBwDQw4lJyIpwxuCn8KmTWdG5VgdE8AR
ZNVSIKiJRZ8twAn340C0gldBh7ObQTNG2hl58mtduMnVFTz9jRnWxzXE7yVNSUNPcxGECvvam01z
taQetAaAZcplmKRkJDCtdtshqKI4dSJXVO6C+hS86tPw0Yl23RqtfgUrzziGpUOzv98Ciq+KsX3V
BYXp2b+0BQ+vK7pSovyM4C651QBZIaysRAfosaKc+aLJBE5oCgCowRHROvUzVhdOBUHu4ZGuGnc8
jgAxnEkDqbFUrkbmVFsLWA1xwKm1qiBvU054pBgZbTRvbpAu3RYkKcw685GQlmzHi/f8O8IAStUG
1i44KQKRB/QcMSH7TcgN98vvu4J/M9JyueOOcB5h7j38W6QRmmN6zAYQky2gzq1RI2lPmc9s2g0f
EAENasp1BiqQBtGNnlyfZeQ+0xZR2T2aWca01BJIM7gH/ZRo0OwhlGoRr6KM37FQu0KmFzqa6oGk
0q1Y8XhU8TRyG9YGwwVsZclMGBp9KnxjTJ1xAnv31fdwZNNT0Ol8CWI7619s9U2uicDB87uibDp3
OHh8DfoDBvsThsXEOKRNue0e1YuYmR0Y+KfzC5PW0hsrnxFD/8bADz9dSUXnSRC/xsc18/gNYj30
jZzzH4TLkO5RN2Ue5QehWJOL3dOeDYKTYy+TbvSaohuXUgTCB6fAbx6i7IzviNwTBtUHua9z7KUC
WcExVxYLV21ArxNo32dTy8ZB8h1WRwLH4KvCKSr4TkJt+NDldt8Fyo/lyN6oLzRmeNIthI2V9xyl
hafxTp4cgQvU3orv4BSaqZNtJ/7KsRH3FoLRRu1XicVnc7uRewFWsPYIPRK8R4m7GiZRtXkL3n2O
MWo3Ui8wUBRykdHHyFHDktjUnDzgZDuEj7bfp1/4F7AeUubwtm8YMg4um5pwfmxe9OzJa1yOnjyS
BAyRTF3Rksz9DNf+HPmcYHzGSbSiNC4qmiEKLGW8NjH2J4bvdeizhHN2L3HT1jJwT5u27GA4Bvyi
TpfPdv+HJ5g1RJpg/dxk0+4njW/uiubFJOpHk/dCO/Q9uhRSLGiExd0aLXqcyUMo+jWgdtLcGdjh
cO/a22Nh5JnoZCt6V2n6D4C/Gki+E/vwtofyig1o9N5zhZBCpcYfQX/gSSK5IZ6Evbb40I/1mqMM
BPnuEhRvMIxbDlWpMGW040q+UfgKBnn8QAvRcY71Js7VoByjLhRatQGAeawUyM/FWsLZjquzOaGM
2z37yGd/H856+wVkJW24sLevDnU1X0HqdPR9gKrZT5gieihGJm7BzZNH00t3XHBrWUty6DFWIa+I
aHvLtbYiCvSwHLCpVBIvzbu/FTP2Pv34JGW9iKu4+eUGksbxLXSu5yDOaOxe4kLEk8/tHcx2par4
nA6pmz/zywe2SeXeEMPlLfF+bwAfpVGK53VnIZo4K6uwH53uqIfRuvV4OvkM1KaAyjaYh84CoZmS
nwGpF7szxpcWW+OkUWvAc6oXkfPSYEqav+bi+kwRkmAu2hA/qLcGtj6e5iPV5KOL/vYA+e06VRqP
empGEJSaHPfoMuFNwT8XKL98KBpPj2PdJHzISONsa5IwYa+UQwzaveU9bbJ1bbCD6AmbuZyVFJJc
+ZlrIx6uqfeKrwAaEcE+eDhHY1bB6s+j6lUZtv207BBniXJGUe4fnchLaQbNPNXtEcwhJEZoSMYc
ft8755bq0mp8rgcUvGi2q44KF+MP7J8wZr8rOhr6JikXWFLCxrZe1I2WAbzCv+sz7fTboPlUmcH1
tPGK0ZywcCYSuhRUQqER9PZDgKDsRvM/ACKaQRFGhiXAFKBw9hLCzEMMmT6zHA+Hom5VBEjYAEHP
DkQCG4m0fAeSAjFHuAQ9//0TEIr+2kmu/eY4dQfHYi0fuDstmnDp32aBVM4D12eGUn1hCdkUItn9
I317tOqol9AzyW2yt9GYfUy8YpeVopgeR6YxA7Ij9rg1RfOtsasuIYpXVfkq6gClFc1Q6FcmWP5g
ZxQYv9A+WQRfwevlnOip8EvdzWeoyGk0zE4uHOrQjcFt8mnBd5lrwytM3Wwl0jGsripdche+4ZIa
pzD5uGlupsdRbQpqfKqNQWshinkMBgfnPcOV07Qud6FYUzorI8axi8iNSvrNsMIvEg5w8JBDUAtX
UWYt93SJ4bdYhNLUUFA4bpIVDNRxDqSGVpRjwEUuZkLB7bpXXcAq3oHxXJ8fu6MSVYlUkG0eje0t
52sqDwhYJ5iOOWfBAXkdJih0Lc3sjhRzW5uphMVWJr2++2uifEbgLcKDlLFi+15X1BeJaRXpWFmJ
s3r0P8Yuf7oyf44OKnDW1NQ1WsvlH2MqIUMHDB0i1C7d30m3tAaV+0RXBVjUdcyhXyDnZDckiiaT
nF15T2zTGSwfYyCvESNpd3uzVjnrjY0o016QDzzTcTmQa03n/zCMCXalWyCWYfrmOgpJ5azQUz2f
noxP9bl8FTSzjISe3y4c9hiUy8i+YsT5yo9lLJTv2JB/QYLDaUvibUPCE3+5IplNgS5neBcOqi5d
TnEb4RtPRtSo4PRko73r9g7U2GBPiBJyGgGTYXg0XwK5rmWzi8bzRTQCie/UEgQoMM7fNdGsWiyt
CHn5XBIzroT8aaQk7LBapcfC4SmOcpPNnZKNKOHwDdeoEdrwxENtJOmzkVYkzS8VSzGg5BajDFuH
u7o+3VGYds0sWMSt/KJdzEcKLJbvlEE8UXBthC1YYFiByfZmza5uOLJwUGoxwwv+k39NNiL1IoaT
1mPJmoDOVt2xwkExAFA+SgwFmCyEWjgNQq1gE4FdNaPm4Bley1nDSqCH61jO/45bP1sptIHe98Hh
bP6SwazWxNGJjeT/Jm+rUt8RohobmBuS5oGlLW+if7pxFUOJJa5PiHfS8fr5mjD4kyo8MhSOLNk9
A6ohT7NPz95V1jtQEIz1bQX2I81EEJQmR5n1aJwtG1Jy4/68ZVmkQ9Dwy0iY+5H2WE2B0YQuPTbA
b8WEkMFlYYiSFBvTi2QmG3JU9WutSBXAi87GpS58c5t2vWQYBRlTrr66hZyf/DzUROH7lgxxe576
I1kjqoPa/FxpmE4NXBZ5dp5xVCL9FeeGRa1xl4R9UogN5uFNCj6drZ7KWOvATiSKE6St/+TJ/Kch
cJ7oH8mXg6erF0b4q3dg5Flk5s8SidBSahXbInEwIN0dZkFtzVUb53+Wag3G02IoyhMjelV7Aflk
ANvYhtHItu+NVudMI94h3oKEJm7jDK9HEva2lGQR5ivZHmuy8JpAWdiXnv1NUTQPIHOEZuRRx6/z
I6a1mLjPSrq6c1fdgElImwZK8zOrqD8WD7FGJTCXs1tJ4vhCuhsoaixuWyyun9o3xZwonMrzv/I7
YG+R+clhTBeMtlmFCIAADujPMVT9W3k0WSECQ5/8fcz669g/JYwWhj13pwva/3dlqfm8bJcbPk9p
FsQhg+I1n4tKdAtTJtKC9c56cGCLXaySfpkV9hravaf87M8/z+2kBvI3J4+wC1/+Ebo6bjPp0RqG
LJMHxKcgeYVjjed6humg3a1jzLuWvSH7Pt7XtsVbMBwP/Bk9KLtJWwViQcDykqGmRw8gyUPWlFPe
uDvckK2YmR6vvKRPG/IJX20VFGA1+lYSubGafgmljui306ihwf2z2AYrY8awt2DVnObgmaeMsvR4
oWFymkdHbJ2keZCEYHiSRjyhQy2Iq1qFL/FOaUjCGJd1Y8ufoTPnEAtpAEKmUjQdRxhCy53E0pAD
niMYsAJefRjb2MGjpARsbGBlXxeqr6WOx2j3uAbUB8ZmHcy0gn/6iXckNop55E2T1AxZwmMsWnTS
mzbJzUsj4wZCSA1C/K9wG4mXLCfajsmIJjcpoYq8bW792m4mctIKiO2u4kEDUu2/OQJFMh1RFyKx
kAeXGW4rrX70WmOgYu8YjTzXr+/DnhF6r2Hk5pBGoaMFw/bWy0kj55/3SgPjjO94jnPfV3jVSZwH
q8BKzW072QtYeGp2lWusnHaFjj6+KKM5zTn8Qb31a4eYTLHxO4K4ft7TuU4sFT8+uEnjpafQAE4h
RvCxS9jJEjIzh/MNNtykKbgoG1sM8CrgivjOXepLD3vSbq7qwq+vYmy7kxf6mg4JhaSCelo+i7lN
15TJv8KDu+2dd52XwXnrFI8al7riG+NAYdcGsp+e7KDJxkK7EXteX4dXw5Els70wTjun+lWiNX/b
JhM4986Sd1Hi2Lqxi+awWqt2iZka6LDSFuop8SC/QmbgKARGO8v1VdR0V9edS9BBwghcOfqXshni
ukXYCNe8w5fe3lbhWQ1D+7oKrWlqVX3JpO3vKaWr9UwghIuKNgWNtv9zZ+YANGd5l6iGTaP92uuS
BngDn9x9HUdUnHucBzVtwKGW5duxVGY5q/rQ4Nelhd9FLcTOyGxqbxtiuTLpt6u4wdn5bJ04GKGJ
hzroGuu7iRsbTaRD+WvqIsw70jsUP3vi2/xfhh9Dvc3k5yXkzVuyAJ8TtJe5YRFH0rLCixUlEGiV
LzkomVYo3yyhIdg3hmtthNiROqApV0bW+5prluoJkxew6z7M/wYWF2YGh4qFOjGmjOxIzKJ1iSa6
QATw4qON3VdqvIj0w6lWM+f1x4q7GqECWHRSq4xQZJUoFa/oXa5rn9xkOlDFGV5b5OOKjiK3egwX
4CKdOZ5zcnJkthQGfRJU8spvHfeupfUwVl7d0vNCaivkj/rsd2GebWkWJO8BYDYcpJcysfkXYcTR
EyZYLBNhNg/4CAgWAdUMNa2KrZ2dxuXJLQnATQ5nlu6tM9IxcdD9eDZ+/ovV+akMatexISpBAEm4
C4PbfZRk5CmBARA8HDYuJZvSu4oI7qdE3QISwwA4nNRr0ZhLGyxDuxWcT4UDl9O0ZiNeePJ91PI5
YPoLIDKjuxT+fQ5FiGMf2tu9/+DUMPnyxu2aE3hFHjKEtvoJPE6x9ur5zdPeFEkXgavY2ziIO8p+
g4V94JOfpma8R8W4fhXsmiSRiHx7TUQec9eGvLluiYrHtLIDr8DIlgOpzox7IYxXCw+ivvnjKX1W
29ZwRC2OYItXjJDGHnHcCpGcf160mUvbFeyQ0TfwzWg3/tZDZ05tyDz9wrlS83WKWTRAKkstHdk6
+CDFzcciJyuefnujsvRuO3y5JWhn0c4Xsgs/u/x/7YyBVeshQLTkMu5S3mGUlkuADXrKN4CcAjok
vV3/WaZQEKd/tuO6oavqTb2aQ70Ikx4YaJmGkQ9Kl+GJd9QGVik7C3Kr6iMa0PfPmvbaFHVmfNwq
zUs37GCr2QqvT4uxII338EVvKCWUCatA/AoZO4XomrBUwwmBhEI+g3CynHsJA1XKVs4Ceu3wsoBm
T0dypJJPzb0mBkwmG5fWn4uFe19OwSNheCSxgpndAl5/dzS3BwSCP1YC0xleYStUDBEPFSSWeDYn
rZURWSD/XPeUDoTz1R2jQPY2AcNi9kYplbBx1IiLotbGVlGyeS7X9PofdlahhhPh0/F+yWONxEPa
XV/EckNfV5cTbiW4REnItxmUEsLF0VHqfF2dQ2lMWU8/DnCaFSwlks3T4lBW54MQRqPzzatcROT1
tRQ+2WTwxMI27HWjauV2kEB4P9G/YkQEKx8SNZ9Y8MRz133irUpb0Og35aNMi1xOohRD6Gum1Vb+
LLKrDhpvn4n5myxeCzTxjjg8IfJIu/JID6oWQWJikUoYSn+vWP24XSI9rI/XlQhWkamybB6uJV52
nllzLcTmXFRZfTeFMKDmFo+B/zMtwdG2pse1l2016Q/H9KBcaaNiKgUhww/czEkGRLZehMYc6Ye0
xdosCGUzfUwD31mDV//z9RfnG4/TsrfEz8ypm4+lNk7mM2iBdto+Bx0wWi+J3QX9PbVt6rr7EmhY
ikIUxDvlxIcKm/c=
`protect end_protected
