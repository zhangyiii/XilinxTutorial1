`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 41056)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMKRcNvzOG7grs/8lZMh3KNjoyD
IXsq0a+K7fwBVl18ZhZ77ZR2ufYNrrwZIVkd/QxkLrHGdxRxCTNZj6M3fyHnaq/Ru/ylm+kMDygR
Ah2Y9WU+WUyGFbSZagYIJy11YfkZHmgbIAJOWa+bcgBPbwIWz3Pj1bqPKZrtPKht4ETfRz82IeAJ
EC49c/ERJE5N5nAWt/8vRyIfpja8CdO+oiWkMVtHwvVFeGwDBBgSbrPQkP1hNfEvVk3sjlpj6vDi
USIp8iGha7zzNGDNpOCJrCwTyACE1/9DcmEeri/jqT1gtk2oKhondpRBmaje5Ev/jzM+18bdwdPI
ommNf7VxHyOpRrbfTiWrwzlFzaORsL29oabiSQvq0Bf8ffsHaAGtOieX+wzIZRxCCnEWAKfnltLi
eLTjKJCdQ6igsemy05wKPbgGpASiN1IL2T5h8ka+ivcdel+LIT/rTDzQL58QZHdhsvmGxqopyjLk
3Szg83AgnQwRBOCAuMu1SFozfeH7b8mOiDHT8j9RBsWhPiyiDHVPZlKVBF3Scl1NR19LVc6Vyswv
isAsvIIzwyLex5eb7e9eX5kxflEru58WgVx0DFgCfpYpGHi9obXtbrSchHg92Whs9JRTkIsW/mxx
wu+tUvYvPlPgZgPg8RPCdzcEO9IdzlnBFnY0r6J833jX6chPn9r+yoi13SkEESXrhMeGHtAywF9M
GiBZNcx0m6MKaHTVfLrYqwCSksFIVxkcu2zcBM8VihU88GsGEwq7Rzqe84EwPa7pAvxjzImvIVDM
eG9FNDJkuNsuPcY2mfBelcP5LBz64kVtH9K/2BntUxYo6DY+YJ5IyzzxccXwuZwyAPqwYK3M1RTa
9byg6IwDCnkOPNgyl0nkVjDWViLXkmfexoBl8je8+mVS5nlSx59HuYBffzeTnuRWb1MyqX7VGJg0
AyKBig7efIjVisvryJFBU8m5uANW+OxftbIMrmoTAX1qaGL0/ESeSPpe+TWSc0KmAGSxvzizQD2W
xGgrN9zHTHBAa2wl3nJE6BMAkGGaTaasjINILghJaMcf19m54yE8kCT2kArpUPSUR34Pw9P339Bs
WtOYIHCWF9wfh3Q1ITLWxSslui2CHmjO/7HI0XAXfww13rFvK6qBh2o1vuRsfSczfXLfgv1Q6IDW
kU/L4kMdlQNhrXEfX+Zj0WKwnlm6DxAwEoKX3muuCZtuAKZEpkRRiMtLAwzIYYqGwjWQqwJmpUqw
BBadDQJ2qg5HCgqzt9UGMmlB1b9Rtbxv2rdP1GXNzOzjHHQFbx5Xr323MLOHrl6pQjy3IDfLXBzp
PfJiL8q8Vgpty/a4gu9RjRRXODmLt4i/99jlqnXR4ImGF34zAV+JyxwoqrVqyrwHMm93SdBGrnJ9
LZjBRms7x50HpUdVGOKHCdvbXt8V+duIb353o5V2BAvr92b8keEWIwNHdl9NgF00O57h1pcTk/l7
xJgiz2NyQLXZRMBhZ/T6/tP0ofoRNK8bwoz7j5d43qnGdqhm+7IZfRFMySqqKwnf7yQDmk4E32+5
M5sKclnDBZu19WXJiHUJwdrmTgxCjvbUSgxjY9Enwzsm7SmcyHIG3PbzDaitEZco7C0i2X/OS4wm
dx/uMDtmpUBCfaLJ+M98J75TaEImFHLATtEDFP+wIqARUCcGIrnK95ee3X3OpOI27KYqJT5RS2xd
kp8zuOUI+zYkc6HjR8L76KuzaYUsPVLb2MY8xDbAcx2KphUKAN8fyMU98WjaVefOuNr5t415Jenp
ZqUdTuc+5//ZDOsaff/7CKlraW8kzh19uyDM5Hv32n/hpq/VpxeEjLHUKqhQEDjyZjpk+/GBuzO7
qxoGW61meIeW9k18uUjHih76rXQ9FTwC9fgCgzreGd/40TDtpwyEIhO3FH8lndXVjdzqDhdmM8en
J8JICMOWlNzpst0ekxnxHasBmU6uhFHpbb/BtqYl0bX6+gPk97M1prs1HcWP+qc0AuxehIe3uJI8
00/5hoxgEfJMQz5FnxL673EO1yQXfRuVqH4oVtDVR0runmCg9qQVZVHdqNz5uoPx7SjTDRhfmG7v
n1PpB5pJ8k9X9Kvf0GHNUFjQnphhX7Mx9zDTy5hTCjitt1wlzb6CGKklDPW5+abWFaHsvU1wAyPu
siVPCipdh40uQMW39vblsv6t7tT0ny/y3r8F/+fia19owWn+o+S9FXDcdxuhc8WJtpyTUDL5dcc8
yzSsUfdMBbkuDVYRSg8ELjFfEbrdshz51U0TZjf+kQELqAtmh1Ou3gx0Ypo4xKGsycaXBR+Gv4Oa
1mnTptY7PJ+y04TDjsDM3bdAWiVFvAbdJuzjs/9gy2I4ZTbLWWeFGPiHZ80LJlnyxL8nTcwS8AUv
3hM7VH17dIqlMRVAl/jMZJklVFwrc+qerGyfcAW3S6ULk5s9er+VvS0+ohPukeVYN0/P5NGtrBn0
24PvF3NG7S8wA7TKbjw/Zu5WLViktzIy21pfJOLrpO/tAjSDPM/KggsviA7ZAJZuRdJwbY86b/am
46nHz0VwhSIJHPJFwG+dhB0lMSJCvc3PUvneKrMAA93o8x4lI4CXdatQ0BNDT4dlANLy2KsYZNy6
Pc3voRSxWUL+b2FjzqAKi9BCCEPP8f9PLWDdxa1QfdJsNbffo/zm5V3x9YWsScZY9rCj4pI0oHd2
NwtxUFN3FVNqQ6fHyIbJRWvcNvSJGjc9sjbK/+ehi42xIRlS0ViWGyoSJP2diqsAVqGrAdznzEjH
Uir2T946hvOuExvyafzJxXNu1ubAGGJpwW7AdTO2y3jdTO0EBFfQVb1Vyv8kaihz9cnNUx234066
HRQnuTzSrmZYk3HaApOtKyZFJuj834WDftJgCjsnLC/lHtev/exFc9I9+N8rztL8G+qQeksDeMmN
jO2OEaqNycuu4v4CMZVvPJyIphVP69txpIbtNJP+npnTNNbGqUhvTAefzFzS8WB0g9SjqF+G8WSI
zgIYwzLRuugc1MF+/B2r8Ml/iGqdWoxDJEo85X6v1XnlAkBp08il/3O2HXc5nyqBMKNkdrR0yXjW
CkpHKSBpJxEWBWk/reTcP0olBlcQuk5ZdAIGTmNOH5fjC2bivjHdrGHKRoKRt92aHrVKpDOLHZ5Z
x10MJfSOPfJ3nnoAdK50gtrEFDUmEqdWfm3akqKn/PagyDDNfzY06n5QAXm4a//w1Y107/+t1njB
FZjkxTCHSAr5NzVB8dVVKZdcuuk44nPSczNqLKHTbjOAr0LoO3vc1YbC1qW5emuM4yuI9PrAIylP
ShGHL9WYn28d++lkMmUX8cdFm1EMm6a2buvNLVw7wPgX32iNZv0vY3V2kw/lgu71PTHpIy7auOzI
YV80wNWtmL+L18Q5BrZO4vqDqxUK9rOvJiVSRMvdrS5pGF7zzF/TpHGwJk1dunr8eo1mo5xtUtjb
IWQISzkspfTtkBqZF9nmxbat4XMw/kYLz1hpXHFGjMwO/KJ4PR9M+rGHCRCN0VOYEd0QIRlzgpHS
3m2qNPueOqlSTs2o+YMzFjw246VIWoqvb0bdh1vEidcYsksbsoKYKKfw0ZwTWztBb/TnFXqQ0qMN
x0U0arsryEyUGCipJ0ihZU0WgfRPcuDJVdKBAfvsxWsiu7s/NTcWj0n3zLJLxRwr1oteho9RJTVy
sN8j3leucFcvv7wWANLnesJvGpXoVqvRSSrDhkmKL2KR1clOEEBNI6FsAsS0siGjP8FOIxhOCWOt
UmL/3RsxHzNqt0d/oCkJS4ExffmkNjpyTYfEMpjljiWCPBdecElllaF+9y+kSeafsNV4EVWTPTg+
L5mM7v7zLtxktR6JSqwfPWLc7+ikd7mMXivScLUVHJsCJPk2uqnc88z9ZfXgc+PQ8SFiwam/eNKt
6mMnrMD/1heInidlcGLJyw7inpXE5CYXQhNA9mo3MHdh/RKFEqBnOOJ+viz7uAKJOqKSfbnm6PJ7
jiIpI+Olc64fFsL1TBrQA/1qX/0+Km3gqO/aldregRaC8uFaT1QlPbaVlIVchAhSuUibA5UJoscb
LnnJjh/CbcGItBWhSHN87qpCqi9GBsQDU1sLyuY3TY3HSGrOjJ4WwZh7WUrRVnwZW7ePvRWe7vBe
Me4hjTaHeF37DzBvzaUDMcbJMBg/UQKj4CHloRkbCr4v1XRdGUYTe88LyccGs0xsXfhlbrDTmaQ3
u4HEsf7bjzKiQxTRVBtBR+QoC/xVEqLYieKfebMnOLSDG0x6SFYtBGaZji73sE5cJYe8kDRf7FQ8
8ObvNNtOPxRyzMOV3fudzqTXBW1Qi9SjkG73hEDXvdJwLMVW25OJJ3EljP9OophFBZy9/5jN5UEx
fHPbtnI8Ktsr0wtSyshcMJIXH9lOCjaiTW2cVxnV71wNSDuqnAgi+q3vFtH5KYtFwLzPBMFLjsj9
m7CRM/DUCmaXziY0KEGsZx9Uz71DXdV/xR8HRd28/Htr1oOxkjXQqliXyZef16cQnpcG09iAPMjp
P7EtmSzh/dLtvjdihh3s4iGTiKCHknA8727uKfnAeY1X1ERFewA5vktLLwo/521K2gQlJspQkXJw
9Uf1rK18sU7mSvu1ctamLxzrpgXlNQvFN51evP7zUKFfR4nEWYTkzsK+1dZguzv/vjrmsVKwiOfr
CA2+7eXjwBqtQp29iLeiyvFTIBBKsQu6dj8oQcwqS8mZoucpATP7slggKWakEqlFVBKaQOSxRuHv
Y58yBTFomW91dKXAhnaEcSyoVMgzdw1Lk/QeyjRGVpP89zQQkzpzDAOsvHWb9qiiiz1Q6fE7178h
bXCvwsXsnayeJPttXkdPj0QN0iovcaGVvECOo9wQ4sdgWWAM0F5diU8fzQB1ZlLowcE/HcMrOvxR
6Ta69JO0hbhCUtbCubu6IuPFjBgc90S0LEWP2V79q0BYiDB3AlozwX8aMmyPbhX3FwsJsDVTyfM0
qua2F972ehtPEcSJtKFed7cQCAdwWmZKIOV09/D9xCbPGGDDxzG6NsXymStg2Ey4FB3JvOr3Kivw
kdBiN0H2UySm387YS6FnxD58O++llEIaYl9uqmBESXJEou9gf7JskFUrxDcnncq7eul3fCZjdcwz
fr+bMu8r0PdGcUFwghUMyVIi1cWUwO/1v4j4Teok/yiRt6+AyPLB27hJJ7MmMRpiDj+D2r3odY7W
Y4DCUqqs4YTCQgQPC8A3HPfIEDFi/y14XW40qiITMwwaknLGLbDkX//E3crndyrH8aFIu1oiwJaC
pfWQnSNXzIRI4iPLsIRVhmwYeGIDtrbmqOLmyaTCVgkD6UvfoceVYPMSlDvbuEewiH5ajr/mXd24
fpZ8I1nJQRShvPSlXHsVIlQNVrCrhBEJdTIGZm8p06CmEziC0rESbkXu1bT/nG55Qp+V5g1mW/mf
tVGlQ576+lgqdEMZFeF87DdfNbAIFcNnAVjPWK0UGEw6JyYH0t3chBFy3p9GpJC9C6dizNaiQLrp
HFiKAYPWab8ntstMRUFZkU13lFQzV6IUeKXgwuEylQbFJ6BIs1x1lFGbsSriZLiu/bbPyBfxzGau
dsypj9Tg0nu1jNN3sl3Zsb8JBnlT0bCq4aTmvyM7qvA5DcVx85hQ4WlIKTfQkmVqj4nbfrFzllvw
PRU0Orgr9SQvVXQqrvau4+c/bkAfA+AIqWk/7ZLpOTRsoDou+arcmDJ7LyzNs09A32j2p0ShgpyF
6mhxYBV6BN6NnlRR0Bs1RFXIhsaP9VpL06ixc/tsCHOB8VK9XK1GLdHPpXhhg29Kuml1cCFwllY9
NYTQdaqz3ygH1p2DiIkhxYyC+F34OXspZXmrn7750zBt004zD2nzioiBhWjHHF1YSFruYM2BFkQt
z2nzUKMFjTycypOBmL18WjrdaqFln7Pei6wPHfmqk9DbNqXFPjBCD6qIaZHfpevXLQ6OD6OppXDB
uGIhpkBXxEQ9hb+AyMnyc9O07E+zQNgIy81m9BOgVqiQ7WxRs2UnWHVIyqWD8xr1DzZJj7EeIB/A
0S7nLIpE0KUNW5u0zjPijmAFHyYlJrDdPz/K+QdfYxgdf/xRyXN2m9iTxSj8MhJ3Q7FVwVWhpXHG
cpZW7m5bZfhR44T5k6xaUk/A2AtzlgKkMx1TspLY9n/7LVbEx5pr1y7bIy2u935QJC5WPcXX1ujF
VHPo3hh+762dvl28En9JV20upvVX5X14+QnLImRyIlcGcEdjoXpTwfLOS2igi8aEpqMfFm6nMpHB
6NcegdoLuwBeSYsPQIsTj8LSLNu/PHJW309e4iKX3vEvAbwjIa0IQSFvseb6Yq1elOSl89sZO1Qr
vsA98WL0w8LfnMqZCcuDZhzAMcvXefhf2kXbJqjduMB75sPM1NUhCcV67UwOeXV+sq9piQGJ16qL
Ecn2Xjb1KeniNAtInNixFIOC+mz3UsbpbOMcPBfnacMPerzP7v6VSb1N11XPS/3sZpe7xe4iBUlx
804AEEufyq5dhEKGY9DKuexeLH2hUyl43+5Irf9KWYv3u+N50Cpm2c4mPAgVjuhoj5qKXKHCggCh
bzOtGxo+mpYPEGwmAWrGaI0DIMaxQnvRloE3n2bAVdqEV6PJ6+xe4/oEgRWX3G+v7i6yF6VjunRg
FXVvjS1W/3HnBsqg2RK0EFPJ2mDsLl2vjKWjadLNj/q/v3zKCbxcIibyyBIK+Q8yPrjz2yUL4l/9
njuvx/RTguxMaxnNZFr+WsS6ZBzhQuTAubmXMJ9+OVFrisvx8Z/1RewEZRy1rT3OIapC/9tpYx9w
FLOe1Gemx2HImZlMADx97XBjTIMxj/FEMLO6fY/yMKotsDBNteCjGL8FeXi4KVe1NvJnhkyQOlj2
VbwJWLuIGv60HtkCMxOPfHVQ6NfCSnQ97P/MejAEA40uJjITRl/HQd+9CqMe416+OX13+/xwcZNP
IbmxAT0dI/TzZcHys/ob91Nzg6EU2UzKWuVafOgHhrCNei7XNpO9KTAIpTaxUm2hnp++NanwQFfX
DUbZ1wph3xd8QqWxDgKDhdJnfwUiMO6W90njq2plHY50YdqLlq9DoB5VIrpUYIEwG2+Uwl/qx4Oi
raQ8KtX6XkrMLNq7qawIU6xsuP60kLk4ywiINA8F94Scup3qMfYn1ehkc48s0X1qelY5vmbtyRNK
5+2ZK+exg6JfpW9HsaRqV3WgT7HxAfjxP5ZCX+eQ/ndDlnjojMRbVoI00OkCl2H3iP2CTH6ro8WJ
Gq419G6DZHwMlPVREaAsx+H98W4sIODJyl+/UkFywP3qTmNG0Y7lg4BEdLR6D3LRjvMEJFjn/i2E
A3XjNOq1Twfq6FPgVN8az/+qCkOShOtNn1Bbstbv02PD0hj9kHlKef3+UUGn6yZ2SERm3uz+1q6q
oZnFiAnRZGe9tnfjhxXxMCq3g+GYIpP0Q5THStzPJ0BuYRprcvIXshE0iNORp/NL2EiM4Iey+7lI
DC2BqDiKkHh58rMiRmmR7NAI0K5Pog2aiHWWygBIw6daF5KDFikEATnUlGvJDsbrebP1L64BZSx0
ZlVRlL9oEHfPu/bIAy+Qw/+0GjkMEUsJzco2AtAvGjpPs+2m/T2DV/yJovCRV4S3jXV0kakaBv3+
NhNxnTnOObnPuYxLOn7SJX4FyuyaWUyb0O5kDRvDd2aU/1OTsSAMae4ukMDa6QmfjGmgaosZw5KO
+iO3yAH9M0DQOhryS+f4XgBKoIxRO2ZvgPSPTUFiMR07NMbpzz/6IdARgtP4uxnUz7V295U50KMG
zoorFUzvla4S2IpxEHyPCusZ/yfnhFXxUbFAC8XUKNzKDmvh9lSQNsPEOEI/wFflKTg7V2+hDoTH
cBXxj2q4DAffuh+Kn8HhK/9FAg6IAHrIlANLut5ZaFNQchJNyxaPpARK9HZviAzPpOjTHuKxg+/Y
SoUqlZCy/vzFX9LVxzFtQf9obGbzvnMWS5i4QL7OyChCOwM6tmSvdmYiv3Q4ug0QcsnGaN+mnCq4
j/ujuaWvtEJojtUneSi6TqYhPXSqtSuhEtHkEfeD5N733M9CqSuI5HvX4u8iljKtZyt9QkEzTGyk
EHSIW6SfKt4BpsGMGLNm4dBXoSQjZN4GL2RccblZKVsB93QkJ/Q6ULubUiDUSkVq6BIRzlBF933I
31d494U4zJ0sDGsjvNwIt+XIS7U/y1ljffu3AXpYrFZNQ7W8XKKiSbhTyKBZgXtGoO+n2oF/VAOD
MwOtvVgs3NaGnuIQZ1IUrZg3QTUxXyPukCkAacxtcoCuEnV9D+G8zwtzEpd3vAG6KL8H+5KqyDoZ
HwZ9G9e0bJV4OXfqgOSGwHrtiidq+4RsQV87Nzdm2Dy40srWEE5DTYW1AVgfjxtRgh9O/AWCScVu
yVTpzIleIsEcp2RiLa/J/MTP0AS86r0V1vAZV1h5sOZU/0it+BV8/idAaHqLh2SMH7GYVYu9bXWn
RxMgYlj42ReUuh6++pw5iglZm2WJTiRNpEwq59/t+bPVdDctGT6S9vK3iFQH73xUDwPDHAiBivEe
2CAwHjJpN9QutMvhVaom7mQqlgyy2R4Ds20obZdkZK8Z9AISyknQGlULJ9ktUKUIY9W1s1vEDZgI
/kY7jS3y2LxGjPH1IxicKvOFeJPzVNDOkX13+cnnw1DkOOUevn0YaCmxHp5OsscuZRt001HMNx4J
SWd7UMQX+ySauRUh4JZb5Vk3HmVsPt4wmG+YTXvDqpt1o8jO+1UVgrYYDd+zAXnBqEwyZD+IE/Fe
AEdXa5lZJTDOvFYEXZ8EAksO4lcz+yTXc5RRYhV5essuOVqtoVS0UKmZppqPyyjwc1gEDvpbE+SE
0JafBSzQXyfemL6kGkgE42PzVKtodzXRluHudwXIgRSGzr+9tj0R1VhMHFMMnKbYm9qDxX9I8i3W
lLIZ9ycEWzHLGeGMhHXpClJn6AkFCn1FQG9uHBuuQwrB9bi0mUiyCq5G7hC1gbSuhA2rqUcfBtB0
41++YFT0smowdjB1uDsNrsummNXybk7wGTi0f9bvu2MuOfQrS8XFyVruirvUsmC9xDPkqgz6ilTX
VDm+4VQFvBrYIGbN7iRHxwmh/OmYe9+yJMcYrZudpH5nMw50bFLdLZ/n2daEjL2w7NP0MUswNxyD
lqxyPS+qOqbfiavMbw77F9pOBRjcO2JLCVs7uW82eip6D/Tm8YFrGOLSyyu/cE/acZo2AOkz3Cpd
rFRzAFKTUyl9cyrWJBWqANnLsp6js+JSyj0yzYmsgivD2aUv/QtlgFuYiDLTX9UMb3J4brLyzzWR
pUs20N3Q5Vw6q+ww4jJn1vBbKXH/taKS7ipdTCfVnRD0tQPY5ouK+YPCKX+W1Y0MFD7BuwJOOPVX
dBf5EPSqypjqrZx09+11lVQd0t4hAY4bNYMpLlgviNfJejXs/S+P4Mp+O2xGd6+6gT6mL4I0Ev14
DIO1RNfMmfYTzWAE5xwTGN8LeMapfKv6Cszf8up0uJNM29K44/EIKmY7GQxBQvwBHWhIZgW3lLXR
0z1/QGMzJ940Y8+N6mRFNoIR+BhcnZnQyWQIcQAgi8CVeJG+3JT1m10ngQ5miHp2PEN1ITcqa7/2
V5QqHE8eQjSBVfPxLCijNgI1Wqvb6ty8HvZ8F7CIh0I6M9A6PCQMx2bLZSkcEuOJRXsJmOufYP5A
yhk+33juy1IjGmXtrIQbYJofImTNJuIfZMmd75b3YAGE7MEct5Kk0CSIw7BEGL3+e4IproZacCLf
dHPyI4s5CZt1idsqvSHIn8gTHtgvmxBqoyrIDp67L5yb0XG/uth1DirVODlblggqkCnBfhhvZ7Ds
hkdZ/9HzVlz4BtRFTye9qkjiCrIBGM4LjoRapONsDKRhApxG4fkGzWP9z2rJ2KvK48qmmh8vCDDx
AoN7KzqN+bhKoTctbUV1ruOlu+4P1h5pqRO6U1XybDWbbVdNFQ42c5I5lBx89/z/I5FDN4KBaztm
IFo2JHg1OOi6UYpKUmtRxy5nOy3Y/A1zIap+ZYgpUAvd1jAbC6n7X6vk0hgjRsgZldcP0hLJwCj1
Xa/2beDCzaTbQSU0YJgZ22qo3DQ5KvT0GuZNZZinTPJdTXzejXYgS0XFowXS7Va4yot85A6f+84d
5LQOQlFc5vYcX2xm7GGk2Y6RdvgGaJkL23ET1KjAWiWgBc1eaWarcsQ4BQoFbLWzwElpxFLvzBvk
h1c6MUnkbRnXCIwNlks+0cfCFVT3K1zhPCxd8rWxhxbuxJFA33cOpr5GjiJNcso+KtnnYWB0ZpyB
6aquGDb0tAtMunwg+oDEohETmn4Ph4stb2ul+v6DUpyI34/9Sfok+QAcRtM0mRRiPOfmy/MS6LVE
wY2GSZfP06uR3M5ASBMhewGjPDT+NI7f4ZxhOTr+tt4LHaoU707djGTFJcLInyOoT0hX/1IfQthW
F1gNZ0sj723myRWVWTPpzA31K7dFazVFfcvQ1cj46g2qvnWE2qzHTEBSbOMqPs2SbEqUu7uEjA1m
VAA5UiaMKjiUzgCD0AFvoW/DHYMwHpu2bh6izjSScph0zxvJzzndkQH6RwCqvNNxWXAj4pLrDBLd
v1FjOdqW+upUCdUVW0ApjLMFXsKYIxGyh1KKkA+Zpi4BK9igsm2zT986hLYG/ioJbaKKK8n8cHyR
vyQMe8gYn7UrbIkMq4ybnG+rTIHM4PLRsdIBvxt6BggULi7P3ArQb6BRzyA/bbmiwU0B6mJ1z0uI
QQJlEGeK79ttQdLGbA0Ogf6TfP70am3iI47I5od9HYLUKVheCFW2XVU4Ts/3RI2pYz0QNYx076rf
qOczO5RVSC6AmPMgEPKciQj2HP/pxi/i037Hj4DqXVUoAuaKSotzPkUcfTmsc8qUbaoVPvLkHtLx
YW4hI2/0UxBRnN9h5PrkaFTPRzwQfgMNmoEGWKQnVw6xiayD+O3tccUJbbCQWuJfsK+iJ9/ohWvX
aJzIiFhbrItPHPeZfmRESYAGRNuPPjdZYX7UKABZtce1pesujJTSw9ZoopDQuVMMyk/Ox6lYSvvZ
yEmkK0rWD2kwRfrCmJ2gkPOJhAdb4wuOTXrwed7d90wQ4rCwuikBhZYjXLXZAsNEpkdA7zslxzEl
ml8CZ+uYG1jnNnRTHWUvBO0XzkHJGrh4fDudPpi6eYXvyLkKGtnujq7DADZncgF5i02AOuBsmHPl
0p9kfZx9Vz/+34z68YU3oc/gB4v34sAh2L+oGJEjKHdbaQEM0zqBOL2dRVV1AH6kpPdaVQRVNLnO
Sggd/pjBoelScFCREskNyuSZxFNspPaYi0+wLZhbrxFTZEofZnfrByJNb7mxy09huB0cO8mSLB3G
e5K/skY2Gx8E9R86eM2vW+dABFPSH99nO0GUildKQFTZPJnS0Ya3ayzsJy6MPRa+Xcw0xAwiGQhl
z6JrsZfo1NQHJSR4sC35ycCZRpwiBpNSvf20jnG4V/EuBZ2lmyPrt5YRv9zvJ8ONO35yIEYO7Yer
FJBQPz0o/Dc86l7G+m6/fVMbpLZEzl/H9THRPwSWf1oEwFInsCcPtzkvXjOhMlESO/bJEQ2YyWm3
BonvOHAWp40BmzoiBpptfr5bU9emYyiowdPPTLtClBvPmvUaBQGAXQDmGN7HMDT+6emhZDizkgnE
fF2WpiIlg/qkl9LBkMSQVgF0dWbWy6/InD2yy0M3s8mJ/8b5nP7L5cgaJ3hY58DD52b362ponB9f
vll1QS0jqwGnLX2KxTzuaw+wOBri8E1MS0VSvOObn+WXT5MI2CmRPHWRuUF1uUJLVoK9jFpFS7Ei
bYb7+Yv0BGvnrLstvzUjWr2BObJYtlf/owrBtEXI0uXbmia8DhuV2LNNoRQ9y3wVvYXcvRGgOtrW
WyZUmzlJr+g/9ak9LS+G51xbra31p4+eSUbguTKQ6VORbOWDtDnyWgkYayFTSQjsinCetq1/Hh69
vUDWME3YXCGOXrDJANlfhtPY+qo0G8erA1wqRIMyl7XoJ5U1mld3i8sr9IWMAx3wMiNxDQFJgPtu
l8dM2QAp++fc4e72I6r8DaoXufFI345pAQMsq0oi+VvBXombLxSbVeUjKcd20E+naEjo0MNuTIMs
Pd0sTlhxOVsl2tApH0f1J7Xol3t7N6ypndb16xKyjQKpfRf5Ej32E6i+iIBexx7tnGmMJZ854ysz
1MR/kmtIsMTM+xfvbvjfVfadHON28mBE9juuchKWA3IDUiZXuj3ywmrpZuRf6rXWBtii5YiNaXCb
NzghSzHwPFLHmS0Kh9e22lNv2OCZb3YzX1TZjB+hkAmEdY7VF7H4p7/QeJpyzl4wK5yxfwgCiqLS
yWxU3Yk3RIK0dd30g8hzxmmGZmm/gQ+idIdMmVZUShmJgR78C9oO3oV6Ley5ZCqcAjDbhanb7mNr
1By2Sz66wCNihzo7z1oNbgEz7oMNv+LwxohZ1yJvIjRdC/SdtdUiM8ib+DFT4tV68vjR6J/VGd9D
uwNtnO4D2o0rZId9yrM6H6MM7dmBIE3jbgr0vI/1aqZMJRqSI2h7hC6qLUqlarpoid6/6FlsAEcJ
T/v4wgcWKAGkQgKRULj5pgibecbMYJzcNBeAoaJ+UWXPm8byEDpSsTuqRr5C7cGf6Rvb+C0Bq3Fh
S9zfnAZwaVAFZHubilZbKpCUMWJPGK++eGY8e8BAvma2J5RVzNjj8OEP5I8PGMHmZpL7F4wtGENo
u80cWFHhe6yOqmSe0JaAqmr8swk/i1fjfxMMMjBL2WKYESbhtj9OUG60Majeh8gg0jxWZ7Mw4n6o
6uu2pWEuF8+sDtzw3kpDdorNftoh5Npm4Vv7/U8/9Z4DC3ei6UK/V4I4BLVpcksrDwEx2HYdazz8
n3Vcd3JLh3sYOTIecdJBErjShLVn39L172kiqtc6pqJjpCRzLkSfUbhMbnKefa6MvtheeWY8c8Ug
KueykOgV3iZNxfBWTialUK41cKbVl3sobw/LP3pGlltqQevFVV8Skbr9GlJB0OfZFjKqazF1L0PX
k31y/pbCoMzvEVWoMYXyKUakg79Nc5oH1dKiOlzXnGfD5H2w+wHR0HDdw0CpW8mOrLfX2eYGlXfo
8SMb/0BXBFERz/h8q7mrMvzAep4b2tdeLIAX6w6/X5B39DJ/wFj6hiKYLH3K7ZnYyXjrnDn8cyjy
q6eyRM12g1ysFjQBq+7JARlLCyx31Uw5nvmZl+usWObGK3odSeg9NEN3o2vJrxJZgQ0O9MiRYpra
q5t5XCBJ3+79p0gKMcENVKm8HpM6LFjfWOihP9Gyo64/W3H89gePgLxNQizy7Mfs9EHG68u19qAA
wVQcUEAwo9085Czoz5SBtDDvTR+Lgj66GZ0J4dKm9Qv4oCmcOGfBdohExiA1L+7m8WEBkYVLmAKE
cKI82kTDkO0eOMGZ0rtcMwFJkI9W0ibRdwPdjaHk2hVYEXTKvbTp2B6pbE2fhnXoGRnPyrF83DAB
SXBFHZdunNdVyCmbC3s6DzFdxOVkEESG3OurGzxq9GS7sg5Y3tLQxnOdDNlwRGGi3eooKUk0QOt1
qpSfFY76NKl7gPfBb8tIxOIfX9oi+vvWlb/mJPz6rMSz0hApq31hpCUd9ZkqVkPIt2pvLtuXRDi7
gIlO+fLj5fHulgBMfrq4CBcviYVn3ZTTdkBJ4lKv5qzteVofvT57XWTLKvKL8fIPailrvYqrM2g1
OJeFUMta+D2yia1Rz16PSSjECC8Su0EA2hzeSmSLd+CKeL1FFv0nLZESzGNTCPx1+CeS8wtMaXyQ
bq/0/ZNOxhfzmYb3fj1FPs1qMcggbPzEpXU7PPBk39RTTQ69KEtVzC29rnRNU9mp7x//DHUT6+E0
6WTDbgUa+ST/Nx2a4OIBv6ZKOX24hWFaX9Vn5YskVos1q5uSj8uEuv9GTMLELdE2qiElsHtkgGII
5RAY/kFVKVGWdSJMCD+Vuno9swazrbnNGmjGiYYt5XdfjKyOn6XpafI9WZbzzDQzPOnG0dPj4KcL
rb+2wbxVPirh+XHljHLJIQM3PQ0QhkE0vXNKyznldz4kzM5R1sPW6FrG4aQ3xVHBFP2NdXVl1TjY
xT5UnPKHwGOMeI6yy73dxdXyAkwcmbGvaWFXDp7RapFSC3I6XUG4PLYHetr1dYL+pMUzMOnfdzVE
15+cH9vgjzEwW51ffsmADr/MkLEqimyiq/c65K5JqQeKjpj9s/4KxqvVv63BFUuDaZbNey70tScA
T37pxoITOXH8udmnjt7lAMoly7vafyPNRpIoXHaSJzQAbfFPt4h6rxC322i1YbIzZ5rFX4JP/yMJ
LnczbjsaeUBV28FIIjMeZnKECsFk4ZdG0Cd2XG9mDtsMw85ryQJTNp3qL1oEoMpOrGIptkloA9EJ
jOc8fXiQp3n/PNDSR1Jou41WTQiRtdRdvfWkou4RSW2j2G3UL1IWDQTaYGdB7+iqKhwDGpEzjGqI
lpd6Wm+HGKVozOFCQrqf0VGNKDyu+tjUB6PbZzHk77NjkInQTU19McMh/xq9wIId0uJauKu3aQN+
fSyouPTEMN5UnfnL38TeIoTET8vNgLTdg4JjcBxOW+uB5SOvZjdDmLe6j5m9AbtjAlqqj0XnxFWy
3HRTT8O00yJqyBmvxK2dYLEMhzAQhCil0y3UT6MQkPJGjnBNRcccjxN+ejGEFKl+NWXftu65TL64
L/uBpLJYNBdJWUJwaM59xRQejsGY6TEadOU1HteeR1YLjWEirv6ikJZLYUZEtKtKDs0Dg9p6whDJ
AGOTC0xzxM1YI1ktSsaGjzG6kxbyXa1qmcNNYSMsXyT1ejSkpNWaZgmbPgLeP0ZJrLhfmSLx41bA
WddPr+GiduCFnoAf/0Vf/SgqdBvVGuXI6eu0QUjPAGc3yicVAXzQ6Dd0jEc/444RNbDRi4Ujt+cv
iWKsTmJG1cSd8g1L2xkmZsD7ttJgb2YjzTi5a3V/Ihm3fNQiIqkmp4N6NvFl4zRad6YV3F1QnMgD
IGb09AJKxLrGDadQHASBHpEz7kkNzmZOhil9xwvYyMxR/wySy7dRfKAOd89DS9t0K26uvRzjg1XZ
+TQMKkThDWwUNhJ8Z3jGBtSjvNnig68lifI8Sua06JBzmneWLLTIKg/fxj2XADe+X0bc+GWSWVDJ
NoWvU8S0HToE3aiRtMJkHZ5uYrYglPnYs5Fqf8avc3M9EtItpFxeCO17pD4PaTNZwmOFF0QHZgxE
r4acdVB/3uRUMu/sBNVRH4m8aSy2sbh8qdLed4Fa5+O5F2zPMkiWGh/kBXDqCRm/LWROEoFWfcIK
xHzicMSHqyRA5iTaW/PbB1Fc1FS8MqkgfvaP0/McuScHz+9a4MOYkTUCVfsnzLikN1cuD1Xbraia
qzcDsGJrXTHz6/BFd9S9/2IcdUv9RJQ8oiXvKxVKPZpfhZvfBkawWdA52qm96WxgRoc+U8wcxjAh
RNe9yYAHSUABxtHP1eB8yiiwQT4NBl0KMImjQGzYc2NoX/8H1szxCDDLT8/3n2tWLcX++bd7Ym2Z
8I/7+p/HTxA7WVINCXEIEy3JoOmr6JtJBNmEIn5jbq+k/YceEiC0LnfsrK8vtYQbuyc0lVPGJ0aO
XhTEqfiI3XSNPZ6lDTaQVyRQULQu43zAeoueb0N4P3qydOBuntXeSXYqWHfPOBrdEP90Ug/yIu+C
8O03FLEelTvP3CkPt2tckl6lllbq9Kziw4jBN9E4ixJ25n/Se7aqv+AgZdl7kLLB80Ev/yXzfDq2
MdYBdvvGBke0B+sSVzNo1GKCd2p+WaPgOFUP4UohJjR1z5m+xCMd4eeHgDDFZWc2E+g6wLB6Ta4d
Hima/vr0LUvRQjZcmMvE5nfxyCVu9rX/dzdDd2Orku9oOVihK4Qho7DSMK5zfQsZnFindfvnXuG4
wqdG8IMSstVylei0Y04mErkL5+IvKjYsXLSPPO+vkvNCPBJTVPXhzu1S051mAabBVbpqXu8PvuaE
TiTOTSUaZGkIzWPFAho/UXSNmwMSEl3WiTwZyxPzVIrWJuboYhsEjW62y/SMbhLCWvsUk5j28YCt
Ay1MF9cFyD5hF19ZiFmciSohZvWyp4BGx3eflOhEQ2TnXurRc+RSxOryfvA8XuaQAOQ/Oh4RY6jX
PwRo/D9W7dSG6qFvtEjTlKEYBBqH9AEUFJOKX/7z27+vgWUtghgUenH90sFG1k5JsNCu3urytP0b
NCIVIG+rqEeUa4r26X6p4/E7pfbB66Eh3lLUT0Kj/6uEsNeYTFrr4hTIvGqXwEZGwAKbbrhaFPbB
6xWP1vDrzONv1Gt+1JfPU24Sbx4EHHVH/U9o4w31edFtR5uyhmV5ubkSO3RNt7IqFz7a8fvwEZTZ
LBWjcHUUJ+cRDVQXkknbfiJmowxCyS3lS9OPwGj1V3ZnA0yLvaePMXOkc1pgYHDdp5sFRSYPjnS7
9+3/1E4CR/HpYiqFwAIzkrmLgELfLW/3i7sTCblDy9Z3UMqDxT2xjPYf/TZeVHubCq6ZsWTTPR2K
Iuict1oJOifZwKmqP2jkyKEVyCCp4fMp5MDZFgrLQINQQe5ikgJQU2SjUkEEmwvhEsPFKuhtUsFE
7q/Cpj5E1MkkNHCL5FnMaPuukPf7y4C5+6mC+GCiKZpNL7aN1KIV+rOKtfZk3OZNQ35V//yaUW4f
qcua2DSlzbs/PMulmbpPwksW3lOjO9Ae3NGaO2+XAqYKE2oYLue/MIdHx+SZRaQgc0d+Z7D+CaAT
zYoQIbxe7pkZC2PwegmQaBBIVqBFqSR/fT05BKydMa5Fnshahsg80UZ1vQ/TFo4VZ6a2UX5Dmiyb
8zGFJGOsE8q7tgbDpdW1U1/gUxEU0X0gkG47DoorV8hG5EXlN4XzEzRnTFhMRfoVZUIBDmwLRoDZ
8Nx39rZuEbQV3WltVHNPzyWaU5GZlG4yBHtCaQlIcbawJ/0SL730m94VLHLtqFg4fNe61MioQxbE
+DlO0e5etfSzeGT/vn6LD0JrfukWYc5Acpuf0AWO1x4c3Bl33wnM+ZfHFcSiykQ7vEDbiSi50c32
yKdqfiEqtnSFfpnNvfKGNvvort7BBiuOghxzNPuW6IzMhcyxtInns93U7LkT2BkXrwJNJtpL+xJ0
B3J/5tfTyMwH6+19dI9VRx3rZ84ddCTp7JuBPfuZpQnHSAclG/hho6MIPuNiufGzs7xmz3FHSeFa
uCOl3S7h5ZrtfhDt3GkBOEfBFvy2RcjWc4FUXett3d7j1wLQBhbO4yO+HlF4iKLl+ZoQZifAJmbW
xoaHpMD5DLc00ofhVllYVcH+I2fAvBW8aQr6oLKdtHVRxZmxK3yy2FHKE+wSFDq1GFMhy202UIQT
YnilpEdmTxAxQ5uIsSUgYB5GbwLaUYUlakgUK19Ty1dcYKfiv0Uv4Xb2xPGyBtB5HJ5X5tdZJf+z
FgJW5FL9PkDuFwnHu/67SCfra+VqR+MYaPlDqrWuiFDt6NJ2lWFy6Nj77RPKmOcSTvq9tj506gG2
uadoRL6isA5h8EVZwjJT3sBF6AaSeq5WZDZRDI9hzitlztipA0rF4inFw1XHNYx72DN8Dd4wnUKz
2rQkPsJs8+hcpElYYGNF6jZ/AY71Ie9JPYsijOl6dmsBiAhsF8ibMOhUY9zGiDL1fanZuSYaNpPz
aDghGDSF1Wh5Bf3ulnnU6bndHaNw6rVYwLLrEhfUQDVcTMU/rFDdrEGJGcYX+/drOYUZmjmm5kHJ
y7lXYzkEnSPsh9NaIociVx7vqVn9njTW/tkJEGUPjl9tujKvgC5IB7gSGB0O1goqRiOveF830BDX
VScbxJtXoxENWDT/wg19QJILNgxJR9xwiAGXFcsTi2AqIvcBliTUFE0s23KMPcqOHR3urtW1xqHl
3wCM2sZUtGflrsE1/ujYYFtVRONNDBhUfBztI+a/io4TxY+Qyuowe12RCElqlKZeSahdNHUEAiuT
zs230sTm6AzhjfI/S/fgJeQqc/BOL/+jPyB+HCnE4StSuv1fjow+HKOWqpbimfXx20/GyAXny23E
DAMbrycnVHkSvZo6r24nsGxTxDxa8Qgqg/nZyKMjmzQChzjs2Z5f6EEdv7H/JKE59VhLPyHTHis1
GCqdTM16EYVDadrC6e87rjykv6R6kOopukCX02qV87/btO9J7Aboe/ZN3IYnBhjn1AT02PHRfJfH
+Quy3VjhCLbSXuFQ8wI3n9F9uEcskXTexVofqQUmURXVSK4izAT0NJUytN1yV9QjluYesIB0bS5W
fEIgl2ksCz/aMr0LFv5X6CFoBx+lhdtCJ2kD8oyS5tEb04kzXEhDzcdq3WAJGVDZnxHu8aGzODiV
7sgdwo1w6IaJsiyKG55KJmvOWZK3sGTZ63kblOYokxMmmAOrMHr1H1Jy3zZ7DqLW/h+wHNdlLryt
sHz6Fxm2an+vUjESOc8Z5sKGLrzlh1PNshvSTPyyxqHnWD4zEG6J98BheDpZjQqoOWQSlguuIWpX
PxXv9bawBram//WefmUyiAZi8652yW02y4AFhZhZf90h4VunaQLIDEKDvjnTdGGH6ICRRCzAS8iX
CXMwAWaI22Vh1Jk9mTmm/4Gblxgxy3OWR4vJvXdw8M1W/Q1BXegwE6rCcltXG/vpFV6TinYJb/Mf
uYQUx22d43Su3B0HooRudBYv3mcyRMknwglamkX++nxMQw+6fO91qK1BTqLPofbA0LISsJvzVjBu
gQCYeYCeYJvRrmraqCmwRxrfBLBEFBqJ421GErZGsKCSx3thNq4RiFJK8vtg2VQuCYpvo1s3b0+S
wjnn94EzkkRvU2sFX7YYu4TSz6qv090izl14hJN8d2bk4P/z6+GmZD4NX9z5gZbtTSh2eK4d1w67
CYqSBB2x5JMhGN2P1g1PW6Vw7IIGbiprCIHvz9V1PWmSS1jfR6f7adhh2qhDvb0IcykK6yh6jckH
0SYvAbM6OR0OjYpVkn89RU2mO4rijlzQT4BbI4xZHEccEWpQSsVJSErPQ+R/EY67OnYNbg3Qmj05
mq3N67Egrsfr5dUPm3L3Ws6wNOJZ4l+RYwLOotT80GQcxE1oKXoEOcK9doais6rLLYqEHrV9UqOD
EC+OuHpx2dRHMW+q/Q6YJWIRKzUKnbYeLtsKtKOVCPwln5HOiNlghCeEp7siWFw+ymQ4fg4Kzj/r
4GBX06GyXwQGPb7HooN9S+AN4F4oMVVVD5ad1SgfIcp9/SgC0yzjFeQC/KLmOdTMFBA4z6UmX1fJ
70Pv5qfY/PAZtzMabIqc2y63NSXTcprJFjUciWovEz6CdkTyXt8KHEBg6XL2iP6Iw6Bivy+Ws9r2
HgtCJpuE4oQcxbdzYXIuYrGyuAjfRY6IEBLiu/XsSSkekqGzXEY4fa1hMgndx9QUHI9ide0Fj1YI
XTqelk/AQFbXe3WBR0+ePMsRZgJCDMRtX1G5J2FiL2far7elPkr9FIfCTV6vQI2WXWabXhw4+isS
ezaXhu6Q8ePmnNiPI+YtUFIxBs+RPBqv8NLplLy9X277/TbazhWMwlBZMEHBbrCRuN+CMGt6SR8/
aYebVJjpTjoyL3k3k3JkZrtuQWA+nsY4sK6pOBsXFtJC7cttXVTg6WY4bzwAMO0QJvwBtm3oDpUS
bfJqacX/zfIf6J2c46aATC+B2sV5H6p6MU+C7hqTCm+WwRDvXLhISPIci80nov8xB85xhYXKWLWu
nntfil1RyZ9rALkPAKsaDrNBKI2ZhydrIp+UlCjJUbVEOUrW9tEU7LkOxUrn+S65VI4n850eNwmN
EWZIHLxaYS9LvN39ckfgyoSBXFLx5Qod0eQXGu036g5/dXqZQh2h3sPE9grQOHZSC+7pu5ug4T+J
02xs4Vr+dgeWe/rfzU6DqXihucPwJ1iDd56v8BCm6xhDo2kvyObceo0yqmMslUyA5/oI97ozF89C
c7KL5raGg0t6pqQKMszS8MA5lwJF8AHBJYHBX8EAccKZRUT37jV0AetRgBWytiNp7Bh7KP2l4Tyr
qKGrSe8tyVYM83rYkgSyAA+fGvq5KoHIbqo+IXFsZTepaFeXoltaoO7AxPZTDBJUwFosPD3wqbMT
K1IOQ+YARfedTdtIe9BedUafKs+AlXWyz8okRt/sLeQ+nhTVyCllCxzAIXNpnizfvgA+FTJGX9LD
T4T3WD4r9YfWC0CyEQcbMcseb7boU/jPI635bDOojx3lixhRPf5UXI52WDNMqcBPnlH/j73dEhTo
LRGNdGI9PFqRFRvUp1aZPVjTpUYQFNglBxbLWqRbRLW+yrt2nQ+ketbvDQPD+qA5mGD+qjKJK8Ia
SH1L5Gb8cJWYhtKWxkNSwsp/VkmvU8CBOM9PvgCmKqitFSwP3VXJkEtdDXa0gghOUzUfYFU1JVDx
fz0jJMz8mwY5uRwR59qoZBr6069LXDVG2JHuWpjXY4PeVEIzJi5P52mLXqQptiYvb5bQpVJBhCjP
pgr/o3eNiYG0Z0JBpFRBFA1QjwV813MK3Ea9XPUR9YN9N2LqltL1Uc1VD93s+9XkdOUKPGfLg9+Z
j9KeCETPidR9S1gD2tFNU7+uR1uY2KWhQ+KfT5olSfMgCy6HSqMKatUqL+k88npjNiKrWYVxUatm
OA1vpEKOuisYeXnxctvdzNyMfpI29oX+sejNpuj1Ent+/9j5u07AvosQgAEybnldynvotdZMxLQe
JfWYt02IfWEs8FWxkOYC4jhuZJ+UQRFoHWW2/tWLn33EHzUWZEZSzMlSNfKHzHqlBnTGlUZ7k9PL
7lxQ6qoYc1tG8H9f186cSB8OG+ly+p7I1AnmTgmoRKAVGmBDD4UKWQm/IVST/viYLCmEVcYRHpVu
VvCtqPtTaVCZq82k2iwTiKHS1ZzzGqWCW2vcVEZMK5W5QpqDGVN//x0IjikcgxIeJ3kmSI+bdJ29
jgMqH3ooAXsHv5XkaLdaJkcU7fhhfeCjzRJ5Fq+kyT3l8PW+NK9pUqTpEubYcUD0sIbBBnTiuM7A
GfD/5oiVNsXHrRK4RNCc5ccnypAsaQHZ8M2LJxVoaNdCLU/8Edn0hwhGe+DHEzw5zfVAew98de1K
fbsJm82/6zNKcDMQhirjuoC8qdoFcelOizvTV5a49QhxoN2WkgO35O1gO3GIk5WjoX4d92f+YjSK
h8lzXugPedtA4bkUye8+l6mH23/+WiGDloB1BSmLTnsUrK8L/siwz/C8uWij93TjchL4GsFoi4I7
dD7Gjh5uq6xN0GkFOBr1OLbpkdUWHCJnjQ5p6sfSlkns6RViIKhBkN8zXEOGA24GNDhm745qaSZA
xhL/sbYZs2JLR6jVnlQ5xpKwVI/r3pb3N9EOc9rsk3qQGEllhjIbus8L6pz9aiVLGoS5eun1oHTQ
4oXqQhOR+Imxfp2U6h5s6iEA2P1uDtp/T8DWhBKqs9nepqZSSTTEzj+6ZBRkjip79/awkQgs1jL8
FSA8LQmA4w1qdnLebdJL+2FgPM9e00oz0dWux/3kr+9GV1DjUz4BcOE1dJhQRhUswX3Szg8qYM85
V4sbAMhWNGpB0xMTJknBJCaSscQt3KFm29bPQUTsB+7oUgZyHu/o1vF4AgBWTafWS8RdYiJ2c58F
ksaXi0jYRPtMimjh8K105Xf+h5V9gVJSOyeXwSA9I2F/Vy6dTN7K7cITO5ZOvkhhYngmu37Ev3mT
SYllhHSqw0u0/FbVg9/DKb9O4V1pn8ZLYveM5Bj/ZI5NrFUtOsBuX6MfdmsE7OTOnSzFm2/sq/7N
Vf58LtWxIXFi/rbPunivayUJCaNquEfkfty05S2INMADgMNfmq4kwg2cGePY7u6G8mjYSeLJAfqj
zCrDd99f1zETeohnrNulyzC4Au6Tz6G5DsQY6rgO+beFQlQp78OV6eLlySN61nNCTJmoKAStSivO
5b6eCYMb6srATXzwdhn9QJfm6YuH4m5FGpbe9088/JjgfrfCiPB0cLvSm7nDY19JaCaja7d09Kjz
Q4VzSq8KqxJicoE1fEJOQkiRJSvSsfa4GPLqOKL6e9eFWglygvh/hYekkwXp/ZYaEM8cUCy8QTqr
8BffgyhQ3TQ6fRVKIqbALKUCGjeTgVxaeKjxb6DtrEqfTGMEnpgeFZJnkFR7d0w1MZJxprY8G74n
jgaD/gCTKhC1e+BFQ6Nc8WgsmMoAREdB624ZgiJSpKr06pJcjqC1BPIPm4M77vyf53YGdAkRTzcg
a59fX+M0GwpiBjeVt/iM5jcaGNsuxR7fu/v85/5cwZdY4Rgyj3jygohRCkYo13Bd2raqIacHKdmG
7TbSeRQGC8onAqpJfzbZt7AYKW5tNVFpH1QueLOVQbdv3Q4aZOWdHthv1/zBozj9fHlj5d7VErBd
aPiQQbdoOa6l93hTQ0HlI8GPf8ECop0dlzgld/0+YcM5IE/l1YKCouOSnKfxfA2Zp8Xd63jMb/HL
oP1Vo8K0iKYoyZqd+KFUxhjfEuORqeyreJOhV6OGjhih7sa02iuNyts91KFQu5xmPekrpTBdD1iQ
56iqIwTvXBH8Kd5zs5IPzhqOLXHndMNygy3F5i/pPvzg4lIBGqOFN++WBZ8GbCIj6NJ27YXcsCbk
lNcR569owMS2ksR7CWH6lXzJYcyrLPvXJmMwwgl0xnv/elRPP3RnA2HiwH1/7cj8RhiM+EOiWkCY
fHdinOBn9Uw5QIj+uWeflexAvJ7eYv2cnZ+GA+0jFCRTUvIjpgQq6npiDK0gDBqjc5K4pRkChRN6
wnXA2Vn+5fU7cplFnZaD2fhVyrgniM7qC9YxgMMI04e6zJWwtkcNFSfuO5JJi1KYMGRaH9LkG4Ve
2Qysom4I+jS90R6fXwkRCJAR60QO5Qm2od8gZLCMBve3Rfs2w9qI9HOblR9RIMHePEGkbcoafE9c
+nF7Yu/CwIbsCUQe2cz92DBqtIQuScq6vMvTkWyBQtAwLEgcNZLIwoDEyDgHIEgIFCBWmExG5rv/
R0W+jW0p3zPcFE+SYRrtOR0rS3fgtxi76HryGrz8hC1pDO/uzHPASdXIqxfmpAU+uqVFp5wnqvbm
hbAP1EESHOXs8J/q7BtlO9jDPfyRcN3vDYSWxY2JLNlmRQYBjk1mq0BmuKNvdaqoHHd1QygSGXii
0ED/ld15YHUYghspLVxSizIIzg/sNhPhna1ubDMZALyxD3F01YrD0zArBBbSCJvt8ZbZ4AVFBsSw
bouv4WaJh/m4yO8+ZMnATuD7O8NBElDyfBpr6CZttdxOcn+T8EL+H5QOKzXPDMg/gOktYFboSS1M
c+sNgEO3kqTpu7YXDd7kornl3jC0CjtYSatGv4VQSrazN61teQiX9k9qLaYIyiHxzo+/SjZhoXXU
yMRRqPyjd5iew6aQe0BqP9RCTqpLLcpfhkkfn9fpJw3V91jAI7iZlq+w98qZr4imw1JrfC93HOUU
pdCKQDp/ROJUsEopCxjZxGl28FeAyWsUUPQk/rIoBG72b0rHicK3cq+7vgrtiwiEGpmcxfJXdCTN
EaYgNnPwP/Qj95PoH32ZXIMYxVnzPhtCuwdLrk9h3upDSDaERBqw6p+8yV2/20HJ00l6lp7k9bI5
ciJsBwx8Vu0G6Ai9SwaojB2hvSgzxJnOoX28kpZbThlnraoVqLkfOgtDjtD31auxiARWh5gdcisa
fgys/89tuhEQSUaMIrPrelUAWhhRBdpCLT8TwjePtE+d0mJR8NX0/qoyut+Uj42XUjpw2cTXOKwQ
Vvkc79p1iV+ODtJAOhNxixJvJUaU+NZnofm05LBS+HqwbUD0faWTW+ZQYGV+ixyJirUdMl0/FcQA
IPgSjn1v+JePklxuGiYVrtU56nt4XK2eZeT5MVUf90r95IbX1rChAz+2u5t+qUC0CThMzzouoxk5
xEbh8d3Cn9Hi+HW5Ipb7pYLxYBrtKcBAZAal933ln+lem73S4hKCi6a/zHsGX56wr/ax9IP0hTlo
7yvFbUnrN78EAwAiZrXxHaK+dNGCfTEMlQt702Qt1Yxy3c9zmko91q+5aNNzONvb2pK/vT6dIAXh
NpnYpcfen2gSP/YHbtryvTBtVGGwe7lsVCLK5q/A+w5x51E1tSJ5vA1ye0Hr8QvzozK0DffX38tT
oAfvZQ84VjHGQFsAwnQGEITvberfT34jd2IvDoayw/DTuFA4j0UXKlXTCYt5yCjX7aANpkG9RXf8
TgbTBBGA1cxzgodRmKFakGEX/b0asFIi6Tl3hVFpz6yt8rKvKFxPwMGKHuzjMZDEA7mG1K75En51
9A9Oe7YcwTfxLslQ5Nzl7OFh9kCwBhsYZPbpaEtf4TWzf9WQObbTcLQddZCWFRdNYU0gbsI4ly7O
4Uu++o6NYax4L23TyQodtnBc3WOl1IoLgkdX4XB/8XCnFWnId3Xv8lOtkU7lERI1tbdJ8+DNC7/a
AomGqWKCIdmTHrgyk3Qx9uM5maY2hFRlgx0cxTIefbHayNZ/qHG3ZVgr67nzBiIJgu7BdHjgXHbx
b/Ftp7LfrBiSXixkYR5l8KkRvU1po3TPHPswLQfODR/Km2NTU/dk+YZK1/v08kxHF3QzQvaMN8/x
iAbYPy50BSPVnvL2w0sZrMJQ0NZaJPLdeZVlIurF2eULcCF9mvhdHmxfPJc0dgvSU/BcJqNExoKs
iS7BzlsMECn6RtvREuT6e2GD0I4ncSb4nCfNmB6kstpMta2S62SCxixZ6D6JEEtU9o7t6NYk9Its
ALntPeqt4vnGJTFtdZ+qGKKlvB2Kho7T4S4VBeKOMvQrGkPNLuxNMwrpXxfecmHdUYPd2erUisKN
cWKuc+v5glPU5797CY+ZYf9z07VOk3kvFKoDmExcCTckw59+JPHMEDmuEAT8KSdcnEjWUdUVcStu
L8teDHAwArr2x6X8zp/GSNkHmMxLDjAY+D2NLwhuj+5+CHB91yYx7bPnxlwSCrwaaBkDVKOUFBUh
I3r2KQWWEyyQ4pp3T7OOdRxRHja/TU5LjtV4m5uOz8XvOyEOFZwdT+8EFaaxR1cZdls2qIJ9mlOr
O1h6eDHmZzTb5wZZEIDH0bdtOpf6HRbIFml/FIWualiPHzhv+R6A9xP3EBtmUDa2j/SANJi4u2is
6iS9RMnGiNbUN/FUnbm0IbeMaiL+/K588zXGxwcbtrvqDRWX2yd2fRQM+6mmX2S1Xj4yMI3xaMQR
5rDVrunNGhIhLbpHMOe1ZLvzqDbGEGJz8LgSpPg1PDnTZhTIx/frBwPsfgePmL/Ur9FW+PJIJ4q8
18toUDkAdl3KzBY/suHbAU/aulvhBaEHLogtRLUGdWpWI3JYAuMsEAeOKFMxu1Q0vTuhoVKU8YU2
M6tTyZ+UB8FCpUp0Amfb5BIKLjyltrW3gm8Obn5i5H0dJ2VSuW2HAUUoDKQ5ERz95UntzW3ZMEpx
80lLF+pU5+uA2tNw95ruIPdEUldkhusn9fq0I4FC55MV9rehFM9aYGYLA1BegFbRoVNZyB/Cvfud
WbFmUZtHBaVxIdeZb+JjBzu6eopTybICNVqnT/ZFPU2ONY3MN6rZCzkeFoS9NPTWsPpHl8xkMQbm
cgagdWFO+kidx0MKjSdxdc4ImmkLfCIIPkFC+M82XpJukf5rKW23orE8y06eQopGA+Kou/Xd2m8V
gm1ueGl4IyL9Gr4zbYtKFWEh/RropLy+5+Az1Gp9N5wu3nv0mfEUTatiEie1FltsdLN1bx+gKZOX
nwANYDqOr6fX+z2nJceR452mZmTl35u8/5S74+0IIxdF+W/ZxA+4f3kIzMlx8cY9uPOKDxsCG893
Y6+FvulrdLhqeg6sMfSQfkcuychipZQq+nkoWPTnw2OmtBsMXgMsY+CG9vrYb1+AFdxLKQY5Lb59
zmR8gxSJ539PUimwjJeruFF1VxAVEmqsn/3sRkQ0+BXpME1i1bvCsetL2FJnyeiwkAY+5JiQEjON
fzkLLm2Sf/RPBxQ6mOlqbHsijYP9HakekcXqGZdWv7a3gWhAkqn5wQq/pLDmoT0xEvavMdUsmGlN
rJAkToCalGYOYTdGjTg3CUnRXn9obMALvTs2Ltf8kmdCl4uxt1rNjUkSrZyvAmEsNMylMRFK5ayT
mDY9MJh2vbhnewxOveMob3XPqeRlbdIVTwi3zkyeAA3JoCweOJ2N5t1CDadV39wq3l00mwDX2QOh
uKP5sUyF/zHLsfl/vpme50WxbOi+LigGKnuddVkYBX17yJa3TxTNdQyAWKn5JyiBoAcPrX9mr6X8
cZ0awtkvzfAROAQhUvI59NAKGVCScIm4+YQ7hbeMc2EU36+a7igafVnftBzT7TV27GEOJDEhLXU1
axIH3fAmQu9ey7sThavyW9q0Rhg6kq0aP/tYzcsUFvchkaAEsGnIdAUJtgbY5H0oe9ncSBqt4ucQ
ue7xdOiSrZWqFcXIPZ/u7WzNMTYTja+0QN3kKdklGW09cnFaqlb47VljH8gdQSuXwhH6fytoBLpM
Ubor65vDbxMadMZIb2ARqKK71+tzIaAwmf4b5Fi0N4yPpMTiQxYG5Cz7pwU+xQ9j7kXUTeb5JA1J
Y8lm6eOK/pdpSxX7kI2t6icmEy3PGHSlSm/lOyvvdlJQ1xyakxH5vpRQvI8jRYk1BEFYbYPz2rE+
xTvAglfD8UE3VCr6Qj2xXSyN5dgUaub1reoc9XwCEztyBvL3lpXnmzPG5x7Iym+5B+YHRYefC5Ul
en8Pk7XxlLrao9DerHSY7sbhGrMl6Cy05SCQIqyv8rapiJ8T/HYHrF1E2b/Ube4TWjJjvK3y9O37
dnvrAknzXYMjqN6FKVlqojUIN9UNNCRV2hIXQhyckOTFblgohbDhi6/RW64GQaVq1Owb4h1khpl4
ydMaCfsc/a6v6E7CbuslD/Qmpb9WBTsjN6bxgliYPcyITfbtsWK1acDYicy5WZK1KHztaE2IAycT
C0TOCY3F/5cSRpjhsmcbbz2+nzXdsarA9NPzXtL/eTmYTA11w8GXnt6H9FE1SlFzQoV25B3G90Pu
elR80wEFNejgAGUfiFCx3FEdyArvkonLO98dZFr3pDx6g4QuLuNbEgIbdgZxpDakfZl3sI9jZ/w7
duRfP1GKhuK0rTDxDr8U4aVIlcpAOVKWd0rZu7lJI+PoqXxOWQ7p3SDDZni+3scEfpI9C6jpMcfR
O17e+ARh/vEASkoWS9L2P32zvT5bE4l0lxEOn2niLMOgZ9pItERK5T8ZBX/fcEUipKquN8d1yzlT
tUml16WkVNxpoNh5OjLWLU3VObBBlHh22UQ2SH0es1s89OWHlN/3oudi/1atzKsZS1S9QD5KPKbU
1wOIzbX9kbIAxnnC9ZHTyoCEcgm6K9tA+538YuF8RI9kumb30tM+bqyjwMCqCEcX0djqfuxXlhIa
9sfpT/Y2TFXatys0pQihnmztCRxe8FdSReureb2ZtG/xuwdokIyU8r9qK6xbZ7BmH7s/MYcbLfE/
2qpJ9JFOGXveSozEFayUUSA6S7et/uISB13ya8Hv4IMQM9V+j9hae/o5j6drQ4iTsR7BQJ/G2Mx1
9qPYzNm4GuMl1Lm+5KSt28iBVjXBYw7PESQe+OZVNoHJope0HGnezm6XA9fqPuGZJg4AFg6Zgfyk
e2fyxuZt23+m2iV8OB5fbxUTbdSVad+IaITEOQilQamAheftwNznDveQaMf+gDZa8B2ZJB0cMSdM
QlxGml19C/LZhyG+etduJ32b7nN+JnkUMFZKChIyy15f2t+2uxFs9ZP9w6IE4jfQmaSFUlZ3eC/E
BjbB0w5gVFfEZa/2pNMlXjjdlv61qkeAF/QfsNlAymxX8qMvUG9/EB3L7k3vBF+NjlcchyAWnMWB
EyUVtxth9eDo1q6lEO/emKTAm/gST61+rXv6RHrmoW9efu90EBe2XJNalNJ3B5xG/M+0oNkTE6Nl
61dDq5UiBqD2dK+cfHO0183PHQGCY7LTGg1mlQkkP0fzQYhZBxrxBc1JU3D6tQTErDFvkzcLUsYP
lHTTnKYyxCNUGhQOsVJeBxorHbjzcj1SjCtOOMTMhDuG2LatKzqDanupw+iJFcU5/NezdyHU2zJC
cG73W4sTjK+Dz0DYCYAptIQIMQAG4rs+L1sSb2AqM7RFwh3lloV97UyW7nE/bT5EJ/zJKri/rmD/
U5dcK3okuYRj+mlx2PYyAk3+zrpKnRph78Mgdq06/sY8g/Rs1KQZUFXo4FPrfP5XJzz3vZ96T0Sq
TH4YEaPRdnfxv0/0gnxuhJYF1ilzihqXqXOMJbOlyEHM6ial0XLebgNaAgxLwzyM1QISRlu3skvX
Hq7tmqronpbkpPYc619TBDTCKWHZTISZOhbR8RQq3etb8+B66c2HEGq6H30ztWOdNesQPsGK3iTR
MqalAYoXWl1vJoM0qkerRi/ZHrG2ma4R2vldOGU+rDwDzmRaIzp55TkYJJoxrNYeoSPzqETuVVPL
ZVFNuDoAIIvpQGPpVdDosW+ZBGRwPBWappRdq6JvFiXVks7Kj+yF4kPhfeveZWoOC09pkqPSqIxV
1hUdRpmSZhbWtMEifOprzuBos7P94xuC2AYXJ+ispZEngDMnSMOWDIrq6JsMKFtkuGimGasjgjxT
53P+shBHhqbIB7Ns9y1avf4Cm6NjixZzSuDn49v123F8ab7t73Fq6syga0jKzS7gR0IY3X0DrV3K
h5pYhpgpvk5jWnSjdz2Me5JjQc7A3MMvbtVLrs/i9aFGAz1GTjUHl2eqWCdcA733qUnacHLJGBGh
1trY9+bBYeIzXMy1lIf457KCrsnoOk34My3ci30LWCExtL4QaSIBErLonS5P++0uC8TNsjzRV0Od
hvuWuElnDGtW9fP1q6v4CQW4X5e/r4RtRn3xqnbE9+ndaazgj2h9Yl6qIXOkIpwjOE6hCr90tg2b
gA8J66dZ0L2QHLKlM8OE61R9hEmj2OnJPbBYaR/UshxQ1WRNNWC1oBrTPrpKgC9BO5Auuz4gQ3rQ
2sEFU5lRSUFssPGc1S3EZSgxxS3rTYVbcnULl+hKyyytjROlzJEjPpaA+VaXdrWHsHSY2hdkzAXL
dMglbm9gs+KPHB+OQwinDvDD7HsTJ/tpY2GVoeMjC+fm4RjTQ+ZsTJA5KSTEJTaf66p6EcrKiNoK
ryVDQswpd88uZhA1J6hh7o9+QjXNCLtEF9lnAitOCQFgWtB7ehgOuF5DSl1tM9/w0eSwY8MSIPUM
TeYFTq6h2UnvQA+6GXl4u8OsMtAw4P9I+/n+hKlYjhxsP3jKHeb/vpQAgi+wEJ0rJhS8dpO2fEUn
KFbeDxDcjERIuZ2i1wuoyoe3GrIyrq27za524OXFUVtVcDB6lQ8ckSINBY23RmfwnyZ3B8N7PiCS
iJU4WFLb3pQdS1UfWeuCew8qQk1PHsv9rpjqAFeA3dVeZLZlNOnt2cTIltV4WEIarU1CAJKdc4tS
ju9JwMnkTBxjQBzztkqvOSzjSV2dWugl3AsmIar3sZNWaZBwKiuq3XoWh6KYkrIHe/j6KplL7xKB
t9b7wmHGBdKsJ58aYMOpCkvJ5qrr92wdJWIyWYgIhBEv9tSRtn+H7uRr+McldH1qTmHddkNzisEl
o8tJaYjOV42xAeMDjRPxS7VJVoEB8IcBfbm1i6GxwzrwUasjdo0N9084uT8b/0lKhi6T7WYt+VjL
BaKTMLibMOYtS3xb1gR92MZHw+4qf1QgncezjfhPZw2sunBHhkm2n93nESbzLaSPGPNwmW6nCg4c
PWG2dM6IWcvFpushV3uES8Ujc/bF+VMpMwwqm3J9THv99c6Ql7acroWDhALtt/uly1w7TBsXdVHb
j0tPREkxSSdopkIGJnLmqwy7jJjHtUWyAK1/EHguuVpzsa364XBZLwRiD7YwKWI4p5c7yFQmGu+S
kvax3pcM/ZZcn5zJ6JwqYhJ3JlJ6lZgkS/mUNILRNiwjG1TulKTKmy9T3rq/xLwqtOOBETs7QZhU
sg9dJo9/L2yyX+mVQPcOdYVdeM/iczB04MhSp7zk5VDya8JX8WCmAZ+M1RR4/8N3fkdFdsxT+uWi
X/CPrGRU2JAZu4DQmMjrn/yQbUOx2jbef5fkQAgKeMGO7T9YwyEp3vhFYlVlpQlcdCsS4VBmIQnK
VB5LFIPYuif39btSMFumOZHmdiEsgTquCZnjSYsSR5j9SJEgD18kI1bAMZTqdyPoXEfPPFehrZwj
LH3XX0PXwiR/prqJQMhPasdNMBQ3G9VznXjuo2yYXiuGe93r+2cVbVp3B69HBmr3F1BYIftN35aZ
2o3f+TnWKb8Rs00TB/876SdzYDO096NbTM3wI1NSr7ExYhZ7gMgma8J60HYu/37UIZPP1UBgSWgy
auMxmmqfWiDwLmwM6eb6yo4xJVsrp8R0W869Wz6I7Y9AjrhnOOBwAHREYKabZOoPVdGHvfu8NVJ+
ZcVwX5ERpagNdt+nBEvwXOmTaUMH942xSChbrqh3ncpQMCa64j0I4vnlLv0QmYOUXEbnUKe3JdE0
I9Rk6ERWHNP/6B92cizH02jXpuxAvoppMc7MeZwTqKQDUWs5nb5JnBM1v6VGsrVx6CQ/Fpl9FFpx
H2HC5xKeX+fVTQavEzdt7VG/Vg4ICS7F19xWsgCO28chjMY1k1mqaj0bqQ8HpQ/zKA6T19eSuZAE
52mxxNIDez64+I26yUCKP1G1hii9wTWd/LPf7L2KXRb4gWSBIknANrdODAPkVCmHN/mX/mJksYos
M/GVMqTQaT2yKV/6ZRncZGwT5N1WfwsgWuYQ3+J8MZK4e8QOLl2EFvNK7GxkKLxIlodsf0qZpnkL
weNUwhyPM0Z+t4egax2HWsy9cTS7tqyZx2S9pNgEWNhSvvo9jDjRlWV16xYeujSR8ZPOBXb7UNXC
ALV8fbBI9y0hWHpQwTBYZQw0Kv1+yB/h0qHY6298oh6CUF9ZUoUy+h6KIY6QpY4k5exIDV4GClQi
L3BeHsKpU4btK29dYqpiHL5JQ4O2lXxOAr2jfJXzpPhA6owAThs7D2t3KO8jET48HNXZRqdbpr+F
hTCPdmo5zCa9u5yfwCn8D0GplopmwKHCQjDRD3QrEpKh7b0FNaVqj6SL9AKNpRu/KN7LtRysj1dF
bpEF5RZeH1I2S9jruyq/zXopWeRAMBbSimuw3j0Iq8SZQGPpD+Ohs9MTqcwor+GxRRTH454sZJuA
Cf38cqXgilFQVHc27j4YEK7gTUuubcroQmXkC99wlur7Q+zSsybeWl9D5NXuplE9rXVtB7U2qXZV
ovq3PnYVVX/DUKAJhZ9fKE7fTcJqcCtJExzXiaGyryduH787cTCyqZQjIwNq0dI8I6cBOZqKYVo4
0FaJ2nDXLeKUKV7rMluBBmLkWtHIGegWDa5jw2z+CYzq60Pf2oV0RnJhuUFYzPjcgpnvc5FTo8C9
nQglR+trzBhLD3VrE6Iuvtpuqyugyvh7d8mEB+XJ/Nxp0SwhyJi1b3XvxCKgHkm7khCWQJyyCzIl
tfpaGPlXtPYMzEESpcK6VyI1rzd87QlLskT0XRsUmY3AZFCf+/DxZYLpVJLZ51ZEnY1t4qxFCgwK
L/YqUZY8Qh+YewdG2NL9sMBpo41SfA6DotBDTIYazZKjiJMIzt+BbsEba+hOLwJQY8RNeds9fRuI
6cc+NiuFhNJ510KZy7zWfcIXuBr6XGlCB5d1lWEGDOt5mQWvhGJ5xBVncOOxhyccrExhFyfLS9oI
iuWrfG5fU1HrM7BtdItHC7WUFc2z7iA9cx8Z2ZOtLWbDepv9wEEprFc1A9d3v0dm+00qX4F+DEBO
NICl9NRlmmC2NM2YTMvGGVh4qRlfQrtPTRUZsa1eYIyUumIsFC1XDCWw2Tg23eWS0okXsoJOFMdt
CramWwwg/O6Sc1L3yAUiRynW3BnYk/DOpIpDdBOwrPbqsSE763SGl6CUj8KAqjLby5BF9CBrL9oe
A/gHR5d4xYtbsLU1rTb9QCl0MyTT7ufizaoqR+UkURba9tkkRCCJyjseSb6w7yrFUdBMV/7DyMsp
ALwjat5qR+D06CMdvn1lFGJe6RzNUU1nEXL+ch/LoWWE7Aera3MtrfYOseUa3U9M6/T9p6aUtHWZ
JosLiEvnmbbRUAPmTM8pvkzAz2guSzHDA36Hocp5vW28AH5afN8GnDKQqxDNB0ApOwFYYPh4W5C3
COWqX68LvoFznUp41yqvAoPDmpta+e+98Il48ycK5OksbK7EL4bGphW/f52UptZfBDcS8ypmUbM7
+2fcHN6Ctv5AUrssiwlmB1T8avU1y+ji0JYfd73cgOzUmZT/F0wRNtF3JpdPANCWgbJF8+e7nm/j
B0tz1QTdBCkZ/u8rMZzfDatTU2cNh8SYR3DVzm38mHo3rJYtUeR/s8Pf9KmhuFb0Kc8XYvt0xRdh
g6ZNjCTooD/eSakFBKLkk5G2u+3sYqVx+SvHIfs7T6Hi0oP9g6AI4ZvSUwcVXy1kFP0U6YoASq9j
2jCz7OZAS9k/thhJxyWWfxoOJwiPyFPuPku2YEVY54/FTuv3jBT/wxIuv9QQ8WZFk8g9UVuueqKs
343IZYTzoinF1Fg7NUlWcG9O62UA9EBNFh6GWcpb3jgUrY2NHDot2ZQtCvK4+LvbIoeXkjG0+HLU
ZxvD2g29z/uCFBa9XiAx4i2BjPmdFeakDjG0ifZvUNivE++fzKYoFRbzMJoGvCoSwG2orjWowFg2
LA5GhDzFhxw9gEAvm5euGvUC7zQsbG0xwUr9RwOqDSjU04vOHalcKz18Mj5sDl4VJOSqnLKzGBg3
mVdtvDOYnz9OrI8VwzcRpZ7laQAY/DL/TXjYMIQ7aSlcwcIiHZoGl8WG1/HlL8Fa+Si9rlp0AGUH
QIMTugjeluGuozw8umkLiSF/OA0hX4+CfqPF5tffAqiM0aWBZ1hEOr7NOyrVCb8DZJCVlhzlJ83q
BZSsF4AnroWCGoZGCkH90AnKYtAKwAftmtq19VNUBnIgNvl1MVdT3ooxzi72HjN3BCQg18Tt59jC
LJB8EfPodPe9MpzM3AOfDn2bln4eY/toMQNY6WNg/SuNsn5IZNgu5Ompeoj4qJfWVI8LXVYLMYUl
mpoqMNk0DrXe5TawzBVU8iclm/WlPDI/D29I4+49H0+B/1peSupphO++33jKKuI7Cg/s7EnmlrEr
HJIEOVGt0hcVlhFCeSOHyJ6FbwFLM69wFt4F/HISHbNSIjLrqEfRgffzMy7ShNOU8uPsqtEUcTuZ
3o/9TJm1/EFm9glLkDpnmAQMjpBeYty9gpDog9d1PAOGj6n0YjstSesnkXiurVxTeOgCRpUKsmiX
nc6izgb6+e9rQ/kgQ6NXH/69+veHO2lAK3AfDvtZQqzTdsSVuUcyzJGi5sEoUOm4uxd4rIl9SWqb
zgBVMbU8DZQRYxYfUd/b4AMq+oIKHDeVsPH0Ec1d1eOIPsZKw/l98m/V1YvFNaeE7jz1SHqVQRT8
R2+YXEFTf0MkASJkP47KgDhcqrICQ5oIUaOjXLQBqPv9RHCXMJJL2wlOsEThyzgkOHsvHCrgwWjL
bNnlc7hELQWz8uRkKXIA8E00Pgjfjzk/p7ZbRFl+06ICAhRL97pWK4eNIZl+2Gqlk+1WrZTL+F+p
8ws4KOXC0GTytgCg1rUp9vKM4TShau4S+tDXAt5E1M79Ao7U5c7QYbGhOy+qZSBUENooMsY+Hapg
WlIubBlauOpFtP1ZjyeDWn9yD03Jb33T4zfVgnUyHxEtkPvza/vo2RYXhs9W91OzfEbkGEsaRid3
vT7d6GSwY6tsguh8a9NgfI7NNqGuokwnLFxzvfXmiZ+uTHGt/r4S6XljozHYFdjt/Nxm0/Za3h/U
Sh2EcR4ODHIVVVPWFMbnAsO262fJ2lDgpAQS+s0lgYp1ujY5btECRy8gi/q6hJIaaLBc8+NHcTxL
xoG9Bu67YwAE6zyyKdBV+YcinXovpKd6gAaBOZvpdjrHwM+Yr9yXC/QXzllCl+OxXKPLhA2D78Bu
uWTyTKLVj0fGlBHNCEKohrm2ezWlPZrZKxUC3z9ugxyiqSMh1icllTSCMJBHI0TlrruwElIo2pWh
chcNa7V+f/L4DvbcLZ4//POo0QrLJfvPANcs3RMJ0AMcuQOeHrCGkJs9TIdu0DsnNCbRRFuCIglU
4EjhnErcIVUOV7tq+BtELnZg40Off3fMsAMMT27fwJQr2to4WMem9ZDvyylGtM6VjUxyoJzvK+lx
D9LhhQdW/vRQpO+fSIk+HLfDyEI0vbPfmgSfh/AGOLD0NjJyZPt3yEPcFH+FqO+/Q7MEaqWgQBau
/5+U1los+Tb4KOy0/9LSDzqhzdlCPpS1RN8c6d5c36ij+BdZOwCiJfbdXk79aA74gjy50ww5U5m0
hsNQKSXuhCidu4CCaIu6lVWr7ndgA4toDLGatnnQHc/S9EjAPzc+slur4eJDyX4myXdLZM7ESmWt
Y7SjwvJNHfT+Zr4aIvQIhKjPJdAdQYJiV3p0oyc7XA2pwNkTrCm37UyWAgrNHwEAd6YSksD2TTJ+
AysXOoUMinhtKRAI8Kwez0EE8MyYpU0N1KsU4Nk4NxKxLRrMucLf3MZw7Ef3ZoEE9ntQ5NaMWI62
qvQcDXOzoDBtKtkTWtNwrfMrtkzKniXpXgYZcPj3ThbKEPpXBZ0o+PNvKm1eZAAwne7WIzWTBdD4
hh5jlFHRGCm12aFghlMVj1GsUlXatKo0rm2MmnthPVbIBr0WL5vskNB2LTp7nDmJkbcJBPhWc+SY
PM53ozFM1MXZ7J+1z+Lsj6IECOHI8l3IF5/piO59SDbWDMxyIKE44B4B9cbMBQ5nptJ6ZRIUxLlH
b8iecWEVa179WkxfUyc0XxtJw7ZHDbMjSXnSkkipKhG9vP6oGV29s3Mmdg7u+o7/QlAWjWTjx9D8
1RCicB4nsj3F4wBSJ6u3gJBSgX0IIWfbNB4anQQvvfFMWvdbZPV2IIM4AQenYd1eZGw3/Lv7IdWX
pVftD6d+Z/DGhhDEPa/BjIYK7IGD7Wfn0zo9WWmeq3HPJ0e9vqoXkdIbJch/p48AAG4jZbyZ0i8D
tJ/L16sA8zbBUXyorFlPIsqum4M0WVsa763olsGRJewESw9hBLxeR3ILMKP2H7WwbduMwsqY3kY6
4h2Mxgmr8mwHXIB8ArbUItc9MCQ3K7m9sIKRgHmcavqr/tyOQG0QHM8iDNKU2/1c2ms8vyaaPlMv
/t5a2UZdFhME9FpmJEQAp/2Hoh4AjODGCUZWyWetpkqCk3j2Ji1On2uvKmDDNtJdsf0ERFma9/0J
i18aUBnFa5NuMJfardtgaRL6mPsqNi4DzCm9LfQAjvqA/KHD4wFhztxPyquVcRRlCIsEXbciqezW
b8B7LpBQvqYs8vzzLInulFr2+fZkbdvqoqrmKx/ukmgx4c0CNHO6mU/+MMyby+Jw8jJEOPIwX/73
LvIwB541jywhvOJ7rSh9Is8hY/xzYXX0G4t8V+RED8Gnp5lc7oZbaxhg7oLeby5NseSR2F5weWg9
KNEf0MJlSOSvyjDQzFH7abupXQXMZNwSQT50ksZ1OVi1lCKq17KCVw4KZAaSCVr9jV+hTk/zrihi
T2ub4F4yECGak8PDZJsZlXuJrp71fxg9Ss7aEWGnFCsNdgB3mv1s/wYZeSYuCXULjXy1/oZY7XY2
3/PxOCOTmCNYnCH98ZGeDf5tX3h1D1nMkXgKBf3H2O561JH3ls8ZfDFmq6OdlAo8sNL4ZuDENqc/
hvgcxH5dUPd+vscdYUkIuw1j9WC/kIxJ2bmmbG/unzr9UB/cCEuJvrJ1DCptTg1RQCbJqXWbxjz2
yYPuLVqT0tBiHyGO8m+5f575gKh4KdiPbZtQ4wbLowqEeJQdz5InDv6ir6MVOuX3W01Dxj7g/v3N
Ut5RvW7P81eFjzYnfN/sD7tP991jJ+JfDHg3t4qXe2sTYgWgdIxRSpr7dWKHInycYWZSSE6hTWVR
4XPCSrxkXZCH3mFri6pKLTaSZBrVcLxopJzQaHA4nsZn/1/m/e7cz+zwZHBVHx7HxJN2oeZ24drb
/AaDj1xuh3h+EmLuapCDLtItD9cue9N/lJkkq6mpmyR0O0CS8LGEIx/wIKqYwB/RFr/d8K+Mcl+X
oO/Zl+dl0MOyDfUcrWHsU363otGpsjMhes1k7Ln4NdzydshvADi1+O2ZzrKDWDX3x0F5xx2Ikk5V
uEiGxYiy9SU8s0Zk44zeiL3SfJjWC8xM8lXuVAsv5IPiCBli2p6GZQKiKKc8aODTvz+M4dXkehyc
bg+TM5HJ275QAKEa0zpR+ystpkqF331CZJ2aRR3cW4UbefT1kPAGGzsiXvrMCs32O5OetIlGbcYz
a0W+PJD7GabL4FAVJzkiOx3ZHIptfYlIvHBSo1LSby5mbcTfjluP8rpryucavIDTahwuOqJkLgAK
Osjkevyx49GZtN2qITFa2aEAg08kT3/w+aq9jl2PPWtdXsU2l6DTUwg1s+0fsjaGx8EXRR+tF6PN
3820cMF7lHNWp1oxROsZE/AdX0eUPZI6zY1aMhPfOIUi19r4V6yj5i0KzDLOENrE3xFpsUyJaGcB
bh7X6K4T8xUB7hXlIRMTaEa1B5qmHz+evHBcJ3VfFEjw/IEBAB1NQ2G9JAugNhvSyv046rF05Q72
1bWHQdxD1SJtWlGzO8WgEJyT7Wdd6Fc8DpZIzBx2j6JEUxoD4RhnjPTDJkXb1k1WnYJzkcCIiB8B
ts4At9NIk7V2pLGr5HxYLmgVU8HRcUDOfVwTcbXFtDz2I6k4/7w0PQ6bQjkwE+2xqHq12cLOjPve
8jktUDF+s58tc3vdCL1+1NiYOv7TVrnZjIue1wa2P/i7rKRR4IzwXQxAGpFDsJkhHJVai/8J55oM
GEHiCPgAVhkhJ7tyrrJnEAO7tT/RcRRQhxx7uapRSZ6QvuKvpiA+dZAG8XXtkQ3uFU+UaJW11FpW
wr0E+FeR3fMIb06b/akNNX65r6iCY/dtvwAN/DtGP06AT7xGxsNRUnI9dOPR5rcOfaQT4eYfo4WM
cgu1KkDcyX0fWWkE5BRbGSSw38I6kDKOSt23epMj4vNxTPdVqoEJd+UMVqwBpzKrJ9OixPf/7lPv
++rl3IMP0IkHG88GWi6BuRcArFXXgHv/V9VdR3ADAsSQlQDR8oETNxUtSQqbRIbn+gIqu9F9Y49U
IfNOBygy6B5ph/ew7W6kjqiSD5tU3uwKZqqCcnhSWIeq1JeZM2L0zQTfwflebztnDDceYSl5ZH6x
xFVH8uySvSf92lMe6KbMWgTFA3mX/2EBdvTyj8x2Q3erqrRYruZWZw6CfCyCUOi5az1oY/Ji6Nn0
/epl07kzuD9hfHP4+JfzAudrRbFsvU/gDMS24sssi2oupyLe8rNmkSqBv0/86eGVT7yzBntajZ9C
seEh0S5XIUng/KRint2AevpQ/f/aYBNUGRtvdWZLN1x+mxlGibrDJdbn9tPUzqQKwHRZkXBPG2O+
gQ8pb1/SY1BSwd/Y7nONgddgG4eVA4hAK9n5aJ2P4GmAG5Mr7ht/x2CIu2LOzGodrRmmHDnwO9Dc
N6kVXs7N5lveOmgdtRl7kuhiAdVb1vRaw8kFrfg5xmOcaYNHG+rHb1W+2ZgNxdKx53bg1Hxpqdfx
pyRbhmp6hIASPioLfL6j/9pu1b2KXzZyR02dnNsB9Ux7JiaWofS9O9ew7MOelmtytjb/lfb6rV+k
yqxTAnNMlVkgC++VxF/7x7Af+oVdFX4RW7mFcKldZY84q1r5zqfz8FknuRtL83kfoYKZzSA66sV7
kY5PwWHsXNjRMOENZd7GxjdUBQ3rSVFX0NI37/TQtWFrlAyVeofpN03B5g5kV8tWXgKjg630HvXP
dUOzJuzDrgGBInS2UG+GI5tqfu49Q7yw8BrOMHXLhFPLqRqTAHnRCKlDWAsBYUk5pk41l3TCK/sG
/Pkyp8CTbLI6oZI7st8jBDhD9mVYo+ZvN356FXAtNJpjzsWOo9P//IltNZcp5TYfj+XeKSmeAG07
RZe7j7Y7tNzGZ2R9sntEY60plmy+4nOTImNalDX59VHjIRzgqkM92ah+pnsU8ULIv+HezjkJq2fY
YrZPjkxEq461xeGwvVQ6Gm6R4SKBBRWegqynWCC87eP0OMnQyuiuvuw9nWQUXSNJTYiD/PSG/cal
F+XUitjwB1+pVES+d2jgxNK+fPY8UjFwzCt/uuMQukrKQHx5HfxZJD8ixrv9oAX/fPDimBujEm0B
oGuH7sfjFg0U+a/w2cr5txLOI8dRuDyenbZAFU3yDwIu5We4caZzXyq7Uy/dSwpKtMIfRj3ByPwq
HoFL+0Z4MB2sAJDqA2t9mEJ/j1zgBNbn7OSOY4IbhoX9kJWbPRNzP5NwNgZp0XuwIfwRYnyWba5G
yLeqAO4kW0uwcFlNcomAnlV9QzxQ0W4jyla92b4CiKjLBqh9qGR2O4kTXVVJ5vcbqovqbtxq6aax
jhw2kxyP9iwPeMkHJZ1Ew+izdaO50NPzJDEGL0ueUuTWYeYBLgsFTf4LsS3K/nochPfEVfLCBZFt
72yPzfjX5ADOkqDt6OIJO7HRU57v+AbQSsAzi0DbJMk+q5wBhFgw/cZ6bqkhyJDnfifYDeiiUh8n
yOmIn+e0rRoVzaHY+svt9fvkY056ktoaSbNDfJIlJF4sY8NrFr5MIzTnsggVXPn0Sr6JeTtC1CK6
X3UYTJX710eM8osJvcGKK78CiWc4nzZAOWLeuvHAHMnzSkN3jV48op/yKeR4AMMQoGMpEF9e+CF8
mZ046OwQjxkQeEjvFRJyCw+Tx46ON321+AMc6T77Kl1axFt6kHANxWHHudzPoD7nKyHs5no/my2G
k/1Sxq0Pp2lSzfmqC4v1pBpshrJERyoos0CieAqDSUEjBVH82VLK6slP9uyOiKsBNBbcMFDmkL+6
dESwc9Hy8I/O0DV1dZ8cKoZdHsys2tFZnav8q20X0V5k/70iWSZSHaljsGh0+wk1EHsCwvubdW1U
aWVB2pY9L1lXVGUF2gHIxfN6GlSyUsk5UTS5FoJgf3e1hOIqMsNRA9r71LO4W+YU5y9CkfcVzZs7
K6KhQojb7DPskGagdy4CvksDHdJ0y20KdbSowMUXWdGT5UW0yyJZrZpuXsjIBKkd7+fQSUm48VID
98pTonYscq4DEzR6PUiDwBgjymdxNgdfRWZiPNMgqXb+6WgH7SsibQ+6tb9WDanidfyNyCw1hH6B
pku94xsBNKS6aMAHjuuasbG55BnlZh1zmO8FEhU5XfCqpOPBxSrr/CL6H05YVq1WYzDEbjcZYHN7
jrzqgVTxzqhwlD49tnPNil7l6mKFWa9v4FgvNPpG8NonlYJxAhsX5pB2e0hAu9lXVO9YrYgsT0B/
MK0uYmPAUJIvp9N3PMCbKynikXlX7kPYbx4m3Q4yH2MQhvijAKKaNSHKxgxpgzSCNLNXFf2bfCmc
7D7V9RinQ3F6r1w3w/XJYWOPCexQcInNCriifgFCyE08a3ahCa8HKwesM4eAQn1QJi2bdDZIfkRw
HUn+8L50ggmCQ0sM0P1UI8vj0d8o8AfKpTPrGQx9cVLkXmg0SekcpX7ZfNNREwZ+/5zsOs22Eh6H
kWPj9otba/jQfFzBy0jz9mjRXIHogE4ClcnJXdHo/bP8vDOQyrSJMj3anBVfPNh2DvaBmtWaEofw
VrmSg1ziWzpZEUoWZjcC1Y12D6zOSGViy18RLHEXkhA7ZxiLvGFubbbF7ophuMUwrpgXz91lVAjc
iVKtisn3vC1r47YFxI8HugHYWRghH7EwL8V/iuHIRYbASER90damvbWw7yTN5gI5fK58hCEW3P0Z
dX+Bz28hS7ekJJBgjTqgiKufO4CcZGXwenkAlduFPhI6HpkIzYMv84aIMHjbnfgSbGxGqPNNyoC1
zCd5cMZIcXG4KCNReeS/zO/Wm+Vwnr9EAFRveX3gRhwMFxqow52vDZ/OIQb+sfGN38QjkpfKSTZN
LnrAvPgP/cgjqKFUbeIfR/auQI6U/fBlALrJ21meckeWI9a5OuJJxsZ5hUnSM6Btwc2fmjMGD2Yq
CTInbaHHYRJb7HcaMNd00hc7jK5ifXIS3obvhM9xLpQCOvR40+kp0G9H9L+UcbmRrbGRa6CnTOCw
RO3ktT7dClLN75pPhyercVH1V1lK7J9xkRRY6nzpcB9kav3sgGI0OFhKMveaia+mh4cYTRarJEz0
kW6pqLS78ckmr8XH9R+B+qpZ9uI8wHqELoG/H+cN+c3aiKNWQ2hKt9f9kvJj8gI+l5OQqWEk13Ur
NjsJ4/QJfaDbG/U4J1VZSV9mqjdwH1jyUmzVVxLwGM83IlJW4O4nX4yOTZVDrXQx8oOVimJEH07S
T38TNBVgVc6RUE4T6dMzjr+e0JjwR99jZi3B0wwC1Uj/ZmoXc/uOC0QZilBPJmfkBU7I6QAdljiA
mvdG5jAxtFfGYKdjkhgFmI8FVdEjmKcI5qg9lW+kU0GECnL9O/QBIF3zf1u4eFrqembSwvNrtHzl
Asdif46qePpaPsGL5TaVdYYi2UgZqrsctl1GllH4onhf5ahpRVte9dAyiQ0E4nP6ZmBduY5eBeoN
Axz2PQBCqFaJpQ+QOZOU9RQb9+9TaqsFNCmAcQ981ETlE6+HSlnY+UJuwgW1sWN1194VTgLW008V
C6CXSj/PmDQqtoqeK40Kymc/wxuksCWTgLq3jXdQdc5s/iMeRsahhETZl2MBROjjeV+QyT9BI4H7
5a0d+3vG14iHVG84VfydR3zASg5TqUSG5MN3mDLKefqW/mRztA65tT42/5fu0Tq4rTPXfNhoP6al
31bbu3AcsvAPVYVcKJMQSepY5t1HZnfHCudj4b8gh1UrBMkmXFh46F9YRmpuPRtVa79Cqg4S2POl
6eSNizxzErtRj5ZHuNq9fHcYXEwXTTO2tTDwhxdw4x8V+1ZX/xxGczS6Ola9jDmJFIXRKCcNlUOB
6oU/tRbzAcEMqMkfuf7at0wsBSyud7s6/4+oYzltsah7gskL0/HIQG3tvUUmXI0Wel6Axi4hUGo4
Z9Qa4xvpXoHq1F4737Bff4hQ5DwtCOIqR9MlwmM+7ADSukLfF+6VVwMD7h2ju03JfFCP6Txr6Dc0
hqpeMk8waUtrzNrE2qdZoHsld255/NXyFFUvJXYazQdn8bfdhfDIkx2nEiqd/BHRO+eLJmSAKhnh
9vOLGQKJp6YEQa8N/tAbLM1w39qbh0bHqmi71Hhw7xvQGdlIaDHvtPZKVdOfj2JXPa5siPj0NfSJ
3e1zlalJRt1abte11m8KyrP2qRzCw3vMrQpLdXCheJgSD2dBPNqhJ7fBL/2itNroQBeB+PrrPESZ
ZMYfdA2pmmP4iKun/hEYk/ly3LNRmZLGMOtTyxTfINYjLmfNUFKnFSC9kfZOM1XKl/yy279S/fTf
wMGnOD2MKIVhE7zkR6ZeUi/dFa052RbLx/BcCFGo47Sm3sqsTcxguFwRMdQ6ehXR3WeaGEt+Rvrj
grpMSQoD3Gj3dNhdpEPdiz8IVxPCL78ZPDM4K4c+XeymwJc+ZTrS0JWMgTrw+yVCh8DomndlcPM0
/Xx7bTnJlNEIYVdcRO0zR2KXU1ooXXi3TrKHxv8uI/KnmEDOC8N6eXJUv9rvHqvM5Zoez/M2qYPb
d4lOVM9IKWcR3JRsg/YlYq92PxgWw/FgDp9TJzeNIiEsaVrlvVSanq/r6j1zMez1r5hlpyR5CHvg
E+3rvX3xBVdlu1I2+WcsNVB+CAY9kz6sGZVHtRs1gEK8IQlmMkVfEdITXqprcn7pLvdFmla3SZFi
VlgKrsyH54r6pOB9XkD1qah+94KxWiS4PA26D94JU7kHbiNUWQDfLwssg0w+/DsrgCmhElCvIQG9
VJunww3DOIFfTf/yOdZDyuIy64K+k7wFR452zNFjxz0vCM8IZlOWHo/yE1MBv3LjQvSyXTrqENhf
eNCbM/YpW2ojftBkreWSZYCSnvj4pojFI30Z8IMzuVbIPDMh7scgT8UvwpLbHscVmCMRKHOhl2U/
0dulN46VRLv7gePRj18EJDE7yLUne53SydPvvfGUSn1iYopLHyDjrR3jojv6+RitU9ec5MWbDFvZ
HVT6KUmpdsm87gBQ40+lMNVclFVNZ2CFTmcm83ap9dSS2Q1sC7Uc9bkJRJYP7Orao+MlIOTRn41y
wuBBDHGdbv46kzMeHBfpbLVOgp0OrJu+rC2284LHW3A6rx9eI7ADRqhVI8B6X7TuGiBC6PeIO6kv
8TvKvwBU3Dsbn02NKjawnmwTio5opcAI8IUMPZt4YIks9LgD+bhlgqSa6WqK3g6f+KxWV4q0akaI
c4E7qgcp4bVDXS4KwpBBwmdWpqKfWjq1k45XWRNAF4jDiq9qQuuvHJh1ivLonCM7mnJFVxYibqLo
dDvOJVEr+9ZwipZvM72HM0D1hTCh2uWZCDFWjzFnILj3q2ubb6epR43diyn1v/o/N7TPj8dMCM8T
+YzI6MD66VOY/9bQyMGOmJan2+Fbiwobbn/Mqq3J+SeEJWTGt1Dj1L12ccsfNe6LA3Wcw0cu9XIQ
5Q+tWgVHEOA5mTr2Kltc7QZKDTA58mgzkJVtnqUkySpqnpww7E/yq/MZ9WQ8LN2GSe3kMN9XPCX3
VLrWfMfIpTrtsQiJYDWw+o5+nhGcMJnbz6Cf9eHHtjBn5R0tDYa6XWMOKcB2ICylBF59A5uSX+Di
OFo0nR1YCtOe8I9O2pdtyzLEdoNxQAQgy7OP9HYfbmjulFP/kLVSnsVtnqvT6jOMAyvc5K0j1Ntl
LZF7uJankE+KnSvdpAKe6LntKvOm48CXO6ikbU0FW6WunRy5ElbR48sSaOr00KUMXTg7qdd6vVBf
ag3qGRCtTS2u8YLBFKMipJLgLJvnacmZD0QHDTnvieKrbzmAW8s98n/71PUH5XgIK+QMV3Y4MOZQ
hIUigrmjssQwgscLAwFXgE3/2fm1FhKRNcHQ1EMwD5f3mHH+tz0yvFAIHTPEXTtFLF875Y+gUKN7
Zu0MQmp2HMhBdUSynWTZ8Iz/Xi8Ku1PMqNws2eofsgd/vtnwUJcGn7MeH/Gj58Mpv9u5rggTC+ix
hrZdRtoOmU/XNCG07bQ2Vi6kjhIlxbKBpnjlrCjaT8CEv2LNh0rmYDuCs7ogjhEkWLPH62Kc1Fls
hKvzOgYjVVf+owOCJ8U9hVQzSPigFC/wuWjVeFtcDzGPkXaVzBF8bhVd4jwwWHfb5cf2aV6oiCIv
fFjXCUqYto6pYqws6CCH5Vo//YhzT2fV8IhgThwru2LAQZbFl4Ct/5l76AxlJf/U/NIf91w+G6/y
9CMWlLHxXMX/TPB3lT6L6V+gcpqzKq/hdPjKe2ojFS0r81HK0eUOadQWliMR3yt6PBaERMeq95D/
sKtVyLjxdLf6SubRMvTMn8mqwhrHAcenHa0veBp+Y5VCdG+JSTWw93xlMIIm/JzTzacXlmigjCYd
pfIuZgFoijJQ2a57NCpGkT9MAgh0XeFVT1vhrqo+VEVc5g5ZITJInGM99OZixJXPzzd/23izi+js
gPDDKIEb2HofzcBEasOxNIsBHm0//pjlxqeXmFwMwzlOu33+HOd9nkTjxpjIYrQ86EIvBejQoLcL
YkKXe8q75GJzyTy2TWAi8UDL08ogWDU0b/NRMZbpbwN2kXI9Fiw69UW1nuiBttOGi5WkJyHJUpRL
ZJD2gUGDRRX/067RQxvPhrTvTNx7vPZFFWIQpYsy7D45Nqrl4OjxUg1Rja50n1ka3DN847plCV5d
LybL4JEj1HSY7jqBnIfFwj4HGvQTV9NPnNqx7LcMWMCIHLSzYF1Lox43FZJSp1V2Xn3yt/cjDlZg
Z0vzjzM2em0lhox5bcG04PWtC/sd8aYhfGqdwbHgUyIvj7uk6zGmmnUNZlbIq96Dou8ITVH+CzBP
rJaTTFybLhDnFQrS4imjmRukIimo/NqVqyY12ZSVwM3n8PP70y2ndGACWIR55tcE3C0oRJX2iyw1
RxTzu2NQ62k7eMfNXi0Psif6N6zLCtibElUoz8L5z7ixztIDFj0cQPE1OZT5w811l9dUQnskPnbR
78fwmF4vR9+yLXHXpW4a/4h+ra1w6UjZheO2NMOsIdhSqkik0UG4s69h5NS8TwsTUGOlatt0WQse
QG5mcwRSWUg7KZRSH/LniwxkZX38UWqd3u1OxwBWaqKEYKmOctMNGRMlqPcLRWUef40zPuDjbAGh
zYF0hlG7AMxE3EemuySMEyXyEfcCYs+wLuv9DIrpvveqYkvvxj+RXjt1Ea8C95E58F3t4b3fzlaO
K6AzDbrYH8rZap/Th6QGAMF1arQBZnTKCT7XPxUl/7P+I67Jt3f9staJGdwWL3/LyljIqzaM40ml
dnGisFDlDokxXbzslfoBeLjPe3QbUo/S7Qsy+2g8tLtVrtq6YmtZ8isOMiReUPbZ2RWxuoFx0ch/
X67/CM8mnkMbSjbE3GcJNj7r6vp/fqsF4NBuYMnSscabiw85bSiJ3JZdn8KiGsrShCk7bDBtuzIk
cGqD2Z4G5k0DZb7f33JpDtW8FHdGOIVbhOMSkZsJdXJPBaETgXHpISnOjrXmUP/KggJoDMvoKU+7
3IVzf79jMOZkUpmkaVdHc/vhEBixDr4GfAtmbMQejD07ze+d4AU2gKLbjnXS4UDSOt8bp3lvpLli
funtS2MM9krbVh7xRVqFbrKiwAA0kT+64UNEibJzQ0fhgEQ5GezUTFqjg7hpXqHZb7gJCkSKJQG4
SY1OovbL0dRu2YSzjZthTxj7784JUUfu2JGheOgBv76oAPhcDvm7HEaoG87ntLp7Z6+QqrA0rKgv
RLqdU2sXb1sCQp4SS/oiNSfEDiP7WUkH8Kdeff899+QOP4ba76jaRiAGxRRg4Wcq+/lkD70nO2tL
OMmwCNGf5/1nxOK1B9OR6ra6kF6V6q2Fha7nFlKu/zJ/O06SywnaiJUQOYrKWf/LEoLdnCTrYMVT
XcTkO2ecJ9VgrUoNy9wnDCt1wmUR+mAwm7RgVSDl1/pr4VYtzqcEY7PVRl4RWpSrQesgIXdb85lf
R5HP6MMRElxIIeu6/aOg8+NRNWzDM1+2ZXuCLxcxb6v+wXwDkkxVaGhgDb3OPQ2rAo9+vGgjRS1t
EMKdva1UAj/R66ki6I/f/7ubVYdfaHWpcTCELLFHgQKRZqbNoi+EJWwLhFbbZaRowRw9u6Z+cUrF
3PaCTpHnu15kYIVdVTkTaxYa7OL1tLkL9RvkqSUttOd02wrUyGLzt4sDbYh2eEstSCLPCXZpnrvl
Xv/9N8FL6Ue9MZG7pahQT4g6kl9nrklQYdgXNoECeJTIeMiyOxrdzT3x/AaJJpQPG8G+18mKqlIp
yZBr3OvL4m31KOv/fTQJWQfr5iwb1A9DXeNF4JTnww2Ls+qVjtpsI3QEMUT0j5ZsmE9PthlYRqRp
SJQva78UMTcvUfPxyCkJAW/05F22j/vJvLR1j/i8ikSsiEHppUmm+G2jZlZV4/XA4F+WO4+4LXjC
2g4BcytTYppiVy/DxlvLVE5oPcJ/KKWr4f/r5IfDc2BuY6D7aib2dhNcLtFM/3nQDKkJucPhs0NV
C5uAoecR7bpSlliHOoloUkZwX5+uzeDQIADV+EQMqmk6Jpxmrw2TmkNN4e6cfXx+Xrpz6styu7Ek
gl7Lxj7/4tZo2xDfVw1QYyi18t6V71JLMZRN1x2D1lzv5J3b48LsaMoyvn5G9zarM3X+k06cQoKA
jDY+Q5r0B/63AQjp+TxHLkc+J4Z+cEhVMNXfRnBl3f5lIBeZfP3beXZqZWwX4LjnePGSAy2tQnwL
HhF2E6jFdAMuus6UxANduytmzn2LY0b7PxnAmugD0+rhZKHpr/+/cV19buvfwfx9nMr3BXro79HB
NNjRutiWFxlW2/sg4G+8ZDnfub8nc+c2vxnauz2kOHuCb1iWmoIq4B7AmmWlUXwCTAk9p8IYwfqd
2oZBDDS8lLT4NoiRGM61TIajMAR9PKGLA1E36zrtGzIwlEIY2RYtV5Y45Gkue5JdBSJoSq4q8Wv2
mHxtlo2sw43zCUIyt7RMhA+IjpcSYKvNk9fFjVGnjn1K+AfLB91CZnE3/sE9Y16A+NyBJi7aLycb
zfEI1MiLGl6n1v4WLPavHqqf2EgGItJNTAM2vca3HrKIlkapCz/SPy7n+gshi/IMZaFMkxdC2J2t
XRwEPu4Kzg4ayXHJu2nMGiZSExCsbtU2whER+S/+WXq3Q3bzZFnvDxXPHzGksgEPY6LSfqwSkzGd
DvsdYdTRG2Ii9uAGaEcIfb2I8Uj//TVWWN8bCSb3tFv6L1BBrhORy9SY1zNAnhkB6+Mls8o0ua8W
ZPHVqmRRTxikSqiW6OLvOYL0IIr/c07TXHNdyMG1syfA78mNj8982ara06dDQ5X4BNhOIDr9sY6+
yF6t/6kntEsPk/k5ueitkTM4FhLFm/LkmsfqUKTP2T1/UcvKcmihcqJ4IriBu+scFV0s5KTqDdse
VBj9/4zaN1tuLyYvmcjfQB2yd7alveieVaZyccLvOdQEG3un36K/Qta/o8/Msky1C/lFr/rUdDsd
s6PijVOd0Nmi5O0s10xQYM1PpsQ9Zx7X4ATDuq3iI8JVSeipIvnT4h2Qt/zXS9QN7PIv38OahWy4
DE73qW/7C9k5BL41q+HLkt5LFIifUJxW5pRmdasreQ6bZjFqK0coJwiUfliSGd/l2QgrgKFHfWjo
LiiR1u3gdGiTp90Ko4ggk6kQnmTYTIYWmgB3wIG7Cqta0O+oD7Omyi6h90+TcQJ1uFLFRftzcyJh
mDEemEg6rv1bVW2ij4cO8BK6nrOscKQkyCQISBJfccQzWMMSVf2TjWq3FjYRVUTAMR3DiyxNkGp7
fl/PldsIYHWcZXaOJWqvjuYh1W/5atgtGG3s+NKnL09iC057ddCvpndjvO6PE1NwPt3oPMJqkpGi
acDo2kSCvWRMtdWYEcwtu/yHaxp3MfOM8xqfUThOvnkXBCQUsLz9lCpGeGTRgRFPKRKYRD8z5QaP
l97vP4cdE6FFEmJep1burbjgFvO/WsApP956MtQJDw8vTZbaB5o1Tn+FAWeOQCZQuO5TLuUz5z2O
1yXBZWZyFuIjNT5ySERGzkjjOC4BFo2JgyFpJWuULvBUz9fwotXOEo0Xz8MlosiEpvweA7SPDv5f
sC6zlPbWkj2dCTBQPhPLpVBsLTfRibKH3lvWDJMcZyLlS6S6R7c/mfhGf+iWWe+Y2zthtJOdlgss
tKVQBtCEl/i9k8U68z+CdqJm/tBqZTaHkfdup6LEYbc6Qjehq6TtEU9lIpvTAKA9XARNSlSOz5Nn
inFSLXBj5pL1Grudm/XVDDXgdxtl4VEmx5NZ09JvTLW7L4UDe/3aBW6s3zMXocAfllqBUHuLv+24
5LwI321WmVX1Gl6pZKOSwN5rbfB2pnTnn2pUup8IjDinsh9HxfdLtQQm1ob/WniU5uqCMgA/MR2Y
TkJ2q0Bl2kEXgqKzk8z0cgV5+tY7Zn92Zc1Nf4CZBgTVu/lbmtwSF17txbACOS4057Tvxj6qMIxz
wvGRTm5dRpTzo7RAmEiUrkfvQFGqR3knjE1XgeK9GgFcMCfSp1HVlohrX7SG35fJtGV75z6GmdZE
RuzI4q/m3NWX8gKS1R92AACGR05Xy1wjxRrktUuW8shT7jkP0c1pgjuBvpLopf3Pi61t5N9NSENc
k6RFq8qF6s86kknQxXq8/S/X52nwz6ULMfv77bILEi8WighaHwgRw26Hh6cYYTpsAnWBQaQbwhWu
nIq82LKAdC8dx8p1XpKJ9izoHlpKorb0FisOJQ/oPCgoCMknMZEegJMcj4sidi9FbLqiU8PqKCUh
9pHlInRurplaEKgRfd17REifg7PnJe4DMTJ0WMi4CqLHQVbC1qklMk2+b/wdWSdPWrJwtcxi7gzk
+7+XJEbY/MoBE8/GZIf9CaRxpZa58DxLMIZUeZaOyYfMmmPCfOlmvpXLdd90b2Z+uVUz5umKlUqR
sFD62JpbBHtVx8ObsUMuv2Nvq/A1P4kCbFvtwGtCIfeqQhvXBTmV7iv47kcGiSKP4Y6TDv2WGxHR
yCfQIIsUCuQvvopW8yFVnXDoz3rPwW/hjHyrqS2mHSCy1PchZuj4ziYGHb9ncP4L13Y49jYO/imI
k7aGPOLPaWIwsFaks4a3//hD7TsZ9b7jhGvTK1+JS+s000ct8QzABrmgivmD3tjQjHHq8mY3cQXo
2tPSY5gHNf6bNw13yKhB0i9xIe5ry1HT5eGL2ugfEUlVdB8FOtiy5fCXwil0T58l0TJAy6g1V0Ye
ZOG0NS5bPtANT3K35xnPH8uH9XsiIUe6hrEzl4PN/jHSS36yjac8rvSUxW/Jr5q8wal+D8WaMe5R
J7UqldDl4wBQKDAZ2T51klwviCem/++vp3EIqRa3E0YNqPxlTy4Fm/lBNS5nZnAB6mxftXIrowrE
WhJkIPsT3U3hjt9A22OTwx1FUs5JZ4LdDSlqMYtbAFawVn7QH5G0iD8K0kghiljoFvPFZvLxMMwZ
ztBZxDDLcH5Ds2t1kbXKXpdnu1Onrl8lwhfFHikjOrU1pwxZzvsxZC9j79kOy95R6/Y4eS/DMfn6
Qnk+Q4hNa0591jD1+LGyzGO/JoU89eaUDhrXBeEm1XvBoxqu3ZcLcFgAizytIRxw00XCnFZjaOFX
+A3iDCS9TZYRQJb/+V1FTM3tunUzeuitWP7azVfdk0LS2z5Wl7e+mMYFo9s18CtjlnN94oY7F/1q
UQ0orjmQo9rByN9vPVdJQZEXMOwetpV1KuZDnc/zgDapi4ZQKy0Qdz7pZHkPEksmqh8nV4rWUISb
fsNcpQFCNnurkxEbLh4ZfIlU/vYWxANwtaO+8breTAlVK7a/PaS71mmLdXIoK6iueZwnB3zbhKU5
tWNQ3fLPtV7ZiMm3dOPY/TWKNB/VhWNRTQUO48X66aWZ8ONPxVxkRTzxSlshnf8xe4zNdnwXLL0N
6kb/29jjr3BLIDaW7MkmMM+CSWq2UT/8Th8l2AnJNrn8MuHf30N8iSCZPRg0oZU/fl9x32oXR2Yf
f2t/vi0C2PqJCu85GREn9jDODwMw0no29FixpIrq6yXPrWyVPYCsZUpfCot99MVwrfLHTl4WZO/M
fJlKI/o5wMQxthzlQZ09+fhlbgm/kP0jaa5G5yrRPizjO5NzBwMlZusfSIW7gTVGdUJ5R7Oq805X
Hb2FspsOqX4Q4eKpuenBjhdcxOrNewrtWv06NSHbD4PMWHG0QvoFwzXQNIS0ho6iKfsqD13ciBqA
m8wHIJa6Oj7rvtYVvHfP+du5OeXll/PL4EetgzCaHXQYP2TfDZw+H/aEwyZ14ZZl/OuO9LZNo3LW
d/tFOBp3NVJCnga1A5b0mYg/e8DowolhcIY0nv3hmeHNj4meEDXmYykmUYJLuShu+Yri6JVdn8O1
SqKtl/OulAvC7mVpwdsmbrPcNiNPGPnTBrNRmaNmAwyV23CvRrUFjZ8BP+0bkTqAT+/hqbrGWVK2
Lg+72aTWgkvaosVTFW71XePriSZsrrFtPZvJ/0Ia9+wdjtzr44Bxm/RfbMnVMpSff3S1H5edCIja
EZgdpeZpjdWCjovW6Z+wDatU1eUlnqgFBc+CO//5IWX5Y+l/rCxJ/+eMP3zYyCx1V2nSuUxG9ILd
a6PPT/MjhCCwTHOwquWG5CjR4ZBCw/pAAIH3u8QJjn9bIIGOvVZbmtG6EcsCSJzc63Q51XK7L7h/
vBuCNLBZos78eBdc/JN4a5AN6lZozSmqZDqWVjK/ULc+9/mcc4b61LosXy3DyIQFnvTg9bPmf8mz
uLscQt8ENA0SSOF7k3yE82bCkEyGJ8hiCTzYx5z/VqCOYRp0krakJUJ1vlORhAldWs3gv4tohLh3
s8HlnNPG/W6+pjpIkUejU7OZRV3DB5qkb9Bf799TfOUbsM6ihFp61ANPp+Fc3mNN9W8Ie38gAi/8
frKV71kWqXt0gA1YtrUH56gx1GqEU5R9a3GzwbVDv3LMH3wIHsLcjniJH07ai410nsKmMgv9rJ/C
K82FY0AzFDktinn1eT2wcXdsooUWmZ1C/ynpOt3o2flZYTwQzckmwu1cMeledQECKd4f6Tvq3HBS
QX6Ux9tXvsjetqPqbZLXK4GmVQZ2tRaCfA+C6SYw8q6T4IUrLdmR7tBSPQuFF30RgCgEpuBxj1sP
PgqEzICYQVHfaWZCD7JRLEFTTDk4wr8okO0lcZmaBMeMfOaJ4fRqkcSTvqSep/p2f/oUBxbrObmF
Xyd3a7xmJyNrt3jBBwm0MUnuVS1QT1MjB9ViS7q2ZfkQQERvy03/hHKrViiouN8anwlGfxMS6X3e
iiHujUw9MI/tjl6D3W1W8JssArx+AnnVWRrFOLy2luIsxfv0mWZtOtxc7x9UGpPI9EOhdMHntnQh
gvD08Btp1IXgPf/1ymHjmnqU2aIcKH71bkjI2gm2wTaCjo2meOSNuAjmlQO2hi5V/s7M0F1g7TkW
M4UNQrTGPqbzAyV4JVSjNl54vUDj2u1+eMqbhaPJaClG6vQfcSFqUFo3vg+Ue0G/zAmCon5uRSFK
LaGYW489/IOWRTSc2VgxjraEI++HXEyDZHSph83JY+Z64gjJb58cJLWG7okNS+zNcmfAuBxUu5AZ
yhs9Ql5rTGFgRVhwlYVnZVzV7voNun6tI/bpJ2Mz4z0akXcKb9YSyg2yL+hkVT7ZgM9jtI3IAtPj
LpzQJ4C9GZPQWvLDs4IZ+aTxFBjvXu1uc7UV2q+CpLwKXfNUqv7rb0PaXPNQRQbyxLifdw2aQl0V
MTTwehc4DH5dU75bUi9yFyJ6eMjcKiM2inJlxLnVSAcnA+2p7wowI4pXpHK4XDe+rtr713+s0Kno
WxWOlIapJW15SxXNTVd1UPP2JekjffNqqk1DJx6z6D0/uRX1vlJ5R9oe/pkr2yCVJwjr77Dvd631
zBMpt37Wy1APXKIsYqEXrJGb7v6aERt8UxryQ89rgpTia+6v8DEIKwKhcLglESMUTk1dV1qszXLw
KGb5WvLuWc/QV1wgwLeuVjckgVsJ2viOxzxYr5pWtjQ1yqPS5L+f/Cm1mfcqE4rOj6uCXk2Ry8Xg
/w3s1der2rggUbm/ZCALpegMRDZ7XjdIxQdZ429G8dC/7PVZ2QuV0HR60VX2gC9JcKN817+8jWZ1
5hOCxrLFGTJvB7AJSImdENw72K0egrG//B1roQgI9qA8c5vXYuEiJEqtJQEmGIK/4izMDYQK+cUO
KaC2r2+1u1BmftAHAfy857ypz/279nxpvh6uCHQDUeV5i+mocdK9zMKH5SagYbmgeZ+Pth1jA4df
5OXrqPEQ4K0JNWJqD3blBHZE7KnZ/XFz1lK88RgP4E1uVjroEfzLPaWxNmpD2h1GMYUVncQlBFr+
UF2itLbRSj2QJ8VjUgdI7xqgq4wFs/lhXxFZhwukrC0Uby/VSqxNQ326fLAE2hII8HEb4/XAKR8H
qsSk3b8acluswNVo5Hme80X/5P5lJaHD15Upz9O5ZyERDre7SiZMjN3LmF7HmaNtQlKtv37jBvNb
mECRXBavOOg0yR/RGxmqfcsuwC/sq/FfzNXT/ETByfnmknKW5PINU79u7Sa/QOWR6QtcQXWIle9n
SbkB6FlMPeCKD0PoQT2nJfNWrgDZa/oYFIrljh5SenypXcIgzGl3cL5U81ZYPGXbLEHAoachud9B
7yI0v38vAduqd1strY16/Ljd5bD7dKKxM0BJJzip5oL2m5t9+SF2+liIfSiz8zYVzmV99cuK/DfM
COjSNzbfnklJXFk/ys9yKsJQd+Hh4vGzpYBsvB3XAN34nefssGiNPiVIlmi2PvrFbNCUVkTerDlu
shg8Q3Gi6PO0LZIbfAdrb0JjH5tJJpMnptLBdIwO9KQgkTWaYkkiJKzMx6gmsOWDse/w6q9m+khc
cLQZpW233TQa77A8a18tQxpRQPDgK5tnBE4CHB2OuqwqmKKYfZKUcU3RgB5gjN6Z2PQTe5asYQRT
SpOwQuc+ypdje9CszQLWgLxNRBLt7d2+I/mIc4jtqn3aEXgZ+rIPea1H8gEwCvKFVM29+PLGVM95
C+eSefzFHiV5ns72ZgKGDasYIMbrYbWSiRrlQfgb0lG8evn5ChiFvEc7zhu8rd3VK443WTM7gTZe
WBIg5C4CiG9qcYbuURrveEm6zcAkEm/m0xijpntjAJRgogssznb/NAXKqCxLw9/Blghkchm6MZfX
YAGD4/fAHEjeq8mJ8h5iJlV1lVdYVW6Cjz3xHfqsUACfx1lNOvQxhIzyrjaj+3kLFx3TQpMYizPL
5ZmgZ52ofV6ly8neIL6+cFTAGeOaDLepVz/TT9iw940/NQon9wfJ43lOZEAtHwWb4F/O6WrvO4zR
stmIAEAYm3bsmr91N9MZ6UsA58/TIPyNDDX5FK4FjG1Z60Jk3EpzhWHeHSJCZFXVFCVQ6zbB2XPg
Rj4CGyprgsUMOYSqbrV8H580yjWWxdHBvFNFpQQjouKRhjiJjttE15ysRhjzU2g/JVios26+7GeA
DpCVds8e/M07aMbBl0W/n6x+WK9cWhx2zGavn1lsg5WNrLJiql1TH8sv7ByABPBzKHI6VHkZDEOQ
MPAg3WRi4ts3qnzy6ntJ9ZATq2HbW7EoqZbUX47AmnPqDeUydLIrFb5SvUj2QOJx2Sx5oKbvDysl
JxAZ0oU0CNr7iedAwVPRxs/P87PFE7/pfvy+OsrkUhvO4kLFH4dopQcNWfRtJ4vRJf6V5We2cN/t
TAHB73FA9hhF7gKuR+dwO5U9DbFLbfUKcYOypv53R3lb3iSZVNfU7CZmltVx+7QqkiMU0JnR5tZs
u4XDw++9iFR8IjuK7SVFY2HNFHTEx9ud/bQn7+xePzxGFaE4zxvSnIBHMexoqSwLDgqCJ3OS6/+t
XLUEgUxTbJkJ2VtAzeHOz1gM6IHycZi1ii9120639n9vzdvbX6k+7tTUv8GA8Gap4arRWwrUSoSM
zdAiXjZigfIZBKxEH18LDGxXZoeRjGIFccOATN96vgqrfkIxRBMTfIEfFK35tX+bi72j/dJ2xbg3
pagII0QpayAMi6LipBWaDVzC0eN7dd7lxfjMhExFDhDwE6tsKyVid2Lc9Ltbbza7/TFbLQcVsh3e
WCv29AIdL8yIXZ7yyUQ7fcnyAusZJFyNco3YkeRLGc5WJ1c99QuTdQYa9Y5udfIK18u5yjL2jnCp
vYAY/EMQELHvlokXvws12GPpi0lMj9pJPWoelmrwXLRQK8o/XvIYMkDk+OKz8nn0wJaw51mhkGhz
KKU+0OPlTagUApEyWju/mySSnZRk9Qzt0vlcMK7uHYxcMAkQv7QDXuI9mBq1sao2maFVdFk/bxf6
0rp4/nAUvDNZj/s+yujrsJf0UtmcGKnesXK+Ugo6jb0KFMSxYHLGZ6BwmfQ+c8WyczMsw6qHI18l
my6ONFbGg8ZA8S1Qwlgqq/NQalUve6DpYSsOGHYGX3opnTv63N95/BovUbpdHhG0dB/MVmfwPW0j
yYPuyyyEzGRJUswxyPGg1Ff5gMQptE+Ph/MMwQDA8Erf/YWMEzAowUIobQBYgxbZfn8bwzQVDT+G
fA83E2EXy1TQIEWvBRrl5H2p68P6T+2nJb+mfL0lOQgzxzLb6o1c49ZYXSPqQQz5C4RjpTs8+nT4
bdRK3aYGkoeRjEtx5UzFcG83aRzjxn5gELp7elrhM9h05J7EBRv9ENzyFZFa0dCnid4EuRc0d2gf
Ez1eDja9F+vLu/AWwr6fOmNGoIr4w3jKi7UgIcMNvbG1FXI3S2NwJnfmqaCYyNIB0uns33RuxhaZ
EzJWMAQIrGluI9T2XhrqpidIRXBNB7GYqDSFC8I0b3Gp+bhB5ROT89RcfjojJGPkdn1eBaefmrJH
19uau671U4KHD+4bZTKLHX2Zj1PZSjgGcmBz1CnquSdnKF/KeEgq2fYP+BVJI+VgobP5ciclWmAl
op3EPp/zMB7PFR3lJy4Cixe2jPciBpuGgAhYMmZdJd8lx2uUlWzajILcJ63PydNMuvsY6SCOPTbm
ZGGICzWT8iVwJtyJjPS1UUUXObNmFpLJmGQtBMJRpyhVcbp8zpnzCbIRpscSCvycErlgvdlV5OlR
eO1qHF59SjzmP099w0iXVF/h3jKvugDQ7mbmnzkn4yxisASjeoCZ59TYpK0d82IKAzXDkWt/5fRg
Pl+MyL5ZUbYIxWh3W0bCKvjYsvtIvIBYKbrQIYf1bsEmJp5e3IvfhUgmoWRX0snlXSg0P3eMjpjq
+lEj1+cAFPjp9H+KR4SrxFHuk4pYMHqosFPZuNiIQjc6RXtTP15Kpu/NAk0bE4UYDS1dDsl9YvPg
B7V6L77iv1vSQZAE8LALn592RsWRRetBWlwsq2sMl1X39c8+9t/SrqTbO9WVI6vpP6F4jFFhwFhP
dsVXlJyk5K/gbwsRPEaA3Vht+h8/8ijmZg87JU6RnA4Gxk91aumrOrWMgBKmIsa/aSz7SIRcA+Di
rcofV14xzoqw2Z0wUEyIMQ==
`protect end_protected
