`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8192)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/Y3
LeD+qw2K3LM++tksXDWlRgF/znF+Jw9c2JQAPXKM9TKRvOl/czmCOhE3aNSoCh1FUwlKG7QK7XW5
1i+Y/6fuS/CW01hotPrez34/+2hYr87se6GBDorysLqVAXMsLY/YV9B7HhDUSw8jyNyknIEmI3U7
WudHo8vhLWlCkMQkDcMf+Ivoy8TEGZRjbwDtOXoE24Tpyh0y7Szqp8vQqEDariMqKoVn6oTmJYLq
2DpWhIEswln6tRI/+zBSleCqwfAdmXyYA/Icw782kOJqC1rm3rVrW/fPVK8K9QJVLjxlLtCOUsdW
MXHfW8zBcf+OJ6M5Ps5WfxcGaSo9F93JhZJwtp16qQc943Z5uL5S7F6uhx2/2/JNEiZKR4nwO6YF
9lApKneiqiV4lMknv2GfPf3Z0yt/epCJ1D6rwzHUxOS1WE+QGHCe4rtK8iJJPU8gdqWBAV0E38zX
DrRSC8OcTDpaHRsM4h45UtUZ7QHuncOnjyjfle45UXlGJHuJmqtQtKoBHlkWLaWs8IxPTRJdashu
kUk0S37b7qinz8QPzVNDizIo7tt1mrqBCLYTAlFjqwSpg+Q2GoQNpEbhhjJSmvYKPuGddRJZO7Wl
OSphxyLgZzVvmxDSH/t87kHgGHsFgjp9dviohojl/U/zWNmgRey6ALjcz02ZkQE6vzh/zBsU36oI
1XLzZdPOsmsFTW+hi0YtW4QXrws+XJn0lDvqAm7a/4zSUan/YXPqgWJAp0UJnu6AAEQbDjLTTbka
rmLtzTc+KBM7Qh/MrR0nLXOt+vB6+4vpyFW6VF57FxmXcsdwTMv34b7IGNAHXV19xTd61xcwO0FS
hYiDkPuuZYyI4HEIp4JXLUgW5zvyHVNvmOFASRRNUBRiTkDYHnHp7Z/O4tBKX1n17fF6v/fg3mwS
2JeiK4If3PXvktkxXJaPGyiZmPmt5A4Bthy7HLbet//JHNLV38xyJ74gKq7QU9oEASiPXGEAhbM/
x9I7SkQ7MIJFc8uqyxac3MnFNurIiDEeYdHyaMERPao3PN6xhb/2oFOdOfTFP1ukLGNEUsk0hPd1
LgkUtfW5A20Gbm2UqEhuCsZlhhN713pRuj/0GuH8RmIBQvAjd/LXyOWfuP01wImCTKOjz7332xEc
vYTB2ZLyx0dZNiESt3YthzquQ30BRv2JZ/yMS2L3RICN8EY6volLZIQ9J/ZWNZnto43SN9PZ1A4d
KcVhHcitoNxEjWlorIlUHZeWcgjrKzRKTms/5Qvq+XK9VFq4xnGh7Oac9iup4UOYCOq/mhqKA4j2
JlpoYNdiV2q/qk1GYiR9lF2o5Ecimhm4F6Qr/f/9tQ8wUUD6qfkiHSEpOGq0Z+43W/6hQ3pmdtRH
CP6CKYahbYpyAC5P664kR3KSyU3BSn/mcTnKBa/6NWGyfV/dwudwQZYVTSGWPphViyNhg4NXBZdW
VpNjfiNyjHV/WD/NL12VW2Cc1vUJznM7Ohc7WOPoxL3rTVqMbdkgPi1PL7rVXfy3t8gZU9LEOkRW
PzJtI3ekd0GtH6hpTLnCd4KmXpUwUPsqehrqFsbkKH7YNuki4EFBpsExEHrPqDWOzpH/kcA6Kdrc
YH3a3yqe7rPGOTbbq8kMXtkWN+YItZVlgy9BxRaEYkXkPwPE5k9IeceOrVP1c98Iv+echFZLGGt9
j0QBJm/V8zqFl/WSHqF+eE2suXsp689eqNMH9JYhg2llYDoxhhS7WHFNPfDyoEWMj1/FlOG8ECsl
8hbPn81Rxh9ZGPDmnWU1rLYxp70uYzLoDW9knjjlU7YCZd0swAJvYRhXsXf3VpO1kz3iv6W+nZMX
Brg1+/LfOSXBphl/YIzzMLzLBGrPVYuVX6U60QduJlfeyJj/jsupLa0YCq10Y7+A2WSQXESFHfnp
Oo1bNau5NhQE2DlB0tGBKT9+EPIslfIrUiX61m6Dkfx7lrqNHGsqror8LWJv4D6YsANdMsKop3y8
ywyUOABWxCDeC4c0Mvj7ZXbQ7mSXzmcBcrunwbWP74A7PloqWvI7iteJV7lKc7ctjR9u2w96DihV
W/DwvdUVHlOVlxCx01PJRop9W1LKbTZpY/0ZzTe7UocPsy/89bc9AcwM4aV8BP8oa3Tq0MJrZOMO
mP8yNtdJbBItrltMSYPKOFrGF8h5Z9v2p0WPw/sstYnkE2z48Rw+6hSemnVMd0wzek9T/E1AS1oE
ZrA3f8QL4jIonmJyBqQNSc2KVR9ezwV6djyk6MGEmqbDiHCADFai9EZ365ggEep82nSHyOwH7e7k
WAk5TUhv+Z/kHNdp52dLfVakxOtEHSbneCdm8hkeGJ7HytHDkfG0EsgZqwM5A1W/2scrmPjhfeMq
Z5gZil+FLHuqDgpnlqk6GwlHJoOLR6TnOa32UQ4VybJP9TMmBagp/su2C8/eaMBKHBuRVk39v7FX
8dhO0ZLg26Y43Dp/r3gPiA1p/bUv+HokNtQflnLHrnfgcNwAFuo4ChGQr1suF+/6MEZ39+YYcLQX
aZIHry63MB6k2POVKN1jUp6i5HvsZkxmE+SYqfeSDdTzqzoy3kdlF3NsS9UON2EiPWysa2Qu1opo
tMApEFghS37Yp1yaPg80jFeZRC2laiYChE9ZVjVUsteBxyUf277ypkGtcghPr72TPqQ1zQtbODEV
01nBZ4KzeBhaYwC0n8+Xh271Ug+NcvgaVLmitcZexDBHRfooei8SXKptlrX0Oj+5f74mAi29Jmga
Yl+J4Ze7y68N+bzIJgr5GmTFfbhcQWOQtM+BOeiDagj3eW0qeSPaLziyW5Otu/hbEIob2UQETk1p
onrFt1MwZK1hw3fcZGOjClWT219Jhfuyy3lsb9z/1Y0t7kkhyoXH0NKDKRuDurkJ0bKhY+0GCyGQ
H38L1GYASu7gN5ku/Zk7VkFeHIldz1l6oisOIKm7UGg0hicb5B93f2Pf12QemWqxMQgJ63mSrLMw
CMUPup5rmEJthSLRCd0m+efD/lITkA/qABvGqeEsm2W6wX+rjFgawIQ20/6ViV26509WcvS/07vv
ZEnU06vBNcQWyIbp5E0BgSx++97eRQ87fAvM0gXFe/6+lnh93OF4fA3Ur6NrvwNsN0VAku6d6bUD
Cit7rG3VBjPMNuFuVQWIuCLBUjf9/npcUtpjl0yD5DmylhnFpU91a5UF6sQysXy8w4dnCA70bGNO
U2RcjxWWqS1XpDj/JaOEMRAHyAUCZmQJ8h02f/A79Ec3Yv2KBu2fYSVGLYP88gzrb4+pqpzaalCL
4NCC1qhNV+AEDzF7cfdF+R5yMolkhoRqv39NTJ6Y6mY6Kic5x6wH3ZIMbIei+tOoXean59GwAB0l
LUkNEa9QZ8t9lAv5HTOAS2/Ci/HIhDB/tHYEMbkgkpSwB+UqeeVCstj/ZcwdNzhcm6XqH8REaPo9
TFNuzi06rbpqqoJ/S0MbWN61cukZsxlU9z4DichFwolak8AQWAA4FVFclHGAgfoxa6M/7WcXxZOu
v0iiejWTZEVsWwvwd+5ILhINtrI7goVh03Ln0h6/cfzlMGLK2P0uVe1gWQtokTH4cN50fOWsVzj+
tvdUwHiCFdPdmX/wz8gZtFQHOeHANn7+KtyilW5cP8FFmQd9V/W4BMfPi/v55ThHGssqxorXln0g
EBJP3u21mc3WPjQtFNFHVGrtzxCkFuglP+wwlroPSRxOma3PfDSQCil/QbnrgkqpsoIY2NoT34ga
kSKvygT9DOQ+HYErUbibX2lXeYIBJJ/R3b71grZElbYoKV9paMsBr+mFOYMLCaVqvWjYCGiIC28L
pOnptsgveWobA3dUBRQgLnNkRv4DlkZT50p+KeeXO7rhyhRrB1+3Ipvup5rh1efxrtyR3FzvtLr1
BXnV3hhNRzRRhJlgyQ9p0XeXYtcF2dNPul/J+4EH1QJp3gitvPkcC060+qzuJ/buvEZxtNhtWZit
R4TSsy5enGXxZjpRRwu/r9aHnEjlGYif/Lavj9k8TA6TjfvEJGjaK2HY35oVHXvWEeW4dno8EUz1
1o8yWUBg++4oI52y+j0gFOptpbuxlVcHN4e/YU7SyJ98TDLHGoAbVd7MPOWjeCt+qUVLra8L/oST
jwE+9JO86bQ2WGdhq59y5WzFx1ifEtjyEhlEeRxIUtzVxstunOLA53+W695eHMMoKu3+Zg53JCuo
88vsp8ROjjTkZiz6SzYcJnXR8OIx4CXqDrQWQeAezD6X3ELWwEAacSkD4Bh21+lu2qd5NspGl9a5
X7o8ao79DOtEu3KWHnpmukTgxKGPpp54W4cLj19p4ae/tpMHXbuv2OlsLCmDaijbQX9VuRXUWqON
JqaalNfUPcpUr8Asniz6qD5tRq/uRIWnpEBvyhh4TtVQv9xO76jqSMCXTMGqcWKhhw9vTwdm5qhi
2/kDUBEVQJtAb7nhZjCEjMvhjevHGhvV7fXhYrP9iRmKYQu4/ULV6jU6GKBZ76IZg7gbolo7m28l
s/C+FcnOYOqo0sEFS9smK6bDqWyJROW2mCYUqCf4oaSa/y8LJm2FlTPiOAII/catPFTvIJT3+AWS
pSFYc6ABLp9p6mau2VSbSLMfdUN8SErWM0lBoINQsNC09okfW30HxICyktLZGLoQULzb9a6q63sa
yJklWDHetQXynpKMCM5K8sG8fM/t/l2tW8S17CaI19PQTjj6ravdorHW3FFiGYany0Mr5NcbMg5K
V3RCRfe1EvPTuVBgbgtfkMs1bQvJbWErB17caWZ5o1D2o6S7oIxJR9yiff50osuMSEhIu4fH+rZV
wm9joC8hJYb3240WD300vguATRyR74CTE5C4hF+vVuCRNfzaIMfoKMUbemZcByRQSenYdIH/W/yZ
o679XDv9mUEhgD1Se0dlGuh1PK1y95lEaseO1othrkmgkZsJvNZsRfFzgqwxMNPFzoGLhz5bloP5
VF4rxCihRQYvP+VVnbwvXWHagmX1PLnEYxwGCpBSTmtZGs5ftqozIuNYyhiGbOUawIK2Fqmfq9Ky
rHTEHGg4CHS9XvhpE2XnAgW4WRXt2B04zFw54pwqPlrHzLiPEbCR2Oi8t7bSooMCM2G67c3IO6BQ
BdwQVShUgGFjdbNEbnrb+ZjqmhPybm6jXEpmkdzSekytemv5AWQQbjHnloqUAuEBerfbXTCFJO8x
MVw7QJUvB9WLRe57JMTsxn0LeQxFX1hDWcbV7IIT/39O9WXTNs3xGnkwliJBqdlCUlZ6DVkJeic1
5QAH52Vzb+fi8FkcilFQfea4LvMJfMyAzGoHu8XcU251Mft6hqUVvvJbHsxqRs+F+b8c2ZOVXg1n
GTt9JgcCChcsPFkgcOKg5f2mYZzWOgqXoBGOJkgyEbVXZfq9JpeSW4FE9S45AFYza0u3wygzWAFU
oXeIL1zCdbpjcsN/fxen3t9wvfbPCLgZd5xxP1HMiYMqDaZVYEpvOzwVx5QrAoU84i1ozcAe35ch
7S0SXfAt34CqLluFc3tuVS8t/J6zmGCbjzKf5GO2qV0wxlJcr23RhHYiaicFMp7KhnFk45I7lUYg
TkgsqLFfLnzAXiXYPPvBkmrTLYmTHc9rrkhmTjskK5v1p6qltKVLhQIcNL5wNE5cOISPfJp4WcXx
+GliZ3e96BUPoZdtmPcr9NkfbnBVP6XrQjrPfAw6EiyBMDtsspDtaCJWXlb66YNbxw9pIlQrtKfq
FPMZhdGe6yntUit+bzyIf0R/1388UYOAOMjE4YBe8SHIAohma9avNnh9pxGm8Jd9LqulrQc5vh1C
pNpgz066l9I3XiorFVC229yVDXurFow+Ujk7uEDwMLpcbXF2bVBRS6XSYCIMdFkTnzHjF/oCcSJy
4hflBWhlhl+n0M6A1/VQZ+txvTSHC8Mna+HsiTI5suCGqZvR60lbFoqLmNnfu400uGYp51blCxkJ
856JSPCEGCveUVNjL7qxETeS4dbr0qFNn7/B1I9mRlWrq5vzhAlHscYygALMr4vmxsh80D0cOciT
WGBfup3bZERvPVku4cNdIGQ6crYOQ6Cf7zWyqzuw0Wd2BXrvjDgvnUGy+MHB0/357TrT4ykAO22X
8wzHD3A8a5+zyde5pXA1mkGE1zvMnnAUJJRK5HUER6dUowINZeB91pnz52btbwKV6BZEaJOSGBU6
eoFu2wT5EPGhTXauJi98YRaB6jM77RjmQv3JcKK1+Vt5sovqR0soCeQadY7Oa7pnmbf3AhI41F7S
hjj10vkdDxXN8ugloERoK1ZolKVK0SI72+BwnZ6PlV/Hif0dqw5fMlw6POidefSvpc5vNIlNJH7C
7Wf6EhKmA7ao4lpohcZBkmVWm6sPQ3Z3mGk5QUPxhFssxEvjIX95yBSIPk8kKe1zjUtKKW1bXNsY
uOuqrGyoheFkBTVpMnLq2rews/iV716MdejY4QtdAxA3Gj0K1qXqM49z/UGg9Bfxz+N7UV81CDH7
9Km3M4eW/qF3+bTWw/mmIZED79jVVo5vHxfjZP1qaF5vkRMwkbE0DQ0vRmP1tVy+F2waeKrdKxNN
2hZUmIJo47OYiw8xFiwECok0VhtWD5SthzfuCKtKqObLPabrX0gJg9UYRaaIvP2gOAAKeYrfiLfv
4TCwrybxmSCAK4QHS0OaPBRFjjWllcFzw1FqWoSz5eQ0qU0D9zH1HT7qJ5nZfRiQF6trYShaHl95
gpHyyNknpjARVnjoWqPkOW4J7JbS7TfVwzbyMIFODH26LhYcOPr+XWdwYjZdXhHW3qJuGlo2WuWl
9apXxaW49w2tkzUk0GRgL54Wl5GZp9KJhxS1pI+nbjP2PvoXBCJopCUkOKFI8xjqTJ3wBI/7E6pY
nx9MPW4zPD9uLeus2PQuA3VmsGRsEVcpgpw5DAzPq3GmM/hjTWCBf1f6nOyYBEq0/wYPqyJJ6iE5
9kT0nfwFr8hgmnpXkjwkO+iUI78jo5XIkk+OqlhCfDJ1AGVFHDfPHpVvk04Rj/ISmC0dEj/ZEmBC
bHpWhb53JbXDm4FjoVCvhJ089r2WXU72+hLVUVMAUkLVOxaUgWs0d85HlG/1dM0xVoKFg/v0K3kd
OJGPhCzt8AOinLGxHwpi8gzT3xIltUm5CJq8ojlsR3UwofQxttL4awjzhgIfLDNb9ggGfgpTfTyN
arNaDrLwvsFG/9FeWsRnj9itDUyNAd8KVf5PkwiJocAy3r9h/ofXszBAPkoNX9B0HLoot2bWAxL9
pouGsID4hPk/LekEPrj9jjALrhxSDLA/JAzXedHoX8TgL9kpINNr0VGCo7tN6JWpNSKMahV5AiSS
0q+Jui31jxPXunrZWSx4W4LaoH882HzK455TkdgfV1kz0zhve5KmOYDGzPbRXLPDa5dDJEcDajw4
J8IOl041ZvF5T/IQVk2YyGiJ0mfO16IFBWJYJmTpwwr5/iMCe6VfD85wa/SO8otSxbrtR9+BSXGJ
H4zkC2mzSO2blEhjzld3EEnvsZXcFIZibfyfp5E5F314OL8s9uy5r8fBxDugwYmbE061a0OOn7/S
enFk3/gtM39qDrtjG6R+SO7R2EtboLC2U1iDjYPHSUZbA0GmaB4te79bNec9sabtST6o5ewc2wId
9+oixhZ4A8auVuqCJPwDDelNx2Jih56gF2nL2DGkr6mLYrUvXqTjrjLYVNjxtWXxkE/r+UYNPs1O
fxJmx2plp5odHJvwqicFY6K/y3C3PGSPyd0jHQap1oJ8d4KU6XWSQHNnrLZD2MytIQ5m3rat7JEi
cGJzfLUlZVJasrrHu70rx5tSiLWtRvGl4ln4y1UwFyqWUYrOgJeCTs6/KqgjCvy6OgQbMIVLxE4e
EMneWOc4S1ypfeHK+sLO6VlnK+muL80O147qr5HbYwcp0GJ/PfeKQujc7jfFNiZwH1ILDsnKxye5
TEUJLXlMKr127ZdRIBsStakKXPxhooq/TXsZhiWE78tYuIQ/a32z8XvaF1Sb+MLRGeLnP1WiyZQ0
EEV7mGAdyLYJBeEv7qXSIsFpahg8o6qYnKfq5Xz/seW2KcO+djQMQFZ8r8uXf0X3vvzPcP6/m1T4
n+7mKGKfArZnvHiUtxJt3QVD5TDTEiHZDKEF7r+9fX42A69FHXpvdUuV3bbi/nuF4DuT8GL7vE/3
yZJzTZyxDXP9JZDpZdEpxpcvfkvsPs0I5N/BFvh4T0Atn+4VOTg9V2xMvPHADjdQ4DUwaLGv+wK7
OK6aTZMVs0lZjONh76Y/zUIZD5AX8B0uxRdZz2d8OzLWkdG/D3X9obAeXlFWJPlr69tgzSWoyXGq
/UjNRFLoujpluNh4xvfs67yWjMJIPwdf8JP7/vl9ZyU+jB+MLrJqAjRvaZdEAIplHd7h7Lt9Lvw8
oN7g/1IxElmUfyweEzZ1/Nt9D8sYj2Nm+E4wQPk/4YW0BewNS0NLcsBwIgvY+6IJqvk7D9VL6EhX
mqNX3l8blV3SxLBzorNaHPGoQ/CIiyL8HtdEz8L8lGUvJLlTg8hWQviC34q79Lb9YCNJa2s5FvcR
givMV6F2bDlN23s+IurwdwueWasHFgDGBZn8fzuqsaETHTnFVapClW4hMS5ALOHKjTKcOq5ovBF9
ZVDUkj7pZbRGdHvc4qZKNArCc61VyYjRkdQbVTQJiDMFOXD2Sm6XD+pIfY0JP+QXiyvYbNZvW0QZ
iqfTLDpZsc/d0kZXuJ1p+n6JeXKrY76xFUhHavr11eQsw271W3ewwaGCgaqp29UCCcYArLDh5HQ/
C6uvNDxhJ0rqbTznIa4Pf0Q8s+TArjw9VWEFu0EJRLldTZZIeW6JwsOmoRIOYJhLEL7C4Yp607Ur
goX7lQpfSHx11nQ7ZN0bdvs0dA/GNwFa8ZJw3Av49RWgNSTRLi8XxX5d+qz0Gf6TMzMVb1OJWuJx
Ak7o3ZYY4DJdKPd7HH6drKnocQ+vq/EumpSU3WPUWTxzxhwQHSKU4CTRAjfNg9m2y7betz2Dw5zC
GbE7A5n88vhGh5gro74bcjIzhKeirSm6vxro/dWKXWx5jdlzw5kjLjyB9MfOlEih17pufIucoEII
O6zWgalqxKMkbTeRY3CEdv4Mf3/y8sS0oMBwQ2ypAufFp/q0jeNWJgiP/A3R596ArhBOgEMJBe8e
DmkFeyZe5XzYnY5/NhOUHkxjkP8vvmCoh7jPhvSUlvToJ0JeMHPMv5rINxM+I7SzdbZELFyAfx/D
IAsotOUFGRFTw8uhOQ7g4tRrzDMXVaF+Z4RmrUNq4VkISOR6GdGZ2/OPoUHNC+MpJanC97YI5vbp
XV9KCtQZC/UnBEMcMXuV4TvB7BJK1mE2UIXOXcRqA4bLZ5dNnHqA3CFWUk3HDF94GP1dA1G1Xblv
W2NnjagbgrpUNgo3PBulbmDK3na3MFZNdyPIJdEqLLxzt6hBeCb40To+T3BM787yB5FVr59JqZTM
FGu7iBU0nASfQ4bqevt8S380Timpnec9uonz1vXCMp8tFTVIMKTL+/1zrAkb/ijODZOmArwpUcSP
WeXjxEB+6WfBK3kwiPBbN0Su3c8g8T2hTik0JJ2NL5MVhZ0+IPEiMx3D6AQgxbnZf9xnEEVaQOYk
gGwE7OCZdew+QG1daO3SeICFIM4v8dlH6CjJt5n9kt2RzjEMDBEeUPyLDC6oaeVfd3Rqhx6qhrl+
L5OIVAMWohFyzvv90dJdvC/CQuH++odCt5nY2Ehtw5dvnq7cdmrH0w0RVGce4ieEIBPVxm4cr3XI
4yiWAS+3r1WuBPFb72/ZR3i7jTLU+PmxnFzOCno8MPiAo8JR/7Yak+7veINrX+ltJqlVdptWkdxh
XtPWrbi/AUOqoh7a6rE/rNxWh1ly0o0Pc4O145RQc62E/CP3HYvXeFKiSKvPDhG2DCmXbJTADhUI
nh+2eOnDFJGse9z0te3f9eTcfAqIRSGJzDNeIZAbPkI4SWNTmMWACPXbM9jwdoXwDwYcac6y3e7P
C6SIN7bDMoGNGO25fxk1soUJiMdgv3cdqAYoxSK8Cxs5VQga7zW0twbSXmOz+7t75uXB+58G//Rb
hR/Ostx2/ghmu3pqZHbrVPkx9PxaJd0AcQWwQNLqHufDmLFEcSqidIPJYEPka2RAMXTrNQiua8xl
VnW/A1RKeqJIkO4gsEeGyaxvMY8U3+MYA5KrJuoEnhDWcg3sO5xdmScy6nbUB9K9kjr9vt+Tox3X
7oSX8eqFvitot0vc9I+XIYK/wLVrb2tip8AljPuWJjL8tGlzQSwru1HhAd0nYVmZHj0tRigPEXHc
Y7JuBpBXmycHoHCid4Q4Y81y9m6yuSLGad1g/fvuzxUvLk/jYy02qQytFS2UK06sitnDLZ3C7OVo
Ng7xWINKkH4BzxMTssRfJxYgirAFSkoLdQVcXGwNxtZKzQwJQ0RWnjWbPBDZqfkqcJ1PLql8mYv2
2TlAFW/noWf9YZZ5CVWKByPYwtmpNUczY2pqiw+dfO+jVtgOM6mqYSauxMEDaP/NiZYXouig3JKY
3E7V6Yj+ebPUFG/ft4smzFJd6wnm+2wMPwDddRqStH+eUIdjH15UZCEsy5JS88v/spMmK9jrrK76
F63sKXmRzQ/rsim3zpvYGMylHTuY40LsaWZqnl5sj9rgLHTdJEakrEuUmf877aIDLHe7h36N5naD
JE8bbBZBJZMSJdaRTfpoH1CtWn/QidlR6hNrH1itn57tnhEf2F5jMI9qCGv1aQGdJu5Nrca3TgvU
Ml41kO+0Fgh5tVRGGGOK0CoqoWULogWRlvNqFJRaqfDUza/LtggpQ0U=
`protect end_protected
