`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11360)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9TaBM/i2ZgCPEH+TSdpehCfiyRo
8iKS9ghH4ejmyvQ0cRxfj/4wEwjVfzJIVUq3M98XHpgzdzbp709gnnYBhuB4hLjzWZQaP5vodSgA
+/UyB5rnbHGS2qY6wy3tYZa2FFiWgGTnlDbwHpYhReYZLtkyyKRvgDjC5RcN8wvY7X57TVRp0tzr
yFICPtQPcR+5WftL+lhaubFcQ/fwA+lUlA34jA+5rq3euqD9s55KVA1km+DbqMR3Yq+TJYNcqCaE
2MIegVs0KLU9eqFfBD+2APgv4aY13tyqrP7rZoDNjRHtgX5DRAwNzIDD+MDm5a+EVu6Q5nEau738
oBs68vdOivlMWZ3AYJq1d987Pf5k8DheWcG6CPrgNaCy2oyooxNWUo85YqwauoRJeIxHTUugRQ9t
/RPbTsuSgjbcNPWbzOmi+3IoK07XnpFCng9b+A8CSNHl5jcaEUwQAt0YnWhtYQ0IpidMSm6+lORw
76wRJAiqebME/O6xT/w/kxtcADf2cCcDthpV82Xi73vS+mmgM5jFuyB2n7asQk0IVAubN8u/AEcc
g7juGYy5avaG17fWnDTuc2e4/dsoHvshHV3XHFNIMDVLWI9FQo+wgYteMvlJMGG6c4/FJUa/bNMf
FpwewzQstj0hxU5lA7AYpe7c24CSvThfvF83AI97uJaoCw+1ZYO+8Qi/zJ3fN8Vfm60N3NjZc3PW
3C5dzXWZJTNeHu++x5UW7sPN9YHsMMuQ5wTN/9XBDi1ettlwiTE+2CqiQf/Q81dzlvfOE6PCIlkZ
V/KM54no7ih5hXW6S6pZQKa9S+bZ9nAkfRpPNEp1d4JEg/xmzVdSweY23lhnSZHr9+5AyOMJXSuP
I3zcXBXa1jj55JD41MqzTmuXxrvjfvDakq3DWEFsiSPwRrRU7M5Bznsjn6Nu8Xdl5n7TJMB04lJl
zdm4rGu9r5mPMVca+PufQv0Ugr8ozX6jesadEbYuGLoYihSyoxDPfJMKj+K7IQH14AeVxp9mVbsp
7uy+/WjXB5zfjlJ+iMN2noYLFO/H75LAbP/OcIsBJlqV1dYLhoa/9b4xoEfhhDqpnNOAUqWwXjl6
n5TJ1EUhQBKWSZs3dqKRhg6l84iBL6wPUUZEveuuk+p4YPX7FmsJstAYzgHuC/qMJxL6YfEy8fSA
hseHBwoQ7VPM4/8pjJVOrSw8CzTm+ZTXtG1fUR1nT0iyLosnHt3o+A53c/YitSeNnzBG54u1wBcM
SNvBjaqrG4f90LEGY7/ClvkGSuHe7y7gP6G0aBfL08oTCPG7yxQCPu5/RssLoqHfB66SfWycHxBM
TrU1OK4oZpI/kw6JbemGKBBD7PV0RysMcyo9c7PQVOkt8aIiQP4Ob76hsnBahrASLJs1i97Klf49
NSXia6RZn6oEsD9Ae6ca6/m27Kdt9yExFTHYmFh8Jl6Xg/Z3EsEkSHFOzkrAuLd9coUXE7Gzuvep
LSFUiQ+EvgIPdLDTntWpVSyxTjlVCytxVVZz/Sej9H5uHYp4I+Au+LO6CAFB33SZ804S+DE84QEh
MW6k7Wh3m+WMVHDZUhMyna+PGxydeHFrbL8NWoJOLn8oFL8XXE4nNNyMG8Ce2v4ljb+M/K3ZCM6t
WqMQIVOPYFFyPIC2xvcTThNsqfIOemgp8szLUeveRk+FXXcb/N8Y85F8CpSDCDu3ir5GjhNuPHZE
Vg7FQAd/hqCtMZepcClUlEk5F0UnkPGoGLXJOY1JghtR3r+DEnLNvpaKaAmIGfWq0Q81lQsz4rOb
saz79NIlEUDFi3M0f4ZOL/CaU/9QnszYYGrFc7EIauWOESWvITr2zzh2o9kP7qU6RWcRFGyihtLr
mPrte6fLtEX6GrCtNLOdZqrfTwv7Ol66L5tEkiOtamepi9tQieTw9Xkh8IvJjcZACnZflClQRHjZ
+LSFY4BXLCDNGlwO6AULIP3bqaYbqPn8mXS5GLtq90Z588moRDpp7FgELy6oYOt+QsykD3C95Vye
QaSjBzqS6jGDT6xJDKxkqdIjmn9ZSqyQAhwwWLQyDAwpAgs/6eqTCLN9ro8eSL+vzYYD+P40hb5V
MLOBFLMNqUzyMCuoKFVOCHhU7r/K8KHShO3Jzj5zlEYA2Is+xMoAcFZvB0Ml2OTtdijAzmxzp0E6
BLvJCgcyerlyXBZxEcjb1+lizHt+EEzoJWkuqQtCJWqylhf4GczLAEVqqFzkxUSDyH3JmK80MfLm
OtXSf0zjeTbZAe/NVDkWY9xDkD/0UMteUNryKXM2UPyoGGrAnLwHCYYFf5eRE8Pa9cpFQH6ltmpH
95G6DU7ZoA+x8ko6wOJGBsyFx9WO+W5tXAD3gHe8FPBMuvHdBbxOLXg7fwpjLGeVUJrFKpaCSyTv
U/rQn4gnsRaQCyuC1rdbJf0/E7tDZFH6F7OYUM7mg8ex/XqRym2YumlvXmh/qXodm/gtBzPDhXyT
RDz2a5zcSNj7gIxCeip/hgrXJjb4bu8r1QJyzaqffFjsb1u27bBm2FEyFlmyXs4hKuZr+AqH8CJb
gHBehITtEzg2kH0lLxpz9+b9KX3blp8JdMXK83Rnn8XKpXOq96qQvpjp9n9Tlll0wFnHAYrdZRJq
dGnchn9gmY1oaMd9iHAXhjG1JaO2mZ63aEXWiaed5KgTE1VwjhC5QbGtXsiAewKHpt62sqaKVpEC
PIJCF4DP+vXbfh4ZY6PT3P5Zo3IhWjg0I/O/H2zcR9iGTbX5EMuWXLenrfoUwMftvrcHUhNRDMtX
F0ESQ6Ipcndp2D5Edrd429X5JWKIKwOCIJ/D9gAeOHRp7R4k7C+fp0ycboiC6zhXVYf7Qr+oubOj
XwT2v07JFAWvdkV4yrKobKwb916zr0ltLlr0uPVqPzxprGonf7WOGfTeWab/L1TbGcWxSmclkA7u
VYUh+Eai91n9n4ZN6KKIaW6bmsZfLyaAybK6PQat9274LJwrlNyVSBKgpI+ooDFu9P/MsGRxNOpd
GXmXdHYlnqT50UtqY2NCugA2Rs0ogrbt64jQsM96LmgIu9XXefGHkW6Nn4123BInomXjaosCLVZR
aqEmLqx4AnvhR4KeX1eYMRTGFNItnZI/pQoMbStK1JwD1HcJPLEYehQgLCDWUDUCYaM4/I989Tyf
Cm/kyc0B9PS4gWUxvVrsc2KI0aeS5HIghP8qtSXAHIb3T0vXJmgu/bR5T8pFLSDLfxE6XkNCsqYi
/bgHgWcsdbHmyXer6XE0wlCEaDKe0JjyPBcO9+MyiCgIvSsQPP+IGAZ82ufatDYNLRAfk4VbnZBq
UrvxU8n1QKJ+3Q6u0+v+dejvEQbbDZ7Oirbf0Qz3QoTPMOfSxfRvoPLJCesicRUy5klxfXGFdqzb
S7uZFF50frDJZCzfTSBOUuULLqOmdYPOHa0wi5awnE1iQNtQhfBviWVtlxvqZRstwOqf/TXc2G4A
XR0CyIiHolNtWxsJ5G2cMnx8FXIGaUgzsLhPevAdAZ5t9ilAv4ueT1/9HN0szIryB54eJhGj5KNB
jrhul49tgpylS9uggczP7vPTEmDfcySzLUjpJjhM261mgyBNEhFZmyUWqG1ptnUBieUwRuy+lPbS
Ffl0fpmAkvycXOFdp1wtLeb7Ql1heXMLVTfAYtPiTqNHy2ehzS2Onp2GYRm7AlP+hrANnaR0gX/T
0Y1I7WlrJh7Pgo04M8KAQRRZhvn5byh4vlrzf9V0v00oCfmioraktkKrtFU08SCWw0rRe0U0SqdY
LLG/IpHiMjqCcjHnjjxOlAOZVDjYhvH1/+Xc9z5OBsI9xNVaCDXsT4V2ohHnTx4Gs56nRqpqDW+j
Hx0HtAXLLlVtOqnu60m8Wn1mqEjLMtxZarDGMXiDiVHWzzBkQLWu48qfb36Ce5WF44IjLTLW2WxR
FufGYpi0jqA6+4lHxmAGUaVeG1ce01lOf8Y/mGhfG1uyNkvaXpQ+vFU9UOTp4u3EyAVBKfhe9e/1
HAZ3yCNbqaSRxUcJzXa0PB3NHZUr8hSBjeLgzNgMEPzqGxF+rG32C4L+Nn2W5B9W5r/TICDk3dUI
qpISaPYdRW20Z06tX8TfZBzgEaq/xO4AL1Uu77k0Q94u9Z8IG8E/5/w4NnZjPgrRCJfkNEtGFPF0
M68kiDs5alyCiDGWL5v4NoAGN9R4XKuGMJHfAHprsXv0f6hw3zkxXo4FcAhKJH0QolimPbL3LYyb
3nd0wzfTrzZmbiIDxCR2gv/nV0/RCbdf0oKVKLEB3AnW0QxP1iYbmXPKoKw2SFxP0cxbfwI+30SQ
Rgm/aCbxk7SMKsMmXJ8uYutulPvnUY24JkwjUTA1RWHVdvlbM08dGbUmoaZ3eOVuZRidxJH+CYQU
Gl2tijaZamk4hbjvztY7Mt2AaiiCjqdNmKyMfAOLBYyfdFGsBfD2o762ROeoIPxXgAqLboeVb5iC
XDvHhmK2AS2HXdcITsJfWMSpHjxgnRFviF8+g/j/KtKzsTpRYB6v0Na0HQCyGjSdmohEiZUm63MO
08wJBN7UsTFAP3wQiX9dYstF7gd2x2YT4dmRPKnJHPmg6kPwiZxRw9pkzuzkvRtkE9kEta7ChKQS
31t2jjqcdrmKugCJ+aIHLugp1GgxE8AmEocT/d0oGH1a8spEf/8VjcjVtTifkUfws0LWyotrfEzJ
s3G/lcCbIYQO9BHBP+/CV7oiyQZUJw5ooeGQSxlR2/A5dXE5c2eeB/T6aeQ4jRR8KwjdKXXRCPaR
1VwvDKs4XBTdGNnag2xrcXyiYoyALVH4orCnfnK9U4C2VdzU+QuY8pwXcSBw6QUqIEaTQO9GU1sd
OKy53ZEXdZ+xq5uJGV1efyfnnpWL6qlk8YvEomYK+9rFO3RMwKRuXVjf9giCbEeGb5SjCgOW/1Qq
kymH6/BfZfzop9WQHEUt1Q7Y/CyE4o7IbMJEnLjrVMFxl/8OO7pd+T6I39N/mJbUuUt8KC0zHoLU
y+aIIwnD3CkHdaLv4ZdLR6/Hmgp2XJS/8JQ+nvXhh2lCPWBewTWsE3b3C6JClmJ6MCF3q6bZH1F0
CV/mY7koc/PpL3pzInGIg0HSX99k5J3nsdgqlh6B0d4xTmdSEdExxKJclsazbuJFHErntJUNye89
fykgJgNyymPaT0VV5nH33RXhX0H4BaCqFR3xngJMDV9jNtLUHvMbuRkBD4bbvIDd5WFWfQfG/9bw
xhDE1bhHLxCOMEjsKvDwS3WQAOQDHGJBv1mqZList8ZdiBBlvRfvTjO+dKatgv6tYjkauoll8MSA
U4SKZIMWXsMW6a+IqR3bTZednNGitSYOSZSjGISG2KTEYlkFYdDABYnOC52cUgnrk/+j7euPsPsi
qHutqO89sqiMSjl/W4E3mToSH+HbmaBDMsAU9zyMrNgm16nPWANZxIRzGEXtA/ZL9K67Agu/EFfx
9vlKTsyH46z2g5oZXJPdEmk+Yw1zt8O9pAE1YONDEW3MZuD7hRKb8UQAhpBFFCqEqw4JWAakWaKL
EaNmwU1FY7llyBTnmNH1+02qi3ujD78AE8+rhgvpFQyDFiCM57H2BNv/n7Gtg1Q6NS5ZA2gjV5mb
H+lPT3+eeODnZ3QeAJ10gDlT1/G89XqqZuEKlL77tYv6UFF81cx9sVBIvmL7UriNFKAc5PQGcg0s
T+YwQ5ODFp2bU+i1jy65LSBk//8SNqMeyRDMTm34oavPGJIKII4zJ2GGFSpR4LhmWZ85qHFqNGjG
As916nuqjA0eeopV5EH+kK6PXlFNyIQtAAtA1rsmoQuBCNVkQ6R54vdaIynWM//MwUJAGXfSCw++
QO6xiFNt1TeCQLcQHd0XGwMPR2HWPZb3tGRr2a0I91PvO8h2JFg7+10NIMUQBOaWxXgwL+B9yR4F
qqtZJ4CZHQzPih1f6DYcezFxKkNkY8vDkAH914BV0F/BkPDtc5RA2LVLAyAMKGzhMUIQvWpDIohk
CUyyG07YpGcuew1Y4p5yOqYs1jHgrItNJyQ+R1sI0ZgN5iAR6vHTQClFmpU0Q/xr/RNQrhtUGGNu
NqiHsLHwAUihmxEHdUtIqRvBlnLdMU+47gmPQmX+UdjislLfsd88/wvjDQhYPLabYetU+Rfs0WRT
1I4U069qoPZepvPfSA/XrxDkbNLjyiMPwMmZa5LSSzYG8/XfjYeF7lFpZkxYRSs0KgEFXMB1icbD
ZepyZAxQmVLSQFTbFrMvS7vU2jiFSJkBA+IteOngYEVQzSK6qrJIYcTJjciENbzVwKRU5EuHdZJc
367OtDtN+ZPp703Y0O8Dvoox45ic/OxKwvcFbphJgfGZyZZuQrj/rRBD4W/M97opc7A9itdblM1p
k0uzA+FiStiocS0Kj85zVxOlQ/ok0Kn54GuY35wjJlYf30eH7+t8W8Cr+WczStnItwXlc69gDiVb
4AX8eGMtrD/Buc1Zy7Jg/7ClPPrizXyHtiQ/RYYwZZZOoq1xr3LJqz8p1QQVHYk4wnL4wx+igy8N
fub/vEb7YI8wHdWzXG9Q/NY7nwpB67lWr/XBPweLp0cb+GVppymRQhzVI3YZDzuj66Pm/+4U5mV6
ecLb/CEi6dtjLnKPf72BbRH6s37/xoZED2/yIjK/pf2IMd86uZIXmksJEaoGj4siKm83A+CHtjWq
ln/yt+xi6iykUQ5UxoXNZPyMji2LkFpyxps1/cgoY3dRm9KAMIfQxFwx6+IY90GbnNU9YFVd7R3D
4z0Di2ut/EDz3k9lQPHWuVUg4/5xrZ4ZcInufuZ8ttZkFHh5NecrY47TEmR7tY79d7GxUnvmLC93
4ybaIFaDyZYQdfVQcVXMcZYpJ/1o+xXJg+iXECaJj4JoGofF3UXZJk/ho0dFDsUTcAsXSv2yqJmB
sianl88wiDytNMLKcVOFBs67tD/lhL7DYqePPXp7x5yhTGzX+n4Lcip7T5grS4jwtEaZh7AMxi3o
T35gvT2CJ/0bW/8upgoCSsn9wVZ7s42BruDsOWHdwP+/nr3OfKe93Ug4x1+bAAsnwN5MfmpRbUbk
FbT0mjj1Q4leipgUHaEwXHDUicw6Wx6aawdATN15v5MJOz0T34WK2burvGIdWqr+irl0QM3RzXSJ
m2EM8mZfn8rH9CA2/PkHrQ/59ilKOFYfKEE7dq1fNPynN9YRClmg+HxZjp4NCjmfc1MztgwrtIYC
YYCIxrKDEPLKED1yzKruh7hGpwASjDSzWsQSN0FLDf4kRTQyiu9LVVKG9ZCituaeedQm4J2PtLot
UxSpCtv6pgwIysdacbkoZyJCJJbiB32UoO7H4AWRlD/QaVDJhtiTLE2h5QSe70t2+P7Z3kRICUwu
EQQVNgMmQP7L+MLLmoAiaLUG4oRC1Mmt1h3kCKl7O5hNEzoi0+2p0XWQIBAz/bSP7duSy4B7WUCz
YTMab/CZr2085cBW4seh/jrAhq2zv2nD/8o5T1ceiR9yjFujLnj0PjgLXLtU5hpK2XC0hu+JsozN
SoaSfbarN/TZ2aBhDwb+4ZGANmaUiLSvFQr2obPyOhbQAJR2xFhavadaGVhS/yzjRFhBhZic5DR+
TLCdnagiX7daML3O3z1QgqTOWSK6U3uqT/Tprqg/8I6DrOoF4YzoX1xVa7oPmY1S2s3pfinpakeM
OfUsmAqYhwWNZDAIqz1tXN0wNiCQMkLqVqIOStCjtqACB56HWNfUHMVOwAu1yFHZo6ISzvObTOUC
BsRFBw2IP1gCNoPsfXOREMv9gLiTprmYJ9euFjXUm6GZiFf3kErl5XCY20xJCv+scpAjcfAy3Nat
wsMOnIm7oWRPdnJOwJeBVVCBNTem+WYl4HwNbiOX55ynZ7tUasT4rhfETmqy+Kx+hzL3cBffiKMC
Q9dFcMpRoSmpiQtI4WSoSVjK8lBeetGgnjR7JaYq5cqnXconC7/SGpJC0nRhoDQ9paw0pox3F8pd
FO/S+9lkgX5ZEhYRZIpgrn8qHJWwf7hJLIFuBGhrsaSF+Ob5qvboOEfV766B15ofEiCl4tCJjMP5
SRgqEreNbOgxKqKPtZDSLKS3P8rJEb44EaiW3WOlEDaURfE8J4ln6xQZrQ4oFMu3DOaQclHb6Wlg
7YBZTeUETGfFAijQ1gotiQlPPwTROybjBmYHR8Fgx6tqrggwUhOgUJ40Lrlr0J6nDJKRodUfksnf
7G4nO3BQowEjliDyx+JwWBGR7fvazvezfU16IV18lAQtVWVS/lH//N5CU1XC0t2xqlwPueG2vhXg
fRsngQODLcFTyiSs0hSJyDfXsPMsn1ng08vng0X5B/XOJhKM+xuMpPffTYx9ZzG4oIRPc5CijKHe
A+IP7Tl2NSMaK2RDbZQKyaaRf0HvPqcL9ZSoPR1JHabZogVPXB/UKJ7QffplyZT0QAfTsCOESEiN
atE6uwSn7Q9i3ljGFlEZqzawAIFkBHZJuKst81pwLcvH8Gbfk58ulJezKR2ZIcU4YNQWXlK0wgyd
w9joRJdaUK6YKlPXQIsOvJ3dA73L5BDmoEs1ZHdLaAtnhWlG9eGYbH2bORpUJnmNBG3TTJ7rdJTt
rL73E6zhUnnkbAX5J16tTYdJqBMZw3ZiSMQguWdeOJP53mNAOB5ax/99SuA9/c+C01rLhfxLPFEL
ppAjdvKNhwiur3jYTBi8gTCvXGTi6506/cVQkajz8gIAxPHTMKgBjxxImnAcfsOTQjzbmpCE8Apu
3rzc8vW4nZ5wyC/Jgs0lPtnLb5mX7tgkO7TuaGs8ffsGioA/J5Zz08HP3XjMLzjcUmZC+9qea4aH
gqf71hQBrpzVOJKzlErzuSxFZ2izAidx3XE89uJa//4bAMf43ar9qukh/Mjt5+ZHzgL7MjmhXKiH
qdRVypxwuRIZr6oFfJKAVz1EHf4KHGos1rTwwH4K5SMU0xJEQlSbkWFtOvQ0SlBTBg6QAUxw1Qlw
yG4KNPHWPmOTEARaJBpi/6gUS4KRtt9vSlnx4AsXhJpYQcvfY2ZA7mVEIVX9wtmeytQbJuMRaLaD
V5IygKp7b6dFmWTXnqqwDX6hHbBCHTbq9GPVSd4b0DejMt/7owyV7UGw0XfVcHloUIUqycW0oDMT
CpHvaiPdzxisbpWyHJ+JZxsspWEmlmtX9f0fMJY14c4pl4xJTbIVOqa0wHYEmctCffzbXESxNpqO
NWseJMkdC8pzzSc3lRHJggdQe0xe+a5JA0XC+vU6F9njVNJij7w0R+GAukbhXQ5GX1eLpNN1eVj3
DXft0oBChXxl5cQrbNMH0U44etj1fKdiD7aqlaeWjVgMxSKue39cSuURM0iP8R1RP/IZV4B4U5Dd
o6Hm7FSxGzxCT5DjezeUkjeFW0beU0K5/93z/aubydIdxRaBkyleeSxoHhVmttrysIjQF25OOgHW
A7+QdROaEBZWCgu6yPicw/QVqdZv3h5vYXnYYCSooiRSVbt2gkgRoZ9e1aCcJmHsTDk+vbBQ2OLn
APQKZK7+p5jb9PV+tPQGCFOSygK9etf30HUt9ujSAv1qVRyp+CZhTRZTM0NljKW4QpZjjQ/+tVkO
9mTn9WcgnCyvHb15euLdKRTKcJ3LQSle6j3KtnglKkJpG8w6aWuixfU6vCI+fH/cztK7cz9BpNL6
O5+kkmW3U4KFhyrZkj9XntfumfkUbR6CE7vg6UnVRV3b6BTR5ZqvWLq/hozCQw6A5jJr+BlIJflM
7hoi4L2hNo4OYy352rxVR/Hptu/Uc+wDrjGj1xpg2trpmkh+WQ3yB2sLyXSupjdbmRTL7p59+Z0G
yCbZ6Glikf0xKsYuS39os1AnBQCgnQ6OwZgjt5PEU175JSLhdHeOm9t4Pk3nj5BWpvWJCY8pS7pW
FLXPAR5UCHHbdPeXMwdYQpEc3dIqrpVH2XX8smq974x3GU6VhqZ9jZ/Xt0oI4Ia2r+RndDI+SeKR
Ekk5hfnpq8YraFDvXOpMNIk5S9o1QA1DMlbPjpqZ8fFPuTPofMeIHFlg5Fo1wRI0tOiFUaGnMtAq
yjIWioPPzLh97Z4B5vsqefB3v1WB2kjhT3aLaL/4Jov754dgsuZMbvCZvARNScJ46kbl6s8YgzBW
2HQXy890OKt8dPTBbYicumXdJCGpBJCeG6B2o+NOhLemumAf/kHFBJK+wsNefef6R4hd4uznjw0y
BmJ9buvDnjPTAw2S0Yuem8ky0Wecr2SPAh6IS/ow2q7oFQWzztVnkLbetyUICkNdwxXlXJ8z0hJR
J0fUqqf40fIM79u0dhtBtZrS4+JfjEopI01AGx9fxFOFfNytwY2ssVONvFiyAWEC7RVjudJyI4N/
qhOuiZ7SuOsHUMlatumBAz8jgJ4D+qyoRr9IEEJ9lyh9fPgxg5uEqcSlDZvvmjzzkdCMwdMWBtES
SyVMVK0pa4IoC71wdSvh0yOUeQPs98CSfTcG3CUkamtn3+Qku/EMBTxLuKdKIooDpOCefqAhUOC9
QZvnv0oFfGeRICNv+XTOVTKM8n1FE7X+75eJUBZE7YuQepL3U6A3kiJ84vKaehHdbZwjN9m6VpNp
UIgBIxasYOBaN+qsr+mqc+XbMPguuBjqTChmDXHropgXOr0wnq7x914THlXnHw3xn8okqGyFP23m
45HWp34POxkH6BbhAoQGXK41F0GSW2FhmqDLBarZEJksyJRUDKcyUBSyjHk6Qls/vdDDxviI1ceX
KIITGdmCsfAP3/9+vxzPuLagCO8K/nex/5G2OHj7ucPmcdRYzAcCfUl6SF5D974VCrK364+j4K99
yjLz/+8CQHh70e9wEFwOSle6Y9GXU2qqV6gZP3//jVMPpKWFRCObEvRSlXI79k56d2C0tb2ixtHM
sA1yhFj8uvXjbBmKTe+XEfCn5lllgkT+9VQ2mSJK/YAtO34Mlxf4yQvJNDSU72CJ2okIQnbPBi+0
1ee7w5Skwp74o65Q9pX8DLKYXoZ5he/PwC3T80EIYU+G72TS56S07zjtfcPILMFwmjSCy4KZmiXK
R6y/IAkMH25ixRRxRLEHkxZlGa8oEJ2AGNORFESBPdHmuy56xICplWXkLjs7ZmaVIadE0UiFnfXl
aP47rTLma4nIqdvrtepQGfjIy3J8MtQvoxv1Yp3uUTk4uYpUp9oIwLfPCIu0kp+CLA8miWTXlvEa
yQ/HdfwrT5dtdwiu1P0BicDUKVDxV4oWShi13xxnsRW0nVNSSilzeWMjX1flfuVY7EVlQ/XsmNDZ
G7/D5WcI6Fm0MGIB/UglgsmC/2d0XwoNkgZv47tL7ZTABZPHt37/LFTIIrwAUnBE/pltoAt7RQER
LnC1WAvxerJgSATZuYT5j1JqqUhpSr/c9N6PnqJsEcbdI+l7V8JrkPznfO9b1Jy9tfFbg9eXVysr
W56Vv5ftxXFXViflR8p3EFECvSvaxBD2LekeBY1y9CvRFF4yALFRpaJgmVWxJpUjZCtZdWmcmAst
4VkcrxlYSSIq7XcxKAVYUxS8nohGg9aXYTf3J8KksMeP1cnmx2NC9g/7rUxIB6CIGReUb4esJCGI
8TtR39fTxloV3MzWk35JMBt5b9Ts6NQ/yDGeSeivgA7oe2C6OgIvxIIAt6+KP8AOZQJMfo/ns3Cn
qto9565JbGHFRsvVkrI29EEwUiInjSC6KVk/06CYA2yQHsGnoHWtVXnvL6nwvAjZ8cRegH8IX/7N
NPJ6KqSvYpXZVVbCKAfRtsv7VmaYqsxDjWmNV5bBx+dyGxWI0zlN7Fn5OAtWJ85Ha9pUdoKAeSR4
Nl1IpNLQEosLz5v3ekAkB81kSTJFQFo5ZSXKUJL99+E7axYOLl4xKmC9efKTHcw6h83SRulUSV7f
6yqsY9gIfkEYNbbdwQ0+A9o1D3EST95S/hIch9dLqdZlGQF4SjFZx8VG1w8GHd4G77pUdm+lJ0sg
Bp73occXbOE32brmPlTO3MM=
`protect end_protected
