`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 157312)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAGZlJFIW4SUFs8ceI5L5QFm9CgKXKD+OsS/le2CP/G2BYsAEZ592Xk5q
sAQzadVL5zNsBO4nOGFOXqfPEYXfoZ0d6OkAdco0Y2xW6WSceJQWBUlIPUyi0bpyAGYY3mpyk9wc
/XjXrKO/MOUvUlwc8biJ+AMJXf8rFcv6QrChztqLeZQ8AMuLdT4o1hWdk9w6W5WCFWZJ9FycWIXv
fNuT4EI2sfz6vXPe/HITZvw0tcnMT+YDAuhLG9sZEpsP16aohnuzjzo1et2QPunApD2RwQoVQ0cW
fdpU7kV75M6jAoC+oLYGhCHXNR62QLEVRicWOsERxwIXE4vKAZC0e5g2gaGra1geAsjhnxd6ecVB
PjxJNpVcagJ4L/1mDjtb+BikQkobuDNqumPO2Pa1aQgk44DKPz8D/fD+xQumQh69D/UVCFzrAt44
OkbC439EnCftY5SKWjq5I2YNz47S6agsm0mCZ0lx4C8i0Gg5X1PNPmD51HtqfsrDOS5BVEqjmAuY
PmbooQ8gS7Z+A9k/VJgZfOU/980ir5NoKobFWb9dIZmgDAR6G5nafMRh3h4e1kTYZjTLcfv/Y1sy
5WNzoGaii9JFwFCVDdDiL3CcfePrkBTcN2kBmvCacG0hEGEmZOi1BgcoBvB6EO6A0D96C32IVOEx
BBFPFYCsAuIgei/lvjHFO/ENaetUimn2klr9oNT/+hMSzflHj3DFxa3j5/Q8htrEimfCZBgOTMaZ
SoWTACcA992CJitqyiFq6lp2nyco6cPuD/7kqzd+ykZtBcXuqc5CEH5HHQgxQcdlueCyCoWCicEl
tfcYaCfuRHF+m2YmF4lq6h6rCpGptWd+yIdV9ksdxtG1DjP/qlqAMhfsCtrcWeFUBzAww9guz8Kb
OtEEzsPJAhsCKD/J9EbrpK+kB/q1aOQImROqqn61i4LbVmz9+cHoe2mfWlp2eQ4479K/R+vi4u+7
YP4nV64sxmYymeCVOf5mppDYqVKWRwBcPo1PHqk9bSyFoBXxFThsWwq9f6Vp6OGrem3QzsHCNhiA
INU3ApuES2/R6QzleEqBbVVF/+iZWRpcYM97VEXqTpCxScJAKizUCkUfXr/QmBP0sjIwK3b+66TH
7+LZGql4cgFNYn9UJXNefgeHgd/w1XmoVRBcKAb65o9L8e7VX0ZHHgNWUMXNxLmHd6l93d6Wbm2e
fBcZyM5m1CHZDqrKUn/LVEw7b9DJyg6Sl+2UqeGavCElYBmBkNJT59Qvoen34yU+BZpTZqYKczkv
KwLlJjqCzGcCOE0HeUNB3pU0sWwbd1sRHsaVrBevXWL2t+a1ESRUu0DFvMDPKO8A5JrGUKszlYGq
tomCEFftKi71eIIc6cbec6rISvzCl1LgDLt1CBrlg91bsNGfHoyWzqa0roiPmhfG8kauParY6eAM
TnrW57z0btrQPSpM9PlT2HspYRE3L10riDV7yH5AFf+5ZzMLgWxniNAYOV8TXLOTZOdq9AqyIW4y
VeCZACsHkWMFHY0hI+pwuBqEQnDx3405LOLdfEt0XndegZ6G1PJo9HOZPFBA0nwNtMEfGTX0AGuL
A4Gni7uqlbhHXIslfBVgmZXxi3q9ezmkRBjF0/1a2WvmGWsxesE8eLn8kXHfAgeYLQb8ZDXzW0r1
1OnkS4nSthNzKisnIL4GsQkfA+6tQFT+XUnLGdJq8Nmq71Hr3WsxqQabOTBXExhqoP6WxFtuszXq
42DkVRCQFIYA6yGWLIx9GOhDrCcKnDPk8NtDy92Gm+SjOHEmE1vFB2NXOd/lJAg4gG84P4wwrJZV
AwSJN6JPY3iomYA7+MC9/PWowOiAo+0C2y96+TTI6p5Nz1PYgYEBg4wuc6JabUFkcME8c9nnB3+R
jjRgksuUSeCIHfd1I0y/9yqT0e2Nh/VYO68WzOxdqpbpouGa3Jl+DTTfco2/R6JyLR77T3WWUrLQ
fc3HuPZIftEwt0V88jhXwZnwrcQshlRkLLQKDNc4E72HKtUmpvXz+IEL4oBgCOib4WL0L3eiFPSZ
VHB7rMye482Q1crUtj0Dt6kyxK9C5iCA+5RNDhOBe5VBACwLCpDfwQZdHmiAER7XFveep1TEn16S
qJZC5bz7CFApFEFDvga5NEEm7cKuJavzS6bGIUPVtkA/RfLEWjG5Ihi6sHq5uizbYavOV/YDwRjN
wUR8M0ydfKbwH2YKIjnFHKkkgjKNFWf62jrq10UXhURt2aUyXZMA9rPLuM4CP1nmQSwMcQGBna26
8YK5zodPUZC3Sxu1mmFqeFMZa4ppXD0f/uMledkApIyN0WXPuC4UNkZBS6vngbSUYU+JFif+8Z/0
uRBy7ef2zlEUBOzpwRcJqsloTNUSRtlCDmrQZ6d5dQnFl744kLEIQ6nKqP25qVLpn6YPuT/rYd1z
pMIK80NPWDeIaM+QcApxVsKqtSuSyo5RoVX5A3CMj7OrjiEWX9/B5GVCTfe/6+P4hwpxR9PhGLI7
yz0wCkLUbve1NsP210zNb2/qm1wB/xMyb9IrMljrbqTRrZ1nMjdKQtXKxAITHfnEyRzEojkFqQ2O
72BZDp5Yst1SafKKWIyrTwHNzJHaooki5Kn/nCLVzk5NDThuv+y6xArANZoBD4pqS6j5IZbcQj3q
F1HlAg2q5CQG+n9z1tmnj40yDHRLHJtzSKHZmefI/T0DXwAilpV2esg7QoYU2s4KQjiPbnlwnChN
zb2ZZ+663XbiaEROr3E3uVxilx8y+yDBQOuEuV/rTjXQsoMXStqVcynz8+24U0GwgOmy45/AK4Aw
JYDYPWGzEpi4aJ6Id2L8aiL61pUSAq7KY8aSjl+l/mteMVsuehZNSnGtaHpfI+XwrEdgd95VE1oV
p8NzPXHCbHTmEGqQgPEKy4BDcskb5O8pRtyQV6hounnQnFlZ68pDffFDk2e093NMM8QWp/k3Xdb8
S/44SpjCcGrHW1di0Tn+ldgVckpAqZmWSLOrurXqYNQr2bAWBn32C7LYiSbD/TnF/oFFY5x/u+db
iKS4YNvu1B2/n2qDp2IQKH1HvGEq7vLt+lGRT6ZxMUq+c4jZnFrlD0kOisSxlVyxZd9ulZFoqQXd
wzDzF4m1SjCycfd1x+MiiRWXpWiiM2UPTc3+fZB8/JCra8bFddKJkQjqWZ5K75D41qf4TJTKIAoo
01AW4cb8V5SLwUmuu0CFyjHJBIfOnrVxxd0eTmqK3zQXNIOw99M4cmAdi9qx27MKQFbwKxn4pgvt
ZkCipHnSXcmt46H9b9L4ahFGY2teFheiU0vcJdk10X1335R6ZTypr0kb59G2h1fbmJr/HXoGktT8
j+EcjAxs0ve8msCFH2IWo6qLlQJ0hxV1mePV7LCgXORdcESIcVTr+pRWK78zbmvFdw7OwbulifRH
QcPyk52f2O50SNqJzj1a499JIb/9GNXfiepP/Q/O4gAM93+/06c53SqdeRSN2ynQCvP2mTsDFXjq
r+GsMdg0WWp/Tnf5KIcK9GTvv7NbxEQ4yXTWEiVCCMKIqchllSbAb0Lpa3iL+RJpCmEGEUPaEJ7i
GVW2BQO+Bmx+QuCauVVZCXO4bo9ZWcBLiUjGLMszjFEeeTctvBVSYb208ZPR/NI7r7lSWUXYhbnq
VUY5MCgGgS4CxWkY1pImUsX3864Yk2p8Cuwl9J9II/Yff4iVedpyOIFsbMkqUYJGoMsUVdyDUCCk
hlWGUYWnQ2euhSpotFQbZOEGvkv+4kIEdfUyNgJd0x4+qRUHZQVLWWASUJfMV79XjCbuoVdYfPPH
F1VTCaTw20mWsjv3UZM9lgJoi9eFp/eUqO/poZoic4pKt0d0I0uJuqh7g8ODQUNfkhulIY7xylJ/
j2DAr06N8CSn4rQbaGITtGq7mzZpL6CBrZzaapu8CAbdvbWnmlIEgz4cREALk22OnK0+oQJCS/Z0
j+H+vly8cBRea3C7z4O9ZBjO2qypTndNE/LmEigw3xkDjMP5kLE5QOeZqyhhG1mGBCmlNP9nDuxA
EVkmSAadQ4izitKlordhy0BhrlUdUlO4yIRrXX47c6bz59MSZ8MbHMnDgZSBrG8HbSObZMbOMwEb
xzO/7fL6gQ+Ci/j2UwZUNjkwOe7MPSrRPPPhEgP9LRhO56jVY95UGuxjXhVkEfIgLpAJ2G2a4ud1
FvMHe6Bir88KWL7pWC2pdRNPPUOamFOGr4d7xwyZwutBGqdpuVdKyG+w0t019+w4XSISeQQ8CcVE
bq506red38rT81k9Z/kSH4TXvuPdPy37xGspvCMe9oDe/I/Ja3fSspBcdjgdpCKt147UGeNwYUDH
hOhBmnjJU1/i49Lu+gqMHVRXrjjdrDvOBfoSOb0OXN85GGfMtPtBgjMZchBcuOem69NX+lMyw5eY
YZv8Fs7iY7i2WMS4m6fcyglLN+sElXhJ2Xq9Bgsoc2qcCeyeQzbQ+QpMFeS+qU+el0ybiqIUf6fj
22DllbGpeh6E9iw+v0K3nC41pKFrNLUMd6ODv8LqHZSiacLj1rUkePej0FhYES9rn+NT+pRmMWt5
9WWgAVoEjBLj706dZp2vbBsspF7PggvLh9D9fQqIqZ1FwrJls06PE7VSQBMNBivTjihtvXa6cnQa
MHmBkIy9jzhW8TGxXCGPA6kA0+16qXtm0xJVk9C8GEfaGH+Th+ZwImEc/NoTMCGGJ+CaEw+PTi/f
CZKBXhVuGj5gQZw9GRA3f5l5ks5+BDCPl5NvjY0Gx+CAmCMsShXtZLRa9QspDT4TB1E1GtyIDYWL
g6RgQH3/NNbJklVpGjkKhWYMZiaQ518/X84zA/JwZnPyjdCEX0KUfNylBjzq53Yp+Pz5+skww6kI
PdVAAin93PEwCKmgL8MAwPhHqWjBI3HwMHsmNcCF9zBTLcgS2cwYkBSXcpBCiyHCCb2QiNg0Snyl
rwfKPZzMOGFj9KZXFgMxdbFaFR/O77kfwSMWB+WtVpukb1wgnIfBGuY7cY5HzYxFyV0RoW5jeB5V
5QKUc6mU/OTkBtXQ6Z8KZ3xLUhllP6PBKKY3KNaAGy1EV3W3gf3ckWP7DnNk4Kr9ZJC2A0Lj6EJG
R3YyDiOysemMfkSwSFePUT3K+vIu80+zXjaBMNVd1w3Vhljrwfd3oLHxhYX21ZnEzXym7cGGSKDN
6Oy/Hj7J65sWGXIIDWnMjNWiDIURaVDrkRUZMsVJVgb2BDjXCMbnlqbiKIwZWsyPiB4xobasxK5P
4ZJ1DaceDAJtydxa+6CgSp6mKEZhFAz0El/+VD3vsZleM2BBpQQIdA1Kp+c9MEBGOotkbGWPnfyB
ZnJGAHzXdzmjL8XkqYRoldQe1NyKix7xrZ1mQhvgdMOAWmU1SBImf03zbep6l78v2MiEXtRHoQiR
EjAxYR8suiFrwQQzBHIfAo1YaJyvYZwcZLsbeXZnxxyF2SW8l5JjQR89fEubgmgfzTl70XiLBqsd
aRvcsqIkSaZGNh0h9eV/IYCDqQ+l0viNNxb7M9GPaoTJi3j06ZYTLz5yppeAoTR17kWikIn+FUVA
gx9piw7eXzsNXzD8041gY9+fftKSfVeWKrmrfmHdXQ6Sd+nkIXl0iGDlzTEMVJQxXeQ3LMtpI1dI
Woo0psJztY798aDkmbMr2OTdxUXc60ovIum612XT0paEoc0IhBYETthyeSM6Tc1u503uzPRlY1p2
+WkB/2CFQOgDZRFiazfkA89HMJgJzgAswj1LO3zhogZgppnO5GC+uNCri/19sBhTXyLkzoz9jfmx
tHE7++5h22qzejW3MGNzPX9yntWot8vWkc+dy1dtnPjjAr3T4O3cv3MDK9VDAxeRykK0t6uETAo0
e3gMfpftIDn5stXUE2R9U6GLHemGR/z0owI9I8YjJriKdlZk9XgexLjQdSwXatRvzI6J9lEcl7SD
cW5cBk5OFf61BZAMwKeNDxPem4Tz1EpSefwL9bcOT+JYpDNAL3BWJODy6B6WSOJ8BBys/nbl/vjI
csUPSBzcFR0/DbM9KPzevQvW1fsAMtum8KyuGv8lOCEwN4I86VoeScRsjtXOXWenAPNaSNLYBxTk
yjujL5fSCOh15naXUCrwFG7WEDuE7BEvUVAvXO/4jV0rny13ymbryODcdLsYdsVyFJ8Sz5lnpKOX
n8d6OVby0Q+/2LwZrwD7zysxuK4BO4Cj+6BDeGb9lXLua3kBRHZFLYQYKNFczOCzB30DRxtWy6n5
k4eHcc6RWMpGz0hN05QiZybj33evwd0dkdPbIejwFveoVhTM9flkUs3oIAUhM0zZdvkqd7aod4nK
7qte/CZCIp5xjdo7p7UCw5rDrgNuc7hFHVrOssH6wZaNrBlvJfZWUvZopg/0cuqsXcfecXrF3AD6
lMqq+SE2Q9qhNtIfuUH12hdLgDP4hSqvbEG1gbZ2ssVeMhDtyzpdNpphpg/hoya1GWnBHTZK896D
MHAjItA2+V/AqmP1eKlcBmvqSLoGmEH9LCKulFN4tedf+vykCBA7Lq/1Xk5Jy8TMcjKHre0Dtqyg
AZvioYu9GeKtEpIJni1+auLvFxTNYhqGoJMyh4fNgO9pbb0xeR/mCD67YJKq9gVZy480sD6Dbfdi
MVdgxEo2L79RLuTfIFTYNSbVuQoIk0c1Jvo3PhFe775JlmiuFmVHepuVGXZLLEX652Fp4a5zuDMq
J3tt+Hni7etmoD5w3PNDlGRMWZONIsB0iyzDjE2qsAY6wxLyhXGB77h9/msmn2/IlR6IbSvOyq1q
CAN2aORgxBvZVvrfVEnNb4zzgaFSQNouyz/pmcB0WODrHKw6vPHb8mvC42/mt69Za6WcLhyw3+ot
w9CJ/orqmzwPhJO27NBaW6/QAoOeEuu1nv4paP1aVD2tN3iiVJTDjcpa4lkcymA0F4NZQzJ/ATCA
b1wsZ7gSLNE08aHkxbuE1rTqvRQmR4IJD1VwSPYcqGoKedubcxCwFx+WaIXvzhjfqWF8A4YqRqiW
vY8SCL8QHc7+1vnA5p/JCWa34vxdnL+42pL77XDKS4KT+LDBVTphM4rScKN+U2ToxwkVg8IDBp/8
s4mwl0cMdq2ji8cVeloTjgCxNE/7fUBYKZGorMSNf8ZKAVzvLXFykysW6DaS2mk4Id/5B6wlJxSj
zuKKa7mGy3C7QF8xY/H/jcYkTr2Iw9m7ENIjZuCO+ibsR83pnwKg2qnHd40jo6bLI7FISN2LPfy+
3giMURZc33jVerVYpqZL8lE3rYhJ3T7cYaHzdmLuYB+jSbq/lVHlYcpn13JDsnNZcy/qdbyaQ8OZ
398N1OX/NWC7nnD7CoIyhkDQL+gFa2tS/5u2tDI1H0cVSFFp1QP0jSHgwK0mbPhAU+OQ2nlHT+P9
RiaQlnRy6En1PZ+ew6Sn+5XBWXj77m3uk0q4EyLbDT7sojfwKZxRSULrivz8pQniC9imqo90x8FA
hv7JGXnn1gMrh/TbtLJaelAcDRjWZd98DwUp58ux6SZ8fZR+nVeys6WOX5vOpcrJS2G5BxzNNY8i
2qXxcJmCFNP0XjQW7/inBTbPD5nTwo2bohyQg0w3y+XQfL9EKClp2MPuVIfKPWTEcKWCft6XSTwq
Ruxw/XzjjZBTCZYg4kPrbKykscMKapiKY5DNoTudJcdjUqJ43VE7L3WI51eHTNKhz1C5iBLf0H0b
nka0JqsRKWEXWzTiLI6KFVVeQ6uNOYT1ISikShkvLWkLpKgz9FC7M0rPDhnGKAmX4JQtjxZg5RKb
aHCwaM5Lo08COeOBktx4xzBEj7JO00Mi9gO7UuFxOQL6SAp3Ch9kb7KiIF83SHBeGueWktXpOsYe
6OIU+VVItS9GP0YNu4BBoP0+lf6d6W+gMYLBRfZSL1Equh7hlvnhnPbqGCxWzX9aUZUblOWs+Y5C
Sra2ese1MMIGFBIolF5uLNW5JpDnhbfTK6yz6BKPkovAjEjxhNrS7UAS84GkHb6iCpDgEaJdHG+l
+n99g6g7iNZPkQRUG2RNuBYwqM73YavMEOndRBh6h+EGGLlMQxtUNPN1EX2NSBOx0Wv7cs2W9JGE
i37Sta2VPM/z19S3CRGs1n2NVJyOutIqMDXxMC2FqumoL6ISu0hFXqNXmmA6aleue7L+OfR7xCY6
8IIoMm3ieQoY4MrwmmVowXEtqYhxFDoNUtHDfL/ENSQCtSq3URWVdxOhmWMPl0j2So0Ucl6ASi5S
p1hxdV8NDuYAkk0WzUrRAfljjZw0baI4pYBpStfwLz5JaZ8TcZHv5m2TDuzE2OULAiiFUTIn5ZUY
yu2q2YNGylx4WWKw/3+adWutPnPNGjyml5yZLlr18qt5qBVjOoosNYhTKKZaEHgM8LOZmO0kMxIZ
saqCOQkpCqQ4RbeaIuUu69dqWvhNZ9oQC6sfXESyQBvvz/1sI1g2zrEXUqkEf8AoRw50Q+1VdxOz
sNnBC6ac5ypkct4xEgOrEuGAcAWH97bBFP2dzX2G9AbnWmt4IStOIbU+qf0YxyjHDgKDA6dBjSzw
MEMMXcFUoF10xXcPp4C95Lu9P1C1QiSIUHdj6dRKUyOlFFHxqkbXgX/21e0OeUGjEnceesWdwjxs
S0ApdC7httsRXUz5bDa4XjxxiQL1xRLhxCRRlnNaWuEbSTNsXZ6A0IS3YLpJ4EhmpXSKCbj+BndD
otBO4FtLOKZ8qfDEqJAwNYpaYW7Rq5Uu12Meb0tmgwjLEFeimjFtmsoy2qCresMtOK6fbOEgFFk1
tuJF7kM9jWzZi3XaXk+FgBYWIfLhIWX8KJhV84+yqS50CaFoP/wmEtsjwONjZHuHf71BmTbBuEkQ
GYxUgztZSdoAgnUGYDe9gA5SP09UjVImkJ+G/nTe6NO4NoAPX6DL9Xrw9WyQitOc+rkinrh1egfP
YiprClRCCDjbmUZuFZgmjs1LXDFqBVYRgWPH6hBMTsIcucsZO3jCSkwo2Di0D0LyB7CaUhY0Ji99
tN0EFYVY2EdSDQa4xZ4rB9xCpjCD+rc7lRk6eA59WOLNawTBjb8JuuKsuc6CjsxVYguQHGzjTYq1
pC0c0JAWysZcs4i4O8aAgbnmuA8QKF3/SyaxFbUJkqrf4P95CpTnqIpqTgGIgt4Pr0peCEzAi6n8
5ufLSu7vwntiYNlk1AGpgj++FNCfBEBZ9efGj/CdWtoay03vESnfV14P1sZ901sUpo0bcy//AfZV
pSOLKgqMixGTJfTFjwuuAKoNqTOqx1+P68SedaWWxYrmgeZtYmVsAV6lUZ34uBJTZW0A3++ekgm2
dFiDGxfToiuiiGC0PPC0tI2KsJ+hwKrPWKofFhXLLm1Dd9SELIXjog+llu26/9vPriNMc/7QUvWi
ke6RUPBGXjWAs+ldQXLso2AzWA95/3l0FnTPBOLuoPELwdCNKQwBMVL9NBIBjdy62NYo3q+d9tvB
1CjSQBl4k/b6CEZMYSBuqpPwu3lWtbwg2ojv32bJWAS5JeAT9eINMgN9dKwbPQhgI+YAxXs/pQf+
0DmGQhTYTGQ/ctOsZlKjzOfHT/thStPDvAFRooY/pQ66FMebjfm+q/EtWE1xEsZzrZBtEaiL/NMh
in5mPdwLX6loF+czlNwaHdAnP0+XdCQfL7rz5dZR6Q8c4H6YEDNUuGf5ZhAXSmN4JwyuqlH3z4bE
TMO0A1El4NaiuaS5QSV3KkRSPVHfTLGqPFUlpsOfykvzkYCuq/uh4TZ5dT8UZPIWuXnun/qyZynX
XKe1BFnyJvCA2KdGba/tsCkI2JrOdxfUVUeguLrQsu8eFT51xbtwgWGsLBAYVSC1j0FH9jSdmSQp
TQU7CnvY+GnGc/M19/sdaqvqECbIoPXHo+EhaNV7XadSZg4/+PcB3HE9rsurKl1kiymr7b0eq23I
hIhbk3jWiPA90WBipwttm95TrDzYLY4Xqc2h72iWU0caTyyZx+4s+cSUic6MO4vkWhPBTxtVAG56
e+WpzleQxxCXW+wZlQB9TiRnsSOA1oKvHKFiYOupJJ47HBa564Ab4xiciu2EWkQ0carbEiy7Nght
0oDxVcddCtSgn2tMOkbBX/kFR4YpaJzKgRW7F6cgC9Wy2dHlCKMulyG8oIsbpGZjrypWY5beQgo9
VE7wy7sa5/XlCsoPAWOgdssNmUTDL0VIp9wTgnEOtNZS3ITd6plShUxpL3Q+e/3FwVHS2dwFWphw
SdxXeeN1cJ9/CVhAijRPhmEUPUnB0ALJjnltjYo6zenlGIMJQ+PXEJOj7XjRaY9gTGBZ+J1ueBVr
XzaFUv0jxocwh0mkGfznwI3oovHYlIPEDOxMsxtbhQhdAH4Jch9kLuqXRv53xu5cNKVmbdKbwtkb
pcjbWFhMni3wNbu74Y0jIdEW9SUpvIJ/FbzJHXNA0cIKKudyjIfsq6lKQnlhap+t6HXxNFVwTDyZ
NpARCw1KmE58txZYnIFvt+FJxlvMPFOUCgkiyHHms7niKEf1Y6ErTG7urF/bN7XsbjcRvAnD4vMO
+kc5/8Ttv/i30c8S/rdkEvyrfuaW9NSnnK7W+OSHi955wH8JCMET7355dAWDQtdPR0aaXnLOQ5uT
DVL/rvDXMUFtKJst5pnNMseFzHD3ABvf0iKcXyExMaR7cYa+k7XWC8Bi4GUI7idch8BJXUe46psT
UdgibbMw849bhOmfJmo0H70oXaU72cb6uBFCcvbkIoDb9NWD/WQmJcAH2m+WBci/6C9vnhDyLjIu
JWuAEyJuPp4QxaD+ISa8iO1u0oeyRQNaYV4Mo4UdkuX5qxUht5Sd3jgndB+usaHMdD7hQ7geZ0Px
4FOJ6rL3w3W+KHZ1hIL3uMQzgfF+h3pB+r8zD2A0uBLLOKSHEQyWQaWwht4y2NTWYJo2zMcnjQxi
dFTK1W9iH/LaW5rLtMcvmnuJmvt9UKnEDSnZq61mjgMwcSZp/0S5ZuBsES5bffPETXxasdVuu6eW
702k4Mv4fVL8TOSUumf3ZQp2mZU9aP3Oz4os02vf4noB2T1qFsgMJOKoQX85OOyNWkMOHj5AQW8Y
hKm/jk9NFLxZV1Klz8se4AcNlI3XjUx/V5ijdBsr78YAEglhXn5HV2vFEtMlMOd76I3H62aTFvxd
GKB8L68pimhqOLTYaQFOrFHgAm1fpZTzDSJKKeb9kpP4/r9uyGVwFB0sz/5o8gUEO0ssAh2908w7
NKHpSUmUkOzcyPx69d9r9fevMKvPweQelMAAUgA7yp+dajmD2of1jvL5YzekOsViJXle1u/l3wuh
30rahSGs7Q5UZWiBlhkNYSOgGhIqaojyJFlGma1aEr95OAtuV22nqlGlmxIqjRytdEKI2HWDqrUD
KynZdj0jDmewTEZfM4h3uI1/6alwrTHZ3upmd2XVpM/FqiK6Q5MbPxCpR9nDu+rYKZD3nIPWDS9w
V52CcQA+1v9AnfOwMVYG7Uhao26bqfE9kQ49p3iTjEHS1sxjLP/3HHWA6EOLTOdcL57IxsZ1mdnQ
rQ9z+AguMAQ0p8Mp5wMQK3RV0MKrTQCFcCJBu7yo2q8EOn4UFaRHPuBtdivPFs7w7OlMfZBQG07L
71eHJ57Jmo7Pzoc6FhWgoOXxJKsuzWJ2qPYBj+BrrojDOb2Pj9iybS1u0Rz7eH5VIVaxy0wt67ho
j84KTXCKGLqhrrShUybTk83YQCVhyKr07fBCDtQcHNg8gWpdKkAEz3s4MhvmIA2sEw+n8Yp9FCcb
0hsOsp8VgSk/CwVKZFST2lYcdga5LCuJsln8UhfnXtLSIYWUmbxlJ9wiEQk1QLIoUi6EyGF5bCjY
gKz0LRH+PWLHK76Y21kQ/Q0PzlbDTAupOPW/QyLpK7leV7JszcdPcH3ppBhrmfozdLZjQYWaRSLe
Xt4fQYLfdh5Zfw1cH8LlcA51B6SU0GPC7uNA4cfIeQNjQqadpsd25Y3MN6P+u5aT8t7f4tGbgZi7
6LX8up5FhRSyVWd2Bxks7czcQWrlx6jLdhxm1kYCylWakM6QsSH/iTwUlxrclXFZixfdfyOkRTOy
BxWuqJ1DKB0uUVbqWyInnr8nrqFYweSKjJB2Nbt/fVTNM837dWZGtC5xjrXgil6mKkNANWUSWkOU
Ejl4vrMWIf7ZVosApA8PCnkvT1Bc9nCHR2RRageer6vuzXjNhO6LieU4ZMnylz//sNDb1KAWBJPT
Aoe9ilPcN3azhqob/+3Tn8LAaQ6luoI3z+ddlAH+J7f3Vj6kcSUmsqqJywfK8unRapUtO0hOeZvr
cYTkcBUYKjKmFXWgdZkOK9cKeEHj815LpCuzUJlQRW97LunKL8jZs0TS26rH1LnVJHmEWT1uobeq
fSTxIgIV/5A3JUBchmu5HGT78Io5ulWbLYXW/htWv1kJG2weXWTTbNW93veCS3w0ZUePrgV6MDCN
YP6G67uYfmhnhzqoHZNYfFj+IJ5RuRamJSSljvvcXysVe8Ykqogh+VJ4+8WsxV2Jy6X7IZPS0FN1
wSnHwxZIBtn4w8iJozwQtXfL6iSqAEajEedYwPZnlvT91Zwpq71scyx/qXc7CrdwD6JKPcm2GQJm
YmljRcz6t2/ppbeiMw6Xm7e47xk6gJIp82J26uwpyeA0whM7ErxfXnsfAhOWExcxHj2GRCS8RUd4
ov5r/9kLnUkvJQ9ISBrRhKQMp0yyXluvgvDzp/WIc8V6HFqXU9TRoD0jEKHbcmmgjp/nMhWK1sTH
zchzRn2WV/2KZos0/0ERZL9SnPwPo6uYXFTET1sxDVN1CUrZAIc26q6YiJJisJPssDkzY4DjVIGp
MKxvWW1q4z65jXcbcuy2hYsh5MuLkAGPc6s3GQqR675+JjQipqvRf995GJRSPGu+deR+U8xBhAea
JHEjkAvSRUA7OWT0Uswv+Mhm8lTKMRTHH4j9l0ndw+PketbDIF40RZvuxF7kCB5/k9iRj9OvzygS
uiA3rLk+J/gh+JCJlZ4Ct0Ls885EdALdNVSpwAGbdhjCf6umjGyzhsFZsXR+q1Gq+arb4KM79GRm
hoFn+qjUQW7w01tgssjriIOvy6fX+BBRZiBvTSsStRsnxXlWuMceGEGojd/NXheBp3sHUU1lJ6qr
NFEZGfflJQ/q57epHqSXukG/4I96DG2km1NHvoN5HPXZs7YkE9Fwxe928EdD3zhPG9yneocAwr/G
40dHI6agGsZagvzgg8JnPmbZnuAl650nacsx68ZPSsuSuxpujhado43sFFSYvCJ3yGQ+VDki3A2f
2weXfjnMTUeqj7g+elyO3JRGgnLHf62Wj1DbRL6le3ELK7Jcpch78+1O8vt9OQ85b36K/YnhvqJb
R5MVXNfyht3Vx6Ym0mj0calzlzewMyeddkJ97rEUsb9XHD9v3VqJgWzYi2mJqI+ctcZjYEI9hb0D
EocsbPfw1MOzQGD9lVZJhrzBWQVMQhzsb0ajAkuPU4s5fZOu7bbVBX8606q9OuiS2+CseWyfazZ4
kRhmMatruggE+OZWicRb49zv/Z0o5qoNP7AI/Na/gzruOdWKvwbh3ni+lspl6aO1BQ5MQUnu33vR
Q5+BE/4a892G9uKGhiCVTIEBBoMKMay1xl8dxtoJkixi20dNNmLyzh2zyxUeqbwFpo1aNbDTX98H
Br1h7708dq425RwkKip6wMI8glWRbrAybatDY97UyNTwExlRNX0lAOOBnXbFBlR36TYW0UQwGVH9
xYHInmcmWsN2lMkqqi7XFN5FDj4B4P/mKk5HekWU+kNMlOAXvyv6QTsBlvxR9UAuZ2zdCJGOQle3
diKUVJBUEqMZ7pjykdGf6nESexKvwS9hHteaRrU8q2CHQ9gRhQpLr5TDVb2iUGqcV5mdSE6IO8JP
vLlFU6WoT+acQqajtz95Tx/0kBexgRq02Y8xMrt0HcBnJM0QY6rQqUN51/ehJJQiE5dp6DqMnzN0
KbfCC+6FoTk/H8ZSCtdr1EPGOVdiFDn7aXfylnU2BUT8IwR2Q+jgs3coLbMLoJi8yqt4fpdM4YQw
lw3W7qxepi7/kNBY6UmUR5D7LwnDZMw7xNCWiOyLIEVbTqifrwjV0dAHCtJCGvsZrZyvyvP5heEj
J3Z9U5SCrW4m9UeuCdsK7mSpiEfNkL0Mz1u91WxlUA92ond++MBe8sGF8VWjEnhOpQ6IDIIHjymA
f3EE/mVF00Xlw6yo6Ubi4zEPgDTuL2FyfC4++nIzwzQ3ec+ZnCqohgVlr0DdS6soO9GzuCGJr0N5
NypOYr3KjF9nUsekBGKsNd52w9B56tCGXpqB31ewf07d2lTwDUVvROB9iqydM+IzoJHZtf+FWh/h
1wPdHqSYv5C97Y5kCA1yRtlMkt5Lbr4jTvGOlKQtGxKBn7HzX6vnOCiogDFhsqUjtrhWsNaQXOhp
LoUIOLKNAOWV9fHUdBsPthXaCtiRGzOFqNQzD2H0Pbv01U49C+ndHQfiRT0NRSdmiAayDOuvbmJt
PQD/lDObvD2LhBYs+GApxqdfj4sCgmsj7PNjjnHP8C8rJM0OCedrtXDzNtxFDEfYVYTaDQHIQc05
V8KxN9GcsiD6b2LVr36T6b5eXuavfDGa4ArjqHtUz16YhpnslM0tBgGOQ2p29rdwbnHC9omPc+iS
7Hty8Ym2OC0hA2uI2LA7DixKzQfqBaGuwROjBAXwPWJhXKvG7TMOLURUOh2sxFF8UnwSiL5JjUaF
kXvwVPiaEe7RZzfypV8JWva5YtwotHQHWMEXUjV4qNOYHc5eT1b7JFYClBVmDLgrzqsSpTxxeuIf
vql+3YHWUuKvlIGPbI2zEzdRy8NobU0x3QGQfhQU4xzitg4HFcPiOElqogRPjTY0VjRRPgozgggN
aiYqhRvTGJxmKy/TN4ZgRd9p70l19w50IhaPZx19JgSZNc3BoP1ghAhfz3RHbLSpeQOgOZ9LBUhy
KAI2G30f9EYMvju1H8GXXQM3whbeVeiONN67WzhP5uMPVR8xd5vY6Cxk27hgEpcd74OR/EteCDbF
v5HaMtCKslYq8fvxUzUyXXrBsmJDKbkMXR6R3MQHlx10bTI4OTjQe28r/YqxPZzGQYQnGpIzAxc1
2egv1B/LqCHKUcY4lV1S8chWbG13MPYdfoSOrt9f3mf9quCzBETrwgSEPqB3o2yuEB4nRCmjLuIl
awVHOdgpSImWp3eSk+c1k9Q7isBLxogqAKpi1FTXNwhbCmKqxenAJmAcd/sj+uHw5HVhPphujX9u
Hu6y1PqJ6f5cwYYUq3RxAQdFCzO6ej8VWv98sNqCMKnG7mcqkK1H9kUjrzaBBcW1g2jWhZgcY2EZ
SGC1Fy4+C+v4f8P4+N+UJQ2yBdelnKWRg6Pmq9ndoVyd0IW4V6ncU2X51VBKgY1Wdz0kUAhPrCg0
hPf+qIHhFRRwPA79FmhyUODW6O/Ve8IiODtICPn49SHADBl877x2GjpBmoi8/VNzxwxGxseY+o7s
sabo07/LJXbUfHUA+W4INw0NybLCPYzco66lWxTWKM+ca9y1u4a5quaMjPDuFdLBKXZbo31NQaVt
FDClPJezykJE7LiKjvKXYYD+9UbIvcoyHOJ+JCwQorXUBJMfiuUsP7PHowHpkf685H/GntyKsb9p
rF40TmXDI1vgod93p3PWCvZUhOO8+oM3rGnhl9QTr8mszEmEJyCbsy+Gkhqec0Lkrzf/pM8PHOYS
tMXXLU/rbNKlg5llcEOK56isf81KkkX3YtL4crITrS2wsrzhk3q1CXC/eNhnynk/JTYCw6b7Q9sK
PHe9P2WHFZm42lIc2bQ1rCTBpLYxD/a+iBYslB3OjuVUjhOxiZ7CgbcioXZPlUHwf5acqKqseUHg
9AY2j8vkLI+okedM2cI8yrt3z94nBP1Zd9WeSOLAMZ/7GnAs6lW2zLOaNfHfslDCK95yqGk2ZKWf
vKFi5YumP6aOhZo7udc1XFv4sdw82/bJlwiX0x65abQ0i7Rm2SjaF9q3j8/3BUqXcDPyyin515Bb
8m/VqrqW81XJfWN7wvpBJo//7oLbimuQWSy4k8jU+PpogTTUrcv2gQ/p/eNlVDGQAEmZT4qoqgpa
a7Rlnt9C3OzKDqz8UAxxbf9+DzwFRu8yLtunXI/rgZqEkGGHhzCOwOoeM1/QoSu1VLyBmFTWjqlH
ctnY7wkubsyLrJtCxsRdsfJfHTVLZ0K2JVfHpNzRNWOyL1eNRQCgJkwLMma3DqvoZyZBE30puzFT
Yfe+P+Lg15wAiYne6NZ4hQpWsPUlbV4M4jXWq76yS3oXdjGYxuJKeaO3lFbBEav55yoUb7Pu3bKF
we74yDlbhC9dIvo+sZ8u/Yp4P+MNkH5e8ZLkexswPbwm3JE8RBsPJjXUMy6q5rpw5yAZMt4Ub5BZ
dlRFnGhe0MT0rIvnijqvKM2dzlpsNSTMOPBp/UpQhh1BwBcAEdUDdnoh2/kSCWmGIVMPCY6hh0Pw
hnau2a/Ybpkgd3gfhjcX/MkSn8fFBpbnN6LeaPquO+Gr4Vvc6R0T6sydjXEQ5fMd/8s5wUUr9vo2
bsoNMZ/H9UBndHNJPanSE964uViaf64z23MpCZEqNzX0mX9B9I7pDW2PKgxna0lmdF08hHFVqUZU
+lIA9oX8p69C3teufNP7zByMHjRbAo1eMAp1bY0+VwEhQh4cZiNdpwyZpg1ukx9E9JlTa6AFzjPI
eYUGljmLxpaWSmNTnDdtsRAg8jweT12jrU9n1e0k3AlRl621DY9Kto2G9ZNttCfRbyjlWSQHk18W
n5BF9nUp/1EqBQ9Z+pH4HBMpINzp5w2T+gSTKZ2vbsyzIQzbuEUt0txfJ01f4EwJoWiqgd46Y9U4
NXEuzTTk6yj+91woo9FH018Y/VFi6Ic1RIkODRXCGQ8wGVDFAMVJR7NSNHf08dMNGPrA8RkoiQFe
1u6wguvt/8QhCC1FoHyFbgkiM13zKmPhhfLhcbeEUgqIlK327ZE2aNobrBcMVXrd/M7DcDXfuUra
qsbY4rjZdyB0VCZoloAm1JkV6KOqF7b84XnTt+Xtnyb81w7hjAXKvxf1QQ+mTfr39wF4mmsXSoVM
7UExyiK+nDlG+2i+fUs4rhMgLZ8TCJQvGSM56r+hQLLD1XMuLSpkZR3fKmWdblTlwdiVMpOCAiBf
YECif3S2khEUCkuhS+e4G1aUnz+wi7Q7fHJSDdmN5ygSm46oImTUqh3SdfgUPFFvhaxwsfXojfin
+7rEl3jsCY0IkRVtKSpKXqLVV/1hc/ukN122fs4pe6ATctSYcMzsDBGImx/3XnhlmjE5ZXmHivZO
ATLT6AU7a57KAZmzeemTn9vLHYTtEZTr/fSA93YaupxSEgOXuJ2VbLKFzc/SLDIPP0gVmmUomjMH
WQdq123FsND/8a7JtPFNXJMQZ/I8iFmQaZo7+1t+blFogBd7Zv780gpGGaQ2jPRCObgBM5rc9qH2
OPTKDWW8nUZ6qu8blltrhnfyg1DLIcsIrN1I2X4RygmHzrrS68CgW2lih7sIGg/M66vHl3MOwWfr
keb7DfLOvqX5EQOnk3j2db9Ssgdf3okm6R2BWMGgEbhUm8R8/2xxVZ1ntmI8u17KL6+32ZFCAMBj
ZaoJJTDDpd0KFGqxj8/UmxyzWONaDpv7xh4pcPa+K2wtm0I3azD+fs8ErEu4QJTqlmrIDxn7C0ef
difGJF5nGMqViLdj6QdqPv9/9Txc11T9wujk0UEwvh2f5FUW1Tybh6EE34xt4P7PPF4S1OiSMKB5
vc3B8HeptidsyN0keNIPN53cyVbkfV8tn8DXvFgAhNGMKtc7DIDVFtM52z58SL9WdxLe92ZNrXAl
UZsnwouMQfkTixXPBgo0CvOHuoyinVA4DeEtkFyKft4/TvXYN/nD6MFQ20EroUV3EKKdqTVTzez4
/4vveKX+j4vPKxzP/p9bdDl7kXO7hCxtl/TlXawweita9Wper3TONWCcWtYaGwTZIBHqjv/I8W2U
LCbFmb6/kZwcVrWkfLgztPPYg+mtcxtKdWmDlqU68LHJ0DaI6WCLSZfFn0LdnH55/TTfD7QSphv8
WB7rDSQmqIJFD5DHPtXbjwINpQChSIH423uRG1bgABkOPTvXm7HIll7DwwHw5p2pb6DR8cJ5SBis
s+tkN2D7LeGz2XjUsuX4zV0Ns7MxphsJDPiqgo/kLu6otl7o1Fcp7f1DbdYH6EMqq7yH7n5msPVs
+ceVSeR1Q2FWZxf2sH75auFv9omGDwVtQCPlwMXkF8vYYKDH+BkdZFlBwzVD5GpkHaKzn3fhcuMo
2h5UcJX+ib7IMZfOlcSCopr/T52uetiEdc3HGqvBGlvBVVQVDt8WrxBDRLP8fBXf3TcIP6u/REjC
FIKAcbrFW+mVaS6e6N88VlzDz6kLO4JRYW0QQV8Eugj2hdeaahkoz/ewDWB6H4rWITcvdmGcRLoq
+T+IFn4YxZBLxwZdnDAd6hjhf4sJ7fZ8SxJfB2WuzgFsA0lgXYut60UxaiCXdatpzq9HHHZQWIMd
52pd3uU62hlAi1CoJfXfB+8u99cXlOo0tG+1x5l4DqpER5YtE1u6xVrzv4RFWyT6fJ90JVyaZ73A
czfhWRHlydwYRMctHv7vQ0igLt1udRGAIbAi3UIfF+KrKtCKzqdPG097WfBybx3ddDFENnFkMcoG
BIjUdBKfwW2aqKkXtgw6IIN6zoU5L/DY03Amltv/4YjPKgY5sYIz6mM+ZrM766XChl/R7zPIcN1/
GjgV7LUfQwYEU4oOR0u5qnAN9b1C35H0dKxFM9vv1jyzlsDdo/H11cmkHBPyJC2cVEUEC9d7fjtQ
tp60UDQz6G67upAy1XBhnkr06orn1MKgsdJURO11fdKEjgsGA3LbDshBrEqxbI3Zl4eIninrJhsA
gnZb6S0L9xXpv3EPudA99/qeaBXv83DI1xBS3Si7ICHLqeIm68J2Cr4IsHy6avxIbzO0fAl8TyyI
ILW10r4nhSqsuh9K+JpZMNbE1dkpLTHviQrtYOpWziMPE0v/RFS5t1SEZgighiwZIx5JDffVnPvL
/E7EART77qGqPV6oF00u6sG5aS3EuX+KJo6MjnMAHKAhEigLF0h9xRLTumddWzVTCnlrPwa7QVRK
s2oCNxYn4ubGMDKAh2wgEGBqWNJ2GEeTY0xa9zjky7sO4Czv1HZqK3sr0r3M55oJIpgFsGdmAneH
mD2H975YMBcU2k5ezrFSBFJnv8G9NkmDS/UYCRcZU5eIcXLiQVRTf4+HDHZOCp86W+UCewjgAkfM
UgJjte8jAaqVZuJ004F5oPSmQfzGILUGKuoiQ5EKWziVDebed4HhsHBxGbVvW7vB3cscJEEC9xDm
AZJeDcEqQEaUpkFZbc93e5hbSvIf+7ZTiPu7+Uwhsvn8XfbQvBG9nRzNcVrFUVEzzh6dncNUANIK
hzVbB4iTWzu+FqWD9odZw+mM6T87/YZRJ5jxFP6cIo8MLNF0psYSqpnwC5ot5aQQ7fcoPQJxDggs
VpyJOaor/5tBhx6gDqPKYLG4gxUHOapyrgCm7/Sb49tkq9cGpnicYwMEXjDvT9a7qZ7DoYLvTAMV
DMQfbPcEnjxr4ZMW6aditPqszzsxgo0xZtHODmrktlUBPSR8iA+DaksW7b1zTWgboHHaVny1MLFU
bcjVYwgDJyvBlqrVFUR8ZNoyAvjaDfI+dxk2P5/3OAqIgTT0H9GWQYDCTu+TTanwMzujKR8Xyjv9
P93VZjEH4415Eat4sIOmQIp3Vhmc4jBz8GnjglSdsZXsMN7cPeD1R2/LuNDGOeJmbf6+FQeKE0rP
Z+g/MmREVdRG3y4f/1075peeKgvM5gGuuCewFdIu4krf8dC6NZpX4ax9GI/i235n75o57vCGagh2
z8pTv4N8zSGPhNOnv/9w3Vg2lZKViWOv+J4g/avOp7BQRySPnNgx9in3JiG5+DBr8QewPmqYmCdn
CRlkucEO5iG1QZ5b8NtguuH7wQIaQXmm2yB7n3/grWXyXaZ4Vk17s5D3qr9r9KrBfNf4+wR2AILk
cWHQZse0YWe+YFY1ENSUUBR7HppLhIps4ARoeSn9XIH5iXk6duftpgv05tTiTfuB67nEuxgM4+un
zq9CSWEtHZ7i6RWIT9crEXXD8TlA6uqQYhoxKo/qJwVOv9VC2plVwj+vFhKnqvyMD05cPtNJTUp4
P28k3qlUhDf9c9Ox+kS2ZCXFjPKZ1NHwtwWbgerG8Mp0CtbBe7XnBAqB/PnAijc/OmGZL9jeZXmb
MDvHqnwtLmT70O5jmmuSlMChvLicg1YreNSpR6C5DxnKlEIaeqg7izCWKtdTylBwkdvoniNzifdI
BKexmhYZ/ZQUBO7PL3JZ3kA3t2CUPen1ssk3+eUGzXYXJeEFgN3qeO/thm5MjOKFXqMV++HNf9vO
3EJHOUBQFfZ0E7BieaxDDbBw8aJkm8RlvSRMnrTK/oDxX6JGU0HZGvSyIvh+klAWk10CYuWzR1EI
wFTpYFfR4WhgpR421P/zaqHTylNMAbby9vvpqdOgCX3/lVQsSgcmZCJt/ZXjQk4D3QMLrcObXoYt
StWR4PNzxDWSVe2IzM6Yn2RGar52OxlwORP6ojmdV7lp2i8RE8BzgaVU64FEXznEiCJWmqhNwtjj
JCu2vvjEYCt+nE6IsPLp/A5/RugmWKpQrqDTrkYwzL+UZ2abAbsbkHCRSbTQCOQZ8nHN2vWnB9Kl
RJJjlM4M7y/wTkiI6BmJYm+9Ml/JKJ/jgTV1BbdoyRCMxrGylDcERzeUXJhAw3SEMbxKno5dUrTh
JxRqkDgOf1n5cPplJ8bPkA44Y/EkZxjMk0ZS+XFULHrvCGv/EaGbf/AY/PFzKcylmvgy2y68iSSZ
B3u78+F4dhS37vUGuLO5++6mX99+kffuPG7GQXmU8AMaOINla2JI6ILtr/NRwBN6uY6gJkPU8uPj
scXpTM82opdqOCc4Gk83LJXc4UaRD5AMsI2qIM3Qmsl7uYqoAE3nkZckqaKxMZqiU7c+kufQApDH
atASLb23xRmWdyOVWp/BVUybibVrBCL4jUlK3lccREIGev0DbVZQpUhf5Jofu6kwNBz8696o7O71
n/LznLGt+Xnzb72gys7Z5n1KjSR+S2djoeowTBCS53T6anaXMzuEujh0Cdo+38hBQyNpiuhRLFk8
hpC4B0HB0iBINPq5I63hV36lRXR2anc91CedKv3WRq+v3Ii9r3yhBaBUasa1IGUJkqooi/yNFga6
+Xe8mJZsdWPWE+eacIA9T5IXODX4xlZCzCBJze9f/kBJe0Gs3GibxEq4XLnOUqhZjCDZkxtZ6rSA
VcJFsHC38Mf+rNSMxlCtGm30IeIL2aKTZmf+xcfa/Go9oeMOeUbcIUVBYZeJiE1WaajW5o8OpeU7
NKhkdJGQR2MUjn040PeMRzheKH+5UsvXgYs9rKyy6EW2XhHYHtbZbol+xj12dcq0FPQMlXbfBmjZ
K1rXWkG6d/pLqMDl4X8HPnrggse5ojhf4s3bVPs7z668B6d0iTp5YM7ai7f37U7+3eXqE/1koB1x
Pe4V6MmbBDhndWXWt6BMlOuZOa5ZXR8fsX7N1MsRXh97SubQS3EQZJszxb4S7MIz14vuWR9gwmiY
EHkvylqMt6RSZgYAyiSmnbny1P4UH8LMLy2azq+OKUy6wedgF0UPv78bKybRMdDlFyWD0uGewI3d
K9kEavEB3uUiIMypw5E6nF7Xn3yuL5vBx9yt1OKJkBZHpK5oMVk6U9uUgtob5PQojO5wpAOXLq8v
dD48crpdj/ML9uCk70XBLyBNNEW2a7vgJNPyuoa0YIIpN4CNjO8nKwMAeI9wag4BAxxGsww6LUG7
281bnbe29EnJMkQcaYcbyFlU7b7LqWTzR5rurATM4sXy2fDH4EINEveP8Ms567x/7IX+RPYdVnlO
07cseJVOWBvS5FY0gqyocTmhRvuiT3FHbd1wCg38zMfoghB2fzNHb0vUJqLqYVASG58MUWD88JEA
RGBEKFCyz/YCabRN69M9/LskkO9t8yiinoRS1FYpqIu15XDHM2MDS6UZ5OHwF8FB/fGtjomz5wTb
9i4ZCPk0g3yjJ6mBLN04Y15AAqCQDvJjcTmj0sFnZ3UC0o8Z5so86iPP6JyQ2gttaATwyzcO61kk
HFqK1RFqs4rCLxE6ZMWTvZMs5mULbPuwUIVk0bJptA7zGWXYRe0Uv/MBrUuBGwibbkXFq6XHOq+i
rlb4sClUDTRSqACW256MfcZsED+DpGDD6zg/i2hMZGQuKjq3H1GUq4Dn6OnNSvIBPAFUxiCZGxZI
OAnMvgLzmdYk8HLX/a5bB5+S5XELv5ciyhjaDeeXiUtqiZ1m5rZktAHlfIn+4p/QI+7scKS4Cqya
s7XyD1V9cpBC6G7jtwWqWjvbMTTxMsQlLQhcYxTyTteWp3xuu79U5GM/xRdlYDMp6v+he9pnuSpV
ZOoIy9W6jycwSamWPxKkSfVhdocKX4koaq+mfOm/HfNx9Zxq48IYv6ZUQHjAIEPwdoGYY3eUqRxl
P2KJcX2OMUKmgsowQtCSwklGK5hbpGOd58nrqvxvbi78sbZobrmJ7sv9dziiZJDtXIFz6cw8EVvO
XhYeiqAmXrJdQFd6udXF9aZN4fmdlqxjHcppREcqX0nV0hitHyyHqbLQLPx7p7UqgypORDEHCnfd
21wEBsbZpSUiuxY79ME2ehEVDBu5OriqDOpQbb03o+2skAJwQa8hxRmDIaQhmURVaWlcgl7zttoW
y6pwJUTEu18JF4Ge9Qvgb1YpiSogA03rLRR1ORVSU+Yt+bHETVVc94eKgJT5MKEpYo2N4bU2bG5w
U3WVw6b5rakM296IZMNtcCKw/uzi19auyRvBHFxMm79T6jTcvVW5F+gKL9xvr9bBIXlqRjg/20or
7z+CfUCWOzoppN0skj15V1Hq/YBXXi5065Ebjl1y+BzP2nNCeSSlnV9f6GJbPyufM1ZxNUE/CEod
LkVUcayhADy7LHIXkITtq5OVpOVmHt4QNkzEWQxIj4aCYYoyzg/qvezx5WACIBWH+MrLn0xh4FAr
FFrcyIkflCbRWA57aKZTbDvwIfTLtD03txsb+RsV4NT5EXMnI1M7mLJ93/XYz4c/zXQ7QmZBJZeE
K4KA0Am/keLaIAP1PEF5IUtRKKCmq/alBQ3XRqS615OElA+3t7f8gCS6IvdVRw1k6EL5OmCUoKsX
dVEozucAs3lHc+fogZR7k6i+/UbGuxYwFimV0KsyJdsCmOiU4G83UXWNx0DNOe6HuQFJGdZ52LHt
811VP5rZE2mZtn4bZ9eHrwC30+eoDMHG5G1WVei7c9b4/yG5dTFxzjYRx1BFxSHuqnJ0X6kLTiq4
ckqhYxpAQN77c8zMRTCa8lcOW67p0ZVltx9qEj/jmHWYzwfW41HytvShTpMRspVvSHgvQZqa0c4z
4BSrl2ooH79jc01BcCdoPAAaOVM0e+b7ue1BvH7THR81JUEIdXWVxO7EH+uR43OMVHgWvtlVkqq2
IIKIFeFp9muvBbxPyMOQgwUHvt9S57RsLGT92ioDzqEWpwULB4hXzB5lwSBZceM8aQ9TKs53BE0q
b/Z/7usS+pvBeUsWoxFlcJ+awEIv9YvNMRt7dzguc+9wMHtXYDITyelf2QvQrWxoNvEGoEjkDsb/
Z/JjdyYj58whiI7DlqanSImLLspHj0vcCr3xJWxiQIQHXYvy70hWHmI3TqXskdKva1BlTyl674js
Ib/vzJScC+I9CGs5BSpfDyxf0Ykus0diHlG4rG+Dkjdz8vcQtFN82huTA0E6RxwDIq0NKABG6Vxu
Y1Mlv86fSt+oF3GR6Uiqgn5fnQJGRaQFBdef8Vx1eMoOA9dJAKiuHpoU6lOkiH0F848dPtyQUSF5
QmwmGk2yT8TEfTlGvAtIDVr9PyqhaXU9YNb9FTkVkITTv1zDzWJ+GDCiikAHg9E81HzI71H7HJtq
Nvq0/0OFKsgfCRsN3pNH5wjb9wZtGFkUGn2q7VNSF73GAnPx2HMQt85ApAXct5k4+rp6pFZCKV+r
tPemvKpuZPaDKuSK3WW1G+LF2AEVMHETRBxpgyGiLy0iZsk2/GIbf7SVZ0devKjhk6DzhC6W6dAM
As9XdqhOGqOtmlhPVf4TYQI2dZ3SGFqiep6VK4pnYVNaWKd7Y9iksv194pB0uHLrp0nan3LZ0jVc
77n2iHce5ZPH3X81EjM5WwA5jBYnel797MhLzh96F3QYvwT/n7m1dj2xPmATx0kruYfmG2HSt92E
dqG9Y9wXIKhsshDTGjXExhpXdsMOZuD+XZ8uaNQjVVHFNmpn/4/JLgq4ac1Sj6iSTEzs3LNIelJX
MLKyQflXkbfz5kW/u6w7YZuQulSz9+6q49YBUj76mhZx2wcAkKNj9frhKjtP/DxOFIFIQDubZoq8
SQ5dAZXkmofOkp70mVIssVvulTlXF2Zlp9hxR4MB/8JC/SO8jQO35RdTyyZmWcl+5JR6ViyVVy9N
8SiniFcUiVVSOfHoEpMkVMMixYc+a0fF6dL4vXsO4XQN/TRKhGNmXsIdVeoINHRZM/deHCzNL3s6
O07UHxO4hcyEUNTaEfr0dtPuOTO2qeLj9+cTgr/YUlRJRXC5VxgRNp5tWgcnUv4oOMoS6kdaRFF4
sEPiNXm55esc3R6CfbJvFlftUSLWcc+kj+xr6TD7vs4FgAC+5AZdZXm3T4q1SNmTsBe83SdWLaDW
eQS24OtoZU52vtOpl1aceIXkJt316dxpW/mNiZm2V/WG+L1wDI00NMOBb/eTUxCz/SINOIEV77uj
w2wYfaBjwXHdvF6GEtiWQ9BpnoYeBTFUkQsT0QtMLICC7xzImKILaIQo4FMTB4mEIZ7GxiUfjTxe
/ySgRwggdUFNDtpQzmeAU/PUwFtWWCiA0Xo6MA3lCB0bjKVE7zw/cPLC3yhu6VJvVvzJeRz3assJ
HKfD2TIZOwP3DBlHz9Q+g/93CUmUqD1Wu2mfjR4MsqMritvrv+dRYjp4z1cZRJcM2Frl/SUCH9vH
VfKYv0dWaEbLxIxhW7+KyG4R/BfzY/FUw+osc9bKB/gGyizB+Rq1m09N2mTnvEHWDa1BbssVkby8
v3iaigSoT+t1NCcck9me3FxvR+FzPx1c4l65M7cZNh4R2CZ5rvaVh5rQUwL7UaUaNltuQT0UibmG
y/HOPYTH2r38dx0fYQeHPXgHH/VSUAdGaT3mJScwKTjlM/Qz63ZubHXLnlRyX2boKJ1NDGePcUrx
JpPkJLTx/B1wxAsOrteNFw+E0kna2kRJbVK5MyC5hOJD3U90s8a2DKxCLnf9UszSxRsU2Xp+birq
kySqWq2WJxrYu1z4qOd3BT34fBek3H0JldMq/1y392MLlaijxBUZbZ54r853DemVixQ4owoD+RcM
BgWE1vwxTUKoLcr6ySk0Lv08hqz36jMnT3jreQ/Celj0wU/bpK0uCm1GsxNI9rnCGPkJTch5Ci1d
PnHUW0zIdr8IhpHxM82RK6oz3Tnd9jC1vQdcdUqt/EJAOJvLKPsHv5zhjjCI/mkkTdRwnwfjUpSu
1oNOMDvIq/WAYupWFT7DUsC2Y298uKyYBZgYW4Faw8SZZmyGjahDkDMU2CzQtF4xOH86Z4rTRRLP
Jd9MxdBry87CsP/npqZ3b2YBZBsv4wCg+Ys4/5h89QtpPWPDN6XOwhm95BOFWMsMN/Ub/kyhdh71
GxUbadLqmTHoen6FQcWPLmk9qNxVLAqQXpWQcP/EATyDvxIcFf2verJiFqqFSZMN6YCbgSywPYhH
JIkEzGtrLBMID8bnrabEEED7Pk6IlrLk9O1vcYHhy1A+wx2wyjBwl8erzil9+SaKSUGZdM3pLQS1
148rfmcXs1RmuTqGZnb3e3aW9J3ddRyc2086bqik7QuL1q31RcaIP8taqeYyBiOxXX3PoGZlODMm
UfNu2os+m3upRIgsSYXeQEuflCngBfWDjZ1BZfDS2nyEtRhtUBOA+UJvIzQIRoqNiCh0jaJBVzH0
ffkzZpfFfASMMnNBd3ZuR1c+3Oxq5/cyMj/447rm/0+W64vi5+ll9Fs1Wt6qZKdx/KqMikKWKkjS
nBPaIbUWMU2hO8m/oOOIKYZa7misfi0cRoNN+awRDne53eg3LiHtISWchD8/HCwOGHLBG/2QLz3T
e6XU6TloIECfzmtKjadjzvM/rDGVSesqQCbmo10NGCL2meLCay0lvDm6GT1ymizM91VkPiDryYAc
Az1HHKCg2ydVFPWcCZYmvsjMvbopccPJPVowfsA/UXdw/SDEzKKeUyHTOiPAT9FwOa7S6swvmzsa
xDOOkLFo6iaIsfPM4Y8+WBvgcT1md0rognP6n9bYtGz44IGXLDgIYkGM3kaY2DzatWl0fqTODa4m
3WLc0dloOraX/xaX3oaZFshYFDp1WD0V2xDMkaPSiGM0iabGzF4pQ1FjQ7Tc4KgO+UDnHuhrEnSl
eAEGBgpUp3LFsVezjJKxbGDaLNRFX99mJxrp4piDGiI2DL+XNfYcof5zpo+l9M/jIto/tDWgljaG
p1dvvXO1AGpByy4jF01HjsJC17FujXGwzKS/nf6YzwVg80qcE6oRyy11P4eFI1OVCTMQMRO9Sfku
vN+lO0zWJmimaJIwtjyPDgpHsGE3BX97FpHvym/YDBc85ff+gtL1CI2ebuR9xWb9Uvy6Vh4EnP8I
xb7puDiZLU51WSNLnHi8UEzfNGD0thcWD5AqaMghAgaZwctXeNnxD4I/upQjGyz0xFb/f0UDWwE3
MY0IYWW1mASCsMr3ozGTe5wHJtqD9o9Ttlna3pHLuw2QYJciQcNWjJ/n4HgztEGuNQAwKLjpOWp4
VmxTQWSDAMPgMbnztq9uHi5Z07WQSSwTvShPB8uJX3SvoVkDdCNsbFhBxIvRDkc6+1CsoE8ONo9w
iYeEvlcOTV8Cr5DZRAhSIRjBFdMUxyoSKP4xe29t7kkZOEVMMBt4rqhGSTiYrKtMR9LASxisrEg+
nk/xYI2mLLxGHcGp2YtLvLj9wbMc9TLDFt9/P8jPBFzyBNZC5RVy7deoPvgZz5uaInwPpiuBilTa
4sgtc9Bht/r9FQ+l0ESYt3jf8nOJY5E2vK7cF6otvriacIDnWP3gZh2l0/5Ki6GiUC2GwEJPes41
67dGiJvzv6iAbrCV03pot6uXDdrLJqkcFf2os0glBlA6E6c8ZhoDrj/2CCQ+vE59SjAHUDYBDDmr
5wzluoUOG1yazVX3h7mjTi4Ciia02Vt8SQ8h14gi3N00BlNQhhkwHiLPfIxUmpymPs9K7bCxUYjR
6l4E3zEBXu473XH0kBNwlJPKk8rqEb5q2PyYjJN6qlN6y+2l66R/cj+dFMFNSySgV5ns2VyTWsLL
8Lqrqi6/X43xHTrtUsoDFxTXf7qGb0naMBcLe6KeEWFcYehnq8Cm+e+xrspmpniTt6U4tV6Q0kaq
Z+IdgyHII4iZ/czvZnvNqcI1PPhx1gtH6vmggJw/MWw5FdwjM8f/x47RSoS8dfKdxXjOO33n8Laz
Oe562oXemilJzB7efRKuIVbF14ian30sIz/leZk5wYtnpCt6c4IunN1gKlQiqrbTy3m4nS/l6L6q
dmTk2dq4MSD1hd4KEoSUJkYwulL97+8JsuZGpsyqjapR1eu21KUBLI0YG3FLJpjNd4qoKwViBtNj
Lz7vHQbz+VY8puJ+LExCWfq2DRNVaatIrTllUuDHbcOXx6rBeq7kLNEV+TlPc0a3GFPeF38orjB9
7EJoexHL8g0CMYrYBhKkMh84GQmRKEiKJf+ldow4NCVGjjjlaXXQaxRM6dY0Bvb5RDy180T6qm6T
4ZpWuPuGyZMqTetv6mWDJYtqa7mNHnijCJOpV8a1I9mp8DpJ2So8kzlHMBgorIM7K4UAJashbenU
Pa09wNhF4tOwFrbJ1iYe9/3hcp/z/oou5Bb4zYDNhA+uQetHjqxXRDVJo71S5s2Ykbau/crPgvHE
vICz0pXlU4hQUqaW2HxYiwvZciNStZKEk5a/Lkf7tMD7tUGURr7c64Dn26TtOba0buQg7Vqma3FB
tUzg+QAfAnLdBS6yvxE5rH8RPEIE6hhaZZn+v9v1EPnqWrjVT2Qm8JsJ7IPFrsCF9zMY6gRh1DqY
0KVIgBt8E1QdIm46OjkIogvlry9AUFKQT/1ZqFPpwrBCss0rHMZCpSyP47UCNsBzPKDEqKqXj/e6
BB7RBsJ5PMOqUOuZ8GlJFTeNZTptaUkfpMXSJX3dNAfMwCwjELYMNZxj5mFEASB2C7X5G2KiSRrH
SCZVAg0JIVEe5Fg0w3nF6BkY962bYCWfgcYv/TsCz0zE0wK1oCpIXRS599Og0dVrK5n3B3FNbTQK
PrT921qlW0JP3onDU5mLyyP36UsKb4eWXsqvQbVfgBFgrrjiPU4Gzmd9TVrzsZvY6ZMq5d2Igtkm
mUntmpGUiljneZjbyEyvmYL5PzijCHex4+XGHAkumoC6v7RZ67u2u3gJhm/lftbODP/vPJ20G/U7
AJViJLpwsHxjqa+eJ68yEOR7IBx2JcshhB79GCx9Fq2S8hGur1CW7rzBVjJGw39KMsRTATQSq73w
DqQ820/+HQkXUWZaDlTnghUPMqRbW6FSKOAnNDZw3pikuiYephddkT2OChCVEwCmirjVuC/LeUin
UJTARbwdZRlvz3IG0fE/i7iVAQ1F4muKhrBh+0rDtVFAwYZkzlUgj0hnIM7CzKl2ESgxJKTxW60e
WkEAwJNUvt79tG7Slku8C+fAI5/qHnTlIkyuYKek4pj6jD7xadpvxQdv8zjywdTRLOgHFT2bcQ2a
NUsbfD7MgxRfRa3bEM1xmVTxzTASb3kSlve/bmzt0Zcb8RWbzKLjTc3CSs2eOj33zfoN4TV/C0so
ttKiX3bKZM75I9XTsh0RE3Tf6GmkDuoSrlumEmWcBbvQ8lBIJGPnIEIwZbSIFEud7uONzbVmtOqA
9GUNvzE9Llrkglyqv+IO/D8cGanMRQSL8QLzAwTtSF6n76OsnZ1kQ7ca/KtTNtofm+Chv3yzg0Pl
cHCwJeIeChj3rA078oXNRhun8o7LBfRuh38IUf1mIdwaVmTMaNr7amWWNdnP5u3SNV9uQdt2VGFh
J+9v3E78rlFf/Ks3l/FfYf8eEjptNZH65yUeuI6vfDLY64ogWTjZ4KH5GAIqMxvNq0/8GaZAUEbo
5REtFsZ+owsWkRzARwDUJWi+pIO6njJMvbf7JivqTLiQ/YaekRzpha638CQznLUDCLhHeyJ+eM/B
aM8fnzVGjTxzV7xx4V9vrJ87jpqxy0dKUOZqIgKgETGArVK93LvUNEn70XDMVsBF/awhMXx84Ge3
s7AF09VNjxqV/kZ/tLU2o12TeLT2QQwzuhyWc8YfSx/HpGROn2j0r/zRO386BA7Vv4mFDN0Me6uT
GCHzkOEAOrOkft0tTmAKKBv4dj0rZYc1T5N1OBsqzcHTrSuwuAIVx0cxSevjvduvq2+jZA3U5rse
quTmI9QMc8B1UR8+LewK/hly/HKpX66ZAFtI0o+OLKVSSOF+7CgqgWJMBcmvT4be6CzXH3qG2J69
neMMHKli4IS6eN0YzUQHBNSyhNox9uUn6+wTVmLgBJgpR3WGw5TrFLw9uqFfA331nUSTCkJ6AJR8
9tsGPPk6WwNVYhFzxxSVOn9gd4o1N2RAawwXd89Y4ZpfJVc2e8SnMGnnt6O+WiB9Zpn5Kg615yr/
pArGJoTFe7Et3taZ31eDt0Cz5XCInYC2J57rAG01MU9BVYLkEW9rmx4YMbqHSf8acWPnzNEN3Usg
zFllT+f4pQTNv/9Mik9KnkETPIkEOyMYZ71Llue9BkgS7IoyisStIBM7+tffCjP1ySl1qcTH4D5g
R0pORFhGSo2QfvHnuez/8K/Sg+LGmTb0pj1M9jmVNQaT0H6DX8TFGcQFfASD8cJqbDuySQckvBU+
Yk7lsI4HNvMD29PfMxZdBa8J86iq4NbLDSmOmy71XxmpLWuF9X8Ir6EWmmJkAzT8J40uuVoGSgcQ
CZadaj7BWUlpO7ewj2o9o+SurbiJHZiysLveGF/tYkHV2CDnxF/PNaL5Yn/TjwYPlC55VJsMjg+s
P+rN8kXc8BRLttVF1E46HCXEJNW7wxqSIn/G6xlTMYbsPCSlpnblCWLUCxe7xrWhan2DRHOFxXwC
OFZ81FshS2pNsj2yFbD5WVkaMc7aQ9sGOuCYChNhuMDr6LExegvUIVTqOb8pCzE45GgcNHSNaRtA
VOR/369zwhwK+acFkx0Nm9VAjgNwh/AXOdq5PICyytc2ghfD0o+Hwo9YL1FodfXCL9wlrxD/85Pu
8BD5BnhwN0lXBtzglR/Xe3vfqvFr21exj54dpwD2bI/wTXkBULem0kp+1eY435eWkBCddvMw+5CV
gueQF58Z/x61QBVSJAwrif/XYajwGIMu26B9WOpTot1WYSCjy2ecg1pIbdZZ6OQhO/7QQES1FSzx
S0NdyZIR9bGAIQkb1sFUGksDyPSgqNmxcZ/xYHmnDURgWe/MINExoc2+3RIbKSqbfpFV0WB4/TQG
DTHFIW6F/yjXsY4qhyX/fN8tmxw1xGnVc9/88P1YGcGb2uuht+GYDmWudNTCVnBpbIWS5cisGX+H
c1tbN2C1XQltMoKo8lxPsaOwIkmwwnbklWLsSkyKYlIdVgltCdpUILCXoBvtiUFhRHXu8bXlC91C
HTNszLLde/qPpohAWZDNddxhwyPuzGPBGNIUq+g4mBitesyu7XCa8j0lEgXqg5FrfGPVs1LAd3vU
eqiGxabrmoaH+C8RjHi8haG2dgNfzYGfZ3FuY+vY/KSwBj4NB6XW+umONLcGo/+bPjxoKaFGDUaj
xea836TIbOCzdd0BEHXzpGbsHKnsgXFCzsjc6mPgzpMgmUDFwEjcvnTJJtXK79/LajKGYS25yKPt
nn01dlN+zdbzH3cY7WH7GaAyP7ahGNbWuMM/v7icqyP1RkoOZav95yMHXAAPEvRq5ooPCI5rKgWE
uuteiAVI4netSjPRZ/wrsphEro9Y3Z5CZ3+pA2AhMF8y7FqvidlgIFkTtQsBJyndEZbRrchrlBIg
7GbxUev1tjyK/MIirVGbUIAzUyDhnVS/fU/oGX0fF6zZwuKdwCeW6Q+Ze8WiDgm7SrMpPCk6MgN5
cTgrq/s1/jneKqAz8Lyp2YynXg9GPA7wtFDcMUIOAPELoJw+RY7LTzY3BL19L/fa7wJmxp0oMone
N4mIPErKRFfvze+6jEsJY4djxahM9hLCZ7VrRSmX9xQTTB+GTEYaLQmgRGLJQT+tTcXFIbRh1m7x
JhgLr7y6BOSmk1wlLVgAH7tyQ5f8AHtaT3XNvMyfPZxjYcncjAfNl3/rMnBwNm4GpdZBFqypoiTK
WMPAl4oXWPARXwuWY/BBzjs/bo9OMBr29j6Cnu74Ar1j+2Do2RzDTIHjp4A6vRjLFgHGN36ikM+R
3DpmBxnsfNEk8JDSFiFtF3sDvTKXo6jjLU1LooN6HmE/G/h6wlCs2OR96VibafNjhnB3VBkASzeY
0Sc6P3dkpaVM6QgjIXznjLG/fL53uISkeYdaAeH0buHyMudSwhAb/761ie0YjkA/zvGplXxH30Tw
QTpGeAneH0/zMnLjxoKDJEvmlSuZioYGvFKZRY8Fmj7ajW6DWI/cWkQEW/7NSJTDkA+H3GaxsoqZ
7ISQhE1vlsozQnDmBG2UZ5/LAKqtANAgbk/ZGH/oO3v7syPqox+IBvnYaVS+POYmcgb1AsQM6sVh
y2bnTrgvlWFF0Qd3hNS5q2VU0IncMGlImHGnwL2Ix9OLKPXj+Q40KuO1V0pwgrQMamfC3Kd4Ii6v
Syep/GAKRHKMTgp6iMBbNiGsl7GpQDXu0DXeXiuUlyjxxP49gUCSYuUIaHqB0rn2oiA7GszUEmJw
I2dOmcpSa5dTw4X2C3954KGCC5ngZ7shRxXzZnd+e37tLSmufyztYARJOB/UY47+eHf/HujB2l3r
VVvbmNIW9J9/3Pv9Sx2DnBAhZKOzDW9mqy3LHfj04z0bDAPVkFgXOilNPCUwqZq6yZ5gFFHkkV7j
XEAZX7ULuvYF4USjRxcrOVN7m8h1nGEIutZZmYGF3bJpdqb9Iy57m5sDbHIkCNH1v40vO1ncYZuM
sUPuHkmG8myL6YVMkUYUjpuIj9CloIOsksN3GwekVo/YweqVQlyvAVABCvBErXY8nW70PA+laJa/
DWLUJkt/PN1IXmegsOuak3ASbdzBLvVAvcsyUJ5hZCndVJ6s4/APi4VJIQysUlXhl0eYtJHm7J+K
dav+ay3kL13O3h+484+3AghbdauoRmwuRPy+rmtcIRXUrpusIoIS/j/zSbwJNVVb78JLIjypvNpT
xq+fJixmjUTczuCeYVOoql3gRVme+4DWyIVx7WjVOL6o+uTko/rkycMoYlwGVWoBrYbLYGjm6sya
XKYG9Ln46wM3hTn0N9c7sxSGRkwFM4EoJdNlWPhsMk4+2lJX+oEZ/yUx0jf4J/n6oj5HzTR2dtQA
RwvgpLuQUpALQbW/cfdnT6mD5eLl0O3Lt9etsGbbs9ADlrG2rDBeV/aeZXmOySSxzTKkb1wiVE1x
Zgc8lPRBEdjY3LXyhuthXgeER+JIIxm59CQ6Vikh/UCNC42YX4QqKN0FAWk8sziKyjhRRMyiTbuL
mR02603u0O94v946AGK8qmxzhFhvZTQEDVZ5iMm3GATRExTHuSCotITOnYIUq0mTVwTd6F6ODC0n
Xc+OvxO7vd79YBoQhA/aFC0eqhCp8nJGZqtzoWJeVY7VtGyaSPdJhXoH2FRxi2Gmo3UBgtvxDbVl
s35/utvgegeqDrY8fVrb7QF3BYaOSsEkCxIL0Yj+F1xAuDIpTGIN2BU1NWT2JfUBBG13xOAV80bY
z/6dPN5cgPCJ0W9+UORt3hj3A4FB3EJQfA8psgFHTbwcJ0js1dRSjNgBLrEwieYJfGC+n2uakWlv
+qkj5rKhcKY1Cm8I3hSK4EKKGS0DEBCPa+pmDiG179EN5iJxFpk1h9Hpbu5nT8wKk3htLsdje1/f
EKI0z95e16mC2YCJI4YEzXucS+1gUd2/lVoNXymWT5PAYCgsahwWGyla4wrxsmWbJKAuLf87mUF9
Z86BtrShSjo71jNerSbaNC8lzzmy43QbrIaG/ydpcy5VED6gBVSqexDaQLa6EDSBZmJLHxAsOPrn
WT8v27HyMDIG0vmnoRRWD7YpXkisqOeXgDvlRxLzD3Bugfjk2MlzkvYm4lVfNN5cwUTxv2MqzgD7
XUMDxtUm2n7fyVXsuMhtUkBeK9BAOSxbMOOo7UxXRHUszqHweSztd4i3BbvRG/3WwrehIDaoCeJ4
uTmPqnQfiHyePTXhc0lFI2Jrlel4oHtVrE4f0J8uv2U5IVMrTSCbN1FTl5VOnZVK/L7/jBlCnLDh
S4jInObMc44YZqXF/puf1jQcXw1SaYskGjGG7cFwq81qJcy2m9jlXQft3bgUSVPlh4NxbqLUkZ91
7YNY93ZUqrcsrgcvWXunhHtUkGZrkvyu+7ETFwhCB2mpfwjFZJpPxcLDL/Wb1wINBlMM6l+FeFUD
Viirh7W1Vw0SUOcqERks1w0TzW9hRO0WWIKP8fvXJmi8dkcObiEOvc5OSeNfIBmIbUBfT3XVukyL
2CaJNAhn8mx0EN0vj94dojS2b6W/4XAKna/1CMNa0soDpmwtct+kzTgwkwrWvH+Kdem7qws/vuHM
0F+Sdp3hVApcM0HGTqacmmBmCqi3bq+RCtvhoevNN20A6bK5LDG9PUAYrY0u5J18OZJTlBypgJqQ
n54YVqJqOSPf+9LjzPAWVtJz+2AgImuERihFjiGa2/yTlgw/KpLIHZq2Lu6ajA0d6k7mjSa9D14A
XHMr6f5bslKrQDpU1BcJgkmqRHGUA/aSuN5TSE/7SSuniO7Wa6UNcj3y6z1JzIAj/72kYkxyZzzn
HL2MziCpF0FsPkimCKRqNJfeq7jeTW1kqNRlIPrroF1h1Nc7EDZ8AAn/V5NKu6FmnPMG7aj9uejL
56rNTS+7OB32OCP/x0iSIqa7j487upkNOT6g+lX5ZSbfCXJ6237vUc+EMCTGYdnF0Jlxx79w6qW9
7VktuwKfsss2E26aijKEqBZmaxlAprwqh+WBbPmLAKU7l0t1dEB7JXmrIuJ0aT1rF0H+XwV4BXos
TUlAnWrIN9j2JUdhs1FB5H8C0jeuFXDaEVoSVu2DuwC3cg8eCcqh/zGYGb17mg1fKvHpi8cN20bx
T6HiBxeH1UVxq1yIY5RS9oTCIhnN8LZ4fmYdztUdHNuG0ZuYV1FxVHMW9qNLXQ33fukEE2PnTwZY
o6JtkpRdwxvSuObvoz2NJTMEI3HOzCN/c+FLbxfa0e8ywXd13ynANkzbR6Iok1A55ZMsONk7ogKG
VQGaqscS/aJ1JhSdXzVp3Sgm5c8+tack/OqyYBZn6lVgGiwxgsEulhLLKGi520XcDPSYsIsF3Maj
t4E9sJlCek0xokHuRoZSNFyNSNQ1rwO4p9mSiaYH8r+KEjVHPz5Bf8UPXmLuXQ8MmGsLqJw5rzuh
HkARYQcCscN5i3P/YqM0Ch2xA5zfFPFZWg6/p9juWDcXDQTonBRpTq6TgrVqTKKhTDsY3MKKYZZK
tUA30FEU7AjfUdaijeADhqjHSzREf6TQC7N89aNDs3gLHo3FLA5VXk9sw8207r9ZOkNeai9NLpjM
3Wu+KQC5TkOJOekYxDEcqXqyRfOKF/OuCnAD4eJrLg1tl2dLvdIuwasHFq05Z+A42VZ7JfggUnBg
ZfENJXEjPHYN3k8VBAadY36HUx8Vs1o+JsuL6esDUc1TIoM3hcWur014GEjsdagvl88e8lDLzllU
uPTJ+xU8Wc+sFA1jKa2QE/eEP2SzPjeGrDbWUmGmd+Oy6vuD167z3dk5gKKWBiV8k4uRLTEvQYg2
ZMUna80KM+rPiITyaorKOKVp8AszqM3dYJQeDQKIZshV3besIsAYgVgKwSzBiF+zLw5cVA5+Q7qZ
JCP5Ox73S+ZydBnilEPLz5/LYYrLAysGkTMDbZSAnZvmA4fyMKuIgJqagc7pFe+CH6l/Cw7tM3RJ
bWOxq50FIAkQQPEpFcQYebN3gPKXDLOwfRDtvEtbGlgK7eVtraEP6xRCEHppZVZ3NMfZipHgbA9a
5QBrvJrf7KMQCtX+PdxS0EQIjcYoyzWbAEai0B5rhKWf30otZtrDxdAVNaLrryX1vz+KSHR9ssiU
TILj1P1V+xUWh/Qu5SmBmV+dw99RNTSg7xJmg+0ax6E8rO7fI1JLXJluKNLOY+at+Xt6GoJSvWgW
CikujWHIpTXS02EU1QkSRSMQnCj0mjqU7x9qwxM7cToM23P1tSNHHwW7XEdiB27M3o+xGXyLxAUo
U1iggxeuo9NWimAshKqsC8GdVhpMUev+hHibKwZCaKd4YP63a1USmALHtqHXraQibH0eoX7ZjC6m
lqk8VoSPplBX4QBu7Ne5f6JrU2K4k6fVYJAwsFc35l+ql0oTb5RyHc5vU1PI+ueZGctfHMurTtfH
Ky8cHnMyGuyWkopFe44TITl/26BhUl3kY1PBFsqVZZv3ufUvkT74Bb7BuWlSWu0/+Wuk7/wp00aJ
P3RVqM4BG7TULJoaOyPQpkAtJPzdXAX4jIthWOF+J4uDsSwGILQscrrxf3OvNNzKsjGhTnkgXDEt
m+HbTu+uM1kI340Y7mpEglXFQUf7xS5uWm/FwJokDSdQ6LXR2KbSNm/rlEs2K3pzAYNg3aQ/vJ88
ctMQn3sXJdm2gbOO2lDPY8+oFsmdUvXI+dJCHU/egy3OVzTH/XmsY+fOR0l9Y2B/yXMLmKkKRieR
AJ9TUhLTS9ubs6OhNeFlPmI4JPs3zHoUQrc7dXkI4ZFNipIUl2udKoMxekB85i5RA3YEahpeBQI9
wG8nVQ9NO/H/6ZIP1benJxD9i2SSYUCHBmovcWVS8BER7GN3sJk6nLwNs0awQNqDp7ILaumd//ii
9kDf4B5fqGDH03FQ6PuZNsJvkIomg2RusfWIzn9bbmV0Ix6GJNvjJQZbflLuyKKJHiFFeYFFCkPM
qzlIOIhp84PgeWeAMV9rNAs7nPo3Yrr3CdDauTU9I+cBUgebyxGHUrmclI8X0NXbowVvMvAb8jkg
7vLJ+ClsUpyJ1v5f0eqekrmHk8NdcXvDow9W7A1FTAkDtZ0Z5UtEkbrVsKMhGkZSOp97hfWKtICH
zvu5U29oRyIK/pxgTJv/RZxuETPmCXFTHX2RxrInhu53Gkw7fZMUACJcl0wKxFF7dLZzwTtzkvv9
XSKHExNvxpEsxz807njw0KE9Fcw/+5z9E6K36EjitSqcpFbq/DMUkJ20qiV5vsp5njaFmhUhipfl
4CuggRIrXnjvgXVkbKTqoh+kygXBybXgT6WnvfSyT00SH8mV4OHxUAn//qcTG9omhh3DJ9IEG1k/
8sxb1c+sNYaqre7zfbaTN/64Ayp6nZlFjhmfzt2iQABI6agFiPk69zBaiWdODQH4+XXRQmqsMBaN
XYWFA2plOl8+bN0KDGndUqpUSLBb3GsgZtzCQ+FhF6rF/iqFuqcg31TeiUVc185hPxraD5ftiuia
ecYAxO9BROzi8RBgMF5V7R12y9PZkmcB9pSZayLPnJSec+BtwWZEhGwR2g06E1tarF7UsZFv7C31
IK+nEmKVlcB4/ZMgdb0nuBhI9Dr4leNuASoeK8xljFakcz1jv9PYJ0lLjDnyfBQ7oadM1nrcOQsB
usFxcXklzlmM/mp5KFGwzAqvC1FMimyX1jrzcPobLuHsCVgAi0qNRdL1RZPEggZ+xafCFTXkMbCC
cLjnfSKNvLxi9f89zYAIsdSUp4hGzUMgps8UufIERLjXXICq0RMUhT9ws9Idlw6zS8g3z1H/Poy/
TZCyq8LToGX3HWf8ogjcbU/2WcZeuB0hY4vLIJTPgC+auLsFp4IJIRYMu9AhUw90gmYU4MQWKydp
VZfwPMEmOejuj7XA/ZF+XaZxp6zEtwZJWlkgxJh1pYi1B7DXpuqWPaP4eXoBjwb9mkk8NM/0/P9B
RhjUW/VgOnwjf+G4jvZMjXDeG28L8ISn046i5JzY6CU2WXsQQjtnYohX4Kw9446tGFeF9YOxiy3T
r9O6lccDn+JGzxq6g6wRZ2W1QxJ/pxww0hhf0CyTP/LGdTx7oQcvvATfHICC5YOyFnXRBkJZmkZL
OG0x7k2SvPoZRrFsCQZs82xzAHT/chLczQrEV//ZVs9V/Z9CARdQfHTbPjzivhuWmNQ33w2lfcpJ
wTcTPnitV+S8y+KSfgZ6XtQorxJh7EVfmkI+uRS7Hfdy2dAyGoOnjfkxhVnzpseL7PjhLl4eCPXl
NPHzG/fTSx/V/qbfCy4ud6wzybQWiyhDWUVRNfuBFKumuqMaSwrpHgNdt3hKyuGLhDKH3P3UtIOX
N+9Lk489mUS20ZJBQ/wUag7zNjIf9oO0pxNBelb1/TVx9VF2mPvd3e0CHYE9H4WFi/p80Hc/dSgu
hqyqQW831QGsd54+tDHcM3HdXY1hAekKza957xajw5kzb1t6NlK3imv1sSZVDOOOoq7YB4jUcwPN
Af974huNrH/ZqUJLRmUQU3LtamYhXU1xv3FfS4+dj6lx6w7SX7FnWHHWob90fn0WBrvatALDEPe9
4VKB6pRnq3607KXbtfXFNKhYQiQcdxQsgDm+5qXyqEohidDC86UubxXX+dO7jfti7fDtaMshloJk
C4MUmtR00nLXWpzuH6ZGWyCszJ5iElRz4wzuBYsTI4YAeT0hMbRfze4ue0nBCYHGLDi8gdjVUg8y
7FPPP+Yqnd79khdzgaIfcnColb469DveWr8DQrE2o8zaUn7snqXiJuros88jXYBgUx3ZShO1+PZk
PsPC0bW4FWhPOEAxKtpTDt/VGEDPlRV1+L0DIKBAIiRZL7Y+Wa84cXyw59iE87rWXCU1RqTgCCf4
LK2Q+ZVIBQU9MYz4GDPMxp5of6yrZPkw1e6jMmFZu2y7ILfmpToLouRaT4FtYNFdlGiI+COEbvmr
BABM+U7s35TcDcdCwm9s/UWd8+p57jGp79pywm2PJUMlE7du7ZWoebGQlSbY+OrgHnhToFeiUHO2
bG/X7r8EMApXiCRQiGj5a3sYt/vEYYjFJgEX6cUyJFrjXxv1ZNY/Fx9PVymfF6OXf5bhWJuzY54A
2nWmi8gypnvaIZHMTT8370fwg1gZzM9fZOoNliNfbUsP1vIgIAqMGK2LuYaiO6a690pY+iarv74k
3ANWY84JDsndoDhjnh0fMnurWa7AzXngi11MCUznLzluLgQtt0azyH+ZDhCaxwRdcU7MO1p1nelS
HHMUmmofkVEi/jy/LSpCW47oYNGwSi1LJE5NFTdCfOl8OQc3aFg9Z2on3/irt8PBdvwHs+a45k56
j6iCYe0RLjEPQy86RQi9mXIpiOrmq1sZB+0WwGsy0sjCNig2/fa8P92O3bA35x0T0+6rjJC5e572
kZDFevfYI/VRlkW7fnxv/03DVfIpC94qnAmD3bIU/z/e29OTg+5cMG6zVWNRGKvEtkoqM+KkAHPW
kqM64ZSyfHpaF/HBh/yzCWQ95f1ekS05TZwitDmnOkghNTbDtrBtr0LKzCqfCID0GX69cSaiJnFh
v7JbXzXoYE/exa4qIgm1vgphXIsjwj5GAYu/FArQkOrDBmg6Tyhp8p9EBrSeBOkeeIkLQFqgjFBG
oVL1qVlSDSNKB7F3wxwRHB33IeM/1UAAHK6h2n2qNbv6c8BBI6btUeIez7ewma2rS/1g1vAMHxfS
wBi8tczLm9980vMVsYJU0n2HASojO+ZaNUpf5HeVMfhar1zTvClm7Ucpgr/UkIFsC3Go4oDhW++X
YsHzNEc6HNOh3juzGUIMvxcyDUaRaSTm1LDRbw2cTVd4Pe3RIwLca7L+PrEidygAKN/JsApyY3Z5
p0KD8YbzTYqdG53FrLc8pCZ3Jc6mCUTvG30mIGyx7HXHwfFCBHeUjrNkw88frSqWg9NC2JyjjsD6
8QBUllMX2occmrmJz7dclbfgv6vDgUyDGH3ABgT4AeRcCkpVN1xbkkCv6ACvqurEPmhRCpV69oRZ
akEF+2YBK4nw97u85rI1pzl1WoFN+cDVFmFvI/idHsJxgMx5wYwHtjT4rB0yV14XbCKPY15uCwiE
RMPPrcACqq5a0sEQKviWfnQ0c9N9Awh4sqO6DcTk3CLYk12LpfM9WQI23PSRgABeD7Eq6dfEP0VT
9cQM48pgJr4BF9W2PoTrWc27JAWn4a6rJHxoth10jfRcWYU9xRu0zFWZwWqQmjkNE/I82f81MZD8
pIDEndSncfiHUch9+oJIw4dSLMe9spbQ6mQrctkLXamEV1eBxd0jmLbEaEGDROLxN11YIqQhAPqL
yFJMQpiN3rliHmsemhXWzNzv9n67n4zFPkk4v/MIaP/HK9amdGw4N28HkzcaBcvgIapkFl1I6R8w
TQRQulqhQL1fTXaUQuiKpAfIVT9otVmGdGaqreOg2ghCI3d9Wl1/hYnuTyaDRSVG9VG7bzH6fVk5
MGp1KDCTa9kSG7j56yggcRvIdgAM0B0vgt0c2IDxVnR5kfqJPopRbref6iqXkfaDWONj0C0Nl+g+
17OmhoJ6gC+jT/V38Gg+PzlUMmS6VTe5tbpEviHVOj+psO/qp3RtnMeojRCwGWSvEry5m/5GbbYr
LiOPvfQWv+RAzfFfdmPFTiW5LRh7t/nHbFAcYdrmCjxGPSzmDhZiqxmc8OBQlEwurAMze4kLKqnc
uGerFovX0X7aAF7wKLT0EE4hoxazgtrnlAGTYySpMkfY3oYNW0mIoadGVtbaSSY5BbH4bs9Rup23
0GYuq4HVAh5jkhBXd6QVg/PaFvBG4+J6gt51JSnb9xWpw3PcE/Eg5jE5wub7EKx+LcxyuAAAesfE
1RSAa1MqsTaI4817PPzhlvd6wuWhng10KsMilOOdsrbt34EZuf8nKWgD/OtFx/FkFTohb8CsPA1z
EIKswTrwzRDlzh7vj2LmpM1i5FL3soxKtywFeqv7rDUo/OrkTOygUEijMq1Z6nEO6xuqfsGL4hvv
oBbkYFx9G7p2E2Us8SnJu5wixPo/AeMazPv7KysRUawE7e0561AudTVEWqt+9aya9u3rb7zCMwNy
0Ig82qUB5+9/wAfIJ14bjE5pY07yaM9xJB0f8oPzJWZS22eeGFSn7TVYR981AMNFZGp1YswUAZBc
EIhDA+CgLCzUpqkq5QeLqpsPcjZHOWU4wC7O2CHqu8EAEBsEo9FgX/CAjb9gjhdo+YP8VdN7wz05
OnAbywojTJTqW+sD/UB1m/8M7v4Sw+LcWK48PwCZA6j9Je+Wk7QJ4z8J3u9K/5R0FQfn3uDjxIo0
UU6gSnf1PX+Br0/W+HZ17QDxV+vRbV+mzSwvUEfIu21kzpfI8VGoEnyUxT9Qy1nSbNKnMAPPYLQP
3xRf6X9d7bvjTwaJl4sVBEl6A66dEszhd1GUVMnXaiQL5mnwE7RupyKIVs76rIpZJYZB7KvXCgG4
oT2FJmTqLyPXHjcMBiSk+LAsp17+6b6kJDvnTvFj/39iCNcnCknP+x3IutvhywmALjgtYuyMzj1K
2CHf7LDVK5g5JTRx0jeoOYs1QJgvjSd25gNroryetLuLbjOZZIUV4fcJFc19RIzSIAVkICA05/ID
JQ53weF+jxa3Gybq4vZAUKgtCab0fLVrsh02h1Qf4FXImrDTF3G/lNVamgmYBtj44HeBXaFLsJQc
dJxesDMow2Ts5fbYpm1NNZ5e283IfeAzqWqr1f4+50Wz3DaIXZL8Z3qoujwMSZiv2O8n5LA27UEr
ciUB2BfdgKyV5CXT4Co8OnEmoHHqIAuYa+c2hOhUxXdV8L536fMNRXGCp/8kF0+0rqan/Y99to4u
NijyPXTI2qvNGV1CJwgdI/yREcYxVjh9gPIoaHR7D2a0VWvpj16jrxxj2MsYc32uSBWnXEkgt7Ag
JgwmsukXsn9iHif49/ArrkYqeb9mnG1G2DCtJnOFW7IE7Q7T/0SaXRdJu5UsfJ8yNm0QQzDI3fWn
XcyFt4b42DBQ7x5JICQgtMdDWNc3En+EhSYbzFvvMuBwJ2I5FUdqVZl+Tnz5eXVWFf5MYb5AUWDX
BVGbVw6zsfwakvNVlwHEmhHWQeFqUIz9vDcnQoUC0Ah4QeeRfi7HsDryKbxixaDKoKix3vFcD+9b
QSvlMDj46UzgATGyZw9ZO5Q6iZevM+n7EVTxcVcethwWEMV7d3qI9phAThtI1zONZO/nxZDA1TVD
pc0Ga++tUMQFBZH/JDCe+tCXWiXl3gVIJsE7LlM+s/DfE3yQfKmFzfyvaPWS5HhqN4U034sm6QaG
NpRcSQHJeM1tyIivPauF+5nxuP6RWqrNJ8G3DEl4C9RTvybmI2r2pPOZaFaNuxEMqk9dbkttKfG2
aetpJZvOYx68oI0MYqplk/qsX6mXtuiz4VPGE3PsFQDe/gUUNmlHbBDzzoU8AB8i5nkTfRbDUQ9S
idZYyhvUjQlNHDN8Sy+/Ed/vuym5DCWt+FNkEiUXiyoJawY3tVuybYDF8ZUox6dFjC2zpGWGtQQZ
7iKGpNCyyO/O18LgBz+dbVN481+iHYlobSHtpSivXYKeqsZF8eUa4hur8qb+MP2WoUIAwMrg8Xf6
wvqX/14TB13dSAtmyxjHcup6cfBNjpER3XNj+SsSUYtyP9aL4ULbXyDjQ3ciYJwHNRrAiEdI5gG/
dOUfuJ/9qbctjYKpreRlpC/7/OGbIjZ336D4gf0qgnXoQ/huFqsfh+a70d4uspN9l6NTDwvdGNsO
Pa5m0+tT01pl0lEGbQV+B3hivO2ltsoqJFmKSEkYgc2nYQTywns8xpxwBtZwqeG6qsTPmz2L8VSa
q5tiEg7Y65hXeAZJ42f8k3rVYeZjOToqz75qzoK/t6w4OslCLhpcGaIobwzxVVZrMkb9RY7G75L7
EKoyWGgsXNhyt+BIch4SyRg/1LhyzEX4cPo3mtBG873xeITkFiBRrWsLbDpxL2B0wl+8LG6hbtz9
1EXlo1DNr0ctqfeV/029/+cLTpML5Sa392oXLJQkBfuCrfxy9Ck4XdJxivuHjTGo49HY35BqumOQ
FmPJefFztxivi1pyZvOQ2G5DLP2fgs6cIzDxUp5TPLVVkOXtU0+ztZx8xy75MI7TjZzlQxOOJqg6
DD9/9kkCc8OpI4wCWNvwAsgyQI5QnBVU6ZLiSBny8p6p1JGaEVofn+SDEdp1erUMkuxyrU5kebAM
ihZHcTLwf0TGMxO4UqSZfoSBBPebW2PXNl+7dUVU8K6RVrO25CfIODWdFq/5c/5BMArVUcqvMLv0
VeVWUC1s+tKawEsyq24cPvksBzn1WbgNGFCp8rtTZPsdquqiD0Q1Fd8iMfBXADvM4588d4e4ASNT
yviVe9v5o5x61BjCIdYeBVHlTGJaekGg3VGuxLmqW1B7lzjz5j8Ck3l7oHWL6WfMT6iH4hC85dlP
SJiy/eQo2M1LXLepISf+QxSa7peo7DwHbS5v7eU3r1IYmdd51XNLr+EwVu0Glkv50xjwrUxVQtZs
IhwsxXTmFCI2mxiCEdaltju7mDkko34xgNSMA8Lty1O033PP6kMCHDNQwzIXWCfxFe1+9V1svS1Z
WgV+B4t4JCAT7tqO/uUDgeLfmSXfK4PSjIDl8hNPieUKiVMxialRhqoCp6xytDByFjwnlNgo/zti
xypk2WS8AfLzi61ZuXP/OeMprdribFFfXlSoQAUI9iqzMdPCakKCEUoS+HTpF7nNsFRnexj+7//w
m4/YNJxBDBxn0CwFN/Upe2sDgYnvEChYtqWk5g9XgHRUA+xMkaEOGa20X0yqxURehlCYS83MgVF+
81nzR/ivr19QQKmVvBT2bHxj31Tho4sDNvfJr5b7YPaxyK6dPw4HJC7pn7fBV22XcznjbY5KVHzy
DmjOoCLmLL6dzD7fYXtN2dfprH/lIhEhJ67EozEiFVnj3O5FxAZG3TAZ13086UfPLSeo8kb1xKnv
MNN5/hswWd9Y4NWvQkCqP+t/JqbT7N73ex0QfrlbBV55fZCdVklYXcft7vHOh4kbtGCYHfnZv1u+
yVI/51jiXtDUv6eunlnoyeN3PsqrGkDzb8Qh1R2GML2gSyPWD5Ei0I/jBUBNbYdn1RMrZNG1iJXf
NEEiMQ2wTPnB74hYppEmUuJ+ItW9PBjWB6LoYWuOEZjzAmiIrmpOAR/WkY/P5qzjvO/3JNdwDAzN
l0wG8goIJB2mffmk/xSyYSLUJEa3SY2eA0MgkcbCKP6vLF9sqwfeTNdrZlH4G2j6Tt8lKYXJoo6c
7mFlr5bBJpOXhuvumx4H9ySnAhNfzPpPVOrHsoojSSUaOouihEwR0FGVwX88ihdu/EsXF3XD3qAw
k+botu9VLdrhdvoj3lmMl/9+0Z+Sq0jJUxkQoO05/Ihdn5czANmbppTJ/npRvoaMUiAWEbH/7dzH
I8rADFiaxzbqIvyKEq7Om3bQULpeiAr4kJaDZl89WMs69elC+rnq3n8H2Qtrrw/4tkqHVZr2TgsI
e/illcMKBLz+kDbwsQi6zH8dSnF0W3+DzO+BIcKrVitw8nEv0ZIGtlHkdwmnbv1Q4Ej+iSHXbRja
aPWU+M7WRzMH8zrOjybK52Bu47auJKt/5VVxWKVrEWp5U/+jTY8tmbP27AtbINSLqkV8Ct/u+pvn
/9IppdhK/OvdhcmSd2CXsUimTp0FB0Vrv6HEDlmCtdkFX51ThUiJPHDqeTseLixJsZPHc1y6ZRd5
YtmFoPxgxQfcYYLWg2LUDwzD1PJGEseHrWO+NS1UBCPJEFXw2m4sDpAVupftPdxWjylFGIPGGehN
RnXCqBCiDyprNwTFIh3eF2LVk9zLZ09CDlsjpdVMAi+mwFHgNv1f1HFSfq9Q+xMr61PtBJHQtT0o
/eLW9ZMkZaZxZ0YAA4c4RhWs8DMKGghrHDuzzGT8z/5XUhXP3Jbe3pclikXHluiuKHEUa/xRSzCW
AAkRI+BJSVHppBH8E/qVIbbDfMc+2onYfFH6zUWqHo2hlivCNQqrGwHQrhSMpmCvSetxuJjQyd3M
RSMZSJgLQRgDry2SsY0I3d1ZNWITGfnx1iN/0itghRuhVHD0SXV0tlGuT5OdK3MshtskqU/upD1L
bid7ja5kj5N+9/ZprVlKrsKiG5wOAtsZRr95B94XVq/TrDeNqxtMXH6As1De+EYBuErMCwUDbxa2
YtzlDvGfPTFpcFRvmj7t6UbDRuF1e7CXxuTbZ87w0gmXpZcubMELYGt3V8bVkrik9Flje87aBI82
ACLjdxxmf56SBiVLdDKL/Mdu0gUO7XG0408E4/6oTiM/jkYnl1IAA9JiSp+5DeJI2e3Vl4rl5CO2
rlfsKXqnNGoivpIPwzkyeTwdZ2uJ1meg+ScfZkXTBLeBCsXD4M2ihAeoqmuVbLFV+OUMHuRWKYyA
cwdHOreerLJTGybFtM5t+dtZB7PKIUzynxn2izTa+f+yVB7YcOEYuDboN7uP/M5Ax8G03LDSOjyi
YTDJdlVC7/y7WB05cEACrrBfSTJ1DYyyfOyKdKdVjsVzj0uEuQ76mJCatTwGahPqa/sSYjyAEJg4
itXNiVyK3AW6zYe4QVHT67nSu+iQTV4ZPgjpiEo9bO15OlPFnMGWrrFhPTG4BLTfsPcfHlET2UkT
M/WQ0iHU7ySipp9bpUi6HaLi0TIfEfevAZxd4m3rcpT7ohftUCFUSrWPunVbd2VtUbgID8L+1ipt
oHSQNUtOX6ZIYI+jZGEBgbMqXj+kuMTxcVoY5DNGOujrhJhwldoMy8NYOAdjW5nJv8afwVh9Zybw
exhtixaWQER6/pRDvxOFgH5IeJt65d1wuHCXOoj3IJ1/HpKnLBFVgwg+BR2kn63gz6LndJC6odwf
z4mNXKB41p5/m2BmhGisDi/yKtK46cYFSQlIwOu5QxDcwk1BhDRLAslMRjRZZOgh89UPU4NJHdO+
Al3GZXtUlO/0X8JYlx5yeYubIjWtVeIshpDSb+YDBT7oqPMXdMpyvTPcPW0exM7c1h53GUKV4VON
2lP4pJNL3GcGxnGq1WkSKy3395Y6+FXCkQfhXxVz6MXzTbQBjTSqMIvFYv2fkFk7ypeKQRiEGDbG
5gp8QqaC60z0o3fhWpYo78AGqn8JLTFahC561i9XPTo9iMSOlmBXHLij47X28CkCbTSk6agf9bFI
nfAQEDaCzciTBHsiCVvxStF3Sed4+ITdt0etH6OzCde3W+Bvj0ZqESZKiI/Unxn4NQZxOlfB2lfo
toUzjZ0z2aXR+AZtDCQgwbnqjM1FXHDw9XjsU7h38b2RO9B9ScOcbPbSDjlkfbbOeo7CHivaJM4Y
5LCxqDpDM/wSIjQ2SONwFk105Q/nBKYR5c9XP5umOWv4u4YtxFB1hj+IS2f9txg5Lmn97lU0YdD0
18ruNhvNZHyo0a8e4mvxmkYkmHH8ALtIfdR9UjYHdavEtfTIuRmIGnAMGkLi4EBS+S3IJgM6PhLe
oIwDD2Ww466xZ9j5yZUNlaQYVFRxOZ5cAm/lKtgB5KyHQ3h32iP6nOoVJNVYdn4O2lpCefDQxiFE
skDws5SlvLopaiIpKNrRl7ju/fG6TzLN2zDEKrPilKClamZbeYAmv9Wa3kH2yHZ+JkEWWYHDcPqb
M6S4zkvW5cRnSDEU86KFh0Ck9UqtjaBaHXlvCnCMB+I/y8x7HJVW+uCp6VA2+pMGw7GcHLRunUVJ
Fzq4flbgOtXpMjTwFVkWu3M4sKPaMoyRAEt35e7AO6J5zSYr2Cn61wI7r8sRcMAapCji7Ex97+Hz
ATqGtjjehdd1xDZ0MNDTFLrctKs52hD49mkzk+8rlJXD6zHmIzSqa0lnwd6i+3w4sSmCHMMX4sEm
8H1YQd1yDBBuSyFCGnMqVO/8DSk859M6XAxRSW+TQ6QDAjalP7YWXwQDdDkyBUbLFQQdP5WhxEUt
h2JeweDupRHlKQDzIUOxXYsCnbP0IIQCd+IZ2VB7o9HlLyaFEXxv/4JdfZgu0N5IsH5MCgjKCgkn
uvGDPzHvclt/EPAb8cooXINQY/Ykdv/jtfM6hUP0ZyO+dhE/SWTmZRWGP4xNZd6FFMULBCXyherJ
auYnwg82t45d7zG0Oudi7kEq5YPTuJTyFCjotay8mNwBq9FWzSUS/obpnBpFLLnCdDlki2Xi5N+V
krnPYuD5+hOC8baOYAaFki4axIZo8SgjjWDGB2Ielle184Z6GiDkSiQfO3kxGvr/JHfvWy4Tl/uD
/XOuSmP4fGSQY3T1DcwPURjigC+GEGd0G4ehNIEvOwnAbmpL08Mgq7U/xEN0oSLGSpOYcwjmPKC0
QGK7NmfD58UIZCzrlhpopWTouIltcDfyNBG/RD7Z2lUuLbl8Vii9udqdRFKYlpmTNtvifFVN1+wu
dmfiGkCi100oO8w3ffhoJ/+FDXox4JsftQpCzUVU2fyd3gBo+uWa2sDLI0gz0jfsYNO2z2zskRTX
h2qBqyE3LhwUxQRFuBIFl06W1Swg/ught7XOb5UH1Ba9t8Sk8OQopiT5e+mfC88ogHz0GLYzhNH6
qXlNScYpsZrDtnj7JO0FAbmXAp9NkXkBsLlV8RO2nObeQixcU4MsODcNUM8GAvWeFtI0ZTV0n1wF
dTyv+A8FgOg+sLSm/rynfbXY1yI3dEWy+AxgCSokfHmIQJqSryx8ZltWdw2nuRWWajNi1vPVKHP9
BwM4g/ZdvGdWjvjjRqbRKP0KwxSJwAhABGujdRomIETdXjHNUmgjUQmWW2EEMUh9NnKN1kOvMLNi
OY+I7EF8w5Sw4qZOg+12xcmXhL00Vo02ygy+Fl/kaOlLPBUBdLqKs07MmCjVmzH5T0PflKgMwaMv
+pTdJhwMMLjjOACyoVvujOWgZXzrcQ3/Qok2SDUmJIIdKuHxU9vTSxddvECqnhJvi5i9E36pbVRN
mAJec2qdLSxgbQuO/lcDuqM0bn7BZoyyEEi/XqsrkZsN461JflUsg73bCZdeJt8lgFV8X42UnTfm
W/VaBg1CeuBqiL01p4ayCYzQzZqaU8HjJQMoD/yQI0NMTzbm22uLrhLufVHU5M2RY59XfftaqBJT
D/HnJ1Rkkq7FuZ4aBvybYtrgNQTSbYPWlz4V9sAoHcuSTfepDSpk4W4M4P6hycNAQP+weK5UH93a
NUjqzzPYcbde0eGSDpWo3GTXJsPqKOJg+jo7yJc39T6xNXHXXbZHHbbCBHrTlaURqMOXAimiKRuo
Y++hn8m2rkBQGQeWLNHsGPbWdVyvfbcSxL4p/DdOQWnHB7/uq2dAqPeYsokO5YAzurAFpZuegRSL
vcWvgbf8ANjq7vFimDJyrfaj8VkIml7nDnjy542RmfxDz6nFORRtPK8Q6O13P53kpBQyz6NTZAZX
nulDMEM/wiYMPKEsSdIzzA/bS0XMiJs+E2W8rULznh11u+D+UBh2QZ6U9LAQaFe9Ju5SwS/knsT1
Uy5WMdZm4UsGRGAyYnVLSyf6rNsX9qeC+SCG7Y4XKDjd81XCEaTYG8kfrc8ps+bvax/3lW3tbRkN
r9LVc8VH/Q1F2cQU1gvr5TJ8/shBQJB3L8RSPFaSppkol3dCp4Wvjr5/mq4ifr+Bzr3lyf8YlwuZ
W62rAt95va8S3FTlSxuat7XEB7wp//UpVXJHiPvgUS2qu0QKe4bslvuer+n8ex2a7ILZJAisnloQ
SsZ8sbJwmKZKImbJkTWRp73K6naiR7chSNg7BtgyJd6fsRaJeWz783g0Te8iWFTfI7iko0tbQZC0
T2KbM9BbJ0UvW89DUwRb8wSBbCAjwwxqxL3OQUsdkBmX9f1yvnuanPf56sRoEIm7ImWIvnnA4eA/
jsvbJpJJ8C8HVfHRP/laN+O5Xeci3dCYNnSdt023ZDLx3NF19kT0zmrAIQoerKFT+SmGFKk7ixOF
Qd6SHJr4aEQoEFNsXh3U1Z546jozBAEyJoeTNLwIaP4npDPDIKGdGLplB/y/sY3u7yB1CLOPfwqH
k1g7O1Fm6nY1dnx7wgWDR5HP9F/MRSsvHPCVGlNG8d0INT+jBS5WQ1KcNWyXKyVe2Q7Kb+MwWXwF
5CrW80jQEkt/kzGEQDAJRNjItRvvJ+ZYxWUfODOtACMXhGxYL/jH/MjBpc1yfOXm/8ZZHkbBT2By
SZuue+AQlApJM3o5zJBULlc8yr77Stm8vuNcmTIVXMpqQCPL0ugFezo3z+5mIkb6y+4uxBJbCfDf
7MEVJ9mWWKdk+LkjjLC6MU5A3flBSS6PeMCA4zBVv6kv9MSJgW1IceI9ic6GOIOBKjfWdogjw7nP
1fctxrFG5fSHbrEWiJLVhXxScGclpsV85QUQAEnfTNc46fyPSbT9rsFzm4X6RmMjfbJ16qB+sYma
/3kebZCqdBejWUJLtASNUdJ7gS6TgRsFzBX96uSnepY/qww9IQ5SXFxPd+VJ4ZTzozxLJi7of7sR
6ZHzkilmdck15OR2rIuA8L7ENbsKJzvYlrq9Tmc1l9DyuxWopT45UPufwfvuGc9PwnptTgirz3Uz
kV9vWVMtzN/NUijVVE7YQ8rlCqEOLPufW7pIty95sSx0aWZcvBEAZ5hmyQMJ42lH0YDs3cvisOvf
ikklISnQ7fW78TOAnj9SBJIsuCoMchuGnKOlZxsOTDr0k3hpvBANdMr5KkObthmey16SJjLH0kAn
mp+dpdvG+eNPak0+BatnNBsxof+pby1gCzpyTXXbtegFgucdllXeEVx+PAA5TwAG7JGT2I80yoVk
4bzwUK4ZIJ5fFOM/vIzrOf5gkWgZeW2QgSMv+D65cZtZ9f2m4zgXXAAL8FcO33mjGxHuuezMXzC4
Vy2GyaawLFOnbJ7Z+wePq93B955QZ0xWHXl+VXeYeU8c2nXZPlQo+NzZd7I18k4pjzGfrHRRLwuJ
kj/NkMsVu1SNUrADA5vUC580F7SsgDj5bNlOQpw1FBsbEBNK0v3Row8P9C0giEvGwrpPzq0gWHM5
hGVh7kCfRiDtOC/48458KYdTA8zgJEWxddUGtETT/w+zjvZfOKzySORS85IHFH/onmuH/8BN4nun
dJWC87xaf5B24CY3C8ZMz/DlaL08GIl/1fTpvBQwuCkBLk4NiOU9jg1nalh4IdKqjIELn4ZRqnJI
Xs/t91oklstWRi8cIunWPM5ISHKn+tFDxfbl6uxOkk/xWapxvv5vNU0EoqyDsvNhW2Ci+UVdzdJ/
nmPPJCNwFkazQArtQXawoaHmlYDOG0m96AnGHlrI/GqA56w9+ManwElhKfCBzn1WuDZw0KnSFtOS
2ytPTmstisUb+kLcr9FhYo9mlLSQZIcVDzZzdvY+GATKwoHbKZ62m22a0KXdRWYVs3A9DwkNWiql
+l3/ni7sFlfL5+n7jWK44aU0C8lLxGq22aPfC0+I+8dlAsIzKdQL2tQKa+6HjWZvirDrhwuOK4gG
q4iqaxHQqmpVGeKl3a9UcM0Ni+2trFRdCbFnTIOUlxOY30RPSpokrkTCvw0movn9Ky3qbY2W1fIM
4eEtKLJ3W2XZyN+IAGuk8lR4B3H2Iii3a6FVYhRtXIKNtI8Sc84XgR0DCPO5JROkgK4T7uKh4cWW
95aQAnTw3nsnywWcVeYDp0vsAAqsBoVfuvilPfqzrxvaEVQUENtF8jdqwtY4xDXVzq0FhwShJsau
11ab1h8Cx4XSMYJFE0Yl0IbvfmfZPaQH04AOnW7vF6By4uLr4Bqr7C/IEvHGs4bEmfs3ufEiTk25
1WIEnoSGg05MEJs90H6EUCImIC/aSuFOnQFU6Zs5/pu+H5NIxq00KSfQaU6erv5xLPGZmfZuY9E6
4HRyt+UB//JztAsJ7OiaINT/t4vWOasRGyNKwpi1qDOvWBoTNqcjNPWwk4UbSWMQ/zpSMILdsfxb
HPURbd/D6v4WJeobOSyYs7qe1NzTzHtIJdwzmm8JcuUReRvg1x3Ws2web16CluJSZSLqbyLxP3OW
P+VokrF4jwoNHX22/4ae1iXyB7EaPYJpUUQ5DKomyTbA3e8gvdDFAT/XNH6mmzgpmn4nthQPdi/B
f5kjzmDoEqmwfEUdhO8STr2YEqsUIdYBUB/3OeAQGoCpqXDwPtoIQOpRQeZVrcYW9m83Zg/LMZwD
aYeIDrhWjera8Bqz+o9kejMFflshiqGnBwRKaQAbKqSlnLFb5pkAwLZ6dw5U757u+Ul5Mvc6likr
UyczmozI3Lv83lNyNaquT9QVrpAOgNTQ8JggBZRFQoTUdbBH0J63z0x595r15nF+FLBJVJnPfAVX
PB/LRRjN3r5Ta4yYUN8pGgu/SoNsvDqwyZ7KnUayA2sznwJT625KT93iNZTZQHEPRUDCuFTNvLkH
Cv/yXhLoSwHs+5+5hBevhnxYY/6+5b+yUxf9gKM9LHHhtnOINXWwSB4SHa6QExYCIM0TUrBWIJsh
vRoyw1djpyMmrTA/EcTnH4HDYkDqKPiCCQAkCaVwZ2/UYjiPggZVQg90Ksh1wwRb1Q43jOXyo9Yx
K6re2RJoUiilC1Mekl23/lC9e4wsDvUJHupJ30qAeTLGo47IRVcrbLQHQ/Zl/atVb/9kxRm3Uj/i
2G3Az+EvRkJrznbFrqDxAakPp05BOGpiFMQg44kPrFWiN6sDmuaKGjSEHa9xq2Nici3nU1BVcON6
hFXlPk3Cq8gAtieI/Q7k+g3pzU8RPBhyjaBQAB1oMLMnHqpb7QFbeMxXh4RcqXx3e6pzw1B7qsIo
HoLCGQvOHzI9pJIQI1B3mZGuSsh93ABSbOGtgFA40XoDJD7LhuUVZcRYGe10to7ltWz56EDZ67Zn
DhpCJ+tDgEnHNWaGy+D+6UoyyHaHGZhuSamAARbDoBqaLavf8WmVOtjqtU4EiKhCoWf8ORGCXdZE
Q6/26+t5SKGSULTFGctLZJOxP58USvUwE1WF6dCuz6UF4V5SHVP1LV3Bhp/VcTMnR22QEjpIPp+w
7Kgtrz8BNYyO+yxTS4/tg3ozYeNDu6xgY+0YQ9COIFxk+upGtanLzqfPWeYOYHxUJXbr5EdAUoU7
Y8r8SqPEDOTeS1HZybEq+84VRXFxiEoOTchhthtHOIlSUtzSur4i6CJaMIlHuCwJElL7cCrj74JL
6rPK9DUucCOGQAOcsiGA8Xbu+VXkMrfIBXz+Q9P43PDjgqBIVzPEB17rmzyOB2h7PhLSi1t2Jp2Q
uK5kiiLmIyPea9UmUPBaNkHpSXnOB7cqtb0URxc7tIf3l0A2uqbZQn+hWq9T301fnvoPQBXeZNox
wzRjzjr/jukaOHv7p5vmlcfDoMV0lcQvFTDNbwrECkkS6v1FN/B97JHbyu/Rh9M09JG/se2Wi+SS
G544EGmZWSHadmCU25955faGmQMTRaFBOWRNVHjlZQsOwonbtSdK5emodOBZYPOoxA97aghS47Sx
r84nw0eOrzBYljzU2dD/mmcV7QJVZ3Dj5DDLX7KLBFYhkqGgPOvgEjw4qQVkXguGX+2EMiHwWdNs
DYNosqb56MnJHn8TA8KzWLtC5eEuvzIAdDkTTnhUstJuyk1F6jl03dVzUPwHfy8Hta9qYWA5tjQx
EpNTAHwBy9nyYhWnztKRzx93UA/mG+KZjiCtOPp0KM5J+nr3xEDMgZDaSocCUNALJjCb9SKIeoHs
Pk5s21YveyKSeljFfDrmPCZVMl6JZKNG8sMfYhmP4SalF+/KmoN4G+RSPh7OdcZZ0j+5nNNOZZpJ
F+vo0dgjECWjHuxiqRhY88MLMe41+GVsV12DFKnqq20F9oD+FqNZoPfttF3TmYTZrrQ4CtgyrTXE
mj58rimVk4gOTZcWoRJeb4bWHtJrZDhFeYjSvvfWfC93++Uey3EHA9G7sE8joguGWo2Z0J+e0IQI
Xx/sd62egL4ZULFGpoYPkj3sxbYi5/3GtEnIeyDddUnNQZT/jdzD9jRfx7/nLKX3YVjc9xwfdqG4
wCYpEpArMqaK2GW+MDAB7Qr+Bl6f1+wFIPRst2eNzw4DAar0KO4P6zPTPpNYT7kGDtGTogNFbHK/
I6havdfiTBjp6oZheUPGfpD7f1VSn9pM+Zp62PNF+lB32mi6UgabsHRr7MVucSDMZO2uPZ2HxazK
Jua7NHKCrwDGGxVvhUe5cILhl09BHtpP39CgNJ9VwLQHQB9KIOxAnVjwRkaDRi3+EVT444vLZuBT
LSdU+pVzJpmgNOe19Oyrw22a3yCfw4iEZZzQ5kCdz3GeinORKABy7tSqn8l/Y49Ls3DLqEb2sDbv
/WuORRjp8ILjsKCTd7/LRurEge11+X+5FNeRDf4bZTVMoACtKmH4a4E1rCqAdlFfVpCa6LnVquZZ
ngbhG78u3ROZESno+rA3Rru6YZL5GOtYD7c+zR/gByV+62HmWTuQwKAW3aRSPuwkYz0Zyl0HCxea
ItN3EJWRtzqkWQeMrVzbH3U7rtBO1Hn1OCwCEeglz61g239FcibI2e5qOgqKw9epWQXTkeAHHkU8
OgDox2n0lyPjQA0X2Ovy59XJYxJ3yig/nbcjSXVrkd223ZgyhX/r6InyOEookpSA8OXIlAIK6jRT
siFRDg7E+JHx1e9VanomMP1iztpFSP0++U1Xxtc8KHj8nhYGpgm8B5qpAh3Gr/bh5TudW+8eKQ4J
a+U2EhnR/QcvUey+5BZDwYPvztTka6jRFardZm8K22TJ8okGNEAKBxeASfDNjgsZGrkxt+Xduad5
gQxnwcuTBFbMAa2jOnoyc55lu1ZvE6npnDcLxd7SHaIUDUk9I1nhI2Ahqd9vvp2bE+6iCENam192
a1nhIxjfKu4z/1J8GFAl4c+KUl+OFsm0K7RysKMHZUA5uQMbaiIfyQhCwtAdUFQc6ZuWJZrzJ2N0
7kOlFmMwlU8m/6QmSrysbL1bkR7YBMaPEhbVaq+jyBjmXLUB3FENRs1RRqVtmrkcazin/LVw/VVz
/hPc2DJLeL2EG4xczI0VraZPEArrsMrOh0G6TJ+N2SAp6kzlEXcA9BEtEIwieWh7L2AFDGUrtoVC
VKtPV6a+zUYOQyJo0mEyf6TZrTv7JL5csokSxYQuM8PraP1VnzigF88gVvk7Y3DmGc51AXhZSiEw
CBbPXqoskOhRxvP2DgxqcGUcM1mtYXQ0O8zoDSq5bTYgMjoQw64TJumhmMWaqFOyhw6QVrl9bfb7
A4jrTmraPx9wdwObTL0RqqQQbPCg2+5GTQs6waignqwzjYmwLU84Hf0PFWKqpy4q/sR3OYcs3n0v
wRuomsvFiotEDnHFVXTW36vG7jr7mfz7TTQ9J8C+0joZL98HZ9h39NueJwFt7JpKcDvv2szWVX1b
UrHV9CC7XcLBnYXJ7k3ZDByT4jFsEon58Y22UeTnQpE55ZskTeybKdh449IUgvV8DRcIp0Gyyuyh
dWlQAFXR7cSG7C/fK9OnoNNG9dAQkvKeT1ufzWpSg7sc4zBFSkTNaVlZjh2y8uXzmgOCZHPuKW4G
pLcQUJcZdAxTiiMTSmswyZQvlFHae6l+aCX349C3f+mwNXF69oot1ggnUnwo41+2krsqVkNW0AL7
3zVXq1DLeNgyFncivj8P3zehcyekW41BnHwjQqlO8p+UyLF6bhpYWjVNPmPghhEs6dspagBy4MtF
VpjX8Yda0FdaZG+cV9KAsfv5vCwBO9fhILYaq0QaDPs06KAmPueu+Dm0pRVtKmwTB3qh+SQfWwvo
2GCrQUX+hmXYjW+wiIZzcR6f+uKKxmanYdb7Bmuqch5AgPoYXQ2Gb5hTDVZ+13YN4PWTopk24jBm
6aTt/7Fdm1dmiXfE7vwxmoXj5C2tTdKoKfHiYtgQmLqONzPAq5qvX8IlHwDPsUvUthqq1TxnMsYc
Z0e+owQCaId9G1cZg+LpYKFA2G/1UdYa+o93eZW1nSWsyFaLBrR08eq98QK8+xpDy2FsTJj4nHFc
TrpelADsChiL+Nd9rKdZ/O9YtPP6ObHkDzaWw21w8whcfhVMILRKNsOViXiod5sfWaIw9LN1ZWxQ
rDRiMJjQnS7h0mnJTIaLapgc1Cj/9gYRBW5f+t18YgrP5+nWpoDW24GGeWZhPdKXrrb1fhAiv04s
7PaSDWUJzraZtCFI5/XkJxNyIX2DZfEcNfuXJ+/2JhqBdK0OD8o3ISrn+5gi9Y0Go+QRxfFtDi4s
kahj3r5o4MHptr8iQT9EVegQ8v/UZM9kJisGJ45DS4js2lxBOPuCUZU5v7ea2zZoMFT6360/hWl/
kS0mMJQpq/2FPGM3Ue+M6gC8X9Bf5z2WwvkEmeEiAzcPjmAQdjozBvrpcGRshFH3/KutxvrooQLv
EUyI3/S4oH+PHbSbZNYdsjHlrbw+Q5pQFK73tZL17CEmBaUhDRbxCD7WHSVtk22OEdtS19Xi+rG9
u2muS9tI/njgic4fVWvoy6Mn3ZsqcNuUo6IIX5dsywZmg0MCEJavgO+X0wYM7IcGxiMsV29kiVXo
6TH3H6y0fN+yzoEs8fXCWzYurziU54hmxGreMy9mAnAAcvVJsxQu+0vD9n+ca+6UQtxQ1Y4JVGFX
kfTO0mO8ONGg+oV/H7hxxroGUSmxhJasa/JawdIUqiERKWFR/7kah2hAoZELAuGa7G3ZmNUtm/D0
vrqi4WupltJcIfrAcSAPW5lNWiP8ti9Rzduaznq+OaELYFWq+7j7B8WPBFO+Bj3IdqJCH50yNb2o
E6GsFDWbjH9fOJEf0RsNW47onb4Om/ICTHmF8pYh8kTUM2PWbKfrKLwwwWWJIWciq/b/pbPRf/AU
CMi9atPqINpaTp6MOGR4JDmzFE82IaCcI5qjkv5/n15oHKHV2GUJwE7yrV+a8rlhTDI6eEp+94F6
Rd7a1PuTdY7iItBeOjEPXCMl4bLTBR6Ms8P1WQKlB+XAdE23DPlWnveG6sVJTGxdaByKpSVhakWF
s5aSzvTqquAStQIxhsLE/h1IztVcQgrTiiwitPyBHwI3hrL4RaNC5Vt0bXArDEtQwagBpAYg7dtr
FXYgE9wOIECGU+LK807XzwGHtgX/r5kRSaeGQcsWOWT0f7f4tL0n2rDkvJ6Vt82o8sOOfZnQAPw5
W5l9sjbcZMr6f/q5+oEvO42VAD1ScYgsyCrz83VhZZrITXcQsmCMrKx6crG0/fyPDeRWDX+7BVsa
VqWOHN+iXb0zhWIAmCPw9N8vvAYHJllcipNKccuGGgYkfGAws9HcByLcyRd2Z85CRZN6b8KuUE/h
IcWY9it6BTnwznwfyTpjVIe1+BRr5PE4n0mZ/x1pEswvVNDk0SbWZWHkfqgqkQmDLEoc9QUCAblQ
jpDHxdgXpj22RukoY6gLs9nSfYW/g/qkEjkbGbDlu3uM78OfwNSz41fRKW0+9C4q7Wq01qktQ/ke
+u71UinZWs8xWfGbzfRc/OtZ3vqI+EcjybuPgCg6IDjAuvQL2psevjw5vq77g7REncxaWqMU5r9a
G5ju+7T+1UV04UwxQ3F4pIF2bswG+SIYwHc989RMpBzFsGUWbL8vOGYuNJ2Xzq7c/ndvFOuEoWSa
IthkC0gxeuFgibs59/X0ujxs7bJTDf7+g84aT55RMdQve9kqeF/L2TWxv54zSEoJtM5jwD9jyMnT
fbG39iM5H8/3s56we9sl/pwNLt5/WenntOxhh/9xVIBjjAlZpqDUkZr50EfWoO0gWlMv7IkXhTVM
OLoOltsnpgmOx8H+W9F449lK5qRQt76MfiKN8g1WzKaNoXDO4fxkkesJL9ygyDs+0tuU/Jwgc0Be
/k41n27bd5p/YYLIBrmvG5Hx5RVT3Y3jjoyuorrP/tk1qlO6gKOOWvBfHy+IZYTDgbgVdkeSm7QB
sXJX+qCL4e8GJdFr/xSu+bAJf6+UP5FtH0ZzrCv6z8JDrsTouwCvj/95TPJWrqxcelbQd72ZRX1a
ltY2X+qe0kUCrpD++MZOoXM+GhhgUlmswxlShadymsDDqjrVOdV7yuf4l3bUEiR+xu6bOZx1Vg0x
QGodlnSC9Tfmb77+KZEkQ42Xs4V0Pit/QKBxj2xIQzIAqmIeV1+j9V/lZMu8a/0P4BvKKx5BX0FJ
xeIqUlFkD3jts9MuKi410tb9JIJGNfO2+QDg0maWtkWrl44se4d7Gw4HWYSa9gNBQn7Mx0m4zccU
p6Q3iu9KKx45XcHRD1QuE/Q63RDnSY/TLwDTi6bLvAM9b44ryh9D82VdVs/bKUarYHz64pr9GfSf
7y3dnaUkKKca1ZAu9pHg1Wbwr+yb3DYN15xK4kjdzM4JJxWXdVJizF2vxzJHx44yC4NWxD/lsrYs
q45385hdpNqME4+hWj3i+vbC0RDmxwNKeWN0IzmBguwOrE6+OyDcmentASuF3YNjWoNLbMMiwh4W
ydOYOdJbYf7lo3EdQc8EbgAl88wXSY66Czt/OgIjk8c75u0Ig6Xdv3oBnUkio6xvDF83/nQZYNvc
SZImuKzMVOS1g29e15/KEQmTAyJ3qbCXLj+SwgN1RVbNR9n6xmGKbESsPPPr47IoQP1fKWZ9Nl0t
FADC89xj3ZxQKBvvVD48A1LDaXso6sw8g1m7CXo2WJU4IeUZo7QiyCstQJExp0dSqfRzqMp4h5nK
7JiGjRUvn/XZmhIl6MThFJ1SKn+TH66nogtzmjGHuz6iydtk0gTzeK/NIamXdr+beXFfRc/ypjzC
yKSnAzBwcc3im4YeDZ7FOZ+rmwmMBNF/2+JtU+i6cq5D9R1fPLZqUdcP26tT3NKZWozqOTmHDi+h
WP7bAEsdX+FXdWVyLZjhajVaslmvKa1yY5E7PEg7dd7p0PFPrhWE9dDgFso4+WeZu+5NbfcrlPyr
jQsh59GydzuVx+IJr+c5QJNWl/aBUVZDsbqjLjhloyqYiWQfKLEgTx1FAHXmbcxZniahQhtR3rSt
7WPFb5iWubRawVB6BckzNxTkNjHpTsEzWnk2pFI55KWAhw5oJbc24vCpIJz2XhNQrD5pMl1H9HCl
spWnGprU5NHYALKeeWrPlP8pa5Lu3Tv5fYxFitygpak62J0KDcqkqwZQ17FdFkHJszW5ihDYnR1x
6/NydZV0rmB32SjfSHKOwUxKJnMBZrpEXBt7SgRBCivQYB6QZXlwmRymZOZVIPfulWYkQkDL6sun
YR++AH8CWWfYsmEvLb2GXfhJK4li3z0D+BEBYC7aAwy51jtUmmNprXwJw6/kWq+3GuMfQYJEi/+k
lguP7SyR84Sa2vohzt09VJZ6qJm/vWgP5W6Go/w7Iq7nJah2zB2bECxzri7z8tFP/9btNj2ZS20p
61Yjh1k7cD8YS1t3Iy6s8nvkmK8h4rBylMncWYf352k4OS7jl/OqvD9uEEqTkcr6D0KO7sRahZBQ
7O3A0dmII0OntrsXVeJlUKQDMiZQIjrhzKbsvQGY8M9ZaG00XPe/0H1GPUJvDMN4R5bnUjrTeiOK
lGZwu2nPGNr7A077Ox0OyqKUMPsMdaK8RrSzNBTxbjjhauFdFIiPbQAdgroNvp4tNePI7pM/crEo
6WM0i9nSWvoyjCJAA1kTewXBzHIkBCb83vSEbdqOU5dqbWR8UYGrQLVc0B6o4uj0pJv+VJUnmy0k
7cpU0luj9zEBXgaD/bDAPnqsbmlP0r3oV2wRGcpPOyNMK219LwGa7hxs5v0FzdQlsFb7r7phC2st
qpxQMM04yoi5Knh/m6xYLvC/auZxQXujaIGPkfurVpnganOoUMCRo4xqRSID/0EiOGc6mlxZWwqT
dd3GxBjzeubx8cHFpJwVjFG+MKJuaQ5c7R/BtUrq/gaCPSUyjGlx3shjrKLW/elHa6+B6rXSey6O
VXOTS7ozQVO+zogy2WU8jppIqVf8uD4D/8mfYLf/RW/cy+hZTEfGGHkLyzx/ujXpcNwQJV/R5pY2
QALEkXUTFXNbE+l0xA9pUDhopi5krjPdu0nibhrkbvR3hqhTeTRJxG9VVa4ttmrC/qg180O5VujL
0vmBsw7czwc1lSKwGtLtB1KZj/YQCgBh31/KErcZ+8e/QThP0opgFNI1eMzPiSMkmuZPPiBO4EBB
lngH19TgiSIuUwy5J8qrDSUSBDDb4y+q/w0NIRboJzTJELD0U5t+BmVe0uGCbVzicgv5R9ziCZZ0
sFCBC5C2BNHG1knTXpcW1PLCTqbIKZW8qNr5EefocxUE/h+gpoCu63nv0/eveOB3Ufij+3pwum1c
JD9quPr/LJUhsNBpOT+gcvE21n7GKVkJXP4hri0sc1j0Ceswg76svgTwj4iNvhyISbkL5U7Y2DaK
EfwKA6cdKvMwn23Fl/P4MV7cZf02s5Ts8nx5tn+vy6I+7J4Ki6P2ASma1l35myLjUrthGitntx2H
08pzpDdm6FktWjOdVxEWhnKZ3Nu5PLdqmobtoKMv5KjDx1ML46fK+yzAZzEUxF3VXWOc9rLZIB7a
ty5sIWqcRsEh0/9LYESn4bedR75gie3bzBo/aygI+Trs2uFqa5q5dVEPGTnTbNhA6N2O52oYKKhz
z6Rfowr3F6XYFa/DRr0n/ebi0MS6fpFHIPVFWfACpAspWU958nuJLJt7ejEy+pYNiJorFsfADszI
Eu78b4jvyKOK5Qw8oyWUMuA0l0TQeHEF7l93x6ga81QTA594Lg7520r0odbXY2UuaKtDa3wXdJ6s
5Oq7XId7ddghZtlxcRR0fGEVCxPvr5Ws1Q+wP00vs/EeQ/mMnYK79nSRN51LCS9nODA7Zy5E7M1n
L4+3he22EgNmQvIucWFtkmaPcLdIaWMMkidUYfXj4daIq8iudXxBTe8Rc8DkwR+9jzkW/Ewznb00
nJgZzIp7mT1E/QENspci7CGL5Q71Pt7Tab4NDfCyMhjZUfOen+NrTxiodK4SecKSXKVvZ514gH+A
MZ1J3Wpw/NeNmHc51igNmnAynUJZ1SrdbvX5OxHO7md4/IxuUzWovqykqb7oPYBSUtAKKZ98UiMl
7+jOWrtcHaBEYgK6dEdB7JrEAVpkaiznF5J97SIXaV2vRkVOz4R31yDDpNEYx+icvCA9d3GH4QRs
62xkD31DGuJXFi6p1SvYO0wT0gkWvHGewiSlyFPZIiOKu4CxFlMbN+X4ZldTgyT1Vp6156bHVDaV
fA4DkjCWpHgF6qiEVLMdXLUr6v6etdlbB+lq1OCs4uV7LpOrqzP6aXqPG72EzFwxfmKqriIH2+rA
eQCvGaxOgxCHAGltGpEgyJTK7YUby2kgsF7ZiTufJH0T7R2nyeu1v8L6AYiv960VfBIqz8g//FYv
oDMQdqvunX0HbC3h9bBS56Q/86hmPeA7vq+ojbB1pI3hE3/M45cZzofks5wEMVFsqdlVzlE4Kb2j
84EeRZ1g4upORpNSr6a3j6teztTZE3cL4oF967H3lUdC/jOmT7849ug+5R8/k9RqE6v/BDKw5A/5
nsa6++FOiHNpn7q3yTke7pdmv05s8VrkcmZSOtnA0z5C/kOaKFk5BK58m8Hinpkyq+DCFzi4bj36
pr59GR52Adk/fzcj5mzRR4QzS3kwZvJjlA1ud2i768vTLTIkBzXN+WU9ENzE6IhS8J1vhQUwWbxn
ObnFZ85A5kFlDI4nSLciO2PQt2kaLYioSHuLkO20RyUsP9N+HVWnq/hP/GlHwv0lrMT5vj9Gr1eM
O/KdnvKA6eBw/vnBWOwbNVNrVXslqjXxOJPsDW9cmxihaouIfO6HtyxPx7hmtsQj954qaq6g31iL
xfX3YLdT2VkAGTzhxEY52Y+sJc8ING3jYFxMzawWW+ROUqJgbIdslPLWoY0IJeJbenZJo+i6ahBL
QACy7JkCFTffuT3M9GDz6bQuuNyyFwmnAb5cdnMNr4jQ/DqLNPX8JTHza34kCsXop0LUgWOVgJhF
xg8NQ4GPKH3JcYm+zCwvwG3ofYc19ZfJKV7KVAYf9p7cDD/aNK/sKmmEJoiMeY17ShVIQLpnhiHz
KmnovSDIpUlOSps53PpLcOorb95PMD3RBDOoDYOC5BMyJMTtWkl4vB6gQ1CXLzWJGc9K5/gBjQgj
s9DkSowoSvAfVixc6kkMTpX02mNMdPW30bP1MQHNZb7CCUE/rCon48lGtmHrAL3Csu1stw3i/GJe
Li8muQQER7rmbp8Tgrb2J2Ppi3fZa+Z/O8+PtxWCMDWmQSIOzcjkZ3fSPjxRN50OFAzsuxke5lSi
Sg25l7+1zYgUgW0a+ZSHAnhDGyzmz54CjQ03kCAo4UiqztyIOsewuqbNWQIym+zIfWQ56os+1pkW
A2THHGOC8mQq249l1HlrjuBMUB7Ycba8LS4CH5EMPwC5dQo4QFBCVtyr3QYKGSeOMiisP5pOdv8D
IZ4UDVlukVKPP2PwPMVY2LmYW0M3gKEurMUCwFHFdpyyRRqyUjmDcPN7r59UZ0w051OnLGHFAIoq
V76uXS3osqNQOy+7OM2Hs6K6f+vy/05pEo1XYBz77WSapYpWdJd0HyXvGVZAWtjHxCT/vClaFv/i
xBQ7NLdPjdhbhwVYeLAjez+V2vd+mfEuCtBhkcTBK64+7XwAjqWPbhR/mGA7kC/HfEikB3SLTa3D
UZP06AwhDesdpGbnBUWv05eBYI6lnFBBZvRuFytiVBcDAb7w75AHXmPz0/ROnAbIEujZdKGvKYhS
ei92c725khlBat3/XzzMkLUBTzWKrx/mAZ/6E1pbzHbGVDfE5IFl/WKHt6YPP62nZLXyQNZzTQse
l3iYOQPrQk3Q7CcAUgwf26d+6zDcpdqRDPES8baoroaY1UYKkH74pIrZ/Ks35G5pSaEN8l5Zk9Oa
SU1uxXKfO9cHYHPmuXE781Z95Yez9HvUqfMlz7ri/IiaKPEBzUO8GCMovAf+HnKbY83WJKu5+x07
h7pefjC/uolz6rOApPxc3BVvXEWI9+vAfJveCpyPkJCZXqpwCnfNhKC7hA+k5vo4hTz+6vhrM1qz
gWf9qSWmNQx3TP7SrswKCUtJSq3HGfESDXMIA8atePb8H7xgxA9WQWEFJe5Cl1rNyA8CqB82ptv0
HAu35ljDaNlKn2zBuDbY3QW66T8lCRwcaz9Bqr9SsU3ZfBxlxBnrw4T90yb654G3v/oPj/pf5GBg
sIg+e1qRtnJ5MXLT8DljSOq6cyoI6JYDZgy6Vw6zsSa8tG99W+dZ/TWdkjDHYPlEGCi82Oo0mxwS
rZ06bcR7YNTwI8C0dfyl2mSP2TuBBX2/d2Ovy0sxZ9sEvoBniS6xEXVP70bfLwjPQeepnwYaCDkN
ZQTJhJtqDOpUzJbiEzVBBF1Nr+6dghlIowGA/8MLNODBIzh5LcgXSb43wm6Hwfi20HCsvmCl3DQu
WqgvOAdVI1Ll+Gudkpb5STpQ5uws4X6R/kVlRZJxNt0Nf3ng74myHtKTw8gS0GwQvOIQ98uNi5Es
s+s/cIw7FhkfHbv84T+nr2usHNqTXLYjkD4bLk+BVOJ2QK0HmXdgrnDcympioicenIcKMRyRPVET
vPNlrhhl/JGpdmAaJC4H3ycl0jZuJwOINZfQN/xa/qXIN4L4fgAnAfSstJ+OrrvY4O+4LP0cj9gp
or9Vqkfs+np9N+w0t5e5v7u+vEQhyjrJG/vS0Drsf+JvaLX9eyA078CEy4g6OzSXjQ9ES637diEB
8BnApzBv600vyUCTAUYHM5qd84lCCFZLzM3t0hEA9accqKm6vngWxcMDR9bFI2s6SnjnG3w758pz
oCiOOJFudV+NdAEBREaiTCg1V36JnFfEoZMgTwi8xUghXz/9PI/zHBCo2pAlzKpS45pXCimgVjRX
y04x8KphU068a/nwpJy7cJvojpR/mb1zQgxa18hWBT0z1VLD5hDnm0jBaDhcvoLcSV0mTAj9IWJe
ZR/AauN4Wy7mX0Vtm2xHk8s24t0Ev2XsS6AogDwpO2iq+s6y5U6OmeOkfk+RF1Pu8ljHDcblhvri
lT8GxLXTDO31T4rbeJXduXgGxi5o1tvuJPp3G1Im+QlthmnaNmz76Ot8olcSDWYzLkQMi0mv8P4J
18+nSe352Em9f0jYDi1TBMw42y+Fwb44CUJOG+Ok2WZ7/exrXAiIdbU2O6ZkDwzqv1bogzMl/V54
FHuZVC/RkIr40L3HxVzLVmXfOqFgDhl7Vlzw1tAlCTQa4s4j9vcaxD/Opn8wDnxPG9CeDz2QSsau
+J/cMQ4pmrgf1i6ec8Jirbp3A2lmCMMNkhdo4hXmjYO9vmhPI1y6Xsp+bVW3W9f7EJ15J3kQ9qnU
RBFNFBYu2WVw2CcDMkVEkytis6V64Hfdd5zB+v9awvlamHY+p8JH6DhVYPrp1ZE3+V1eNar/MwK+
dN9nqRaWAe9vbrW8WmTSKsT4Th9OYjIHLXZFt19RsTmkdVvz34ZALkjZIHgKnIqxhgLDiUskcFeF
OtzDkIgFKWYYRVonzrMSKN+FgQuBeed/R7ouVOfoqhlGt63vDx7juG3FV2Xpu8XcU2CY1rxZDUqt
vdcZnDTX1QvhcSRhOzD00ys5fXFus08GGho+D7OpyFsVzJjXBsrey2RiU5u4UBVjFns/J+h0uQBt
o8gCD/Z7orguvLNPlKiUoImdCMTgDuDekmINO29X0T7Ah4zVIgst/VsUxRXJDONYTrkRPyaEJ+ZE
BF64q5ZhoefMtHPtUPnbDswKEyGXvbx93D6xBOUz5X9PdPiJLC71LPGVS5kHUwzM8U4lKYYuCp2W
k9RHl3jzo0QXTpzw+VE8i1lc/9WkWiufQczj4puHYWzn1bDSf+U+UgP3pGxqxJxMWW/007vOrreU
vxW5/UZ2vBZU5m+0Q2NXdoA/QD8/06q/0qt786+jYTy8qV9iuhNMXP6PetQL9C+uAXzShq030T70
KPeAlktpWOrIvECJ131hl68InvKOfXm304qiYqUvf8uclHohSbu4ccqWMVsG/HJ/tC4PbnP8dUWU
n+3AEgDnKZUVkBKmMisJ60653PybFPkZmMROHT/T/r5qhePTvBlpzZg7aNR8UFdwcQuUfHsGrRlE
j+E6KF1Dq4+Kq9xD/TtsMXW3lot69LbBInnn+FtOJzzUlflCV89QNRyW/VuPFujEieDF4N4a3UJa
GsC7nMr14dZO9WB9Fbx0cPIgL3sTQ0acgnj4jsMQfBoszCaEQHwICaL2SiS/J8bjURbhCm9JvbXA
+dmhX0m47dyrEWNuUzOQTs5Q1J5nNuCRlK4g3VQSoqxMmow+Cfr7QuilKWwAK4G0h8LAtQ0NEt6l
wwaDT4Qh/T2srDiYuBTxt+/8ntE+PVBeUo3UBERz5ZRFlnEPNpV/3Bb1pZbsEGCOe8sWyLx5HSWh
wP4FVUOHiq16f+JtQp1ruTNGQEzpthsTusdwzq5gBsQVD+efH3JQRHj7D/ydotux1fwgR0cKS6Xq
UuLh8skkLzOIKI5k70YT2S894bPgVWZLOaoSQndzYdF6oGtNIh8grDGpL257VCs96yFZYnb6nK2K
FCRtyplFfZe4195Lt4c/W+oPKA3SEco08LivKSSv154VQp2MlESi/RjZNuRcHfD82DHOzw8fYnlS
e5qkNxKunKb/o2myYbPC/KDtTOcJBJOM6VV1HqyVY/hBRRHFQQa9mdpOqPS/ImD63xRdtpiCuOk4
KynTqL3sXodjLL+0mffbYumVAi3AiWVNzuvm6bMpAg+hoMAwnxxmF2KBwIOF4L9z3uY5364HIDcm
t5ojpMnWXEqjb/XWZCB82c8UkZkSoypgAEzbZjmaL8bCWJZl+OnsaEDNIfL3BFrhAOw9lyt8nPed
eUb3mO7FijMgt32cAfrspq/deNXOeDdTw9BJqQW/NHVeqg9GuuCOj6PXN2+c2kGXWaQ1Tt4l+N2l
CiVc9Wec1e7PuRVuR4R3sfR5Nqk7tVOTkUuZFsMMVL9Qn8SVYq7F8ymQX/+9zx72bYCKwV3UtMSu
gpDvzZuDd1tYOek+hGSM5c1vsWaVyu1YqongU+qYkqe45WE5C6QU2lw1M5FM48xulP3NIkQoEWlc
jyl6MWYQ13cmZkcxZZ1vQvP0rYEmjxX5FmOnKP5RrCqTE4JRc97sK8aTTkGOVSc0iZpn6nHZ8nEa
2JiSrB3jZPzxgZRg2JNY/OiDi8w4DKVmZEYC0Cr2D6kncOpoQ92/dHOjNi7RioRB5EUXZgp/u6M4
LJ4tSvXYJDQqQqpIrfTqHCnQmCGiJDHC6Mhv2XdEZ7CmH2FJ7HfUTXvvSgzrjT4I009WfGXf6MXl
plagTKCYCj/EqqXPDQVQfruFp72OvEawAp3xG7EGOo6dCyZ/JaXQCVL8IkIz3zY/ceqH8RAxsSBM
S2mYHa+o4WuiznK+qLyk8jBJk304bE8jZyYvtsOs6IDTTnIs+9PGjLcbVWcH8HGpjwpUMwqTj/Jr
bpXrGmlZlqtzSWjgar7FaVYC0Ht1DDkLjPciO4FSIZsSq6tBThNASIkXCRm0R2vQZ5XBUOfszift
3l4LOfeQU43FaDNlNVtR1p5TMWw7CSE9TViU3DofftTKoeYxJwGF025EMYerkpj0S6hj5VnDh/s6
bpSBaq4iT9kzWK0Zb05/AYN/HZrmW2U4/0hEtMKl9WIHc3TzZ8o0pMQ+8GqXebeUd0rHixAQwWg2
1FtK+bd2lRQvxz2AzIWulIFPqQMlWGczso2P1sv/+/BD4eakaW1tBLPgoOfq/fIKQU5u1AeQvTtt
s/+GbVkqL3dK+APDbcY/KD32vJ7byP/Wuw7n0qd9TECJU95DeRFDRH//BYu4GfYUoojRYgO3N9Hp
PqCep5VX/Fnp/wwtYY47lYTzncjJ7pXWQX/cjOVVQQxUnnk+dABhboTl2w/atjAIL/dJ8O403b7/
RfRcKYrh94VykhlnG0/Sk0TlWprJ/+yusX8vZ5ugcEmvBOoKsrzEmkf/QACmUPcMKN0hncRkiRX5
FzgelbFkaNP69z9iuZcDlLZwAh9E58XPD54eAfXQuI6skzUWoOC8pWhdkF5VjU2Ms8CZVq2T43Qq
9EsbYS6h0WX6+ytx13DmsM18O+dkIh5MVr7wBry8B6PLjlDAfIj9ivwvJl42M7hJIq1TB4XOw9SX
CMynLuEF2GwwTSMAuReyDUFCVYdBMNnbJoT+tzPbvzIJ48jSnHVcLhqp3iaCdau9nMNrJYxoJQzp
M0bI9zMhr6ZN1NvlToZzz0LYKZElc+b+8xVwUzfCDC35ruURE2bAOHUU7iKy3tyJtxZePk87byn+
s4TxoOxgLC5mxYQ0soaqP/TpjPAU1tdeHJV98rYkIn+X/7vWG7ycqk++g6Yobc0OPxr1Zcgtc+VR
hJ++mrrJkX6ObmFjO8BpWicItWiLGRu2T31dvWUICpbzwN7qWj7NH24jn+ZGajpTGkb0nhGHkOds
zk5cpQ5JeOZVg4WN7DSlVuldclQHgSItajF4/szBvNp2GczCBRDr0qZ3+LZPKMBaAuiczCD37iio
rIIq7mnPSk5B/mA0BU6yEWveBZTQRdx1aDQSNFn4BFqkYnw21lEvJZySg/OVq1tEd6W6VRvrZhim
jhutcKxHhC4zxguqj9H6NwD027cYg6f/AtINV/7odNyMVgtzPnJNsi2gt6AAwieX412K8kx0QK5r
CI4M/7rIWd2DMU8L/RAx2m82eAG8/2EroZD/UVlVywIzQ0P/vp680OAUDROECbWY/Mixy8iRe+dy
b774qhtZyJYbFiFhI6652AFpQlcCczfvQHglks+YzHlHEkK3CzLKZ9ia1Cn8DtvsZiRj04HuvaEQ
pRtYtTv7eZXa3XvLu+j8G1uebG9tj93qsYk/0VhigEJDcuBFpo2njTFHF34Mw6OgNOBIkeU4DVdd
rrv2ZR9HwuyMe+GmPT19GMmKVMUO1KFm6CFhOyF/kvnOVfl5P6psIf7nwETA9V5RfoWk7nI4wORu
NN50l+ZMPpu8aBWKGtdd2uEpg31CIBgQNv7LsgZq4MOHljUYQsHvxahvYUfTvIrydC/qRTaQd2xV
xxcXMr145IJ7nb4F8wRix0ndmlgzk5lzaefi7YI6p5zaXJHUwhxmiyA7MXx/F9bKPDvRahRUMWs9
z1tkldwBy28dU7qlq07KkA3AQKa0+MEzmBnlxLmBJ0Bugm7HaLNRJst9Gu/ymrifllRjwRyXTCA3
KrWBbantOEVyn9teUQ1hID6DsJqBRg/1gW9e0dpNNIwRiHXpfn3ppCBTQcgK9wfGG8HZihoDFld9
ilUND8gBHTpbvqrlQMN/CvVx8nerthbgksia/F6kqDMI5NM4nILOYMVXenokQwxhHJpRFeIN1FQx
70Fh24Y0GAeAnJGhZUE4zzOZ5Oi+qgzphJZaPuRPgSnih4vIcxMBzio3LgHHDvIdo0zqW9qZRa7K
ESkmTcKhhJ4sJkXy6+0f/8lRh3uIuu+DIuye6YLFixHpPnZVObRq5ApTqg8SZlR2B1ZHB/dvo6nj
0QKLd7Ghlk0zucBPMDnKpEqyb2TTsaG4YB2D/jS4oShiqJQW5tIPQfAnSrR8Tk+2bYZnxhQUAMh9
ICHv4I5k4USdy9NOePwlcUZOJqOypd9FCbOlG+N2OjYVU6d03wRiYZiBeePd1UCYLeKtXfDwSlOd
blTZ5eyvFIxgctnURtTQHlwSr/yBLOrkRrSlDJRvJkxu3p0ZA1FInRvdNRS6xQzzedXrgHHuLYOW
IbH4vBxvozBbECA3B9YVP5Fjr/Z0J8fwFibIbgeJ7RZMj1RigROAokhaHNfoSpx2qYOIR/dKX39H
0Byz98LU36HJ33jrGETefOuUF1Z2pcos0gQyAUnFqMkdp7Q7xzUVsrohg8G4SKMWSykvKjDU1/sm
TowobEPaZ8352TuJruluYgRAjfo+/cZj9gP9PhAlYwD635W1C5H/pgewWfV3qa/zQu1gzNkBqKqd
NNoe0BENRbSwU7VIt+OYEFShuueoBTcmD2b9Y9v8wvO+/8zmtBUanf985OgYXprCZ8HBIl3rBLri
/3EugcRM6X0vtqY5Y69tt/6lbDClTEggo0Q2D9g2S3wzafk5NVbGT4fQXlklFnejqtT8em79j6Nz
Uq1qx4VjYR9GEMHqL0/pp/VqdBruNpI7Qb5lel3TcNaeKWayV8POugKQHvRrpGgcsK4pFvJMlGqJ
AihjDrjkKxs6mdpf8dgZGFX8oT1gPI93T9HuxD2fAoBccWLCFqJJr6oeaEP6PZhnaYldrPEnuHA5
8TtkjKY3VYpWwlOKALqt0yq4RgC1RhsOkeB8d5wfOIsqmZSIuhFOsSkyyGk8IKc07o+acTz5u7t4
j1WWm6G0WnPLu9FBtQdfyVq3Qga5SvocS3rJZVYUrGN5zFQ9FB3ATsPtKgF7DtzguJ85dx0uDs3l
l5AgCN6tzXTTME9VuAIQUoLJbKn/Ct3nbGdL3LXaC3tQTwow089deCWHlvZDV/ZhurI1u6ugIV3X
/tcdbJ4/BOQ1RXPAE4UGgi+lJzgByJqj9vhZoJ/aDGbvaMf0IT7CFEHJKkhg3lULBX16yshRSP/1
nbRRIa/W6uOlIS+jQ2JZCGY90OPiqH8Mx77pWbdfgr5NhQXm4+te07lKvYdlnBR7aSIun4Y0IPsZ
+pH5BNVbW6cOGfOmTl3MRppR1UmCfHd3ZjkskssVnf804FBmeoMopd7SzoYCGEay742F7iWgZQ+7
4MFEiNxCHQBegt7BMMIokAsLs8E+yMnuIgBdyuWyqq4zUNJ1msLNexl7dalabq5LKTKD6Yvoudrv
6WkNJ0k10QWKUzvR2PgkSeGqQo+0FZ6aWkE4ISNQoYTGPg8c91o+5WvznPVaza/VIgSeUY7LTMZJ
raJ4Bb3X2akss1EB4ogqXWKYSzxBpOKOddZYrfGz29p/EX2wZ98RPCFbi7cGCjRfQ5K11q/y+yLs
69q65Qv9t07umTXDzlteInzwDUvTnJv2pcD6e9cre9rcefc50DwukRiIKNpL7PTfvQJraSIygTHo
sqhJkoGQB+0K0q9dyNxL7KLgzrpIKzZqDNIG/pwoJ49PytJyJjf2fFsYbKdlgTsL/g7Y8el/Tmxa
PZN3tHqYnX14ZboG3Vl56d/QMoCslPXs0K8TgqXI+SbipcUMvwLvQWYhky21HvDRZvdIvvO4j1AN
iO4ylr4AGE/OUybwy4A7lpHm3RWJYAhoQvE1Xo1WfAL4pqQbHd2m7KLBU5ZB1wtKo4fhD4Czk2aM
2WTCFknw36oQ1NyEBb3AD+jfJJukBJuitUoDichloCPQcbRqG56TX/Emvm4g6wwE/tWBnqaT7NQh
IckexwLddXoY5bkOXQUHyHWL/K/+jOcWHX/6mBt8zJS14fvsJEhpf0TbELsFdB3pMVqVo+dJcs7s
eWc1I5ZI5XjrVYuOUB8K26oB1a3fwwpQGcmcKDvjIEHd6bd9Ura0tJmN427azqeCPLixabET1613
Up8NuH/Xa454H+bW3B72rtujX8D/GhzqPqqGd8ORn//dsuGOz9Hn1Sk/BMIL22aq8ruKGdCb4Qcx
bVjF9krgrHZFWSX1KR01HmI19fJByZU8YGDbxiUjuU4Daezzx2vrvDPWxUwxflZCtzTtkvXWbmUV
LVS/KCmAUu1nWRDrdI5+B80jl/y4l5+XPD5+Kkqogmq1EH9q6aPHmHJrlnWgfejVQP3YpY4yQgJC
dyBDC1wiWLEJBvBHyVBQZwtNlEzaULCdk2wFQz1kwhwOAdVFKNvISH449jX1C4ry+t0PiB7aNQ6x
Z0KCRhPnJSsAIEuD1HXiKbsNFaQJ4Onq0U7SNx6VEFTfqecNd6fl5ZOtjiE4GH99RjF6XyrFE5x+
HNjtcxkDbixOX/P7PO1Zkqic4VoGk/GOiP75KeVp0nd21cHde9r5TqCDXLvWhI/o3fO49VuZI8+K
n+az19uJAJ0LkKT9GCCV2RYN82rHIQayxa1RzA711icqtUORjrwkna4f/yhDztDqz7YhaHGpBbwZ
trmC1S9OWS0Y+/poSAmC0i3F9DJtkR+FfQotzNSTJn5Qet622idi8Kz45tu3KajK9xbFFJSoSnDe
MpvZR+ByitYKb69xYQGnnSd1VdtuJRRK4jGuqtaRcIJwkp3ig9StQtOjf8DXFzY5A8rBV6WWnPbw
QtDCi4TyDcpvtUno9Jf9LEYEzHbfCGzPYjczs+n8+z47yxOP33tyl1ukAm1rmIbMS52XutM2Hi0t
tCfzXBmnuG6H31Pev+qmppOv4J9soyFzYG7HYzUmP8HAnSNTbBACVCRg0sbIk53AG8FLVGH0BBtS
Wv+7zyrri2AgBXfjZhACjdFmUmXhZesY2JYNAAMv2UllS9G6ZJPl39KVBQTzdcHVKMcYDTa+Zlrv
U1ImhVgRcQhcZGAiCu0HmZQ4FYa3CS0ejjmuLMiMz0KHr1swYLzCgae5m1b/4VJbMJgdqjXpbRix
9w2u3F6pVM8sP8EVon5tPI1m8pXJ4PrDI5ij2T2FiY5KbPkWxqR51kwYPsSokt3rdDpJ4KylElgi
e8I+ks7TVgP92n1n8btWM1yOSNFl7VA3n/a81ieBazuevYU8pi+u0uogQYPhmajG4diYLIzvqW6b
X9Lx22q/lBcrvcH7+GlLE2q4MXzuowlRFG3pHVKb1CLQeKy2b/tDPwAXf6uetHFAHqkwLwirQtBm
rDaGPXrQb2xXDjzD3w2a0jo3oi/Ok9jWeznJuGVqcHRCl8uezxLWb79kAmVaY63NLla31krCYZZn
TswZtJCaMfsR2lg75Sl1YBiTsuahYLLrFafBQRr3MMVsg9mtD3JQubDGpBPdcIlHzvfKa8iD4Sxf
epvkEHbfnI5df/vGvSGecKj2KdZ33uxDgozuM4i8JLWh8PUMVRvp0G+LvCe39qbOagixUKKKURT8
w5uG5E9i5AEGpx5s8pmhJBIhs0ZTPiWZv3XwlTn8SzBM/Q+/JosLiYwrMqbW/wgJdbNvBosnVK89
RaokLq0lk1Vizf5C2PMhr3EypnezY+Ff18GoyGt10EokcQlfurUF1O/QCjJMqJ5pDhChKlw38nrG
OmF4B69y8SRseMLvNzLwaoViIACRjqYpF/Le1dffbB7IuTOskd/uUjphKWQEMqBoCPWqQ6p+prbC
kZA5KZ2+DiltgDKWBrznm6VvT9UsGoPdlDszlqWpTksqYRKvv90DhSpc6oKuol1ElDiq/dT7kEy3
8jBvkCCnX1iMjrPzeYYkbgtjx3W0K4RAD3AXGE7zBK/0t0ySD7EzH/1Sq5d9sLLqyMyLGXWPCo/H
4n0A0D5zR+IY90X+ASnoPmBuF5uBKXSnv1yT/URlNDAXtgOJU3r68+jxbJzdNV+t/NfnLkZq/6ZQ
2Iie29IY/v8mvPoenGc6o5AIBZ3JxD3xcS0rEYBgQUhlUN4z6U271SrZRKWRFhDodX/hVIJWc7RF
yvJ/NTsV3HQgFsO9Neqp8oktY674IfB6t1TKKbPNENnVYdET1gUIb36LtjIox5T1tZ2hXgo3KBmK
Kb41Q8jXqmLhx8tQMuLyE/4Wn4IUxLT11QJiFVXpd9ZydDX7WcmJziw9iIpeiyVPLLr3fcjs1aFz
I90sEHO2IBimZzpKA3WacpEB7nC0EcSP790CVagYL4VCvIGUkA8VfMjDtADWr7bci7zqEM9M163x
aNDZ8f8eKwRgQY8y9Rff8yurYHIbOkff0GAvdbsgGPQ5h3ALNCNtoUcAytfCNapIKU4cMn28h9lX
lNT/c1XTn6AHWkFnlTyuG4ovk4f0UvaCbK1dizTMsAnWDJLrz5Y66jKWHtx91tYZ4Hb/CFvDyZLu
RBt/yQjxLDqoso+GLFoshaRFayhCUGr75ID8N+7eJkV5WOWNs8rOVk4cDroK0EUv/eDj/u8yoIFR
RkHAphR77exi7ie6mxbtejkdie5OG2eLYEWC+zUwpOFRILP3ezhV5nQbfMMt/pwqZfls3muXdiHM
ldrXqrTdV0M1MOnpL7PunI4blU54eR1A11VprK1zVOfi+FIEJktowLPXX6EL9IanahE8v56MfQvH
lQjb7isluMq2EHl/fXfXui2wJd7mgcUl9/H5HovSf5LiayTUDFU8Xz4h2m+toSCP9czA+ev/K6TL
dxw1SYkdoq0za1PHlQXbsKib2MAw7tVK8HCQMie0FaS0FfEEZHvxPegYHdN0auDh5PHomSZX7rWa
5XgolFUQtOqkOyYdCKPSi/t76OcaItQ4LYhTkBElLa9sDx6hhe6l5VrMO5AgbZIB8YuyI7Ojg0wr
vZt7N5FLsJCOlo+VC9Agm6aFfzNzsGT0eFn5pQGMVPR2su8y2T0DeGCTds05+RGZU0ADNRDuhhFj
aH0Vi7GRfx8VcxRYExZapam7NyU0RMWmdjF+h5zSi7yKyzpckhsxPfw4pAlZMA01rX+axajWQI13
ljOOJw6R3I3TVs80lnsMA9UjXHwc2QKNkNiBd3y/BaB/A0/u9wn8MNhalVkOkgTPY0zgdBvMyXjA
fMkL96cUqvX4vxTH1CacbTi5YGgvYqdy1G4QeHKGVBcCjG62YyHfqd+2pdSoM0DzLrt0CyT5AFEt
xjozsUHEEUcpgW4yi3rRU9zlV9RHfQF25OcDHUeAdNfddnx61HI8bAfSCClOJM+KR9Q+adACtRBl
n280FSPxMZW1PsDvOwmwJiYce/TO+HW/u9HuVnpbFZzN5gXSnEmtKZ9wb7k4eWLbcifUrPPVCByW
gHfmPf6nxAloold4cr/Afcat1IdokQKDdYxmsCH4J5K5o3yQeMmfx8Z3Zz/wkZK9HVOhd4JrltIU
aumitgircAGjVOIeMlicztPNVgaLP6u74IbzE3FMJ7hs02CPjrMyvAszg/Lfhbz5TdpeWSLf3/H8
0SBRk5P8hm65RsZfncZsygVg8mtk7EVcMZWZWvSJlx0MWy1DBcJCTSCY9+j/qk7IYgu3GW5sG+OY
Ye7gMUAWu88PmoaODj8R9zYRMqanSZx2ATbbcEnlrw56cubawqd21E6U2mONjDvaOiomR5DmVU+/
QDuQOn55m+SFYN2smYR+jyb+UWuuilhwQ6gN09BWT9KejHvGpRDs/dOET1J1Zbrqa6JSEEiPBTeL
yWA8cPnKg4IQCnqADo1wojmtu40mH3N/86mJduczhXELwetu4ykrG+Qxcl4fDu7qm8jk2hsgVeX4
wZRmbLrMy7a53EzTKUyl4S67nRhTWjSmAx3GROVoCqmODPsIsXTV06sJ2LCiZP/eWFUkqOG7lX+N
+7i8hSeyu2zHE3WLroq5ub0O1cjWZU9s9IDbs977EgufrJPbm7kaDj5Ep6BAuFWUjC3qpmp6WyPa
WItM19AmE/eUg0WkWWoVUl7SMbh2yDZ4fmUGupdZI6FUoyQoM5ZSKLYwp3ri/7hGFpOQQcG5UI7X
Ovl+596jFG0p08J5fMA0bCPMRGm1FBjBQaMwtu5HfXAdndY2S/3DjP3NnfTHMKHDx+RJ4bSvbd57
xj+l0QNk3RocY5LZy9vOyMeIpHKNF4yl2A4ULCu3fRqxXqNrLSigDL8ej4EVdA0+nz4oPQQ5TRsc
5N+OvV9Xjq+ni80G2JAostGEWuDPDWUnVxF9T+FrqpXmL8blCZYiimpVVOY8EptnyLi4ercy4apn
e76kkC68Zz5chnnqyGzqZI2rOEhFR+dHIBq8cfpDJmIdASoOyJ+vUMiP6VjB8YIaW4feYfrKnypX
iFXAOl4vA6YROBNRniFeeiGobCbd6d+DicpLrDtHT+yiIRQuyrQhzfN57pFreV/NhjVMvQjy8LWS
7K3a+L6W68CipyMYi6k+D8gGt+TAGz01qFswZu0ksPoSBxrjMDq49F8EZBY7BDWWSJUhSWrQJCkS
jTB7qY0bwda6A/E8buIFuG1RpsWJUY5AaLFKmb5z22pvqVzK4M6ik3XOsvOyT90OazCejrhtjnkN
VypMxvUqkq+8znKmOg3x6y1TBXe5DwCh7EKg8h3//3/saDdcDz7eV2WoH1FhjuCdH/lYpdmbCRc7
S4Uxb1ub7j+s6uOqzEmuaOjmM7Ir8FY62hezOrK5lN3MdRxviAM6aDZNt2+u+hGxPEriryyezrdT
ww7eFX9Sql6cQ0VEuaNKrR7Lf4l4XbJXEdBdTCcOKRST6k81TB36odeQkJLJc9v5hAfJFZWpogRe
lhPgOJjYIMqh8KryOMzU9Ihb14mK7nOwWn0zvMLFN7nrqh44G97xJE4uR8p8gs3953CDlNx6JzUx
38EjlEb/uh4U9s+fGTAHh+JPtWnuc4IeZll+g0GCU/4578/BDmAfceMfa224eKmLvhUR4XYEo1ch
Qg+3sq9FoZeobv2wjYn6DFr8F/RiNiLd0tJBWW/YEuo1Kp8DxwGsP1y06Q8GvwVv0TND5HSVdfT+
eaj3LCzpSiSx1UkcqHOvBYPVyVZdlF5mlvJb8eL3B+8/C7eMXxnGpJAWk/KqJEC4Xj1yCbaWBrJ+
6z5TTIA8DIosWzk0clOY4VWLqMhXPrjiBloTjxdR5YJtelqBnrR/FXziuiTMX/+pDpwliI6FJOml
glS9zWAqa+FVyOe8rmiFRXQ8jbadOS0bxyZQHJECQXLSEZFenvwJrqozqVqzUnm1ClrVJw49dcUg
cJ/HLuxHTdfdIQtta1+Ei2Ufo7zInvYwkWOW57V1Im9cOlYgnLnnlr7QJ99yQzEqKt/zC9my/m11
Kute/SpZLeEPw++GKdtuSc0M294/0AmHWBZJrK1y5B33pb/yzKuAIvfOVikmBo0v/OP4ZAbuohb1
RW37Dy3FEkQWvpm5uuJqjRH6Crwg9ylb9ApXpiGMnyEDXJZWR5cypA3KjUue7xKJhvJnVoKiaKo3
nFlUP3KGevM+fWsrZur06FieQYYaz7RdhWOC+vE6CvJbDX+TGuGvPMtwEWAzS7FWvcTkFLTfUQbl
bVKUgeAD/77jQYymTMzsKMlRsKL6IxE08VEDHvc3o1Tt7WOpBlxlt7kaCixEQYVshzffhuW+hTXX
fjDFhaRUIiX4wgr8CnoYEY4rSGdON/PAdENqb08z6JqRfFChEhgoZ7gy6Q39Jn1joMrlGRlYb7Pw
fxKAMczCbTv8EleLaBKvCFrdSQak6xctOBmH6yp/DK6D13FETFC1Jpy2kHFUwmbsZVsDIfr3E7PB
KhN+nTOhZ7sS/a6QMBupP5kBu4RAIaqIpTg2pTRNbRXIcYkwrR1bTMmNUXyyVrL7x1mM1IMGXTAF
yhJQsU4ADA7NKvkU9ZGKpLXMTp4SljyIy2PUofaipAR7MQ2KW0CTHMnCkdeAwRRj65KmSLMI85IT
wtpfezzIfkPzt5c8ii9z8WuMN4LMovhBMIK6VaT16F+zlU/ntf6bh5Gh0LRVaEFXF3+RxMh/TygZ
3f4nEJyPWmumnh/QgLppFLb7zA8XjrU2AePR6WCJ81MdUT0Dvo0sS+Md+L5F3MsUgbSaczemWRuQ
2LLf73xXsbH+s7vUmDdbpn/Xg5UARhJA0O1Bog8XfjUOgvvzi8vLPGbnm/YVoLRO7a0oAcpUsAqh
qaC7IVaqpPYMQ5oOyKUkXC6sT8m/aQP1/JT6A1bwRv1aoW7lwfiKyy/iDBpEQwFkqHWrpBtjH52Q
IQ66z9S9MS/I8ZxLou0Y/7k66KjjVBOz6KGcErbpPFoJubqXZstZs/pPXD5cqtKm+Uf6KHse3unq
XRi0DQwb88QGBe9nrBEOh1f4d8HK0y4HrPDNsApvtCIVC2mE2xf6W52/y/DWrevbWzt9zNURiP8C
/JACL546DmAObhYzTLVrqsCnRk8NEYYOE0w9DPPIHtxYwlWv5lxrxckE2vtopj0+qo74IvCF5f2l
/qQwrlqpyTcW+uWJc+elOIveUd7+gErfuJ+LdcRqA4UoaMXyf1Sb3OuFAmNw+CB0QxENy+8nYM22
RA34whfudmTKDcwY+fjWJk1l8YvUlV3njlp4Iy1MnLowBQgXYZmszXVmREQ//W/poDLpwBZ7dqHM
V6iD3CZ+Io1gq0nhWP+S6260qZzjrhX8SIDLZDDBbEztA3Ck11O9WWVbbafZ2bSi5vzfW4HqQosQ
kDx6ZD0YxsfFbmNRcFBHK0hzgZz8G/0L+P8owHT0/xnGcQdXm0XbprNRiJnpY+IKdCdreyYzYinc
Rx8eG2aoyC4wPq17NwrKwPydLl37BuIQgEkayKw+IhSUoLpkHDo46iA517bkZH9M8bM1/TN9QwwQ
2Wgi3WCRKbPmTMZ0GT4qJ+y2GDZsId2Ee7A1XjYrilAd5t/qQuhN7RWu8EXau2azblKzyzCDYNfM
AQDUn5LddjKSb/IBNSAszWbBbFiAm3v8G1WSUUyw+TTR4iTQ3AtUm3iZy4M6///iKHYUZaVV4Tre
eboS+gzdieyEZ6nHc5njjcdGr9jnFX+TBFJh1jcU1TAhIFgRc+aOrSIw54/p2qZdOR4v1Vc/BgDL
y7e3ycEdAmU9AJTsbGG7L0OZiiS8n+a3zLkwehyClMYaavTrKGAZKk5VzVk0Qo2SE8t7pDq0uzc5
YxLSLGzDwwFbmzL9bRKCQ4ALmNZH5i8jR5E/rxRDFHd+qggDH7JfH54YQrJUizJv7b2jx7d+bpdE
SkB8IRvnKZVAEjRwrT7jCljrIsNfINhYFMzJX7RPhdJcplP/EATBUca6c1XjXBRwoOz+pC848aUe
IbsFRMPA80tWYMwQCQv6I4H8uzzw55LpT7HrhJ78bJvcpBKOa9pyP2+K89oUbbEIzybF1iytbBjO
R2b5lyumYlxjXevJYLd26tdIYwuX7oy8iM4TE7KIyk+LnokKmud0Fj47QKwlv+kZWQcabltub9Er
uTAn52Dj9Kyznbj8czXbH1RgM7wvlTefoOeG1dYaC7a7OLJb/wIgbIlHDSKY6cbYAlBIY7oqj8Fd
7oCd+EH9lDQP6XLyX4ZIPS+SM4ApiVk2g+CkPCAPvnHs95yzMpPul4OTaUFoDYQwd9nnOMgx4ZmI
1gUy0FiDAi1+AkVA5LKdjPZz4HqDXrmpsBbpggCdMmQHMvmmJfOdLaVrk+qgS+IWjR/tAN9P4O4m
kSeY0x5WRiKzuSjfxLAwjuHHr6pnuNnqVXwRv9hSrk8vONc7x+zgcZwT/EFhJe3QbrT8cYQgjokv
HfY+TdOKP3vy96BDbmdxfruj/Y+U2wabkfVA2c80Leru+3k7XlBcsEIrORTKBYQRSGCq94Y5dETk
05t8ydsG2ysQJg0jXZsz0omSAnWYj1pzCxRuQ0A3cJLRyZAP/FTeSpUnO8l4gLfn0dlIN2Y+hu20
l6PZAJos3y8ZF8/mFcNraGAQzQpyjVUfhFu9VVO2jboKP0bYWh+PFsOhUTlc12xm1fRUkvGpzGWL
xnHV7kSyotOhvHL7KYAMtsvAbYOH4eV6QYEX2Hnu6g+SVLfoHAeit43bXZISn3PHCWBD21jRc5kM
4uD3X84sHw/A6Qxmja/OJa4kjxHX+Lpkq7oWZGJLN9mmrhHalmxBzTH9kr6WdDNjCfu9SEv6bdtD
U0A35bg+ERJimlBPfUUy7kC0Oepf9aiMeS57MVSBqRghdYGNYVI28jYae6UeJ11tpH1wJDvXc/ox
JuD1AYR7t+LUe3t4i8IiiR3p/ViirroePAgxIGkUC2TN7qFtrYYsdyX1DXOfPUaio2WyeN4gWCBP
th2nPCDTkqUki+QIEL5GUtWhrZemBpfAWmr1Z8EsMoTC/I3hxpamcPnYuoSnHjBNfj6F1gD+nidU
d90eAlFOyisBHBSYBIRL7jCNfgXEXPhKLaY5lnDweS8d4tNSJB6wcTgcN0OAb/UA6LZiemYg5zyL
LxqDGsGMGHOUlVRcTtc64QHdoXubDjz942qQavPoOel/cWw0i41nuvrXJcCm9ZHP/JdzBpezTUL+
1482FOqTYbA9A7vHkE4anXOLScDJ4shtaZjgGwFK8YnZ6qElzFH7E+0deZDFxiw63dWKEIkTwmVr
FLOA5X+fJ7xbs8lyDQPd86QkScqToNjSnXSxLrzmIil0n56e92CXtDqhmfKb5PgVizDT2s9ST9KH
QCI4DjGN6lTFi6g1uqUDhOsXRW4ZV5UB5ZkR8au7bAhnV3KlAOtBEutKhFZ/j/YmQf5i69VkIW39
sZ8Qg2o9wYGJPaIej/JtIJRGoh1KRFBETKNGy2qLF6DOdmXsiK9toNSz0mgrDO4OpBiaCcOED1ZE
O6LEnEtxLt/cYcejfxc2Xwtpvdw46NB639r8DFwlovWtWd6yisHA/kuCZgTIMl7SCioQ2GDfi71K
UzI1FI68qR6A6CU7RIjPEqMKMXa4bi51S96sJdS0SAuQBJVaMJOFXP/Y4jXFI2v2Gy3EInggRKfO
0/PQmCeEWsIgvLt/dDYo34hWNIqLx55iqqhBJkF3/PhMxjpUg8XYRcxP6FSwvq24Q/mvkd/XvzY2
4Q9JmpMUtdv/EMPeRqDJieiQJBhe3Idzy5aOUnAu1zbmg+8JDaNrxHoB4XWt6kqaGKIsRoboYIH9
+lFRx5KHOUoFeT9sXF2g6E2GFbL7JkLyeM7Icm+CzIlXcmNNg+b4RDvVfRkBLfRW7fVZdc952G8g
O6QZ09CmZzeFyxSsogAQAzHO3Xs3Gzuli0nEE+0lCGRf3JeVqk4stok4ucwC99NEnQNFZR0eQYry
hbNs2H0mBDE1jT4mlz00Ab+t1hmRXqmrFHw2pDJNOw+IWNlZM/8FJn7Hd8vSzmgLog5mdpNuuJuM
Xn7KGgDrWiVQ59vmpiAcHWad5I90vVRARaheBfiVrpFYkhr/8unEJTzpmrIsJsuar6Puw+GAgKM/
dGpxmEe41GLIl8mkrLGToNxuBDgOdWH3Ux5mm/SB6VE2K6aEfXxBaZjeQzmJJ40kK1nZei0dJNfG
kHlopNECLEgl4CyhsqnMU2RLPcwC0duRzHkzZExy8wGRISxy8ep7tVGRNTNgQXuAMEh7P/UNhtCo
0otr1gLXyQNPhwJfm4dmKAUmcBgfEjIQRNf+EFAIpSw/BNd0aJO+E0Seljx+AlR9GEi3BAXgG33D
pnTbry4Jfj5YaZdufv5G6sI1V5k03xH4/SzlInvXF1YoVzW6R77XqgEshVvgcj93PCpKSLrytNDE
da1FEcUGsiwXj/cTtU6/vCKSVKXG7yCfFlk2aOrC/6q8gc4IS/L7UTTjlDjLhpi2RJk9IzVlaHed
0AYVGczhCamoUWPowmdjMKEJlu1ZyX/epnOM4i1t2apR5FLeoAk/sATuzX8JASXI5EClGoYALczL
hv7Q47PWcGyNiJAynGcJB4oP0UDAwyQwc9m0/Q66GWG8PpBWLrdjNkVXbH1cuFyQcaO52VzmCVhh
L5Ek6l9fH7h/r7zEla2dLRhflRUwBljjY5ouixUqCeo0rgxUqlCNOoDTdh7b28cz2QTz1kK7+IEb
dcI746YiEWHTHQnEr+lLAjPSQZJcRKZKcxPxqa19H+79b1a7KUnZnLIbnMu5ZkiYCODjbYMK8qB4
J7xhM+DY1xd/mUglxpwTyAmcLoqzGcGDIxkKlNuSYrfjNyW8FyeHlbuHFzbdgEPQWQu+/KdekdDv
wWE2tOgGKtWa8vgpuM3yrQkuKoiN5duudbxwsMGkRYUXaBCRtDQcbr4FzY8U/iWimgzdmOdiEfu6
Vclqycjs60G+dEVS2fEnVwfU4XoGB9xNhU1m5McxCKPkd9yU9CS5BURY9mCP+oPXmf0/LKuGtIcO
orIEXD/9/nQdSAJDt2PYwRUxyacVfInZpY+7VuQOpn1li5v+sOQzuwW2R7ZSPf7EorAa8lK5ZTXH
NS0rb2RYm0ym+CGBat5c15AOLhVmHDEjgw5l9IrVKipmEHD6nVWRm92oV7Ya0lwgCvzpbLqGjTst
pgLz2AfR2CcxIuiMMdWBfPIoE0p2xRkcH721WtuXZBfv9sq7iTHBWj6OZRtLrLjYnoODnid2T4GH
pcUIIKxSspZjZS3cFCjQo5XkFRghGh13DjCEa86XW6T/myOW1D0bEawCDNiOWeXFd5eU+Ti7mBgI
3dsvwPs5aMAxrQzv0LoVq7sGEsDxI7pzBSc0KmNfGXej91B/QF6yKS6GQCAGPqsRbRP7+1iNmSW9
QRUNt7Dt/SoCh2wOrBTmeTqnn4a2KHWqwWr+t7CFfgZrNiwS6SmfgvorVFVc0eGtMknNIsJmC4lp
68mQpwwdocdbM/0P+OOK1Mh6QvJRVTlA1pEmC+U044yDr9m2AbnekmrANdujYKUHh2Wnf0XSZ9Yl
4UCcf0dNqZtaYLIDZaUhgfb8eTMqdc1SgPLN+tgAg1cbE7lsrwQ3cZJz8OaZMGPHYMFTx8Z0lDZI
cFugRFvdOlUbkhD0HoURAyl8+foDgWCLNenWbI5uKmqh3i/t6ilNxgmywIxq2kNEqQcuHMRGUCrt
9ZK24XoETPAtY4Qhd2Sm1Gb+Xc2SsnSrJI51ECEXwYlbwyIDsoTXlsL1SCmEfb0fIX6yMz05Xdn6
4gKwaz3QF0bnPiL1dUrluc6oqmegah+OgWzNr+avRnAKxSRpuCbjMKiXMVrNMCpDB6e2wObMAR83
dCBuB/miPns68i4TBbrd5+W0sywo0utCojZCfXSpOIWwXjo/NkGjjk9UueLwge0AFVW63nn4bYQr
/pynna0xSPtr69mBRZkQmqulQukoYlzJvtHCHDn7AQmzcM2MvaNWqMAt3nEb7ywaWl9np6k1Q4GJ
+T/SANwX5uUWTVqFbTe4a3cfoucysKAOHUjq4ieAkb02alx617C70MuKirVObDurc4QdBtgbdar3
wUwh8VueUuNEErVqAaQ9M0QUwCIeMdGTZyTpcZQKU5hkcJbSFsZLzepP8HI74IPW28XVJmneN9z4
7Q9s7BqioQtkgcrkAQrrmFSZ6VBr3eIuE+/kxjwKJXpt8hhwPBYUzcbhg05Nr4xZ1vg3B4ejIZvx
T3t3Z4rL03wBkzPLK2IWI+Cp5e6xJCg5byb43AWdPmWqgZniC7dFS6MiDVuXbgVK3w66rtYvjt7D
YA5jxg3+uBP1uCaEgkWu47VRw31NWchcCBZhea5+/QpJqAjlkpMQRc3Eq73JSiL7MtHmhgXZY2EA
b4Y4uNBrB6wqg6qQUToWD2kga1Xilul27MqdIJZgpjsJJx0yVnT65yRgsdUBbfQqsdgfpiEXms+N
tco/2ZQclLOVaXb4SCkHBrOXwAg447Z9LA0JHVjFaNR/xLdQmz5UVVPrzNow1wP6Okb5EvPjeHHQ
83meC86qgN3PxV5Hk6uosHYXdHJ74RRraqdCnj5zPALJwGzk5d1/3aZHTR48+j3z46SxMIV2A/1w
6r3q4RsGgIgaEgLFCUwGYWOM9mITKUEmRKi0kUbDh8z6bHs8Xz1DvTJg2EziMEjaon3C00dy05oO
tApXnpD3vpCgzoA6M4yvVBLHhkAMJK2G4VQ+NWGp5w6uyah5dmZfPDKcAKSjU8tKEtpGUtSesbsO
AtTexR2pXUke0HqEa2TjBZkhD9+47fC2AvGRZa6ZRKYd4E6ubNdK5QrIB89v4TWsFIYrUoOznwQR
i8GT+z51PJZuB+pW/eScZwJLwfD1ObYED1P11fiBm+MWcTXNm163qdYWJjNgQXbVRqPEJL6sm59E
pmwBErURNIAiJCTbkptcOVMdth60E5K1OT6kuGQ5Z7jvOWD07jmihaTVKVklTd2vi5jkKz7rB3kf
TdSP8Yn2okih+pgZmmDMljq7QgJ+ikQ7RA5gn1QE0BLMBFCw/rAT5BhBisKlZnBAePTbWVnWFcoJ
xWPaZhKTQB2cgPAxXHr4DuUZG8qfRjhs2gBxudxuhoul3v78J2EuwOBe7GMDgEe9TClbAI5kAYYd
cD04B1tbKYcy9ZitwmPy5on9K22xH/QqCk7JS7kQ1kTW1RwXudj89Bt23xtoXPK/QpzaqpNMpI13
h1XNl5ulLitywlZ/dsmT9o9qtGSJV2Fll1F/rZOV61KfDx8ZnsCc52gVm8szh6ueN7wiLpvwAg5b
yRUJHxULJzIbt5Yztovt7dGW0Iyy2r0FfACZSrIpO2Uf6qjpwhPecGGJJVz3z3fcFarsaD2pv5Sq
BxOZqUb2rahSVOTbknU2XuuufSMjRbwWZkELtOs3OrUIjN2pOp1up+HkknRRx6hjNDylvCzSRF1m
3NnMJ/2z/S1OqytR6+M/5CTSsiFKrlSpmAbqK/4An3OxDRVmL4QBBju+4Asql0kmDHGOLnzYWK8x
hVQq/twGaZHd+hCE0zDT+Vo5nUIq0DVjThkkPbk1UGMO3inAWnReUsj4EdMsGe0tqC+isPm64PZU
/z1tOsk6jpXOrHWBqG7JA8UVEsVTXkP9pgUJpZ2fcFnLetfLMnuji+xYo+noJFAQJ4MosDSQK1Z6
WyjSVU6gJr8pdKfPSsa+Zowhbf6rpxqYJb8fAByQ5fE5HUhlHYhTiD2/F2TbgzzTwdnQ438EdMQ5
tGSN1o1DCfKaE0AnSPkS9tiBQNtJxV9AoSdkcsOS5rk6lGNwDVGmD3O4uE/G0jHd3z3kzI+Iw2oL
OxmNzJAjTpxxA/pagJKe5lRuhvNYwbMm+UE5S+1QtAE73ZkfAr8OAVuKSO8US8q8bvp5RUEW9Ao7
l7Z1UVnbZn1Wcd15PtQa6lUWsqcgecwZITX0/FoLtXR46Fb4kt4AJVr0M1lpeom72NwnrBdWaaJp
U3Y4w3jgrwrAOBJiKM6A3u9qAQuQY/uE/5EI94sHT5BKeZ0AxHbXfvXZ6HTO8hw6XOxlE+SV3qWC
Ge+D6eSRczWo0AYJL+3M80SNZSg/jL4nS8+ZNwVEW/9vTOg92rNg3gxS0rLxY5iWtsIq+9+/r3hI
x7HzP7MPRKj8+KVacxZXqDfWmR12RO7Nx3jUvKR+F1aC24ZCnZ8pZLJxs/VWCZ1Bw5nFWnZ78U6O
BXRIE7+nkQ5cbrdKNaqQKlTq6l9I+1lWxt4a4poL3j8fYkxC2qhy/djluLYzJhy7WHVi8gBs5LlG
fpDxZnt9VdZIYK3ERoeI6z1BItrRepgIPCUTvfVYUQnksIR9zvvZYt9ivrjEOTczh1WB+YBa8uWX
rQ5PqtjpwmYSduUZWC7DccttX9sOhFsQqQM5U5SPIeq0/S4DdYuN69QRjackXQ1DIv78q5mEWY6I
CTa3z1Z6gLad1LuwWL4dl7xE0jKBaIxfAXQyTpQXTSw4ecWShptSQztUyxENRX2yzjcWI3rIgNpV
ubchOQygeEdRx3CxZnOId2DQnQIgtEETaZXVcde1KH48Nvy2cIUkokG7JBmNXLEOxaO6Kv+t1V/r
DvIiR5lk4SBVRAvnEwqE0g8JDg17Y9ySCX6UCzMDhUhh6xe4ibJfXAO9PRZJ+dcSINeYvn05Pxna
PjzZZR2PwGFsiyl1OSXm2Bf03k6jaRaWysj4gEeVRwQObj33yPI926EmbDxzA74y6g24apHbQmB5
acuQzpgsei16VPB5izC+6hzLtHIYavmBspPxU6E2VOPfnH+1i7YxXow/GhTv0NqsymCvY5nVw6B3
qKYWxR383jm6Oze301RBbMh4vjw5aHkyA76A1sy/7iU/T4elgEPcHO/wjAlNrO0tmnoWXQoikNJu
h5Lsr0SH9mt7yZKSDVvu3Xt2bv8Rg4ubMkgTO13FxvwgNmWvU5BQRqdg4rYSyP1AZx+hY0LockaH
LLsJR1oP8m9TfuiUpq1q812kg7W/mWzocSk2tEK55naKaiSdnHEWcnG2IZQiUJY1+Llo6my8Z5tr
DODDp+jSM21lXzvOTsm+3PiluRIrsL7Aq2OZUWSa08LUhBkBPpFTlz2TIxs2DM0jj+k7OpcyE+YD
OjyBzgFrtOG5Wmpbu/T+J+GNmBy+4CPbFzj3bjzJC9+Z3LhkdftuIhW+UjsEt98fSIbPHE3U9cOG
31gt56eCKB/JfGZ5i/VXWVIaSitIRxMf/9MtBC7noKyuL5mruJCyBE5pkbbFTAtsYl3ebC05pdsd
ysMJltD4HizojFiBnlHhiPQuexFKIsRc8maCaZIrTWnV0jQkTP/6X9xYT0tGp2UtZY/UuPJWndBy
lv8s/YOtwJMPVgxHL6pw/Q+io00jfA1CS/1w3OVJYlpiV8ztEsGbf0Hf9xTROM4Ia2UtW3W2N25I
Mwqy0w5NSaLvWsllYEW3TLeYiTwK1ZaHJmvzBa6Z3FwR1GIZwq+KNDgGdQHa3QHDTZV9CeKF3hxA
KaTu7iSGPCxJxdhhfqT44DRrtR0K2wNisJf4qpvQm7WQfAo6n4HJmyPWWMfJfzROORL6DBDQjAFy
QpeqYSuol8fZSpYNWF+jBFBmOORCkdjzu7KdqQodphh4H0LaEYzmFs30TArunolKF81nZRpxwXWy
1DW/AYBotsqxupvuMY/FesiQCulkP5VmnZlwDZeY9RszTTCqSVX2VoJgz1wbPhDFFOS/T9SnsKit
Ac1p0Pax0O8VHMvig2G97gub8TM2K+GDpIMAxqA5LmAYJ0dgBeNEWmcIcILXQCUDDbZqXrIZn4Je
YO+8cTO0oxAlRJHksDC5gwP17gSou5aq9nHm7KKBzIQzG0ZjpNT3CpW70wbxlaLuKQPks4P2fEAM
P+ads7pA6eTaOgLnmyTDglKCAmNhTAzG79BKVzz7Js7yTaO4zHiUc47pjB6qBmnFE0DGs+vZm0UM
25ks0lqOQi/iMXRrjp7JoHfUgz0+gug8WjAUDUou1PN8zSR5zG1wqB3ODsuI04vsMX//wImWMwI8
8AJjaHKVLpLCd6wnY69WN7AwGq7H/f9mW7TacvKJcRJMSaBwf5cJ0fQ6SH6BRZMkgPVV3+B9yszt
gM5gWN1Y5gYBC4gzW0SGYEBjt6drDuHHSbBAIZmedkPDoZa/q/9RdylttYllgXrY/q80st+M0H0R
Z5hKIYV9SlA11JcbDds3WgTwunjas4JuYeZCAUUxClS4SEq37gXZl3GWmJ0uOcOCY04poMcNzIZ3
bd407CP9ILRAhKihNSW9VtCJU5609KtkwZFfE33FlJ4cUcM4gg3M0Xsvz1qzY2IVbgwu/uuB4qQg
8iwJbf9+bAZ4FM7B+MeOkMA5j4e1Wd0/TpABYgShcINfzfWlruJwtgluARf6OwZMEHqp6sBquvu5
zbdALqCTFRgCySCdWSMrM/audyAdaiNJJhEke2P30EDPjmj2GpOuBQX+z+UKak3Cd8ZnwKxxhWTd
gCzQi2SeYIrjbjgo7Wd9ibAfq6knZCIUq/m7I/KeclJci3sjcZ4ejj/Tv82C/IOEvexQV63FhZzB
J0mh+OR60LyLkCrvlObNa/RzvCVDxJXXs2WpOytr2eH5/Zbqpd3JVFY8LR1P2WLAjvSy6JpVD/hp
XFCHLpO8cvMyRZYjcDjlBHHLVfSWXEjKyw8gaRyRfrLJ7g/lL5H8gJR8SyKCRsPqaanwh90+Fy28
gpYhBm8rHBPwyGzjcKnvpIMs2L4OECZ4c7Zm0Ht+5vFWq979vJqMESPCFXKoZCErJSzbc69oBXpD
us/zs5pnPUlwZdVKp9CmGW3yj8J9KUm4Ue+YrkF/lY7i1Xcwt2AQZp5FSaehD1N6kODrTRajOudE
FIOOTfVzgUUVKm3Gs/zBdoGak1ws/FYJjTkZ42ZOmb6OQ0v5VGIOLI4taGKMr9doEe62sCaGrvxR
o9Xs8Hndg3/lEBcl0uAZZD0SIzmpgJ1gqm0jKcpmnZK09NJP3qn7DxNycE+mllTpQtQpe3Dp9OST
qNYDAskHVXihuY1SMwT0usx+oCVTE+JD0wibpyfjFhM2F33a1fz/jO2axxVCMw3haLbfs4NuPW5R
HzGqk1gamP9OnG40KT9oeb71kz0guSyfxaB6IqgfSa7MKEqaNDE52cy4geNyZzu/esNTUMOToxV8
ads54X/KqVqo1zVXV6/d+dnb+CIG4nKNgK6T2s/82PZ6AAXwXMiZRWzH6P1LLZzvmFVDBwXrwlcr
PM85fHm9PFbeQWpjf817M7L93SLgdg22GrRpTo1t0N1zPnXfyLorXCz7Vm3CotRhlDej3zrbdV/h
i7EszU3+SJHsPoUwKPK3LQcBk/VRIt29Je+mnqjGU5qaHGeWP9jaXDjz5e5MJN3Q3stMpc1cCbd0
Qn42fbasX89XxvBir7nTHhCEkBk7PbXdx43J4fDyjWBLsc0ZsjCHkEq5gxSZ6AXHE7bun1f02ezZ
N4yoxkQtGMvbB1CDOt++Wqy3wnTEH4bxvRjKf0q7s/HLD5M1TDmlbM7bhm2TCCQ7dDiYsFmSFJMY
a1gYcB/jAhLgfk3/C/oYuH8PqGOjpflATRbUi43qfzuBqa6JjhCS7WGpkwYhiaV91eJVXqS5coBj
tb51yj5tvqfMWawyu4TkYHIY8S04pVE7c0CwKvdMZpHnQIkQydZoL4LlA8qCP4+0bV/nFketoHtk
nwv6X79ETatzno9o3ePzA1cCfpUZ7rA2FfxjrqlmMhGEkx7Z37lY6NyYeOfZw5ibA6g9DsBEFRHa
xks4k+z76nKmsJRAVFzxe20g4upoEjXytQB7nVhuO3ePI15tcT0OQsc/ZQnMmV4Q5TePRpPhpwpI
LU1jsEL0TFNUSAGjb4FaUJD93z3IsY78lyb0e+xrSULWElK1c9zOV6VT9ha4BKNapKHpwbW6avnl
J07/S86WKD3UvUd7PgFRKaURiaesomKQN3Gr7n7DEwx5cdmhSqP94vs6v8IIHecVQYqPfV3+eLil
+6movJ7L6MQvsaH0gRa78vsnVXSHlzc/N53NeyVTjaZ/Ey0/ALjq0sxZwRKJ9xV4AcU5TGgmrTi8
L+m0P3iplBQIXanVAIoBMfu5R0J+8hMCQOeBuuDsVU3qeTyxWh5RoKWCC0fFWdOZLZgBTr7UF46H
Q9n66IKQ8Nb6Uh98jjTYweKUTA5Ga87Z+bAAuMMqR2NzJq6TMmHcJGE98qWULQOeA5Oe0a5Ydi8k
OVmjIIxj5Mds04O6Ipn9lUIv8MfXG9Zx8wO0JxcYr0ekYkibijIHOGDt1qikQFBk7in4b62K9EwM
tAMRv1NW9GL2YE+Sr5HInZaM9IZbFn4r5UKx7o5L+C+ClzlO6rgVfXmJdvEr73qYKdFdYZT6JGGr
K3TVgQ5/3KlCLmR5uyMPwfusfwlN8RvEOE5/zRgezKN4YtA09V96y4aMuGN/5SQoDqDsaniECZqf
y3yDTFSchHru94XXRqkrF5FsKc3QG1RjN/hvM1ciNSsbvcR8++7A2xAtL4LnfLZQwsDmdap+BZ/Q
SGAiP4PEpWqpC7MsTLVL7xT+eVPj78W2FgrP10oVof+lFbgmrI3IgCHN+ElXvFP6P5Yzt5V3UXwj
fMQTzVQbm/tb2KJ+Sj1GSbRuwAGAXBsmY0i4CaJQij7q8xLY0si8lD5TYo5psk2zSl+s0OCSm7U0
vYNVC00PBWihK5qAwQRloDaNlbDOO7KAY3nmif7LdHViyliGcWAlgtqH/rYZN0VEf+l4wxBCtN0r
fSkvQxpo60fiZrZ5rJqTznmTSnkatAZbZWK02l8AcNpSz5IRl//0SQRAClRRJWrqqpqfCqAuONr2
HW1sipMHkK/W2qR9ONiSAWhhC2dKY6GVTu94uiLoDEAJGJarEquRZfrhnsmjaVe2bKyP5NdmPs9j
0LT7l6Fwa5VD6krLB1wM3uIL/YAgdI2RkIUsZbnVGHWcbbd0n5uDnWghr0EBp7oyCQIMn8QWO6RJ
TPqF/o2PZitGuz7CyIzzb5RzmdHQDLsTATi7fndopW4hvNY2uK3RhPpGEWNj8IlEjbf4FE6U2rai
STLNqWVP87Zq+x679d85ZzuNAOkiuVWvkOpM21N3EGsGjdmB8+ZTxV2aFIDbP4mWsYDiRHwlExTF
9duMI7Qr7GLHBsKxHehZ1lrQV98UPP5Jk3RMEA04yY5WNjSkpYaEeG7/VFAXREVEKHOscqaM4vAg
xOZgZ3yMyFyibvOdxh5PdlTOtg9e3ydiuri7diplsoWQR65VkF6IYzU+Wcj6v5vq/sybs2AR/c1g
LClEiovCUK5Mag9J16+Ps5qxyA24Y/R/7MU3QLVRG0K5/r0ePAFfgIOyMEhYpoHVWPYrkYyBLUFA
1tESdFWGnYJ1dQ2pT0dBsW0GUlumLDNmWTzOVtQVnLS/HU7aN+mLdMv4+5EO5LpOTdkk2S/Xr/j5
saI8DNhGW7y0dUH77t5salFxJYoH6pueJipiXpY46FF2jeymqCCkqw8v5TQRADlMUvGhkojbthJR
tdbfS9ucIL535geAzXcuFXD/jol+rWNXKjQRJNfLYa2oeNhfLWJkFZYLVvQF37o1YdoAVcwmAdLa
maPE5RjUHzF9HP2vltltF3HGKrsZmps9tj0Bb4X5zqG9K9QxBlH9BLZqwDxf0ZvH2sJL2fSO/jt5
Q7GuSTLHM0PcQzQowWy94R0hIpfViD+2ZNjv+LoJgqgoHRp9NO/YfA/zeWY9OpjCbqGM7mfbHoBY
/jjuPHZJnQBamgooenFvRpZWuObVfcEsHV8nyoVULnhBlZz9ibmPMU8DenkG0Z3/rsxo1tVsir+j
byglauYULi7G3ddB6Qe89/C8lPEhdjvr1SKCfHe7fPIma1AOt9CF8ZArJ+ztVtrCUiwRngi/gisN
LC7lZkJXtloMSVztelVUDNWevmPPivqFLraWwFNyZ6HWygSSxjx5aPSo2JL+nrxMQ8FNXc7a+PJx
eNOpv+cZudm01Felh3zf/ukmo6m7FiD3JqrETMFf/8WVyJx6Y2flQBuR4eLPGGSkMb7x/8F2D85Y
ETeXdFppifsMM91EGkpYDSh8iGcv2MXzbixSqFi1Xg+L3D9l4vgVIMsrSJ8RbxrVNhDDX20RH1fz
wxmD+6HqYT5sRp3P9Z0lm7cr6Xy1WOLoXxXqGKPWQvGJj93V1yq72tu9KyLr+WLJZQ5tgbBdMLLT
FuM2T6yvA0Q58DpU8SBdo6olTPLFuzaN06PzDAMz8ig+5+s90ia4wlo/F3zACdd28IRvALvIglBH
oqKZ5Zscf7tdat3GTiiaPPk9tTlYq858XGijPk5Cjzjx49nGqTZadQIBgqOEav/Dy3wDoVz11zuO
dJo+uMcI5RrdnYEtqEeDEflXDTPxvpEbYJTvpblHYzILDc7zmQgFkmTEHWl57anmVgG8RLSo2ezL
XPRE2WT1wcvD2wBGhqT1DncQ/8xy0Th2J9Xuda1vv67tPfHHZRkHIJKSbw7goAIzyl4/8LT3eLEg
Ddxl5dCcrRgM8JQF77Wo+aQo0a1Mlhmj2hT0bnP8nPEMylgVY2KV6QVPV+VTVFUlUx6j6pYtxCST
e2fBcbG15FOgnaeiURdkaFXvqqFOfF+I42Y2St8FlZwY+k77nn5qFy0+uWlc5z0SwoXg44Ybt49c
5XALxaf4PCxxCBJd24+TR9th87cR02j8hlzxc/400sUyf9s9P7v3ALxiEEWvTS7PvxKJuAmH8v8x
gIzcw1UGgcZ2HdT/S9RAvbbHBgGHU7zIz0txw2dgXHS3Jk/SuZ4/svwLXDnB16Lkif7rOGsh1B0i
ZZKtcnM0gGzu9yel1bkMrT9KL7e+lr5Hh1fcll1sSdqUu73Jipel0MS33jrBNGXdTOpxNaRdjMiq
uWpwbM8N8Rd4qF1sjSw9bP3oBhVILjU+RuUOPxzmXU0XRpjooZ+99H6+sZLK/bLA2vuHNt+qaQVZ
BjRObb2DKfbdhbIsAO1053mqavFDcHXRpWXzA5jDUtPzwzc1RITKF03eI6gjf+kZ5XK/jAynGYWC
LqIcxcg6Wxd6XVqrijzb0vyX6q7xrjgJZKfVkGc7zJlJuBoKaN0CTI2+jyDOzoy2uxHoxDTrvhTM
7QiDgpYNKsYI/HO66H4USzmE54vzCUgVsn819pvhEjdhFEl3vxEIKAWif9NO9gSfU8ihNwAkvRyg
EKpamDDbRnnN0cyyKkWU6tmpgr/uaM/wyRyngH07gFWSNYVYINkWjhb5kGpj1XjxZ3HXlWzgyiX8
jnOg28UhNh3DbQwRCg6o2SE4YhWyZ2dawYceIlHgU4TaGZWRItNzcY1M6vMddghRL7e5eNcxt5pO
7k8wcm0WRfGOqBMkc8E435DnCiGF5dC9los6xArGNlNmRaMgc+MtPR1EuOYJSlGiL7zhgUwoDClj
KHrEQamy28tO01Yno+4BJOq9VfgyU1UTddbIBbkEPlEnoFr46PGF+BAjaeGoPpVAyw5DJfNcUNvJ
0JcF2diL4AGUpRENVYA1sBH32WRp6U1o8pH3aYIGNZMo84PNURzTnMTv9g72DV34LtrsJRHEAbPO
uBNk6WjUAwdNv4jJsF0ryzQOj058hwo1wzDtbk2GiyliWPsnQPxhaE65+6LABummnANUeBTuTnxb
coXCuhCAzUJe0AtlmkUzpQo+KCYvVBBIFC7j7we4gJzzIhZKYZKvz8BMvGO56yVzSbhXz87uP4in
Gr3u0HA6A6fCbpgT/L3vsxomu4kj3wtZXko7eeanlPYaMURO7C/a8ap2/Yd5c1qNkgjRHb25WH8V
KAlP8JgoBrJyUwUbtfc6nUfDR7uWMWv/MB8O22a0pBDypKhSDrEJkY/R49DeJNE1M5AZC8fw679L
UmqbS16JJZvbgPFPAZhZBdHivOWg1i3EMqj179oV+FNLEdO5C0BkHtqUWQuEFCmFdM4KGFqgLy0I
f7N0P7AQtUdLm7N5b5Wqagf/fv+bl/Uop4RK4qGkhUOkvFC8xpbHEL7n5LzyctjY6U6dp2f50E64
5U7GIwrsR6ADcyaUW/AxmHX93ZBIedsfkyEVHo7/usyGCSttKUmSd67FST02tAycJgPcqfLvEY4M
aThfg0MUufPu1Mb8qjnVn1i71FFMFJPMkMSzQQdZdEMPIo+RWSEUB1DyR85p/uQCP2UvVUTe/d9a
EGSyv2i/mOMB+tuBMvMil65yfa8qbxPXwp+DTGzf8KoNzYPCJt6xwMlFKWAZpPAT6PcFVUJmPGed
40sNBiYh0vhIe97sUDOSyCCsbOSUkFdZYzRypJ3jyFvKT6NaFFJJMaFOBtvRQVG53JYTVv+C7SJm
Ou57jQTCumGuqtNwDsYFS/kpikCT9MHMG0TqBWCIdhq0huT0djf+xrze9Fo3ikixAndU0g+mzyHX
o7IND+KmspA51LApNUs5N4GEQSp7LGItiIWsU1WprmArKGF5a0MYsi+BuXTv39E0NruqZ7UO2JnE
Bp6AQepgpq9klOmIVFJxuf7be855Kve4k1dfIiIR33Ld0RxsZ3WF/Ss5gRZR9dyC0IoAR/s0AEwo
xBTKt8QlGnPxlzYjxFAQ43Nft2rulvuGs9bjb1YDyoU6O/8HjYjB94RoL8bF4oYmWMocyYbeXiEN
EZEXxu5t45gBNjn62kyoiliux+KfE8zcBnJLMK/Pb5bTZWw3Z7HyCdLIV41wzTkGYsWvPk/YFrJA
42qkcaJMhPu22SBvmo0ddQ8tLRdygzqt+jioITHzkNh/yOj7JqVbgfTYQ2xkZvieTChaCyZ/r0Dc
Y3lTtlkRghvn4i4x85kK78H14UvZpwmUJe26WQWHeNH9DAt44MNWC/x5F5rMk7kSyWZDw2pewNCF
wCk7ndkE2RCR5P/mYpgMbfYX+nNFpRa/kJ/tqrwkhyD6EBKm11l+1aHfJUWZ/pDdtba1nDNLDEXG
9YhqXCkDiGobCu/zvYBHmsNpW+9PwexNhil7FhFcWeUpsyXKfXaBDpqiAE2hVp7rL05u+J+/Csjv
mvK5jQMNEvR3i4mIOMvLWRgbq8ucx2auVz6CD+cgKzq+oT7B9YnKBpkS2ZOe29J9klpJno6MABfD
q/KlQG29ebfDGRC5kQNaYIvXsMFWlFiJp2U67z6dK/LERU557L1pJmcKXHVBC3LBvAjw48f5smpa
Q3yxQAk0wN44iNEKlwvvDxCbmEo4ooLWMBkwj/AQvAuOqv8TXTkK1YzLsdVaQyQOOsLW+MI4niQI
0g9o9WDQPcZ57dQikPRzqMMGMyvalN9BtiWLFlZbOkZQOGJJP2j9lMd/eYAadOxzsrltBdRG4Xax
QbxjiZMKtKX32nue/5jB1TJiUiq4s1Fv36zJBfXFGuDJdo3jb8YxUdDIKW66HGnOv4duDtas7s4t
KBX6N9S8BrINHHwK8VEv4WWwendKdS1yVYKTVXQVWTaCMU54SilxKnu2WWE2ERZQpDyHCprCbg/t
Q1Vfq1li/n5I6tclefSFhchQLJQxLmEql07zV5nCIPHcZAEe53zxF5s+LvPFypIwX4pjhPt8Ybkf
0/8IAib6f+/p3UyCPHfWcKf9my1VJWPb3ILNEP5cR7SuWazKguy5TGIBAhsbcRAS1nw9xcxBUejk
c78lX3BuYVNwQ3JDTsVMEE6x41EPuE1n26R4qhqQLZfOiclndvYmUw1bunKLF3Q9JgUkdQaAk0Zh
J2l3lmrrKB9qhLSWwq2kP8V3iLTqMmz8c9y4IDmVuoGM1enL3hVWT7xW+9szMWCeeaS7AJwdhTf3
QHazFOD4Htq9IVrvHWxb3Pex5KW6jMoeFIFERvzgysSsCoykNt+hw4l9sRTQyQE4QG6cbsjnRBdZ
rFR3yl8BHcm6HuCKCQCWNaZDT0dizE4Huc067YgMwNHH9JisCay2q/vNUjbrH2TKZE3krb7WS3fr
ETfh4VXDWIeLQmGLc2GJII1+A6f+nD87hNxQve1rbpDWwzASDeEEsm/XX/9kR0L5Kb/z80Ufgm4M
i2ekz7XJl8Ib2EuyM9e3oh9KwjTAhwH5fZV2IeRtE9KeUO6XAqfRPPNTXjTj0JhNeUsH/QcNG1M8
yN2WpX7OxdA7fyN00bnCGXc15isDdp5SNf1+QLmAo0xn3jNHDFYDG28H/OO5Qr5+0lt+rHMDA4i3
ia5Q+ymASo2HZJ7AHC1mBnEwuN8lafRI+GqbEDvfcV4NIMwjO8WdUzdNEegXTO/mR/NHN7zILDZm
9H8YBzNOg3dx5CvWIDGplNJ4peQNZnE0YozI2VjXD+qiirEh68fvofpnDKbs/59LFWzN4yF5kO/r
etXCkvz1sCXIeZfx03VkrI6gIQ53Q1hKFQPIkAKWtysLT0SD99mWxw/gnfUAmtXuE7VqgWedeUJ+
jc+/s5c2nkYJVSza1uTrmGCI6SSbB0tm+Mtg7R/wYwi07S5eKmQCGTdaXcDCwZQ58iJ/kg6Z4648
+cIRkXrqVxjx9Cq+uS8wHW+1+wkV3gFpxziuOL97SnOmDs8ebBK0jzYvjVHvckhg/58URM7AuHbV
gRh+3O1/5DNSLBnlRafIwwdyFDs21+jdnx/MuiAoBFt/smLH9bsOWZJK63xoaNeyk+8ZSTeEk/1k
XRtpzLND/rgatEE06/nv+5vinB07NHetVZTWqOpv2+OIKebV49GltKqFtffILtRQQeKBnkjl29k9
zIw++6A4l5gJfVt+w+4cNPb8mnX3qwuqT19Eju8FTrDOXaG7TW6DdGZm1KhWU2+uoErQxJCAU1uZ
fHCrD0cAU4CozI9adwebX2x0ZhGxp9JULkPZ5HfpPN1zW4WYraOqMzBejl/GGp0o7HXiW0UpxnIb
nuTgjMaktgXqsvs1vJ8WKNMbq2Vg4yCAf1ZzgKecJmtOCR3w3n6tdDxz2u07ZSZfFZnndtzLMEdC
qojZdXMWH8rxO2UvUAltzY9UNiC1h4zeGLmQIQ8Xoo44oBkibZ+2JEyQv6AypcuVxqXmyDnmQ32M
wBp5aDB5GPjBBumOTeGU/LI3LxfmcGDRX2+PajNU8gfIIHM/9gP6TUaujCnVLRMBkLcqNVVkEJkk
Ec/7RLIHio1ncgAjqcah0EguDPSn8HpdDHmmicLZtOad/37rJ+MW2fpn37fGeCq2RkKua/s55RTp
vFWtVtYTEESMZPKIYGiTWIe7CFEYbzCz2eLCBgwVYYEJbSRRx3K+vC5NqsgFlbmIRXls+FMkkvyO
sq3Jd9l5fDRzLz4RiXvK1pROyx7oAujoOYpRcP+RhgG6J3upUWD8bCst17y5Kv9B496Jx5nwNGFI
sfjX7KD1vfYZsrJMvxjPfo3Un46tYZHbOiQQne3vppn7891TmsxsawAApdHKKGBQLdFNIiDqqbBc
0oHoAuTVsikRPN0yzCoDTAmmEXI73RH5hz/Kmys536DvXgOaPf8jO515oOnXzfwyZtFwHwOKpCrQ
qmhRzkdQyiZtEHC452Mwm6f08UF60mUmsphJCalVyeaxr2eCBWnis0yCaGfRI6vUtrrNEh2HtFPH
tcnXrUcAgVv2kEuzSmu7wobLJeTZReehrfq6jNhiL+/AcC4aCozOyLhgb4Vm7uVa0vp2cY/O7Iss
vaEvdarfeGM3LLTJMATiU+CPwGyjKZSpm3eiqFYN5Itr1//Mq7GKlxgBFjb6K51SH8XJuFC6GXEH
d8jSsFQ6yAVB0/RWJLuULCpLso6wL2dlD8hEQd0JWU/W2ma5VtPy/5wfEKyrfIWjfzQLEC+D+KKy
gnw+IYbnszjUR6tTxZBw1FSLe3/BQ3JJEk8E2jVP87UtMwiyUv03+3z2FxljYwO8exeRxlRWi0vN
bEYuBFnV64MAT6C2da6XkFGhGzEECa2F6aUI1mF7Rn2iKU/YURuFVbf/0pbpqOnXY7zepNsQYH3q
cCYudOlV/8Z+388makqexPnMtgbj2e6LOKZlbLmV8C8WjQ8NhptqVqRO5kOn90GUqqSIQCVPEAXQ
YzB4f0GyvnL9gghKfM6sTgYXpKzdFvI0CToz+/DXOzhIDPkP0KeMBEJCiuksrOSknauf2k7HLeMx
ISnRSYVJhBnd1ewjrTa/Ty9a3/LkizWK8DVT6cB20aX+YQ6AeBlke83Dqp4XqrC36JPZwqsi9H+O
O7ByxbGWq5X9wAAjnXH++6/Yqbm8D6Pf8n8UDeDD3xloxxZxiNMhvup+B3xWMwYso9Kz1NVqQJ0Y
nebHplm9UNKmkZ8Z+J76lhRsriFW8Jq2PzPMJMrFHRAPRv9Xb7I/xG0Dkob/L5zJV+RvQ3/nQWbE
p2XG9RNP+IMW4RpaEjhUmIvcY43jUy0F1t8avM2QykgvYYDCtykgGZAAJ8bfCcgCk/RbFD4fJOT3
7Z+ww8zNzVWqX+/cPqB1pn+EgPCaRYJ2rKNUFpiujhtdBShV7GNZKnYUBoTbemtrhh50KM/mXa+A
Iqq5NP9zx04695/pQ4CQA9lYwGfhOOv2/5dCyiP60W9F7Nxdyhwlj7mbL4jdG7zEkjqGMM+R+T5y
ioYC6ZdrS5b+ADKnJPDI5wR6i7qJNj/Yu2xtdBxT7yqShx3aNB1rwDscjDjmsSEgNeXyRqIgMjaf
ueHeYfp7IHEaFT05fxnWsN7dFqZoDyK0EHLRYJd4Bg4LjQl0Ue66/pmrAV30FBDUG8+F0w1LNYpv
ru1ygfyMEPRenuYgtpG52de1j+2PR+xZjUjjHBcWQyiX0Vm/htsdtRok8WKRyW9oUH3Z8fArWMJ6
E4FNf/QVnSbGR4GYL1RaCjfHaIju+MRLm7F4Y1HCn8lJaak0Y5u0Jt7bIvsvUbJwYdtN4RaC7kAO
gj3sCmEYRjvP2Tlq7yDec7f/8cuoB+UMYP3+wYZyLscGUCbLVDloytSSzN5UMwTHsTwlLY7DwSnw
7S25lujRA9vOFvJN6d5DDtLDYR9hHOraTM2bwFDsVVVSiTaokUZ56cUOYmVdosqsYrkSv5q0ZcTG
YsSONlUA9wwW9DGoQ49nlfh7Mdq6rmo/geBq6Kp8tP0DmO+hRx9KGgNyyfy39X/To6BWCasubp9p
L+Z7uhx6dAM2QEIZbAIKRf/S6mToJc8uhmMw4urmTgbMShm+TsARIAB9j1MPFEmB6+yNuF8lbzZe
1RMH/S6Yy1+14B5iwz0AnIIB4UBgq9FzQgifZOycNdXOB+efIF5L1w1mxKf2yHbNiOdTU3d8ZyDC
tPas84GgZwRHkIfK6o2F/O8+DX2qU/Kl4VgVT/LOCPDfQ8/DxzNtsANUDTluHWdaJOl9g/n/0jYk
RBJ9EPKLZrhOheP810tMeIxPEzMmqOYb/4nbfFGRFb+urhj6hpaa5B5OsOxwJTElAEuN42zzGagQ
uu2kg3wWs1YA6NU3Isoi3/BFzd3aWxqINp3wnw4uTukPx4n1sc8uz8gT9VX92rUSrY6sDUNsoWRE
tIvl+9EL67AE8WkJcQUAXf5WdvCBgWtVU4KZ7oQLILxAPNAffe7XaO5WVfJMzEDIbPr8AX6sWWFL
J+X3ZPsqgBvp20cQ/3YWsWm3A5w1K4e6geVOOt1ZJy/VwUJZfaGKKA7Vekxe+iaap44dV6xzW7fs
o2j4YdoFLmwDUI+zy9pLVPX/ocS96OWJevQ5K7TXPBSR3SISKbAReAGuOUv+6f2d7EEWlaaLc4Yl
Iy9O8FoZbtrbE4rwCplMFjmc4lsXYjJs60MOmkSgobWWFltNNrAP9JrnU1YaL5vQpb4g/xFOX/k7
FrfEqR424zsY3zH1zhe6BkDS132NJEl4odKQmeyQcyBdsZtS+TzndKKDIy/r6S4COzM+qj6XTagw
j4vQ8Oz5JAiF+KxdGQRHch73pJTojQ92MbuoZhbSJGCC4MvYuPsREjG3Tp2FjnKQ9WiE2FsEfMVd
HQ2JP3PndOWeLcblQB5R1bn7K1WMR4F+iUlqqwRUoUD37aguCUofkp/EGMeLCKiO92AuBcy8g+4B
HyEMM98NC7Wz/HLxqGvoMU4MPVsG6c2IeQFbJb33FgZvDVDQ07plUAHssXlS7iTcnn8nvzPNYkt5
uyX/CuDE0JkNl1SQyTJKUf1uVyTYe8pS0UYrban/1sS9MD3O1IEO33C6dSBMxr1dY5qSODK6Wa+j
h3hPfiJTzRslIhAD5ukOi64BNlHzEzK9YDGqoZGoWnvKxO6YdHLpWQpV5tYDzrOwwtQ16791uSh3
TwULjYCEa11CnzB26xUmk1ZQhO/SmQDSg7YuCtgQUdw+jZ+UW3CJPNGztRLv7WbP8jRMRD630wIf
v8E4Q75iCQ99jKj2VwknLPbByzKhYXwBltT2xXKQoVDH6LJ6xOka6+hwtGwlyeiBYWSzsnW/uumt
YSpJ2dtg5Ujwl6YOZ9zOmX8cXe4CyaxWcQ0qYeJhizbPJkqT3P7SecHnmGzMujjtJx5QewAtb4hM
3MbNcsiRcXlgkrtCtocaeIUyqG5guIAGsy3W+2jVXcR0pW+xiPKGB7JmJEhAlEAqwfHouizTylbV
N6c9BeXYBu+XGzUt9Dq1ZnwHMJPnr89YcffocClHWoElSZjq3XdU+DCAY7oX4E/wd68An7Cr5my9
bqHORxM+LbAgDiYAbo3HSHCwbFcDAYxGt7xdsArgzd7QQAWyq0pxx0wo9EroShEs02ynoFXh+qeZ
+ePE57yO/mskXp4VXLuVH97y2pP5O+b+NYIWY8hcyKiykm3ZMAB+9hyK3G1d70AxsKSw82CHOsxl
5YUFDaupQVrGs+c7/dpMZ3TgZtYTjId2xSWqJixrayoJUuaHCh74/qgBvA/uD786gg56xjK5d7Zo
FzjV09uwYVZGsmhvsoz6yJXrxHprw05QyRg16zqKms25gHKw7LaFw5ckW4I8ovzCQVM8fFBN9Kzh
QDtIQJHQ0BnuI4o5TOTdPSpq0QGUjDgTl3rly9eSUA98H/bV6AGSFBvKbahbK+pNeGANYEhlCFTe
d9rIISXjj01we22lRHdnmYLXOsJpejo9EbvRhq4STQ8HZ4UL3/mLndTveZa030a7s3VLTSm7mJGL
uN0NE7k70LjKk4bwSlcIYxRhk0HfXTVE8lPlDAdmg2XD/g6ck8SoTiXlTTZ2e1BjcqdkRYRT0PQi
6TnWM+6TKzkXFmjY2bAgbHyvQQKv7I2jz+WJ47gwMQiAAvacRRcIpD/adw0dNnCvtmgtCy6V0n91
u1A1OQwPcu5nLK2+7ivdxA7wd+gqj0VhXKwvdbIc5EWaCxK3XGV/z9Uu1pLMAqPU6mPK7P+dqIQn
SqEcFsWlwfuKYMc0OrxcCwuGltxSKHe59jkLJJKD3Yr+FHTmldjU/9nQDLSI2GGM51EcNcuEuclm
CU8GvgV8VO4pJcxRvxur9dOUzoXkJXdb6YGCSpxF+Dt2m2rE6wefaFqbbwwX7RKlDYAeoWzcssBc
NRql7wFHY6KOcTKXEWWWLV/YHoa1jeTkoNoXCL83ngEBbPa4oUlbjlQW38VOVx1BsLFAFGj8r8RL
YyzgS6k9yiFhbWKZ5rN1ziD6+eJaZl4f2veLiZZf8Tk3Ks+WDEKl0fHvi0fYWkLDrTikBZ3V9kh+
pdu61SNKkjLVCWGTE7julx3rR67Rlla+eldJdOtmOfQLuuzZs4MnDF/uQmNntJTZTfu/FcE4roIm
yIx8abtIZevxulVM1kq7ccgZbmieradYKJw+6fRdzFWvEfP4+yWM1yoe/4glC1ZIKStDVQY3FVF1
5Q915FlHfokJWNXhUyHg7+H+ZKOg3GfsrLUtVJhxLprQhwyy1rVNXrPH0kvAwbf3pJ6kJvHWu1KZ
VYEXqRvXtzHlQSsMBniW89wQcQphBqRrBQi7iiI2N1gbn+29PNmGaBv/TYEzBs9iFKJ/uocM949p
5eG/NzWo2YLo4hwLmT5CVGnceLSChxxrNl+AeoANbdhSvVuGBaK267XpG8bu037BzD4jcxGvEYP5
e/mIEEMdBEvRbGmngUhmBkntNInHrEFzDE+olgVthz+R2bvm6aKId2JBHZ1tv7lYxVh00KPR1Lhz
SxM6xX6PTeIZObYUpkp4xuoo+mOp0jrtgbi/JjRcD9eT7+zXJXs7xBYm0AWdKtFIP6g/a1DgY8cL
A8qYPieTmlKyGNTvvwj6P9HvgbdtydtielHHeSAw7J2x8HINq6uFuVjRX1f3ZMivAbnpt1gK0EWL
8DDVvG2ul7eub/1wjjX32x5CckUyKgRw4LMNz5d+bqmh4YAREFYR9caNGazQdOQXHkzs9/9HeTEc
550ZbgcrKMHL0b2tuHjCzATXQvieGlYwzO1OaMUBS0z+nG07KEK9X1hnez/QSXGGCPCD66J8byVB
JNvu0zWSfKzrbH1tW5IijeryHT0y/yLtqIwq7gUD/0jtbVtTO6z4FCFVv0byMEtvfuONUacFikpe
yvl0D8sOWEGvAKWYUwl/uCG8ayE8gNEnkqp/0uGjLhsWT8G0dvYOsz/OMzQBN8LFo6dVePHVRgox
ML2p6mW0+gRwcW+Yme7fkkUfsE6qu55rQwloCuXXKo5MGzfUSV1KoO8LaxVLuCUjNT4wB283Sax2
S8pKymvcwN0F8JBRs0IlEQdqCPbP5ugwzWq1EPVAYS9goe0tQ6FcyAqWTiIQ4jdsZ1NhUIAfMkru
BWdZrwZP9F/H4GxLwzYg1+8wRjHSDVGnu+JNPacZHmVGGX9DvAdPoza6nshFsO0jyhBQfv3oH612
tEw3bvY53K/9qt+XNY3YMJHmDXWum/VSewn79nUYFD2cQaP/Kvf3FvtmIVqoKXfmQ6XCUz3w4kQ7
H1NMOcmcXW/bjxps83LM8ph5wxkg7EMMwHazMWXwcBzvtcEtKI3NX40XGvxecFsdPoTjJx0FEQYB
7naN8J4H7cA3hmZjA0RCgIRWX9DYtKWABVGkVwCgKG6dcWUzK4d1VtdFX7n/+saP9Y2oIbAkMfU8
1pqR37dCwPJA1IeHAZxtH18s3COyMMXTl2Bv4U3p98POY5fkupdzFHvJ2jAXyojd2BwTyCyN8swg
IYmzXDi7YaroSAr8PBB76Gxatanr6/yNbyYstYC8i9310NkihAw0RUOiYmSOgXGJzl8fvNZKpU8m
MrKKQCqtprkPyO6aVW1pIphuvgc19f3oaUo3Y65WQDFyxM3d6csZWge/zQgj8yZA5ZtPnvoS3CRC
SBQ3yIahHaq8ilcmRb1rfYfdKdpYSlN0J2sHRwns7s1HpTS5QS/sNaka+/knR0VvvibJuGWjPMOa
AmMII6E4+bfBA2FeExhE6qm4UH2+WRRaFbjgZ99YV/d8DAI/6eQzKxHM1kzVzux+K9Ptd6usT9tw
QZxpa79rIS0AHGXAxAiYOYoEHfh8bzsZQNLDwu1xoG+mYgSBaMQdvY0tfzoH2SBb+rogsEjUkc0y
BkrksBr1ZdFkMVC45IMKeumTqHfRZIcmxUOmZldf8o6BKs3KkLAOSO5Z9Iv4QHrknCZ2/CuTLt5r
NQxgZvwKRlj9Xeq6JjSucNfCxQLhh+hat8v+aKpzi7od3c0+Nh8FkFoRP1/JK2+COsae5s77pBiT
nBh7umSGG713pauc2VoVhtUzvp1dKUtQT9sJ2+W1ozSVSbOX5NpPo6qnRAvF8PiYmaQdI9GwZ9PN
myueyCW4u8DgaYuWOoM8inH2FEqLsyp5FyA27H9dNc3o+PGVBx1cQNQW/y9LY83VL+SV/JjsXLej
uDpOC8vFPMWFgJI/j0NqSwLlOlHmOyCVoePflmDwmEKpQ3AE2Av1jBu7Q+HW5XN34V3zEXcnZfwj
B7wKkwl+vxlB9L4ATuird51Rv4eM6F7Z6I+DREUgaY1BT7p2lUDWpH96pNj+CtL/ocHHVTC0h2ye
xZq7ko37gsgxJyTiEkge5OjXYeQyzXGfz9r0jNw+2H3d7UsDHOrz6fb7wcgmfpGOJMHj8rttsgOD
YJrrBOzJOr7oKURrehYyJJ8iiaOjSpKlyjHlPW/ZbdhKww3i4XR8CLBEyVYo9MhlUuuwpsHAlSYu
msnp9b5C9wdeJ52qFsuEW3FjfX5VrYvlRg1rccRRsP7hAegVL5daa9nZoK+EuL9MEi9w/c0/BLsp
FM9g6FMOf/3ILF5GR/HCrF0hMBcBZlFXUnSGeuZsDOBsIURw17Su3Mia2n/1ec97wpcrG4d7r5k2
qEIEGa6SgwNnl48LsoroTOpJCRF6C0sQPS+npZ+WH+KZkF4UUErrYOXZiwRfJZBWj5nhqmx7w0ij
qjPrMZjJg7HlNuLP/8FtE/344NyzIqCd69ZH1w9IqaBHXE0C3qcxoAwGcTAnj3EJ4qU4BWO+sj+X
iubgWfrm7Xy90opDhsvTBGGNmD/dN2HR76BlHS+rRBCoPrFeVnuKsdzMlZoQfGkfizGYBLoFd+tN
A18PywsBMYxmRbKF/6ZhSUpWdUfzN00CiAbI4jARWE+GYY1LJU9/AMgtutU/IT0LjNLkqxMKrV2J
SCRfdW7/NxIYPd0XHFlW6cw3t5ZJg+s+YtdS5iqwxfgCgDpenrLvVaXcORIHZYAaMdB8LvfyBIFX
qSxRI226r0trwHeOB12KR9tK6OiASkO4L5op8CMq5e2mJKRi8l2jTXZDV1A0NnASvFmXAF97uyEf
/mq7ARy9ZVDAqAeE0AsLgjlNs0EI15gMXeUIte8bQeizQudcfHYktJN1vCqMp0TyJvSNdy00ei5o
6Yy//xfX1Haf2yQGAZY21l1WYGIeAvi4ngTATYg6G6iwIqQJ2bFPPi5WURpAgJZpuDM6ORzdno+X
7BZpaZB28E6bDXyBaeQaZeh1LoTOi2qEEPw5OJ7CianCFhz8qQ3fU6rw7a4LZGNFmPARg/f+SKZc
zoT44qIG+XRdiiKWQoXWzwrc8SVj3WjzNX7MKkj3buwmUpph2APpZ/CX0hspoEI7FMoCK7CyFRwz
FUI9ol3wTWE8iWesxAtzYnnnw/EfmJ0Ko7fzVZgRTqnRTtTH8kPld+nF8mh0rMv0axKzQKP4Uiup
tNLZo1hqcbS+HWpoylbKIWr0F+loARm9cTNzyJOlLJSWgeaVFoLckoaConmK+w8zIiv+fEBL2VoG
wcxGaHAfHbXoHA3hRxhrlzPV+Ch4kt3xidvhwuwrfkRZ9K5n6LCdYtzrwvqPtB0WZ1T63pR9Fv1b
UWIc1eR6xnl7ohTC8xdcDB7onyCFsgxdh3RzcB57tMqlK28L7hr+i8voQVxPDt7vHGuv4sQUTxh3
uX1KVAEMaDMx3Ju6sQUOsNx66/KzRYhHYqlVkU0IzCpD6pfAo4KOmkb6hwerQGMqEnuV39Kb5WsG
p1FGI3JPhXEQJ74VIYZ80oQ3DIbsRk0N7I9Z2Dz20CXtr3/UF/SMBMsBuRkcXZ5Njflekp/GByL8
uURSyXlFD1KSsBsWKCfOXNJVpFrqxgWbNzhdHO4BlriC30sWa8aCK2sTiTOpFRxzekk1ToKjpJ0x
IOoRZcik5s/Uj5OyFmjvz221D9bEkandfqEHc8EVqoKwoDUj3oBZbFhJsQNFyHG25iROV3vg6UCS
tliTzeftOaCF9rbfK4eF/fpykN57li7lHePIpaY1HRpmxZtXECFdybNLYC6pkB/bvy02gWEwVMsi
T9QxMBTsQ5tbIi8tu1OF9m37YBIW/YdQg+JSnT19CGjxY/6wcX1X3UBe7H5RuByZhKUn7fHaLrxM
wd3/p/9vnxtXKQVud6F+yXMQkHcRPnYKE54mdxudUDGLI/W5IyrWJz+ypPwP7jI/3ZuwisfePJzF
cVk2vcss05iNwWoxRdfCXrlLmqnLeHKWi93inlG/DMBdY1SFpsko5F3ujAidurOCGSTv69VIcWUD
rK3cLXso+xeGIIlnxHj7RW3JQIJFiERn0Bgc0j+Xm56175mNzBibrzGtrHsGtv0CeGVowfGXgfE2
MGU+XKaIxydNGE3+VxB7hiRhPpwCBXmpINn9rpXz0ayEQEE0nLSluOtXEhLQyECqwrx1ngnL8/rd
ZJb+g0Pn+4bl/eBRjAVE7HEXuYTgTDvLQiv3ymSD3DQQxS0y7DandNU5z2bE6GdRatuDADxaHWoc
WT2l5cNcvRjqqsTg/UUdpW6D8RVjtjapIQg/+2vxi3NjYcPdXi615kWqI1CLXbC49T4LHpjpppae
aFmljSEm7I0rVvCfmLB23J1dJRNGup/WPMm41N2lubtPxGyQWaUgX2akRQWHoBTJvA4IJb7R96iD
uURBYqOsZ/VDTDfrS1iKuYCHFLcPR+OrP/yykEPHSrrDiEY4yxLpHFhWwnRv/kO8c2oEdL6dp11A
uWiibwowgWO8ltAKybfUSmt6d85jIRIJ14LknfiD/HSZSm2TLMWI29CK9CDzgMK2nNlfGhCMPmlS
DTAfqo9VY/Caw2v2kzcre+qwOk3d61+Ctn2jwAP1yQYskfmW/a8wwnWSSAnH5ptw/7PWjB05ziKh
CwiF9Ki5/2eL/wAmFAIW/o8tFkhTvNG6PDEYPF4ov0J+mVWVQj2YfAYD4wVkwNju/CaqEnSlKGf2
zPdVG4uPt78rbTC0Kt6xN/sbG0fpKoCmL0JbWhQtD/O9gkWixK9dJTNz8X8gESCpYHrGrkuKE4XE
6In6vigmiUeJVRYupToHmh7or715baVxZS8W3loow92jlxyhopLxxogVaSQKFy/WTzPJiARGVzq2
0M6DnzziVqmV+wVw96wEDoRdzMplm1MktdjJXWs/lPHRYRswf7szGG+NL82h+u0CvuQ2JD6njisy
MUdaBzRes5zbpAwvraGm2fEks3RLT72XmliNBYyC4oajDt5GQuDSNLrAHx0SgqyDn4oo9gf8P2O/
6QeeMCUMoKvNHpmIPIXq99JvqSLtFl2Bs1UASLqotN6BObdwvEqqtpl5XkQTSHGlr9J1oeaUmSGs
mKgHycxlbf3cBWp1oyBtBri0JB+xFVU11buESq7PS/uHkWKxeACjeaU0AiajeLiGKB+qNmBTH8QM
6auacU7Q1XtMo/2Jz82av/Za7B8+BvLz7b1qh9lBG7k5cMHaDiAAPuwfRerb0vHAyH6TiwIhYnaW
yNH1ODhvVqj1YPqY6SMKmxT46m/fZOyMt1/10LEBc8OC1FolueOmY72jGuXez+XQAPxcAtlXOoXK
i/EsmkxyBUBD2Wx7RIqlsTbTnDgfWLXN2d3bq6ptNG9M2S5IkY3OoA0ubJxmuyOCWyWT/q+wo4YB
dioN0fEUkf8C5ohaSbK/nA61YSPQ6O1eEIbqEZSrYlvSncw27b77ixYrIDz44i01LZVvacDZGI4q
68oQlF+HJZs0P2qLJOwDWTe8z8Tbb8zSEwz9gKEFOfxTfVQgA2q7M1lx/aYn2x5882LVfSR6KAmX
KTIBHRkZxygsET4hzLb9Vb9DAcw5R2CsJa+DVYMlh/LcLyVgvTUko6kcUGVYAVW8C9tvqwkuXOPi
bULCF95RNOD4KlwC4bcOhupZ/McayNRYIW7SCeyiJDCjX1ANd9t4RvTqrq0fUembhAhCnSvp7258
0PFyYW40o2FEbszxzIpm4rtDgaNjfWWVeQxDSACIgFu9oQ11YVPkHJf6StmVbReEqzW1g28GB+gc
/IZLNYJMUn8iBsWuFF6ykQcrSRHXruTD9jGeX2Oa2elcBjaqshB/VeEM7iQAouWsayE9N3g8xss5
4OjjVe/7AOmLqrlYQuECmK/FWUq63XQckyWIP62N481zomL/yTEfUXl+sRr9eg6exzZZYMSotIuX
s8mTXXoeB4a2o51J3K4hbWVyit9rnSq1JoJKb6e9hxjJ9IuKG1KPdlIuJVHvwRaVjGUHhMPIp9Ay
SKtHbOl+QylKfHftMP23wZaUvMxvOrQMTT5mOOKAuim/i+s+yTX25gq4dNV95TSYo1aFnkqnX3GF
4JrK6HKg5xXZy6qOWFGzF6n9FWopKc7m+jvd2wQ8P0RfXMh7qERC/0JwcjGldzUUVVMRZ9bHYqsw
EUPBMetdTF//SZkzxob+qXtlWTp14Au8ImS/kS31kFPzEM2915LZD0ERrkO0Y/vrPH9YB0v6Nkqp
snIaKoJ/23PWWjVq67aKKn5MYQG55l5XofUKnmu1IhFks4g7PKcRumZfYiz56YsusI5IoDPYy1+f
6mRIGz9ljX5NGjZp+EHJtroCP4nDZk15E1pFz4Ujivg2CG4rpbXBco9JXqPhdeY+AtXSrQoAYLRO
/mBHJqIsj8+EbwuEFbLhbjXshrO5NDokCyGn5KlQY1XRtxROzGqIUp6zJJhkzQ75hybZ6F2YrqBc
IUvOaZ3k9Xe0xaSTK2Rh4l1gTA+bJ6ogq+7Sv/YVyWJRtqwzHdI1I9sHnjwmHKZWIdR05fBXbn13
PpJqeN9T5lR2I20fvyYiIWQ624dDEReDp9LC36MtxKnPDCe9AMwO4p3RUEgLi6o6+1L8En980Lnb
TE8Baw/oUmLd5QrkxDzmeeivKWe/dK4fj3rUqtyljvwkLf0oSODRYNn9XLlR85eoNUpJBrpHxXmL
alBTwrwgFgqxNKrWhNG4UJGZ1xN8HTZUrvcwEeiMF27w/7uZT/SaJpG8eC8I0GOUwUoIgpiu3xwi
5WYSPOaK0jdMt8/ElEa7Ocw/gzE/BVzShrTk+NjsfyjscUEeK4qHK+NqJGSqh4osrsmHtnqlsKbz
TKDNp2L7PDc/n1FrYdfnHAe2lTWBNaLRif720m7rrlHBUdnL7Fueru/s69gDiKHFGLFpCnwJ1/vz
HapVrmhMHzdUdRUBGfphM0jt248y4dEhdSeIcBHNG7jLFXMx7SZ7ocKCaZgJxPmJY2KpDc5Z3c4h
GxO/rUc0l2y250pSOpkpsbSdK0mW1mn/qRuD4mZJ1ELt5FDacCrnwg5jxJPcRlRllxKyHphIMUdA
1G1H5tMPlSByXMM1HIi3NKlSXuF5wHCdxF8f0yKnL/dMs0fFVCRX/YGwTFuFVoNZo6bl639rjUhS
BhIQowb1NMiWWydDugnbClMxjvZYnRp/6gsv+hbM4GwLODi9qbA12phS1BpJ8pf0m9fg/0kvrd4Y
nEECI+EMIk9+7X9bJjBwOWwl17h+shZtB3TRvG4K98aUSXMj0Lo5hfix52Nyt4XxPIodH/1PTuZi
wEM0IDNR1ZMC51t43RsnydOKQIae0QpWodz+kGvt3m0o+OkzC9r/YKSZEdJxGAMNTzfQHcY6DuSX
4MoD7sfC7rQ3mUNQdiZbjhlz4qGLLcr0O/7D3od+6Ea9x0eWuZrKILkQBPyvi4U9CG/qp0zbtDxF
01U7B4+z2VBKQNzE9OxcScaBOVYHksg6YzoNSlD7shNB44XF7R3OoM/VA6IfZxohHcjWxDTzxTgk
HygSBjOZQKkQRAwoORdc/sBeo7IGpaV4dtTuMESoqqtSEZwIKg6T1NrPnkDlNkheY4aJKKhTrtui
nrvdrqhtTu0yIAiwRf5QvBZSz6vN+zMWKfx1unu8U79l1tn+qJmBkM/jM8WzoVzGAAvucoZgKq1e
NkU6SWfy8csGW+qX5R3dnddnyMHtnKkmRcxn1oTXo4q6pWyHNyp2MBUSMMeSKon5XjgmObs0beDB
ymxf2TzpE9HeXSEbsHJPRNgLqgoQBRPnBLY6ZFItqQIgZ+Yx9m2TZQJo2bo8+6Gw30Ad4XW4yRZA
QNS2Mo3U8cf/+AF6lRROBy3jXvxpBlNrfYqXTVXuJ4NexbLTuvrRW3tKTRsX/ImUZqzstDjQyN3O
4HnFCHeQScAdQFWNc18GmXdXXKxOCARWc5S4OllYYj2qXpOO4mhBYhYkTjzvpyjV/Wgw8jZ2i5uB
+ZZ055OwhAMgNwdEvP+52VWwxLyVyzCniBtaFYR//ry/7z5ziDXZJCkvEJVMSCOTppuUgpM9UmnV
kocCEMnH0HvNrWdbnDdgsRvLFemLRR4pfDLYZrGDSQvB5fjeMlxixrU7dec7/MLk8uQdmFlZq6Yg
XOmfXrDCY1ByIkLfSyeiyBaYcqkhvWiZxl9wcZE+8c+khlddBhAzLsMVK36EAMpDZDNiWl/o+Ctd
/baEP3sWLXYRi5bSlEJe0AvsBX7zPPKFUCAXrQ6mjIkBs3ISoPD+wrRo6o0te9pfvasxUAO75p63
WNM5N2BM5tGEIe7plAbii11oDmN0L/hQSgXU512yv+wdSTDDkZhFyFx3MGr9gjYXdDHOJb5Qn6Pu
01OR7YpjCKAZcsi9huYHbx/y9JoVohiMzLg/zouTervX6XKBo4lQ8wiYLc0J3OyYhgBaIy34GDpo
UO5Wx6KztWmqsgIxle1ntuYIo71yuANNf9MXdko5UieMVHgxkvEElJx2EeZAFzWGcX1hbi2IB6xJ
hnmoGHbslxFe3wry5zulAsGZp1cp4NA41PyxJy4gGELPN4+z/CYiU17QGBebahyGMxwCR0GnxTAV
i9l3vEVdcVvBVmWsLoc2XMXXM8zHUapGIvB7AAZBrneAOfO1agK0imTsGWBxkr9gO6/DQfRKHFkl
8WFOhLRAM8OxR9NiL79eLtJ0KVAuhmYubRzZUIK3YSvPtSPwd4or4VvOvXj5Isndj+oTPhKr1izB
r9infUOZdz7dfCPgAcQtEwYQfBkczyTSnsgGFhe3Zxwdh8DwAWEBbyeOH5/9547pAJmPqKGQ2Epz
WPGQrkPq2RPALSYZ7ofYGWEcMZptjLppNwZXQcZ9+eFduX3QwO+JbTSc2jMICKZ+Bn//evnMyc57
96r22zYssxRRLynwzLtaT9VzdtJtUxjus8ool7YbTBJQYSaL3pvP/YZfoZ2L5WnEFJs08E4uuO4/
HE8bu81diG6cXViqrnrv5gYm0Xb7OD5OgBCWrVvCcep+ypAAnN7/CL1/60e/6IUuxgq2Mh9Q91Lz
VVZ3NMQCq3r1S8NxLyAi4JczIDKlxHjknxo3tuO7L2JVQp7oLnOdujdmxk6KKNSVePyYxJ5HQlHm
OmtvCwEjeMvjgR9c3to9Wa6Y4A4iKdYuYEaEpsWGBtVPlrFuhgmS2y3jHvm5PQQ2toUwWmxKDt92
9Vky03ZVkL6zQID6h7QnW06gDPgF0cqmMmvKEugXRJbS0K+s5Xauqr/+XMR3wcAj0s8tBOyeoSMm
QvkHFgzzh74vRMTM2W38FIy7SzLZXbhoJZI4v/JZcmdrjRMuYSuy6jw0T6q3DZ3WpgD2kAKrdxKS
MnTt6YV/KMPTceV097z6BCTzaYafzaC4H6bcRujva2vkW6cc7ume2qgRgO6ODAtrCeoNupNSpln1
dsIQWXWRWVFqcKZeZg8yDg6e31mHQg5cloZI608xCTjlvAtlC3V2su8w1nKDKVgOgUowBBppOFnd
BpySYjob9696xreL1MT5U/x2SDzJDjcChBDN5whWgYu3u6G9hj0fIjFP6rSbcnts2VLimtGod+A2
wFXohcO8wqGWwv/7vrp5KvAkMHN/5paOVMz5wJSOh12Sa3AG1/Lm/8CumyJo4zGc/sgXEJwahaSm
tmdh25z9yoeeGAs8D+ULD+ZSzuxWRacrWLGedIRkWxijuf4ZLq0m6C0WHCS9LWBCVWiIBnhwkMjz
BYjfm1PFZQDCtt5WcySAbK3+2kM+rwj+xOsi/AKZNkgOrGO3UslVFO+E7Mb/5l3l66fk6wKhK6sz
vZo2az988xTeOa6FwRDCftWXzfItXwj1JmRRBrEohpvL6zq7k32mdY8nBv6eWq1zAQhwMW59Ruk+
qYKN7H3oe7MofiBYkXxQs3ZnXxErZQMZJeZ5O0vP+tYTW7ExdqqGGEWYL+ZpKbGr2YovC/xdGhQ+
+iKMKmDqOtoZmlLynhfSTWmSMgSlBbUUVwrwFYDW3I5iWQuVZsGXdzCz9roOJHludfV6GE4BUMEb
9Gh+E91DZXHKP3IWGyp8QmWRmcaDXbPvzrbco+lbPC3gekds8ugrr3U5Md1j15X3T2zH8cgGXeG8
D/zIzswhFoVXQ7kuEI0Ne58EiqGs4mE63shvzc5RZnfyqzIO9qy7nUnYsUx4Ko1MIb4A88vg0ACF
glQe9WQQuJ0sPsczh87K9MQPozCvPqQnGq+8Twl+3PEgGoC3PVhpQ2z4RIci3pocz1mCmvIJcKDr
E92Y7M5z7fSqTBJwvuymfp3gd1EraH5xTPwkIWoJuIbCqKV44hDssEuSz5pp0Ngf2GqsyZRUmFDU
gLMj0ajxTvc1CxuXd7PmTPsseqweFoQmuiFWCoFWO3JMV1Q3grSCyjn0m7B3Gv2jRp1//BxIGGMl
JsN+Ugg0Tpd/ABPtAfxVDXMEKg9M8GjMuDmFEO7Ia6ZS95gJs0Q7k2ND/EGO7tTujAA014uPtYSE
siZ8FF0WQu5zzcpnNCfbct7mzZluEHMJqSYEhCAWXCMJRvGY1NfC3Y2TpK8KTzy5wTHhrj/sNG8d
kuT1aCs+2+7F7oteqzaYWd8GNY9t4pP+82B3ye8qCmEZQMEb40hAEwR/rFAsU2MKEYohvFmWE4YN
3MR8LmE/05ar0bI7xtmKh2ZHkQr5f3VauYYql+HwiJJbQDCZrC9oqAMkTZQpN4QGgdcLoo1oY6Ew
e5nkcBu8HPnIDSwtMbxzcUxR8yihprH9yJb8Xc4CB1jYYppZraJ/va04n241yCNAv70AodmxRkzO
6+gJjSxdw/a7SpffuQ0hCf5Lm2ckNfHPkkkKVOCONo/o921qwUAE6iiLZnhb0DBgt9GZVT4J0/q9
S823RK+YvwlRB4nZ2Cjx0jxoAJ8m7Yw50QjfZXW588EbIcZq4NFjBCx8Md7VuTgIdka8pazfoWdY
EZnN5Aq8TYRXsuuk822E2mCJ9SBIO2s3oPBW5bOf3vj3u7spN50KU3SQH6lZkKEbPtCCOZEvLKje
+fMRVRY5r/3tum76mPHcoK+l1nVKcnXT+1QPnQEafil+BKT5i2JLko3OlxI2KzaGg7G9B9Gu209E
xUVhK/82YcOw96TkaG/QZ04lwRt79vZnDEIkE0kEGE0On5R3J5kI4zAPtVxLrTKPWOU7cIAa/+ye
Uodg7ziiRFxjmJM1c9QJ9RaBcfC4tzv+vvlKj9UNgMVq1YEf3kDLZm4Z0NDzBCeC+Zyjds15E8+u
b9meT8kX6jcoVVDWTorE7+QGj0Kvs8rgljktaR0BBS/moy8Tn7umtLBJ9iYaAS9zX6+HbTmuhPpK
QGTCt1r1M96Y7jcFQtXGAhbOY3MUAylsYn2dkpG0SmzoRpOfnGJyMU2Dl2FbeWt8CY+zh0dnD9a2
dD8niiqs/RwHKJ/CUW9WGKdkw+//XX1hicEOpOS9ckdYkr/xKJLtKl6Zb/J9D6/1NCt2WM1zLZKG
N3HOUjmzeNDXTKV+5pSUPNNWaFct+CPmwo8MlKiPJ3pHySoCApZOyRrSMpy2RE1xxy1vVq7SPxUd
Sa1UGLMYV8dGAULJSSslf5CKxGdPVSNFHodSMFwoCUob88hF58nLdLLXIO1hqBecshiR0K2Zg45d
71CsRmTvXXs1XtSM7Q9uCoZWtgwaX8P5pZZN73So4+zYVaEws7RR3eNreNOZ+xs1MpwuyRktQ3Ok
ShYVGblDbR3uCWre6snMvPsFrFbzD966RRNs+dW7hOJLGQ9CXkIPm9I+kRxRtTeNi8VmtbyDNV4t
8xJinKKKQZQ24kbF0FGMrveOreq6LlZmtnTqgQZWlzpLXON/hqyK46vpe3xYvnyIUkgq0c1DDYum
HHTa1TYiNAvei0veBwJ0DnkR46/F35XI9nmjAWHJeg9j6rfxbmyjQAXGbFHchaM1KSNDWc31QMYA
GnA3ksYIn/d7A/IDXpNwHNQzW+yJgtoGpndUvTaGe6wST5ReU/Ksond8g6LpYQlC8jtq57fvGCzR
p4gA4RAlf7gtq3CpoL/qZPv6mVcGfXt+eb8AKX3Ddr7NyD/82osHyI3XsfXE3gnOcz8OGysTYuFc
aCoELy+XB1fi+ywxI28TFhUSSeQDwj5l1SQnibsOKadXe0aHnmpyyFREBlfBSTjvr8JxrVLwSde7
zkaEnCXfVusop+k36bSbCIOnz7wQHAiISF5vLwxPgSUchByyoqTKd1ik0eyPMC0sSE+PFiHZunCj
nwpr4VZ3VkvjeBLilW0XiPUF6VMswBUk1GZ+RNEWP/+B4bspx5wsdWLfgoR76VZienXfvPjIgBO2
hfM9KCJOiNl6/h49pZR7VRlS2eQXctBwyxzecxk6S9CJ9yYOlfSsMx2tej25Sh4M3fzCV9iQT9g/
/3EdgVlq1wEmEW7uC6A0cn4z7ROZKlAD+BaSUAehedGEpRiEcnwWqrjiLoOh6DlMrj9xAmAYk5jk
7ESZ/vS9U1aFdLNb/avS7xs9bl9wNfrgalR/2qvKlEGPPFjDREiRXDdGedqKxMCewDmvLlG/BFnF
7jJuxC4PC5j0r603qx+7c4Bf64OIDZXR8wgKsFbPhJWrmC85b9UyQJtk9KTMSVLWBStGk8T7TLnL
SXrOWBvwO/PD9QkGimZldiIOX89mEO+jrx1OJPSJAZHQZLaMwgaSnCqEBBLSpBrK7iGa0GUu1s3C
Lw8wx8IW0ywqG9pHcm73+9ZFaxHNW6Hl1BdLC3B+sVsUsPWNHh9k9oce8P+rMOl1F8zs6eoYc09z
ryD6HzwOVv/YorkePGDnvo9HIKd8QGGmpWjtWNqpwW/a8GFR+j0Ab5bMUxXln8iLKJYZ6fCAiKgz
J0rlPUoesU737j3U082QSVs2LUsgwts0T9qYl7RM/kfGzjPs7mF8F3coL+mz1ZOsxYxa3ZYKvIKe
7BeROvpXDET2ptW8hogzzVfczO9u2n5VpGAEfuO4QJQ1UMiIN+9N9C1NCCoN7AT7m2d70ECPtooI
Jd82sqw0u4l2GtiDGAUjwcegLU5TzBmbLH1Kz4ZxjsDGsADcqO8PL5Au81H9HvOMS4ipUuc4DunC
w6zedwshXiJOQ6lEvFI6yfDWdc4ljP/cDXU24CP1Tg8ewineqP1s5IcXZaUmpt42+BXcr/iPtv0Y
w/7KD/ehHmks7+HuIlVQaDHFEOUMAPvHrHlZS18QDJ6j6AC4CNQdgYSEe5x3lDM9qS0XYuD4lWk/
Lsl0ZgFxRZZsIr1vH6Y+gaho/kIgc6vuHr0b8+aN2QUOvj0t5uO600fQ6U3oXWqzyIDI0NKNjF+W
ukN0fVnIxEbjimt+POSK1eCcmmOhkEtrqoXj/yK9XCK8P5nwSOE3+yRgFN2vwcc6cLX7Vzwlh2lH
hP9huLGSRNwZ950IuKGB3A3wzCgekjsN4CzREeyTg+98RmJCeT0jQPxINq8iDXOKv7qk/bp+NJdC
XsVd2V7zAutaVfRpZqHWY7r5b9NnaDpsIUESarggKN2fzVGH2zvLFgIgS86vXe/gp1F7nu+6ZTRc
bS2jAGUVtIyRuPR0Iz4pqEwIkzl3XvmKBEbIH1RrK5x80DgZSTtE/oyg8eyEmUV8BYBAQTC9Eh3L
vKLnoildcvu+8JiiH+qSNuUml4TvU1r3qF3Or7NKe/J51xz6ZaMZ8Db0B9N4t1lJe4s/vg4dIZZq
hhbVSA67Y40MUpGPe0wfNx703ujm0BrBjdM2QKCxcYE8XAKyN4dSReeYaUEPdpvw47vbNjpdP2bn
akYDxMN+TBmP6dL/nyt1zXHB7+0debHPRugp7Ks0/3sz2Lu6FzYhzgcA8GIhKVv0R5VTgJP14vS4
YujsP3vDLpEUqN/4Z2xnstS7yXF+kcQPCMF8TWZc93qfh+JZBGxC+kkEgELcTqNKMERjng7bEF5u
7amF15KP4xKHBzmT+NV8UoAAbTICay7ZsGZvKtieWWVsaDcPCvX2Ow1QNnrU+F/YtyV1kTjPnLtA
XzyE11jshtVQLSYJmqZphiiuhRE3KQQtAn5ny78RTGGhUvpeBAKwpE2Dh5unAN970GF2bwMenzmu
N5iuyXII2Ql8oGH/TKB4Md1Z4aWSqVhSdmw2pfC+G76sJBfLXs928CzzkgRJH94PKutX1iq9VWqX
Sfw2VuwWytlYFfSbD6JrlZyqeoJMMEa17wBvcLtKqdKSdsq+IbIWJoeRCHM9L4fq6EmeKroIeS9s
UUVvXW3h8kCbjoheDw16ZuzmhJMHkkL4OfCfGi+6A13rNqhyXLol/DTY4JORZxo7/czs+VbYFOor
dPb4n6FmCsE5T3rNwywCOSgCokv7RZ+1zaJIgvDnag7fY2gKJInNTVhUAhCVwUBZ6NwCjei+/lvk
nMwFAliU4OhUbibA1pbfXmUcemAjSwQO7DZU/QFXtjWIbJMpQzdXbPuJee7s1dDU3N5KvIbSSvmQ
PuMT1j/wTHudic5rf8thv0vUx9I0uKACT0PYEg/yieJripOOyvVz2N6HMLTHmTGscvbS2O0cL/x0
y+36g3yaFUsTHv7rsk8KBeRh3BNPPa7JgEsaGOfqiemJoiyH41cz3OW/ZzxLmQcnUU+g70ib1ggC
5utJM490R5f+PsQSP485LNRHukwn3PNKcIOTJ7lqn/ifL9liNsgoEERfWq5azn/geB+bfdXwc4sr
eR8hLjQe6/K17VonJ69xe02giFortHWQ4ODu6ZyDj9QHEpT/sP06mnOAqwaPAIYJMOsivMhky7sk
pzlAZrFrwVtdgx7M1eeSg6tUnY8YAzsoNRmnh7y5tyA2brPNGT1mSvveLk1l+fJqXt7T88kmVRA6
LnmtbkbTikglcJ8JJvyDhYO0qqRYuWtIe+BLxzqqV0fq5s6ia6tmPhJrAFbZYtf246BESfUO8iMF
6wOEYB4VWmNkBAHlD/ll2xLS9P8SKkughURG7U+L9E42ZIfTPdoKdMl/7PNivnD2jksn4ORTE3xh
IbYoEZ9U21SlrQBZ4xwPLONBWQAS+XvJHLaZCqW79e0mQRsrJyYFrQaQcT7eMQAZxG3xb02izCRm
8TLuX5cmwfTt+Oma8sTiWHm/4BWP0+JMEwZkP89KMa1+OnpeIuomJ1CWL7FtguaHOw0caY+7WV6N
5jn7HwZd6GGhO1g9nJnJopWAuy+PRyvcBLUaG9syRDiyIAVi+RGF7H/kIvMCp+P6XGtRJr0R2jzm
VnVwU5dzwLnxMyebuYprgFrkzTpH9Evv55y6SHPDOjjf1As2lNJ4yy18YiQwISKjzpVzNYGR21ee
EfUA81T1ytbCMMPAbvt+AxK2NP5hBMx1hC7Q9Fqtp80D/M4Jrgyo/hwdrHdm04X0N3q2RO1cRd6Q
K0D0TSFpR4BvUK2gxg6Cg5uEe6TPwixXG0JzwzP02wawAnqDpKHG+OUIBLj+9kytf40RsG1wPf8+
LcgzF0F2QxrFMmeEMHjC9Zgp8yAheVhQYhiP+xFMEnd4wHK+quPWRFgHInSD2uRVjtmMoZjCNwhu
nXFitdgGd8H1YXsOmGI/liKU24McHOBducWLECmvy7UjUys4a4N59YZ0a97wiJN1APYxWBH0n67Y
KfyxgCTKncCH4MWHeHiIrd/NQTUX2ttKN8tzqMM++MsugEzIrvm/Bl37PA2he59T2uzBSi4DKAKI
dQGxkvnkaX02sFR7UmUGGpJRVOwzBxYYU62rvuNGO1+DSjsNGUkoPN7pxsi6jD3kXv8C5CqEt/pO
Z8ptQySUNfhVpkHBKKueFNs9dppQReO8hoClJnfPrZElAqocBcIVI6i1dkxX3ivDMOd17Z9L3EWP
AY9KQ+YPCP3NyqPDaB67J3smx0w1DwrimVeiK7CP9+6qMq0z9UOzeYFTTzZdddhnoXU5bpkyriJz
WE/o9zKOXucJ+1DGNc3Z1iN8WqugTurETwO+dE/1j9yMQ0IWKzbwWGxwWix7OB67uccLiGNehwAI
zEvdLdaM7LN+M3OqZbBWQPwWHERt5mQWzeY74IpxUk557AJPZo098H+oXXlIFazOagyqtoqJwAqW
sgWxebQv4DVwmt5OTQKDN8fr2+scGs795+2ID3ld5MI36rQQ3AjBSRZ0vlQ/37p/I9LOG07lr3ZD
9wRi8H7nRnOeXark0IFDstPOr4kY8Y/+9i19Dif0VIekiqU7o3rJ8r95BtBNaP2HaFnNBQ5YpFVC
jWveFRAQlhPzqUgPI6oJvuu4yeIv2XLPLm6z/+/M9XW7cZmj7OJSiPJk16e7m4rJ0O7qu+ExuiCC
NWgksWLzNJDXAIaFDFWqDMXQRrr+PBDoPL7I3mw9j0gGC02h/IS0V/XbR4Oahn/GENdx75E4U2bh
YcQqmfGov8z3PTt40g8UnPi/ukm8YIM8fbFjIEuWMD2AEhYgdzMoDk0I2e7lTildf1MhHzU43iua
HwHAY2WLr3HLm27xMx4DDuuxfA4y+OO/HCa5cNbq0PTTGtwwyeYyBclom2KUfOvQgr+x4+VhR89/
XjHbv7dZ3mVO+Z/LLqoLmCaZdx284joMFFLMt2ClM3Tn3xRhEALQLYVEZktl8eVXVcORSqcBxClM
93qADnLB340Y+tQADErfmsHwl6Y+gr6Yx+/I6mTnUqUcCgXFa80FQOIJMuPbEoExwn2Ft6rcsQ3O
in7tTDH/uQHCarn+JLo6gpzzwOk5poJWTRrVvh0WLyj4SbI0pbmZPMcHJiqqDh+ZBDWU+yiqghu6
VEBxdAwAUjp7N2ImpwilMUkiw+2OxfTk1FmF4dHKudfETpjoDikCsoNs0/TlcqjfuXxRnyLaj5p6
qi3f84kiYvkRr9hVxSthkT30+dONT9Rj16Jo9Rv1WnMLrd8+q9qNDyTRlUE/9L8muuYruuc5Fu2A
4JgGIbFJPNPg4dkr8gxasilG6U17vEh++PS1ZVOLkRlTSEUl2sSxf2jp5i1H5wzxF/gOHagDuYb+
R9JrxNCBR6Bh2ZK+t4+KM3teBULi9K57OA3SI7TjDRyiKaY2h3EQRsyVpx0sTAky05Yj3dbut5X0
C4THaID4eL124JRB6eqMJbNxGLGE8G262NbEFSqZTJW1Q35+ZXllid/oCFSwXWPkiBVXOMy0Arz1
8YgxCkx/KlT4EiObElA9oRsGsKN1LLM2nIIfjhl/xoF+ooyrfxcLfJZoXKO0FWgweJZORM+heDmS
ul/vZDDhIIfXK8BB45Lk7OoDR/JLERpntQHgyJbQFpe3DBN9UrGvD7pzuvfEBYN4JrtgOKjPuQ0S
3c6tUQ2q+Z06SY6dRfpktgcpbg/FIbwexkUyXYKkDB5uU6bN1gcUII8iYLogQ0yDsdVOmpgUJovP
D0/+vZ1Vdr6Satt0qTdpKGEwyWvT4o1DeMZcsKzOgsv+t/IhPjVRpWwIuHSr1pY3+ytVzPDMo9qM
F6TRyrOaOkwiFgm0zBhvljy5Vqde6ShE4zTtf7LOxOeK7T9iP6cfn+BSVaPBVzry6V7e/M0E/8G3
ZrYpa6/3WbHoSR1EbbHRBqn02uzWk8vWnRCWyMwIdvckGoyGU+KqroOCH8HknFqggi9UPAj023eF
nSOVWHi5DOoPEcfbwbZHnul8dPsACGTf8vThilLhVyRaxNCweJZ+C7AacyR+N9e6HuutxtVv/eZE
vyhEPLovhwvjtVAvyb02ugq7uQ56bxaNs+zRsDEifTymHEXCgwkJcjiQ/kfZp7gce/WUZjMqUrxf
cWEAm/JBfWZTDIPDTghs7GTn2XjM0zX47QJ1GXcuNiVZbr6S7hi6pPAFkwvGrUhSRJDPH6bzPwZ6
a7lLIoGnen/HGvv76Bz57HXkMFGW0wVax1vMjGHfu6gTI/bhSBWkVg+WYa0iExSm9Qdb4dC41w3D
UJAU+ZjhdcJabnmkxzmWFSjioZgnLPujgxP4rUTNObZPey94B+gmIxU3Sf/yequ2PRkOTad2k0JQ
pDhSjBaGLNf+nNFfKZHUSqHPvVF55tezcGMSe6DuAtSRZMxnppLbJPuKXD4juYaP0GzuvvbXb6kI
WQXBZvISfAjaBG+CZpLxiiQZDic8kkn92RwXx+7y25Hz7GVofDZ85yaRHLVEkqNDueLNsweU5x6U
zB9Ns0H5c149jcWucIweAEonGfCINerKQMSRW3UGouEdmuPPSb3qP6UC83Ct/a2TzR7xVfU0NbCa
08/36HuZ+bLvo61HgIjK2HGQuF22hQO4RGamf0G5qGCYXK2FsclVdtxAObSinLf8YunDCWzpFD+E
yeK8W86Mopbk8Ln4RZM2mgDxqiyH2mFcJSnV/4sH2rEoQ8t/wnJPkmztmWxhx2JAWrG6+Qb2YaoR
sQUkVGfIVMJFzjQd9GIQFdehihn99/y1v1AH9XctGwmQbngNMf4wzP049xpG1EGh64Y6v9Lq2GHP
0Co5QXm4crG/bEF5Lw0/7w4od4r8pgbZBdgwGPsmjdgFKJf3OpKNjAwmAiXFxKBX4GTVXXE6T4ee
QT7OISUFO00am0OKk4n9IUXEMStma1gBEjx2SPpVQi18ikEfX6GJwBj4lloQ+2JJ0/hTz268B35c
mGruqz49BVLtV/1rzkFb8JCymRwhtrIJJrDS7Knrvsv6T6Lp+jWhFuaIoKoZhuUMlDbL7Rv8ofKC
P1S4pgjcw1Yj1+fKzTRg+yavQFWf1l75pth/+B8inZjxMSMi54a8sxeVPCH1907xKd3pYUq3H2rh
QiHfqX4uNipoN5x/lXZXwwFDUmqWD18mqhOuir3JRqE3FJmzX0FiJWm1X4Y6W3nOdJD2CGotgf6I
vylUN1GOUpmVHaxFdOZZI4dhfogLl9Mi8dEeT9AKgfGZShg0+fKztoggxqUterXGiUhloHfGpr9+
U2cRbvfhquaan3VrQBAcvkT+evrhjvBjnQYSmVgRbgOE3g79K4XkmNQEF/dbcnFvAO9LrjLzC17F
MqAniLemIS8IeKSCEDA/6cfLineQdrqRIupeYDhWkqym91G4CkqBx5wP8W2CwJNkhCulK4sylHy6
UjaKD2qJ205ot343NUYpg4Jk9wJjr59LaInd+hO5jsKTj+qJE3hhayqT5LZjHEXuoXGLG9E9zjzx
yLQWoZKNdkmOB5HxO3vqcskcDjFFqP+ulVEC7jvjwArNKrKI9tO2pbqpFb1ViaYFddYZO91s+UJj
A5ol6zvjNg92Eas4w9mATOCHVRHMIKm4cc2CIZi3SOebkQl+GGdKGpIFV45JJu6EFujhVSY66G8T
DSHd/VyidpYgFQLhot8sin/J2EFvrLCsKGoUSIWLRoUWr8dss6jMEVit1CtIUhKBWAswjjuhd/qC
THOZ08u6L3uURRlEh41e1o1gQxCJa8LQNpFtPvJvvUjhEDxu+E53Q93RI853nKIkvGB/RfO1/+Hb
tDvPPVdyx1PpBmIGv21mBsAUQWqrycdPGrowigsuYgfRI2KySJgG3dKKbuhV6HA/5F2SFmIbG8aX
FvgrCaxvMuhM18M9kXb1yqJ9YS09SMPzaE0Aj+bIDwo8q3k9rJeExOkFOCjaBzLkoJ+Td1Oo2rLq
1R3KEmlxzqy8S2wv/laY1vClYBYA5glwieiElmn3oI7C34dYsm9Jqs8AoL79wrce07HC+Y8FdqUz
WY/3RPb/KnKtDOa3Vh1PbaosXxsIq0qokVEg8tugDbfbe6rrqnCImuu0JhC87W+qZEi3fVPNxGcO
OZ7fNjau5QXzJr6rOLv/P9+BdUs2nPbcs6NJxoIKCph9uMuolk+9hXn56D32ZVLMV9E4O8xjVH+9
J9ga1zlXkcTMtSlc4s+AJzcNQ5Q04J06CcVTqOc7wNjgGVOCA+YCRgnrPf18jMhQp/s9IEkJzl1r
Jjp8y11wVPSxERZ+xkLclylbHEirU9WBkzTTU5Dzfa+JXxKBQFNfzbMTM1DktBEiG91nr/tcH1eR
2/ESk8+RH9Rs3aXIjMmRzaJqDT/AstIgEunl95ARQTwcD0S6WlgIPkoLZrungqoObC4zDjv6NC13
7pcmA9JU5E7i1osb7BYXM2N9RCqzUo6+JgmnR75Y01TLdGoWR19wCH4zkavK1AZi07Eo7LoLweyv
Xw4324/0MmtEVLZiYmYRZY2JqBw/uzOHMKarxJmxljLRo7t+KWZTq3PT2djmA41J60h4TrfV2ER8
d6lo3GxP50jFQoJKvMaNCrL2t4wxdwx3HzhXnK7cvU2cKjwXAaMybfZR2i1h7ge7v8tL64jLxdjH
S590rjWlt+8YVlksbdAwa6Ay9NVXhdvqFw62z+PHegpHLLkguzcwyIR+vGS4rjOylXKyklhbBgva
hp/AzGs2m9b6rKE82ngvUvxk/NYeND1h4DqxCbcX9uYhOifhxI6+hZUKp7P5nZn+DQX/6Qxx13GQ
BDQMGGp7kOQY/QfETto4EMaLhdx7OXKwaaL6qDcuTJKtRgFrUTDlL40LWv4Z+hQdrAcWQAbX8eqj
Cd0vh9h3GG8IgiZ0ecasv+GF4WGO9wHn5vzmy7IjGTPeeYFPNhAIIaJNmS2tgg85AelWPVnuzt2d
I6hTIxcqPnR8Xv0TZQhbCuQPWDEFT9J6ei6VYzWJ2qx/VqLdCPp4FWEdu1HzQot5mTStFT1w1Par
VWku6IB7vejN6sHv+hqU1MC1Wx7KGGBm83BPSzb/X/rzroEEhHGp4S16a1Rx3V6gy+LilEg7xcO3
963fKknlyhMyGyCglUePN6NhWkhetB33xwr89NOyuy6p0H1RJEqBSCED0D6uUWUF8NQieXwt8mGL
OymnbuMGJbAN9bK9AXDR6bT9HPuZ1KMFaeOhiPtewMR+FvnOjX6eDoUu+4f3ArG2F88wZhzM2ZcZ
JguC8RJd9YNyDSWZU9ydp+VoQh7B3rO7W+Xa/6CFt7RuBi0rKc78Y9hpbDoQh0QWYUQrypH6bWeo
VLuuJUKgXMUmcbm98RCwZ9o7VFrlLkoT2tFT3JkPkihcd25HM7jVUIrksjUW02ilfTAP4ZOCnCxS
s+yynzQ3VG+TyB0Al8vfMw6/nWfHPWjwxnwvDj7LlvMkd0zNKT1yoomILF0a1OGB5Hx19x4o/W7v
JoFI6NwNgi9GF3jk921TLJ4WlZw3XD/gjo+Zu2GhqmS0PIo0Gz1nBS7qbYOZS4AHSCIVWFVCmTUs
GwHn9/MF9LwauPcpTpGkwxhmyu6uOlPeJmTBhT7SxGAhvwp38dU119erB7w2AM4KVIAESFzrw9j+
Eb9MpvKmAIAN+3iXJFxFWLcnyA+1ztn7+vy2Ls9DPwvsXBt5FyWk/IVpxO/nkjiv9bkAZtj9uihV
pG5AygrJW9l/lCGbC+x26xcEkDox/Rr00wqOZ2xk+6hEc7VQAhwknP2AbaSgwuOjJ3ThmPXv6yIS
m0anxtBuOSRHAe8M1jj02t8yW72UMs1MLPAJAWuX9h6rCt//wfJ4dxFjT7SimJMefD791Pk5+5Zp
kP+InXop8Bf+X1IcZJFSkt+PD9tV+yXHM6oXKz40R/u4LZ+h6rC/PT3CaTtKcUoFo7DGG9wVfKQv
nlzhLdYJ5zgK5pPsQoljI+9FeQjI0hcIssg87X7hhWfcVH2RT90QHSEd8CNLxPkBAR+ONxOdzXJJ
Gp8JtDYLnRhAh693ySNjsiY0G9fD1DR91PIv/AC7IgGsNnWlc9dXSBJGEUlbPjDqQiaaoQYHkX+T
8cRgzGgcif1JzLHrgNHcJ7L+Vi1Xvs0IRj7Y2O3uOheg419OYoPrnDCdg7b9puMLB41hooVoXLl8
Ws5gnNBABsco8wxD7LbVKEnZvKsvY6K1n/q6fnPXVx+1KKzXpvIGQ00yQ2VlJnN5qeRR0BNR6D03
TbRyiHIZ5sWmmFXgRTvDSTcKq4k+8qpQ7tJZJHGJ7XobVRw3q6x3GjfOtb0BhguawM7kLx/K77bT
hvq9dkefoWECyywzji70L49AANxbnUdI5QJw6HLFnSgWnfhZHac0gY5nDMXGLjrc5k0ZHwrgAIHj
uZ0Y1G08xoQK/4JxMy/ii7kROwld9r5pUzOlTdJfVoWy4riQ3+lYOo5mlgBNH0qw1bNSOu6gIcif
FgvtsflLcT9atUsXab46Ft0zxHBlhvypMSWgHKvLqo0NGAHqUvoV9wGs8zGGgimqMIj17O1nw/84
LdSXmo9JvvkXRhDJkXAwgg4WIDnKof0JmEcSQSzsUmIg/vYR5iUESDbvlXDq1HSRfkSF3JcUR2Wm
YyrGR+N7CSNdKc6ZVzM/SpKgYYGKtncc4JF0z/9yr0WgPpCHAGPp7TtbnKdf75+LqCymvXHkjEkS
lemCGINLtloT2pxaaaLw/ujKK1XAUziAH7WsEisBjmJFaC40XQE7cJEvvttslJk3XRwQEHR1vvvd
FAEpBOp1bsNkQzRVF6dRoQ6lTvKKwz+3ziOSWvKIZKPBBVLPVvsu8q8hU8PNgD8LifH8MvWbpGDC
FZe7uwQCAnYdHuU7nMh7vAh5yL01ULx2bSYzaoysfPil9r9vHXTPAuDZFpBjJ2A9oIXGntn8wqUn
ycz3y4lIwpVMdD8TxqsNfRMSNYjSiG4p5dRDIHxbs7nXzxQqqC+AxlM4Me2Ce/XsXzR6JNQQocDR
5amOCSJ+aX9FzeMhMNAFp15W26GafGAf97VZE0N2xPcGhMrEtNwE/qx+UwgimBzHt/Dlv/rwEHq7
ITFLD82WF3Ctsox2C5IZVn6C7ytdnij0yqsWdYRQ0zavh+iheRAG9o+LPZubHyib9X1M2JqWXnqb
CqUU8TqD79OUu/VX6vhuVYtBrfVPOpUObPH8H5lmLVxqZFX9eQ+cN9ldodcjLqQTluxmoJYB6c8/
zYtajU6lSINsNnXD8bzSD3Ru5U5TwlwQazDaXy/vEZmXH97xKxKolRbHh3Gfasczw88Nz/XMWEay
WmHci/KXAEga4VVvtS7pCklV2FUauFeSAr0dEtyikYNGuZ9MLDl7XvdFNTBQUHBdmmAixJsqDGna
pQV+rFfjNFre7IPyFgvcJ4Aaa1yg1lCoDpSJWVdBAdrgxPiLRj3YKDa5gsKReXBJ05DS5BsOdnyf
pVQbzyjIfHp/6o0zkMVUt68UJ2gn/lQVGDyt96FNoiWzdKiy+0IInOcl88r8tj8TTX0XIdueDbBo
OER+dDM7J149l7wlL6D2ftJYLLrY0nDsI0MeaS7fnWBWniygTrosDpeWVUp8HgLgMPcNTSal3nIa
Mu+b2dwqkCGzPbW1MVPJrGcaQ5fNk/gHyQGBNkL0y47llLklYcUr3qe7I0up+TPDFYpgRxyIGnXn
S8utUjwFDJDverJlpbmt9f7X4EyUWLU3xUqjr+B2Gp4xGivFa9jXwVpSHuVaqJ8yDmm8DcUc/rCn
4lZXe4V5Bqx8nh4HrhoDfpoeKNe7WzdbghOTqcSM3dRRX3bQZ34c0UsQRff3741aiNy8JwuVTLcl
vuDb4tW8iQTJZ/QqUO6KKdNP+WlBNxaboz/AEvEDEqqaAhvEqJj8JZnAiaoRLewJJ9z7SJVSAtH1
USGppxXWpWuB/L5osp2g9w7rZjzOlZohxxLqu2bqLA+WR13RevMht/u+wPuWZYNf5WlE/N3oldEN
mcfeh9hSsLXoJL7wYsEw1ja66ZSYqnUBtQruqj8M0OLaXYRbYs04bz2u06vH0CsrCbX6W8jwWxUI
yor+9rJS5TmMpijbZjUFMQq263jhwtFDf1OufUGWzvNoXUsbFsj9hR1xs/peC3cAUkqShCLTCHvr
SguSLfm512j+vuG7D7qoSoOKjyrW3Adc0x1b3n/eDVSiv0YoX05N75H0rVNkadGz7QdJQnt3MS+q
SZTGHEi0PlPt0JUELYgLC1Syjvshfh8ayYNogPp9IdYq3YpRzUxGBGZlM5e6B53sJvz6PGkdMuEd
a7qHNozO4z67qsUICiOvk/EpjygV3Xf80bBgPCDm6AeUVrgJrKEeTPQ2E1tDTu9wKKZONCq2xI3D
kb5BJ6/O8SLn3FlFErzWCv6k6AdF88IRxiEPVl4OoWVPBQCTkbPetg7+UYctkbbIuVuhnQv+E5vR
s1ck4SYyCfUjHoQjB5fIEWD0Jx05kD7cNaniqgwMzlK0VwtAkSIizPlukB4jLMowUiiE6uv43/hf
0W1LlyfqJBm5ydQgCmaa7EDSLKAcYhVtPWO3mftL+zrpaPX9gBJZ3PNdxJkdy6RHpMm0VIiWOItm
6vkAdUHgX9NMFbVMt1yTj/ZAJ29a+ajELEkjU0C4OZdpBBrc+uQRkPV/kw/9oEPUgDGIq1TZ9UEB
XLd7Vya6oDQIGtYwObR6Wl2D7dGQLXiaIZNRdVxUDzNsqQIC8dIMY9sS1MkI9RRyV7W53IuqjzuI
2NtHE2Hjnqz8MloORV5/aO7Mim3RpGtwSxHwdfJt1INsUb7ZIX8MqwycY0JCMdhBNdl+dVUP3nwA
witERSLrbzmQsHdaLb/Q0yKILuaYYTm84kggtzzuA/ST6yNjalQ35C1dnXomXTAeZ7VBcPOdCZ0W
V9YzZwiwpVlSByJo067HMPaINkWH61/sTCWtlDSkYgy7tBTS+4Gb2I0IFmPNAfddhdXYBZNS0XVT
/noKj3gWihDgrCPlzds8qOOo7CccZ7UqvgA8CeZClyi2v+4sLrR5p3N5CFEPW0G0PSbsFqQkJ1Hl
4iitBB4SnJvea1TSYT6sxIbcxrwz9rrH1+3XyGBMe0gC3HJwF7ScS1g8+YHoD+OozpQH/y5AEwFA
ZIqgJd0tJqMiK7wwxU1bxPtMSINCcMiRhESHJiuMfhn/fb5jV7+7lTgQYoeqYFHdyndhqOl56+1m
eCLn4d64qG0+yBkhP6A6g5kW3C2gvN6jbfDiGuIz0eAn+aOnUHWY2tjgCFJ1o5W/H9yoZC1gdFya
bHOL0UVhQDobmJx6U+aj/E5z1uMDagBHtBtY1zk/C88fZwrWRp8IJvS4UWOAFrlgnKkrE/nTQuL4
XRGUovBhx/L3CebgwPUq3TUsNSScBQeBgUjq3gnwDaDU5odai7MplBY0ZW1tVu7nnayRdefzZboK
KfvN9Oqk6P9oW5WOKDawIhxJf9JBA2A3TLnJNedZGJONNaANTtMkR9bcwxs7+chhJGBjtQ+4gasV
v9S0aCHeKsnqnyEXCxsN6ruvjsVtdpNugGf9zbM9T8gZpJjevXSyQF6mV6nIxPEQBiKSToKUB5i8
JXeghk+GS+LgTuJG4Ke4vkP/jEZFu6gjN8k4Cf3mhQhddba165JO0nRUF4e9u9bh+t8XnlTsoQWA
aVSWaAPA38CDQfYPhyqgkGskt4BOvnkrSyEaC1r6/cOLfSB5I9D4+AS5Eifs4EABcOBiY7RvYNkf
/1FING+sRk8PdxdrtYL9d+vXLzyg4FIWqlTauMd/KEHEFPQY9fNuPaHAc0oTYUJ4CxWqdNktdsq3
qUtXh7PpYcs+lPgV/uFL25N5ABrwD5CM41uFdAlWQlfIQeA1GAKN0Cm8/1SWelAVyL/Mg1ChDii7
YxhYoEDISa+Z798R+kwl+2CLuQKlwy8CHIZ1/fXs6eEPVbXUcTcPTBT3MBwAquNL7PhkoRlgcGls
jPIm0iU69lwA8qz0BlFGje/c04H/RTUf/B2JunVkahLoOe3uWF8oPgLHVaIL3tymIq53tmkuHzGW
s+ySySrj9viClssYFMvpw+7z6Tyjb3lhiNyjoqTiCCr7J+Ov0TXuz5F/opIEPG/y684vrkXXYDos
fy0+RuFLMoVdWI07NqBPhQsyNebSrzLpin3XQuceH5FpUkpv8sh/QXn1rIgVAQgCZBZwHSvKLBrP
akursr8k7lVtVSGgDrap0l5sAcy2LWq3vORrAH+hA/rZiDKDMpJXlJ4b8N/+x4ZTbO7eyJw8HqPn
zjjF64A8rH/rczVFnea2w2aDk/hRehb7s5BJ8iwL3hTCJGkGig/Cnr+/iAfWui/MlsCx6by2/pVL
8k+forTgCbNGh1AMbcQj0v2cFH1ZYFm7yRI3Bc8ZFZcqZLs1f1Z0Yybi7Bmxgsix/wqaGZcpJ6Cf
hr0SwNjxheSX6OB2a56SW+OV/PQE4KhKOUFZKKOQL/E8ug42jktvJjNZ+Pe7kYaBvS1O57orN3NI
cXhLr3JP/RjdxCVSF9LhN8cC9QUyeFkOAxmVd253S9lbS0OUAIQ/KnzXwGEQx9b6mIuqNVSJEoPE
lYAJdG+Oe84r3+RKF87MhjeOjdufurevTWTC/AdCBEV9KidNDzQfUJcKdITMGUeTWcJIocMpFlHh
qA+MHa+EURfMYU2MGESCiQVGpDkO40NbCqNSWVC7Y4zq+ArSbFsye8Mms+VvkfFuYA8KuV1H4EHg
urp1KDkkoy7Hvg1/tzcv3XBv8It9cQLE27SYtJ9Xfjn3SwJ8NEsjK8B2usMx4q6lFB3aOIpoZ0Lh
jrGstQfOsfXOj7UHdpMHGCAN/AO048XFHUTJuz3w1LHE5g+sfEPYiVSVmM0ADME9cekyP9DtsMOJ
ShkSctchlk95TXzh2xBwSb3qBmXxqIu0O2dcJK0lrR9kMRowU0TIRDmC1JVjW5TYiGvEvCziq+eJ
B9cSVIsz4SAWLbQ+WnLE/gVW1OPHcgR4sV/NAzLcEPBVmN/WxvP4fa3PZ+XRCweaqh1EScLuvrjF
sU4MO+9M50iePKqYyrfRELJICYyVthMOtACPydL2ck1947aCz2kDudCDdSFpMHn7kAwlKfxtUx7N
N8Qj6hYKtjG07ojld/zro9Lja8fR18ZqrCNSSxKsSLen/Glyo88gyBCPyak5eZC0A9rDr6A4QWKz
JBRbrWWE91Gs6Io3dsC7aJ3APj43Ayj7jtrKKjb/pNObnKkgKn9iVQp2FkjOuUHU//LiGbLFsOit
TDVpwBmx2xvouFDiPHgssB3v8KxSEjOLyxRzuOHtqmH1SyhhsEpl5WcmLfDjAhe2I2MyuRNu4LIG
HcR13PsnEaeb4PlV5Qqpdo2yLrofLL9VSU78xGNydwsIahZnVkoFCIKvmAEZTWGPnYwrx8bMwPx+
uyvha4xUZcsklcp8vruAD5qIal8VUHkyWLMRlQw4t05uLWrcCPI2oJh1NO3+gTCRi4nOzf242/+3
wHrIU5ebJHyx+93aNHmXEWod8mrrg5aWdYD60AyFZIapuCcQfjC2GZImJ4LqNoPDTgJZA/9JZnO6
vBYpywsIO+9AxytOT6D853eN7oFlscK2v7B2+uda1ry3dmJkLxoUQ9chNtTUodnqYW7eb3eJHm7J
ZrRdrxIw6r8Tx1dQNfSffY8Sa0pafOQE+AwXBHeY/X8FkeCuqX0mo/XfeRKNKjgRbUCD372ERCp1
S/cqntqB0LmKXzvU0PdmP4mjtfokgxmapfx3JgRDb5xecK/juQl+Y3cCtJuBbtnr69D3syHqqimY
Mdrg7NobAvPy9AxSHqnvkguTS+QdaCFcxWjL5LixsIUwdCib2njaKc36BMuqZuV0nZ1fiaD4Ez5i
cNxPdV4ytlTyLbAbVKQgbaO/57pXutj+KTkC0h3x6Q0Rbk/bUNH7YLMm90v5lzlvFJDQzeEq19EZ
korC/8ZEKrMP+uQDjcOeeuUGfYZQI3FqHelaO0K3U2pyQFuUJ2vhWple9pdkRArFnDiyHZatHf9d
rFSE+3KPd948xWJaXffGfJpHMAH0CHV77JB0c5X67Rv5tD6cuSPrPSpAEsrBW1skTAvfGLrgh6tQ
gmQLDWkc8v0JBb5YtaoC+TclV6Q72RanbyW4GbnpCt5M0wfUhEs4sps4RfvfLnFeZIRSX98q1/IY
rtA4+Pgn343aZmhnUx+HIKJpe93FuTFOBaog+6Cpemm0iusYxPHXMJe9JiVxGFiAZ0/OPW46hdjd
jNI+noFg+P7pntlZEOFCMWq+BG2HrAJnzaPRCw/eJ0vi9ArYbQMitJxMUMK1PE+XYgYCcPRfEeMO
/f0c0kWd3A0LaQTTcFgXGceKDpnCiQrqp8zR7xXbPJwdrWXIAMQXwm6ObbK1y7Ji1AxpFzv2ku83
g+1uOrWvNGeGczpss5hBTKTweRwZLUqOSsR9SsLIm0EpZjo/6XJbxoqfyUYdR3+Gup0nAi7u4Rp0
GcRSKZMdjcygEqErRgv3gXUWvxt+oGAwZZjceDbtYQMqCaHe4FNHsn5KECtWD0q9gCo2Y75Wlp/y
5kwxYJf0OL2PMex+tde57ZrRIyZcz7aY9qbJAzcHtUiNopsCFZMJjSvFNEOkNreZkz8tLr2rG81i
KcIVDVtn6I+XmPZ3+9pangu1yfb1Aotnj0R5U2Z6kpDcEFfQba0by43IJEwFV5wLiEf6HueAlI15
e64SF8yO0dApgAPEBjR6YMF98O2l5MlHjTNl8OKeLvn0HQyLrZTqZeeN7uLUCQBjKmrOd+M+Bos3
/IddHq62o7+tZeLOL2tZytWkW//7GRFXAPBfZo77+SxDKVbPKuY+oEvq6MZKbCDQ4GHCOMJOh/RF
tae3gyoYR8dPniI4QzlCfzGHzj4/NctN0VSPof/ECbzrdI03fCPmwp4hySMg6O+RpJ1z+cGguCpt
g7n/ZXYIMCWzLUxr/R1vqVzGS4ZK9BAQmBxRCMYU4jdGDTJaeFbpXUJfPvbajaSi+bzvFBVtqfGB
fSItonmtg5HAboQOEBZLJiCwfmPI2kCKiVSDrv22qIytMH6CFC1RT90KluieG0T6NlBFy1rbL0YF
z94Dboc7Ekg0G/yfnNn7h64J4aR5BcMWOte3IK/cKZrgAqdNtRKo0I9HvPQcbP6WGmdjgbzSvt59
daiAdfVXfFMFoeo9DG5euHKMZItwpQIF/ZAd35143e0JFsemUkH2WZC37UHr3YF9syGCwrneyMCn
GWP1eYMiHoui2aB+0KBPYqHCucbBo6Xydu484slzrE5SfImnE2dIuP8fUkxvDR+GNeCdVO78HEOM
gqVUyAJ5Efi810RE6pqyWyVAd7bw8lby4n3IJRds9p8o1HsN8cNI0Le9eq/Ari2l7OJTn7KhUenc
8srnyAXjbpWr7C4AkqewPYZLwVh9mW07JkMIM4QimT74P9/aY71MWiHTPOfFArmA53RiA6Df6WOi
hCjIh2NONOuHyivOfE9H1u3glATvVk74IbXkI9olYaNLX+xpLW5R2ckzgCsFShmD93TY86P9dbRn
LGWgq4RALK+9ot3QRwzaPVOVfmzG6/Rf8pv9VpUb6ZFlo4lAUp+B/mPwYDNnPGbW/SiUTApLP2Vw
swvItpLXTARrZX+tAUu6gLlG4Hdztd/IH4INI9MbVFOH28806sBkdRXppcVlOFpNAmh3mRgHXgn9
HI3texZmORTdvvd9V87YKDk7q8vCADoGfQniS978dPQE8Qx0Gg6R5/Fw/OpDCycG0Si4CbGiA8p3
mrDI4r+28IyH+P2SmKYgLvJvjP4Mciy13RtfY2tqqYMgPQC/XQcqj6FGMpreRUmAJyGvf9zFAXZ3
W8DOZWXAhx44nkJ86BiuERN7tIuPtlg6Bi24cpjToztEJce7OC7hBdgjd/1ztnnjc5f+w+t3EXG1
FmrPnjk8/SrTYWT+zB0PmOEh+jw2U1deazYEajD/Dn58Ky25WbLQH/EyYMhSe/8GU8RbxQ4FK+Dw
Gu5AGixicSUIKJgU/P2jfQTfbwW4MnNuD5XOt6MCm01vY03r/9KCEQ9pLwFNkY+OB7oysW6TIMD3
qipCl2Op+ZsSt4O2csB6Li6VK0iWReRBEsVDAvnLycs+w9QN2HZv9zclq/T84mHJLdwSfYYgXVWT
8r2BMPqKgevuDtjlj6VGLqPfcitfpWTI4bVVOcpKHwm2ucLWM1/Ai8Ls0LKsGcN2E8taNaeWzYb+
JNLP6d5c2m0AJhanX+kZtRiPUD9tJD2MW7G3JNPrSgAShz0oKHZm6/H27tSzy6XV6jg485x07APh
2zGPjkKjpCoNgmd8IZpOOCohIb80TaTWrDFfDg4XRn5l6/ZkIuFDk3x/kg1oVsg5W4bGEl/RANQh
aZKifEi08vIS+XLyIBp1/c5Es3E2UQcdK32pLryP2oozJ50JmFNfNqfvf9K4s4XdSTXyulxtm4e1
HO30k2IsKVSlsdHXLSRU3ISDDzgv4QVo3rPls9tePZxq/KK9ORPQ/ysgdQkh7Vde8rxT/eVp/PuK
7Bmv48b9+kjykVgYcR860Eo9fBOD9Gr9GwkEvSxsSrmbb2MNM1Pv4Wp5JE0FPxKiBJM7em29AFKJ
GGu5phMrXndy3Mgik3HqSK+D9vZF2OsA3MQcMc/SNJrFEmCIcLYy9tV6bvddFckVu5BZ98vsquac
e401tYwmtskmZj5gM7EkcR/nWv29YjLU0m1/1J5ht6/G0exzlyVpNBq3/7Ghlo8Rx8Y02pdj9P17
dvoWL6VSx0g9sICVpaIq1Xi0fCB7w6DQo3bWF/6jySEuDu3sD43CKlr4/yiNSdAwgbqLw21U/rcH
mRxFElvbEp7UQD2nEldYkgP6+VpbGsYSdZHCZvzA3bV/F6PgTM9yH/XF7rg3VCdYEOTM0866tc/h
zg01AisMWLVv5aw6CiJ3dZFQWxuvIxn1McoYs4RbBHdJXZVx1ZJIt6QTYddLf3uY+b5pWn8va0rI
W2J+prZqkbcsI8zjfddhJ7emrVI82/3beMPDM4+GxzY+r13rB2/kx15ked7nIjq6Ca2aa/P6asVl
w80kKPjBveAImEJJg2XpYFvWz1dHkrP+Y20f9HJxuTUk2dzd8QKbECBTL8/Iz+Pvnwqm+r70emvF
S09LRlhlT0W2J5T6HxY8UOD3TL5tnSB6nziXq5IN0MW6+Gg9ZEGwgTgU0qpd74PDS+P1tmWcMhlt
Jgc0OZvX3J0hjGusocMgaD8AG8/jKk2m/woNHSt5mQzwnXXBKKaE0FFjuwS7yY5FYXYP3bEFJfaV
AJPTiymxdkbudkC6CyYiFQZx8tgJI2T5bwZSKMFhFEblqltN2a6tY8/vo4utjAVc/nZax06rbi+E
k3f4NJF7nwdEMn+WgjDtZlV8by2ySuPw+YF4krnecWd8Wgc7nlcU0UwsEiI4qvT3+ePuzwXeKarr
87KcczRc1Rs5OGBS89bRTLD1/J5SfMW+PlGmsl1FHRKoZZXxPRSMJzTFqvXbretotMtcTOsCqZAU
APzZStbN8RYR7D76s+qeTPSi2E1d3Y0dpLMb/4sOLxvbBlFBIHms4uw6BaRssKpXGj4ZhxPjG/Am
bQbSwzhvfzpbjpSrDiVsjSxayT7NaUMu15woiMZVi7wxqDw5CEb5R8lVaWXaovh3dTSMLRABbbaR
B9C/89jJKNdon+a8a2Lz9wFnxPq08yHvYGA8JImBfRQPwsm9cb20D87AMqrtEnycnUIsZn1amXRD
UPV0TIB8K4BDa6YGEUOqCDZE04aYD+lw3aSc0eu6na22skb6bLFoJXWFb9WrEXrmi+8aJhyhYCBs
qXJjxZD4zXGj2ckWYFNltWzMsLlzDAsIzUgt+IJU9bIvWcWs3uLhdyLHiAGOYvvAfKHHT3msrfHx
doFkoVMe6TloDQed4R+qSsU+CyrPl21p2cvCsj4+21FqIONgtOAFpPH31NpIJaZt9nHnKDPR6LwC
L0djgD1DchCVRTet5hEk1RkQqtUxu39umkBF9b5NShvrVru0zcMlq8dGEllRHVu+J8QMLNa+oeoP
QE/FBiKc3dpZAMV1lvE7HsjvyRYNxgWrMiBnMGFejGKlxwLkg1KB3eRFfocZmrQX93f530XlOOZJ
G7d49iEeDtMbEF4GJ7/ls/ei453VcwfdvCyGC4YNtbdszNT7QoDh3LSspehYI7nWVBij/2/4ASFe
dZU/0bh8Tf14XoXY+61mE1nlmQ2Dy0XZdxgT/YyJ7o6nO/p4mScDoTS2k+1rGm0srp3iIeEYCELH
BG3RGNGJAq3MgvrhJ51PQtTc+vWgFYM99RkbTJTXmgaQrgwb8waspFc9S53yvCfQlJe2M2ITlFnb
eSEdhVInMNlbrePJ6QK+pdcOb8bDue53tqXR2kZnT4HeaHrYBkDrNAw4QLxkRNjUncee7sMjogmM
jVmDFTo4XGR5GCua8LJHyZhmHAEMc7cPxPfHZdz2bsOFgRSNU8mOy04WMweptiR++PB5uieMWc2y
szqXE/5co5JTbZlEnjCPakmLPBZJ3ZtqcM6qfHR6QBamsg9Zhwfy/IHvij0b0oP2WUnk6FQGFqJh
oIX9QabU8ACJsG0fVZRHSmdpdOKzrDKVar2N34z9fgs77QZcnfWy7xT7HOY5tyy98OCtDV3PYcZA
csmiOXmCr4sUKQOfkZ3V8M/oW0KYRTn2IuRasBvwJTf3F1SAAaYrXX5APqoa2myEO7dPYh+eb9tT
Spbguqp6S4v6jExFg3HuwfpCZTflFI40GYxw3qZ1Ql+J+XgVTMACvN8hAT64pFfenMEqaw2JA8cL
83B4ThrgHtbELPk/wGsbHQH482O2NHyQi5g7IXpL+QIYwuGeS6F7ZsV57VbRn6KmgPlYHbqCEgTY
aEHErS5xnUbBGJJv4HBZjudG5m0W4LVIoHi7JEmLEyLdFZvjTTIN15FiXypCIg/Y4xQh7xEODE2e
Kk0O6edyl+XGgnWRquTbRnRTU/BqXdxPRs/GhEs4KeVUtCyGja0HRigV5G2D+rlPKY+uLlV4/07g
9URvx1vGiI9fh7s1bIQSrAcTGDzpbQIfb0vS0kaT8ohCvOnu2vY0MuUR9aS+0ZTAVXO5vpnYtDys
gQt39KrVI7wZUGIIugHWChWHGpcB7+Qn0sNiSEYFDTPCpJaXvXr4GikIHzkMJ/tKtNONWUujJvxE
1b05rpSsfM0E2QWI8l5XJBzQgHSmVLhOlganJAitnZ0dgfmRI35CdXz6+DX2XTqGhUmRJLou6y8N
31xYZKRs6QL3ox/LYZBWqLsYzvLWVlMkQugExpdB8+BLzDVw6YGdiqSGV4NWdQlkqc6PepJQFWdb
vYmmMqe5NybdDEAH9OkTOn5AVd9qsjJlmktFmOCWSytTlFPVfrGSuVoHHzaNc/kpzTWl0XnepO4K
TGbisQisP+uuttbxRU2tGsPBzAIjGTtZpkMhfb2nU0vfK3a/2phHfzZYFyM+cZKh/Y9xUWgL/DPq
AzbtfW/y27HgKwHU69WuvTiqGU35FQ9p7Twx+8QK77/K1Bi0seaX7Dpmv2PYJeGVrV7quDfVWFU0
gOgh46nqFHGJ+X4jXAvoQbYfdbsWpndFd+0j+URyvFCuGfFfkCHKdhyAbCuI4Z8p4TiC4QynVVlT
FCDCovRjG6FehHjOYHzQ22Qerfk1Hq0CE6X/SdmuvbOYnRkYMPfjmt7ZrvkPEdaDRD+v6yo+KhhX
ZjAQbvriJwol6x7fvYkECnc0lgu1d550zIMKfT76H8so5KYSXymSPhkgW5aG15kapmopjpidQGV1
k5gmGDID6vX86FrYjYhyiHsxLRpub1AY3nkpU3MK6z0Zup7hs6sunlHY+6HQFoVGKV/9UId3OEqw
dO2YgIqAANbP7Yx/JW7AkQ+mN6PQMd2+tsaRXrdCrLwTZV7jzUApF5IoZWrw8l2YGTWWy6KsPv9Y
f+wG4jkCeo81Tdl9s2MenjBBWIZdTNM2HBXr6qiRsuLNIvP4IDht2ogtFahj+byr/7zhsH7L+bDu
NSvI8WfZk7riLn6Y6nisbJpRYOTbIEs3/0oN42A+wjAyKc3fZsSN/QM+3Cbqf0zK5Qw5dHe5KH2J
+2ZwTmVFjIKxH5s4lzwL8qHzIYQ6aDAgXuvmP+Y+j+P3OEmp55HA49hI8iGbaxJxs1CaNTC/0+ik
E81sTZkW6WJfVTZhYryfzx94Z1XIintuuWAPkGyarKtiPwTEvI9FpBDAi6RuOZxJx7xqQSAt30FD
BAvQ2QihJ1hdFew4v9f0bJ1rLwptDA1RE6zdjkPUtd4+T/c2UhVMsUUs6qA6X+2GJb4jXkJOk9b3
ZixLVvqc0ktu/j3IHcmiQE1PytyGwdXz/Mm9Sv7hml4ZunzdBtQl3+LxHhlHMlcABnUMa9wHMyxK
qI+YTGVQchH9uQbsb3+UVWQLgWiYC87N7FCCA2/zSbiOnX3wim4b64BuRyHUsm/JF36ZznGcFZ29
ATz/wbyHmTHJkri0QwdmMSNhH8tCRp1qUqBjKv9hgS00NWscvV9jPYcaUD/GvrV0YjzRSiJl1wFx
GP6Dt6LikNBGeaU9ohW2dmeLmAITS/czgO2dUMikXmqp1FItyLCPmxbIJPxnvIRJquh0j8TbAVk0
huKLrRICOL0lrKGmUnxT+fLnkymgjfFz98vlIU6ZTvPbJgT/B3AicaXTfQC9u8mf5/27JaiA8Ajj
SR0B5M7CoPhLPg6NmybrGiA3ILjP5nxIf7YeQ7laHibQ7R12Gi5VRThMZ3IHxdqGuNb+q2+tXxuM
1dphz1+tbGyr2h24D7NJV48W1+SFG+E3hteRJ4k//B3DL2xNBoyg+0JM8g2O6x0Axgm8wBbzkOb/
bCdSiSiYGDu5/J9X84dFh6bTF9uLVoRUyAloXVpYNmtnxttIbqwFxWtrOiElzHdHkJtjZHOwzZK5
NdAoW22zCEUhnL0WTmBmtF14q6D6li1aaja7PfM4N1Nxi2tkM8B7HAWB11iWiLpUmrFQjQrzSpex
ttklWpNn6A+HLq6c7IxFW5fkR3jBELMmwNxm44CwY/ln6hb3kxhnNTuOkXI7zzjDL6vvzXB44XLV
SPpZsEzIIQ/nIAVzJSTV/GjDWAVijvOeTu2u+X2XFtiiXcMMrhzlrXfg2fAvaSYmBER9b8wtXrSH
BByDRdq8vTHZFn8NHooojI+jeSQTSZhplW8QSq++MXrrUil+h+3T9dym3ZIzxc8FTYKJ+q+aTdni
w+Z6ryDE2YKyT5V+EqKfeORtXgUGKUa3DJNgMctdIpOzso90LpaqYSHHxqI2ekCelpGTYpH6m/XB
zsAqK7kjLamdcKzksKa/zMwOLuHkMrUYAbu8FXe2iv948DfEbWygLTs5a8OwGJ7FvzKBBdg3NFdg
OFyez598WEElRTHwrA57EJNw6evkbjDqdtyiTKNvSTy/13gfPGsEOUpg4mzLoerbFg4Qep7+V6NZ
4/4yAc0nk025uFzhCriksAT4oaIJyja8qW5H+EL/NMZ4y6SMe+TpZ2eOFYe96N+DFR26/3qIXxlo
5UalMmaEmuGFISf1G+IqqT7B5+Sh3O1ivcmFCAz0MYzOQLCEV8/nrLUocRy8tl3Dpz6fd1u77tND
9R7pKT5u+dnL9dU0o3u6ER3oYw8KbPtbXlEHrfDwyEbXrfPnvCpWntGjEVDn4inrp7Ojg+4/rGpK
p5Maaw30/ueFv7ctjTcYveMJyN8/XCk8vjjzpMxIiPSYZ8pxspngjEhj7n3ZXFIHvur8FVe4/6yk
tqoYgvtl3ue/oKpLyr5EN5Vc1rj8Qt7ws6enX85NTDTwyUKRDFnVKP8hIRgLrcvttRcgWm/VVUnx
qO6t3gB9iGAbI7UVqCDEjQ4Ld76GREMwCIH4Mqtg9gzjryTlKLL1r2WMwlxLbFF93JMpC1HjdI6Z
Hgw2q1BI7NBnx7Y5WxDW2WgGLXUm8lA1SoTyfEHkPssCrWtXkRJCsy+wlMmoQCZlMrmwN2hP57Nh
KZqGnWwQiXej4DCb5Hm11gZ9/4aGao8Sbs/hq+sGvbiAT5xk5xbmor1ULla29dTEdKkwLupimhYb
iooa7Iq1clgPo8C1YcINrLKaMIxYxOEFwLMWBcyuBhR6LundTEC1xwqk/WHkv/SIaoMXnMxj+4Bu
qK0Q6kK1oUrjZucsUStbLg97FfnSChaUXVZMlO7Zt98BlHQUpQ5dNHyON47Xfv7em2wmO0IojNTL
2CtmyZtcVqvA5vVfSA4mCqP7lJPj9gzn5XrSLxE+8nPOrN9vYBsbOwl8QKWvGP45AtwWG8ahOcjJ
VPAZjq47/03MPrUDY9pKIa/jiOmIMTqt0XH5+kJFbr+q//B3kYC+DDLtd92xmAVVWWFBhxKY3J1Y
9FXZkRLPK4PpE7gN2kESGTA0tZQq8nXqpv859fspSTlSbtf+nTaWt54NReftxDHO3rOkSxBEUORL
fGw2VzFMMtwEtO7zTuNsumX0dGOhRSAbvuZWIWrk36aLdBaURD/kq7HSI9fkih+qdN1SNv3Csy45
XSRbahcu2xJwDErvK8s/ZmkzFRH/ktzeOOpTFc97afY7QjEn1dUDr5AjjSyOxKqHygFlY+N3nXSU
uVlym0hzAL5drMUzcILvHB5TljB/KGa8fQNhr72Bi2ldOo0QPjNIHBheB4CcvQo3BJpWVrxOV6Gb
uqafAEsoIDxk1U0iM3DyccKBnPbV59bfoKV/8nkdRTGdh495mHqvaVFOohiLXPhw67ltOnZoT5HD
o5G5jaB44L0HEFdMw35uGaAbOUqzKckal5S9GHvnlGA/duFz86DdDA5V/NHfUL2NtG4b0zyGbmi2
wqlRWT+oAdOQ3IK1CVXNId+6EWA8OHHryWDTflAoqTdyTpLOxZqO81mUy+wv0dedvEKwia7BK3yx
IFQcj+kWw5pxBJLlK146BHRsp51gbKRKmkzTdewxT5KKKQ2sKFmStk5TyCBPrFcF3dFnWc4LrIuN
rrbHC2KmeFpI3Flpqt4/h5z8uMvvAARRp7j2Ej4SdXDoGxC8VixxnwPrFIiTxCdqpnI9sl2xDeG+
u7Z+8hhg88ugFfqJtgPcwMgv3mo/OcNPFOWasJiIY0VXijhyg3F38p1Bg1H+EiEOI+x2hafQbArh
+NZZhTqBgGGdpxEs8KtcN564lw1F2xt72jQA2RXewY0Lkobx7dz7qsjvw7g/K3mbnVZ7Iq0JXPBs
w2gOh+gDgWBfmaiSahAQEvUKAYL9FTF+HtpJXNPERg9AfDValiaKFghRX3TNHP1IcItXrJhfyi3k
thWG9SYi1XwSGpbZ/OBAMK9hpXZ6LQUDpKwqq+b8Suolzz56wuhxpXwS2KxnwUs6iinu9kflxf1i
1IB6heCZx42vgI7RAwvR/udyu2TgjLc0HIYkmmga2QfFdOoQgZfU+A3uL+dBaty1nG69aXtTQW7K
5f5jbjnoNLiwLLEH2RbQdYOMWTRecG7fJHmEQwsntfwMm7OYrD0cwm8G+SK3gUkF6eKkwUjQo45/
biB6zAjFvgIFfc4oko1RiQ6P4Vns/Qv1M8a06a0Si+cCyf5GJA2VVy+FbBHgjdTup27NGdf/2+y0
86hISzBv9syc7llLdynA4XBV2lvVT9BQ3OCsm9qcfAZYr9zSUjloXo35iquw5LBwcABhlU7FmT3h
MjAatVDzT6B1OAUNd6BxEzu9b8goPsr8kT6gj/RwFK9/1cZmAUk/0pD+KGKNyi3VTjJ/ojtBwOoU
/pL0PPqb/DYwRDd9HLebYkyAlsM7DOv9+pAst4WxcVZIvQgnqPTiCHmoF0AreDnKOW/3A4CpMB7b
cgIfe9KQ87JY05C6w5ooqNq9gsBwMgkimkLn7ie0zX9musFW0wsOznAHUTe+/f5VSsQSMT5Go9ep
tEKKfT8zvR3tSTpKSo3NKufzMiGGWLSKMZISlhO1s3EtMA6TK66qn6u1nLi+X2ckonsZCxBjPPhh
nXXCz9PLxz41Y5nQQaA8kSLSWWEdFymZu9YtYq+PbPAspLwp2T+8y2gpzP9U7d54W6Zn2jCxpxz8
yBGOUWJrX+1HK491CrFvm0eEkTG7qrah0PeXn/OME/N9d1q9Gz2/5OnQV99dPlTxWifltw+Mdax7
SGSo85pvY24TzbgZL6Ng2CnrcPD89f9wHlpuAljUBHBLHeXkSMPPiH5eaOefyIDH9QbVs2tU0bc6
j4KSBQHzPHjft9fMTJIl89hi+O5Uy6Do6XChkxs7MFxZyMBZRg8AcYFU12tBcwLTA5kpX4YROa9t
MJQHMEX4yVU8l7yjuyOPAqJxZ25eHdexMuzdSKCM5ZRIMCh8qmYujeTOSrxocsk28NPXqJucmmN1
94J+HIIsi+s/HyN8DoBoT7z7OtETdtaSAhs2fuYS1cIT4PywnsESj134rpnD+lCmtXMYSiyzlg1q
UCkFsJvDFmNnqq2ADxJyIIUgNoXKfcqZjIiR9fWAuWJgQ6CLTzodW99sk5GMRvd6rpamPGhI+L+t
NFPPbnZGtCdoj90r4hbb2Gh7kyZFvqxYQOqn1ZtlCrfRx6C99DaG8BCNoS5H/9eVVf4uv73ilnUI
1CwDDwJQJBV5tHwRaHOAt+3jbgWhhboezCyV5NyLx6v7NVwVr+sTIard8hY5waJGLKoLFb9hSVfD
Xb6hK+cVjSt1WqDgwVNV8HJpN7+/JTv2MO6K84IEAQkahE3S/yumfMao5+M4LRYHxmmQi330QlL9
qLUc1/M/tpliiTMvNKydnRgy0faTegtIEEaCu6KU4ydvyoT7PFfV8MrcWhs/hGgEBWeqpwUUedLa
DA2vKZJ7azWrDDRFEsGxkbCpHjerMEGpUdwGxeLRreytWz6AbaD1fRRTm/06Tc1tbaOL3SDD5Byj
Z4MYcY8hUYtF1EjiEo8oq0cZv35PStT8/G63tFdFS286DjtkVD7VIsdt14Q6i+Ht+5vQpxO33vK4
5X/VoRL1AZ4RtZjQjyG9NbmtVwjhSLdfcIo8Flg66UqEAXYUTlXaGp1JsmVel/ZmSIaxyl8d0pmv
YVgg/hyxo2Bdc+0nk9iYlG4x1/9s5uiFHOxw0QQ8rbGVsemIlyKdnki/vda/8JgKp6d1ObYYsytM
DAZ5W8KRbLigAw+/7H1Rsuqvbg7IMe87zwMbmL6jp3ddq4/8bFtgZZWRicSv2M3LepWbuLM6f+D9
pFjuUZIk5jwWBI0aAwEPClkEFPwRr8gK//BzDdSGQ2lL/63HQS9Y93qqw3tbLaafT0q6YxsN5IKX
UkjNpMZ5PAJAVAE9+MSWZD2z5RihS1hXldcNi5RPd6Rv2dmkshqNys0GcXHYXgLM9LkjRnriHEUM
vHnh/xgPJInCvihu/YF5i3M++Ax10uUfG0kBBS3QfaPZxJybqlcwk8wdHFpv/1GCQ+EZGwnVvRV/
r+XZc3YdV0WEQHO3+yAZ24+TM8uSOBoVQOzb6vxgr6gidTBrROJ8SxVDW6ihN5YefaoE8vE20MYz
NgrPA07WwIxAZZSzO8IThByHznC+z3AmUev6tI0rSqX6slU+Nf/nvDx0Oyc+G5pqrRWiw9eFy0EG
hJbHXMObhWxppnUKFb1eEbI7IvcIdskpBEB3kCjReQ9K9weZZmCH7a48SJ1XTttrCOgNjGzGsCgC
XOWbqIHVFPzweW6NYySEWDI63Y1s9RCIm3PazT7FuQodrw5H+ic0U0emD/t3IWf6WcY+BNauRShz
8Jh6azbyTCalysncgvrpXnorEHbgi9qoTcxSd7wkS8QF95dceql8jOurD4mcK2H6Rpry1tbwBbx0
u3IoOupMM1BmiQ7fq1IN6hP6FnyfXfZRA392BO2GLABrmLYom52YJyVUyMfrCc1TRqjucYVlQFXT
r6eFxSlBtB2+tENhw/K9Be7RG7DlrldFPUgcHiyypwwOUUlzNRpDCZ+qiEN9gwk/Yz4vuCXwQhX9
meokqv6rJtOiCrcUdEHi9cPoAqFV3K7/gJW1izpu7E895JNBf0Kuv+Ag+eI2MAShkA04jVy5z/2I
ZYw2WgO65gJJwXJ3YvWBN2HmH/vpwhJR1tC1t+0hgGFkQkSauKCKCXn5zxxlsrrghUnA9YlrQh32
TQT2sMx04mFbj+SsfRVwcKTXrnHYo17XmArRpmEZCEfYYovmI6AikmD+cselSz8m463FWQGpr1+k
W8o8B1gDRE77fXZu2YBHsi4mwJpKcgIGb26L7WKbZR47NROuaTzIWcrVcr8AtViLtbZHmiylYQND
p+0ixT+lU10RkzPdjI+rFT9BJGiwD9YHCV9P8jZkI2OlREoCGcpJ2VUx10BW6vNLx8LWAL2IYG85
AfMEaCYpLCpytr0R7MBl2lT1KMAib4kA36VwcpEd/QlXHFgd313N5WKMDgE8q0nbvVy6nMIFFqAp
KsQ+OqYztFxsCltf/qZTK6C4slJjag5PXTxKTn1ll+ZOh+Asr9mloQn5NBTjkxrzWUq0i5k3AdQY
JnyyGy2kersduB7lztWcLF45VmroLFCJCRY8zirJr15Ohc/K9zruZoGqdrKmfEEmtZgvJYGaGcsB
WUj3y6W5MyU3fdTSSq13ilFyPphefR3hX/MZObiVZX6azRjGxLPC0/kGtCjujr9BMNvKq9oMihld
86nEcybCVGo7BWumA7fdoiv+zS4+PwzzSgM9iUiUkmvhfsqokklTxDJVgPsE35YWhuK99bt41Lbo
59zwOgYCegujQXfcHhrwb1evuAEQSHitAOD/k0NMNOF6qA81yB97cL7VgM8j2xENMrQkLt81rG5g
z+ta3aFpCWklb0hLxw6rU6bTXaBBP1frF9982b9aykbYy1bNQJUfkr9w3EPhQLfpFK6Fc3MytyzO
vvr5PuBq8b8ZAEmx2vb5c/5My/TcFtIBTg+c99znTk6Xw3HbWqRVMbWKX2NAy7Hr5s87wMhYdW1H
0NORnAxGSyvhZLf1+xhT5su7Pi7+I4zreY5KrYaeKwbKhocI9AFvTlfn5an+pJ9so3zbvJ7cvylc
5M/yJm0EbA1Bq1Gwsd3W2IJ5cPncvE8YHVbWRAoqOxa3AGeTPayFSvE6fMr9wsuTaBoBHfAukOZQ
/PR+a35r8w2gtQyUu7Nr1joabUfXuALnuFVJSG62b7JPAZyNFt3wyNbJ1RgtYtMWf5dUFh0LO3p0
/Xa2XSIGhuTd90m38fE+eHzhjqRqlZzqaRkk5aTdT56QxQlxjjqYDUdKY0ZE7XWAOa0rfWHTxwRH
t1yjI91nak/Ypu3hf7S37Kj7UEZQyPmxBaJG4/GVpaHTyec77DhjOxH9FzdldjBO5XkyOZ3Y+9U5
/uMgS4AL2SkASbLH5kI7Vk3qp9cv3N6Opz9wrxGgo6j3xrPYOWWhDrMCh9ySowhxLIZNKoA+IA7l
T0jYvsymw5MioVeh6wljPM3dYUxtUUi9sSoxEJN8M4DCGuNYE1F0iv5OWejX71JuuAex2cgNwZvU
Q/tDei86kjb/pUMBlutW/KaeDeq0Q9Sp7hI8Z/iiD+ipvmMw4eXFWU95Qe1dAuELy3ZtAqUZwEzm
iJs0uAvHFpuLgreNYml9P8IrPLxT6OnugZSiUspd9A3U66c8NnufI8ESXipvbzTUtYiXoADwgyw8
OknbUi5rYdJwdHflXp0wf2xOtJfcGbkoN1Wl3XAuXjS2sn4w9gojEauRbgEYIIN+JomQYIbAI0ZX
mu8QiKNcoh9wAtkoY6aRQfPXJ2gZUNVGPkHvQSd2XvAuemQjzM/v4SwL2JP9evSaXq0ONiHN9qFP
Qgz7Tjqtg/HuMVg8RTjn6UROGLc1ScQ041rhxyzxlpE4VQperng7vefwH/7JOf3+T7EY45E5NlMm
+ib72lKId+b+8n+UppKbDtmm9sXzsB8Dq1fMQrfD3cpQmoIR00ssDW+/eDJgiIJGBZLcReHdPQ3J
VPpoe1z1Qk8nGGg9Xrqa4uuGEJM8SojWypmIjQJCzuq9btGpsqcE94yIFWPtccNFHHJGDW4C2o5J
LAdxAZQqb2aU4WmQb/dwC/PwhaHXIAryqUsr8qK2GCBxnGnJfh2hoCxroIR0a3RTlq8ogIeMLlmz
6oPFhJwuHJYkwxollUFsuwWnj45MXHztzAJjl4Fpn+wJpLSDbf/rRpvzfuFs6+8GpEogxQE3phVZ
4+iI9RMBO216eGJXJ44f9Gxj68qojxlQKADPonVEia+Rkt19wsEF2KPN6EZGL0ZH5/tFoeBMzLYO
C4DpyymiIc4VHtX3ae7tnOngGpx2AlOnTqNt2MXb8uIgWc1vxwryMvPsBQSPEGlV0d5U3CF0leT8
IoCr9zNE0QJqOwsnOqGlb3Q+DB8RUXAlFJdRRCROYVSYwSX5jQDCxkE1TE0QsobU1uA2vaIIqkJa
BslVxI4uCDkJFjFA/5vubLBv2JwRr8X78lcKRBuqQKEJHzvo5X562JitKt9UWIkSZop0GCgQPYUx
EQEYoLJ2arX4lAZynM59AhthTd/wGP4wC+8gHKMLMuTeyzLb2r+gGLEQxyijuNNH75sicx54eyaN
urP4SVtn5FPS8d1oXJ9qR97Wg0Hfp2GLh5PaZb/+qdOR0UfIMZUVH0xHUSb6oqw7/knuPy7fPkmZ
jEozFoHXT0rU1opWuHcSg8rLfb5Qe7tMsgScATuJMRAgRckpqulINbvTE1rgFFVNDmZqNkxETpk9
Kdi6wCNt3OZq3ezyI2nNW8H3L1kYNqi8oFHAh9h2MD920CKG/MkGgAlMM8RNjcUnsrAftaFnet05
Zoye2MhMwEnoIzxsmNm5ktwqiNcXMaO7J68Sqi8GCkIC2r0ZTUETusMIX63tplMYVwGNigqXbtCj
z/Elc9nVs9bLM4N+AqdGfnJgdx0LFE1i4nlXT6j+2OLfVRNQqPnmVSj2GockIri5fVn3vcShgHen
EpbNJh26p2MygX3I/DZ8OJmZqhaVf8FjO/gTyNipX1DS4kmDdfEUhugVDxBfMk2mYuunVPwGT8Q6
jhvASASq3/1TAzG3MpiWwpnihGr5Zl3F/nqLS7aoRWZQLul8KZv9eW0LpavJ8m81zulNyE+AEc4n
BKRZOz+qHl39KjUHom/TJvD3KvYifgok/xpzWFbAdVo6cE8DKWovwe18gRo3kWbP7j9cTPhRsdsl
Nu+uR2kkeWVGXk+NU57PYOwwNFXWeOyAxLAEmnkgiJKF+/sSx1Odr/Z657zwpIOtZTY2mjCM0dvA
HhOQz22XlXWChw5xXcT4RiWyNsDgZNOyAI36ZvUmHtuVyH92+C6Mqx9cr26uEybBAGLcWfYmCvNd
9vUGecwG4OYMClJ9QEqOFMBNLUEbbED4ZJNGypIj1nSh9dGXXG32TJ42mLbTobNNsaVT8o13PnTg
prbbWTlxGJ5pk7FtENPaJ/EeHHLWqnSQ06iEARqHcLBL8OjXTWvHduF2HIfIWtykUv2j/znGgswb
Yo5TKy/2QPHm3Uk95i/BBmtQjku/uZYxGGKWHQ+sUBodWejf/Cs+9/5Okf9jRRlA7RFWaup0SILn
8nMqAkMxa8qicCRrV4r594DpMChBURu4Chsq9Jcbcy3+25HnZNd4gJwkfeGOKlH98vsIzwB8obu/
jI4PpcqEUFr3ZV40y8S/cSFKu2JlUg9s2wMlZDmuzwDYtnGSqFfzq2m4mzZy/8QFbfQOMv619bsq
iAZ6hTWrglOGRyl0klRv80WPdK4SFU1htpC92hyWfBUBDEk8MVzyBaATcho75zq3p0ZtX75sLRPz
jHjcq+N1dRfa+JxgpQd9aGNqZym6L1bljAh5bmD9JT/OlJoWR9L92LpTZQP7xFqIN0fHHpdM6vx/
nBz6enfdjrTh7koFnyn4IvK9D4uO8ltOUCOoxjpqHvej24DOsExIO/QD9pudaDcO99suuaKf1JTh
YUcg8iBEhnMJf1Pl4y4587Zt7/KeVRMeQaZgEaO2DPOMXazcKt0BAEBnW1boceNfwSXEDLF1SClY
lt5l53edukZoZi41kTf+tUat3grGHunwr4JOoPUfecmi+035AXoqIu5Bk+8+E1L4xdBvR9P4xkz/
wKe+LfN//DyFA27zfZg/t9DEj2KH8haChIAF3QmLZVrmcbdtWXGhropq+z44kXjmd2o2IpJ49c2c
kY8CG2xr4YaBUbdueUIKMKth5ygbE/cQNd0yk2taXnXOxP1B3ZNN52FktrPbTJtghGkbfodn6Vgg
9U/OFgen2urMlI0LAuyyyG8x9hpRYkrCnNF/F/BN9m1u0sPlMXN/2vmz3tf7+6HKig+R0v5KlSpz
2qeV3m9kP7mnEciTiUskONkYbY3CjvKjnhDIIoPeyoS/gstCLjKIZidKZsFQULBYQb7tlTJpgH6a
Bz+9KV+WfiT9J1AUzU+b3DQOeqRdtqBuO9SdkGCRujXuI8RjMdMLBz1+qWkbJVcCFJnCUeCwepQ9
fXs6LAb+cy3g7U6ciPv7qj69oEez4HUwbRGSUkWMOCjGku5T9zk7/ItfZW4Dyqq7CxEf62SqVrp0
c5Rj4URM1UJYuKj6Kjtln7d7JRX84Ce0b80gZo6RQ9qZjVQVkV31mg9wp6uLmM3QHVov+WLhnDND
cVtIWEC7yG++vrDOYgPafKaXDBiorsdQXSF3hb1KiRnIKcVh37qfqO4dv3OOzNosXXqgL4sTP6jX
NJwh/aN1lFOdZDHjXvLN7qDPZIijtqs1AT8QkWL/aCehVjKjmKFpC8XXYqubeOv5T9TNW1Je87kq
Zrss4YHyDXbibCMXLk6SAfWGiQJh+YJNxWfbr51ULvNCQw1KVHdurCCyqrxCfHcU++ntMkptPCR9
a2b0hlGDoxQCvUuLhURh+6KPo4DJizsMqwrb5BITTEzdO1/sST/5MFv/g/iDR9eZs2qDmfrT5aL7
H4TMNjBfvON++fIUcShCX3JnMeN+Oy0zceZ4sIoVBNeSLUNJGgwHLpipv2Ex6UG17gE1UH4b0gH4
568MXwG9H8ggyjxolClKJ4lB6cMyrZ6FyNhI1aMbH6dps1zi8ZJrk36ckXZJmkzOAGhR3pekDo77
e1kzgrONaHXPDDldYvHonwqgXHEanKpuJGLIsrBp/TFfFSgWOkyr3NWiHQ45jd1J0eQ7QEgK+XeW
MSBEeDZC2Ki2ytcLBkBmGuwQjOXieG/RXjiAdddyHKgPV/afMLH2rfTsGqV+VGVfU58WAZ5K7MEW
2IpcQ8XsvzFgTJ2HWUTHXispmglgdXvvseA6g8C4kIDuNBw9/VHrp7OXNa04X1xAqnwQ9BXQbfnr
NJ6HlFiT2XBmMxBEWtgHQHeYyUiEV7lxPgBxqsagRdD3480nucJpB05NDETKiEk5auIHwdyX7frY
Bu3GyxwTSSKevBBkzexsl5KbPoy2hKUFYQE9LXCsjBHWI52/4+suTEEsLzoXy237vUN+GtbA2y8K
L+dIV8k5zp7V/QAyVcmeGdF3+OeGdTrlZBdZchlwzjRbyOTum6lvf3Tca80KJ43Re3uhbzstGs4D
3jjWtjJ2g3/UDOD5rDtIi4SR4PGZgNCDYu4g7szguCoFsL+qnJLX7NLVPdNm8vpEm33sbFzaB5GY
yTPaijogG7mJCO7u1+Wj8HDuu8oxG/zpgG/D/69dSaBcrFgQko8Npqk2DRm4hAUVmUq5bVCgj0+y
FrUK6NBOjzll+ANvOhWoT+9zA2KwSGncH4WBLVjm1HMPNSPOyhpWkO6D54xDQz9bOfzgGe5GeQyb
ZaL6UPa4vnbzaMbpE2CoxZ5yRoNT+n1+cnJH1ZsXOF3fckf5dXcuX7Pj86Sd3B3uODUU/mv9MhvI
9xPdaiID9VEyIFvAztpV68ngLg9YB53xHvlYDbbnCzIhyCZ337H1dzAawwA2Yypnx1v2lQqTpzVC
GL2FTSFbt0Jtb3fZgnqgJiGRJRVsDhs5w1oHJaUH5JkhbtUEqCMwGSnsULeMyDxmOu9MyPxcItOs
TLpe5Iw+MNmJh3XnHQL0uKVk6ouDvIyCD4XZDs/u5je5ml6sxCvYfaZk4mFVz0/iaLiy0/bm8o11
0MEkPOPFxKOvdocAlheZiTx2UmvIdo1HVn6/2V6Kb52DjALiSMtM0AycLJ+CCWaP1EB0UHq2U/Sx
km2STCKPzmbyRbJBQkcgpDe5tGkqjBpZjqPxIM/WHQRflMlMLN7Uxvmspoc9h2LeFUgZ7oEWLKhq
PAp+LzFyALJF1fQJ1vlhxkITPErkSawc1Y7JwkSgbHY6GbjXPZhHJMOfpEFjFMvhAXD9rG6q+0Y7
WgptwJVSn22/G2jP/B6r93F2iVfeSKAnIIR2c1ihrSrCfr9Eaz5hh7SHXpILUyNasOR4BDysMf4I
eQBWvcTRiA2UdsrXWP2Z6nMm0OeoY5q6KWhaN1vJNmZ28DnIbVVIu4ImtzOkKxRm8ycplODfqnN9
ZuzDVPS7ujlnkESZMaDlIJJeu7oM4qjz6x3B8jAsv6wz+ur7zk8dW/KSch0YkwFRA91S466CnFrs
/TQmCG/dP/IxedTcQwlsa/dgz5LC3/kUj85vbr/GAqRPvT0L/IL58Kli/sUoPD8b9CHAeHWNIe1U
jjKc1ZrV1B9+o+MYtEL0bacGcOnfoj4wd/TGyyF4mHFc32JIswyro3se02jSDgddAmYE7mGrrjap
S7M/8JuJsK8+n29tHTsruDVhjwH5ukZzyHj5jn+s5gffy7zVbZuoTHFltcEGV21rTcOVzltYJL+T
fUQkc7saQDuIJ3ZvgIrlcW6DyUHRwDOMQOmNrcNyfK1IvlHa8ptYeYDMJxB0RiZdxLV5KRT4lXGU
NplXpA762EtNPqc/EsOH8G0L4i/ukZNt13k042avcT5lUR/Um7TfHQ7tmBdCJByMEvXLy1l5Srui
sUPHSqCPZsQFyri2LmHTcQlqxiNx5H8TZRl0lbPTU31nsL4TGl0tkGn/jUc8k6rFTa6Gip6o0ZSl
SCb5QcbGQn7IaSErB5ijAbR2RfDQKbqEjumRLM2qEJ6MieEOFmC9tbxJmftzHQZFSH+I5YpiEtmC
RXM56DMDuTLMKoIQPblArbAHjSA2wLVyODild7FRFrJCbG87M8NOFFu3HgyjZLqav3WvOkr0Mo93
0mf8MoX0ZS0myQeINhIVxgOLVzOCN/+asu9Grgy5KXeI701l8SXQdLeV6IP8MAHbRRdDE6VcdmEl
p2QC3V6RKdwgd8DT1q378RKYvDUq+0YfJpHKl2g+1Infuu0HgXj4IdWZAsmYSz9X8cj8snVw3kCn
WPwTydaQalrURFpBQGml7HOCReruzE2u6d8qk4CwEgyTUlga6xdoJGVM8TtaNrz3fDyOhlrMcuxi
PEX4N73zoHoOQntkY5EZ1KIxTmthwl/Vbnsk/jFCKsd9XSmFHrVlw0/1ZAo+m/XzUggo2Cw0rKpr
l3TT5fystU0mTuozmTDxCj/2kLLnzWoEGnJaAm6RwgzL9p9Qq0XxTcx9EqOpki03Di4XaBRLH3r9
YyP5Qg5aCaTMsIHlsK2RYsBgE8ym+rGO9IOgdRZOZ7cCq7eIo0o7nRmgxKBKWvci/I3a5Z99USee
gS/TaIgdnpXybtehBEbCcgf8ojhDwHGmQV50SjST8V6b9/vo5jrm4x4SO38bVKDYQ9km8fnGfiRt
JfL7kTyN1/xOvFDYVLxqJBclp7l8qQM6gYtaxuFNDsoWB9//hej6+XwRWwkWCtY5El4F06vlp2hc
B4/Udv+H1usVf0/RnWnNw+ipaD4vqfJgRRo30Tq0PmgLsjO3Setow3WQeNIhJj2W7H0atsoorWkj
tA5C6KtHAepUcMkrpPCpeksIgzynYLq19Z2r9NWMsjVyxiWcRLTYPsDDiGu0PhoJpKPvX7U0Wyx0
aDNwMJh1v/EvI19GENVfIhcHT69WAWiEuczYWYTe5GCgW7xnaE8BtUTjxQZCvGF01FKsFSeYkFUE
bOhMXVf3YyDnxip3v1azfZg2CxRLOclwHQ3Fnv68IK+TMlWeyGYnK5clWMhFYNRenTLFaIzn8Nax
eYFbfvB1CDgqYBLsKyw8y1O2NAsYG8/7z8gIgXGYSPu1Lszr/5tOmxkH/ZSsRbVPNzj5JdfM6uWa
lGIhFcrEUJy3IkWQDbdcWW425LakQDcqe92/nDMzlGaDHDEvqj/uCPO/ZTaRUvCJ8+wwFBMI1rGT
RbJDXbUb/3r3jUIoLL+vwY7vXXActp7mHTwDqWvxvdzNXvqTZ4a3qrc95UALCidgPBzwDHAmxwOn
qsL94+MtkuzBxc969RurJg+pLUlxvDyfYRkRNg05MyuRoEamF3uidqpKXfqgahLuUSYG8pp7Snr3
mIRrGDZbAMxwgUZ5rttjMV28beDyCkS9nRsnXfPv9v/sur9big9Y6VYCRuB3Xm69KK90fJEiCE1l
pS5g+E8p5kl4wWXbYzI3AYbZ8i3p5q9zGQfbdsvF4ZCvKKzii5q2VhM6cGGLjY5jJ0H7dbe5qniD
+uaR2Elkuggs2L556qlSuTxvgnkI909Dwx/bJhGIWbF7WUx5mvAaJqm3Or6kHK8URhlZmDB8GplF
OOuz0geOrOzQpUrZclv2txz0w8DM+ior1RVFzQz7s+8NO8qgAsyHmX7SnotHHonZT31NHVZsIVRb
aP1bsgZwpbfcJb7p89u7rJsIBY9sOAzESzGXG/aViji7zICDu4SNOqaaK7T2jNQga8LTeJ74sCk7
1CqBDybVGK8SovuXrTtHuKTjpjBWPC4gum85AA527ronX04tKv/4E59hB5/p5vRwUkbYC8cVFqmL
c/fk2UNWMaMwnEA1vXLAGOPk9uUMdF7ma/VK//wuQ+J4Y+0ZEn+hAiweU0lPLdcM0TSIeDcE1/n4
WM4U3j26TC7lNVL5xP3Cso4fBsMiTSfEjJNrDX2Tik6jPoiRskt6medRc+6RAZ9Jg2KZLLO56aty
rNUC1YoGAQIYG8paYDy3PyL5N8kwmKDbcY5TsjI5NA1IoElCNXGAzvxkDWR751HrZGUObtYLmpGi
I+G8uxLucuQdXPJ88gQef2I/OaAyRp0Vuv/8xXEsFkqz97p9sAYexyfSnM0Orc1MTAiAMI3CeAJy
JUiIV+HSDw6LSAsXKxP7mwzStznUlVwZtsMxT9GRgMPqKW4EHv+U+8yqprGzvOqhc+k9f6JxkLrZ
AHIl7P4Z5/HZOpClhgd5jqd0lL7gbxu2c8wgHo7KM8LosR9tHHOaB0zLMBTWv39p8amIhHHn6I77
7SbNq75NqS5JHFQk9seAKvu2+kqzeUA+oHK5ONGLXeL8zrAwFqkR04SKXFkhHfJY+xT6VhoQMDRr
hKaZsh9mmirgplzG7juHS7a1/UuO6PGmTpDbtPJg9hgu0gGn1ruZJ/oXazKOJnNVTj53FQ3LUN7n
yaIJFPAyvOkGPMTQzwhdcgTNs2JnF9GyOmgjhQ8vcBfZBZFChraU2iik3lsem/NrwSkQRP30WJLK
8dkPLWWTGULiPMz8m6o3KCeMKinuwNolBuVEYHLfI5mcMEi3bSFvDjwnYEx0GChKlWetVuQtMrDF
yHR0vGpVbjntW0pLaz1hQZZQePULfZDgHgTZJInu8eD3JgPBpCG65cCr+KTbrKg0JHlCtQ9jJaCe
BMMPVkXXWHETPVRb2GGqTS3ih0seIa9/MfCgO0dJtnjEnRkJK5vNRqTQVxJmdPnrciFlmBSSZppi
Kow9M2tEiJ1ldkZ00V+PaSlcOsQqMXaHrycmD+nNpu62EOoZy5169c/e7u1o6g0fFFJljrUFxcZe
TZyCmC7EgdPmCklFbFoxKbpGOc7jXwol3geBiy3fG3v98L2QoB3hgjufV7NTwKC8I/S+wKGegA3H
dDM6l92LwWSFwMEijTguwzDedHp+9llL5EDm6+/yAfSFcQ1d/D7OYOHOYWJDhSHHb5kuk/du+DU0
uYZdUn9nSQzIYVwODpYAjdnl+cuox8g0JHJLhAA7tFY1o2SnvPxawDhkr7nhofFm0wvkWUvDpahX
hrjUD2NDYaRp43D3TUmlSxEnCAS4miUInW2/4oQnPIvHzo+aeZwVbYmkYB9f3ykL/oPw7VjBZafW
l0TqRT6sS0H8V4glX2H6FnyFRkFWCAvZWFeW6/t8X97jYM/VANFrz0koePk/rJhMjuPM9XdFfFwg
rk+ekfSX9XQ+mJrkUtJXY9ouZhamY0gGijVvXCbfcZOo0eB9KCWHPUOlkX/UXuXNJEvkz+Mh6Hj6
bFpUxiN2CUIHlTAHR/MZPGv/h6GEan1AAeKZUytpwDDG3rSSbPfdTRclQ8D2uDygublKDkLIbOXi
843704uBVHf3mgmAHxX2m920vmdrT832foDBJE9ktMaO1/Aj6eUCXIhe12jh4BQ9HonAp3dlNy+J
tTJSSfTU6inyf5A6M2jFsIsAs9sqxKRjihRMSEc5bvifjqsdgGIwz5oBBvoJiyOYy7rW+GeugxBx
zTHfA7p1ToKbe48Tpx7GhGrjhaKJogdFTYf0X13OV6rDNl3HPURhKXYkeYh16jIB5m5R7eK/0V0j
hG45UdQaF1sRNccmZVP4Ft/9jV6sZJ5w1wh1dWpuRo+GPfW/GTmEVFIuMk18CL4bgB1KHDLQLReP
2Xxrf0e1qw0VSt6YiG5pMr6rbRTBJe0PIAUIdlbHs0nrC/rSca+d8YyQ/2iog9hYspVk0p8Ua/wF
QeSOcaISjRj+WDdzHDC3yJbRfrX+P3yn9/WkV3IQmfbu8erNRwP1EghUK+EnxvFFyxgXmhamybDG
6Dm9/MjLkXR9a0JTu7UITIBD31QKwKN7aqHlRE5EY6mMCrZdijOsV5r5Jwpwo8ONjGE+SamDZVV/
1jAwSgsoA1T8mIdwxFZT9poaJZiQTmJLJhyijjuk6b9/q61x4xfKPwHbz1WgP9R1YIAkXA85sF6i
xJCPpkgCkGcMlYtIhdMIDxytVOqMqpOlVgFdvWbDOik6Xz0CAnU6Vt0Qz13PwuwEjJ7jOILlKYzx
SgYLCOZFItBWIWE/1ClVi/9o6vJ8kP+15UJO9HGU85fEk5WHBX63JO45B6uVWU9QC16nZ2YkVhVj
kwyaI6d7iGu+zhSsVc83YdNGkJG1AXXBxoqPN/xyO8ylIMzkomBCRaJAhX2o7KKVa1Kl+pF9G8Tt
1nADBNzEoGDJmYz5tA1Ku1zEualfYVq7SB6MIPFmzqzuefaptqahWJFx7MZHkmueDlh3n2+re1Fj
ldUytx+RYjSwssD4QC923h70L/CG/QqQy5f054fa/4Sd2jQC/D22jXsQVwDQpJ4E41Ef/gcvYPTg
teyc1BgYA/TanVXqQtDNqQwRcm4ht8/1+OtC5RuEA1iOoZQkZA8DIVswgwzylpqs2sFu1I4oFCpZ
v5pjy73/uhlGC1w6uXHrrTAS4XjieHSVhD3V4exKMhOGHTSHB2YiDfJzUNNRewcUsdX7oqa8lpIS
O8f9IzmkbDYVwEanmm3ioT9k8LtAR/Pj1yGJCkVckb0KrFN101T065Q+WpygMA38pcOEr9e8+48d
u5/yeKJX8pFjvpaEp2oXBvInevA5/pmjjxqw/0va6ArF4RRJUPRI+0Qx2/7uv8TXZlQpTJrVNV/+
2JEjcwD1UAyjnZk4Nw3clRMkh04RRvh8m0Q/jnRzR/V/KHhHyLv6JKS+gct/mu2T6MOHNRaL5oun
G9pfQA/oMzaS5KSViNYBLgMbuw8SSKQ4Nn73bMedpE4NHXhp7m+skg9y1T3n1Nq5XeN4G9Bt4ou5
Ef4OolKEeVOVQiI45Ge6S6zDPeWQL9GJBeBZ6ynWsFrlveJ198L4O+7V54PyIESMqwjnF1ricXE4
mMgqPOfHeNqoosjwiDUYs87dvjK1WTnzanmK9FJMwn0TgyycCOXFowATGCsuD83im6NtBRMnna1t
uERGvoTr7BK8aX+h9Z51Rb73J0AXp64ONBK07bXxaq/m4Inu0i3IBteCAgjmTJ31wSBpZDQBX3cX
p0dfzRWTb/G7BZckESOSdxW1aHnLcgAa2wZ/kvVFHancPlTUud5NDnsY+3T8tiXWgI/pjiHiFHFB
10yjfxGc50OZeg+eQ1YzPnw/gdLszvu5g3xp8l5HA+T5fZcOLIYSzM2q1yzA/t6ya3VncoNksKt7
aBywgkCnd02yTCSPMs0eA3hPjYVP37LF1S+Gw0TH7yil9YJC2fv9TJDDJyPGv22vcsf93DTFJ1cl
df1d5sGifPqwBpo/Q0kC+f8ris2fXHL4183i9p/DAARPXyFNeE2zlo8E/gKeFXPfrtxyfwBcIG4i
IzkVwbFLL9ZDGYskFnRZ2s/o3Gc56sP7sIuXTUaBNur7xGcZVQhgy4A7vwbBK+FRVwhfUVX6Cw3W
ZN9+mVuHtHzipecrCjSohkFvCRCsgMcwE7vE8cBfdhfW5yhS8j65eGuJKY/PtC3HgDmEEZB26pT1
jv3F5PH725Yr3Wfb7Lfnz2MQWQ2ttxmFjANn9CXyLmIErR0hsaFyhP4bozL0MDuMLih/drY9+6qP
DL32w5hnscxac5AoSnx5GaigHnaNjfr0pHrzzjRxpps1nckt+1GUaaPDwnGQYDP/uiPzZJDaCgPJ
uvxh4n3VWfeaWiwPakGrJ7PD+r61FCpZTzJwjvazmTfLCxEz1CRcNc3BbVBUc3CkDQE8Rv6+T5ts
Ws6aT+4J1JzSi4bc9HdoTB/vOKROZz77b0iC8Bxv8NhOlsfMetklo1C3GcROyzifUxFo5iSiRVR3
WVEyc2kQAJlcO1Yad3lZzQ7sic+iwCD7rjFHcJUuAgfZabo3G4/k/k/ExzpR6kchNBB+/rlIq8eP
Gyq08RFrqd/YXX/RLwwgRiD3bdkfje7QfQAmVEDbmJ3MKajy3FlDkRjUs4FhNcKLWDBPahONQXGp
mzS1p3mS5dhqevmJ4ldziH7g0agEXd5JG5AYiHWXAQB/OPKOvpA7TZ+zum0Tl8CIPqks1ak/E4xs
RKG/Nb6n/dkicCvY9NhSxJg6HSlL2xfz5w0Nw6uOaPjaK8KdZFD9RT+PClJDEPiihWMIlhYXhotG
57lOwnZrvgJjuvmZOJkNPsIqv9SaixKXd9eOzN+WmmHxG9iInhdWlxfvGzrKT0c7iycTqK83ekco
w0fnq3tFfRpEbMYQSuAb/mZcbZzfQP3paXf8mNpihxQsUsO9g+WjIFfqlijYD/9+cmozqnvg6OEa
oxi9YNFDhWDNBmvTR38Z2/ZZ8n6XwXQcOGZy+IOHgn2Cb7O4vXj1671Fu8iINDCCGN1NTgY6UOJQ
lBIogx9ftTqm9b3VdQUV3UL/ODcsHqHcmJmbMtgtHSyR5BHNl5zkUcsQYnQucuUKyclhp2EMz4lj
It66/OTJORIvpg+yGmgaHnyZ4uDMD4ngOUhsaXZgGrhCio+ye45o/JVXpntgmCcJk850+QJOqo4Q
1br0hF5nb+LIgN4Uoy2q9ZjaLWnCIBEXpK3Iaum5aykppp2YkWXHjXkCb3L2I7Kt8G0QIyWnhCrC
mFzRR4v0AjBoG6QVLOqn3r/XQfya1k5qYxIcqkQ9B+uVnW8HKA+s8zKfjD6F7arlqzAN8CdS3F5S
nul2ck3/g5yoICzYfRdAl9hSJj9vXukze4BKoLpFDMAuLjIt4ejnWtCWkn9DUvIpJTY9pcWd7ydN
a0ssvIYdtXRASIDTldngWj4/90rGMz+cvtQGhyuEwP21xa0bhELo7MrgsyAKlqSMVFE1HhLZnZlW
yDui6YfavKKCYq2YRSoPTzDSAiaYTLm99mkuoqWfXusaxicGt9J3jXq3TZyEA9a1V8p1+S7Bzw8K
1D3oh2BuY0RSvjnfQinAKWOa1J0MkicKVLERlWlW+US4fQp2NBEK6jxZFDNzKG1RFMfzcjWTc1wd
mQqdlAJMVRKbQwY30uQkhWVT8bWAb3RE6963WiVNTB4osRs4CxIgM6KmEN3WL0IMVNA8hcz8udNz
rUT3wvg4eKpCzvP6YOrOjybpma+/I2TzkDl+950kqK3+D132CDvJ6frdcAhxEjzXu4i4KtA9/JAD
a2Hpb9HwjzzDAiNoe0PISR0t6hbRdOq5t9eo6w1qwKLRe9YFPYwD8V48prO5c/34lmRVnN6q9mjk
IqCDVT5Cx0xTk/F+FsQovZLufVD0SqFtaTpCle455ycZsPkjRxaTo9pnh+iFN8nzngpDKiDBGabA
HWmThyW0E/dP4oxdFqk2g3JH+CiBXzNwbQyeo/3NnRYd8KvyIV0jzTTVD0WZZMTtEOE7kbWXu7GE
nC1bPLJ+yODK6EVHyvrTa+OkkltL9l3BulWFBm9a5hdsqSFouLRTDsiEuEua1vBJ3bzN1FrzYA4b
QzVO/Qsl0I/4gImRokYXir9G85pt1SY5xGVtSzXpKlyLdX06fJKVNAZJveqtBJiHn5I2f458bFGn
/NiLYcGeUHm1y65ok3KzBVU7KKlQLFbJCDBRU2Z3cNCbwkfVulm6PeKCFMmb4QsQQTpkfsIPxh5Q
09OO4YXVWJk9hFl8gMQUwzOnQC+6upUmMUP+0FdNVe2Y0djW7KYTu5qnbj/edmAdFLlOFKlax2Bm
GnROP14W+DWtE/dFNz7ruKdGUW3dldV+Do+87FjUewaeN24nJZ4lebBEtcCvc55HzIInTxJHpWvp
8dkuKvE/PW582c69v9HpErE2OtY//L6gij1fP+9oCyj21VH5uDIwHojAUxd7i55sxz/+jKsHxu2X
xV8JXvxtdKsld9V5X2DTPQJ90rE3pYl2OgevLcA0WOyi/O55FXJuWhRycOP0pNW7qPxz4XuWyDaT
SkAir85rfeZ+RT9EPq/tb8ErSj3uJgG6lg0LGm0diNs8cPuGpIdMHZG/dCN9vUQAvgPMVI8Qol7q
L3qVFx5g5s1AU6WrZP6i0tYWTgxQwv5AIbmkoYp1+wlNzuGzXS1Vhjw5ohewt66PSs+1LEqOP6nq
fD34R151D0So1cgDTjwCGMcfueCRu2f+X/2o1iEJdD2KChRqHqIIv+5x6kkCD2Jbv1Kshqzc8OVA
Y5F+hVj5nQw5iWz5siG9rOAGWhAvbj/FmMqwCjuy5prlUsbkKyPDPikwvJfZcQ6rampMeABS0BBr
01SPa+QugV74J8gLmhr2EWLLzSLweFQx0GjHE7XjY/MY7mHIp8IzQdCviVPB4SAuHIf451t1NFl3
NGlJDZlK1hVfjPIbm3LZXItvJzSXIvYVV7xgizDiT9rG2efEZEAYlzkcTqXB32aLG0I6/7tKldEk
hBdT0D+QOA8mCOxRj4o2DjNEQrBasN8RU1XpZTnpg+uB6o9Hm95PrNQjuVtdPHMc11VWsOQfYaoD
34aCo89tIB/Trw+DzXNWt53g2P9zBqGZFfXAuUcdT863RW5YCsd2FNUIVVHKHF85446g3c6Y876M
/hUh8sGiBc217BKzLxd5FL1OJVpLZd++gBjJ2qWep1fMByWZbJ/D3JnyxTye4Wu/z8ui9oAqbXYb
9JCi5vAOPIDAiDFGMbfs/wBUxkl0D0x38cOaTQKacr/dc0aFEzgMo2Sody5E/AtkDDwehuDPLb7k
qbD+Ysu+0VCLnRNdqvF8I0C1P3UW7ycUE6mt/36wRMYj8IfHoPC5R5hO84D0ibWJt2lJsOSv3aFB
nodmsvc8ojY3v8h6Fbt0FyMFk4BAaphTPTRbmir0HFOG4zrG2jp9G4UpIgLdWuBKR8AP8vzy2ShT
+i2eiXTR+KfhInVGjvLDiB1wsnlbFo9daJHMmgNDUjQrIJFfvnCUY11ZP08oO8fhYSU3c0vXafoh
ueGgFqC/bK/9vNl0ZzmqGISbA8N/HB2q9bH81vngs/yikz9kM3Kx2MWRx71AzAJaEtUejgeugqq3
H4WvCwuR04u8ncQ5p3UAeJFl3eDtbZJgZeEIlnNrd/oEyU1eD+W+aWkswd2NCpZI1ma9Gki8VVZV
fviV5LA0xaj3ZmBGxq+G/x9ZyWb+/IwmxYJh7P7KLTppvp0P9tp4V/4/3aZLSphfw6P0kmfMRVK5
Mej+pQ7pVQ2xeBcabZkKfCxeU/BhFBxZbtfMpe740QvTa1dXNCTmhCmhcagDjMEoRPXPAHEtooze
ByvyCiwY9EA5FpkKfJx85wMvtGnkhJSCB0I3u3lxjTBZ+qeyk6CuAlJm5we/hXhojKK6gVGru6Pf
auPcejAoNN5nXSpB5IorK0hp62g5WFSFsL1EqT2681CAYkigSY1leumeU/qnnis90lg+NX4Jh33n
Pq9TEyZeoz2uGRfA2qOmupt+diV9UjmbBFNZRZNFlxC6vpZ9OF0Dk+DtSQNM8yWXPwBd3TVdacNr
JvGzWiUvF36aX3wnuUYZcXMUb8gvkIuUKvXu6bJhYvjI9/ElmMC0DctOhjBxhv9qCaSZR3wr1bnB
jMIhPsz7OQQsFnUQLjsjTlh2PipmXUZ/OGEORB3jaiGc7puUsa9Djiv21GdWClOtz1WkxKI2oFGk
LLYhHgo59KnHC/RoKmYq/BIz5RALzbRiZHwDUOgxeheNrdKtQSVShwH1dd177QhE8jWnQoooVM2q
Tc8f6iBm24nUAGeJfiaoJxwWw2VONCZgflgek5/Q0ybbYWmHJStoGMo5Sq/J7n5MYJwBg3PaBySp
d10tHzrk2mEm3/pdr6LURVy98TXIyiXz8a/3mzGS+vCi10Ce05zKX6Z4RmPnOr1aNUWrCpWS+tVi
nZ3Yey8eavSxdVF99zNmTrH9GDM1NxeHk7MuiJWxp1/xkyqePPl1pzNAfulcZyctDZv63taajxo3
qgvK++35xzRSzUf30B7jjxnfo8XblgnAN2idIdZX8RoxQTIM8Dyaur0hkCVHDSbTZ8cVz8q6J2om
0JYmIQR5ZpXi8pLFMDoltJhIaISQoZmXlwLZqhC5RTN2cx5y0FMYO1tZKJ5feWUKx17LmwNBr0G8
vCsUjFQ5dLbDueXkEEw1RlQ6+O81zLXrg0W/61fOS1833XDL6QRoFnhx7nLo1kzdYCZCke+lq6jU
tk2v592UKjoN7eBQ5paxV7230xU4IGgtb7HBRz8gGWqvjKPtmBgatstGzPMcCW/e/7778tU82nNa
W+tuhp4IRj20rTd6oUR9+AD/ypcWHVpd/Mx+gBXjNncBP8KbvseMe976jqlX30YlRCdpPK2HLEyw
ZohxiRzcFGA/JnUL6Pie9q6TfUbWcbbucW3Db83rNCYrQ5D8JkT/Di+6oUrloZ6Yg8cRkMkJFDS2
w3IqvED393DR4CfbnyigU+UIatJYAz0fZK0rDeG88S/2JsBPuVSJB2OyY2FQ+p3W2g2klI1GyYh1
ViAOVc0VEA1wxjTR6oNgwdt+T0h5owuMa4Qi9sugGYQIoWnXI2ykkdEih7unTGe2z3KdgXAskMOl
mrlbjCACJx+IYn9K7YfTzdKJH3A+w04hZKl7PcNOYpy5PrN9bHLijmh6/wyRVmT3/B4Oz8rGS29U
x0nXlXgRiXlQ0aR3ky6QHUTSO5NjIk14YNvsOrZ4S25uoF8qsLaNxzXrCE6wHf9rsOVGl1TKlSRQ
j5eLlIKDdYWE8g5LpCCazPg7yy+KdlIYA5Gw9E+i6AliArNGela5DSBy+HV1k2AzygFNQo0yD5iu
vT/Ztr8mG5Avw8H4qnlgHCp57zhStmFqmGuP3vy2f+4nkyZvheS5X/DP/SyC99LQjVI0TcQ5LEjg
nzSA7yjbabrqt3MlRyCWSvvwpIgjinAt+/u5aHw6OPYKQf3EF1E0uXyAud6KNgaTHKNzeWW7SjOk
J57PfnbyDW06ThbsGYoqq2WOplqtGlHNwWo96JGl5zbr6CcX8vVcejZmCXsvlTpobD2pBNkaiEdY
uT8+reWUOMFuAO50L2FIQDrJw6fTeTt0l6qL4DjJXmf82XGDH5GiM8p9YaAm5N3i9bM2C95yRwLl
mG2i8po2odtN4fTc7pTGczjm6wl5ZKuhp4bnis0WNv3n98tS1eNb5gV3kR0oeRrWmtkoHXLjIFlw
yCMf5UJXhwXRRi4NTFAxBZ1qKJItgdvTCk+w0pd69u9Z2k8V6NdpkTV6xG7IU2mSIP677KZlnydN
lyumHovxWYDV70GEhwAY8C8qKQ8xWqgCwrZfgMb9EYkN9pxpdqtSaF8GZoLH78wITdP0TQqOxT3k
vu0MH/FDShu7ZWlTJP2K9ej3+3QatTVxz8lFqai2cNTHkDMyuIFJ2Hc56IWHnC9gW4zV13XoRW7a
kdS3vipw+D8FQZ72rJBqON91R86O55Z7m4Y1QpFpu/um06y2TwWnS3IsIhe4M35YiDIHgJB1yE30
+5oCQOatO0WBmNWdTanTtc4Jn3Lro/7DgoXNIftREMq2d3B9cHW+mA5r1VNPBO+SA8pXUXxTLQyj
cGMAotS0HScRiDpPJOhmRErW8EBYKttN/XgddGy8FtdfysqYs56jXh/g9E2HbazDDcw/Bb/0uLe7
qwWiCOjx3cCA5piFPCt7dlBdfIDcXvVPuDn1x47tNmuM5CSSjnm+Uu3hhjjcpn+udrKd3w7Gkd9u
m/+JKtmk65N+3/yNRYnhJQm90Q1cB2UUkFlYMtiWgiYABndJDPn7VkI+xRhFhEI1I2McDQkm+klH
RQwRnLqQCSl1KPEZsxnHJleE5SEK7x0CB9cDwb/tLauGCjNOGBnMwGz9zyvPybyumB7um7iK5ZYZ
I5mLAziXMz+RUGEs3r67Xpm7x0F7BOvrI+pJFtQSHsjMaB/EsB/LajEWbuAIpGfnbigFKLNWgL1c
jsdCTa95P+icDWo4s2U7E9MFHpJ1O5erBb+11LcxE/FKCM+i7cGQVrs4A2sezrV9xmClSLkylZi+
qo8zuA69JOdWzNJi+ioeiYIEsBgTcDgBMeEZL9XsMXmRSmAEJtYOdI+LmBxF+jo+Qu/4l87hsIEg
qZbd/BlHmKdm+fHT/H0cLHchrb6lwnfimuMJ1nehQdqk+hxjBTjmEhjRsqoMdO3gYObRVch1cWUV
AgmRGLCW58VzW6COKwRNlIJLm5A/z3kPBwb3fMJZhbdzCR2pt3ZpvHtnjKORb02zzATXG4qwD+eU
ooLGYzAph1y1UIiYjYlnioSYATJlye2zJLUMvQU0h/z9Tt8ZI35ColXbzgOYbUEX5djn70zOP1K0
WtSfP6bmKOaArBR8V48YtaRyl57ypnbt66K9/QXxsUF1qdNPl34y1yOQhccrkKmyN1P9REp6gX65
bNM/VqNaCAyONRIbkEbO1l0u8thrfaOGW6U9VO187K7MWUH8iCK5BNqhOIyMnrGolrr5JvMHX9Nc
+OLtH4LT7mwanHvvAlUQRw3EClKQn52nuB5fr53wb80gey0Tlmm0IfRfhvu260QJpbiS7D9upu8i
58XKFw07puMep972sh2m7Kz9Bs1aOtNTWX1gCFz5StsZxwat/yRJgbtsB85D+JqBHKwEG5ge3qgh
S0G7RJ0xTcUBOhvHi++9C12QD1IgymNJEN0lgwLd3L2HXigUzUy8kFnlzHrMwE7DY0HYlzxWHkQA
8vjqk6zti1r24vjr0Us9a0wPJWpii7rdSoIjU1Tlca84UMgNNahWIRXphuKM/BL3uDenylTTqxkZ
0A1cyGTK4psAzXNdO36BNx8vtDv0VuPIDO6nAHLCGY5eYeFh8uwbBqaBAuTND/wXULLrfQG991Fv
CuKcNrt+RDusy1ZG7gKJxP3XT2Fa2XMEVqe50Eqaq36GCrJ2KSxdCvGHyZJryegkDNnT9507s4LY
++1uMFp1xULVqNvxAH+ouJq9vFjmx8B9ESZVtdMrnxFf/WzT7Ew35J6I90q7bLQRv25B3nm6lzbO
suggZhCDyLEXnl7pBC6YJ1oSJ+6nrZBdii5YkH6gWSRa61XY6Rn2PQNx0F7T9X1Kzgp3hSDK2lk6
m0YKQOuGsMg466gg4gl2KfO1HvjLTff0N0xNFE2pV9Jt0CvjS9srdWcSirrVbnsBbiWcRUxw3Opf
hGfXXHAKSO24rR8XyhMBmoM/4j7+9YyKEM2RwwCOx1ajUfiyoYO++gtTetNc3JE632kTU4GgWfc/
kEKl9z2s2uaqNc9YOkWS8Byg2RErzNi19tGslcq6hPe0n133puVt+9cg17AYLBaMY7cWv+HVlPwR
c10RbAzj1EkZXBNIWJvMn/lrX8NbNZtFd3Gzmxmz8hSEi8cDp2XDzGsIKpQGDs5XoQdOApVqrxmL
ZgBGXWTPy9z1hb0YlM+H/BDkqPCNkq4OOdwcsQVtUjLzG4tRCOkbBDwCt8jGSs16fa8JQVfBrIt+
J6F682K7+oOGL5NUJddNJK+CJfPX1Ajy1zw2HFbIYEb0EU30ID1BhrWKU78yxbKThiBwil7EuYxP
jFQswXGycJtRs8OfQY04/GAhE3u2MJwBs7f9v89QACtw9uGC9D13mu6YBEUWhSDSjUcvE2PrE2m9
/Vt9nC2Ra0ShRiSuuaQU63U+ZBTQNf6GDAkuI3oxobdTAM1jYLm/cUvNAi+gMFrk0FoGhqyxa+xp
fNBTArUR7dEVAPpQUefCprSp4dTift1wlnSDbLx0dnO4GD90osrPSd9UFNWpVistdRamngQqg6IE
Fwl6GS87xEX1rLR/bdbeRn0gYw2cbGgyfPpAkoypddFHFnH5yNXZarl7YaHPZt9csBNqzHOKtpWj
H7EiDAX2I40xHB7Ji+vRtRbmRVRyeUu4Ymr0E5O53UeuTdwIXZwHOQq3LZBN6Tky4eafO4dynxE0
j1Of2WFda7zJMR3iI/ZaXjMmlW+7kho0kml0HR87hMmFJB/Um8go7VlSM+fUEapOrKf/8uKSTpAW
dqwTwI4/CPZWHfeNUyKInUYERnkJd5bo0agb/ZIWMk5VX8DjYVHExrcyserpO+ecWv5TAtpvxTXi
NPaRv17OoQJc7RY8md921BSIeoKk2I3Z6y1gYrTuyobmBM5omCB+CLLTGFn6vfJHlPQ2BdzQJkuL
unynmF9kA7xNRLkZ4kLn3zk0OK/xDC4NNmfVRjg1Vg9pSZLnsmJYQ8lovc11ySC4DGyM9tHPNBRu
dtEyikYx/e8cIOKuMC/0wwBhR1z6/sr2gF+8hN8v7tlQEDJPi2dEaEqbW6kwUBEEYjMtE/azfwCF
pwuF42VLB0O+CQamlYvQkbac2QomTw0xcsxSP3qclGvGGCA5Zv1Mogd433z0Xa3xecKbu2NBijNe
p/w8DaQYP1IIDkiGtyEh09geXDOCqPn40vowlqiltJFqoEgme9jOUvlqrL8mJ2ELvOVAKwlEcAV1
nreMqRTzMAsH32vj2s2KMiYywC8hYos8lq5l2veUj37lKN5SWvPHrM+Joc7jVGpDCO2ACjVk1oUz
3PM/omCkNGN+aCFMqFNQ+ernrEa9FPoML9DB2WMOFOxHoygcH16ky+aNcnC3BVQ72xSv2uTLPuh/
MVosstfl20uwmhQtqS+9BO8DMThhhGYIx7ZldeexGJZizPZuGUF086Tycw9ud2QA6f/XRbBjBMwI
3/aTILwdTfJCawJLlXWfl6PsguU8U+pxE8h0TccMcZzgr6ezpj5iMQ9h2QEy1t/q+l6xajvnPpiu
clHi6MgWG15+q+FLr8SnvwVNjw/lmOZYXowVtTNQxMbqsF0ZHVjNv5b4LMHVWz1QWeXDn2PJX300
tuYPZMoRgDfi8oTIMifJUeq61ArBJwbu9TPCrwvt4+DwLGqVJhocGlWwhQTHKroIaWNA8vMATdQI
SRCtfIZ5fTLr26ig3oTTag+Ouc6NPW8j10W1WBeyxr2uAKdZCcBNdp7R463P7TPZP6ofRy/vwmCD
M5xCOZ+jSMZCYl1NN8WkgrUBPWszMSCXnI7aDb9rCZTKT7vi7hCKL9wzATX7bP6l98655vywuQDb
aLqlcfb0sx9f7GwTZiwB+gE8MQfawjRGZ9TzAmlXErLml12LM8DowSPweuLHS53BhG0ngAvTsHSo
947Vgu9oWUInzOFeE2Mfyq1xg3ue7TlqoeMxXAgOgstPrCroHQB3K3DHe2l1tlYeSaBEmX5nyiBg
EWa/Ep7tRCk0ENwZmS3WZwBBRC6xWAK1OCvT9T7c8/vuJYCT/PHb8pVF9OFjyktDPqCTJlcSgSAU
zXyHhGUONTu7JOmxY4lTtiacCoDxRxXqpHoOFCxGk82neYqrogjRU+2Rx2aL/spfwi5YxbM9ETVv
MFOHJIl+Eh35CQ2WaTHUFNRedfW/INRJ6dFeFsjFLL6DwFidOhYZrZ0+h3IPcw9owouwT9TWoyU+
xZw5RNtnELf8GBvuqVxpyh8HDsODxBHqduohWHTFZz/YH/1P9uoHA05Qd9oSNvXdnGmywcTynJtj
jkMh6T+eOV89y1EkvYatE13xvXG+McR8BhVqY8EeR2bgSOCuaAaZ/+1RDoAO4PCY8CfETP7TJi7I
L/6Axop8OkFA+DzyX2buiJYbLXhhtkDIEQw8FeWe19Vtn1J+xYZuSu9Vg1w/n3BsF7QBPvUf+m/8
nfvQtlWb8J3VvPSyFo5wHEO4thoZqm57Lo6v7gSe+hZ834YAVvsV/6tdxd5S5TRG3m5QiPcPaTof
fsWDxd2c1WVKqJsDR5fqPAbvqMQ6PRda79BApfaFfA8OIXKHrn6iMkfjKcbFSwKKpkhDzFy2mwSb
wnn1ncHferTTAM9sFXU2la5t2TiIAGuUAnOGPdXIt4lTmEFWJ993eqWpeRS7AEWokusmY/DikBNz
B+FhOxdk6hs0u0xR/SpB3T6362Gtr7s9kwZyaZ3nT2aTsFnwiavirCVOAAAQ5zxzIW7kurLjntiQ
sAJJQjdfZdba3Jqs/MoxpW/keaPxRGgDiC9Qa2qJppbNrfThYuLBtxcZugeFN9NCWT6XIkYYy843
zrHJpQ0OUM2qPG2nM+INEDoPDxlmKRLS4OZZvA7o/ieD4OlcTWQzi5pht94IRR6fZJqF5fqyeXCK
kjSFhCcHOuHm5bMdllioozdoQTSAlaS0GA05P/A3D3kLfrQZ4pMclFSxVfyrTVLCYAxv3ikfHZ6U
7ZY9T9aQUqpLq2ezxrz/7JLLLZjr3nQIJjTJZWcX4rsLx/PVflC0+zI9gftNHEC6+pn4mzZD6VAs
LUYxZpMH+ilykILu+W460vo6LOE0PSzsDXK0KgSdeT/Nj8vBZIvP2AszAAng8A5rXw90quN50j+V
uPjmI5H7i3WiqiMdC13nWGKOBWdtIRVJWwI+CmByA/VQ9dXkl9tOHVWYJfa/jkilWSFU4QteX52I
5B4cLtcGClbGxNajfdwFiFoMtwYQFdUBZC6uOVnOoO4ONqVPIwQZjJ/tYSaEWqDDABodd17dFquA
hamUER3nZ9RZNf2BhYQWavsBpPemXjOGUlw+No1j0EHbcfOATdiC+p9bZGoZJa3AGyZ7HRu1sCIn
qUtj6mPZiDGJtFSHP+6n/hNzT7j/Max4v0ApLAsABJHNgw4mJi//4ATs4HgH8Qo6++GzIPUxKE+v
p0P5rkDRMXYar06bFz7vRG+T1smo3/H6WUVkrYfxEGIfeiwTjxa8vdnC4b7C+ebqaPlhxR4IQBqu
3bgjyC3ZNUZ2BE1aWko+ZLVe+DBmPjejA97XzKZ0OwuQw/ACKPObfDT6HAkzi7661q8CBmAOzUZU
x0W4Let7TH4Gn7J9HvEosOClyDF0j76VSkwDxFt18vU4qLzbIyOtxvYqMqJIj4XkHwUIQ/+vCBLc
aOn0/6RQ29Qw9415lLc7ScYyjZxLfkOqUz7CUQ4mrzRZIYpvbdG3mUjUJIfBgHBhErZEoXJlOLi7
TIgXD6OK+sREOtxbXLxjxQzZfjZ8kwAW/2iFDo1znBb7hYNMqsQnYmBAfcCWNaTfFwWgpOszyclf
eM/aK4PO2XIWYpbaAFUTWJt2WF5DJXdlq1zXF7hcLZbjQQ+QRn2z2ckx+i3wCC6iMxdGsZAXt2ok
+bAozftpgaEMak+HoHAz436q1Bs2RoX27qyr7yBR5vht+YaIg7oHkcEOa6Bqt+Jr3TKyox1LZ69h
vsOvPY869zCbTSCr4omfxfERoFm1ch6lELRuFZtt7rUOO8f8Rv63xNlDUhew2P8R9mTeXhfQnahR
y4YtzFw85pm3O0jnabOeeaEEP6hn1TU7tFi7mKiJ18Q5orZ7W2H+uTGgoFpoxQqGnyrjN+LWu3SX
Gor5S70uAOMuSHVJiEBcDxuddGQbhq+8EzJsEhLjSt5bWFABPwLOFLfDzvXZw58igpEIKUW5DmXn
MWqvB2Z1rVb2EPxAOcVcSKngJaDCvsDGM8Llk5E1QRrmjeI+TjYRleEXrJEuqaG8goRaj3DQJid7
Hdkd9Z6rLT9YhkJv/NJf/8RZWbMnJYvGQ8auYHfxSclGfMMzgn0J7hWVH5y6bsbLs0lJzwCAdYVj
koL0l2XpxLNPgv4NJbT4S5A7SXAO7i0voNKS+XeRpesRT9qvkQq4nMlqJVfjeP4xqZa5g2+hgTz5
ixaZNXJJJo7lX/jkH25njS9+brwPrUd3MOS3Sx3wBW9yAQHbHu7cl6o565cOiUu1cORXFTHNFioE
rmNmqt9Xn6RJryIceP8xBtmV7rsNp3JprTZS89/kbeOu0WuesZC6iAiBQMKXuNwJtgTkXr1cpuYj
BklM3qI2YDe8HsAZvdysnRFQGNI56n/ETxoh7s6dHRfSmSrsbSB/PsXJvtZflTedNaZj1enmagZ/
iPWXBnWGMlKCrK9PRY5jEW5VEqm/UyIDh814Qom8+shoeG27bNKc0Ob2yp+OS9Kg4h/T7DbpS/qi
4mXRgz38WcktyzJ7ZnC6uHCNZKu9f66Xw1vDR2c2fQehSsoB6A8nQBrQ1xEIKREP0kQegVfjCQus
5dyausiy0yRu5/AImhY0gKQmk5TNv+AL646U5NfMZDoPKdDCSIynj0hPWuC464KFvK0Sv3ikgYOJ
XmrA/uetmDBr4yeKeGwBX+3PiZMqynuCivorPKplAW3xILPgaYL0AUZn14BY2/NhscvyZP0VR7hQ
YOMtOqEn85v7mnvIl4bljiEkHtvCWBlMQrFZlXxWUxZqxyeGZZMTec0D/SHtt6EP9d95yFLF5JbI
S6uxPLkb1PJ+PozrQssHcW8p6yL9hdCfvFt1yO59cALJmywF+YW02A791gtu2qiZdBXKWwd7BERG
0/DTg+JVZI1kvmB6n+Et+EBNKtBG3lE1GN5eiLDof1oxggTi9uMDFi5saYIyhuQtokhuVJPbMclz
IwcLXtqh5fHeWdKgqaOJOTq+NOXM41Kulf/ckaAv+sYCWO9Iug5OXRNOgLEqrBisqT3simj+Saas
0VGsvZavVP3ljfh5gggapdbEtTFswHyc6OLlf1koWyk2Zin6il4RXxC2Zw/OVFocBwCXOFdAf2Ly
HMmwUCQZJFajvb3ug80Km030uOZDSzFVxPNZvS9KGGzb5WzK8cNVMy6ghkc+srjcK7/xiganE7FF
O0OL98ztPmwFBiOq4gGqXGnsWqKfr3cOD5CV1Ypl6UApst03rf5lUgL/gdLay13DXoza+BdD5gQt
JSC7QE6Yo2bXnMNN1k8OP88PGcOoAE2YMThUOu9WcsdWIVdi2iDejSAdRx5rD1cCPslFgoo5C5MM
BKSz2CZCe6e23S9QIWaoV2ycxv+tD2QTRWXQHmVkiG7O0rn91g+uuXs5OYLl4ixW8L6M2UUHoEeu
7CVAyHiHAnPidzrJTAiHkxlxWQLaBQolLLx+B7kmuKZYhP80Y4Lk05i+JztzVV65nCYSDtybgfFR
vmB+TGQkhnnCZhi+khLLXTBQ3I6N/9iC7/vbP4mD2Vdn74860gw6Xr3iCkn32zIu5HgTWI/wPYDz
vtSLphUUanDj90IK22Azz34BVctympwD9TMtivsDdTk/haLa22fvKz+RYO6p07qDA3oAZo2vcNvH
pr8IA4RxT9/PM9tKd6kjqPRBL7BXlhOivPaBD2N4LDSWkUYJL0O05J0aeuKedIceMHfzFPbIT6+U
dVoGT7fL/JurGKkQjCR8mEKHWIpYoyIv7bSUEP/PZHhXg0DQC/LyZGgBeEVBAuNLPg2c2MOqH+WF
SY/meLYbFPp7g4YerXxdni8gNu9ncglfA+dqolJJyB6fqu14ExDj1hLbaZJCw+58ml471tfp8avF
MZlPndckqzmpcd3i8kyAZs2AFtT8uAkMDk9RNN7yaTBkxUFxsF2TFiS1xqWSCsqbYzCGGaA1m0QH
xvCWDPpO+Zb88c/D7ltn6rBD+0i9rUSoCuu9bfwmYuSo3R+aXYY5tSKjiCxAjj7biIv7Ka2vlql1
jtJorOswclxotc/6MkCETZDs5SYdnzhGPIV4pCt3XIbX81WBBTURN0JntG5tHU4DeWyk0qLJT49G
Y6SyPFHHHqDj036+P9SxPNsXwF/xAcznqT7Z5+XvoHiw5/ld2F7p4wWsWqEdyxJ/fEvOT2pZGmr7
FxdQCNYkdnWT2+xsK4XMMoaCVu+G2TWGXkWZKMqEmKQ3dsKIa4FM6NnlG2ijM/k4YIdbniCIwyHF
im0EM5MZMWQo1k6zd29M2jMoZ7fjNs8If9omkG0CT1ACDMMSzey7d7PX1a21d6ACge0BaL1yEdzJ
LDLLRiqnu5zkvrl3cCd7aQoPdoU6ny3mW2jsPFLDdDsSOhZQ+Z6F4mGa8hXDbt71p0Z6Od+gHy4N
V3K1iLS5n00kRf0m+EXzFoy3YQ8HsOBEoy2rRQHdxxvb8nK3wYvifEb5/x/WjKeUDzmoibwERxFk
nXY41xeSW8pwu8fWbdb7DdaQyEE9JeFYLXZbFZWhFcFKj/Ri3rZ0u7dIGOE5RX7TlGw9XVAKZ+YE
xxk73N3IK9HY8v0qNPh3dx08dlXMdK1lgdHZe42BtuaeAm2yfDsN8KU5vOKFZNgeisLKxjOYJlil
dYV0/Bm0jP9yH4GR1aJ6r1OGaBnZGmG6G/vYx84mjOsW2i+hof4R1lIkIviC5zRHOZyQLAxRmMr/
KrATgYnOekyNQtW5nM6HEcSQBAT3LXaS8eMTN09/bKDEhJguZNGl5iJlLWGobA7u7Ji6+DkG+X74
l9rb+QTtI1gELGu946JHEC+RJMBC7+EhCOK2wm/fmWXjbVUfRIFRoX/2X+hPE+/Galj1Ih3MDtjz
+GZgyYPyeY89kcNnLmBWK8uErrs9nkvMV3cTZR7Org/lxAMg4yEbLsgY34Fhknasy0zCOQ9gquxj
/wk4uk3grgy/aw4yw5YThVtxdVBy/m3jVRw2ICgReAFaQGrOpk1Z0yRMLmkPOQXT4ks5jPytSlk6
yBodU3OMalufanqbZcLreropTIm3BEHf/Cx5EcJkdYmxBqhO9WvW9Ikle5e4mCqLDDFsorZU6H8O
AmvTsJ1fbAtzCyqEENvyWKujh+CR39DQIu9YfNOzpZS5PYmFNnch3xEQpAU9y/717HwLP9uRmMHL
sua7KIj98LUQAOJgqgB3d0X+X0GF8QMKU97NCoRBy55sWsik9wpbXL87t+DVDIL4KkNNqWjMIMB0
F+OLapegcnCmrBjXeIukUIDSyNhY4XILoUJnYLKabRg2HCezJFzxx5mU/NELNzU6veRQUMAD7BWS
cHz/YFjLfQro8N4U633J6LhMdR2MHXVsaC7w1RER0qyguAut/JiQjhCrQo3Cr453kUR+nwY06Or8
K00NPX/HHoFGGQsWYlaqWaPyfT+8X+V6JJiyQxD/crp0HOg9++ycXZ3s4qE7CbpbmIHZvhn4QU2X
Bmq0OXnQ5CpC52OPgxFFH2tWPCwAbWmwm76M0HA8AZL/wRBQhEav+WOWfkDyzc/Z3hHbbkkK8qIY
xe1ZZDSUBYuWJCzHcsgrY1QHFzpxKmltsERWbk+KsSVyOUsmTKTl0mAmAT1j/nI0H7wLp0piVC1S
odNhpL+k1vxN+J3eTA1qr7aMJLVORSq4WivE20galRd54V/AyCViiaJi6espk150dcsvRKyD6wmN
6T/4Tgha/X3aR7olOrEJFyotzKPQ/Ztjdt2KSARXzE98ji5WoeYHLL/6cZfl+wEvf2I8oDRFfAQl
uZ1hB102dVI9E/+vkdurjiibfjU8qb/5WDeQzZm5RoPXEl+Ns0Yf7Ar7R0DIJU2ReOd7Ac9/nJIP
rPTMkQpojCQhhIgWMmu5G734sMmVrgwMkSbbPAY8pnuMqRvEimiGMT1nssjx95eb7b/Z5kUoHH0Q
2Co+ix4uBG1DJFi80jTNwo6WzQY69RtRRKijhTbGPcVC0OOgEm/JoO6svLdBxEHgv3c5Kjv6pilW
GEgXrUwwHqaqDA5wWFGHllb4chYYB9nfIQHhveAOHqehE6qBP5jn97v1YKuWtavhadV7OC1sRT3k
I1NDBhqql4WuP+QkZaH5AyxRSMnhOfOqKXSUMkQl7Cy3uNrizwKB0+SL0Kj0T8BL7R3YXAD8uguX
pIHxOHCkZSiYS6axSOupH3fqIESpX4tsQeM8nfX5l735c/p3/7bLrg/LwFVm/9BP/HXYR6taPMcb
h/mydfH8AfZLNpfyLsv9R+5MHNlqxIwa29B/1ioUW0SN00Ud7h+m5hWz6BQnVP4PSEP+nCytzZJ/
JN8kfnEFJsemLb8SJbqGo1+kgoH2q4XRsCbGE49N8dyXw8FKWtKzCaP/wD6M0D873FTBApENiBSU
oXhgweqbKvijYQ6tt7qVJVNhk16Kckay+YH2xwPnelzgKYYYDuP9D/nkspG2MKgLQY5bJOvIf4Ko
tQ0fxJr0K9Rs12OyT30mmCoiv1GpdIKw4hklVF7WNVSLeoIUk8jZvgUmz/BddK0mKkzACMQGLGeb
/QniR+0YoFNgg+YWpGHECHNMgmCGPRdPL9y9wk9Dr86+oIPGAhmCZGM/RLbfROlFK6o4lGkJjcYw
zxAKN4hRV+vfoYsn941Aw5ok91bPcGD3Dm22XsFhms3+HvDB5W24uoAl/gFhJaSCuR9oIBfc7M56
sxwGB9ZvrxlqwG1HuQSj9Fnup8ZtG14po9/7hQB5SKgKUrFjRYw1iKKSE8ggVilYFo1wHwf3Jmiz
eG7x8oEiDdGyeXbVPcfg0tcIaej//2VUp/Pz3WdNgCPLzOaGgQE/yU3d6nEb6ueXYYZJltNg6c4m
2FxcA1ung06V/kY0OaOlbQ5aDRXt0xqs/ZadW0gmhCunNYiAksLOwFvHKNCJV/gMjM/2oBDQxh0s
zpw+EdMu7cqUc0aZKh1gJkiVl9qd7jeucEJcvKwdLfOfX6v8mvmMxMKzh7DIy4DW7xpCTccF2vLy
k4hMPoUr3kCwonQjU/Hn5udgTrcA6vZTx25AlHeaDir8ByUq+b36pyfC6KqvzOJHgCkJ6NlIPOkK
X4opf2qoMSdKjaN+oBDDt5w+0GjaWaCqryqOHDyhxm+PthCHyC0d/hiqL3hr/A4+Gpc2tBT4vSr/
jwwPIdgyFPI42pFfkTaY5lli5ZXa2+68mg1HrY9NmK+c57l3LzGpPgzz5dIM1xrNEbugRv/nU0PJ
/qoMKgso3luL6yv+BHXipn7LooZmoG1dKpbHS3+wEgSgP3qA8/+YWdwNMOSwb5VxEMYeC+KVVVLh
0T1iFjgzHDut5uzXav2WALBVvaHdVuQALaGy604EZaFznYyIA0VDCQc8ljL/JA8D1ojKJTkkS/g5
xawnErGL6GQmvT0THSwGFWOQakCIMPspkFwPdas3oRddmV6kGY3c3zBXB4+h9S1+TiqhGsyReL96
sxFpzgp1lX5umczvkWBoSzZxOvJlwEynrh9nDZyjRbdQWSiaxIHmy6TheChqJsrHR0BULO9F0/pi
T5Gn0JZLNni+RKuMJmx5VM5Dm7C2cUnpkSkXa431MWoI9qiNiD10f92STO5QukTXUUXplTkJFVqO
J9npIqxbG24NIo6cm9MDYyfPY3TjzNu5dD+33uwxfDItIM7ZJlK1VS54pk7sv2u9CPAYMaygy4K3
Ys725yiIg1O4UQZQ69P1pUC/MSjG1xyzmmwrf91H67VBFRkLb0IB259NtFonEyG2pbEe1zaoUakR
7vUJMy4YvTccYGpNiDIRNnRpaNhe3hPzqEkrBkdz3dKCmE1QqJ1K6LVVRJY1MXRYxnmG/Nql2iLg
ziVcEGziK3N0n4c9s5m6QQM2/gJT1JZWQHBGoN+GOhyF0/1LcJ0ErS4kP88J7/EXOX2A56Pmd+CD
0r6LdmuS9Qhy4he882hazALpQDOeE4KhWiphmHQAKLH0xirkwBg9gmkrPgmGNYwgFHMNfHQkRXir
EmebVRY3hkhT50bzTFMgL0DvSg+zWlbrA4yOhGizUirRVwnHfn6llN3LoEwESeTaIRWhXvgQ8afB
v6A4wY1Krukv25P1LwwFhyIVChttqzKBAcZRG1g/gCIYJpg+izkeOS7gu/nzUt9ElZCAa8u6swUS
kp1nWLwTkOyAcx29Ph4pw6Ivntd/oYlAaKN7y0MZ7an7rIt0cCqgIlkt6QmRUlqcxbrlCnMi21qa
/ARr5+TSYh0nsCNsb0lYbSt/9sea5azfmyVeBSWLrqNlTr7L9VPLurlY+ItnIAmHYzX5zFIb2jBJ
P5AwmHenn5NiWP7TI0brZ3R6A3cI7a1attPnQYNQmhXDWLEaEQf0DGsjfdmOk4A6hXCxw6nZ2XRx
1/w3BPINFdcvEs8/vn1H4OETyQ/Be11vPauFwlFUutyvxO0P+eOqnQis/sh8VaYBPvsR1YEQ9pWI
aPWkVvpC/PXqeJB9C9iKExwPu+0NPXAOwj95NyIKZbTFB9gSMwx3pdQX7VJMorj3MEBb+cp4NbZc
ZrfVdA0fzqM17Gfh+urB+SWOVsttbOeEsDWOW5DyZJizlNINX5Fxcp3hbPWhDGYZAZVmfAqW8E/R
O92DQJ/l7ux1KgvhJl/MFgOHlzL5TF9cXtPFnAhWW4ngbldywJYbnyd7Idp3StG6T1YkI49IxOHl
RzLfs4X8megIoqJBLXw4c2TVoOJ5jQ34uvyFbrYsxdiY2bmv+gokNoQ40Tx3JJizxOHokP10ONue
TsFmbuFJlD7PxkYSOPgkM4ZhaBRC0wCogU/zanKZxLAWuOiluF6Xy7YiHSnHCMABRRnFUTRv/7ml
C9GK384HhjylNDMqpU+lbNcpKWhzf/ydAMmJ8ymew+J2dfTxF/VIoXL8T04UKgVE5rRrF8yWaBIL
GhfLABLrAZ7CzMLkdBQYp9L0w5VzoKm4sVe7Yn1fGgOa+FvzpXznkiP9hPw7OGlJbQnaQ/MowmuF
knVTmk9kEIsZBKjAkegCyOcpZYR4/WoJWRKsH+yPEaubkqSXFQGLw/gyTBFCY9Et8bI7hnUSNIl3
OkHxsqehSXGqpAWwQirkenHX22SdhWsVfmUDXc7jN9YdZnkyKrRvYrl4INPyFr8XmnG64TFmYxa2
PmwJiYODPX18TfCDh1f6gMIVTMNzzMfa5nMwqbxuKmZysrz798wnOOkvB75VFXmEq/q4lx/qu8wE
STZIVawljBjgpWCKRliFq2UjR5ud9T4GDJ40dQNe7OsO7BhuZhlue2pOQCJJHq+5Ryq8Yzpk1ZrW
EDZf6h+J0l6FcUQMdD3LJO6w3JDFMhi2lQ0Flv0bt/zHcTH/g7RQnOOdIa2orCK014nW0eVrnSAo
PQy9hkBOu+KOg3joV7NfrK28t+F6vuXpYO94XMdxaPq+7BUnSBCa1yOwTvaOU+lB7pM3UYb49Gqa
ClGxIA0ZL+Cf2x37PnnWj6Er5YdMY6ftEAXlRnkmvKJu40Yaj5Zu7XyEKBieJ4GV0rwc3TVqkJgx
C4IYhe4QcwpyIBKUll3odMOKsINm2v+ZhPnxbhUxFWuedGXQlQJ0qUZTeYDclL5UtzFkZUiVRmlj
8IgQipkT2mWL2I7CmB+8sxrB56vAx46ipeLxlH6ILjri7j2uyCsUHnxjAXxNKwPLPJhO8zYMEJ6Y
zD2QT9Qmx6jWo+ferUStVLjDbHgHvhusR3s+lYJpKCGfZKOyik7IhAoZvpxdRNoYkwTPnQ/lAbBE
bCQa3FTrRI3Pw8Db/3LEhpN+xXslSz+MWApcgV2RGhyP83af8U2fLJQcgIvalE9h/uBr2Ua9Etzp
kSJjVE69oWWStcrDtah3l0WyQwNbrgO3Ow8YsKVKG5TspaoCj6Ea0RX2YqowrHxiRTfOER7RVbfz
azQz7+ljqxK6/9wGmIbFkpQkXx6KtMLuloqAW3jzhXiqIJPi4dNLWSBGgZ3SvHIG/SQ44Ee4Rx/b
NeWxoAMaE1/rzWLWngr4VTovdHZQxJRuG9+RCaZW9vjfPCKSC13Poykk5xpZ+F+RciCY+m4yhDkT
keO6TUzeaEoQ40zENfJ5d8fQ8MF9r4FkwEAmS7AK0KXAjLRQR0YIc+XfHDI8da6F5zdoPSZpGSg9
M7RnT64wcOGff0IOaFQJ6SPIT+ANM23Qb3RcAKTaMKfSW74iyQYrzJJsAXlACob3rxLOTWwP4p7w
bRqyon8Mv0nDy8v0cgfYz2GiLcccpBBeT5owoKhPuGuyfOqeOBpr2qbia2peeAXnV7rbDXr+cNBv
HJ++37O4WzKhBQvSpE8vWGmhjETiG6sbD/f1LQ31ziNG1X1GmOZCoqm4XF+ciwzPB3Tw6wrrkdou
gRfoiGOgHoTUIbDDApHH9rq5qBHxQ5BNT4fhrDOQoVUes518KYyHDhWXZo6eV7ZU8BBrwwk+D+LK
JwqBb/ddinHgNwXD/2iGGDulrBFMf5qPlbIEmByTSR46+jyMlD1gWlSATtRkLnCRd81mFkhor9N/
LUtpKmIlC46/nI6bFOPCK2QW6k85m2sqTz7d5G/RomZ/Czf9iyYSeFR8ZSjCo9ml/wbDUYWc6yJ7
CQ7/V6EfUhnu0h90et7+1tfduum7F5pRD3Z3swietrbhA8xSHLi+0CyFQxA6PdspM9SQaYjdBhe0
IBbHMroPjUP/YuYW71jhYzDIy95uLNoQo2xiaj9KsyFw36IJPnv0QGUx82ldbKYmybTP5S8brk0K
OTR3RQI7RWmii2L5g36tgmrmCfPandSnI9gfY+hsEPVmar/gzUDLhnA7pceYxyLw2OQ9MFZrfOV1
EyOQKrWgms1KOa1WU9Z2u3YciJNUMNDcSbJTVMqJXkzxtiQQnYkxzWWMTY8jYCGr6mqt/mKIMqbf
Y4+8gPazblElmrua2Wo64nLycON+hp33U3YzpOfxy+eR067+q9yE2UELsqqH9QtuytqISibmS+j4
TGFoX8Ts8Le1UUfBsz469TpEdnPEeaUGJ+4ahPcNTMisHkP/lnQva1UB7nk0lqOfemZZpnhoSf+s
MaBNg3W7rP7DEmX7eBSNXpNn+16QuRrWAZZhnyEvhRgezaZq6aRiOSp+3tC3HUrqFcdWS5eWRa6X
Cr2IqX74grkK0y3U3LWWhAK6raJGSgFuEhG7Z+2+8Y7yE6R8uNledBc50vhCHs+tQ6ag4LbXOat/
pNl6VMQuvEmDNZOdDYXMZBchKHYVh4gAnX/DYEiyl2Ln80GCowglbsa1V+uYnZ1h6McBN8HHMGqM
3+nr5ZSNVU9AcmIxM1GUnQUjvJW6le90+RsbTmW08jTvl72FgK/gygO7auhfZC+lqApR1VBUU3ua
lK9AT4wY5nphZHBwkaZb9RuSnX1r3nSW7HHSFAeaS66wlAWqQCMLxz3dPoq/C2a86wjU/Sn0Za77
qg3imZ89r7Nke86I+Lx67YCjLYEoboVoyHSJNkKIEe2MSxSW+Yv43LukGTFRazJ+3u/Ka0kYPwlp
YqmmaN6Hm5QhknjZsaKa+zkgmbkg6M6KL0WAQ0BU6IBEFgnREM5q9AQn15VsLQ4JbIGcVn09FeMV
uwDCL3QjRKsqmCihtQjeGUakdNv81Jdd+JwYMJm5ZYKJlatZHXlqOegoKqIlosk4w/7w+0F+xfpz
j65UXErqc1zAkPHxyPWd1TBKQ7I7eJmgyQZL1GoXWFumIrhC4OnhpPlcty+vCFzdq1Zj8kcQ8vZw
Gy3koX17LOwpCBCkgzHXsDx/LFHdAExrHQRwgEtILZPmiTDYExOqwtiXVcbf3lCrFnAgCowL+UXy
CN9TBZ+7rxg7sb17ihEQKx699lqvIExXfpgKRmGcE91Tb+y8brPiSmk2ROWCk5NeIs/YbzkNVgbC
Uofs4jVpuMivAJgwPHjAGrUUX+qPnX8hELbq73hOWHbbOTYmVU+M0yO87dWTYTWcdKHYeegk2ve4
eLB0nwfKa34RKa+1zkHERH+UQedfHeHoFCtlk4kcFWEfRZtS7HHwADWlhIzV541Zv0tXITmnYD5s
xzrBFtc1D+1bo/QJW2UbZH5IPuqon81CeCLZYOj7eEEv7wQbGkebHVQW3F9wvyXv1G88KdkLZrDt
RKdmnDLuts1qcHNsCAF98XJ317VGZWIHFWnpcFxUcEM7SJ5bEmOJKT6apaz/ORW3vQHixj3avyT1
foMmEcXFEpN9TpJlOcoWpHhsqo3v9OR1bh3AyehDKP18dfFcfRyWvCq5C1ZUbL4G/NFKAY0DI86y
yppFlgUiz84RRB9gvgnENYYykGuPSuy/IUIwnRCTPg2huvmVOsqBJPyMcnGzguv7EklLWKrzoRCF
67krF7KVZXGlBTo+9YCsDfNrtILZqgAZpsnkGpAvmKNNVZVfaetmEoWiFpNyMSd3n6lUMFpX++Xl
wxLXFuEPFLdR6gvhGeZvz/jt9Np00AWFakjCUZr9jQoDdB+25THl3BqWRbTQjScK0R5d3yFsb29t
x8AC5WAvDE+NdPTjjwJjiF7htZrNYEaZtvtu43qq/8xCiPsoroB38uuKWtOWOMN7be78pT6IOMm7
/HKsDA/1b/9UpbFQJYl5WaOEnpE+n/1mEIPQ3/1jz1OIv+lQq5RMKXrxFrJPLVaXKDkmFlcy+/zO
NTqgFNQRNLbCafzToGuPm7c7aCJ98xqQ8MzsYMD602mb/l1JfyqZaDIQf5wlAolOY4WzYgKb8ziO
0cSycdrEUNdPrUTg6mCB0YLFZi4xczH+MHOIJlkrkSTCjQPOQBBLhzQDmP0DObTr+V+V23bOBd2i
sQPO8i+H+NONDAnZjVcDMkkeeqTO+BkJ54TAo3we+mpIt5FTx+GYzGrQX+oNzV3m83ZxRPhgpsoG
ZhYLfwpyEvIQB4F+kcqWrKBR+dF0OHmi976HtIVxr5CYndQyXhsVdwg4E85TfEpM1HPJ5obsgLo/
Pf5k8YwljKEwbyzCakQ+0z3UIFefOHaibNiqylgzeLf7UZRHNVlznP0BHrvg1M71Rka8WplV7CZI
YZS0a0R5OIMnKW/sg54JXAlaVlmi1OWMiLW2TmAqzkE/LQM5VCvBJFhuj1RDm/d49u0JjK16UI3a
gmKygW1nnt44o1G4XIEldh3y1HpfDfrbsjnnieaHKHWKVt0pIOjPgkC/NPTO4xyu3M2Fp5UOLl+d
rVL0n6aM/ru4fhTesROFwV6hrEstfilYZxsavoi+zR7FeNUIqDNQLjIkYJbtwhHOyIcTE9AS1Hp2
sgArTn2FxMxui/N9dbv5tOnSzftL6HuOdS0i/1W4nsgg8GCp1M1+Kt0BKuy5HfumVgDlZBYDdQce
PWNBQUv0Sm3DGZN7H5mF5rStMQTcukBIsXyYylgpsaDTgSZOua1UVL+KLT/H3wL+cb1zRJgL0j5r
Y8mxi+Hzz5VNoBJx//oxEc3lh1qxBt1Dyh63ON5P+EjKq0w381A1VIROxZn4aMxFiuSkCRevr1Zx
6qVBDtwzVEJV0QuQY+zEpzbAN1OPkT35cbJDD/dY7h+T93MQ3iB1VpaBTy6vTO8I9wfPAddrMvWS
s1Kmm1xys/zVe1jW7gysuLIvPTVVkA/lPtUXFUaSAoWH1eOmMvgTmAqEYq56RgHrZc34YQK1yjjB
1G6zLI3T/p7E2daAd6oq5znvXlZ4ukqIsSFBVvfQbjtmDBEzLyUI9JYHS+RajiIw4k//EFFHxdP5
BZkLkAY+pqmJg7l0b+pCQfieBE66GIcaXx5Ix92cj8SxHfrn3J9/bYn7sjcy7ePCpnfro9sUfrDm
j7O6pd7ekxfPOpnit5R1AGHZefEXOQrJt8qGw4zFXN4gmDxPhq7id/rPJzNmv3aFHlmYYAW8p+y3
WCQ2HFp4KrvrTUPa4hPdfTNTN+zwvgWm0NJK3S+Ld0ER2CTDMK2785lqSR+yKXxjyKiYsMBFYfuv
yyM4cORPBXuFdscM5vGJo+wFeE2In8I2klP6zWDWUsnXD2EhzzivGVIcj2Mncajylrgj07KRcB3B
LWHRK3nmr1WS4d9gTmeNsPEB89IPACW5JBlFbtU/3h6+JU3wsFTBqIlrGlJvLfXY09Auh7s/yJpf
vWjkUCQqktUUatQ8OqSEskcaZL6XurAqlCKfy8eH+WuQRLdmt0jK33hqHpNOoUBwTfB4vUXfgkMa
26NR/6nYP+ti8JpdW6qxvhyfSl+jdZQMrVEuPmkmvvcxzfJ2o+qc+p6bTs7WG4KQYUMEHtbfSK76
uO35+P1B9By1aYJXSWJ0cESUTdL5YDJlE5jS+oHqR5miJkSTxPgxqkVmGezGbmetONqa70FeadVu
VU8LbhlSAhAHkEefzgngG0NyaxV3HgNztkf/bjGQqoepYjvoElJk8EMc9HXN+v9CJ87/XinIQ0Xc
CksNhZDsA/nZAHmhSadq357DTx1qb3ikbjXLvw37x55w8kEni9xgt5nkjPME/wShsBCg0VjAZ0lU
Cr8G8YafGCzZBEzNvc7oUI5fPNEkCaRCWas2IA7fHX1aaBU4cTmcNqCumSNuIusbKkelt8cQ2QUS
h2xNSA8BNZXONeV/MO+fw06Cef1drgWF3slMmJlIrdGlaWyTxm6c9Vg13xaeov81jAiyFFW63m4N
2raUH6avyCmVbNo1JJeHmZkG+u18E82txvPpzy+adDmjmlFQQcWe/cyk8cRfsBMx6SNgEcQeh9ik
6N7IUe2uZdVBzVql379ftaxsKgihLuCvtzsdKFdzp177pLEhXlSCE/1HTdtUoCIbE1OE7WCFnyuy
b2u3opk6+7VXZkbxUWktg9J8Gw444iLeBPYBNpVLl08EVbZVLkiRp7P5MfLv61GXxiDKhuj6n2Fx
BvKitG74pOswr9RETpxpnP3JxPpUq/xFiPBxfRkYK7oigvVVHGo+CTyK26ahC3GKFFBiHJb+Uaa+
b4J2TMyTCS2T/dtgxoz0IC1NXAzaHj0dLNBKNPH3cIKUXMxoSeoh2quHcbHXa54AaFr3zT8PS8ub
vaqMMGRbjVuyEK2V8twlt9qMNsioPKC4fvmc/n9CLZSvDS0jWAk4273mB/MzFv8WpAZTIHbjgOSl
Azxk/5A2iGXi3QkGJURXfZEhTsibmVwUSlAQUHydmMq/OpeDnjccXztKdFdWBtzecgnATmrlBs3G
whYDsrp8yb6k30+LRBfO5MTzyHQXWEYbsbRcONyPqBQ4GH9t7AmHVD5gqm4/eMO3bEERCrW44NER
QGLnGUK4OjuaCdNWltGeVXJcjDNWjid3V5G1UP+bHcFvfFfni3oWFFLGCBjKQZjQeQ0YzPgP43nU
NdJ120/7VwGbJ9eYPyH2m/tUa7WtZmCShwqABb0Ekn9QWSGZWzquqmiTljrz3lgab/yUrWGrDtW4
022zV6HjOeI82ctgp/gOrjyzCP9mOF21+i/HCv/oxUbEKxEwwfgU6HFuSNRoTuJwnCeTdATNQjPK
VOnvn2liFZoHSJdBI4t4TQXDfwK5MUag/8nffJMfcKLUlSRXls9u0hhy/3Ods9rmFSJH+A4GvCpE
NThVrMoaGywcoXGsJXzkKsWg7U1Erpd80h1L1l0VFEZECKIBNSkkFElWUCoXrWmeZRS87ipE66F6
vD9qlkgB1XzLMt8bkPVvUwiTGVgiYK+ZzEedfB4BAY/jg3YQeK/VW8+D6NmS/3QP4gcKJnYFvy1D
zLbDNDZjqHvtikJPw75wfhc0GDzC3drJiJxcQaUMRMrfsMeUwPHPHLqa6uvTIC3KjLjzAERZ+BK/
K7IRtLpSB+2ZEQQqLaVJY/ZTBeyEq4OR0WYr4ZPRhGAWhKFGQEM+JVqqKw860NwqEdLMlCr4ECtb
TAvqMDFCCX3tUQ/WPRH3hCy/+1YnYXdOWrigC7/OQlFEPODtYDsJmJVM2AHlc+PuPEp7SzLcLVwa
3Qk3HyRWCD0VlU2qcfpDoKmh5p2A8xdB+Pcgrev4k44A+MgnjI6ae9zCzDLn2xF+0JWGLzidrvmK
PYndinrTNuQ8S8HjkQG7G8WwkqskahCO+0h6JaaugRF38Rp24Z5pfBniVGweeNXAsJ04cMIUfG1s
DkpGRQfAixdnMZZhYy/IGg8FNkqq+Z/NEyhBshlU2JoLLIn/bW7YYQv7gTx5QodE7+dKev7lhjJc
8ZwmST4JPyJhI82+ak2tYIE4Gn+oav3SUkloU5xKWj6BEUW+0fEIa/upgTyJcIyM72Dmq4v4/6N1
OMlnHvZ8WsZz9qbDwZ8AWEZO8AKqzaFoz2kBf+KTpos1z52W8MNdXR+PHahHaIHroIieOLoMA1mx
LMNzq2bECmAKxyVDhuvXnI0PJhHB+v1Xza1qLAqaH3f9lo6o/a+rc1I0z0UEfcyBFcp3IizqAq80
eDJQqy/S0szpFnw7wk1JWp8I8F1+e/abT20KU1PB4J9GQF9GL0QpJldav8mC7NpQ+P5cHnKFbgHB
S8qkP95wjKHEbaFl8VWH6TBodPFycz5T+mnLBM25Zm4zk5pTVd0jcpXVqgrz8SQtQeVz73aolXHy
kCxIvheBoRtr9eT4H+ZzTc7isiN67Y9OZeMoMaVa/P62MxuwSAcqqfa/MABZYQRd2r+715Q+d5Sr
koM62zgdROUxVh/cXDUyNufejzOfAny9cMWz714lqlXF7xHossZEv7Bs7yfFsp1iQ6EzPpBuVehj
9I6sp8KufGoL8ItOPvEKruGGLKJuuaI2fbBpsHMn68C1ZlFuqkD0uFp6I/9k3MAIYH+n6jFF9eRk
WFgYMd+snkjrjZryshr1QtrK42SeDyS4TmX3cjXZMeHn6G7Yj//1t2MCI9l17362KqdfT1Nj62sG
zESRCTyKL1pjU18NRAVCuGPekIlwDYuKonte8A+oxC3jEKrNCEXOw70vdmB4d4cxZRYTtag5LrDH
31iNk9VMmZo9CHefI3dQUe5diKVqXDrKXLbGCeQPEisO6fLoQPIIPWTskXhRK9SnoYTg12UeNw7r
Qs3YK0TMClBha67gQjC+m+IQMZuotOstd+DcPzld86YOgdAHTHdvPjcwM+nOzHrTLp/3+ZWplP5V
j6G0Ddi1zrgucARxNsJYpaBTEsEnTuGn/gUrFS1duVW1PQFwJEaTT+Q9/EjQSXNaK+jD3FEg5C2n
r7+mWsk0y+xLbs6C4DOYeEZkN+6DtVeHkqLtg5KW7YjorBJLbIFY3q8G3gwjiQ/Dmz12l4Fv1Asf
JBMI6vUQfM1rbu1GkciD072RXUTH4MYjuhoh6u2NcXLQm0xEigfcNTasNTFQ2vjdRrHymIzPlugm
lSef16bDuIBgjzVfSAW6kRLm5pMWnFq8MuEtMlZ1eK2qi6SAlioWqgxt17S1xNePzH3vbycXT82G
IcVqfkQE8ZnpWPqyfAFH0uaL+SyQC+T0UnXiTqA+XmGygyeBeSNZSEJpoa8hQWGc42whPOIqHaIO
bPEyk/zQXFNE+ZtlusCugWlYzPlewxjMTdKtsVRDZnGwJcCP0j06Gh18PYA6EoDE4xpP3HQ0UcEz
QOI24Kyrt8LLOSnRBHV9RzeugH97KnCkxP8t+KWY9Lc/wv8L4lWCy36nyG606jQqsHzPlMQYmiew
usPFQJNIPR2VsRlQ9Eze+zjx7sJb+aOMg+RlwRwWA5x9QgdQdt34MPrmVmr8agxXQKDvmH3UtQYL
mYzhHtPoZraon48tAEZd+1VfnGWML8IOGG90NrR+zWirdHjO9FpjGSdfWTB2odfmnEFASxMrwd2M
eec36A8xP69VUeqzEovdRtk5oHAqZc7bpz76x1CHiCpnJbh4IyG2/WXtDmV/dbRiyvIsL8l7USzE
td0x1kNVv3Zuz2+ihA/teHbvlFP0JzgOx28VClO20RiVVkd8U7+RZtSXYY6WE6NGX0/nMdR2Hvsk
F9evj6jHpmmt5+4qNXB6bb2L/CO9oB22UZdDmZpij2Ee4EtSyzSBfsOSNDRntqL6wJvjxlWHOBHd
dg+XoXr8hpI94m7pTz9Nk9GCXla/nOeuLNQWekUHQdvyGq9qWu8Iq8r2KmXs+OuzQav543pdbPgG
sK9j9Dp9MVohTRGah2RKPE4PEXNIywR4u5M3LiEN9vmTRF6n8h+Z31+8gZPo/38AKNmm1gCwu6Dm
8OUlCDoU2KQVj2y5KGdXjA0wIK7alaQe7ShFHpC6r1rW60f+T4Uy27JoUX+E73PW1isxf/VyI1tO
5P0aub37pyMkpQg4iy+LDHgIzAZvkB+R7J+wue+8kBKvzQccX37lT07WlpO7MX7FlbpXvpLoYB7f
3IfhIS7PnDDc+9pEkyfsoFii7xjFLRvAFFNQJq5ehBXi1TSQoMvHx89iD7lzVkr0216sWjBjOJKl
PpDXIJWpMLFBvAHzvdOSdPuERDcrIUXzZ/8tfUPTRJ/p7xpy+YayTVJnE6UDalVi6HGZtxPao6nU
DxPCVbA/q8dazH6ygkiXALs5+s4pwVGeKwzhV5pRAsfkckc+MeF/d1GNkztPqdyNvJUWrG2rpRU9
cTz16KJf6XD0nX9LZKi0YVTvQVNekuV2j51KVshzKQ+1khry05vysEYjpZNE0ftoK9GftjaTZqRa
TSJYDopv65OzBohgus0Y6R2LLHX29ggl91AMkNd3Ph7vVqdvZnlcIBSfoJYlMjMIRMPkSypI3RbR
z2pd/TSf/fhiTQod3U2FdyjiTeMCedHIwM5sAYOXtJ19NRvyyIZMUq19bsLfOG3r3Ch+fWewKV9l
6GJ2IVnBWC6oegPVeD8BoPznBwEsP/LU0E5pjVa63EO+oQYduA2TLU2TnXUAdKT+GxFjSg+ussQq
aBLhg1guTZWVl18bIEM33GM8JnqA9wgwZHKiAbqUbZ8JTOozDtSqOE/cDiG5KSbOITGV6a9GgGUJ
XBNhliU4jYWSKdCpFAno5QyzqVsTQ0xoHDZ+0r7xxsYv9sas7PTd9eG7YWWbRbQMkbc5TrIf1kKp
zEbj0085PsuoYSMrFeo2C56JLINok7lgSgmGmarGWUC68tcuLUCP1XBlNHmni4gqy012zXa2xnjq
+WdUXjbuLOSTSZwBFQqP0P/E9qXGbAW+w622h3L9KkKLD0y2SUuBHZNQGJDW6WXsiw4B+a2kAtAQ
LRg5ck891LOM/rwfBLiSC+bpnnY3TO93IzlhZumop1tXTM+GGmtSYmS9+bfcpkT4Yn+OqYm2P5UK
izMmTKmp+k2BqNSpN4SCcqLNDVJgDSiUizF6AqHFMzulcLg5hvbDz6PTLm9X3NiJ8sBny8cF/3Sw
2sS3dLJBg+EE0APKV5N//Py8zotSb7e8nk3P8iQffz6EDou44Gxxm98rc6vSmVJl6jpeRUWFLmEX
7HiwewuthcB4CfIt4puRUY3Km6FAhLqY7cgT0OPSZLmab57iqR1wtzNVJH8kRvo/w778F+CEQTTC
CtXnMd9TdCJJ/9C00KNBZaIs6ePOZFDvUwUMfiCgiTfsoJDOhyhGJzi8dortiFTeF8cxTRJPsm12
TNtXyGzbupk4Bg9LnNeKaqrb5dZZ2bhTknYJybBAuae0Wh3zK/sIwVVR5cDyWj2eN1d1P94/wera
W1Hb8OfiygWKoc7T/DGVL9TBIpvdp9bM+4K+VNbm7gT1Ibge7s6FpfUV7DOw35d17//902ZzlaSr
lBi98G4AAriqWu4Do6+ZXm+KBZs7r4IwHEM5JyvVf1vVlQQBfaz9/kRXya7RVk9bdOlGsJJR10Eq
yk9G/68KLh9u7EwUsGYeHMW035jbWd0PZYJywz8v/nZOC9w9tOzS9fchBTA3J6DSjB3Z0/X53CXf
cwpPSstzNGarJgJOLryAsQ16ucI9awQDkX8OFtnHqHmz/39Cepcc03IT4uNHGNFPSD5l2jWLM7kv
TwriRstoEcR6qkhCp7AmZRz26GBuYPqDBEwfNx9KHZLpBvnq19ZMI8gR8szl0NlS7aqVzDjbtAJx
ZHGl5rnVmnVHTDm8d86GX7VV/7mcdXPxUgKizXg/HnmcocoqhVcz235SJLYBLgvErGZFNe/rX3wV
K5rjkEc3UfMfzh3vsJ5Crf5jZk6xjry9V4lgnrEIZ3egNEBUpZ2jgeiadvaDDjEHHelR0OJhFfCv
5oHBJBm7CiF3s/AMisZnyUspSkUK0ng8v3kshhBp2rS08my1AteTVJcRLxiutimTwVUPFPDDoCmf
TB/y0+LTcFlaHHKGUyvq604URJwfN0wEpTMhm8OfooYSQI8UzABMe5dZcjLB/4myHynTOHF2amCe
WeYzP/7A9+tfEH9ZSBBm9y3l7XXtWjBr86W4O1tgCvFJYQU/X9o2jKSk7C/RxUIsWJiPMfiIlhdC
P2QfJfkQM9qpVgExKJlIE/fOufaONHssTgoRxctExIBJ0ngCvQzqSs7+gXNP25nWziiBEsIXSmVJ
Qfzdj83USdj6/SKy1GF0jrk7bw/OaRhFfR8Dcmq2dnyHIFoNyAfHMeRtCjNQYb/BTtAjHr3l/A+a
guU3g/u5OXCllLSg/cPZ5MdlRaIs9vmo+RkVDImz78+4h5ag017hytQgBqBHAK+OsDPvO27KrbOP
O2nugiY0Vki+JZUD3naTl846LkH7mj5FmLDmVivTFes0HUkhpIr9A5tfWZ+ZVZQ0Cxkd1pqQaz3H
xceyEXqsWcW98FVOK2/CnpfIx0KnoiUkLX0TIYEqbdKBWG8synuQti8vu0LHxcovOeFrFUzZ5kpj
btC2rcQe5MTHF3+ysL14iZz6YFnIZRKwoB/0Ih/I4ngsvWCVxakrdpiS97l5K71G1IlsMkEx92Hu
XNG57s9UBswawdCYTYBAWwmOAsUIebc0OObxizgVpTT2VG4eFHAwdCXNgms7XYxlXspDOIDpCRYA
JnBk/kdpZEED1mlDV0Z4RKOHvKOHJ6XOXEW3LLYxRbkv5+pwhRl+cDyD6zOn/iHMWXdMgz3z+WS2
nEHt0CgorPVtWVZOsAQXQ7lUaTIOL2V8uvp8+UfD0GHHKqYNZuNDu/w5XiD1qIggO2heHGJMC+oJ
Nkyqng3fK3UmgL1GXviz92SRzgvxRcVg+ZoW+xPc075YqHiJRw33MJ0KZeqib4fOVg3uhJrldv18
D67TZT+op/KFpLuTwD46th75K27MRGVaklShTI/KWQhL/p+WrXTPa12BLhdFnbCEhjO34bSVOkNI
mvoXKYtkvG0MAZf+w4CDtniFTIMGGuGZHyLwGf3TlEnkfQgFk6wnABtcR7XKmtlDM82sDXCLDOxq
SjMo2lnizcMeqIpVybMmTU3KvJ8gGr3IaZzQQehbCHJyBA7U/bDJ/r3S7qyqN8vZ7VRoss2/M4Bk
n2ExQMLTq4NhlvZoGm9+NTV4HF+GiAxNP4QxbubgnQoQvM1QZXsc2+zqPF6XOBBJlbLAnfCqrDMM
d3ObryFlJMHf3a7xuYmCSAAP/XOP1pl+Gb1J1nLCp828c5TSJtbaiwmBwstuaTxUJwyT0h557Pxy
XptzWtYudO/tIkyy9pHOlufg4E1w0o0d68RwZKqxNGVPJj8MjyoIzAvxG3jfJzY16B4gHNIFSJbm
3lWlxuobNqsazxilTAuBdslG+YlJ4q+yI9CRYVNADY1SmVROSgXnYllyp4YC4vwFBKdQ1TOizSXG
htkjmD/fxWyxD1XMj5mGTrREXtfxPkDyCVXT1gAS/ncAcfn+XU2ERKQMXlGCC03osVqnLWsDvKvr
VGzOnhcCufiUQryYGR03Dh9xYhQpxZRs8Pt6ebuclTXp6WPGZfx6O3wPfYlvvXIGKJ/1V3MTwo2j
bE8DAADmpWe52+mBxY3W/JmUTuhKzY+5OWJRHHSN4o2C+q/NG5jryrwNrfgpBzNTWHSsdmTN8h3y
5RI3i9XQZHwsate5A6ydm4S4Xqfc7kmV8dRyw4ZtnjdW6NiGRcCYxHRyiTgO+JYT+WFjBYkO/gi2
6njtv+SOvnVyTfvHUpZa8E3eI8C8gD8J5pEcdvGnoXyzNGcp/1DevVOyJOkT/YZuPbTJ6fB8Vcin
tZaEnTvkg2VspLHi9cQz4qJC//v5YArmYTpDfsN8ZmIupbzq+1Vk/EaG8Noqc+qiYaG1LcqUChBT
PxKfScIGAABJJ/CRwgwoSDK9q04z4zWHZnQjkQUCMhLM3o7laN4lpBYExZVDl07jEtGjPh7dFKpu
+wjdW5nhauA8dORGtwh4RqXXDo6vzHV/avVEXKDbEPMnyNaTHX9wxEOHeWEEh/Q+dNSZUaMLLk/1
T/wgBY0lF11e3ORhgjN1EyHOuFu9dswPlL+PGtkjpjUQds/EaO0GkxukZZ45/+QgqRidLC3U644H
h8gUJBCKPbpD+wC8SYaib0Z1iGcBJroMEvooiMN+oqwXx309oRV6YxfnWH09GQzn7AWlVvj4iF2D
kDHsZKsmIQheMpzZ7VOqIu4rujm1vaYP5fH8YVau4py04hbDYIE0XH8N5safi6PK+iNIJsSxZx4y
4lGkSiTGby5KGOaeD0itr2+Xg42wg/+/QLRYLfRHrd2faSMA1o4T3fm2t5/Lcp2ZNqEZIjCCidPc
zI1V81VExNmdXHaqI0glNDw8lYkJsu8xX1XhcPaHLJssnz3nSLIqBbOZEt/LDGnZ3vNeHcUZ9V9b
Y99ymkK3NPPyLmENcqop6M0AJwyd5A6b3+oo6xrqrKbpq69gA6JFvtlN4f/omSVNqoWoH1AmWrcp
i1SmFK+mnvmCqJy5xgGXemULgbnQLa+OT49JgcVdth5XLHVx/2jEokVr0kH76ugbg5DA/RF3WYUT
YNtTbZ93wXlpdHWd2QGSAGou4AITM8mw/ss4/o2gfQRlAh91w3sP2wHdN/0xhc1Pi9Ug/f4S0pxF
HcIssgC1BrLhHt5ftLJC/9U7Op6jyYJWNcPBOoeZ5zjjTNPiM3DrEWaP2lFFwAoPJqwFJZ3zv94A
c5kYr94NHJt9QvoS2SYbQnzK/pVrHx7xH/6QAo8iCN9/owS82dVMQZPOXYigj/6iBHlrjsPRm2VO
k7u9DmbMTJpgGGPmjQJlP05rwDGzFG7hejsYbGzktDfXOAKH3MwtlFJTZwpUWiTneDpwg9KilgbO
WBskbTbKKwZmaY96SxcoAQOiM5sHeDJaDSUexKX8uCI0WHTAPu6WTiWzvVfaFDQykk8YjsxL2+CA
gQUnIxhQyQ5iD8HvxF/nrhXtUmVnKnyrVfqKjHfUXu2gbPJcL3AzesqAp6ut3OY4ACAEX/6kZdzk
32LCtxegsGplVyiyl7uAoeX+A7plUheVRRKZklv/hzIv1lKLy2CshKEgy1fcnhOCCgpWBZPk5D1Q
51+2JyfKqIT25QMR6BjkMNcnBpJFHL2CcaATWILS0QEClcpq+PbIY+e59dlkx/jm7z63knrZkmdP
RHzgaWZWEW/nmkT3iWPGczyzggxl9MVxKPW+yMdlUelMbWaeawZkM82rcJwJyEIii59vLD0bFHcb
JnfbaigfqTCRu5ymZiLH8HscwBT75YzzSTjk1bo+Frx1hVyCPzlzqhv0/H61ToklGtlZNepnbz5X
RU7f+VoIxLmlRbMkJgtOh0zAMn4PR9MeutlgNBFSa4XZX97KaPCxHadXINqutTccjy+yJZh3MdYC
009yRSpB6eJZMrf+/35y/P+96cmY9xr9QiYKpok9EEu5wssth82eWmp0HxsXdHh3CtiCT41ad7lC
EVgYh9qLrFLSuLGs3ydpgYBYZnvtCaXOuHTgksNzGPjzMLVN2lFhqz3QeUNDM6g/rqQjcUTyyHUW
x9jrLRQYw+na2DvWa/nQMbgWSfBg34pyCNZ3YqghCKidY4roRU7tcelkOjpjKyl0RkZNThqLrUzy
2EKicOktTLx5gCO69vDKMQIQnge8aCnXyoYtqLr5jP7r6bGWq/OlfN1f1gUufXuC82ESfpQr0t9C
97M+tsvjN8KplHqhTURvZBSZVZ+L0NpW5GXH0gRZvzDXMnFYXMIl4wGnZrL71TsF3pYneTZbRSLp
4S+Gbw3Ab5SLPPMtUu7dsuVJ019OzONmcDP14WwOY0qwDFzuzSKsv4iJ4o9jBpSuYY3P+dBAAUqW
SkC0CMSS3dndmFe6Yb6Qt79u8SL7fOumcTB7GH9DM86r2rBKsaPnhvdzgEPiqB/N5jX67tN3cgd0
OhkWHXO3OVhjQ0A3V6qD94O6RLvyRTln4Dv7BFl/ZKA2I/3wNH2yYg6oasHs25eN+aXZzWOPrIFs
zE+MVltZPHvP4GHvagYb5enjKTlFMKEiqoM6+N2mabO4VEDTjAbeEAWCZp8PxaqqD0Z0ohYa8CQg
Kdjwv1wykc2toHaZrncgZOnZgvkRMdrp/SdJfGLnl5Qrz4/x+Nqu8er4czRNhwIrlSsK+8JhbPf4
/Szwtb1nW2bjynrfXvF79p6okJJTIG6KUAgvhbOl6PLXKXRSVZd6CDUPwsqYd8yrDMcLZeOn0l5r
jkRWHreWLn6wNI+2FyS2SC1Q+lu407SUWfgr37nsbuXcKtViITQ9Ki5ttiWs7uBZjDod8c7xsJyj
bDhdRwNk4WQkYiEv+5pDcNOVTXfyMdQHp5AKtFEMyN6oKdm1uiaQjAaa8jezOcBLY0FOFvFq7fHA
siCGBbmbvovlshtdQKrCnfZ6v3xH8CFKw5ggLHKGbkq1cWMoKeJfIlZjjuZfq+bImtCiEM8xu1g0
x7XTAaiXw7biOq5flZ+2/VqxYMm8ht8dw3HTUFYwoOGOMrfHpN1+D4BmzTkFdrD2g57SeaJJQIJK
2B8yUrwiNfyY3WOzWJSarG7K1vXoXxfR2nwhvmb7g28dLxwMYwF1itdFErbXXv0vgN90FrqUldPf
auBvHrCNNfl1oJQFnkm6zcM7Bn9vg8Skm6bUME6OHwokaQnXtxEw5GazmCFVb3kaJ+D3n3mS8Okt
B0HaKOsQobqQqRB2mYmJ6csjQB6meX/krfAwNM6QdbMuUDD3+xy0JwpaqF3A+BNYrZQHfk2DtZX3
xO9nsAOtjUWugPvY2AMJ+sBegaCROSgCxwA69ZQUgaTyJ/aN9eEk5nyKHCKK2pZ0ZWTb9EUMvb6+
wkm3qt7wgbs9ukJq6ERxxpRXeUfhMw6eOi8N8wRBU+ESqs8DtnQ5tHIeMqGee/WSt5y0GK5BATo7
PNBWsPbHBPvHIJj/cllLlT3jqmiN3LXRpUC8c4rfspz2QLvvXbxbecv9ViRoTfV+hf0+EN7K3aV6
6MVXl6/zsrAStIMxGp3ZhJo58KXmQYwRLw7xKCymk4OuP0wpp3gST42sIEHXzuS8wz2bCs7tjb7e
rgTJ77PBo0U3f9A80SUl9TUx+VksnkJUjqbzcQDZFI1O6E+bmJR/lniJBwNoIZIWjM98Mf4gppc/
x4ZetQEZMf4yVlOb1bO+23PwtV1DFj7RIOySicSDrVk3hie9vVvC+TGa5iOTFhVsAw7CgGa0IeON
l6WMfFgxyQiHQtJsmIHyuXF2qACQ0TO+k8GbkSJ/Cp8iw7nRL3YZEtvA1CnLR8NzeUoiEUxTZ9aN
YPO8zYVfO2fEERup6Fo5fDTWgu6TEc1UckBU97lfybGerrP3/vHD9kIhuRyyTqRgIn2oBsUxb0hQ
TvQGZpM+bxxzB7c2lh+fkzR1g5rU3+NE4pOGCQClG4HNEhRQh/B99h9fKzAO9hz9c3XeHJ78StYl
J5GapAMqOW9wS9qnmLTVhqg/nRHv+mbkTB7y6BHjItsp5AWmJun0caSxG1M0iLhpzGb2P6cERXcv
2Oib2XwV1zVh8SCCER//Y+oGKqhbu2MH82mJ5sxZfQ+/JyGfvafVdc31P3pZ9eLgJrprPOUoiER8
GyinSoldo3/tG2+OOP0J985Bgh2Iwo+oJZYB8RYLyZXCTkZXRdG2Z08fCAA2/DCV5ffP5nWZrtlf
eb+z2XuqHOLyyCV/ezmyfEWrArtfi6345XA22oK1VlNCBCDWgR5BEslcIkJtVtg/GGwmNStR9S86
3T82PdVcKPbVTW14mVoPnXfau2g/5F3YjKw+UsJFwDmQGp6M0eZU6QOuJmlGcWs1U2DK6JZkEuVr
JgqUkh3tP4xg5Ii4KNzPbfgTY+q7e1qmGleo5h7BExlxdJiiYAJY7yTvL3shZ9Ojic44BxMTDVsi
Z57V5oGq+BfMrV5aakLwrftV/BNTuKZvF1tVFk/g+5bcO+lmSENb2V14fhG+qTjpwZfVe2LYXtHh
dSd0zRGdRUVSG0aDYZEQ89dK1sHOhHLmBPkJuJNx5eumoJLCbiumLEzeStGdIK94eFGMgR9zT0kD
a264urCDuCdCWcdz1jblSEE5P3T1YW/DGaUqNzNALeIxLgjy01zysUOCWJzDCLq+LkHZ06esJZDg
gk9mL2jgwkRX9rtcwcXB2Gsivi8cYItQc9LLDe00krQ2snjEQUB64CSBZe8bWGyY0MYGWU4ibqPg
TNIsHM7I8fdPdElxotSrNSkyQYr1tkH6aQnrzHbZqfMNWjvAUQ2/MZC7D13CDdKKu933jb47yJtC
5E3ND6vqubRgzR23nxm0faXbd36duhzc3Bb/NgXe3aTC6n+2U8dF+NKmzadtvIy+m1Gmd0HsJbIN
KN93L3bQWC18k2EK0bAUhurleg0YKom4kZ4jNKuQ+DY7lY73fDTCfZujWHFviOVzi4uBcYsUdq/S
mZAWgoMwCUm+UoxMQAB7UX0cnJqwD6IMIR/OpIvLvji1Y5pnn0pHsTsa1nO9WNJiNKoV0D8+dNzu
yoowOtuDlRgdSV0WEymXrqwNrQ1pRFyFBDHGX2hgql5ZcEb3K2U/3ECqBe9VRqAJqUf2hErjWOJg
vPLQsgvWRHOtTAWykdqZebyh8M9niICF4uJrAElaClpZxqviNaM8jvHDiTA25q4ECCZ0hRC7Ocgd
bfwby0f8GnkFR+1upOHYQqSHTM55o0XDEp/tm5+jcDt4b+smh86gHyRmwnS7rovQgUAQZepFD5Pf
dqbbWcVPiwW5ajw5tyiuYLuUoVjYr2arLU1SmdzRjep/z6Aeist943kMPyauge+198l7SUEMzemm
Im3gPieEJQkBVIbQ/Z9v/9oK4kvx9V7nl/WzadcBJ/d3rHKgENHxB40EYM5Jt5hOKr8697vKtjKZ
hU17KiTRu+3URw3TH3tBKbgqekPmuFKE0GOjXkwBQhvg+gRFBb4DShh1wE/av1Z73ppTPzSiuPNP
31+ZyPeEvuDmCCt27ulvB9Syxm6XKrkal1B1yNUKNPSieUpJeq5QvVePu+zD04mJnDBVVjJj9CPS
sSiWPKiJ8zU7fXJShWn3fOolpJe9ZTK3OyAfLWWcv5Z7hF8irp3IpRscobhB9kgnYj95tiaSJs/g
0McNZ6Tc9tV7MMKyt2mQpzMcpUpkepA4MIo1AYrFDdSeIv3a8hNXQiJYmLdqVcOSFBlVEVFlgeyo
0lQbKQzVMO+cmEsOCNIHmNUDc4vsFF8q13H+up2DM+LnELrT3v2VgXS6ClEBkdwo3M4QO97dYs9Z
0nKRWn8bgMTGpNB5Rz2l8xWEMusjW+PT1JtPCy9lZn1B0gYLB9vX4nst/tZPnFgf6tcg1w2qxF2U
thXjQPCogz5tXSw6YGNa4DnfYgVuJuY7Ly457VwFSkwI4TaqwlNGBcOOaH88dSm0pEPaiPUgCN2t
FV0YqQqRlwVxfGSeJ0MSMhAaDELtp0mk6bdjPM8MfkKIG8U4g9UdsEvThbAZym1j/zkOTLorTVKb
k+cWitVbO1flx3ObmHII99KxXI8VN3zFKPw7quCPVcPovk6MBIT47BA7xYCvRkxOHHEW+qcdN2Sw
tAicya0Y1uZn+LC6BeSAm5CofK/vEDXEx0ofj43DylazlvuokHc1hLbDsmATMM7CNuzaXOCsaed1
NRtyA4owgLwAuE96E/OP+uX9FtsfLES4qmoeQ6/VoatWc4DlYTdmnHYWRhW93PgOrSa0NSVWcC6V
bvr7dDoPTYNz1l1PgaZpyJLrKPhpPe+xlq2HgdsC3OpyUUZTHBAgw2tsmRVyg4/aFQomxsG0wbBY
qtpVcJDoXjV9sxQosjKp1QlbQTKSgPgeK4Hzsv5xNjeCGULKxnWuWP3sSRq8FIy5zAAggsWKvPKc
rnGuuBz/7gD9Ew2RI0j7NWTGJpXz/hDT1s73ns6oM91yNr3Hki4GsIqmhy+UH+9/fAa7XSHAWHZS
nSWguFG+nq1nlIyERH4a/d2bdpDlG1vBjfxaV0M6wNoCReaT9TGSgGmjHm11Bjl2obvVSfB6uU+/
d9TgWEl/RqoGxrc5oj8HsOiBOBGyzc8xzyw3/tmu3vPpOxAc5FZ/sETEnX9Osu4RAS+9gNw4C//r
cFRAqHoneCvWxBuFSkAIEBaNiW6L8OkDj4vwedbP2RvbeXGkQlwmIUKPUdGG4iMJYnkrVzV0mU2Y
Pf4pDwvyyj5Pf0ryVbdRq9VFf0AA6qHvOHl/mrM2hPU2jzgdJISkkLgWspr2wcsejFmOgi5EE0Gj
TVf1UBqONsFtVJJV76yl7u5cGZC7FSeQOATgyvdhesfw9P/QRIXtZBNoKEEOsyJBt3IqZuBxlYux
yBcuMuypMJYYX9w9Gr1o9qDlhyyfQaW+fNXRSO45eu2tzzqYCLAM38CZR+txiyERou8q0IJwN6UN
emNJjdKuWW619SYoujuYqrO7pvRlSsTCZYT+d3mQpaA3MOvlBSPI8j2G3uBWfUjg5nGyqYfJcIa3
80jbrTSuykgG5VxIq4LHfm3KhMhtGN3T4XDWoVu/QLQaytjUdysWUfcTLrqebqmLPRMjornVTqmi
USH3G5giNW+6nWddQlS6LKQb/+S0XZ+v/FytYYdILzxpBLczwIVp5Vwvzmvf/iRVP+KLaDYJ2whA
13Tzz9n8Tc0RvWKUxZgx1W6fr76rguh7oIALu2LpTPEAdDjKsOT1tiD0jArIY3j4nqgzdhX/8J6e
ohxnCBh0MWV6CBdVeO3u5ga3FI/I76JZqYkyJZqD6uESY/rzpLKWUW0vpFmYAj6vha+sJBDGfHLi
C09WMsyEtgbOX+g9D1dm8hqN3yK5E6b52EfErau5JoJTrPD846CtuZLqRpHsiZWOczW1asdBLerD
c37QtWJWIQfOz2Xeuy3FeRHTVrFck1FOxJd+eLzpvgIOswvnfnYCigQQJsdt/JZNMLyABqXRi977
jgG30OkB9tiTUANnTOKX3MHo5vkcBolLIqaO2J1Qtzm4IXwDFPk5dPbp9tXKh9XTPJ1ecnQkH8gR
kjJLBZEvDZMia+cTAPe+U/+3/tGRibbodWL4FXL4MAIpLdFM9BVQbq1l+rXEOj92RkQAlIbOL3NI
5aUJ7rUb2TE83lpN/nNWdKTLNNZS+32jJZ3ymp0Y5NuvobgLYG2HPdKkm1XsewqkCG6VsbMKpm0D
KJZxTjOeENv1x6l3liWp6lpzuCj1NyYDtIDcCqLuKeGSAmSFgCvaF6Ba+kYA/tYoALi/JPeWTeVv
jRlAvBkg5qLBAZOz7Z+712CEW1L7DGvBIUKxX5PBlkQsOlgHb2R+WnFDYlMb3BUsn8vnZH0WfB5o
EsifPkyUNnP2pQEuEmCpIj5Z5SUfftcr90krro5lnmZHQQpuEm3d6iNxOgGmSUyw2yKSSwbJiqCW
+FYtXGLGTLI+hU3+ynY/unVaLVAbEVrcptsWrvihHCNECN40tk9k3T533VsnyVSKD+91VLU9NbxN
AFapd0v8/3+I3tdOmyde9st9YrPLNj8nMGg8u2xLP2n/ODhlTVCVrD6zI/q+c5LBzqzksZ6DRvcP
7tsWL1f2dXuB5WaAXeUhOYmDT5ObwFyDcf+k0Wndf2aB+jBewSdiBFR3GT4WIg0hGoLOEgfVRiLL
UsqmoSncS85kxQZN1r6Z91g0Hp0lLcj3yx58ElsKaHQhzVJoca3eXPSxGT9ZmUXtA3QjRCoF9eEL
yrjsIAXr9GB39rjCPjctsFk8yGzjt+YSlutnTj0r3gC0VHJZzlIWSpRhqHi884+0KxMb3xtdGHd5
uPNGtsaajSWK4iMhGkbCnj7GphtISKks8ZjYS4nMUB+D0ckrYnAqjUwZQmdjYAulZsUYMOiqXwgw
UfWqcipd7MxM9X8hOtAOSpjF8EWubWUxrxgw/KGizDbLmWhOlZ03Ayd8jmDn3Xr57kS2Qr986fhE
IStz26jzAxMCe+TnJGeZ/MWwwXMKZ93zLRpllTeq4aJGt84FEBSrPyxpUYitIGxy29/hMHJiXXdl
yX5hqL/ZztyTTNGYDg1A3Aq77K7HjDPif2S80pNwq/GN1exJy9LQ7lyNK9o4rH9MnRP3LwM2UKcK
/y/D61xxYSKyxIoOmgiSMhw0PyqCGaJ2M0dPuBIb5GdPmdW77ANxolMrVUDL4u734lUylZgyKK1T
Rc5mhlAgDquVDAYrc/BN3L71JqDh6CR+HOF+dWOesEf+syfijLwb8ldE0WKOLW6j9FGNPfID6aiY
IyHC2l+iUQkT7Grb9MmtbJkTUkmCnK4tT9Sux52BjF39RT/7UORcrXDhWo5ot/g/nh01mNKbtWT0
dwvqEtv2+CSRnkxeBHgombx2j4L6x0EMU5Pgn3nQDt2rYqRtEZ0+tj6TcxSBQB3K5BLR/8VUww9q
wIRpgmeupPyVAZBcBbsrukE+krffHIjKuWnsAY68rRk3I9aJmCfOtGBhQAOwTjFPx9lqRB0Aa6/Z
FbnD7oS40Eo9PrH9AcegSMBAfUQ0cb4Ipid0sCWCfaA63cVT3L//xwbgng9wkEUEChXTFF5hxZwA
HBsUelVT4FZIzd1lWlwbOZ3hm0x7019DHI+mh8CfcErYgT786ZTohiP3awGtZfz3g9fT40/MeFX7
0JfdBZLaiVekwroRgmshTayzIWMKKKMJxzEK2vR4S8hXi+qaOMOkKl5/bEvFj97Gkahc7yY7O+HG
Ltv7/eUhzOTVh2M50AJTBMuyaYB+1POwlM57Ntaq5FIw486x8D7YL95G+8fFb31KbEU9UMpr10ue
zJDUDS/j/W79odDbhkTKRWsvq+Ioa16nEpsOhHFvN/DxYxlIE/J0d2oyQd3mDPnpw27QOeIIUWDq
W9AQszhScb8MzEy37OU6JBuYjUNYKgq2XRePeAFA4wsfpNjAKFiZBIMqfUWEik8n5Ggv03XCWNVi
TfW2cfFzBRRWuvarrF/I7bSJXRDVY0JNmPrhglZdK3dEr0ZbdwhE5wjujKu9a7ZMq0o9ByLEZVN1
MuD5OqmubWpKZEqzU0U0u4hoeddsnJrfnqPlCaEBjbdj329z3A9nc7LxBPxDpWUMVXuhCf45nGja
xDmiMuVeLaz5IxnYM9REAFyJ4hFtB3zv+XWaC1OY7gZ5+skpZCWv+ee2LuO+u6w4Da4WQIyPonA6
WGzk3c8VE+yV9y1V7chbpE8X3ifeC20dVrxaOmjIDBAJvhefMt4VOKu0qbmcTSeAuqXxVo8fNblL
n3U9nnGBKG6BMeUUr4tnK7/+vabMxv/Uvr3VeCJnX8hcesJLmVLuq/9XKaLBZZd0RP9GtwSFRCM2
lnIBxY7ahfEPT4hT0Ps3z+8WQv0DYVpI3YvCP8U0ZENOfByOU7ZS91NLxHT8VDBGAW2nktKlU1AH
YP2JQ8u13c5qpHlkXboKupf3BIoxM9Zx6PigXC7O4xS349RSVR2OP7D9d5ktI11dL1cmtPLPvC3L
WbH2hhBKPEcnd7qLXirNh26pGLLr+WNZrdMCPu2BR2PZY2HI5ULpXjZS6V9uP+qYQrEkecnMCvao
LVAoLm2l01itXpFrruzWALq0r/pQzT0W836Fg5YZ+U3X/MLVt6A1S04p7tXc3FVd8aI/U03a8WGq
bdsw14742CGA1LLl/XkjeCrk9MBgFqeZH1MsC98TPI/C0YIjJ0+qhroRbjX5hec0d6y97wZhK1M6
p67rGCD3D15c9KZMxREjwj7Ihn6aASy2crDxpcrrRKwE9MEgfHWz9P+N8mkaAREW0BGVpteMcvt+
YrYnKsWZgtbPu3AoeZqB4tIgKYc00GGXoWS0F9EjEMhWshm1Rxchj2J79jWcIecyqpYwrcdvxiSt
zwMqso2XiFH6MjymiGElWEFsV1HwgXVEEYGF427O1f/T1LD/3hjMlBGuIdqCfSiG+0f2TJOJs+ye
tlr/kPTlpAu6OoXeB1TU8uZ7YgN2JIal7M9LqRylHzobyISpycdnusq8/r0KqqUP+IV5y+0/f+UV
+wJ2cOEpbqEPjOBKsA1iI9m1lbW8ozb4Eq7XquC02d3n0at866mzuAzaf8iX34gDB/f7Bo5CFnEY
3TstYYhfk4SyO/OFNXipmImIG/1jY0tGlcSeDDGT1LVDoLh8i33kL+iEH8/P6VHu346M6nPUOjUx
SMDWeKpB83lA09508hHP7Ah+1F1cyj8MP2+MhKhCaxZh1LWlvbJD1dkFmSO5rqwMUezgqKYm+ka6
1kd94KlmVRTW5JO9ofz8dQ4xwXhqNUZ1WP2MJySbtPIdKxLIkIgo/20Ar7f3O33hVQtjW7LY8Yvd
NVtOigMFBVjDjN06fsSYN2y8s24OHXJeGM05NxH0DEXa8oP5P3s5zcCth1yN7X+Q1dodGqtdhKx4
SyE6OtcKZfq/5ZAuKdIlU+nEGlHwQ8XbqDtFDH2jRgR4cDnUYCwm92kfh6QclxqZysKXrb9U/3D5
Sy/yIWxQndQHGmWjiMV73b8xjLIEQwDbeKA553XWT730M/VV1Bn17YShp4hH/HKqQM60KDmk7IwJ
DVzJVDJSXMhozR5Mfmsc3mL/LnW2PJxDJ5x/IWYJl5uR/OtDjLy7OPwG7V5dzrJ5pAgbabnzU5DP
rWLbqOE8m0gIi2gnDNAxveix9Y4YFjFSMfniYgMnAA2GT58qUjA5xzVsXlD9MxslrS5lEpBqDf8P
XvmTRb1pW/l9Iye6EmEC50RFikQT+jJGkGl+fOdjp7LbOvePS6o/X7VOhIZMeYQQqwxjuGTEii3G
BYTo8Uv3a7F/aLsgsPom6M0bIGJ7dr5yoLV4mbaa6EnEK9wFai+jf990nvGgHPUt5MaZ0Gh8nUf1
63t6ql2L8pGA0p1PV+u6XSTmYhxDxyC6ZOxhWBQyIItvqQMa/zwcD60cooXYL2Fa+IhBe14k2WaI
kQefJUTDo4JXkSJAULCbAavbDqzyg5aKxYE8oPgqBjIs7drTXr0sqc0GjSKJivdbV0wIl/JtNsML
2javvBJi88qivM5C/9Ty0NEusqrNz/hv34YYD5T3UM6wuzAzAzXETGRJdkZU6cReCcBk/2+lf1hu
iPrZH3IRRWoK5NYKJC1KnVrFY7R0rpV7Sl1S16ZT2yLOMebkOluz0MCaUp4QHLdvnpxKGW+BBFPy
0eGYmbWibNP5KO3Qao0W0Odka5+t33x2JhgSAq5m0H3s3BSH76KXiOVdXZyTymayXgb34wht4aQO
Uah678kt+l0h3aGJEjf1SEfCsvL3avZMcAow0qY6garqUDH5+3Ca0BupDMC9V6vGhJM8bE5/7yrm
FRzifzBn8JDs3he8vuBZUnVZq+cBQFa5doPCJ/5zh03RpIRls3IdmY3n5hMPx92VJcTwmIj3JGAt
0FFmV9HFVEyNd+USHf1spwfVkSakw/zSSsbEO3hqxZe8zVTxVcBmDyQOZdp5pM1NNIakzHcQJHu3
41uWYN+XFT8JtB+yg7VXTmJyo6wPw8j0StcvEayXmpcI+YM2xEptfVJ9vBvJWQJF8eCzrgNcOPSu
e+qGQ4m5IeETHaQmQe58liIAHOf9Dp1L8WDyM3M6solUKN4hfvHsj9QEsfzqec4KvJmPFIW8175J
wSr7eAImHF2W4w+Jff+W8vo5K5dgny/bDonMkNSRzIVkaBWh1QUXI655Whz5w6/Um8IN1i2UoQZr
G/cJMw+bXZEK/GCwbqm1La5g6kQHgK7+A4OfMgK3iSu9U02oHFlDgyhGdYXSa0L71NpQSwHD+qwC
pEKHyC6KqsMChX5w6yIj31Wde9m65UnjbrKDioNLqxpwolYFYHFA+sWMjtEWmwNO8s03MinQzzsl
twH9Qv8prIDI/Uac9aZEUyOI4L3pnNSut+nV6AqtvhQ/kmSqTAjjIeIEWNfFHTjX3tuXdftfPqVS
TIxXluwhd+4YBTu1GDX0ecvwMPWyfATH7Zz3xQY3ob/YU3bjpOXCmrgLnMzeYftMoE2zJ1/6ltCs
oFnDW/xFj+Wlll3egYqGi8d5foIvLUmA3DBdjHn/4IqXBGkA+ffJ26iICXg3WkXfsYF+EemBXsSd
TzLKKPBwILW94D2aa9KCqsmZHmrtxzjR4M5fxAzc2tvf0spVITfRrcVjvqbnwc5aA7LA7rTcTGu3
XWKyzyzSkIB9za+zYWmomCulHEQC79qwUoVbNeK+Wgwz0Y55vmWAdfW5ybioeLUmI8vlreUNDaS1
A9sgzlC3wAqlF0j1BFg947uwsyiPNmTZclJ0e4k/WiOTn4+iX9hXnYR9iZg9K1UODiiZCRwE+QwB
+lqSjI2kTlNtnVO7M5BsMnRkT9IeJaSqdJE36EIbk9dBsd1KCMJq8UttVI3VGWT0lrT0UBOGXps/
M71thMMaHKgattIhC+Hlmh/ihiE2Raie1NQCoUZuU/+DTPQof4Pis9Ndzwn75tx404Ig8HiopJZQ
V4dSPAdGZGqYPo6X6YS7jXhTeAg6WX5rnMFIrIRYK62s8ffbtN8t/dHY7OnSxio2vu2xY0Zw6gNz
09eHKQgd1zCXW7LOb4eVtCFWRfMaNjy0HWHjlhMjo9i4/cHfmHGgUIkHly5HMNNb3Q+o4aQh5+Li
9fW5hand5tSbrTpcpsBQ0HNwdF6S7XWLMZ8/DJu/JO8pObS+dhN1jV0fqDtUN+NFtnUWB0EypeDd
Wj0e+kYDjC8PRyy2HDZxsfGwE4m6uQmZFFdPA3jmpkEKqIVzddMsVA/2sqrBUghKnkvQhzM94Mrn
InBBjza7CpVPCeW5FFlRaeZBal+y4lj6ctBWcF0rgLFckJH7sud0UuyOCA0onUlXqs88eIQUqHnK
vI7ZYQRj2bUQffNBgXlu88OBWqFMI2q3CMfnxaN2m+4SlaLqhCBdnhPPEE5IqK6mVmRNxhThOWxe
VBShS1ifRcXbv9/VUB7+ui5IQSkyQOyUm2UvhJJYWSVF0WdfGAnuzJSgAgjZrsDfe+3EBoO9hmMq
iqW7/G4EIDgPUyqRjq+meoIvJS6DPsZ8VPkMaU+zGSAw4s812e60DhLUMKlOjgijcsK0EJGkFX3x
k6Z8W1TZyUTY2CW6e0elsrn5fqjfv4SjNROiymNllzZPj9MKe17qapMEqzbwU3ke8y+rdXmPyOiz
OKzf8czInY5Qu2YfWuIoWwVektY7NFnWbhFPHYlYB9crsF2KKTyB2T2f0SVJ8f9FF/kXEMVbASDh
ROgzZ2wLIYmaOibXY3vUTJiUz/w5CH/Bqb/GxMpjxMcyPjRfJlqVUsWxbM4AFWI9nsTjEd46P+Wk
adroRkX8M7swFkNCYWpMN2KhDYhqXFz4B48lK6o1kgXu8mZC6WcHzog7kW90flGQLToDcNp5PiKg
UGS9u9Dp7mLhbvVhMzwxk508hMGD+YCP/Dtb1dzcmiUI75WI0eF0Jm8Is+CQNcLrd2MMAlWHPgJi
CXjoLRPkq9b4vc2WL28jg19sNj6GeabIYSqZGUIZ7Euqwu64gS43J/MrF5ty9bTpyqJhQqG7TFaz
gVHW+EBpDBnuKPuagrLF8jweZwd8GcBAK8EoOyr6Zcv5yqFwRI6o3qaGdEXAgNUtXPbCKFPWhUqo
9ZSxyHGARJfjgFvUh77sJON3iSTdk5K++it4Eq8gqHyLMcNA2N/NF0OjtRrS++PRKsmCsbslI8+M
PRBhGQvyqY/oPgjZ33QX8W8BgqSYaV9PzSXt9whA6RvUZlOzoF7t9OEiN3JL5TlsntMzL7yaARMq
fYWblKjSg/mTShoIkxkiiLFE2aVHkG+0OCAHNz62fGAR1S3eEn5lTYbrrcdIr43MTRa8i9XJRifU
cSrs1Eeyk8Kj96Sisx6Qtp7MCJaFJVkBnA6j4OY0sAvd97XsvpOSHwT1Wi4d9x4iENQOKm8g7fXu
Ba25zbtcLQojbsD04s9cdD/zcrwPPWmr6QCZes9em9UD6I2ZrMSEx79d9gLymcz+M95YF0PUYn0j
COc1G8HcQykk1Zo4MrbKtzRdnvs7FPSsGdh22nNmxpDIE6lJ0YO8k/nF67k6aEp5IyOPNgPeD2W8
7J0Luhkypl/RSu+ADtKybXLkNOSzLu6DUY4BOQ7vdIbcITGSozlp0XwXY0WBL+vYyAAaRpr6SdHr
jQzGTM3cZqH1+y1tKCIhZJ+6So2cjK+GLCiCrIIp/txvu2u3DXcJEVAxQzuhiaGG2IF2jYGMk/Lv
9G+9u0Hpq4yurCxAzl/hu/94I0C8XK1J1OcxSOy9TqEm1YV0U3SRrLRFDyZ4xjH0UEmrQZ67OQQO
jBUet/syF6CP60nyH947JonLyWqH646TBbSyfnSThOR6TEAdJfQRHRmXniB0B1DfgDajRyzTdsOK
caV+2HWSSEYY55RTauVEmg+McAe2jW+oD5LaFb5dMRC6ZDfT9DhIOy5izsVf47L50RXtfOY/uP+3
l9umWEZoF8JXNlzmQElUa1Cedeu1lBsPATLbZo1cH4UCezSyMA3FsOgpkO5JpN8ECyDxE5efT6jc
oMKx85Kh/OboFubOQEpL8SQl5dgNxAd/KHTD/4iYzHzVv5WgH7KMP2zNango8LqtpPGksAx/qeGn
CymfZIh/obSIOefRNDJLIl4YeCE8lO4O1cWQC1U9bQjA00PlLAFev2ZvuU6/6VOrJVIY77aq9CYi
uk9yS95ZNE323plH625MKCsCFJhToTJhokBJS3lUizx4uduS0Lmo8EOwPss2sJV3GDcUVSdwaUvm
CZ20mnCp27LtDDi2hkEI2zisWVpwGDHq7aTQXZTzmX6tcTg+7+CzZEME7Np/T2Nx9m2mFPgsEGqU
nltIplHMv4qKvapnJloyrLwCYmoWfswAHuhXvq6LFBjbHN9qFiN/fMoq4dWtaj9vD4QxH7KBht+j
rNUKRgPeIu+5B1u5J7Npyi1aIZsUrJLq8TEPvV79/JwdZdTmo+0GDRK/x4eLuufEvzlT9W4Ol1dm
t2wXMXTsEt7TB/utVaE7Xe1NSv964oND9VNBsGRnhCLE+7Ij1thKPg0Hkeoec3Ed2jAUzts3OVYj
XxIZTF+ZE+92dJgLMRL7nahjFnqGTXw2Amiqa+4FXn7Xpj1UsX1SrNkxL9jsCTI9hcBRkoXmb6Xl
mVgv8N6pAl76TL0UhuwAUFyCAQsfvO274VsG2UnNYaaDR5w+0JiTJTAZT4Piwo+O1GTlibjbvPuX
EiFBb6oPnVqYE94zkP/0G87hX/i6WKyQ6qAYb/cPybuezTs3zDWghpMtYHxrMSlDO1WlM7fzvj02
KejCFuCJT5OEll/EJEeZ+POk6v8KWu/CxFEEREaPDCKsvLj73ipRbeQ+Bi9tchr0UVqUFtcBTdxa
Z3B0IGM6cPp0tVIwu52/lUDtpQ702GyLObFzOuOk3ll14elzXb4ciN85zgwjpZLAsVO9yf4D29hc
olB8LaHkfkj8dEf97InvNh9Niwi3Ix0YhDToP75d6DGao72ygjOaRC0BQ7G8ivBW8bhcGKoZcsYf
ZALedoVMSgzmryIosg4EHJsiEGl5e5HZFtZbU6Bu3mSo7VAr0Z4ZaJ4QkoAungBc6nGchM+Zz9Qq
+uoHFoLBldlnhd2pEkrpuko3+ZSU3hYqfZ2EhJdjT7u4TzB3haMjISd5YmDsEwjJHHr4L4AwJGFY
p2mk5O8BxQmMYcC2DtQz/d8mPIqTG2D6wIBu4cJSkJaATf6ob+QJpvYyMJEc6bT01f1FKk07me0A
359lMsOCAb1xJYGyevH88/fim+MnEmTsZ/eMdarCw2cMvDj/iJuFW6sC3MqsWo/7yNvwNE41trlr
gGy+/7cGqxofnH3AaXq5JIgoGyHwj3Cr0KYOA1BMoXGfTcSI9F7uwFLDi5jwASL6b7+rzDMOa3fV
2EcKaR/ku0HGeSEJb2P0eeBrYXmbxGtb96C26uNDfk0kvfy7rtQMxLTxzl6n5H6pQR1ioQlBDFcA
LaCVNcXsobi4+yQGJh1oTOljBF1QnaeD4VsE86/4CxnJIxgDkhimszlJextM+7hsYBolIDiyhUhX
VM6qhShSf9Ajj9wGt/pheINYel6aHn8vg2TYHXT5ohZOK+mqJweiCHK4d+mFJtCxfVML2WpaxBVA
fKXWMAqge5oyTPzkDTGk9ByxWutm7zyX0O1irNzbWl340qvTdaVcCZ3toFB7B8k2odsHKKkEPAaj
IWqTThje4vWa4FiCeGXa26byx1o1h7592qK9Mvq2Xv42oqPgxDM9N8uODWzQcICy7gk1dGy51uP2
rUTlPrOQjmjVM2Gx2zw+o49sRvDcMkYdaoXG8wy21QNkX5iVOXHBrzWdEgjVX1+PnHXeB8T/IzjJ
qk+sKyfgKCfVtmKd1VAHwA4VviXZ/z9P98MlM5KmsG1KJdb2Pd5j0u+bFjjYGxrASclRd83Q1z6a
Q9sj07rfjJmGeq8zENBZKTOf9i4+kiILf/zDtMAnAOXIQ4BJFm2oRB94TFt0jKsDquFXDX7jmuqN
Vas8C+Vidt+oS0WaEltfkia+jdE5u2mwYE3dihfH2+BBnkVSvaGI57dpBS6Ri7H/s0FyTZ5xo8hX
ABgBHF115v9tVeiaKA5RnklGy8HxXWpY8m0+YzsuedW68QcaKzEXIlGgIiSlypS7VPHfXZNgtH4B
pUmkVrGwUaZWedwSUNmUimPvO1oFxOwVgDivYEZOT4CBgQ7V2RdD4uQPPY7A0BtQ0IreRUIO51Qm
WA0eCdxZjY5xxskk5LGFDnfQJRW7Z83P+ydjppns5/ulOMiCDuCBDTwV1NiTMLwsNpOYUj3ZfQKb
N3DjhDACeSBw/KB866f/c9u5tT59wIbViNmecqwmIRb+cUxfCcMVMqRlIOJJdKd+XsemMOo/UKvt
yz12skkVpWl1DuXzPPpn+fhkooAA8JbuYyPpzGGx5DMa1CbmJUTs4avfaFCFgNWDbh85v/78i2jd
2gIEI+w9CVYoRu8+qJ262bmSrtufWovmpH23WcROLrZXadrHZ+E7Gl2IdkKZ3G1jC8F5Onrup/jg
X/8N/DtxMkJlUvp4z1UKdDLIyLqcYxP/PEgRWLD/sXKqr3NChxZDDPNE3d3XW8U7qvVcWhqp3n5J
YS+erSAK+QjHYdpCSHDKspm/qsLBnMFzmCrxgbJuUYyHNBfFWM9NxN56ehmSUxxZISp8YOS1dPm7
MCy3IOegjup8QCK/ZamLHUIQAZHeRwt54n3+doFngx5xHP9Kvb4LOacJIH7YkWKIty0Nf9eQtfIU
5WkzSyCShTC3AB933ra4nAwX7q+9jwugCauQfJsob697a+wbIu0L+7Dhll1hv9LYMT8B41d7tDsj
YAjI6x1McWg8u0AJpN1fyS50RJ8Q9yOjOXkb2oWxH3fk16pTjWKXfD7/QtRDd4UMpPBvY9+q5v+3
1o8YusmRjyl1bASR2yvkv+TCsflgNxMrALcDbbJj5sFfgmF+nRvBbTaXw1eagAqF3dFpvtCY2xXg
BzXmtLrw/qt1KKXh58MzA08t9n0RMcO2yokGvxcpD6bKMl+9NZ9yW0SyI4nTZv3F47AhzEeEjxvj
Rpyf1Upc6nJ29l+1cjN5GZw8Bv36btsqz0EzXmpfrL8hM+cWQb42hASFdFp6TiY6OnfHcGUy5BS5
Ep0lkGZKbIj2q5nWINT8rRc87bBq5Ev00Jp0DMheEs00l/hvNfcJDCjms97a4+vtKoc9umdHKSZp
eZVSPgHUUDAxhxXIbY9NoEN2cFu1xDDnFShUJ9KTJwStUzxU3gxQ8Hj5TqTZllzTA5ROQpsjrR7K
KUYA/8teaO3Zv4NDVZanGq14IhshAZggtt6ElwQfOpLSvftAE897ntUyV+vLaJCfcgWHFlBaAkNQ
Sawl8zWZhgzizMNMuJMWtXS/8nQ3SiOHb2o7Nwyj8Bl/gMIqZ+pJ/oZZOV+mTE1AHPFQJwK89tTE
jmGo20m0w2XAXRFRmL4p9Pr85/xIwAQ0PXvTTJBy5QWLIMgXJLEFE0DRDg9BIWDnxvWRqVErCdxj
ZkVEqfpVsgvoC0zSIs7HJ064KbqQdMs1XtVEGtwkekoDR7gK8jQLjD0/mUTu5fkMc2hMlgejimx8
FWKOKA8jdTev4Z7zL6HfEJsE2S1YvBlX01VKLB14eNsaX3ODlByDTtQkO9B9umsMEYOyNiCc1/GE
tH5Bq3vzEeFO95zXeamLMvREjrdG02ss+uPJZ3UFEFJTcMBB/QvXIzyGds7O+Hxd0AZ3zZXrYjWk
abxFd4AXzTwS456kC48p0s9pNSz4doS3QNrQ/+LB/2X8PPE63VryhnKS/sESTA1IUApWT6xGbFik
ATDyyyLJw6i5cUsnE9yzHd711SB+Il6EtMroSMVddL68Q4oAV61IwRt74QVTvq5aa5pDPQ11lCxK
MQOI+aQ2Uu42BG4PhgcNvswgJroI5iJsHuUYH2ElgyxqlInoeA4+lMUNct8slM/58B3DQYTdpCHu
GqywiS03f4UpWxZKeb1IH+qGasI8ossVHxvKW87IR7EEwTUZF0B8UI9HvOAF97TDbmOoNKkEpaM0
qR0jI1gnj0Di/zM1g7JD/iWLjCuQiCZKax4JW0bQJO79+wqxOHQIfZrLp3O575LWYnECP6L6mdNu
qRVDATKbuaytojNXXAdy4LaACc68IuUcsLgMgtqOrxX8w+NO2EM+K4vdi2v/uX0uWKgXmG+/2o7U
F8Qe67WCoSWhtv6/Mo2/Ai5ZGdKVhqBOhfaUERFQUCkzVsdU+zQSAx6rC7hNyUB8p9m39gqxXd37
7DGSVyiM9CiEwIWt7biLojj8/OUeBsxdb3FYPf0HrSX7WVPjq+NR+WCzxoA02GUH17ZpnBGPbfi9
GDgwgtFnT56Mz2Kt1Y9QxKzzhin/GKhECyRcNKDAbh6TPbPjomAPCJKtlqxuj69RTGmJpX+r42NP
NPZz5Te2gxhR3aUKLOjV1A4jOuKwg/Nf7NjDot6zSC0YTH8Wb0eGkTTC3Wcq1zTBrbF+KpgdR9OC
7jkjYSmstz8DcJlBkOK8AJkCfo5aoClkzvoqBz8ClbZEqVSpc3WVDVWGBRJgwYkDItI6pkAa4TFA
VO3cfEp30QaxMY2hUTlhVzP6v1Bo3BqZuCIP9s8i8vwwubnqak6grx8BC2RWxaOQj1ZcLq9Q6oJJ
ktXe4mQmu2499wtT7UzB+xHZnwGUwEI/A1Afbgn6wGm+RnfBxCDaJA8IOapshwADY/Ycy4wT+L6U
pT3eolaff/aPT+tp+MeKvg2DqHf7lLyXT0q+nDRIPofbJPN5ia4MVn1xGTvZuSxXASTEVu2j7PgV
aB3DjFSz7VOTQjwjytu1Hyc+9smIDLSXnsJRnBoCQvtDe61HrP7GgMsbI2SJWiRvOWG2CRfvHhRR
2Ui7uNLzdEnRLMYl8O1T27CigVCBQl03vMIxvJ/skpI2ivzMomA59syyapPdsRXUdCxx7TNHwzIA
uCeIjNa0msjUyNozX7K59AEFHZ+17676Q2HxLsSNCLsDdW9zFTlSTQO8eLJ5ZaJY70OWNHOGF2At
Y4G/fhDSFD8qhrjmdRj5GLz3yZ3Aa2YVbgL8wmvWsG46bt+vkiXW+ZqjEN6ZgNl+wnLN9/dfj44L
2IvZVJtvOcrlOE6gykqY+1JqFwuJUUBQvqA6zIeB5YG/nD66QymJP5kEr9muTvtJgxxRnXQzeYKj
Xy7gyCyTrk7K0ZDrOvhYarqJh7FKA0Tm6ZssfDw4glLaMBnGhopVQW2Af6A4tjtciysJh0s1uJPZ
tdy5SUqC40xwNb9UzFsAc4yOxAFiauej455T+eZk8aGYwYMlPY4X39SaF3lIWztRvrjbkwX3FopZ
ge9WuKtRtnvPAmKORlHqHat4+6dBdl8KFZWMuIhEbkZ0AwWnx8r/E/HkXsQybStSbs5Fo+zjT3N8
dX2GgN8Kx6VExxql6tPkHk1FPyS7iNaZ9D+XrhRqy3/sfr7id+K+pwqIUj/+C8VV8Dg7RYWRSl90
VXiozA/jZM+nzvY1Rtvc+Ud/xeLxMEBISLOG9vlwDZCnuPzgoWagSXZR0/rJnJpUMetK5Hm8xvUU
4uqwkzWiQquumlfbIeNIBB7a+weDTsgDIoDUncgblXBbXkY5M2ssk1VE+QrjY4+l/m45sj6OTVVv
NQWq6xLET/ndylbAy2ZPis4Nilg1D+DpFreT0/qsRQjN+PDLPtGTwOglATRIDcexQ5LMXFnsEVwI
OPNamFwgYhTauyK3aYobSmBnGzmAaTGDf8TtQGiPcfqAGmn3ldkneKkBZm5pkec1fXpm5odzahHn
fGHoahZDKnjbNf+lZ+dfjB1yxjrLB95fgmnMNh4AkMmd/Jb8d0ylxGTfI1EbrkLQIjHASVKc4neg
+QwjqfU+JviIIOxPwq8/7NXJtGjXqY9iY4NziHOheCjyOiL2mpslNPYNmNLE6m9hVWue+AGRrMHd
eKUSxT8MtxPSobcjAAB837LZx2UudvnwvSACEIIvbe2/G1eKEnQOFjU67T+Nzj10Nhg+cYkLPnMh
kZmECos2r6YoOFzEZG9SMM3Z4pIZqr6G+zhkFi9ARQRJpnS5p+s74qk6LGNdL4ViauoRzHPigKzf
50zIupqlHg+7/Fvuzi+DtCdaXt5gFKVnZ9csxMA3ep9/3VBtjrBd52d8YJwAMmVy9F+NzXT4lawr
diOB93zqGwOLML2vA8zr0gYQGsJxla5jVcmggy0EaudeGx0LzItt8pElH9c1vtezKllPq2QyZrW6
/SLiZhBnGCSrGVRffq4p7JeJroEup/KQ3AdG1AzW4T9WQtNxolmtub7aMutkjr/BC8Uwta8PDRNv
46WtCViLMIS+VXjm2FuCiK+T1KD+VjcSsqRfdPJJMK4d/vcJgTHGbXi0ptDU7usdBhwyW0eePaYs
+QYZrvY1R4K/BenWYB+Zq7eX6uekHYfdMHn2DrAhxlV7owpx7lUE6M+ZKDqGdEKec+iRMheEmBPy
TpfrtgwnTHvDnLmAThVBgFcOGWh8ikZSSK6JT+2hFQo2svo+gSlcUDvDbsbNO+W3KqMmGwlX14or
u7I9BL1QDZj/vjn3yVfmMAK3J14LuMtRKA17hdTtQy3KfG09vc3NqggcwnmrMKbxiolZEtMfvUoN
5LzwWQ8f4mzwtN39WkygWLRm5MN/7HMwVsUDETpcqPOzaQ+JBZxUOsXMBZn7vIKazUNihwoGWVnV
+xAMfWsYsrNRdtO1yy09/ZR1k+NlCpviNQtpAImOn9fUavylhGfyf3LMzwcf+nPITnOSYcIs3jMM
p74plTrIMnT41Izzf8YLcfj9kCBmCtpGvNKRUVEQ6ff7stKahCfKxW3y99coFGbcwKBFHvc11uOu
T4KW/zRY5/F3pyUl8cEb2vTigNB/db98BebLbzN6oEeOIDp3sZSxvz6vLsGrHAKr+LIuysf5dfhL
XuH/ddxK0JMV/vCYSE2+HnIPgCp/aQv8rv2jbb7BinUAwsLSS4f3tn24kctxefYGxxn2o9LYn8F0
f4IifA6h9AsrCOtju1u/n6xbuZiOLknPnM4yD1jbTsvCUZwLmHmcwgbrjbHKB+TLKV5oK7xGP6Kv
dX84DeYQarru9MhhcN04sot05rIieTFY98QVsh38+41+ExKSoL+Ucnz2u1JvQUtlw8mRI/CMPiu6
d5gzUtrC/RLtYiwY/UCPhBK0Xc1BJxOh8OSuUbp4nQn0/tx9k3JixwktYLok17XZLP0TqKhU/qu0
sGaTLTftRkn5eOxFEAQQtEAKI+FW/s9S8KUzU45ClGdt+yiWMwqh3vsdEyzsrIQb2pfz/ODwuZtB
AWaNZhR8I0ZLojn4M2sqz9bXRCQF8q2l7ovGmvtkmBqJRWrsfGkSM1bgGFA134FO/mBvSz2mhq51
R8++d0B1Rif9n03GViEr8MKC8/xD0ku+t6OGq7rePTKsW06GzGwO23EZCbaY2CbpLBJwKP6bzDbe
cPrkOi4i79XCPsFd4ajKv0GI2U/iiZU5b2q4pdg4vXvv/nN+TjCD2KFwYrJLin0VQWKYXpk5chJj
pqiHxGV6XWSNSMeOUpNLZ72TFFRoMgrQH2DLDr4V8iCSKd9jvxus+dXfdCFGN51jLd0E3Qz4TulL
4QVlAbPFwk96sqqYqs+ZksgxqJaWrh3n260IcQUnQTuyoKhObHdHRpdXuobGnHB/8MkVV74jd2t0
kgIQEVdlLevT3sYZmeIvx569k6WdGoBCayfsqG9ik3WylFX6M/q1pYZqvM/ts57l3+L4840DQpAk
++krFWtXMd8bQ0TE3vsDbmF59hAWoRUht/cFBG8DXRPCcNDK/QFs4Mh4Kn67ZbyneaXWRmr8Qbay
sZdIDe0rWfgR6+UJkMHlbd4HEGtDwBOya8Xq4ccD4BxTRIjh26iZJbbmSLe3ordm8Q9f7Xb1pMVy
n97h41WmhUg6XCFFSAh88Jo2K1WJ9Z/t10tITXL1l7KOdE2YjAMudZDh8qrTxvDGHcgUmG6SqNOQ
l1cYXxp8AVUSB+cATCR14e7BilVFAAk1XAUT2XXxhPKJwkcCOtZ4O2m52o7VgMNu/Ai6qWWQVQsB
M6nl9/E9tD3wNtyq2PyQfYvgai7nJpy3dwhrXsAxIJ8Di1RWIaEp1sTjDbh2fnLL1fzy7cWztSsf
D4NQcwv2svM7HDrhBJ0mv31TxiKQDHssTQ928Q+rP7YZCY147ddKYEo3kf9iC226Nuh2GqN3IZP7
eyzYzXXGEmyKDpuLLxdIFXdhrhCA47XhHH2XTB9ZF+CwFgpOZEiiCWL+4HNUlb92N/4yklOmZvIZ
P+nNt6kj9dnRRoVb025zVOEq7+MJoQikWT9puNEU7TUWlo3fd7X5DUiM+k4vcQeJhQEptzjSykmi
GUopALwDLNkIqK4SpMIOqGMTKy6Qz00Ax1pU3cFORUxvHXwB2nBBl/wRRXTM/EP8/8mpadg7Hrdx
dRIEl9JzRT3FuzHKvug4d8VuPWTd1FN5gJIHRa5p6tFGw7iw2TNzRiA45y15CvT74AOQEBYPPa9N
XdkPkhuZGYKzG3vCY0iuUA0VbGqw1ERkQBLNOEYXAK0/wH8HhHdeZ+wvYIkjTrEg2FiJ7zWp2IFa
+EAGkvlS4OKKAQn4ui050A1ngHpY0sHwGQJBc1WO9CRZgmiUq5aV7VcuPGVYyHKAmdZjcGJUNe+c
49tPyZGXnQQCZHeGDrfsze3DHVxczIfheC/2aDiY66VoEHZMwTH76GIE5d+B+uB76hMur3155dpW
dkT/R8N22bqLvJH1uHqg41KSe4b8EKeCDcsDsW+bXecktsDlpfWhfXSowtUuY/tio0pbZhObGeXN
qdpo7zBVlan2BDKOor8DgI5oglDYGS1qS0HrUsWnY2h7VNGdFu9xtr1Z9SEKL7SKIPkaC3jJVoj2
B+LvFsrtSKDkPu5tv4uGpxuMQCu1SBjxM9eZ1mRLJywzn4o1KlYk4zBAfZ1lLCLZM5yV3aUpXTBA
BuWqwLwmW4ODQHdKEvI0jyFryPhpEQPxIxNX/P4TzdZle0HL2zgtRc6fy7DZPxdWh5seY9FAxajf
65a7gQV6SBJMIDmNAeFYMDL2zoZ61bPNzuAN2F1g5F0lsM3w0IeoeiRR38Z+mpTvxlzQqYcLBg3o
dylAhce/jzlLU8RvGA+2xJ67Ihkk3DYzLeIwcerE0Pk4fiWWsszU2b86fXLoEVRdpn+rZAXn3ZC/
mnryyLQXulqXi/1xwW8n85MtHux4kKLs7PC87W1MZOhDm8A9V2JXasAuGqOyDopAdzRRlLAVVfjN
VmSe41g4n45kD1wGeYO+7c5Gt8nA06YtLQ0bFt6vaP4THtJeg1sYZx7nujLfT8hpy4rSNblvkHIX
wK3hRhQ24t1NPzwVAGkN7Vi1JRLUv44YOzfMeI4QzKQMYJnLKasE/iYTHj/1QlI6X9ZqXWMn/UEZ
OrAv/RxG7KqoM2Nnsxyp9s0SXwC9i7eoH1GsGItZR9DwFYD0QdoZs/2S+Ith5oE9r2Iat5l06ybW
PzB0fEd0GYLSoxRMPoTes4l8eFGazY95cYhfw08JeieHSg9rQRie5Xtq4jq5o8T0KfBaaXrPiS9Z
RMHy1JCPpPuLU/VVG7bRzeUZID+yFwx2kVLJ3bvC5pC8pAwhJp78LhT5W3664pgRz1nuAel4Giy6
varibFoThep+hY37B/IKCa8Mr5TMoXEQIhJoGmU4fQibPw0J6ZNsB13pJzMZKI6h+rXSmja6iM+J
dwMGTM0syRLDWYU3C+pU/dNol2qIHEuXiXo57AaJZ1jSxtmQqIAB90tqCVtbT+yu7VSbOXoHIxJ/
S128u3V9jPgeOKMgsM/hGHfl0G1Pr5vY5OiP3L7zQeSeqme+smufMK4PmFjLDe8Cn9baANM06IUt
TxfGoqx5y8SRl4JyQSGo/JcUz88+ahhVI6qwB0y4FRHa5rSC01iFAn0T7ome8DjI2HSc6Np1COJh
NejIRGqWQ2WUWw248TGfKgNxEAmjW8Z9fEGahTuvK9CDRkT36/LHJaqIgw8vFjCVLq06OqMlTZxl
uQ96HEKoQZ1xyk7fiaUfnm3ozAxfA/5Ku3FxjFIGv7gYyoe3Xhkk676jXs/vnEjqvQX2JbsQNV24
txZScHadVVH9dueOqHP8F19ogV+Ly/gD7rw/+/UDZCsDrXA6wLv+HhaVZWeJPzy0pMHO+eTxBSbj
V0FqFEqYc+fb0w5APUz4V4IVpW3yVzGU3Grf0JmAxV9U1FT3WQ0C78N4wsCNMD1fX2zQ0Q75XGZ2
OIETnnoQRb/CfgJ9RPgJuf5zDRYYjyfIaQw0gTj6sktdX9X3KzPbYmSJRfXIjAK/wMt4fHW8blRl
mIYHlqa/pkCXNz/mYBBpbHwd/C1anpfIvwvqKhpjV7mHynJavnBskPuieTMBMrGQvtPSzbGt4grY
RjWDj8AzOXY5r/nHWnY9KltbaO5qevvX/Wq/kYJqMRnt0pK9vQQGiA2M0OhstonKEBSee0MGeRtN
h2QWkOgqDyWuo0mtJqa8ZtjgoifDpmANyZrAbpO4L5oBLmEb/q77udKhSJXQz4GonUuY0UsOAI0C
3VWS92xZ/WLGH2qa6VA2uiQjA68ArzYr75ekTSF6vJ4O3Y5U+UFORyvKPO/3WMaIwsiGCDXUV3I3
wuCcsq5aeNHkNfinQuSnOG81NaQWHkfPG+Y6jeBb4dQ4dK8Et2AYJIWbJp4p82XkH47q7mdC8dYK
XhO8zV2Oh7DOQf+GTUTudwfHHLcH2r6R+Ltdpdgo4whM8b1+A4l56lBgzeP/F/ozHz0rakul6/r4
Q0aQMoeHhR674G4P+ZUBF6zUeHeb2y4ALFYnK/8b0cjEde8UhlPzk/As4hb7fUI51M50HBvDm7ct
HAIc5l7EEgo0krSSiR8zPNMBFgDlbSAvzj84ZMoQmEx7kbgBgX9+o40r3JhBQbFEGtNm89WXAUr4
rQG9dpdL6TYB/ZUUphnC2DSQD5lIUiPcLETSNecY2iGkkqracYWCF0g+Rcf7Ppnxcx/OuPaAtEJS
IcywkfmIg4bAbwZdiIZ2qkbZ9+RfeDrTihldWC1NpgR6EXP663aahvbv2GDwTI1HdlCQTk1iCWzj
14GHOBgd9K7iW7E0r0pddYC54UsxCIlGQucnHRWDeCNMvzjOB0r1t2OZsi0UvR22m2JMdNAc6XHa
dh5u7P9vv84HmVl+L245KK582EreBvmHxaKJ80jzAyEx1potFkjklRDX18hEk8Axz59efRgZ7VN2
T2e3nrrBpUK7CO0n5Vi1f1+4fozgXKLUxJxrUBccIevvJzvZgSVFwBPwnHfx30irc4JKn6BVXMrt
vIVOjvzcD3d6xKBpFVrmuAQ2EsUwejnsGXd8n0SlB99MasqzQZnyDbk62K87+tFCj1hsnbYHqvZX
bgA0rmkrw+In2piQN08Gwoehc5ov0OeZwLWlLlcqh0V9MDrl+WjyxomRjFx/acROhHYZeGXiprjL
AIBfjG+wFPzN39S0TioHzUMhxSXJOx7jBpDpa9tLo44+RtVlTsQTi6NDXIJwylQUhK6mD93rjCEJ
nLW3ATnOf9mfNXLWSL2FG2KpwaWWLbRtxgFk0SUVcmimxuJpZw6CWSe8pmoL3zjkdzuTlmPdLRml
cWTC5ORiduILLh5skyQ7Ej2gaJq9nVgcxBwBxtLR45IV2RrFTprZRWo9N7wjOHVMX0I++jYQjUuL
HwUnwm+Fvty5OqH7ferdrsaeY2/XJjnCxmZ6zEUUb+c0sVqjPvxVahxIt4UTKFS8wXNdwAUyG6iO
JA7bcixIhKACH2B8vTzZ1DM/5tdIN09ZTCuFK2D4EAwOpROLrfXF9jxuPwxpY4HpN306NaE2JH2a
vrGaljEdW2gZVy+gAIIAxi40/L516RdtXV5reqWDiAX8fKdn2lvp2HtltEAbhaGgEoB4Px1MNZF/
UdcxTe2nPfyxDYVQWdrP1r3wn0cbkPNZwnX/f2kbPK9sbuN7UXkWo5qiyGawBezhsTaQRaa1TlBT
Ws4FDffddKsTbQRK9r9JbB0v1VJV6lBAnVWBEb9Dx7XOuM6TkD2g/nvSFo0Qy1sNTkDcshbonE6d
asqiZIiYTRBrDcfUKWEt1MU9VqKcEtYE37dIXSuC1Fn8E03gwgm9mPc0ggn79KIkWKV6Dc5E/RU+
cqSEQKMp2u6/mpN4RvZfzmn4bn1g9A/VoNt8Cf3rAxUQ/Ay9fCAAhT+8rhy7vufAJVKJ6kEzhbhU
++AI/mNMaIznGtO+oaaQgMvEYtWaj1jVN2bwNDFzzLSVFjQnttCEtrASBcrr67tOTon2ty7Gwl55
76ZJubkvzHBlYRlPUOGbAQJUs+prbLoFJe+QR6ppJZhwgpChj9qMvWb5dtk4KNGdgbcXTcopRFN/
kAZUZkUqyo6tL6d8QsIikZboCG02ermsYF8DDL1aqdCkqNEC+MfHUwjKQboPxH9/E2Qogqzu3toB
X5fYiuB/RjdDdUBOEni0WzGZiR7vFo1bWeVFUntFdTtgyo4kYSiO+HWOnhnEDvIgMcaAn8RhuSZj
A0Nt+aO7fdNucS5seLt75OmMHOa5Q1f+FhYrAaDnblo05y5lz/v0KOZ2xlRSralLYlaS1Dablds4
egnqE3f0cXEnUJIWWEM7AVgMsHIMWrfB4qUrzDHOI29TQMa4pQCNPJFt51hhsBPOmPjgn6HNkFiz
LsBLK9+juPhxx3O5EwhOqrkgqzWmRJR94kE//ejHFgeW5CxqN4pBsTPziSBm1y/++q3uyc9j2xz3
hMYwJ9+X7PhOjwXFP2GPh7WFibX5UxZAil8cm5bEIyjS7VF2ywHq7Kb9+nmD3WwW3ihlb6Trvg5Z
hTI2ehxbVRnbgyMgfsRW+TUIDppPWQPJ1Pp3HzGsD05QHb7myc8JfSbt8UIuoc88+olkOKm5u9cI
0jtomub/O1VXUPBW49Z86okye4Wnq4PLS5PZMvM7qOhz3LcN8zLtnOYbwIcraPokaieDVR34n+Z2
nSA0vGkWCcQh8WMhhZD/0oFu7KSVj/lhH0FpVo2Opi0eyPTG9TPLh0tPgEsRyV1X4l+cdVhVn0dz
alC2UUeZZaXkJlwor67O4lqyEOPJYxqMpH9179XQLcdTqEy3fjV3gkCvwYSKiZUtMDkbCo3qI89f
XDaaQBLRQv8APOuo1V0eA+xp/tBBr9ZytlFUkWYhP9BcBwLZwDf+CSWImBnrOqBPJbzd0NSTDn+u
kzsj5M8lZoYlOUh7nzk6PYln9q0sepwB9TpKCvjs3DsPaK5uRGd/KnfEEIgWxoHxEmfwpawa/v9w
3Rf6qjFFOnUZyBhgpIsQIVg2wdYhfa7wqlLCrWtCempWPzWCDwEH94xFbWRWFyOsu3UP/Njh4YNK
DuCrb/TnNQ4agWrmdgVykksdqIkWUZg6nkQ1NEUqkewTMTJez/JbFDZ5+/cJFDjU9prXaEMZRKGW
7NFrkq6nNfln/ozOibGC3Pst1+a6sT/IVX7TNEQq3mDrNjXggROHGiLElYrfnkn8k5Q9NZoBIHyP
wYdMco0C01ybI+AK7kRPgJ06Ix/c4N5ypr7HnGFiCR4YcG/aSg2+FmOv15r42iPPEO9y5w64g9dO
lJ6Nh3uBH6qVOVlaAKI3cI23Ug33vJUPzyhbfBxnbFuuTgaGehEEIyumKbLJx8tZkidAgFuOWUyP
VwfMk4FqlHQJTOFAKTmfxh7Wy6o8U2QIKhZiiNHFNv9YX9ZLJeKh6WwaTV5/I3XCjbba7x8z+G9A
Rlkolhjddz4+ytP5KkCbL79oxVfkbJVP56KVs4waYpG+SHcWhR8PO7hR29f2WLdvRA==
`protect end_protected
