`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
apc1CnSO4+T0xR0ZUVP5/vK9/mRe3Wp2sJuEVvW+2+GND5pkgI2H49+dTGseqdM9G6e2afbk47ka
VrCpABwiaQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f7SlyLV9nmSvqRCBSsFRHrw6gkFzGs6bg4K3McbZAPIQ/zJdiVM7Dc/Gm/Tv8lk3S3sKHgY2uf69
hQBxDm0KM11s10OJwjja3SYnKnNJZAaq6y7/9Afyyy/P7atSjGgcABH8nEyeQ+XCcIqEpYLT6o7h
EUvF9D/ONa7s0EJE6Mk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oM1ZoDb6aiWXXQy6a2GvOT4KOtd47FrXz/3g81u3MVP56zMR5GtLt7ryWgUn+rVf3VK7jzLiGQsM
w4MmQlFxy3MpvOd70DRf4eFrAO8knFaX8NelViGofkaaEwXl8NifzOmN4azyihdDxkszukClLEIK
SYUCXslR7lplKdOPsIjpOD1/Cpik+qHl5enPARNjAN5Tl6UL6EjV1qD68MYLhbUMb5jro2lgTNge
g+GoLkProEdkEeWXwqYRXcxxNpUVviYnaaqWEcPZAoei0kmDtX2PAvaYRs8sMIpXALSIz0GuW8DF
HyKVPa1XbYk6yBXiFqhGxRAcVAbrOv7Kgm6Pxg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RSIm5aPJ/tfv7oec9MY/ZsD+wv1orhtjRU7aQhwCXt118o42kowoxl328s/sJBbyFzCw0dXsDB21
6VgE9zya0iIr5nIEPfRr/74p+jO1YStFYlh+BHOPG4dIS/d2dZaZgN6dLkUeJV5xsJJx9zFq22iE
2CO8O9i5JJYI3lJQWyg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pnSKQgBiazZRJltZY1V4Fc87kxUj0Hht5jEcGbZ5u9DDWvUhOczLNM9CZh6kMav9h6qXXCSedMp5
IF7vxEfVCpdGdEBSwAZwRG5IPGkYiVUbYcuSJ48MlSe+d6AT5qAVDKhchsA9elGf+EDj3DMPaWs6
mNU4zA0B6EZ+0JAZlxeIr23YHgR0/H78dxw6+SVqdPMF8mcA05Pwu2ikVpqrc+RnkdtMILOREiOm
nWZexvCDDpkEv46NGoi+HeJTwqnDR2aWNi6ji+ox0k8C4qrjayUh8fW6DbZM+eykbm1KRK3XlUOV
zsKGT7nN0aVQAbFnRiaPXwpIdWN0hnIE0CdonQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103072)
`protect data_block
YvC8HV0/yF7t/AN7gkDr3yiqk6DKwknhJjY3ViBB34d0JfwqPE6LJVw7rXiA7yrCX7mqBUKocCcv
ryujblGgAC8HZURkY3ywe5+/gyeqpNzIsWgvxY21uscbvQU7a3pH3B+QsPKRS0q2ra/jwUUFAETu
A4tyKpwuU5z28CA/YKk+54nTNOJaJ7/jzLskx9G8kKOZxrvB31lXYb8U6hRB/nGim7dvPF7Su0Pd
K72GHw1zLmkDrsFcWuSYyUDbOtC4Sv0drnuwGIipehgM9NWv2Pl5nYB0xfNnCsIHt07bQ+jv3ygo
eJiUBmzzP7ifKWn5EICmFft8SO+PsjyqdSNHbJumBxz0sljwu7kDS+4EpS2vsfmsM86jKjOoY6D6
aCb4SPYjVo053Qf44WO+lMt2uugslMhTzFz7GvI06otMmiWj2ssu8h76HHT6H4LvuF5WFj2OYMvm
5SZ3aR/wPENb0UdW1beJdkDCkkLV1MsXQZKaAfWnhu0jEA+nzI/4pIipF1o9le6ua7WqhaoqZ2jh
4tV7nSBuoP7W8IvQAuPWINtwrWAhAuOLUKZX1D41INgLk5hIAah3ZdwpDQe+foXUzXFOvqNhnj5G
JFGcVU2+jAocEGMR2hbCgR/koCSrjfb8aS51FQehabLJ458uyF9/cWejfqDSdg3pK8CVcclCxTHt
2/O88RB/naqS/c86qRNtG3gnY0oPkJ2fkrkwGYeiKizkWzCgNj/Ez9I0nyYgPbW4wR0UkQTXIz/4
Qho6F1wf6yX6unsKRR2zUEaspE0Ww4/G/0N43ViPCuNaJR6tLuDSVulVWjYDZZIWpFJG4lWp8ryv
QLtCLYRewCRh+H7kheZ+v400/H6Hy6hUgvcXIbmGWq5voQmn990VF0Uq81rEztVaa18iq91Vx2oj
/eSXD8EplgyVgrDM60GjivRu/FAriWY/LSz/i83JpoZHwMmleZ0PXZcnb7z2009TAhIpP4V5GxWf
v8xxyLczO9FZU/MxMstEa0LIhXrxNYGshgIgjfveIAGhclJBYqO4cYB40+NTZEbwnDISuTpj+Rq9
bxMVNEWV+YgbSI9MsGC1UQJSL0FXIA6yTqy51Su9e5cWc27e2/3B135pre7Bg2VLkFJazNKMdp87
EB37w4WIa8gG8MPQ8oQ/o5X95tieDQz3mdayB6jqGRxHstpjIQKIkB9hYL5k8EMlxOc4V0weWj/A
Z6/vKb0lXpfbK/m3p9vHZI9M7QWu9+fsViSoEj1hCUncpCox317FmStZHP2sug8n2YjZvYzhoBp1
KHN7Y3/iWwcFetFs8iCrQLnFw6BfuuY8vLmGx5vez6IejhTpZpEMxGbYaQ5eF3a6cq0UPpISGWSn
Na0Pvpid3ni2YCn8AuXKb6e5dDVgF8V9SHbaQHZfqr2x/4+lJP+jsXzXOiTCzl4C2UG35JuCGjLF
c2Ol1sOHCgElQKylfrgZdC9UP6iHfWW3h3gRAT2/DkLMEoWcLwKJjeJl+9M720RhSmtdWBfA0h3C
GRF+xKyzA/+NiAvMfor8z4PmWdxxchhxmWJMN2szAqpLNdG1g4sVH7mY3mQ6iX7U57v1ExtRUaNR
3wGudG62uN5ykmCc33NA+HdT4tV7zHysKVlZjlzL9FjeV9qS0P7nx87cFbJBCdW1OUvbEWfl9Qom
0kji+st+WFLZA8fwf5nSdMYdSnt4aFcAX6MkYLIzGmcTCCSQ16MkxcVfdx1LGSjQabWLye8mljvB
hiT7v4XtREiTeXecs2+qN13VXA0iu8hy6dcylM2urYGWmzsyyBNhLrkj1jjwhLbIfE0N1E14BIN2
ScGy5VcFpdNylb0thiWKbpwPsDi+EA7S6qAWI+b7uJFo/thrSeqQob7km0fR1uO1P1aNVMRYbgAp
brFascqwb+lLT5Y9P+C+2gQYaJuh3K+dCOLjK7g9kDr59cqMI8u2e3vzwtQ+yZ08nYKSXoRgY9ng
b+aR3pskW2eCzskYjv3RoC+21h8APeTupa4jmKa130TFk2Gotgmzn7OvF3ofDAaeK87f/34KMzdp
hzsuRM49YJ72Myzv8hd1WS85gCWgRnCXNjKunObCpuxF23MZvLIR2mhY8slWRma+asVYuWSct/J1
0j32gi0hTDg3om/HR3hIBIDbIhZRomB2GihxziOn4wfqiJITY10+PodctG+oS+bTD3Utn03QNwJ3
SwTdsar0klV4XgyPwitiMJsmxqTFiGW6YNF4myJGWb3GlCIQvncecH5Dt/9UWXbTmFEr6CWh2Ddj
jUVbnZpWzTbyWLZ0tbStIp6DSvoV1Yzm2fS9duHud+UZtCwiZ9iiJN0mDPcvnQ03X1VnX9X0a34W
jZx+Ue0YrOtbsJTlSZirj75LRZJyTML7v8ZX5v0noDZN+1ZPlqllAybo8fHKtihhg+RG9qu6RIJn
pJ4UPPxVbSvbGELjzxoTmJ5koao08cuNzNIc3FVlh/gLoYiv7uLfbF5i0jvu80fqbf9JdkekGiuK
OH3Aw4P9/9bs9NUh+qC5n9U6f+qapqi6Dvys2x1djTyBYvjbx9+d628C197Im4QZlbGhJ7Fa/0Js
KlQHdUgf1vsHRUe6OJmv1kOSd99PN5xcsp27fG6Kh7sNmaewcNRYVInrcTMoHeZPIhogkCGwhZOp
92EeJO+gAJTFQMhPEl2VSpVeOqC684dR2czAIvJ6eQTUsD14AC18+7pIocRVhl3NsgHmY9eQLX2c
UP0sWfDZNrQr3nVQINETVdBkuOvosEFOJDYz42gTewT9POpeJRNam70Q1joXS3jC3qVHiFJ8IM6s
k9moR58q7XdWb6do28s2qI0EMr8XbH9lEC2ospy//xGb6hcIdI/uHcJk1fKDIRpRJuik82+0zKrM
jHqIK+IbaagUIDg0BVo0e8zMespAjmxg6iE9tJdjfDWZJa8EkZ9B32CxfpkSEte14ZzYVaQbbd5q
tM6QG3WWQe7dZEeI1IMVSzragNOscwWSQaFV4fQoxol0K+iylJ4il8aI85yPTN/hSboObIte5yv4
C5V3Vn9oT9Vjdy2lgsO1vPxB63MgijepJt8icq5U+Nc+0jUSXJc5HLm66Y3+Xsjb/rpwf0YknfGc
pEYJRxqH0dR/P0Lwg5Wxcrn4E7YaJiopzpwJJiLsMY3BStOSteHONI0Bk9OXlBeXF4Jr4mIy3muy
pMadaIWMIrNmSew11FG/QLZ84FfDvcjpN1eSuf7a6zJzyNsa364guhed5idseXII8H1Cx1PYq9er
PP7wRGLkTXjavwZTr4UpV7m442WPEYoc1YT+8oxrc/Mx8RwW2POjOsXH7yndJ9xsn9Se94gJiFBu
nS5oqzqi/OVH4QkrjKpv008lA75pDPwT6d4YnHoP3TUa5zBad8mMZO3p7rGjE9l5UmiLaf690wN6
Fl/8Zi6thW8v1WNvcwtMrMNXPBkQDf9P8sEBUoyGo74yl7QowliA+3HsnyQg9P8WTjPSgjZymDP8
QjuNG+AX3ZzD6UU72oyqoZF7/wG6f7271Ek3lYMGNLVLFLGUBa7pFhs+hA2wAt8p2B1zihGippC7
LOVYukmv8Q9rqH9yX7R1IUODhQIR8VGRR//Lw4BxFAqol93OxVzENef6HlqV78LYFX2SsZPK+hEc
FG1dtcE8uxhbK68dlllih/D84ZyeoGEh1NeTxTpuPYubW+ztLRt0lgwhlAo8LM+53U54Hz7qI/tF
30HBBc7mjdit/NQxmE8Z+cggIv8B5gMRzSRQ0StPWB8ga21nbcBL0jo80M8kqh9zOfiR83lh6Osz
jLcYyOpvKuEZ1UwJOSn3RWc4wwNsH3Wnt6k69LmnwKDkusDplJWQrysGdNOEmhNa4/mKOHpKdqpd
x/mLnIJSRX9W8KauB2TE9oGgxink5xQlAmGYhu/ot72ShO0clCYJAld1Ab0/AZt2eIdATkR1PRB3
5xhhKSGk9j09E9yraG3pulPsXx2nCFg/JtJiLv9K89YgMvx+VZIaaHwk2YvGoNuFGyMWX6RN+QTH
CBI7Av+9uplgZtxx1t3y73fUeDbNrbkyZCVrcaN8XcTkGowpXoWLwdjxSb+qg3jUSotSXP//mS2A
PgTB5ta//JDbmS9u8blYiJrJ/sbjNrFJ/rVNm7c6gE1ww2GU3IW/6BpRrbIHeuQORiwxUVc0QvJS
RfB2fNWRe6UIkMN3tjh4AuC1jMNsmPb/BhzeOK4+G75wUqiOZpH5jR3yxke2o/0VZRXQwBizUCal
UWXndSOulr28ti1AM18wDsiwg2CC7W4BVYdemfE0cEqUAxVafrWgR1aYgcYE8I/+xql2a9tsA6AK
sDUUDsgxRm0ULRcM8wTgwurIathM1dIpc1qaW7fmjMSnBI7e2FGvWF3XFzeV6jnneU7yZL14qClY
jylnPjoZJdyN5XUEweUrlDG4x+WNgWIz19RM95Fa5obfAT3t2VTgcTi5J11I0TIaIWCFfg7JT+MZ
V/RQERhHq8ujXqQjfK+GQ0uFfAAfZWVXZMp+kjlWKGQOs7zblKMY5ROoTLepCOIRasH8bX7oPoyZ
Boj1j0gCkiWIkSbD03cxqXQnHhwKJExE4urKkSvZWAEflWgmWtgceYKGx2TOjE547yvfS7/dC9/7
N/osOXGFyhFhr1LmfwO4Vr9iKuSJFjnL3V7HpSL+/H1Tzo9VhYFe3BYMfvSgWaNYc5m28JiiIcc9
ZZdHSm5B4jgU+JARbYTeHRGOv0kJ0Nba5Pio6E4RgqNck3a5QjxncV/RCW5yih1uBjXt+SSahWwP
pc6U7VgTE5MDfNriYub/Irc1dB43Y+BVNvjl22xcURvsVDsgvSokM9ySU+8FsWI48oLeLsh/ib0R
eeV+TkmCCRWzK2INF5Tjsp4R/ObFQIWtfwZWWOmFc6idB2yBGg4rlHxNyQ+VzmCMBAkLWqo04Qq5
82q58CYFoAEMzwRa0ZyklULpKWYY/pzFnvwqsbolyrxF6uF5mGWQwVHJilXxpgIBhrK56P6pNZQV
MHC9YUeNes95gaeWy9SwZuNI0vSxKr9UcqXz3E0u2VS4K076Kl9XQJIOIAurl8SMVOh/NogxbmF7
gYX++2PLo6+CVjNHTayqmJHRiwi3h65wbT0Dooi1JYKeMK11oEOYuFJuHNcCrAEg8kFzArsn5I2y
nRpKRUOtZqD81jpkk2II3YqZNOLeosNOTgw+ofs1Tuf+T1AywuaM1R2M+ZUMCEiIVEJd6q/aYAUn
+vReUf4P2iicBr4t5NOKtCSdrVqmvShDf4DopYwzMRCuivxHsPlpYYk4cL0KoO3SmJEn00fdoV6d
pJmI6Eyheoef8peZdYGBClT9grK5iNcg9bQx8zCkbLTAJ8oLdIivTops2LKEEoIugdk92Pi04b8a
w2HJsQ/1ANSFf9fX+bgMj2ueP4gb1zpFdZI4qGu1nSjNJMRGOCiuUHKJHdlX/CETTa4iwxc5g5lP
+ueCxHe4GsdJO6RYJt2XYMIHRO0PpwsNVuVOfXtyXgfzurM9MuZjh0X6YP+DsvFKblPuO+tpPdRv
kmE2qggmdOIhJ/AkqFH2QXHLlZJRZ2tvfW7QvrPR2eBmNG/5b/+uXjPgPD4o4bwfuHcunpJy4Q2C
U2uiRjO5aa6eHcGPvYIikqblHOcWpB7bmAcNi7VP/dKuupnLvz2tsh+3KjGepVcNvST7zpf6sM+V
QstdEf8HZkNUdy0Uxm2qGkWit7X6wHo1YOPYBumOcTzOruXspj8an5DweNg+B5d8dpWd2TPZTDSv
O7EE+nvlsxRzIz4kzGlMTd8RHSVsREofaWYSp354j0s80d57i0/q9/eBEot6J2HyDdrTqiPcyUhs
YLGIvqjMamGB+ojNdebMRek6RicqHBHAvMYunbfTPEst/SGNvA8nPAyQNfiBbB1QgXIGf6axjenC
Ltq+bJmTIWcPfOx9sfmUyWWQF//XhsH7+W4GdJM7TndJpvpI2RgX4TE1Z1l14XqgA500x9n27ikR
a0cnIIErk/o/0vFEnypF4vHp70oTftbbWQs5TiQ8KOmfn47+l6LfWVB8HDIpa9pr5LbM0A7jZPJm
iNtzHAXbDpFtXQdVKU/zqUTuFCg3q/qkfQ9iQSCvS1Kz5SG1rpSB4gVELuXB55sKNB1dM4MtasnF
cyn+vLUBTDMg1dYCaoan/8p5q6dOumnpN25Bqb55PQrSz2tWgeW00RlHPIa8wC4nP5JfSCXnf5NC
ubcPxobV8N5pXwGiTfu+RfNmZFXnGkTWiSr7OeJrFkVkUKpDPS5A6etmRs4jBhvrylI1xsOnjASt
6CNXMBgBr0Lh5AnXStG4C67r8Jhul946waelnhMSU5B/wFQ9Fua5Wo2kst63RqSsB3KXMG4xITi0
qF+urATjpVMOwLS2+qbqNv6eu0m2OSVR8a21wW2DJk9CtCr83XNA2sXT99IPHStXBfJoY1p8hjcf
ZuFsqrGsbJgMqBD2dOziQGyePx1VvLOjdbu1O0gSWz7R6pUUhZhdytSy47A+CXr9zhCps/KNLZT+
vs1616REnGTrBKzIicmZ1W9tpWgWn+8Kzen6r+rgNQCpNnw3fjtwa22fkc1VAMxmp8+JN+AVImXL
g+Yu2FOXnfpNffDJeC8IduMJjWUjW7QNHRz6Ij9R7Brr0Sqg2KrmgQmugwlwulei7MFvV2h/ef+V
ZvVG3TlhqhV9884GEFMsYzLArbYvuW/nXJDRPZarZ/8p+rgqp0uk7BN1Cyj9fWWBo6fHk0alDq5g
bpzB8E6a27/zIkvFDImiHUCyA/zIcGu1vYAqYc5/+Gwc7b/Ev4Y7vNgIUhtzrWi6sZrGfwFw00QQ
ZaRjnP7Tl9jnvOQM1i+aac7A5bmRiYb5/Jbp/cavVAlU0N89NXOqDl00gmJNgRpw/59zwCUv9AZC
8sp/Tw9gfnhygBWUU47x04M5SR0h6YGvPk/gon3JMXRk0noN9raXGx6y+c5A+dBJ5ByRuEyRsiFX
g/mk3KuJmO8vUs4c2igsdq+IxAK6SnJOh+sodIxVY+n6GtS9YBm0didrfzPd02TOUQHuPtJlrZ/J
/mIfXlG9F8Y6Eh3Sxd0pCmGnbuEVgM9bHee5VGmPsJfmKAZrMk2v6PCddJwhrmtZzF41+1pCmgGE
LZ/Lu9dGfoi95ONjLm2plp/s8FzSavD0BMmlfidjBbh8M33awQa2oGhIaXZ7dznCTildFzsBdzAZ
tN2shR9IZsbKmPou1zycgyWzHvEx9B/oIJakJBMKVAMPUuj+SchoCAv2fFe4artd7k35jQRtJ6kg
GNbB84z/TKqEk1cWjbmFHO+T/cvtosNczsn3b9E62yqFp3rRQd20AGrkRsXOB2PK0D5Ikg3QYbTc
p/R8IJqGlwfMC/bE+fwlCNmd1OYx/Lsb3lf4lGrCiLs29fxvUjG+CtabYLh9QUOeVk9I6HwsVLPE
gs/5GRSn97G8bRlnbBDLPtQLXo9PYMdxGvU0H6h0FBhkp3f2u6hxAr7pJ1/1RXvqpMF2dKpJXuIu
/879B92iH9iV6tdNzxU4o6KqXOVxv3aEJWV8W26kgnqF0CDzwua9qKEA8DrqCpcf7RVUFYE96WE6
CrOdJcY5lGQcoPEq+mRIRh9dsodBB7dB6X0PLKybLICncoc2CixI6f8YCCFQgnKpbg9sha3/07YB
EYL2UUsqEdRAGgjaCxWHKcclreZVdwzfUwsxJ15AZTOVede2EKwOWk+5w6JmblK3MvFHLK6xgqTl
yFwIZ4bjNAdpwa45UhEUF7EqDc8BN3ghOoH96XKID1I32MDc62nzTI/HLecyQVLqdqzaiCveW1ma
qImh7pWdt4zQlLYQ7+DwkVCrm2mCRm8sza3Ygwcp2iY5khmfwjRKEk8GjQHY0LUUX9mNsBLJhj8a
LJNMu9U6JRL+sw3UVQgazIwYbixdDuAJInU66CaYzKkdj071tpCfuHga9UdPGURb/Itq8meJnMfo
5XDVC+034Ij0NhmJBQGnBl/YwvKWh5XFW9b2vgbG65BgibAdec/NmdglnfqCqkp13e2ml4ZuOJZz
pl7bkz09S0I8vy89hD7ituSKb13Sh9QUpEeOxvPwgFOpLgenGlSI0V3p6JueUxGzpcmVzmkFVhLe
3cYtKxPH0ECSuezsPW1jZnYkXZD9j9ZhuvwGL1mpeggv9riCIwnpS/tGVal/PANF1e1SzUsfcuUE
IIpsXew9j/MJ68kP1Po0zjBs9UyM0c8jNX7qwnTqkhI8YBy78MKXCIL0asNdc+aniun76TPbQ3dp
WJPTwhUVSH5R7justLLnx1V4v905HLrfoRZnTGa358Ju1Iy0g9AQvg5lefVYkH5JLeenyHMvde5n
6iYGfiD85PiYKiz5H6fIRklrgsRgAp6wdroDpOZoaVrpsAWdLXvmUxA8xw/myOO0wPREG5FcEJ3+
j2NcPwz+L+aVdWAuoIHkvy3e8bkDArfFBOcnCrmWMIIcE+1MNWhvm27mFF5PLSxBmrYpvjeAxPSw
WSsub3VcK6+pZpeWujgtntoDzcF9BTolYpSdVtjRLw39HPIdjfvYYUs2r3+Wgm7/DLMDuchdgeah
VbkaYuWCMO7+oCFxLLoFRwm1F75kxEWYG7f90jBQ1jNOqfwuIiKYmuA89DFo/oAhwfKrFBvuEjSx
yYoxDFMljMHlFT3bfGswrgLa20+EkpgPZ3uaM7QiN1dWrfQfe+EMBuk89xdjKMFmPSZAI154wjCD
4B2mPzG1+W8HA1lBPw3+v7eSne8MBbLVqgFGabhDVBqdlgKN7UI856dBM3ALdCEkcNaZoL6/wzTI
AdMk7aafKG+CqU8z3v6hEgPUm9jf471rT+wKs+FPJQC8hJN4WAN36QQK+tuSSRDOvK9sf/5+DMqp
S72DBg+dUnebzxUw9GNWGS58p+SMCpDrKz6gksYkJtT4ew36KDpb12wqbbA0uHP/GdoSRGBc4xjo
dq3Ze/gV6mG8Fm6m3yCJZSFnlFL62QwbPfWKgjzINl2lXFtuMBd9+N/TLHThB0ixTOwKDIImakGu
xEkDIpWJVmXWvCyOMLp0t+RGxGXFM2FE3283BuZp4tFoJTOkOy9ENcXmwo05Z0EiFj1j7a6E4GVj
kp4hm/Pbbwo/C3HLfRAH+Vx+H4TEtYstAQVOb6B6Wtbx+2zcCN0HZoXJRptWYaQ1ZU7TD3QcKLXm
16JAhlXpFEMmedxoBFYz6iklQpkL69d74anfZYnKTtJxtXFhNGP1SxMECNReg9LlqRYBGs85MmQV
Z5K5MfdfaAm0N4oKncJWs5zmNIhvBTuPaqnvIPYwBlht/dOA1d0U6j1P0Df2v1vb6nrwdmS222d5
a8W0GjtmlYG5CJ9mpyQPCzehZP40ekUbOoi2M9J4FswuF8EVBkhbQ2Mbo1eT3SIE7kDMHm+yLz/P
JFwtKpRASOvzgjjdpx3gReX98TonX0d06pAIx96YddcMXNxjGpg5YY2CjHbOG4uKGatT7ZAMslIv
VU+huOG610du4XWXl3Fn4PNP4/YXgN5ge42NBb75vXUgYACjk5ze8HruPz3fgTrX7I09eYaIYHI0
ygkhTIJi98iiq58Aiw6w80DiOCPjqPsyu9DIMuSgT/j4mh+zqeV5PtFHuFKu34IkFPH6LXP99Cw0
PLJceFCuaQgB/LOM7iTsA7jH9iRaEEbArV0ee/MT90JuyDj0uYlwYQXYH3/VwctEszUCVuqpBqhz
Er7Hxi27GBY5OQf7iMXdC9MwTGfkIVRYGLgPAdugJEI2/QRzh1Fxkrr/RD1aPARm4opozuINzRdm
YJrsOci1ILvvNiPurwkHt4QjKrDNrK7emKk60VBPIFtJb6+IO/CdbTV6a+6aM/uSEcXqoysS4rup
SXtXwvZreyEOYVbvJcDjja5HFL/skk1kN/riLfrYedCiYdqzmqYi8v6P+33+zqcoYFauOJt53iEU
VdHJnNZkDEDzbk14YeDhO24DtWtwa5TInRQcdxqX9c28/XyW66ZYmdF8EMUyOvGO74iDL/jig5L1
Wj8Xm5oQQlS2sZkfw7Guc14TyvV4r9YLU/V8UqNG7QNutBmdFy/UNMkg8KyohtkfH9xPpJ9N+Ggt
0FF70ZGSvZnwhHhquYYodv+2eZRGJv01k0ZElijTXgdi9cwveHLGzjdEeydvOS4FHy3BaUQuMHxi
bsuTT+g3dpArDCay+T/nIAYoUIribpnf1JiQYtw6JvWuP4by8NyfyhgCLDUwN2nnxB0Dus62Hkfq
1btbpHsctq32V7Dp0nkt0RKQPzKyaxuTrsOnPwJuZQoCm/1umFzEeX9fCVypJZzP/jjfxzGLCQ1q
hKOBWHQhc3tf1cflEqH4c4DDhmHDORw1gWwP+YeYdWjLU5Im8fl365Vp7IhpGuK+wSnDdN2h3ZKP
W1DMo5wmQ8Tt+Mm6/rl7WCOeOtTVAxJhTbLUEEknawvjOMySmiDrPZ3o1AUxXd8md7TkhFRz/UhM
t/yAVrMKsJeG0LyMpyjcC67eno20In3hA0egjGx3Sn/5wfr8xrmpTZvlb6W7BHlSejh8JZCrq0JR
r5gFvdhnz3kyTmJCdoXMUsbn7lKtrW59V/FcdqdYmwPgDBJfZK/2J+5jbT5tYOR0DvZ5w5M1uq8i
0k/yrHjK2QtFhjN60oxbaJZjhFR8EgT8s3J4DJJIRfXaWwQFQPEvz4SLLLpH3dTBXcAheUxM+MAl
q1Sxp/TR10NcsOIKBobia6BKJA8M4yN3wui6f/AbHkSdF/g4YuSCpxRh2yqw2dX3wa+VVrnKliaH
nHg2cRya9mKpTnlo+GimSHNlSBU9Jnn9RFaVXwIgSoAPHRGCLgUck8Uuai89bZfebnXt+YiPbg9o
FpyK4wsoXht621V55FQ/8L6BHvDXmpMx+97h9R0Hu71YnY8f3qp3QmJCqqoKeDmGD/dqFMEHZNAu
/QtRQ40lH2thbDnUFG6hydt4Jycs1CQziCY/dTK/kFtgjpgkYSlicKTRBSFLSI1rU5xWjY4en3TD
cQaIt8GqtXQsxwX+5wD7ipmWDA7ss88zA5wNyr2Y5/2x/ePs/nT/dsUBlg/f7fAAHjL/kgcHovg4
k30RvRlUKiWJw0IB5FxPrMrRcKVIEvbA2qfH0bPvNYqYn+YNO/vGw/4FTmE7cPJ/w9nnIqN24IOQ
Slm4mLfvJ3nw32a+reEyIrVfjKFVYgXmSmZzhDaCJJCxY0qqNIxKN7XkLcOSVubHdLUnMPNgoKXm
lfR5dEustjRVbf8a171Ty2+YDWEd9DIRWPgrV8wXXHMG5AsFuNVrTEGflQVGEDhNAPQV6V/TvE1t
yf7qJr4PxGD0q6PpV6vBmEqAxZfGIK+aA41y44QwqFmpblCETtzfmUJL7Sth3Pyh3OOae7PmAuYw
ezWfw0lP+2ARaVnUO/BSRXU8ee5KiafFCvnzwxDv6wyZg7DHrenjV6SFm1jzZW30Qo3mPimRaI91
kVKqdholJaN6Muvq4vbQNJwKaUCu5ckMXaEIuKmG4ADENjfkLEtNVE6FPbdHYyjZVIN8Y1Axm9wW
aidyh5cm9ReNSYGZx9bDn5ZtFkKd2eo3nwYcVwoc94HWH/wlSjvFWVio9BUUsr3HMmA0zBohG4mA
GYh7pFv+ob9+S3oIgs6Mnx01+dt7lg0SmA0oewaBBh1wdxwg0XnW96ED5HLZMhzTzviwbPtgi/kM
avA2A8ZQg13zRdRmy3g4b/h/CWAAPbOJIwARMO9VesDnWj27LTJiK0jBCtpo9KD61lYTfMXq5qMe
KmO3dSfwOljIhKPcKQjXGsjjo9bZ4ytsGJ3Az/DCccREFl2l6ayQ104y+yqZFHWuSmuHJ3RZmq2I
AuQtjNXdl/MK91RjQvXiPZHuW7/POwimdlj+IoSotSlO0kecOcZPRZ4JJdoKegvpOTxcwHGYDeDW
g75WXEKFwY56YIsDhGOxpoICePEZWOeGwzPSOO/sq+S4e/HSy8hpHaFHhTJ4HP/D37MKGUK0Ushr
BQpQyypmB38lROtK5Tk4UP5avg0r96cF6ScshTQ+2v0HnhxT2QvzUpS7cqwoUbQhgHEjmqdLXV7u
iKlwnqP9Lb+Q6MPdmwGnsdPBTrLqXjO7lLYqx9be39lidQE7j8xbUapeRQdNvJfuSdemjcjF0Mtb
61epxTaiAyo7RJtPe+dkcPNAqbWWioYws2zP4yp5lLj+r4Vpr8P4Hzg693/bGfihC4kj+20U0zeg
VodF1K+wJa2eRZb8SSKTVOvBHd6BYIbP2LUMTQBEgxB01P3Gwl+GtuZ/teCbuJbsch0EXuUeQSYB
66f4Yr6ULkK+Yr166IZsgeaYJT79Tm7ME5cnOGilz8UstdSEKW9Jrc3qR6bXbOQIHfFPjEw/6xEO
lzaToidWQ5DuhIcokkfZIPHgtaabjDZwkOtC+KiQK0YHWRazAB/AaqfYwctmUpmjLDJfNS81P4Mz
mXvO4dlQnEayDPoqoLy47yeDTKb4bCGXG94/Rciy5OcKM00nis0lkMKukPZLnoFN+idTeQWerEI1
CamC/8Nc1ob0IyXaiixs/CH0reMCfLuZoOyNhCDxhmNTRoak+So1bUmbGfqg2PjJb1uVtncWTS/6
JKjUy242FkPgryqunV4nTK6bhDwlmZo3+JTTprQNtbCzDMCq9Mm6Xgl1Skt3HcyrHDmLgMa6vQvT
nbi6PixgaZE/KYw4TfaWKYzG2BPiYWCvLdbEmGiBHuR5FOHid3RRQmMxJiIxzXzBTvnAO3oBcSbn
pF+I9yj8qMbo1GoBvPFtRjOlbcqFwPbNx/DQCxTj9+Jut4/MU43fDV7rcrbTqPD64vsmyzqMITls
uNqJk6ik4MJwn4HJZ2iqp+zmIZRISMqrLrEsozJ6CYYwIyGuXGdkvqj7OnWgVLRU3+oLiQD3eDUS
jWQWq4KKQ9NifpGTA+FLxL88VUG0Z2vQgnRMMyODAPQT3EP5Sl/F3PZOCzTFATTuc1EiarLUCIz9
ZfNc+O03zShzy8kXTqdIVucrTUiX1YDoEPTjb2cnzUOuvvwGgWjX6HysCJAf+XNVIWVSyK0qDC4y
xdRuE7AV3WtLSjuO2uLIYlRALF/oGtdomw5llFobcmw/kW/2Zx0KlHdaZUP0O1O9+oG8s1RTsyID
2UwcUUj3P0n6NPKdv+hQonWEMXqLNjB+HuYeJvnmxDMrrE4YR9p4P1UYG/B5IgtqrYI7jjrg/6CT
LDOGOoPLo+WWYSjXpWN75cuXimhWzXPU2JVMlKMsHna4c7m7Y9f48pO8DQKsFgrRapD8CAoVHXJy
FOfuFzZ7pm/csN41ifI6xW6b055G2acmrcsnhjTSnmAh93uE0KGiH0y8MEHcrLZtGN8/dkfR9h3Q
vK/fFeFRsumiGqnI3/QdjHA7MmQf8UaQWVlBeD3S2L6H3lPA7UhXE7dOj9DjFk+N8PR5ppCRBwza
eN1j/hEEAeZ9fyWFBMHVzMnY6SzlegZhR2dEDgz4lQQd3jpAYZyGufDuw1gEBcpkSCFoy62GAwK6
J0zrjwbDjMwm3KgHZSskqeROoOizpyMIAe1z+5B2O8DbI4JIHnEer9ruKtRXhIN3UTZID/y4vZA9
5KazGEopGe2ahdk27ZnOkgQ/eo+UVrvLh0YM5F9tNWrM16ECLLmKzioG9G/cylhxGmAkRbx8pbn3
fsofs0xWS0lwzhy5W2+3QrZrPavhhAYE71EXYwcONQXFW961a1fo9JaVPliBnW49Ehv+gbOgYIVE
qcUQd3p7wn3sKNluBOVEWXfJCMt8oAlKIy6GGnYrkDuCSDh1zAKOJMrLE6xvO3oTW9VoElXxZTzS
yd0DGCZaF+5JL6g7h92441aFicTs64l6ulb1kZUkrCHFk/XiqCCCUvn0DJQC9agcKgLriTlH1hKV
QJjIooKFo32eLGkYKe3XVP4Uk43XFiOJFBLGLtyKV1jBHznkrHKf/mqTcWzFbrfUpbquJSbJyoUc
fASWUL6lzU6V9g6qNe55pt9GEte8hvP2MJnHW+clnplwz7DjUB9i2EqxflpNdNeS++qGuDKdr0L9
dkH0H1Qx+DeJm9S8oxqS5O6zdzUGNEabWF7JNxRl+qv3enGuNQeX7uHadwMjrbKGTMZNgHQgjucG
NTSc12tFfyS3hsAUcnZLCbSlP/At78Kpm8esrAzpOxqpbSHtcf2QPNbR/ojNgFLibh3PVqa8fu76
GqPEMp96i7ZgZKnaz0AjT77YFfTf2XcUvH/BZtwsHuP/LTSr3TCaH1BAzqX7hIhzzHcFEUFneTMt
fsNea7rV4OK8FVrH7f1jyZtEJ2IDMcgO3G1FXGhix1iyZZOeQObWFRtunCwhfel4U1FsAY7s886q
grbL3U/cA8ePiWAfkycub3H6HofRPyW+Uuo29ODLhESAURSm9/amIbIhN6G1sdyrxAL2s9NOUIEV
cyHVWvzMlSrk/J4BYR+7dXQ09T0ScuTWzlmnOGPrsPGWewUzM+NvTbQlc3qIdcfVEgzR8apns+vH
MaXjevQcR4CYwyLaXSJvXbPeSOqMfFlt/Glv/nHDOdwrA797JN11gWAvhp/b0Ncs5t8iNISw/fHw
4vn5zyuOnizGVae0THrT4wN2zHNgl6gqqgx4/EGV1aDviiebD4pX2t6x1BOx99TsG9++YvxIjKz1
QOp6t6j/eggFJ8NbtNO/qVIOHlQzXzTkmA3WxLdRMBD+IlrMqYCrr3EXl5J+VtQC2RqD8MInwH8F
QwzLEs2lTdZdqu3mIIJeb1HEKWvZ7f0qbdVnKi+uRKmA6f8sl6mBKyjHAZ0+Co02K4Xtn5blG9//
B+fKQoMJV/w4GVdCNNLOBBXqkEei03LipYLVQup+p05cDjaHjQeknHTc0W8PEvPbVdKyQZiV0oPT
OoOQksaYk+9HCFA11xgZwMkWS9I82OBh86D0XRVat54aZBZ8xcqbLk2p+M4MBJxJbTazAJF6I4ze
Pc/g9Tk2p6HE+BSkKFpZ11pR/eNGt6kqkNVSXEju2kTFd1wCEYz8UNPGtp8eOqpStZBJK/vm9H1u
owl8lw98oPYYxGUTKy+F4BrZDhxKvVDyQsZOoDmO0S3p1Eo8jPu6KIV9uNB3+IwuRVsUsAJ+OVZV
VeVOyHZ6325jzum6KL3hzVwZLYrBI3OZ+oORWhE7XWIOBIcxVAzxb9WatRD5VJz98/A9DaG3sVpO
flkvvbBYpJW289SWBQg63Y+EFEVXC0sx/vg+wjDXAAbupHUjg29//eqan1hUWfd0foPRg7jTEr68
YJNXtjHbPESmARjsYFnu28XiCCSGRwyK8mNQRKjAlY6gWA+RR0wtLqWe54Ky91Po5vSLJr1XwRJ/
s4DoVhTHlHR2+kgpzuo7AGGriF8ojEl17Rv9cSiv8zoERH2Za1zSbCmhRuSORWhcOU/Ht+5OWTdl
FnHlZVCn/EtLHHYRbt+AMwyqVLvntiVJTZG5egbSe7fd1LDF20odamohSJBTM1kh/gLMsDukcYdZ
1oeoYK08mkiIM1THUQ/7a2uJtrCQgYFS5dL/vSLigpWIWv+2fQYiODtKJCI4nuLDTEwFLPavKbrO
1R/sOx4ENiTJ024+t09bE0DCgbBnOTatfXkHmJ24xFSpJ80m4PFcAI5Hgb0+p0oezQGRgrWfFPn9
hswmQv8+DPeKEVMngkalFgp9avMTT9i5NYHQGJ6QOiyivmZ/CXNxFfjL97tVLynpqSFmCzimaSxk
s+HaoMeUvMqmsIJhITgsdcYpSq2hX1jH2Ri2wdMmPOJvE8xOCXpoI68S64mipVILD8jFhxPPT1pr
N6o1JviIhUDyNmIAYBQaRfTTTB/7wC5y0n5QETwxvy1+3MWavYQEZMJHOXenj/BzMN5bW3F7cmGR
ywnVjIy4Zhb5V4U5+CI7FQ6ttaZdVtrVMcNTkE7x2hJiX0IbVRM442iVn8F+h9kOUpVE5JdJtiJK
d/d7iFmnzq0gNc1xymfBRziTE48+Yry11jEorKjETwy4iwjeB3DIhZCDRBHH14lk6eoX7v2Ij7jG
2EaE7Ltj9kmB86T/wF4JkKLkF2uhKKtMWJQ048dGlmLJWyq7Bd465GrdLZ5CU7f/P1aQT/jtfMQS
w8oE7eUHJHiQ7ave65RZeaKcCG5K37FZf8SSrrx1g+/gAo1wFTG9jl4Tm89TDP4S+aPExWXdNqPf
63lBIU5qZCDmC/s6W1ydITuDVBcyTXrZpmPU58TujkvX9aZYCpkKkUWbyDa1UY8Ld80MZkZT7SQb
m4utXLnhbKxj1IUs12iIVJuwomG/SOi0Hs4CQGqfnTIP2VLOBFK3j+CWpZo2T6jz739I/nWQ0G8F
TAwmUr6fN5lmFLr/TIOWhKSRq9Dc8nvrBCZa8Ci58Qu0u4x34fXj+LXuqRaXsnTVBaGXcyZhZ2K/
N0uvZH35jsUJrA+eTasfLfxi2GZqmRsY8CMey6ps/2FssO8mAgD8Dbetijxydn4KecB6y3J2ADfe
cgLXWKClJWNAFynymqSa+O0LjvIyggoWBN7nuSZLHTG5LHEl4doBoxeXtqIwomV0PINWNdn6jWl7
I/c/mMtLnNDLGwCdmBXbiOHSjTPAtxfOjinu8xWPYYc0OTFwmhtv+Jw6E9n8SjM5FeQMf60+6IaL
keDute8P1Y9dmDy1iDN7wbdra7c4JySkje3IKJSh6dBD7x5wPGcOr5jFhe9iAcO7zsmq7+ojBFeO
jnc/5OuonpnatLRR13RToSGDxlltFS1TFn45vCcv8FB2LrFhLAmtdLJxyIq1yN/mgX33V45J7DcC
QdlZSQC2QT2GVWYnWtRmWDignW+udZZva8lUSgA8nmQNPgi548OFqmzin+gE5KtzMTTCQVDHyxZ6
a2FXrSgqN/wADmyreoS8jIUBrK20X1YEIjw/sdwd28GcV2IBkfpGH2qR3K07nAJ9MhMeSDChUhgG
SGQdf+6rekk5eSDZjx6M7+GNSXvENfc271y/jFrPjBprh529x0nOKECiUzdFZujUXkFF0uC6bUR/
jpPi8VQS41TFXNAOKjYr+hxV3497dZ0iAIgsmQQL3bxuc2doumkavuVOXORnY84xG7SG4q9jNsHv
nziKG6aS1JUGEoJuFEZdrLO+/faYl6op+xdvO6PgxvO6IJwLOkkO2xpeqQ4Kcfrwd9D2ZErc7qrV
RUYv6xg/LLukDxoXPoAMu24F1j7+3lk9AmceKrCKHPwF99yi0Sm0jzpqAaYpSqgz+XeGElbczg1h
WFq2ZNBZX3dqpShwTBuDyKgkmAbiNSAf2m+akjPqElPQ/ZN1PWoYnlij4cvtXK0QSctgS6dc3jHR
1jTFYo/8rnSWU2gQTTpBb6BO3ku2/GjA9w0DnepoCzSJ+JwcdwtjkPEMWZD8IfTEoRWkXm+80ps1
gU7k5hLeqjHNIjrGFsRMfquT+qd/8UdQqZXWqBxdSXZ61lt+JBcVTy/7NREypkIMTYMdH7oFCMMH
GJjJrkBmaYpqXOwpe0H4QyN0UNpZf27vEMOZSshHpwM+aJ+oDTh1gpM3k95yN6CHhtj2Wxh3C16d
FiUAb6oJqjgevpl6DZPv5X64/P+cVvV4A2kXUzhSw+Fq84n4CqlLtQFHOlwWWA5JOqdbH3uJwdWX
0dPO0t/z8dPoHbCKs4F32ftzVhdNIUPp45N3Rl5XCqZ/UuE+cYJiZ10ZeCezY8Q5gBx2CG+nSKxy
R0I+536ZRBitSTvtqo8cpem5TuNtGRTO/Ux0iGkEtgiznTeN63vfgPupbq0u+4tlZ1YPtz310z0w
pb4ivUFinrzQz4wD6U2qpxzJdrFVE2h+LbEv1O6HcMREIC+mLMxELA02rdNpGl5I24TYLdF/PZo3
frG//uiQMz9kLU+dDiEMzSC6opGtSCk2qfE9isjpjbvXUUYBiN/otJYGDbC5iC6yVF/bMfGsxs1P
bT6M77IDZG7dsQUBRVMy4DlH2l7X9UZJplaXCFqYfhZwaBBlRTUNyEr/WMXUVDSiYw0+ForRTdFU
ZHv2lTXq1G8xRRxrmwXoBdwU7VcmMgKDz2+4MN6PpqULMt+GigFjo70LfJ2SV23UphxB0mHXAf1a
ZcIBmjtmejL8vGz4JJti8OtsRUJ5Vrdp40W3ESi+yfNH3xmSP+ojXbht+DddMVjBphUGPnQYZ/k/
q+pVJtMWaf+iRnC2jDiv5GGZzxInaCyBHp12wHKrXlDrjfZrtu3TCE5o3Qs/8ZPfXoUMBS2ZcfuS
w1mYNv8fPh3v6FtuLBlabBLpIlaLJSPtSkxuIuyJY+YAsRBNFUOfnL+xdC0K9a7bpImc1VaO3k6W
DwmR5cKVuca6LOoD5z66ICgrfuAsgJ6zxsaqsYOCQqH4ARqSdo6maNJBzbhp5S1amJAp988u4NCZ
t2qBfQoiwSzR3hoiPGf9Fr2qXSOElO5n7xSpnwYPG9CPANQOqaquK/olEOOgRQQlvJ+hgArz0K29
R4EqwLvWhR5I3q1j/FZu2Jn+i/1DQ5OwQs9UwT+3B4JU4+z4GTHvFGz85KeZsiPaM1Nx3labbaKS
Fihw+l6CD0SoFvzAzFQxt4RV6udJeJytbwBBdioBjIgOr82WGp2P+iAQTmY0cS73HAanULrgMoW5
CT2lPFfSO0avpogyeQE7zfRsHNsrvr08lbX56+l+POB+vQKYAOlwFubMdnymDQ4MONiHkCvC7tRG
WXyjE2hEp9pnU0E6juV2On0oBqEDtPHpyGe+K3D53ENwCMDsgt/PjqAz7qg/UTdPO7QcGOY2EHIL
zXxVoYYYMheULKFCEzKNl9jn04eMA5zUvpIOhyR//cXaMjWOmh79siGEaHq+xIxM0XWbL9VZBuV1
ki2vjb0a/Z6OaUDwESkZA4bFP583/96nNzVHyrtpnU+0W2pQeCwnC4IDIkXGaKwg8ZhSBXNW5q75
Bijf+nqDYkbA283ZCTmhq9pRK5AzjJo9u834D6GqcUOgwwLZE6eHvAeuYroBKF9EKnUZbCHGEn4N
bk1q57HJkgnPZUdG1HqyR3Z/nW71HYXxBNtJxuGr3vm6Uupzgj2adGcyLtrpPgxKoQydRM19JsuL
DWKWTDQKM2/Jwjp8WAZgs9RS0xa5El2wanSwqtV84PmaKXcldmDAdlc4HEn+fzASKz6e/A+a//xq
aRfMUIhgpuMYPS2AKZSd0bBosGKnNMda5GEJYNqZzhfydDsAxzS+4HGzV0y+siYt97G2atPTHAka
eugmMlnvghVt5S4iZdaiczVPxzI0NUm81vJfD20rB/lqQCOgqKjpxRzU5muQHslWup04LYLSWNHV
kBCAeKEJ/1ao8nXxFvttrxrXoG448KrtZUFSyqTJvGozQgCxVrR8eZQNaNkbQ+leNrbRetpIO6Cw
JQ/NASPzQcfjSldlWDW5mdXzJ0N9m43LWPPri79qWU/70aOVHam1VSGTfLVA5WW84fDJz5ynwQE1
BGDr6b5Ty4IOsmyNrvxJQu1XvepX8sc/01B9ede5LcC5ZrBcj0dEGiW1OtlgX9zyZ/3fhVIOWl9n
0u8CmXHUUESO876R6vB4fTMkTXjnWI4fRrf0Km/U25e9hUN980LBgKDQx06v6M0MQ9Se0i/24a/F
wqWyr8R8nK8P4K0xPSJkhY2NBEPav8/Hrhwn/5QWBW/R086Udse4csXVrrT0imnTIzDLi46gyIUJ
XusxdwUnFeju18aw0lGL6sGGPOMdBHdQ9Zm4OQ3/BIwwc+FTWLeKwlPwsoMSw4yreCoeaK3IPNRy
7nnImnchVr9DjDYeDA3qlYizwIk9XAhg9bzLWuxxAoNlit09u0nzGbrdblnabwXYGqEw5LpD8vpo
PmcMOnVbCYvB/nd3Xe6OTnCPvGpa4ulPdLeyW10OOyCMQiucJRWyYh4ApglL12+PNEG8C2fd989R
CboR9HglTJR5CagNfKXkq557gXPnMETj8u54uTjdSiG2KKRdr05ghL/HdO1x0RDeXsP9ZZ7Tq+GZ
Ml605ZCQGhkO/qqvrdq2pbnOhHWZ8bT73V/zL7+ZzqBhkh5DmccWOjYJWilI4mQ1I6f+xJzxb9eh
OcGhHW9ZL0SnY2xciFARPSuBkhY/UOZIM61rtSYKNC8THPoSPxZRqImiofdaU5pMEmQvWjLGPZa6
/QDVSlgVcgoelrTKjqHP7+PUvvF59wmjbciKeq/AfDikxHtZiVlYxOnJe58d3EX6g6OT7j9IzrXs
+hSX2zmtKWTt5FG2Ce1oYU2vaNnZlvQXGECgRBLV/UAJb5SoK0FjJKEh/ZCWa6m52H822JtnSiif
ZwFm5ah8sh3Zt442sLhvGX/ZDeHWT/7H+q1sp2xv3ftZMM6Be1n8fXbgAJFECJwn99NZjRW4qJ6G
W+GYiz66Z0wdtJZHWuDBuvvvLFTxOmfy9n/Y2XNynzOb2gjenY2LtXs/ni/v0TLtjDj6ZwZqf1SO
eOmkHFdE6IPa4WrakTup+LfdhOS298TFcsgzofUp+d7GMBzintmWo1RCAhEZ7U5zSGfBaKHkEjIm
RAXJ7AEVUqrs2VvJEoY1b2EVNjKdsWCmbzlzKUg7sBS5lgyoyq2Qh1i5pKyomhcRS0EFvHkTlsYg
Vkgb1tl50aPsYM15jW48X9L4r4rjm39mNUcgaCyBjfxf6gEKZ7UCupnlTqcBEQ75MEdmVG3jYGs8
DA7sP+aKhs+mv3FdrjuBSmWOqZKhm2xnubvFjC9ddZwundSUSDWC5UrmTCihjW1HtpTL1C3iNMDc
u7DLCNVElXL/DMrz7Cakc2jziC3eK8hFQMB49alkOocUzVJY4wpqX43KwnkStrTysZxVtvlj9DfL
bpYGPcS2ZA6BgyD7/x6vtkHscMtspmbo80OWoOydPX8pwoq5Nd2ysa7bGDz2soFw5iC4hJIBgjO6
y0LKWeC7BsOIl0p103k7tr3iehWe7jN8kEzORxnxpKDsm1pTKLDsWdxMdaYin/NIRUEWTlaxIvhj
dWWWwMcDBv92slF1LVqVNzAgzayPNmOQfhVfkBpOPPipYKGUuu21xnW40hsZjNicKE1IKbwtW5Id
O6EsSuhOKGSoROjf9fTMVJe2VRHtKZHT7YKkhKbur78O4z+cta6+1gGgbgJQHl6P9QJhdXcNJlxC
Ljlt7KemJgGpNBmx7e5D4X4u1o20nLG9ctpSETNZgBxK7UXl6u8UuYUnCjlXmYujHrmBmkQhmuhZ
Witq/r6b6GRsHgsRAwRSrNXW6Ntlmo2kR5cn7q4+IQ3/4YcORf8KwHCAouP/4l6R/2eF+bbW8jCP
QZa5/La2+/RIFNe9EhyTOA6Y92l7pWaYbPdAqpkl0jHTqKocAiaf53uE9DUj/4rbbvapuASXKNqe
BlofeFqf5mVeak6u4ss9ze7z8IoBRdMh9mfgHQuEupyFXc/stzY2EEJTn0mg2fqTA9BksbfRGzYu
1yO2zjw0tXhgio7TpvtTVVoEiEZwxf46qKwyXJYAYeyp1sCyUnidLLyrqf5atR1wBiQ/NZWHHDpH
+6njGHKdjJDF41IIXu1nOwhx2nsW6VvZtDA3zAwrjA0C6+24XY4vx/CZP6TZe0ti0Um9p+IfD2tq
lTJeaO+ZCi5L4Tf35r3MMOvgzaodSjm4MUz15U0w8PceZ6MecxA9lT18XVI2iMYxPajvXIT7ufjl
zdaKnmYJa2L7cajkRZlSTUGRcfqZ8+FCuTnlTcYFGYIJbbaAtL0t2r+V5F/6LrpXJ0BBbBvxUrp7
4NBUEE8AJF074o/ZRnb9wJVTpTIEV5CbdJAAYUX0x4NJ5OLsYMJlq6nAJIKtUCPGLoFr09Su9SQm
jTUAfCmJwJn43Jmm+FUF1pUjvAFtskK09wtUl5pNKE9CnxouJmvJSL9pTfBLbYHyxBwBgSoQF4xg
RMXKKT3wiHEDa7QlQYkR3+2nE7PvTEJ1LNx9bkOqRXr/HQYdcrEg4P9eXXJZARw2p5KHF6lXYR7I
gOcqVR5NqWy51q3EJrUUidMyAuN2ITdrUxBk8A6Pfiyi2cE64Su++jIV1XGokBRYXYMlL2rzJsKK
EnfV61NTmfABfJePg1u3ekzf5Iq3Gg6A/cxR85DfrcQYBRr/Ia2IqkZf3W5IuA4CL1inmGU6bwsY
FwdGGS+VcdvG8AIpNrr19hpRUjbqOx5w6dt2GrlFnmTJgSe4EGNHkXaNEzwvEedTuNzEor3Qn/mH
NgIEA9yzvpGP78gIIUBmQiObnF6PU69A9XD6e/cCVUj1iy+jigY77WmRmErlv7C7dYbCbJn+3F7K
6AhOwgQELkR9/bw6RvLxY+znbnJOJKxbrGFLRim9ZWZW950FGqIbVS65H6XcbWKvppvSigv654xJ
x1I5PLMYOviVwyAELCAEJ1aybMDJL+3uZ3ZkDadZkUnArRNto0ynz4JCJA51XKmJ0/31Z9mnXm2T
FxyGtChzM3hNPEPO9ppGGBaAA685ECLkHYeayzW7FPZ3hGpOgWxXr0kMxTSP3uD9rEOoCEnPwU2H
l7N90QvghF3TTW3iAOwnU+Q+XbsUKHepBZ3RVr+hHfOqk9tSLlm1Ntj87Z1InxsBqnXbhN5+RukW
Jb0MIOGBkvuQSjx4na2PG8IHHC306i7ljn9ca01oeWIc1Gdp/VxiYOXgTdlfLe4BAa9TUatXvjB0
E7zw/+FlrL4UH4nPAzl1cMQTTJSvfwtkR2CD0kCQDqAAqA/rOtE1KaPmIyFsQanJSMJ3C8hE/0Ow
4iWD6Bi+Ww0mchJG1/x0sMo3XpULrHp+wsE1xRhICBHva+3WJXDYSdMWpvg4DIcfbrZejnJ0FPaK
DwI8qw8xk522Ny8YqIxi4qHM6x+r+jivVBqgmkMC8O0vJjM1SRQ282AYTfOaQ2Pq0Jwfrni25aCF
UvOpaGxH/8AHSinKas/b5/cjKUW/0v+Un4afzqZL0eTwcj5DITt7OPKWlOBDtm37ceJd3HHZbqN6
i8m9L7dEiGRTJP9hXV9CiMN//De63Ldl6r5fqyUDYatxkIqX0VvDJ6BfVOVc0r4uxEDpL1ouF4lW
P4fC4W3XPzYR9a9IDo2HMbHebKtr1UjxN17f3F38yM9l8TapqY0lUeeZ9qKsRrF+7JyYWYtHAVNJ
dECrZ+Q0sVftH53zAU6NbGEy7DRM78SKc9bpSPCaEpCHIt15TaPGsS3ZWR1pJRYYOxWJzOTxl45y
XbCP6QNZ7JGTDQkim2rCICHPxY3zH6ZXVOpnJIxNXUqPF6TleTBoZV5ZOu5ugbT00UllCLfKDtF2
jII/U8sOU67Y4inlx7CWNHl1RqH8U83sR+VN++Ew+hEq02auOEeQ2eyhIggVidwwjR5C5q3svBrI
6MqyprVXvj8iT5mHGLP92lWDraQ80cPF7UUYcWomNGIXVdRbTnE2MxWOTJ8s90cHDbHNgkRhpUtz
8Dh6nyBmZIY+Gm6aF5cm1aiq85Sth4kgw2G035ywVBEkmNwSU7xe7btbUOZ2lakE2LJUVr8rOI63
bF+qsvxWUDfldZz8vn/5BoW5VKzrNEPUzhkYzCygDQLo+fqVNBRAkIoaABzDAY0c2rN7v3GK6yMC
tTSgyII7RtRJ6DXY8nTe2ScjUZ4CQZ5ohWz+ss90mhCE/nvjeafnO/9GTG51YG2S57FE3rjMez9s
s38he+nn5uClboxLsLtfQ+ZKLmmrweEeiQNG99l4XPYjJDkBr9fMQCCfc74KHu1E/KxwesvvD7yh
Pi4ga8MdwONsO73OUiz66kj+PjW/AzGR7XkgHE3i/+xZTXMz6MUmMTzHd/tfrrUsRaNH+JF2V78A
o21G8naST3mDDPK+9C/l+tuaW8pzUciUlx8fBvuRNcnAam9hCDd+ysn6SHYM8IAE6QEDuCENj2Av
7e4JDuv6jQHM+Xa+IgQRAVxGllzqSD3T8uxtCNGa/leb93xavW0EAlATeFAJlLbLfq+iZwGTg/4j
1tCN9cBkEqrcpBO2Tl3pd6yvwtl5deFpHauHi19SpSQ5kbBdrUIZBfwydXVctu1SnwPUbLEtbGhl
XNb2dJtc+OqOS+Hyf1aEDSYrF9fS8lSHLZrjsMHng4dNDlKJ6/3a3UnhG0COhGtZozqFdU8kqgBW
gbnpcsz2lTy9ZNWww7I8MAPeNC1IbBPQi+rRuA7URXDZUPwZQ83g+bVBsv7y/aOi+Iz9ebSsLI12
Y93AkHGul8LTGjJjF8t6K3ylRype79ydvdDyOtWDjsyaBkuv46tIgQPN9FCtYv/l+NH4tSBUTsb+
aOGfobUnXJo7AFsDn5/ogMacRZr57Blw8Y22S5cp6BovlOEnmtA76zdgUgvPRICYU9JoZVrK475c
nISO2lU8AEh2WLs2yyRTcPFip/KcxT69FWY39S+s4qksJ9LWjS66kQDV6KM8XC5AM+v9XQ6iu5qa
+inAFw1qtXST4p3Pc05O2pHCqsPPTWK58NwfDmfKDclS62RoBwM+XlwYNNk2Evr9jD99TsJOt5RY
6EYm7SSgukt4Yx7q5JK8k8ZeyG3XCeiHAEHc8PnZgRnjl7CA3tz0piTMeRJ3MzmZiK7YyVjF9zO3
rHdXqO6yLqXBxLHlxi6z5SYlsJRjdtFnKTZFP8ZXxF+3Cm21aL5ynb1Qy4eOdmzC+IRync2/hLJy
GHn/kwUoXUm8G6/RQfKDQVNeXEEl9wQVjreD42IuDuSk8R210L0YLmW34Ti/xivZtI7QydJ0yh+R
MN73egq1PPQqPgsePFPX/EBwQWjXsQzpTMM2Dh/VXpl/gL5ISDFttth7SdrLA+jN50vji3HKIoUW
3bn4eBSXlzbkIhuwZu54IGnOLsKa5Y4A9I6a6NMAxlxzvbJCFYxRfIAX3hPVMFhSF969GEpCMRuF
oFyAO2a3bic7bOfDDsMiN59BjQndlpIKgOlTM8gdoojHsGVeJ1shrv5jKCeYrtVcfaE0phDpnoC2
P1qDp1gpkF263cE2lN8x6OVIAAASyYz4tkbg4O09E8F6U/l1jQUg+ycuIh9HgNWUYE0q/acUKmdI
BUqPHlkyjLRBKhj1lnmSBAzamymIFh88bBfunJeoU4RudIa1w5cCjyTU6CeiSGVlnIj7JIkP/4yB
/ZprvmI3+Em2jjNw3lgiPouiK4dPk2LloHVesE/KwWerQJSa/SIQOJUFcQMRLcM3azok1OplbGXs
WCeZJYfCE1bocgURZ7IKU0DjQWO53q1Mx2h6kuOl72BtMpWBYgdLFYdg0bYyqnf+uBeQoLpi0as9
tWstAyH9ddCYReaLPKau+6aB7J2eiqjYjHjJMtc8k06+035Ird3dYmLO1SvG2bV19+UQf7P7GQtu
apW/BHFzYNXaN7/Sd+Ly6qKFMbLzIQOOaKTbwAV9fnAqXcnhV53TRvAZDKYp3Fji1GGJJB8txCI+
aSc4UiuFJMDcw/dgVRG8TPhNLS7nfiX+t4nzZujx92ingoI/VhaLT4vgd0+CfTIeMdnrjERDQzHW
Yabo59si4TiGR8tuU7SqaNpzcunri0dDs5XY439XuWVa57tLZIQhSevKZhqJ29XevZZ6oFkv5J62
b++U1KFYNaMLEBUVBQCOy3uFTVGbyXG1qP43LLasoDLPXfk1D8MSY13NamMcWsl5r183OTgms2wh
B0Mv1EYXv4Ycz6HLq2Up4BnCR3Fw15/ph9BlBolSrC8tdftxGVySa9nT6orLE2dm0IOloJiN+iRk
fKOHPAvxswPW2CVgu9MZtWdjvbYTM96QJ+41GLj+6ywCRcHYNyGTDt1qGtdTV5l+XPegdP9pNKaY
oUsD0s4C34hldyh485n2RnfEORRNYi8cvMsMiiVpxKNyaDhxbizKCQPj++svCEt3q4WcohX9c0Jj
VGvepn4VGedNcTFZaDp7JU39PyEu1MG3T3I0NZfBfYhsCm/KHk1ywpfJSwaPVaWpxjaQldeBgchl
Szo6rnfgkVOU3ItX5OY5Tl1tCysMJAiY+Cos2w9KIjPWTa9Q6TgC84d4W87NTRJfLUzp+PdmAKYb
EylRJylkOi3j84vB9UyXG+ISR5ntQiu05q6CBGuKFpQ6qbVSsOhfrXNorUCvJl5JbbR5FWn/74PH
tkHs87UyS5Oq36M2WNS0cr6zm49940XUi6IH6Yu5oCvo72QBC4AgqbHoVdHEc7Q51giEOrI8JCJ+
MqLOEiQAVm235RxOtB7enkhjqlZtjAs0FBmnjQ8BA/RhAap44nG443ynwEqq+U4yvHO/QdUT90Fs
Y42fkfaQbY2SOG4QBrooL8TEYy4kfgyC4INhAE1lgQL+egsz0C2LoVIi7THl18lWHCwOPDDWG4pQ
iE+67yU0kkwghdVfz98K5bvQ135ZIUvdVX7CfNoJil2BI7fl2OUWCfk94Vlzv7XGJEt1kg/SJ9mH
rCs9/Z9VO8kVRbQjOnWJ3eC0g53a9ZxThgvttsoGkNu79eo4Eg/duWgWRA+I9/pfPd5Dbd9gg1GH
XCe3uHYEEQiI+BcwEIdGkb1Ja4YnNbTKaqNb4aHxwmQDgaKboLMsqVAiALJ9mUOcmFqRIKl20NGW
/Oq13AFwZ1Um+olv4jKssur2koZAa/FhmqV/fcZN+mIKywQpE1yfZ8VSLukLk5vi0oeIeWz1XjBK
f9yTzj27JHOd09wgsz5sC3Iym7CmQTSgAYndJOBX/6fT4hO16dvGHkIv1PLsXAPEIB9cAp/VgLm/
kEaVerUP4r/eNMlClRWNNnMwj4EdhWFkTA4u6eTWRQ3ku5amPGtNSTm80hsFEEhAhFf4XyGboCmR
D18NdOubVHUmGhjiHjeb8MIIS5zwcc8g3MpMm0qS97GFIMDDDUcT1nfdNauI2z4CrK+N5nJrwJ+K
8HiyvjpZL26yzlH01fUYC1H+bVUGHt/g8aEU8zScffXt+hyn0MlM+plG4LttvhOrOrQWpXG/f8w2
kTKh9GgaHdJBBt2D+1G7mI8dlNQ6Vb+ZtKrlELytquhkH5e29fmr7cHQKC3SE6Kx6gL7q2TBnArj
FUDia/jEfIl42qEOYAZVCz0YY+0MPDWpc11rBN5Oo39OGCMD3tf3fu+Z/g5tZUXRuw1QUN2bwfR5
EXQeTOb5FF4/OuVuOLZseAL6EOBQfQOHVPKbVWr3jaNQIBH+JO6KDKaSqkF5aI6h6XAEwh8hT//6
VEWc6zX0Ci0+Zl1ClSIgaqDWq7WCG+6SLaAIo8o1jgFP6tWYGN8gODrtvBxwwj3EpCSkpzOmkbOG
wurrxYAP29zNKfhgNCSOawqFdA3Cr50cwXO/Xx+65+ixGKNrx4dmDXw0DijdXg5OTfAdMVEmZYjF
aDOzKbW7JVXguPBYiJM5jEwSVRYaP/QdJ1hUmbxA1dp6LCJTx30649vXMKBfboFDhxllSUdQOeE0
PpsBD19/S1YLGDgvCflyNRMOiVUjlKa91BgwPp02BaITrxbiZKKroEOrWrHR8IjhbR7jTVjh+ncI
o24Qvl0XxKcsNekvEQfj1NZooaU3PsVGxBA8PxX/TTh3qzJ4Z75ZBnYsrYv1qP/3tRDb40ZULj0v
Z7VE5jK19EojjJh1CmHQCG9yY+hjEoniuKJkUzbRrgKhZrNyjpoIAnX11lxbJb8httu8juFMkM4H
BQ7sgBNewhpj8FRB4gTJneDiKo2vtUIgZm89yXwYu+mVyqT2AXS46boWT1WNqfONQkfFJZVsIsvc
LCHNyI2yeVfW7qW5rQW9mIRr1tFDQpn0KsyiyAsGWEsoRf9+tH11jCtn+H0zwCYhLPEZIU8nxi1L
yAdC9eFF8puGl4AKwUHNHU2bt+68wc7FxrfA4csXe0Ja26oJTVuiwuWkO9/lp+fyEW24wIfeDUtg
1VdXYFa0KBXg8syaXyHQjkihxNNxu8628BN7oJ4XrGuLo2XMQaZ9EYibwbtldxg++wuviC8mEy3w
QnPMH3I3Kzf0dDBMWkrl0q9sFgta0Es/63KEabWzHBF7bPRxdJ/OjEoo2X+Vn2ReplA2OQjbpMFB
LFpLhKqo9xbKyltpwKwWSRIJfVMR6zK+XvgPYpzvzZzGNwZmZL0fKxAgpZUMZ3jXCrPXqRl7gCf4
leIBDOjl1dz317+7qDMFCbszTMuoeUcGc8caVNvovkts559i1B0L9yCOx9+xpdxNU7290mwMg5ji
K2xsrRXqOxIYoUi8KUS9mhmcI3Ft9MOmfgE40lVjTJMOmL70UlU13iexfDsjKNTnwh103U2Fv0lv
Fr6tStPsSyeNiBUXMBBT1wdZTQ2brszlRQuEpiAucbwVjEsIdVAjdDm5saqNg7tgmx2oWv6bPASq
tQ7EWiNGiX9DyVKs0iVkkRK4y1NDaQZIBUozyod/1HWeSmYKN7/uPL68tQCyAECy3YvkdQmlUNmq
9IdgMGWQnz8irAE3kC5N4znGwp2RIUbO07Bgk1UyWnPXfGxtOkZtW3dAj0X1rrnzd3MvXSZNwS+o
NBgA+7qFwbXd2LQ/6fq7Hh2srm8fNrxccpx5/2R9hPy4ZQXr1bcc63UfLFbr2I/l6yb5o1L3VPP4
HqT9SPrIfNxTSyFBUCkja8dTajeH4Q+aqgPRcM77X69jVwhG45V7r+0zCW54y+LatC4BByU9K2up
vzFfkQbzYlx/Ic6RzL1aEw6KwLaJd81NncI5TVFrmH0Rs+8f//1aB2gNKqtQK5kcJtHdtyJKyw3O
7J0b0NTaUlp0aVzMwA8EumkV8aeM3I3WwJsPAbWP2CWZp2Sq8dPwcKW+9Rx9AXERaIIjpzWxbL6I
4W3c5oDYt58RQe6H/wpAo6Y/kDUjnnVYnHByLkxlm8I3+KtykkA5N+WmHTfGGK/7qS3aQsGt6BGh
sshaZgybUh+5Tjfk6xKq8dRDPO1MyFv1G2lIE2W0JEmJJr+MxP0vuwiJ4dh7anQsvPUaQD7A80dk
fdh9XJLGBeD8/rC03HASCIhZuV/a0VHA8j6NJ12EvFXqV32NMHBP+Drts0dA5bGCNSDHEyI8h0Mv
KyFLrijpoZvrd6zZ0+YSqs7yWswghQKfTS2CyZ1i03wjHuWMYksJzCCsUrliM0vT8cfJO8dwXQb7
MSmgZmgjYgyAKMlM8jT7Xv1gkD+BcW2oECm1jFsZTf/6O0NP6o2NAqPAbRzS6J6mjz6u4f2t8eoE
yedSoCSjpjRQyji/oNTn/7CccoOtR7iVVImykEXkzBbK9No//tD++L4UwtcylyhW/iUIPJnCJT6t
F9XpkvxX61kUnXrA4b8clrgfKCaexWNyym1ymdI7IKPZQzweKt70V42b7RJrUN8+PUaLl4JeijQv
cLGZVRgJgRQdQHVtJMpg1kju9phBJlUbPiRUb93R56iyDJaMnw2d0IPMOzES51IWO7NfhJR+KB6h
SUZdTHt9xXtzLSTzqYehJjBrsW41/9j22uKKpaoxGWjdz1qbFS7BlNu7M9bg3OfH2Y3xGh16mfce
hv8qJaSWeN1dZTBVsNbmXrLr54UtPyWXyZ3XkA7vFARxeT6DsGzkmrIdasFwQb+c0leYeh8J9oc5
NUlm5xmZYoKH5oB8ikJa9RK85JwrOgGh6k8mKLYxIXEkq9NGC3ljteRUDV/Ht3K9oBe9KxnJXogF
GAlYK9himxDRDsQ+09G0sTjKS114TZdFFn69GeQ/BVfXr9sSWt1WbGkzVmkTctS1BPAIMSu7pSuV
Ffx45W0J1ydUKQeYPOX9aYh4TbkdVPPGtLmURS4LEaVRGOBNR4aTG45yCXAa01Wg6D8vAVBY56sQ
zbc+FWy9Z9lVfPLFfPlX2392Af6Q2vd4KKWZJGS2fNE1sQc1P98FuHovc7J7RMcGBxeUammHi8yt
s+sA3Phodl5Wff89UNeS/Qqas3TUuwEolqSJNmSODGpxZlkwMcDpn4tm8aqPaXAe+2KIFr05vQjK
43Zag8GPSfOyTooZXjF/T31dFxnw4LTNr/0LWfvJQ1UHfKgAAK9PGdHtM5icCtjKOR1s0eTmxecJ
+s7AontyHupCfc9D+jmiCt1oQbVwCM+hRSA+skLB0w4kIb8YnVerzAtuvV28WcdCsinpYIlNJ1zj
kH1X33TVAvb9j03R+HNCRMFtuikhELx1Chl+TEkKI+NMVQo4RHg4W8/Avs7TWyLv8SI0WvMdxFgC
n9MkcXVddnTZ7Zkudcuf+qDJBK+apqSpRyvD6/WpsYxRH0ydxhw7dWnGj2BSKKfgVPgFoy5g3Qnu
XArs3IaCM578+Xx4pHPFw58RHFutFe2dpoqsQTqCfWHea0+6EQ9SpEODH2W57Q9arLDY9mBdCSZ1
obSMLgZRJSv0xGaKKLi/U2wCbT5fMR6V0Uurcj2U6TkTlG7O9yO7eTxDmujwsair+iiyr3eqHJ9r
ZLRAb1CvuIhTuiYapm8sg8oqwmwBWxWS8EkzXrUBuq244MY7kzygHeh8+lgB5/iQsOuoq+knb4mG
MlYtkyAFamhaYfjgJsW68fTbdcAEcsWJ6p42BUFOJfKKxcedA2dYB5r32tNYJjXVlhN4utmim3ym
S+FDgDhSZfgl1RoAdXYWiQxh05H2LUy2psC9BaZgKJwpGVkBAWPkBXOZ7Dx9KO+8VhCmsrhsfxUn
Kh1wBnC2VwzeE9n5Wsp5hpwiekkZDFlNudQ3NORs3FSi4tvfyD+g4wc+QKsfk30SXa7Se4nMfCjF
KdzoZNYW7uXpKeD7aTTshd7gR9IFlI/mjJKnmJ81VgS1Xwmeud1qrJ4HsNOgw8wXDHLQ/csZEh7+
5DaGaCRjDl/XSqjrldNfDRV1/LmnEU1ym/UWYPqBw1RjTOwDE9wBcTIVYfXk7Vi2JDbauz7dX6mQ
zzn84J3Y129y2fo8zAu+mxbP8Pgin2TuXyDrKFLPoSGr0aVBGfEjWB34GNeULSRdwJSXfJ+SrIF4
9JksBVwBDOthIySrOdPIRRAlDZOYn+i/GbcS3GRQDE0VJL3N5Ey1rx2y/ezD/Ys8INumFlxnFfaK
kzCD6eibxpfFk2Sk9UPYbw9M6cTSp5UgQ1hikRA4FIfEu45ywnmlVLbdsMk+q/2gGrX9MapH7dPe
A51X1opG2DSJ9cVDSpPSk6ljDi/YYWIuzhiCfzwuyNGav/eCECg+JkznRx6U/Tz3Kobg93AIWc06
SP7xAUXklL9p+vZ42NEkPykt3ZMh/My8JKilCQ3oD5aRWdIaWThPLi1eMojcx7uVsU+WkBNhg+4l
azO2uSYfqeb0v7d8FQRiBZQsQKknQJc09LRy0jARlC2soUjr9HQC20cuYzYp7O5tt+LlgFwd2qCn
4O0c6rpyGsWn2dqGX8IOCsXC7pdTljZHfKkz7VpN9Rez2Yv3Sh13wD3CDR4lNWOcAxzcrIvNk8nC
NVFc7BuCsPnvn7rbHuc/YrdA9DxAoHRTgL89y+fH5laNHBYNFqwPw5mpMCT7U9TqclDyZo8wwd6H
BBc87RCM2jJlcjYyo5Nz1uut8JuH4h9BN5QA4LgknnVIaDjbQmzZQ38NxvOIzAu0s2eqOii8Ii2m
WtynTjzN4G0HITzyX6YoyKr2Ind0Kh5IP7XhEjMz2qKiaw4UB3eNcGs72exLHXQ630lMMyCI0qCk
6GOEVZC1PIzDjjsZwPsPcj07NaBHfbKgnfEqX48tTt0kKnYJhoBvAe0YmmqZZg6hbT3JWDd+MfBe
m6Ueb0zJ5fuS1Ul2TN3GXUPAlSDZhQS04FEML3gVtJmCLHyERrI3UIAm7C3UjsrZEEXU97Kv09r0
haLJklfrULUmMI3rVv7eNHDJUUuq3yhis6XL5ZARfLD33G1ikL3vqlJRyTs8Ky4j1OEQUFkRwJMc
Hx0w7nuqushzSYgZbOHG4mbTCCy4Li1CgCcqKHc/uYGM+93t8oBuW+SQitn41QZQ750modNv71rA
vY26h+eioUIIxZjJ6vM3Li28tSg9Tq17YVO5iMJCTHtYdnqD8pZJmUfWgEcME4XLIuhn2xLz1vA8
nqzQXnMRZWkMiDL5CVgQlX8lkLj2rffztnMmLiN1A/kEYvIaZettJJsDEEwhLv4ZBH4TukqCwHwE
5n0j6XsTHZ/2S1Wh8Q9amLWmZKbZ24lmHG2M9xmbdnwXz20hPsqWCQM10yURXhvwPz7gPLFZRxzS
mVlSd9pTWYRgzV/jxqUTMNDFIE8Vm1J16jgjKizLwrtBmpv5s7uXYrEWgob+5+QuY4GMqMIDufdH
QHswpS6geVcSstxvMDEY9Lse5242GKuobBOlrZymGH3UYYua+kRu25VP+AflIaFdGKqfKCwKapgS
DOOsYcWvM098Sl8EuyjQBiKFGu81J4/A8+tsdca06vopzbksqOGX4WwgZBeOqF0ETjQWM9UqpI8Q
x2EZlOBPGfytIo3HyhADBuGTORPeE5ci79mDfYtR7YRDRDSqgZnSFUwc50tcDL+hE1GxcX8rFJOD
L6qAgiaBCV+gWGfG+Z6uTD5Cb97WH4/Ck0rncEZOnENHmzK3zT+TBh3EKHzXGqQnqN5IPf7EZVE8
CZFTlDjU87t2+EhYFCxQG9yJFs5xjrXXkh6nrhrbTiwtpl36yZk0SQswFkgkevYnEoWDrSJaZ275
Eag3fWEzKKooN03wq9WTHtHD6ZXj6cgscXPU/QPjunnBpiAE/AzpWVI2V6tq6ZULAefJZJaFhFYJ
OUlT3tBCbxxxEyqfo8WroM749mGsvPMvujbon9AbYq/KD2MZ5mFcX23aZcWWw4kka5RmPNOvEaej
NyRfRPpjWR/QovmhdCY7mBmBjJdKVuPu4aGNT0mnve1eBUdhbtERP2eeCNwMdwWMFyMr1xUUnIQu
lvehKDskYkJjGqPbp2zhHKQhFgNAbZLT6iAUrQ2lWCnnsliXzMV4Fncz1e8bU2cBNkgzOoV73UpB
jifkP6vYASnYENr7AW0rlaN0EuLb/oiODTu/0jbG8aNKZMgVNdYiyGVr6Ruro9GDiL5oBKDOgRDk
dhGLf5pDrE8i9O8C2B6WHLn46hP2W1pt+UpC9PlmKJ1IiSDMxoSHsPWzrLfFf7RXDKFi18ZMbfN8
EPZAv3z3AveruUdS2/AhgbZqNVeNS/Dq6kSWxLLmquxBO1h1mIfWp+gfgmE1fEh7z/qhRRcHL5Qj
rdUx8pzOwDLRZuPFpmD6zuVD+OZevM1d1B1luZUOyLpOL9wKrW97ZnE2j02fc5JSX02XHNmbt/V1
ktvIBSGQJjW8xMPSmG7qb1LwXPamf0nkdSnNhkQoKVLEMZ1LaZGaQmJXZ+Uqqj0WcPz25BT/yBL1
T+6uaZIkwT2yMukRi3oUl3U7r7YcM5RdNgOSQh3Ar+wbtbqB99AtTdlOsSN4N6a5rzOKD1+AaXmK
qzWCL00RXC4KL9BhQI/MU5TXUSdfTeh4hsIShR5Y+U9lI4n2JjzuO9AdNadbv73eEw2hl7VzAx1n
QgUyuh8wf2xsjVKdLjgoWiSfMCXrsAd/k/p77AO56Hds+GFFLBzQo86kaJtN7sMPqaPsqabKieLD
b2v0Ua1QWTki2zssRTwFEssSA7XUVZY/vrKlLP/t1jifSPqJ/KqySC8H8cQXxTqVPSEL9KKxvSY7
0rziOoO1+ZMTFyh05L7r5shHAhQubcbIWM1jQB0VqUCgB0t2iTP8IV/FEezyDQ+7Xqo4Tu6IDfWF
dX71wc1EqWCkA0LpVBmQqzO5ZItnAveFV8a9+mdabLFs3XwUJbMLAkrWEJSoHMbZNTmiT4ArWGrk
PPazXVxg+FVvvAR2RzjzjHkhGV2vy/XvPH55bhE2+uUeaF+mPUst8SjwNy3B3ncI/LmMOUAuRWiU
er6oUWwCn0tnjBpdZWApugl2aIHUcRf5rqL0HnbgSaw8yHK64Y5JEnxYIN1OJicjipgMqgpYgorw
i1Or8JfDf0a1ouiyO9JlbejFAMP1ibXJAYLJBfnKx8bxXAeEVquBVNZI8Tr/3ATyMKOptBEB7kTg
H+Us1PrLup7EzP4mwmQvc5Hmp7Xe7hmLrHrRT+gU/L7ZEV6UCrsyh6hFjuL1+sbW8RldbkY/jwqA
5dAe5CO5qjPuwpdq3BYmFM6i7ZX7wFCqgl2KSTwmlOYQOpmWCu9xR1IDUNny3ZAwdBp5LVhcyJKi
j6/lUXJW94GkBX7LUOsddzF4jkrrU+t3E/b/bgR1Otj1clBetW1rkauveoh6+16i3Vst9o4ohOO3
d2H5+AQb15sMnGdGACOdBKlSiXpuaoJIILTqtkfudc+EaCzk9jPKR13qQBX05XQlnEn+ZtOB1yKR
mCxHjkEoODLBCThnIDDOwGWuKIiiOBS7NNhdymzD79MFd6H6vOWv70P8hD6V3RAck7VIztSd3IGh
LPsgW6pivypFgvAOIbcS/VyM+xfNfzFCQcoSbJNMSEt1dMNVZRmPWoEMD99cNqLOzW5CZbm7heOn
/zR2dqBCeulJsf32WVTkildues4a8qFVhkU7Hagqxt9aXbtfBsY5v9n7LLgDmoM9YF8xtcSsMMFt
dA76B3b7v2F27viixOwl+7EWs3eiqyIDrOTFWrkFD8w/u8konkKbgHF+dOQY1VbkFdFzTEZbe1GE
VAr1oa0I9GiD4Y7HGUe/M6DFIrtk2Rev03O1iGSh7QYoOalBF/jh5OtCD5i9IQQC3PQ3ZS5ctY9T
zFto97pFfnRVL6XSrKGjU+bcbT3RMNe7V1dfp3VbaNcqyuKEdZm6zCNFOFh0VcHGAA8xT5E83U4u
ZlxgBYi3ToMlZrXt6h08NLg0O908XrYBDOi7se+CxlfzntSg3JJjR34OFlKROOr64izjyATpOt4i
5KLJKcjaPvseQhhV9InJ0hNZtUo1XKHbORl2B4raWTMb5/YvVLxCWS+kSXXLYSEHHuwcYFIZxKTb
Ot8ar65UHqdmT9/E8cII2WjzszcOW13DXOW7s0vl8lP3PmnG3LPRHwbCOLZJRzptPuA87PI/A42b
ssh0qIPnfW7c43YJizyz13c4a/TNggTKie5TmZFKlHTTnw+p84XUQo7Gupe6baZYuuSCsIW167HO
ZKbz/ZWIneXpqPxdL7+a3sZI+Vnk1b9DUot3PYSXcfAB05uDhj2G6IragxggHsyTo2BIQfoOVGTa
Er2hGY3Soddc1K/L2Dl+SsXucBxFhj+55KnXgNgQewsJSg3UL/8GOEbcbhAy7as3X9tDQ7YCYu2X
l+mzVoaf9tB2cSegJS1bx+9jfN0MJK0cdodSswcx9EQ+ntweEIVnJg+t1zLBrKuV5sG3TXSsSkwm
6Tw29YWSqCYwdZQmp5IgKCmUm19DlDH65+f6YxcDxaLeFhEgWCkl4sZGPQCO+16WTBpt0Ff4Rxmw
ffCz2SDLEf2nUMhxdz2Pl5Jsb9K+JAE7ksZRA+ktibc6wuu3Fzw4Kay/Z7SE3NrOJZEY4EZKFbfy
TNW3MtG6zagRtAMAZauz/OjpbJiCSMyQtJQRuIdenmhDdQTwu8cGlUtQzUMaugEDXmD+WkaUBRv+
ezH5YnDp8GMgXASAO1ck4l3k+kytU8lIEenrZjkOhnFJqHSe8TY3RY8utJHNmCtf53T19BT+4rsi
NESfJsJoRDzIn6TjQuJlEi462i3+Zg7sVPB+LzhReN+HRE2W0VApj2gwPXd5tjqpyXXgnck9aXNR
MZ1EEOzmYAVrJJkA4xjKKcNxi2HSmdpovsmL2ldazXk9PwvrWmb1EMT9Yjs6q4P0yeCKHAb1AQV7
brSLK7aVEZ8IEnA65MzNYyATm5Htjl5544yV9Xz+UA3Zlf0diiGHz4yDGJF/9XQzvyzixdkhzdVD
XVzZqCyLFVXEL+A+NG8sU+AAoeKch70bzXdThaxq8HNMUE4f/4LOl8tV6Ptv54AkI36uLmNijn/z
0sCGTB7xmkOhhFRDfWW9sUhVgIi+oRsCUCZxopJmeeiK067ZCp79XSHPdvL8DoN1/N0wo10dtJ7Q
aZtLkxoO/srvbnet05puFc2gG38gINYAym5ffHPMd/e4qYKDjCWkQcXqpjzPbnbZlZ5KIug2kg8A
QH+cpggk4QyCfjXyFpzo6sohrYKJJPlBS7C+HcsWNoz6BSPFhKMIP9tILYsU5sbcCjPuB2fGdqcR
mVYdGbyXgnyN9ZKjZu3qQLUqbq9NrQ0JNPOCB8Bf95zQYnTJoRiKiSJQb9F9Qs0A2MbCTAxF2/RK
H4MUDD/LOnW/y5h8dm0nBOnhR81BQp7vwIGnAuFn2CQDKo1Bekv1+3U2U6B1b3EiRy2moTwSP6/Z
eB/lAAmURrTGjYkGpdHXFxPGzOqcRHoRQ80ruB0r0RunE/LqWrFQA1sUKnYhpBpa17FDlqgN3HMe
vBCPk4bKQhX0E5VHo9TB6VeOLAtwbPQeFHlIZfWzhe2SMOMiqktZW7NxQsvwlDRa0aL+jf2EaVJ4
ntLfcqlau52CJjBYJnzSWVwxMqZ/KH1kR0yMLQbg/IF9iiVzHjiUBKaKD9HEJZl+uyYft2dKA4iw
sKkfSjcLlWnQd2CZ5FYAYcrKvaExaAh5KR+t9TdWifWxnsb6P96qC9yLwIqCmwaVwHGOUqMbtpHH
bM+QUaxWcQyLyLWS2qBQaGMho5Uw7KccjVPIqAfPa4WkrLtVhqzurnHR9PKWjnjOHI+LWfeWJJe6
yyCCTHRG5/fiy2RtrcVjnNfAWcyioMKoFVQKjmBzyAuz+RbE0RIvYUbNcH7WfXsplzoC10fNBx2E
E8KN//6fmHRIzCs9wyURcFirCZKzdOQnNah0EFNLGaXuMcs7V/5mL0wmBVeK04IlVD0q3lATupGX
voWbag7zuarvDKqkfsonrM/tsdHM4hEv1HR89+SYLVdVRk0wROOrKKW5Wtp9uydQb+SLyxsyxrF/
Tj2IuRRBg7W3rOsn03QABGtagXn5DtDCb2heaFgyMwyek6bcWS5C/E5Jw3XHV12s8BgG2+TDUg2p
TTn239W3Ogn6VOhOF8VWarLRSk0C8+PkdUqEHsTSBjT4JpPRD3vTnLqQnyzRm307ZhJBPfy2XsKF
vxLPfscHM6GeGB8nmnMt6ssQmBD7gTatu2vmAYg0tA7OtThCB5Gn2jyQqcSqejP8Y/lR3/W2nElO
lX2A8m/4+O7tMwmMlqolHls5S89Fl207eHbT/xcPZZKn4v5jkXdQTZ5vwH38u/XWeTzxBTp9306k
Nbagygv1R4whIp8dCTKX356z9Rzde7vySd+t9Tg9kfAmNoYqAb54nauADtiIkezHKsYpbamqz3F8
wJKGZaupapKtA013fvpMtMNnr8EgOekVEyNk+kJmR5GBPDm+/xq1uzVsGasAxgdrrYWmRHnPyXlD
ba6PDBUhKh5mP/mWmiqozPnRMrZ4UocaZJVrOcV+QJ+DXFZaAUhI4p0s9+kz9GSGalA+FBo71H6U
NBHnU+3S89zIpcg7UsmU+B6zPyE+3uGiFiq8hi39HSsdurjl/cLgR074AQatFZSQWgwgNuIZuB0z
U/WCOY+ebiaZvpzO8vbVvTqvUZFDkoNcW/nsv44eVokBNmJ0oZyIe95AGZE6bmZTuryeWiRZzg9O
cPqSnj6SWKX12PsSI5Atrt1avgnl7t7/mYGL9IJiJfQ2w4xc2NkWCBj/txSasP/IaGpWIvdIbz52
tUPlg+mPjdQUvxPrl/V6dQXSn6tm8hLzOFFzquC8Zha+9SGPyJHdGjFzV+QLQ96wimRrpLqsPAzx
y6DvWrBRWBAZExrKahPl5yMqQIvw+lk3yZDeVho1Npv0vF2ZKeAaFJdg/BSLFvg2/tlgRgEmrTKy
hwj4J9py4TJNPTqLPY5IDi6AJIBo4idVHooBcoEkneKsBlPQk+Q8HI1wQOG59m+J/TaW/BUcFajK
aZBXw8DLOXldb4NdeQogNsfKR3aAePiG/s8jSeyovWnwuEm/7wWPVNo/9B0bITGGEDcu/EdoCZ6S
lWdHdgE1o4WktMyNlSVolJSbdFLVceOtjwUkHL0YZNFOu1xTVPn799tHXt21HCLsodso5ufegVEY
tVIamLIGBIwq8jWZGpFkotdUNSyczKv/9VjMqP6yb3POlLH29Y+Cpjh7xddHLyIJvJwG5wxSW0Tt
Pc+1Eh6NpUVgxXUDYnTsGn2VJoGu0YDeAQuRxqXmtFe8W3Oy0E6Tsgu4Qk9pm1z6gyJCAOUoO2AO
5tsVFryj5C+euybmZbIqJl7F89F7h3GdQtrVPrO1UddaANvx8MMLZ8VnGPBYZbHsaqCZrMsWr3PT
QllkxFBq2V4aGZSSRm8S+OhY8lpxJupe5JisA2GB90Bogzc3OuBa/N1aXEP5vpCqPmdgva+Ki8Ru
ibSvzMpRcUhMfjZ9JRn5xw6i6YbDLeGOw0GhrACsW/1pQ08Pqni1k2Erx9Mb1gGsxxIkrNMo3sH1
5OoT1z3c4KcIWYZLhvAQpnQDiivOidWathm7Qef6I+w1K7mWJ/H6DBgoAE+Wyz1BkIHF3+neX4Ry
WIYtjBvzyLNEOkiZ4CoYcPycv7f5jVLxFX+UHu5db6IIzQ87St7FM7HfCb78VLvIJv3FZmSJzJdo
I4T27binj9laQ1SJ35dth0M17H7fWYdTeKTqVeOD4jiChaQfelMciyA/Tbv/VBFKv1cG1YkFWJ3V
9T8Coczue+/Q3LcbGARUl4P688kgq6wdxQULi0ARzm4mg6yqN8ox4pJ12O61WiFQK8J/dOhot5ci
1kgPiqWV9t9j2GDZPbBAueh+qBxQgcY+y3J6AUAqJcRYw1h5cBEA/BRm5rnin6QATsnlgdPM+PNN
fL/Z/QWBP74C2SrF/1SiP8GjAbM7jg7Y2/i0JcMRB4E8rmHNNCu7aBoFlI5FATY9XQ6RX6woDsRd
UuXSmVmNo67QBNEIfwA8caBe+albuFp25nJFI/Eol+QoTRoBfPtAYy+JTHtp73GRDMD9AUcoUpaQ
NNQCrCK+lAG+ydhd+9wZD5zwh/WG5KIyV2S6yA08Vy5V5FBi8F8yfb2RbsUh+8OvxlTi9CF+KKK0
mhNMZZvvVkuvyPJqgLFme3hrH7G95HXAXIXWy+RkH3E5YkYfbo5+kYQPHH+lebfvsJwZY6KZiS4y
CeTGbWkgX2RDebBiO+0wAzhEy8VODCJh1zW3SJDQwb7DHCIyNqLSAwo0UrPU5wJKLcsvneCGp+1o
zkbW0YQXpsen4XnqhtPVzuNb7GRx6CWNhjSkQ44soB0mQLvw37Yv0j2gR7EJaqFimiY1a9YTeNGR
vUI/qKGZ4igPQRrSKWSTNjESr6hB/Rz1Xkye9fhJixqEQAPUvFqLjuCHHmGGOJmkqxw5RtcMTi/G
qEUbdCnHlASz71sfp2ZLXp2fnWMZIv/DGbHX+EQMyUqfyMMgaMb4oyVJGewLoUZo39rch3Ojnrda
hNl/T+gRjmN7Od64DrDFEImbBTNuu4I67YFkB+Vu1f7+TngCa9kqtMeUMk0hB8ddOWh9K6nBoS4C
V6Cg1AMikkhcsRPbqm+RsFspWHdUipdb/MOPPhglwVW/rRLhW0CCXInHWzQpTDz3BSZOux1J+cDY
iWqpEJN9noi3OD5zxKC4dDHGrm2cssSI/RUTTMVdVxJwjNQy71ayz20lgQ68iGT2dQCrOlFsKMRd
GurEwxnlFqio2YxSwtQEhl77LAVQ1mVl4LaP8XCKPnRKoAg/VbFwUXCC900nqvJpsUFp7bv7KiPF
lvXXcVLfb3g/OXlk84v7XeuFM23zW2R0eL2/LylFe46r3uBraswnhFfqqkXGPsrG+Ecc8X3HQXJJ
gJLtYAuWk+NucLFKGhcFDuQ98TOovD44qlPWETngxBAJIctUCJfvcIjCTOu8YXhIuKEshvC8KoIF
yJDnHQ22CTOQ/niP1+/wLPem1+eixPEHwrFclvQYLb7rOVw+U1E1iB7NE3H5TAK3Bj/65so7Uu0y
Tk5wId9v57Wig6J9AphR1XsAbxmJeXERXFAnSj2jIgsmLVjzBWDVGngKewSYrET6ctZYqWPK+4Oe
iCKVE6LfHEPu4OjKMgdZ8c4w8lL3dg6kgEv/nHPvlcsPLa19HXkhCafw6DdTay6eSB69GjRKBC+z
YPH7SEmuGCsuWX9qZR8V/PFBQhwfroLelkU+u8mm3dACqfMe6+tZkdNCkxOKKlG1bllIy0BB6XIa
7T0krsxh+cOY6wpgj96kH5TxCxXipHQajLBl/Kd1H+0yvG+lCrBUJTLm3ew1DE08brzCRuVL39tK
eSfyQYbqRzk9Q6RC1Et1asO9GcejzGfqfoZ7EipqA8zPEHJgckzYvgds5Wk3G1M62I+DRMClZber
d1Jqxg1P1YVw8sKf1l3ZR4gN0KwpESnd/DPNS3DnJA7+IMjMKM3OsO109neGnEQcaS0HR/OFCLgb
NyJ6SDMLy9gXLBVx536fBFIHUAnQuhQQ552ziG0u6JOwxHdqYH030JTXYtiR3snlbwrBVSyPPvLo
mo5Rse2Q13gLef5U+f7OeZmhpr4z/Lx1F3FX8KMA82nxe4q9ksVS5cJHi55lbFlXQCD/p0jG/QoD
NSPUtsEeJO7NWcAG1jPYUTLaE1MWXeRs8oid9yZLgXQkmrWtTiEA6WWRw8DnKd38pCtmjRXCZyrC
f6PpoF1PRWNaFsAHH2XrpZCkqQuGb60u8IDL6wfJTl1sW2vLlgGDFw1aj4ppyBj5m2wFOhCFDfCZ
itFU4FS++Qk1KMewWFxe9JcbaRWDL/Zm/Lv5KLqEPfYjgBjE2TqsbVgrWol+UXM11RLRBDQblC/f
iVELuUyUx5MqkYHfkxddY16l9stnJgZSfZJ3ACRtqHtIu5kM9naLlZz/YRL2euMV986BeRCIzMTY
5tevs373Y9I+6qIoMpnkg/fhxCL2YUYhCnEZ0rPJCGmxdYD4yr+y4IoqnZDuvq5zTs7Q8EMi462o
3/GTT61BHZ8c/VLfD4CFWlev/nn7WMjL5oaN1Uh1VjvXRTZFvkdTbQuAOHAMnVmZUKUcARSzfRd1
7WQFDDGDn9kLdER7tqEP8R0OtXdgfgoOzYnppTb7oCRRx8ybfat6iLxLl1tkLOf0xnJcL6DXkG8B
A+WiThJCFUlWHY9s/QMPNwxnSEqaZptqHYTK0gI5hD5337dVt55DZGe2lv8pmtVKN0WhV7+0fNJA
hxgNg5pqQfrgWq9SviAvYoB8cTPTwhyH8J9vifMH5/wlt09krkilOCo3yN5oE48kA70Qr3XwXQtr
TcaMNgoU7Q9pQtmHZUXFrw2o0EAeWRH1ftVPxAK7zps4sR9bTeiUbaFheyzzKNab2yRSKaJ1PDWe
SsyteJBAE/NXHorq4ngXDfpVszPU8GvnnZnLvo2X8q3NGX3UT2+xd5JmM0lAtOHsHGtYiuu1ozMv
m1fUviEo2V6KJphHB8zz4jq6SGjiuE/D7I/v82cS3f1rCe3JvSmKzvtyT0abqo9NA+xQhItlnnAE
c0rpluqs14+FUz+zSvXnR1DSj4XjY+xdw7npJ6Q6p0n+LiuFPLG3TTS1koUV1iOrn/eufw+vXtVJ
0VcXrK/Kd49+zEMbNMDvMwyIHDiOJe9v+FuYxBpW4KA8dsUP2xllL4ya6EBqpPzqYq0HlGE5ILoU
wASNLcbElJGRT/lSdy/Z9zecCxWwUDf8JVzJusujUN8VZ1Si0qujIPr6Jz8fRFB4PwGFqv+reUEX
p5Y2E9SkpFLWRAY7lKCTbSQfLwuTbwaH9V+n18QhKz1ZdOM6JIS7EFKdyWaT5NIgGDWDol8Sf6c0
CyA7jvYdRMhKwr4f4lNJKcLodK9Z7uSoZiTZwVZoNtEYh0Sh5Zy1uQyS1qK6UWkhJ+FXZ89GlC+2
fDHGy4VcZW4RXyxYPuFBuWa8qY8dqp7SMIPIelOidiidb3/8854CuzOqktWsL+h1AqMZsTGENJ0g
B3fff7VcF4U5YwkYocyHS3u8329xuoG48qhVN5mXMLrSu3Xd+6GN5+9bm99FUYpLlerP/1DP/0G6
o5Wvm6GhB+PtW8y8lKb07g4v06HlzFAqbL3VUubo2nS8vBjPwbxFErQH2UdNgZP/fujsW9M0WDZ0
uRt/ufKCwQQ9ObbTNfClUiA3QvV0dt+waNqXi55JNgJZRLu1KWer5Cc9XBR/JktvZTFXvDZ3Cxvk
c4Lv10XxciwTWqVTyaZegkmXwfAX+wSJSlR90TgpBsQm/hrykWMsAoQkdeMyf9u8S+4+eIAe3lqP
HnoixKx/e8OpW//PUr4yfwHJBxtaItc+051G2JWZyNtef/d3ttgtadV5P5+C8Izm6VRNzJs+ZGBx
uT52AZuFVyS2DX20pJgzF5Hok/064RXsz3vmCqi3D8wotXA0PyNOg7uU15yalM8AZ+HChKpoZUHS
dLRLovGo1H09dptbm6EmdJwvTNwamXwvnByoM8PFsTbtczYe3iMHyIGY/2oNWNbkWyFNCW49z9g7
iPDiH/cky8njrWAkcD75zeBiqldeqdiEds0GXJOz7IekuEGxnezXvdemNkfFm606cVSIYNeYvBMw
2274VD2EQN+mBPzi6RHbqLlAoX86y+GxlcOIZhOdSF21ZfX4hXlgpvNm3Ac7RI+NylUMcbV09LAV
F0C4GGUv6dPXyj3zSZgqJZH9cZGg3VYg+mlhDIScYgdREbCrGBvNNwpqBnxxt8ZqXERkazAc4Vhs
Q3PZtdpdpJiXDcT4RIY3gBOgUQOGYY4DBnsHnHr4/e62vxKVRMGQC2/4OPlLIPB9wsdkeeAAcYwN
uylOQ9aZ49VUFeCNpEc0MNXErMHM/Ag2vogCT4P+fM4QjnyZ+PIQpo83Y1cF3qy3ZfefKrp1nOk4
cvEWBpRfkhnWtWBKQ8UNrB3ImQ4ueXAWdgK9kruSXHrfMtiUP9Pmje1xNs9IkSxNWsGFvuwvkABp
WaZnoLdvmsI7jZFgg5MZR8j0cNrmkJQazbbQLT/psso3aav/6QnRZE6eahr9V266WSFfhBPc3cYj
ZTQHGX0nwtHuaXkkgYJlgXRamcup9aUmi8GZpdGXowXQzg2c/0bzRHTcx/zCyvfsqghYgUeL0uXL
lH0b/1nzzsjOvzw3Vykr9t5Cy+Y8/hKraqJxxrnASgrhm3Kbkx/zCQ4EYn2GfUMIGjipDILI5O99
h/1t8uPgR5s3Q9MZOtxdWUUpiugukiUy4csCOuklKkf8paG9dr3S2ggykCjHFPYc0RgcNcpyUYxf
dwhTwejokEFVIkkvgUSuB5ptMLReLKpifl8URS1nzo4wUDYICP9/9arJPNtWXBUO0BmWGMPcPsIG
DkgYtcAyGmAQT7/CXoe1e6qyCuJfsNpKJjBZ6tiwo1vqVAGbsg6d1FUG18zFLmWeDiqP+wxaLbkN
6rUR2DvtCp+K1A/1fG7XYvr40IpDXoZ+YSUPT5Sb3HK8xKDUXdoQpK2mm4wxW51X1vg1I4KXRUrb
yaTA1LH3sBRnXWP6HtxluOMenvXLooRUrcwHjwbnyzysRnxx8CMlPuSlDlaDQquM8f7XtzEHPKlN
04O963mY+igHxCwPpeZW7wcPilKD+UsfH892DieM70BN8FGogV3D1DWwjWurS2Z0V/I3Geboj5IZ
Sj0syEEk5Q4X3ebfOOJBKIARHf8AEow9nuYiXuWGhUGj5VtzU0TbWv/frmzBcBihfA7fOa/EIcFP
oa5+1a1QZYYlylw3pfrjZJMt//dAkvx5BL3eljHKJpBWC9tRFb37ke2SwF0m7n6O6uXbKMPb13bM
Ehp+W1fTs0DpPiqYRBiRTp6U2ipzIOTfVaQLM9QXvvj6ubd9MSrp346I5PbRpEFYodSt/Ao5tuRJ
2oOqQrLmI5bXzWFrU8OJUmPMk4ecAc8IOrWVjJdIhIkQBCrmJC8Tr2UWcvKBCV9f0aMpJZ3nRIhV
5T7uAhGyEDNTsVfxBw6L/GYeKqv2cE6qaWuEnpKpPHG5NBt+k9zR6E9/vzo15d4ljU5Dvbyp8nz0
GQmWjMZTzXKlwkY+1CxPi3cREArn6dyLhppJ2K1GI86/L/ejGFeuQlvl12QLarXqcktL3Zxe1b1w
Cd8hC4p8KAJVigH0rBedvY8NFFVtE1SdZpWnhh5hGpnAV/gprO/m15fPy9XGcL6SxQ5aJqCiB3PW
S1Ax+23g0kx7P+v8KGkVIxKtfoKUdKToIf370qmFQW/1A1w4UY7DmMa+h6N4GfVDGqGHJxgqTfaP
sH25EmelZeQdl2DzgOfHsUj2BuTT/Pt5EZ0JC5fpM8YxK9eKTxt6Mt4+hEDzx4hogWabPRd7eVZU
SJ0fSmEF0AS/cP/Ezu6NltEQJNcHuvk8//O7t+kTKSDka2pOQclNH/tzOPeskECQQhpED5pUTTUI
6eqQxd4Isc3MvydCPpnk0HQhkbK2aTh83OJcgibjcdkLW/FXtFDHxeq932ICEvYxyGkiLmE5VbdM
wE7lByP66kX09/otF3qS9MED1M+5n98YP6CbJnNOr7oOa9BxiAVjAjTOlyL7ObEb3GuhpLyjL0NG
G/ZjQ9aC9WRWpJqaLaCmLbIRFJpgD9KvXZSDbboFJAOQJttdTRglAJsS2n40LuFawgB9nwHdOQLC
175REsxlX14lO6xF+zC7FHj66q7BSV2NpCkD6Wni4GkFPnllocBODYf9Erdf6PcyNohSrVntWhkn
WP5meNvnbKprkBiEN3LZAVlvUZG9YJpOVDPO+Jj6uDMdvl5a42dCf47fyH6FQyRjfkbzo6Hy/cbQ
B9ely2ysnvFAPDMvXCCb1i9Fv+TC1lWX5ve2uoV6mVnbWnFMJ2HAZFzPpryJf5oQBSbShfSh3qnI
UNxNVbcVQr823oadFlv738kPgsWIsTtPzMpf9SI3iNzblY6XU8NWHRBOBpgjUi5uB3lHaU0bkLe3
TP2RcpxgQK7r3rYk0f7UMOyqStOiKENu2uBkMWgsdsNQRMUaVqqdjMFNS+tl79ObR2bjcHgD8hzC
j4UUG3bVKUUJUQVIa3YlE5nNYb21BqdZvTNNUic+5Z1FFC954H0xl3tlWqnzOVHAkIWgIjtHiByl
Ja48WNxAoaCitF52qKZokTcMtaYMGLrSSIDCqvkEWWuSRwGlmmNKARY8pFAoQZAvusTdHhYOgZKe
VMw55YxPzeoNM/Sgbats63U+AwnN9eEgbnjy7D+uBGG06ZmgvnNCqlLZG5Lsi6G64/wt8eGMq+Ip
ZO5fpb/FuM1BnRcc8wO+Ggf5/cW+bOkWb0wFOF82HHki7A8pH/n9OmUNrARQtu115QZbQ4qi4TIo
cidY5aWa+eC6sgkCkZq8G/tuBGksRi357jYc+76JQ36SVOhqhhfeXiYHp61pJuXuCYTaCsPatiJw
oj9tWAds8ZknIjS6e+QFE+3SIc89YglFWivgD+FFb5pCO9F7Flp4xOXf5k7oyVtrNar4Bm27BjxS
5Sn+qVldyzbfeMcmUhjuiHQdPUfPKvKfWdWWnPY4FbD6OMmc8SJYpQEbhNDRZZaY3+df1t+7fgeL
M1dV/5qWldzmqKXRAG8MN6jNUEnviLnKt7IUB4D71PfrwqLRR+0Mbs2dd8nYfZiuk/B6yGnFEMAx
7DFdno5yaRJq8jAJMPTQvbQAxw+133tsxoqyiNXiQ1NGjJ+hZNjkiKFqnPbes9o+ZZOH8bWNT2mD
ftGJEBUDg8h1ZuBEyonqKH8kDKXkQYo+cG+QBaqwK4t9G67Pehk6Taq03Z5QlNioI5Mg97dyjych
YUOvKGmlJaghmrJSAJGzsqyVJg5qbrkV6e+gGKzUB/mVi/Xn/dR8nSBAAP5zXKwQKxXyAJlXxDMC
o+be/qegbneLt12a/g9ydJyUCaVswPMJC1+JldMRaczVBJ4D2v6JLizX6j1yXr7zCq9arj0h1nKT
LOx2jD26jozzmgSSswUofEVSeD0g3Pj8/utQ2t2V90BjLBOnsMXhsupkewlo0rDtkjY5OltNmzPD
7QlJwAOqKVchbqNRD3iX+1MkbumMad/IyoaFcQpqR9TNXSnueq+Kl1MIc4azbVQevgzI96WIDIv3
S9U1l3Vz6ZXWDLxUd7jKqR5GwDbQIrdkeco7rWX4UTQMyZvBdyFfawz1WMhXycOBShDY3+EHE7Rq
mSVvPy39jRkKQpYV74VeCeyVmybu7SylLviVLl/MNq4eBNHehUcSj+VNMErlm9B30g13guDuUZ75
uHNGBSYsbOBVDbbVLmf9vuEneTGAdjA/2NB+U0Evz/zdMQRwL4DRZM0CGz32I81KscH7aPKjTzW7
n5TuqKhTsxV5YA24MVt/Limuk/cD1k034XO2Gap6HwVVBcqQGqvGdlBnclwAIzmMm7Bvi9wTUWEW
aZlD2bOnmSJycnd1jubcOO7HWQpPiXlJMn5j6xvIzAI2+59Or8vAPLGYMVmQnlVbnx2sAWFIYID6
/VoWB3EY5aGI5C6QVyvOPJz08qxqdBUOtraCO6fOR2txoCwDaUIgnw3eUt1kCosfSM0aEVLQTLAE
yM30Lbj0WcXGzQ5JOkqMmFhnPoLJmb0TjbAkk05j8VVZqonZB6X8p+tbiBa8mLF9SQhTAHdsjHCi
fbxqMNFJGtWwVr8/WoJ1Sv4h2diD2a+cbNDXgDoSTVGQaH9gvGyY6JOJ7BvjFljFMePORkdrm2aL
Ep0q5/Izv1VFI6pXqCtwp9Hz3SCVcNf9QL2YSj5Qj/vFSCB8sU1NrAgpBBC+dxUBnGDeETXk5OBL
cypQcFBqUBWv0rSu/nXTZDQzlaXyMjC9YZ2nSGtOjwvUmFp6GCzkH9TE6AV9BVEnilkl7cuQ15YA
adag3wNLry1BEFjXJ2Dt94qZEci4ER86ZuGtn++I5mNf/mh4ndThLUhbLt99/xpN8c8u3YYa/xSh
A7wHCYje9s726+DDlreJWpk4VGFaGA30An9yWcjLSm8r6TWrwXPG8BhQAp4jDTb4UbLWAste/sZ7
jZ/WzaNf2Q0iOW4IqYkHHO6ypJuES/RpnwHNIALMhUA7ZpyIbgdW7oOPsHnrIvCMsmtfkOXRGmS4
zbhzU0YIqmLGdOHI//gjvXR13IKfgiyLmvuWtouyINthfdMCo15cuMTB8YR98WeS3tReGOQAyzFU
BCsJ0+gjF5KcCssbg8sM5rkfuhiDeJ+mZqdOnGXAY4iMB7obrF3Ojm5CG6VPWC0DYXK4lR9TrUmN
1JU0ut3d+yIhFFhuJka9OzoN+xMcrqtuEIFcyb7+zXbpoGRXEVDdtg8hdaqUbK6r+3mwXr9gtuZ0
1iJdtEDCfXHGuQrbhowsTuyG63deqpRnX67dUQIs5R6DD9eB0RvKKphayRgjJ2Qb/VPUVNRICYJl
uBegumLKZTtZIPXDYEy13Xb3wreYYfO8OzfGvfIaRxDK6RV45AU8+Zv5HgYJB311YwD21N7zaOTx
jRhN49HSl0uwsOnMGPgRDLnv7kAqZas68EI0cGIollwhATrJRuy8Qi6uyUHV50N2ey3I8yunabiN
LIFSK9XuCsJLbKTdd/WkkZ7qyqJ+wuqI0qrPgxs4LGxKzH6iYXLWLfjEo06wPv3Fxm28EOkqYiRY
teWhwcbM2QW8eJoBZDuAD08YW8KRAIWC8qAH+H2DCuiWGDFqiPMXEJ2CsT7KCGh0vCITN+q750Z2
ByF6dXdu29Lq88TmCshb2ftjRaPIWxpWXTxbLa9Rp0L9g6lKW3guKZSIXhvMFPP9g0scApHEYbdM
QlciMff1SIVn3bfeUFVZyqG4JLF+nRa/q2UiiPEsU+DtQXm6hCWo2xAMbyYqpTw4OiZcYMynGtqj
PL46yLGJdQfo7BQkhGFvXexx/GaAPzq4YQMKyVeXSLJ6apwVDPUaASNpA/UPqx/s5Pley5iM1Dh6
8WaEfT3PlVD5Yhv22aKuypSwKo5LIrUKsPUnkzgxXqK4ueBL9IzttCWKxvFdb2g4gxr9KxBnYi5M
4xH7Cl7ILnJmXUppSoJ3jSKnxbb3EZY6gMD/WpzZmqqawNIGYBgPoRNsINOnogRMOQi4wMq3sQv0
CjDRDIlGjxdXtdzpDUgqZm2effREMu0ZdX7EmE+MDr7CD7UoPcftLxFDtWbUNwsvDjJXNdO40SOY
EGOm/Oj9sPnIPPIGI1r2iD8tnAn47MjoFJOZtTUbes86D+DIOKmpfEunGkZ/qq9lrNHtJiqS9z/Z
5BTBQ43utLf6xLj+EZ5ZinF9xrE98ZkpxJOs/mBUjQgBHHZymh/EqvoLHr0XqyNco3d/KwTCZ0nO
Uca7pPKdGmypHDeNvIKlbO7892iDoNZ8e6Y7tsc87cqjXa5whoC94ZbhjI4Hcwa6wz2DgbmLO0vr
DurCeWkUR0QXYRW9k3H2bSc0zUqYA3PE89emOzrbSvSfeb/6ca4O2ETTgvcsxxbz7YxQTIFZRBu1
ksrfNrxRugrmilC7/0G2REC9yX/553s95wPJGV5VigGysxFyVgI6V8FQYlBNSJlQogzatges6K4K
VfH/rH8D4yzLkxWMNUyNt/fZgzNiAtnRwVMPqWbsUYe+HanzdHDtZmKmzoaWXo0vGS3pt72PEdNZ
yK/aqDrWrycH+vo/c602K0Zjb0Ocr90VgBC8jAEdKvTqpq3ZC+FYcIzVs3h26FNdHQzhds3ktoC5
BWDLAR6Mm6VTeJbqJtz9yTJNNhgCYnm0Xs8mycjc7XTy20Lh/VZHPCBtnT+pKDxHDP0gX70ZTSLu
9LBlwYu+WaAsmXiuRcKKHcq7n8Is8Z9d6/BPzfLf0iFCNLfYjnJtzbg+hBpwId3uN60NWxw7t1vY
3kv9PkjYY7Yur+afSB0SZkwvrcIVbOIn/LeBZLujS2P4RDENFqnteix+3JifUoptC8gdXUrBLtjR
lergRm3xjqk316QPc3zDjvqgb1NLl88UPmbG67+JWh4Gso0gTfKNJK/xnxve7Gy/OkpyYRztXZQ8
4BoGP89Zyz4V7Ho/thlrFmYVdXjxh3+UIm/G97udYDx4cJYW//wFQEugbJ3Pp9PKVYcObB13ueRk
9do23b4qjt3FRrlVhkv1wMc322CXb7TsIFxVa5Q1sX9+R5qIYfbEJ6K/BiwZMjoRP0ivVwPf6Nhw
QMQV/LAYavSdkD7giXe6g0GjL1i7lq9x8zKpJhKMMNxS6lo5T+qqO+2r5FUq11US46EdVOSpD1aE
p9LsYQsATL3DuKT3LV5QbC9ig+pcquKrtrHCvtK94qksZvl/wIXDgBVaOrRu0z/KtLeXfwASK/z5
sIRzRPdRtU4vveniuLnK3J0x5W0adRrVjNkgif1wTFh0YURtOcl+Px6/gmo5i8Ii6SYwOmta+jCT
LWeBDWGJvGetcM3P91PUBbXN+ugVzHg3U4zlBcrU0X5mfPizxIntU5g4uVKg5ZTSsxvkLqVCz+Gx
M8kXiGHWxhsm69EREBzb0tuKBT8HoWy1x0rmk1VxQ0oFLnejNzzduSdHfYJ0J/O18n2ZU+VpNeiu
SQfgX1axLLypTSjP9itWTqShzTOSjcztGMSLCf5B5w9F1OrVK2EisOpA1bg0Dv0g2VLXGhx/tpKJ
fl8MdaDA1WQiLCcYd/GOo97tj8Zh7RLfbJco1z9CniKrcTjA6Pzpf3WkKOvCJQZSbcwxRK+DAKfx
L9hVKw7s+jogI69FeKX+fO/IyuuGP4dw/Ow0bd/Kjs3Z8BjZaQGMlG91M2GQVFmX6Ck50knXZMF8
184EJ0RcVeIlkBQGUh5r7ccm3+uoMutdC2xix9VVe+OILwxlkIS+d0lnHlRZhozV05IpQK1dNkKd
41z3P1GtOnr2foUS/jmpv1g/qF5jjLWvsVqiWrMZ2KpyugB8b/0K6wylOUXpTqeIg7u2gfNfsYCn
Bq0vm3qfhzQOwTHi2uKRxJOBZ0QBzyf4EqAMRR7GUQyAzP+Gid4rYk22V8xEO1sLyCr6LlVeRTDW
sXTomHL+r0Oxy+LXvXLOv6fZUzmafhVdXhzQjmWmPPfKbQP+z/QE2218ISBfuFJPOhVatVw6dzBj
XotD769ZF38Cwjays5nGGrnldSgpTurGMLWKh+AY9+9ZlgUmTOmiDfyg7q0Yhy3zMOtc/ipXmGyF
beJJFcIL82JGQ2MUgEB8tQKOrJr04HANkyR5YOdi7QpthGfud6Cw9B8YBV0vlGZVKzEo7AhntHEf
2woVfah+OLySiCtQpSiDbfbB24yQiGUy/hihsLX8GVSNDvPYVP9efLQV9J3nYR6x9FjwMQuod7wW
eXhGRSzCGn0c7r3EjQajXnn9yx3QxlDm7ITgd7+74Jgj1EV9dbQYWJzM4gU/7D/Ff8O0fM6CWkfV
6QzLFg4cAwlJUTqSSIT8gAkv6tVvvBsPTUY4Npug2ktNwpCj/lulxNoi3/KUx2rF+AplA0oqucZh
k9LeDRfiuzO2qOXPC/GXJ2H5V5BZjFIhqk16KkOU0wfR9nX3hz1D+PmQwFeKLIsW2h/7uoXgMvNl
s35wXkesXCt5VZ9ISJc3Y39D+MIacZvG4akEKaemwXneaHLbwKeJNvzeXX3ph3zqCPtmkeQ3QK8T
Tfm4GuXz87gVrqLpJahjRBli+sLex03jlgxTR7zM2iQjedySIa7DtB+qkSQUOuSztQswZ/6/O0CO
Z4J/9weY7wLG10o1ODS3PCZaY7O3hWJw8l/psL7iwt+/aT47Awj5kBX4px8WGni/FUmT7fUpS21C
jpyU3gTSbsP5NzpbJUIYXOSEr5b/o13/hv8KXCenptZe73b/jFuF98KRSE/RPG2ju2V4VTj17kJr
YPnR83DOol2bT7H8dMYpQBVuKQCJyhUtDHvVZg/un/ypYlsb0zfSGMyAku58tM9+CgFJB6ue75Cf
i8Y3KbFzYIoX2NsRZdihmi9lmVniBBLj402o+FI2/+SAC4UC3/67HTyqPkboL2wovrVHEHoLqFpe
7klLlIzq4ElSvmAhaHLB9jHBpsZ8loobU7lKNjXS2BsY5ItZke2ZFYClFVwF64U6rs9q0XR/PvoD
BleVvybEUXbusKkV65H0spaxTdfMn0/v7pzbt8xXVgpj88bmokziu07L8kmY48E5lxoTGsetYBj7
Rk2Yb8v/HywE2amfTzj3b/3gRYEpEaiKAPNC5kJNsmR7K22FKNXOVn/3becj5qw6duLuvohZSEa+
EpzRBWha81bxchDceP0ZxEXSXXuLePxpXW/bQowip/ep4MpPjx7xTFlUILXdtKzV91v1+R+7pkqa
mtHD0T2HTQYsxGqkt5MAbU4poq3ebA7ra7fbBPk+4nABzjUfMJPqtGQgxaviSTTdyA4doVEKPTnc
04TlVeJFL09c1sQCCJnBNiUCF1C0ts9BYq1GjL0SYUSa2otXndzSUoZhJmZw8+ayOW0fxY8ZXyvR
mn1cdRg9kv/AJMo8zgxQE+6XBK5i6QN+nFhDA4fRHAfReieXg0UqR/CGH0tkvySGXWX/jVTwOEOb
6zIFgV4jfYjfWljth/dMdnw5wWmLelNwS15RnvyTZotte+YP4gZJZ4kGFKzpWpvWGVT3LyFavoE4
Q7m6XJHRhtQxc2djV3k4gWiG9/ZbJgsSG69uO2MpZbE4cqPxwwtbL2A5g4bioPmL2RSk+uxnu7bV
Y2kuYb58u+bPyNspE/6f9kge4QD2nnlCM9KNQ6cvBFtjUtB4896dT1GXiyr6RUpQwIiZ/cvJW6Ko
F24b/XlO8rt7pMoKtBcQyztplQmprns8xvvJKqxCVTbYGZLrAgIXTxiGfeFNKOj0ZmEDsHJbAnul
UNG9XA4zwnFzS+7EenXSqnoqkN4nfrddZhi8GCcq6NLII6JwpjLqey9RR0ogR54E8dGIFErHZd5g
PJ9eehy6bMTaoZzqgon65izfyIa4x5VDchqZDqba+aPAQvN7O+Cw8o1FVPmbqZ9U94rfDiUp5Rf/
C2q+HBqWbgMRJYov+Mi6gODrQUFn30FkUNQU8/Gl27bwaH7yBlTjBw5pCoC5MnGC/3bPQ6BMDOQ4
KXkK1v5JSxoWlYut+k5pQnxfOGRGcL5nmbTAf5WdZAITBBCJi3jaX5mKzWQqCb1j/sXeoxlE1qks
P7MDDoB5jcdw9zgAi4ZJqLJbDtRzmRgbGddJ8Mc33KP0Kb62ldwp5eoeaUwoHcfapjBPuAMniuxs
zy7a4UgZEOmUxtn2AKbFxlECPR+kxieP/7EBNIhKaXRhCveqyKe8yIgN37yI1RCZIetuUjL84WKV
DV/0eY/pRJfGIIbc3EUCsO3tYHx4XKTXEWCLebkh/fu9fOP4PGdiDDh69SNu+ISd+g3cuS+DlsW+
nQ2VO+wEyGA9w6+Sd3POzZWMfTuP8ZapRQRvGrzWiYNBAn68skgzhOkP2/jUo3cmbUbilkzCGkEM
qiFOH10iJYNAPT/RPbk8BFnAGzZIhBhXsOqRxKAh1V/VKt9G+bov5L7ijXe6V8+jl+iPMROUOMDf
OeYRhG+RJJ3MnOcqtQKThBbtfMs+N4iF3CNvqwYKC+kKPYUn2Y9ZgWoistJRZWbUhbXA5c3a14li
Nk0h+B3Jwfvjq6tkOYjjfHjJzotDheEkGM6cealSGJGiI1at9crwGVJ+61IY0ySBQ94BdBrCz8RQ
TsSd73riXrgrOmG5vv4+fKpgAosVQqWn18Zm7sGnUkuqG3iB59MJ3LTV//RdLh+ytql+5quo3OQz
DMo70MbjTIAPJ47zV5jpPXlfhcL9nGtldODROoOtFwFquMIfeIc7utBf74duzV1STN3rGkHuHEDF
pkyU9Y8WUDm/HgD+o6C2h9xVoOba3hfUzfz9V6tjJATcxWNUcRWwzU1GfS2Umt1pCIhEzpa7N1sd
+Ce3sHkJ4fIHxOf8ZxW7S6XrG8P4YrRY8KOf3qxs2bJcD/j58IoH7pnleUAYcs6C92uvJpyN2M3n
usYyTlY5NRqMN6eq8iIVu6zU1+yFgH2eCKpHg+kYNgPPnNbBORSIXWRf4gMS7jcms8rh94Z/Ayow
TgFGsymwmGhMV212GCLSHRtUwr4V9q3cNIL8OdZoFJvjhqhwFMe6GF51AQhltBC7V72EYHow52p3
J+0xwfdgMXdEvJ6+SjrQOGMRzgnaTDUn6wIrc/VpJia/CTll9J6elSDraNA5k5T1VfntdxEKJFmC
EMS5hRJr7sexPhC6tWmgZ4nGX/Ryl7mHqSmFE8F+/i1+8Bh62mlh/1wwjruuQ6QYZXaXv1H0rOfj
zbk1eVh/R72l06lQGi2yPPgUX4tfTbVDEK/IgMR+hiXL9S8HJEjdYs1NiOUg0LzDTh+O4kzg0q5M
2XGeuSLmCp251hsQrgGC8w7q2iIZLPm8uEU439jKVVq1NID0u/yVyfWzgwGKLpkm74122BIAvdEY
8bIEDZGusMHpXeqYUf/mmb9OoK9etPitiAzvMEB45s74RmGk5Jfw/Au1QoeeDEUKjknoST7u09qp
IVJ+sovHpYjZ9AVicvWb5jjbYwx+BVqE6z9eZpJIAPErcGQOITaOjbcpmGsgqIJ1cLRPvUthzXNV
leQdPafw2VMJY0B0FmnIj9jc7HqwXefWVcnYpg1l6UxlnSYjl+pCxe85BdTlqhCIiOhoza2Tvs5q
bgD7eVRqqEdm+oCZj6mQfTPV0WtEZCL2b85bNwsBk+9h4AFb8gVxsAQB1xiNtqm2DNm2UyfweB/w
L5i89ZcjBhqqyrKqcN4B2J2jym5g3zdG2QjAq4GdMAol0qQjSyF58r8oFxOoBPysLQAot1rLQ0WD
50+2AaJU4/+35exe7VL6QueASYMv79wJvDeAsVjV59sUPGY0/UOHej1YG7XgVCBkmAreZOZRZ9Ba
wRD6biEBgVcptC4HvzxECDNdVsZrF9x56vq/J58bMpH3HXUFd77MDQC+bTDx7FPGqJ2VHZsHOS1L
R/TwFUjZxhQs3gpYJG7/E7LrJ8HTjIrJrEsbPKoo3XHczAx8Jhjx+xn1fjNDn48OmTTjy6adCHTO
i3t3i3yDYyQhuF9aUe0RcG2yhAC2hjEsmwc+vUjnGDDm6JfOR3lU5mH5JiRZJnR2zozVzGh+LoSj
Jv1yUagVCnaOI4Xb/tl6D3JL/Dv+IRfKMSLpvi1Oi4SkKcj4VQUZp+Z9sawNW03vFNlchfRLQxV0
BfBJfDgMEhU6afh/Dbkwe9Icr0Bkp1NemT1kPF7oCUQ5XxZsiqmT3HSNvWeh52Q/aIWPkMshPchq
haW7YuCmQElvrGNQZFitKGtcaoSwCwPVW0+fGeWLKT7M9wjCZa5fLvH0jah/ciuHIIDZX5d068o9
iHzlP494rqO/NdvFrOApRt1SNY9Vw+13rz6XOrMFZu7s20mA+mS3O9EuJI1LOQsw/58ij9TMozHS
qXtID0cIvyCUhOrwv5sBUR7mON8kJ0x9nwlLM9F7q7fhTU3CSIXIQm+73rrLw2oeBnK6uW5K+jpu
ZTxk2CLOfH3xHkBqNdDoahd3IWk+nuL7aLwVjTadicKqZk8k4WGHjOWhlEQ6kYx0sU18J8KGtme1
V92GcxdbCELmoDZsxb7RCfR18kckrzwa7lAcGU1t9a51a1/4Jv034xi5Qg1Tg0Vk0vs+1dJYh6sx
xfkDiTs43od/D7Yo/PVXPfomfLMp8ELanzBBDCMhhRrs8p76qPl1zyZqQGGRaGoCRKVr7jX9/cJW
3lEIYyfM7GNO0j4GiebitSEUMP1ziiiAVizfNJYHx/pAjkz+LzANqFUAn6IJ+IbY4Pl/cnqL/OBO
jgHSsUZjSupC7nuq1FNJsAmIuaho9+Lx4SZZREzCpfqyvehvzaRuatq97XoeSvP5n0YA1ybWlZJO
mwXe/U0OulaobSWvEsgSZt/acRNlqxFHH+5jfF/uqSHZ5Je14AOQ7BnLlI6H6Ri2VNBkVEa9Z+16
S5pF26MxW/NY3ilp6xftsMHTGdVnK0r68XtCdm7P7GCka9ApFadUL6ccWQzOgEtrEhfg5toUZlD2
ooIIZp5YsmPaQwtiLZ3K47uot5Cau4K+nO2bUSS/i4mNEGCa4o5YbijiYkWuyOszW0KtRh26IYY7
r4Ja3+GKe95GlboB97BTEIsr7IGXLaCnJ0n06ABD82ApcjFVAG6zbqOa4fHREeIYtErQSSGoJg20
w0WKF1CbVPdIAQ7tvBM1w1qQyDOlslpVLbngo3tKLL5KK32Kyy+mvOpGRKlz/GxeIbtNZojeRC/4
FP05VqxmHWjl8OwvbY+LZPidGAVvW3lOiFe91uvPfuebC1+ekp0wq1KzIQzZjkbQmFuRvMVMK7G+
TsFrUh7sKnH5AjnKkJPjupm6r6auPSfQBsjAY2t40+0g/8a1Dt2xjhEa6iobbh89VHMTbjgK7qSs
hjK24USAu4bW9RY0W9FXJPb7l3W0zVWRlzA0aSWKR9dV8HFuPd9TwJuA9Zxlk5cOsr1ZDXGun31d
ATGCRTCPRWOs/p4jYn8pyBGQhn/49XSNMF0Hs7DzVlMyv4ijVT/NEcL6KHubT+AIqb2GBHTPAvI4
AkBr1obk4MBwt9ZUaww4UySRrjAOz9UvV66FC1kLgKDYS/VumU2RfpmL5BxzYXOYWIXBWqMUCuoq
raOIu0IqqFrY1UWfKUKk3dS+lb4wLqK0AAjNwtcjm0ezE7VcQFBe4fNR8Kn+kbL3JyxdzftNBWLF
te9qTSxuaEv/mANsoKeswhNOPX98jkxIzOHC90ScSg9uZNqQpOUh8bH7cgKOO+k8KAC3V0xwKS6V
7iDPQnGHkDoXeW4RxW2tuF/WHrsCelYeHpVzuKC1DJfTzUUIOEgFLfcAvqGz93XGKxTQ6r82TEAY
9irUgCzOBNX7MrcPVO/TCaDkhrjgbvOQJAMgVZ0irIjrHCBqOaqlBsD7jRf7EFcUzvoerXpfTM7l
CBM/kvo51VmXUz7pdXbkknnXyVDAukFtGgvoezjyYdln6OPKr5dtuLKW1ABdKCOXCD5FSQdaPYVw
+6A/yyKyEHe/u7T26V2+mk0wR/oUwn6rdZXzYaloL/QPUTFPlemK5vnR2YyyDuM2gSYfzn8MBOZo
zGl/cdLZrFbmV2hwPK0OErkjNTlp5Jea2PJoMMMOkGUJrxAgoBld+3sOAOSLTIYNWtL0MhNQfpNz
woph2Bq+x4RqEBhT3J+WcRirMyXo/Gb7qpsTvtJY8Dkzz+oQoQzYBEfPyR/ui7XFJJM8+Szpdjd1
JWAR1tSKaNpAxD9Ma8v95BwOR3pGjDkWwXEWmS8xsRlhcO5x71Syo/MxjQ/l5WHPJq8yd34HlLph
e3tSmp7d+nC2UJhtKxJ/I9t4JofF1Siki9XaNXV4rHiL/7sxhZTIZnhnM+oPFH3rsEC963CharPE
YRfFuFxgI16oT1+iE2YIMWgkv75uZZiFGkIPO4h6n2Lc5Vq2tpv6nYpAZQonSbbJzaTqotF7+wcz
H+k8cpxu+f8/Xfyk6gEd1lldAUy0TR/u3Pwg9Qd/tCs+kAVo/N+HYIoXbOu8wnabyu83F/MdH4/D
X0Gsb3oey8pKha4SonVpCAwcAI5AcnBRmLsf25yP84l4bHaY4CrxR/Kw+QG6ZPxp+jPdVVEp77ta
Mv0aL3CkdG9EY6zFBvkXBoH4NArUq7l6WeXAyRgRR1LnQPGerYPp7N0NBZ1pirXaM8NqnfOz+Set
bpzGnLXoRcS3plW1Uta4NsRNygUOO/JumcBLqy2sus+xp2lgV+QjV21edSNJpdmjHd2eDue6da0+
0VDqASGMnGhk8CNnUUc5+nqf0Dpu/37ujIivle5Yx6hchNAv0RzxmAvgkvIyAJlBxVqk0mLDtHQ/
vY+PF9zttuTOredZMPTiI65UrMoSxbbMr6eVwW1Znd7MFQCdpQBkVBNpDhukQL6aV9Hc2qJ/4fjW
s6UONvj09gx4U3T1t7Hzjj0/ARjbVOzwH4xIg+KUZ2ME7oWuLR5PaicKgIdtgRsKWnQ6Cno+/AxN
ODBT9Gw2DFXtTEp0MRCgNYf+eA01S0yuna9bkvtS9efY1s5n8hdyXa/a6Ib3/ddu16OiqoUP0w6R
WAblKad8PXe6ShBeC74GCsSf3cct8am0t6AdvxMWpoL5fk5khsBEOXJz7UnAwjXgGZl40bc0f6EA
tDwzYtN+rua4R+oA8J/3K5tuYICH1mDFQX5m1C1HxRiwpWr9AIFOV7qb6+snQJmf2X/gREl2Z5Go
Q2S1OQq4jhe3wWaOEkwYtqorvRqViXkCeSdWnPYy8xl7sfuEPeE+d+b+fOyjvCeSInK/dtL/zZ4w
mImWJLaJbwNrf+y7tsLN8OPvgollKNYV4Izq6wDlCkj54BGL6EuOFdv4+lQ9A8o2lnlLnrdHRdJO
ziXqJbwRMpmysnozzxLHB95bR5CmvPFhU9Zv5GI9KK/zvyNmMta2HB8j48HcjCNMllRw3Wf/pTPr
6XmlmSFyvayw4ix/x/hwPJ2wDUlzL+M/7zunZbLhFwswv/dKiTWAEGN5LuUyIIydyvsHU8rkd0xa
L4/rairSiIN/VSyaLLvBwe42N5AtCoW2OMbjbjy3aTsFPRROIeX3ouOaMCg+LaQ2JUYNPwcFbzqi
Ks8od3AStru9gLr/44qDo2EmaW1tM0rvwiEn8oXpHrYs6oVaX7IVNyohMbY0vOmPSdHbU1fwm91j
2k9wdSN+GkTUqxHIvnGtdmFMRGCk+HoHGX5Rm55rSuMP1pO0RLDbJ5NCEC1uf747S3lHteDkhtu6
5+TXAHDpM8dnSPRFS4REBQyh5+H47dcTaqdGBq09MFe1X7eImSyjnlGxg3ceTQ5ZE4UKVzXNpylF
8wWcmzYmRhULMW2jL8BErxvaSwcuFalGVrTDUOP+tmmkWIYkLzJL/+umHiPA43IqdJTy2Xmafb/6
URk6OE3yQ1jkPBPRwXz5ZkD17m40Wt6uEAGyGlcBhaRF6dyKVJ/nhofJj+SEKz6M4jNfUj04vQkP
thJOkTgBoglUiZAs6Pe84da5aL0VTaoxWGPnWThfJ+HHsE/OZxBTnymfdd5ehIirkWakmBwfJ20F
bd8coVWMmPYD1j0AEdRM527mbr7Tu04KNP/GV3EiRTfH22IVcn/Le/S1jaWQlkFUC5TOiA+qLBYu
JeAjgRkMUb3JeTAiDet6YDj6eJAsoR1F6zqau7NxSHVrHyHZi0rvpSCMgJORkLV2V0G6xkzZL2Xu
xfadZZ73HdpcHHIWdWTlKBAh4WX5j40kgkc1+Gqo7XpmGAUUVtKucw4kFFk8VvP+bJOF1hlFAYaf
rzErMINmD+M4JgRevG0RQLCM9yhfmrWYgEf0JxJQK/5lCJnSLqdB2+HvRYiGKo/92SOr6w0YvhS9
TPPK+hxlOw3K0ZPFij9SACr+bMoyQsaKGR/JITjW/8XL5Bgtcu7w4S7XqcKINekcIvtm5LKKbGTh
H7ZvpTdean0wssDKnbJdyXB/kBo0HVkASe5QYYqLZJvd3DIQuxCtRjjdAsw+sHSRRtu00rqR9XMj
YnXicGjJKQYuaD1hcigYV1Ewuo9wiMZ3LfyQjc6zcXkX/abGFVGNVXr8xLgEt4Yo1GYSzY3xzRl4
U0oO4r9GK/0lpKbvjHm8+ykCrtCCZD7lqBE9jRc40ayMIbORtAJGpgdux+24AdXzrD0tNUkp8GU8
P9BN6vuhoL3W9s5QHIb/WlpHOu6tfU2DeeuUR63YB02d5/oWreoczfZohBbAq/YxPFSnnKtYskg/
01L095kMPyXqI8eZZDa46O5eoXRrFijKprGEQFBgaDZfuw1+oL83kHNYFoIYx1iMuQchHeAN7Y2r
z91MTv+Fabx7WL2u++vIe7dK46a+LnV10w2ck7RV27+AQuWq8+244X5NuXbBJltJGr7uWq/k+Fse
axAHWkwNk9EX2Ch2SZsBRfg6vhXBIP6gk8fT16YKJS42rsVmTykwtAaMb3O9FCMOM75AF5ulmAMB
fpRY22vVCVpuZSWhD7hXWfHKfd7FQFS8NpE4SRkgeaKJIqQ0TqQvcvNr0443tjY0/awM2cyRXD7j
Ktl21HQp4ApKeu/X/sIXVLiheKPJWEo4+e4tFrv4AbC9p45EtQpD96rlTZFUaTa7oddpQS8OsgkH
yklCVTdAHZcQXKD7GgkmgVjnsmD2mpSZIVkIbjr1Yh9/GOaAx3aSShL9cOzpum97cnoLPgih28Zp
Nf/0Va/C1ZdT/i8GshiXw8TxxY5DJ4QPsQ+HMFVTTI7xCyy0bMNPKa42mIn91DPT7EPdWR0kRTQs
QPFadpBVHJ668NB2LE/bcflJJ6EFVa6RFFMkALZsgkW96tbMTKm1USmpCiSs5kYQOMivt7mb6vvH
sFXWeF/YmrjJTBUw0k0BoOxdYJYr4JW8rnAdjhnWsvT13NSlitD3v4DSVt6+AlOJi1nOE2LW69zG
KzyWZdfWqlgIwEQloGapKpD7nr7BD0DWjONpLlex+FYcx3JrFmtOdVC3VVQpzDODxEnGmF0+mtsA
nnDpOUa4RSFNWs1E1UBdui99nvAbyzKH6pGZnxl7zQW5Hsr5pLvce9XcDuh/0sDhTbC/nguroX5c
3UnNfVsOhwtMyU1dfvnZ6OzqSgrA3mCJvUJnpjmCrUvGn01zOdGsemVIGhCkDhKo2pqLHSYBJq9G
KJD9jm+x2Yc4V0Ig7btfTgl3HH1E1zBH1nKdc+/Z8Qu6BTBveuJDRBZdza4+GmVEfLuCPouZolXu
aqEhPJ/7Y0Mx7NT5V5qjxTfK0KmjTlaNr3GlT0qOSRhP6Zzv7ktZmkjmAXRpg/w6idAaFkYso/LI
7rCksHQdt2pP4E/IllV/ZvYKw4TclY75IZWHo7UTNylWZ2FswcMC3DPY95qbswl8XSlPEeNKLtSG
SxQw5vqaZDg59E+xWYE2wZnS4/gz4d2BCDoAIQNYazhER4V4HRd15AAZ90TK1fGv32sTaoS/2pVu
s2+fVXPqNG9nvmW0R9sCWzwR6stlltvCxsA3rsTE27j7E5OeaxmDGw1putixBPY2gO7IMr1h0x10
f/fWcA/EAnVc40iL1j0vT61a1Z0iLO/3ZBEvB3gki6i9pGaIphlmBIBdvfY7mHvyHvNLNOClLikb
b36wTvKaVjWfBmJdJU6e7MWHSvxhazhlloLu7oi2AyTL2RGRsPLDWMzCeGCESkazgJuNK82vXvKe
40ODGBWkJjorVf+AvTo61TOkZXFlEITSVrDLCiIdgyj7OdLsU8R0bVjj6L4YvMY4QJzfu4cJPNbr
HrY6kJbH0IoHkwV+TNnRGaFqUWC0pvXw8FR5/VTGfinGXSXEKg06jUe4iWtMePlTaTDILKSZbQJL
e8N9NsNe8r8+xczPGKGeE4wwdGUbhJFMjbGl8Ii77zv3eZD92qWab5zPDPBPi019220y7xUdrQus
xrxrLf7Z8DYUOv9JYYLo1BtHTpY5iJCzgB57C8kEKbLjLkIM7lQwijJaz4dyC1jOdz8P8gq8UgLx
B33Rhy/zksl2KBIiVN5M3ackULaWztCQo+7mXd/3gyVH3C3j0VqzMHs4E2eptzl8lRfVrPB3DeWO
0rv3GbkSjZrSkP6NiYoRxuGRiBzGb/UpQvg7b6VOAcDTrtYLdxwNr3J3oKYivEkx6VnYONWuEvI8
fM8ebcQonBCghGj3qlr9uWiwXJsiIw808VaUrmiq5GBpgX7cjHJp4Me7GnrdiY9X7Gp5GNQfEZsc
yWE4oZeuECh8lobtzdB2K9FD7fXuB0eMXc3Bhebhf5OuJFKD6wG9JzIsn0sxcBe1Ca5/Es81qGBR
0nFWlnK+BuCoi8MfDqZOOZoy4ytb1gkplPZa7YYizm0kTm/DsG5p10F6E3McCNGicWYS8MDzRoUJ
rismdKEnpoSiTTC7TEHk4P4fGz6OEq+O4Z4Gzt4j/9QRZNuQLiGHUNWOEOmoMGpZcPX/emj+fkL+
NXy0nyKMA/0T6iy/VHatt7FLgnKOFNRYrT3Y43lkZg7ksGMKHGZlkqdVcPr8+56jli6FoK71HjYc
kaJ2voPa6tD/3gYn8stHcYep+rdx5UdKgjNSCU9ElBq6syv0PmSuB8XiHeKJ8HEjXvCopiWoW+cq
X7NtO0iA+YxdKaRx9zVwCbmmOxO2i8bg/XCdTZVfXX7SdbG1l/hVqd+FS1/le+BbNQPwMmk80F23
n3p2tkJOHCtwCTiZWYVkgX88ICySbuVkHKsn993GSlzfi7x2So2SaKJM218EaRQFfMEawzSO+qwc
m9cY8/h4IUjY7q9rg0aCd/anISgYcQMCYP4HmpIjfrxHr72eF+WFzrwPl9u9ZJSgNPpOsGhAYYGQ
UAUZi+DyEtsUtGkNO2CU+EMIIFjTOnLvQLvsHKftnUDf2pG1gKLd6Tku/YFHxUtdIXmCcRMMcay0
YaRWqEZYQixM3lgFtYm9sBysS878rmUwqMIRy/iZPgMtM686oP6jdpNiW4GHV2LCwT/EkpNy/eck
2sFQJiBP4PTEoajFeGlaidIHZPsNMCG5Qwxw709RW3HjcnxxAmNUaWi5CMMCGkyZHKyScgGC7xSV
lAF6qVlu0eGLwjCqqD81Sk5zfg93ugS90O5ja4hWoprGGN3kdWvAByAuYPZErHryWfOMCqEAjxwv
I9QpHxZbMv8GyKWsuHhdwj3HL1OuXnv6QB9oYjmgAIkEJ2TrjSkQtmVYO76b8dGKy3FxYkafQUUu
M7oKqXoymX20atQ9ASiB8ct375rlf7603qkzFEWw3bai+Omqs/xpje52lirqh4dNR+MJn6MUOfDI
3Ibt+Fjlekg11euNPDPZkATL3CtWHbo20tJgjgxayZat/PsRnGb3BHDWkx+f2ol4ADJNw5hpd8Nq
6Fc1CetpflQxIZxgcungRy4fq7a2ihk8qcawPYVURZZC0Ire94Xn+krnOECPGr0EA9Hq3h+j4+5L
lyHa4I8SlmSN1hGHsv7+cXINygJ6sFb3KkORoqAQ65kEOjjEmH9HPDG0VKSjRL7jPd/sCdbfYRAV
aA6gnSm2bhJMJo4vECDB4K5ttc3uFEtuez4HEpWnp8t0gITGNn0DRMRt1s8iI8P2OL5HFEv7/Agb
IYGzQHbNv7eloiqHrIPGTOzOYzBvLqkjQuWVJa9iPzrbfB7uaDkzhQZj4c70ZZJNKT+o3i5Csk1M
mCw5qvmF5bikYLRyt8NBM0GISsQsa6oSk7G+e1dWJMGiwVtcUgQOuHVX+McgfnqsPnnt9apoosEw
4ejkoh5Ru4F4OgFYDPEiNl1W0YptamL2+lauf/mV1Lv7E4m+/wedVrz7CLAW1Mfm3CAKc9U41rAw
6VvREjwkF7RyK4tlZACawRrvzEhouvG0KI/N/xr949Q3lxYR36GTVtQgXBDM+cdVP6ef7L4UISrZ
3Cnb+251mr9jntBR087XN2i3LEGQt86mp9tKBJD+IPelQlXeuRrNvBJaN+SHbI1FmjFZBZ3f3fna
0M+y8EXl6FQhkCQ8mWfhVgREiLYA+9xojdKST0+7zrIwac8nxTzfmkYXwxloyl78O5y5OIBAMAc2
TfRHc9uxJYqpF7vBKYwzRRP2Hx+epRgoSMKLO+KWW41UiAfw5sxtALwr6dLqscrxUe0kWh689IWk
iJF9kgPb3qdGx+PiqBZFgRJJ2uOitUw1WlwsAMb6JMNL7MEyHhpQT92WyDanyGQPBQf8HI5790B6
sQ7VcdI9WGpt1n6QmwyvZF49YhqIxIr05HqoKyoNCQiWEDfcH6MdTWGghZ6SqgKbfpPF2xOjTW7h
Fc/isf2x19T95UeUScjy0ujzGreQG+KEnqiJhSzrd9vF6omR+Kd6QXmvSptv0q7j4PueECLiFLH8
IcfzEc2XaKBCSKb1RR3vEJ0uyrOOzo7S04hvQIFc8cs18fTwiaJkpd9U8UnHkzLemNeVHgNRJ96G
sbXA2VknY/6l3cEuu7z4O5GpAoVB9RsYF2wUysnoAs+dh7UbMjopCNRH+QGhnz7ebtK0thzDgDVm
b6LAhMGPNaf7iRj22jbc8boJJYHY45DK7vsWmR+nYvLoX0zm9tQmUr0XeFTU7VztpD3iXI31fzDt
4p2xOGT0+AOhw3zBwAcT33kmC+1lH76reVsC9m6by96lICmHXPtDwgW1shxah82XeNcHIaXEkBao
Q3SwJMDKtXjk4Dt3WTp+bBRRavby13PkVXV7RsPeAav8xhkr/rirnmfX12otZsdho0xmR2p5OIq4
1KU6Pdm+JyZJwHEs5QEpChwUVV/nNUVEBp7hqHJ1G6Iw82UEx4+l/+BlbEv7Je8cWsvZBLpAfdAJ
RsB+Y9OdpOvZhTzJ5zg00KHNIipaIqgVtXLh24QZgZ4FNByzc5Up4GF1DsB3SUP348v5gDUtKUku
wvqELvavV/3V1nk7A4bZ0yEkxm0pxWb8AJAr6aXa++cHO57e5qTpe4SCvYYCCiHQ9cOGjoiwmdqY
UUDuiwPIAOczlWk8XLuVdyFJt9E9QgrWvmRGLf6EyD++iY5pUQ2TYLfDcxzVVbiJDX0f3ebPdYY9
f5Cm91Y2qF2vYz2VsZJEBbBfCtyY1z3+S+e8Ib+MV2kGEPTQw+rsJL/c9TbRL/Ac4nFZJ5TTsVTS
ZNHGYZZ1rM3atyl3XrtQVvYiUtcHjHx/8b5dYTAM3hNE0MTEffYFFMFyst2dqIcMKoN5qMayjB2j
oz2jkqQv5WeSdWk/rm2WdwrFBuWIuTsq/iv1JPtjqznBkQOgb+ClBanoQyuCFS5nsGm8gorGKPQu
wxG3PtfsL6otQBN5YpLSp3+G2QpPrIAZ1pl38ueuSEFgB2skKH+SgDgm81NnqlgGYT/hPpvsXz46
D5RN8DUoiu7JRGgpBEslK+f7VFTHcrspkZ441SVXbNpAQxeyPmg6IwX4hpltfnUz3ugstcK4AYks
M8Qrbhi2zwsC92wFS0eiUQDxg/gC/YRa2wxXs0GtEeGHYCCaqNHVSpyR9hw2duUnE9jD/nQ+4reC
oTpEZNEufdISE3lr0q2kIDyhJ5xc6E08ueuwW3sTLnrFdhtsvqhNRfDC5JKAA6W9wVF+lgIBtJrH
H5rwRiItNp4sD95hu/dqJ02yPhzdBtFPNGsWLggn8m5SUjeh/AOQN2be/N5e6O+NKfoIU6KvL7Q5
kEDnnF+zolA5DJM9+ewFcHB4s0GHH9wCxIRvoaYReRly23tB6DxIJMw8GiQkTn7+4oBMJT6opQsC
UIgX2uMkdBX2WyDVRqE+i2uxtUMpc8mWOIeEBr249Lnu5JNK1guuZeminDyvFAm0S3S63/dD/fkR
RBbKzV7irbQaeVA11ONuMrY5fKmn4muymjHZFwLQnSQUvz2C1sdaH1ryVBGREhNMOg/9corg87O1
Q2k8EW84dna/6caD0eNubwpXum3uUvY0xt2cinQd2zkkx7yiRvK9OolpXuoWUYcY4VNrtzd0+Z+m
sj7RoXzPKm2uXijlW3FjRr6kAD94gq0xRuQJ4fqEHaFqtm32LoqPR01EoaA/w4PePHDSgwUpkM1h
OChzSZxr2NcTzsB+fX9OeNzI3+DIlFkzNHAYoQahkR4vXuI5Pw6E3OQ20x2WubMmtp8pUCV0z+bL
iZHRsE2ooFPurmHjpiFsaCy41dfeBLIHC+KWr+y+Yf9+nSAXDE9rw9kbXHI3fDhyZ0EcysqR2F61
aTu4B6JYPFjuMHcZEuoucF3TBFncum2rx60TNrfZP1nUJfeRcUo2W2vJSAZ12VR4elR+mRpVNhF2
Wz8UfTeXrgD5FdYivwNO/6f48Y7v7k/KDGGnYn/uQLhBKL/QAfUGTb7dLDWD/Ft8j1bJ+GPPiH3c
1Qsm92vVg2s6bE1xlPsghkNa7tje9YL7JSXPCqogk4XmruwH0oF0MAT/b+jj2/MLcFSMgqf8MLzW
PN+L/3WqnOLRbJnWEXZuSc1Af0GX1HBtQ7Vk9tq66fTzcZhgj57TZmlF5L5La7yOudnlY3Aa4kZz
qIaHPAjJX7htbQ+W3or9sS4Ch/1xdO66kkFfPtfoBZdz7rhYsCzqAzj+JbWFqNKrNyCYjrEVmF5h
cCw7VN4AKDczNcM2HWNhgoraFF4G7jckMjKbhERsU6Cm5ZB68xVZo2yaXrcvIx6vxbt1q6+LMpVv
HozVG9wv9CZ5K0fn04JGSM0nkTxtDGzLptYLrzIaZHL47hJHXfcIiNdolnYSnEm3T1YP2kTg1bgy
4UixRYG+R8IF1OzrKLzK+3OIZOeZ1C4/SpvpseFASKFhdA3naV+8Rums18kfHS9fHi38tKqJQdfS
oefHvwnxRjAzAO0cvJoWsym1y/v+Ha/IcNTuSQ6OmO+F81JbMV58B204usRC8b/REdETWjBk0QzN
s+FmyDdIAwQkJlNORvUq9iQsLQbxJoqFaZemPoDkRroK8ET9rmBpSNsr5ABbmVXVhNKUmwXOH6lH
WcNiAq3WFU61oEpKhphxtbp5kPg1lI1ufd9ft7VkHxHA0OB51SVJUcnvYgXvnLbzw41XzPyj2dSY
hH6I9WwLaUrns5yA38LktYF+FLn5memOv57W6UAR10tHuqyCQa/Fge8KrHS/PCrFfbMxTLAgO8eg
UMTIRG2uP0ADI/WApve6REF76bFK6Eh50ZqXQH4r4yZN8382rLSurM4JOa5mZqzj0hOAhmABktsz
3iWJaDvVdSt3uwEvB+nbOV1FO6fEqH8gRo3Eac7bozet/6E2Nat27ynzoRQ+4t5VKfWt43SEIc+5
Z5rNq9GNGWG+y5xP3Y/HAPdrqA70eg6vJidBdd+MlGVncaGIiHEZejJkqTqp3IpdJ6sRDp1/FcOB
uWRM18yCoRfZmoD8nr9zPynl0EpaekHJux7WoojOenu04gq6GVsYDM5MW73g3G1SCaaWoSi8VVwc
dlzBkF7eaYgU527p5hDUxiOv1cigmPaM2FXkI+YPS9zLyz3bvk3Jjwc9m807eg8vbwYl+BEwBuQP
fFMvD3sPy7GF2hzruKmkn3FV/YZT9kmqMLiv5MvseaMUX/XzR58MR8a+KFShr2B5Awyh4LtsuC/U
JLpWqJtwXUPxjsNiNa63i0OeY23KrjzA+aVDKM+lCEylqKSPiUxFiz1mScFJG6qOK9FcDJw7fODC
vL1C5SC3XLt2yl33uXedFgvvghVVV+CjxuGuVXzy4fduuWrIGTq5h72kwFW88h4s5tSk5dDlKbzN
15B+U3da9HmLoYmn3iQ9jhsBd6OYgSOz75d2YwCKDobaqWGNcF3Yv0pjdMgTVv3TWW3FeUKDT28d
d8hDY8L7E7TmVGgMten+Au7xHHIyt/sw4e7kx23o82nZGYoyBTRv1wvz7NyRYD/DKyygjj2uFoS8
iBh5Ajmya95A+pAVNFAqBjz45hQIgOqQSyRh7VLv3D1r8N5eFMeKPQ8EDmq7d7TaDYX1dK7KTwUM
bKuEVgXWHOAoTNwWQnfSWBNKayjdqUPdfIkGS2HDLAWrdE1MPhDfJkRo5t+pyUkLeItn/r/FrzX/
r9upQ90V4rEJGCpi2/mrortEqdXbLWI6j2VAVS5s0EAcP2XJrO5SdpRft60Bh1aVV0iBUtkl/+lj
bwKefyjynkBchCys0NeSu3XZA8tpCTJowWVO7bJgtcrc2/kePqEgA3RLDIDwig6TcJiAvkylxN7Z
0u13rICtOpEtTWkJjWfPbZsBzKmtf3Nuji6CaGByKB9WzCWxZyg7OR3WSeIXcMXEzGyZ/VmcK3nG
/acRIF1xaTc1OJ74bOAkyxW5sPbDql5k7TI5630wBbnsVXZmZl7XkuGkRi1m+A2QsQHaheDNkR99
kks2OwufGezZQ56Pqy3t2WkCxbE77bjNNTF9RTYNTf/mfAmcGxbYEMW9HgK6vifU6EQLMzeBERm6
910jzsM3qobxM7poHKajYq08cTG4/kFZJAlT0Mp8mLE5C9t6LO8l4+85dkn1kZj3fzjquxMIGqC0
Gm2BDE3AwpUky5EMTxywfUs1F8ZKJk++9Q6yE8a2R1zdr+XmR45DcypRBpGqIfoDUzLuy02wzgvk
8MbdBaNl/iLfKR8Z0MwnO+PlWdFF9nAHAI88QZPVZEQlJUYWrpsvqeuZtdOx6B67fmhNo6tSIczE
NmhmgMgSRNCwR1X7PeF636esbBgutn++BtooyHXEP7eyK4BjzrmbxMenw9ElfjDtfv8Uk+vY032W
wS01D6Ke8qpG7kRqaDwfUQxQoQKXhzeuyVBD+0GOJ1tFx6SbfwbjL/hLAfM74DoAWrqB7QABZyYa
GG6IVRjtqCJd2doF5xs3fAEEPyNiDHv9AvcRAeqzNitYx+cVjk870PBdkPtlFbWWbW0ftu26sVm0
TWVNhuWsM+ZSadSy1BuKigGBrcjASOxChdJCGHsiR6LBLtSUfTjjl+4/6Cqy/htVcFI02zWDC5W4
uiJ6HTHFio7g14Y3yhx9RdC/LI1Qolz2Uaqum4gNQi4goPJYcNGgcaVqDaslqGzGRHaLIQ0RNLbL
q0CcOTu9Y0n+DgTKqycJ8AuB0r83tjF8kAnLcIOsxuDmhpolUHNEZzqxkTj6CNgsGdi2Ii7zZkAb
1R8Fs0DYlIS/Yl6nWl3xoxsFilHuNbjqzzD1sw1PeBGWQkDCIHewhCo8L5NAucuVn3wZAuIfYFhm
0ve+UFq4Fqf/was+jc0q1VjmOUOl0JsXstGUUzlpf/No+Tk1epz1grDRh4dylZRZE/7KTyrASmD6
HCWbQ+treszeJ02bv/doVzez8wOHSxBnCYGxxEjdZhSMiUq/MkzNUmVDwNWceQ5Zd/3MkxvgEO6z
T0VlzDH21ARPU3Ig8Ox7dC95rTCnY6qo2sPaKtD4rxyHmRAEmsCqxDxGYie12N1En0Eg3ikRGcTE
TJbzfC/4JpaJmcqnuUzsx3lB2VNyM3COAyYakLoaf1AGw3C1y0mrmuWlv3Zvlp9UCGaCR7+02hua
dNBbi8s5OkBhWAEdK2RPt1HXB48C2XRkSaNiCHmdIIg0S/X1GYNEsTizoQxx7qBIlt7ryhDASVtd
eOBY6ABVL04YqWzQCZ41WfkdRxU9NrmYCHJ3tFT/zNgyZNQNfgQdKvgkpddf1nOnnQMj8GcwaHNW
tC2Vv6sVqvI2soSZGtoL9QArG0CQl1E6gYPaTT7oMPN9a/cOxMsa7mSyQ3bl7j2+0JI0QzPFD3Ay
L1PAEclKYXqxjGYoAmBaP/I1WsuR4lfwjfQumD5oaUm2le7dzS+qQX3ZOaKrhgF5UTOYYhOq9X5k
KvV24PaGPnczC6vSxUOE99GB1WYTwCl6OCLZtHI6XJz06yY3+ncRn3JWuBk4ybEyR2jChnmDtGIZ
N2GLPrsBCvM/pC/zLtrFD5v0s6DYtxJj9UBFI05fjd1JKQv+PdgY9PuT28l6ClWCutIvZ0O+tStF
YSkz+cCBWpt6T+HgyFQ444aE24gLwQApeo2m4TboQ/iu6bXQg7SbFrQwRqJ5Ra+qFTzZD7CjOCeb
l9VKMRcEZiLv+V4IY3AOSoUL28iauebZjJSqCiU99sz+H/GYmkm8KsrJhmmuAmCY436IqJ4QmCJc
tzL6lVouC9defknq/EQKjIB7T2oacBGtYtMpfMGBttt6pJ0fdymcq79db2tPZgAh2fCGnlBuaLJ/
XGrjrDs0+IDZuE1PJtgIfZnPpgSM8p1gvk57Bb3ugvC7i9bl1lpsjGxJX8f68Z6Ivp5dbO0KfW/j
yzGo/XPMTvunkVoYEoc7BLZwTyTTT92nZXtTw2N4Sjkc/jiIgxxgYtsRgzxTf7v4bMl4/rSJP3UU
hIwSLNoIz9eHxa9PdjeF+vwgF7qEIDutK/LLB4ced4XYLcHpdNXwFU+2PIz98g68vUm3Q9mOPO5S
fZvhx9Vv8eDSZZwHeJEVRTC8WE8OUTWvUw/AaMgWOPMcAovzUpvEcrTlkMXtLRFzcihD/qIWTKoa
jAlDx8Xbad6m/9f2mryi2EUC+OKAcNZkQTjPpVvrKqPpuujtTNSBAAAa2DyfC63i+VVZeJTwySSQ
yKgjurMZQpZOyRn/q8c689RPx6lyA1N42lh2UcDwZg+/2yE06P1ctszQ4SZqW+Tdz5/D6dzwtd7s
KAHSz7s1xWUjY/Ad+BZFqG2APPLRls9aqYemnmWjdtvJT3HfiVmVD/kULMB0Gv+3MSeeFdGCQ6jZ
iATT1H4Xdgc2DA4tg8oVIsypsdgQSZdH4TpSIJ1gK4SDD3uCX+3+fmoQjavzh3asXRrc3wuXKUf+
VX34Np79+i+sOoh7qzelZuE32WxMSkALt9C6H8lGoSe3R9SsfwwmEPAqZl/61/5890mN7i1IkjXs
0MU9US3AaxdBPFtU9jNgmO63766HzpgHm+pZahymGGbQfdHN8OppJpj++2EDQl/5nzWnuHp7i9Jj
9lnrbfhHF/9OozD9BkCVJ2UCaIfYWMUFTHdcndD5lt2UD8hpJrpxs9k9SBiRCTbVR3/vFps038zx
qg4YMnsk6uaHBSWYcIaZNYzd/R/ChT3opEW0gxiPR0p7YkdKgPTXBBvY+LILgvxRyR7ZMrFLDL4n
sNPS1AK37pmuiheLHpF/8GfLLqsAxC7kWPqtL2D0vkafZYNDzthH5UL/Ar/SK5Fh/9wLqFmWHMxG
LiK8XIfBqRzUyRHFh3Z6WQz3Unrg6RJ3IV63WUu2EPWKe23L9p4Cy4aydDjoZN4XNlnNzv/EmLVB
b0XZRNpA8ji40QP0xrINVMzaIsXsoYljg8TdVLKfxknmARs1VgMrA4TTOJRSZa8Wvap4hoJ6T2To
fGsQH4b2tHUqBZHbvgHd1loGYQMkPS7GQxlnDHxJPTx71Nd6A+0Nnvl5dln86kCCcBTbjhY4FSX9
b5SzQmZyKCvz9pTj2oEthFjMTBIFgLVhobSeQSDtLr8AkWNrytrpFVd49kPfFEQleLtWCAjxzNxp
M8VGjOrx5uv0GfCAJx0pdeD9bAd8jWe3E4o4WCEaDkqKiBCwXk4Vs2KeY7dE98e6JhGVEYp8a8PS
wGJ1wliVcIsWoOzZ7/WdwN32y9687CcTvLeNcPf44FBVSqow5PgJXI+LWdQcutjcQjE6HcwCEddF
oeSLYrnnjMKY5K1dAptJ4UD2QWBJp6SmKYk303wjQBpk225/mrmDMi/mLio8RdcxZdrp1YOTkuKm
Ste/BpVx9/BlXdzQNulrCTrUTJvfv1ZnKtuFosUE3vRSIapvHwoJ7+Jx0/LrcrUA87Ap8ufwSKxm
RIeUtoIQBaQSPkQXy4s8cNHbGWc7iRWPL6QbFvA3CfaOhXbUf8yZFXQqTP5PW14NarOoP6vI0DoL
vdSHcAB17ipl8nSXqfrdXdx/0yQ/PvBF6BnTdm0aN8utR4QSnmTsxm+oulCKPf++rjX9DWTvT9MK
Ak3JmKl9m4NviNUVzqQYI8FIBsu0LGXuo6N4lLUOzK2bi/Pe1ckbx9htJBhHFX2YBPmd72khWBHJ
mBrrbFyBAwlfW8IfibUgUy1GIij8gOBnALMEX+8GxDeT2uT6RqmyfbNhiyqX/CFd1j0WaogUBhAb
u9BB4o3qvTPX2vLQZ4hr744+eQuFmfG43v2Y7aj3N5L1A6KVXW3dY+pRrXCZYktEJF1PjoA5MHQb
uIqeJ3kgnwzdxiRTtk/hAyXY3SFhaGHyTyR8Ww6Hc0VHt3HDtynM0OsQa3OLMgifILdUwgRHV8ub
v6rUZjyxtZ2Uql1JcDXV/GyoBQmT0NSdi9003wGN45gnxC/YmTGL476uMJYdnz3u5EcBa1sH7uSp
QOIUDQiKjNPb6Yoy5ihkoMzE4P11ISIFoW69TZ21DqFfBoxrUkfGaEwWycgon5eROE8gCecCK8l6
2sDTZKSJyuXA98Z8GvnHQ/6TzVlnCzbKykfBLCHrZBAiMPAQqxzN6ruZJYtgTx17EJqINXwoLaI6
XEPDFJ13Fyrgp5t5jWRh0Ad8CHhnuNXJERu7lyprb0r21hogQGfy8mF4dOp3w2MOCAUVZPxVGIIm
QOEs6uczp8EEB19LrF9rxWusri89GLKcuXAy364EWZjB10B5YB7LEb4Xepz8xJR3aN5xozOHrfHo
CrMLN4T+XT7c2DOfj3j0bGKO4fyDJecyTix8/5IMevZGTRM354E9aaIuIqWTA0/6w6YG6yuyZTL6
eAOVqb+C5k1nF7GQjvDy9ZtcYKDiIVLyPyRBcRmC/Se2+W6/f+I1waR4TFaZl2eHO0zw9RYfrto3
WNakjawjzZ6gJHGh8gLwDLytnO9xymqRPC+gvLmPN5nJd17+63bawy8e/qVGd40Y9wf/wWPMS1NP
ALPoTUPQt5zA+4YpbhCCfxdfKmo/iAc63MLVl5mKvDpO3mDwDVaiyo5r4dUhGVRJ4KQQfCyU/1wL
ywuRF1GyaXE7nVIJn/UhOTRULJrRERX8wEGW5Bc7tbHzjCyTpxgHzEA+dQv09cZbSbKpfQRSnfuQ
5Hud5eifoL2AUR5vDMsWjMlKBvHl2tmziP3XyaERHQukq7VJU69OBZm5cmDY6FtMey00nUjMS4mf
wxY/re4uVGeeSprrmbHqo3noptOyk1p/fh0myoS92zrnIbpuG0x++3Mx0fKFybmgKXZa3h9/T3D5
igLjaPxabNbimESQ1G2fOY6ZXe/AoDHVHnk/5x50qgLKRUlHQ4IJln1SLQzb2R+UBX60iOxg86yl
1or6ECHQUGl7da2Me48tn1+pYE+2oqgzh8OU09VyFSRO3bLphi673UcVnCuge2LQh8tz15/43SRd
emtrhNRvAQVnvByGJ79W9EnmC8ToiVbOlYni278YCaJU/ZMOMXh13O56uXTl/chwx62mLQyF7EId
JXFKmHRBBX85WdOBBWg8uJsglPCPOLYb+n0ibHohVZ9vC3fAG4kr5ed4Ew6Ouqijzmh5SxwVvqkd
oAvc3zIfaTv95vSV9he51lrGcDBmMzLH2bvCoSNaOJAksS3M+GBI9P5tnpYVS0aqxqECqwtGbrzF
T8MotVTrAJcqN0PrH/JtZd9qrrpEdf+eAhVme6bD+k0kKvYiRzUaPDdiVoOyf3sAT2huOUnAXUIJ
odCrzve29lBQ7ETw8b6QsQdTwj9SmWcF0w5ck1F0j6OVW91ZLe0PdyYo8IWXt8NqbmEk9tTWv3AQ
q9cnI4ahvb+x6dYOhTCCBYdql+OPYDUDnl8Yd6qv3RRhjKHDXziDezuHBsUryBeoYG1sdvh1s6oe
fr85orGx4CucgKNG9WwuSuHXhGkRPjf5jFFReos9QYwEken6jr+w7ndSNKqRroW3lE0Q8PUyJjrV
mOJc6ERiFSJnzR8T5MM3jw5YrBc9Zq9pq9tDAAXoVKeCMaF7l1VQcQvhRyBAf+6EP60SabM5J9RE
h2WNMOHySJLeDSVCDWh3AAtwgjS8GGQ1dkpT6bPmacMoCxqYUniFtXjnIkA92YwlaW/tg6pm4ysC
mlFAJ1S9/NGFOhQT4mk3ZK9nWiUGjKIElqx+pgO397YiWs+DdH4MXLu8CrrjosjxGKoUJwUB3G+T
JyjBIpn7CFLaXc9OFgjB1Z1PJELy/TvBfeeOis7fnMa89TrSb5FyLO1JSuZJdiD/xU3LC4Is06os
/pWJln4EpYORBO7yjIR6hVPzaNw5XPlSgF5/05fW4Z+NQ7rodngmlD5QVZF6T/LtvZ3O3CrsdOMS
rpoU6f1wRHVsEK9y80jt0/b6D7ADdw2YysgVOC7yEzxkXYG+a/Ybagircv2uCVHkCbd2To4Ab+/D
EgESdwFVSytCEgPgxGeckPhSdq+XCBKPom/5iQpS9nSujrh6BBf72LVXYsr4DTAAMnNnhUK1XEDS
Apqn7Zs6b8thwERIGkeV5nR+q2I3PBsCGghtjxJIKzpxtbrZWquSzG/erwkoNXlCstb8oC9iNRxw
Nt1QpR90hdu/JHwEFm7uiRJe/TiDmCUor+a0LYJAVZwY0C9JTtOFtc6QlXqfm77S9FvZ/MvAaBOA
OypdUpFELxxU8oTrDTd9n1H5PelCX8v0wn9gzs/sKT76BzdSLQIyr2p1d14+19obCQWsb4Oh1tqk
2V8qhR6IaqGyWG1+LO4hmkLwOM4AgzEGqnenHCIEqdOniJDhYonW0k+SP0cASiET0B8IyWu0rvRY
Q6mqwYBbkNtLotj+jHmcFAZDywktt+VTDbdj/8LwuOsg2NqsrgsIXKGCXrTD3yPqbumL0Zssle1V
ZMZrawS/v385vn+h3NsHqJo54vS2NnD+iT2whzXwGx9nVvKAKnd1s716qXg4j6Ck+nsWUUVZK/Mc
Cpmajri594dqA/qRyjND/etOd+eui5uoD9qlKoxDevgN1MypvE6oITq2JhHSBH8TZffK7gFL/bkf
IyG7B2/aV9J/koIVi7rtrovE6Ck/DvH2toJEpa+fCgpQc4c2spdIBG76a+D8binzYHetoepKOB0+
gG55JdQOeuMYsiuKOxD4Gk/F+q0txzZxHF5+vDOEqAGr8kRbmspi0/QvznVUUmGGi8TLsTQKgdV6
SvG2njoI/+pYp8mE0vSA/iDRtxrl91s12sgbuM24y+NLZ2FU4R4/nPOspQ+UJ7eozFAtw113HIw2
KNU/TNA1HUNLZKb+/DylzIFqEaOaHQ9cPd9dRoEwKWnGtA2NC7V7jqxS6zAlDgdc+s5okPJrpIRN
e9jTQHb2s4NyzPWnmpubGou3XO0CTI4Xux+CQN/fVGHt3Fa7m1uDxR6ABLaV8XTo6dPBhKfKOswX
0aFSaZ9bLg+cLbfH5A5fhzJ0NiAtkN0Zx5cjCJovSP+AUdfUaXanvOjY/YLCiaKzEeMbmSz+SMYE
60Lh+vF8j6munuC+m/B3eyPeZhi20zXW4Hes8jdsjAVuLf6uZyNHkKqqI2hU61gg/kr11Zkzs+6z
k3hnbRaCumswH/xTz+IHHbAEE6WkuUWnzg7s65skTE+GuP2ZwqLhWUBJGqFobWGkjaUHNh8GMuwD
CDA9YBKRTx01NTi9CtYUlU/oKazCtqOlEYBGygR1fY2EMygtWGbx/8dbr3Ojnn8JIXEW1Dhyu222
ma7sgF8Kch4tXebUn0MgFFd2LnN+Z8m8uJEn6mLkgwyCIJQyO7gA3OchKrgWunB6fBw4TRws1g6Y
T6ItOwi+blTEC/fVxWvi5TwPY5peRtt0NgnqjV+lKxMzUsefRXX6sIhNYL6whR3o55ahrTiKKUtY
iIrvkm05AcRuFmVw4LNSfhJLaeSWNnTtBd0Mfyk7gKpdOz5Bhqs2bh4Ih4HXM56mBo9Htx629yaT
R6YcO8ZA8ykoIVgHaqDmb9vdN/Q8LoOqGGsmzhDckSFWDY85P32qDhLaFNHyxYUyS4GMzeixzt/I
Ys42DlaYFZRdsPoK7DvCyToQu/88j30VjZrBU5dR6Kx7uABTewhgyOy1Fb27SSlZfbWcwpMhPIqc
3sobbMojrtNTX2JfF9wysPFXNWJQ6yUFYspLprNu5CLurWf87ETEDS96se9OxRgzOOzN5gN6HpN7
WtdhuwjyS9iS7hRPep5q9Z/M++OxYWmFlHKoHMQQYwQmqFkRB2fB2ilxAzBLP+oy5OU0AMQ4I4kt
c4mwsnle74TzYbnCRfV8MgWYpSMCVLQ8uRWIfaaANmcmuQ6ibMdNJtKoZHa/wIDB74Gkk5gMfDIe
5n7Y+DqPbP+mmNfnwrT5sGV0lQywssnk9yoqEz7EyObesbv/lhNWI6ZuYRi33zkRqO1M0138jkP4
GsPI7gAn3JG20lbqKVyumVNvtmfHlw8QyITV5dQEF+C+uwpI3VLY8FaKxND9AMiUDZVeX2wfLBEM
YO1AfM6mWj7UGuVVsb0fXmQVOpbJADc5EJuyWlgl4dsJj3aIBbuF50Vh0e92/PJhdylET+bNDCNC
YPeP9+ObMmWMSqgswiyiuFQkH55e+yMuFPgDpUh/Q+AiLYDd6i3pYXphp2Mwp2yhiphkDbdbNyD+
WucYdX47jUrwSAN5nzIp7eiJEPwa62dKjdYi+nH8ZecS752Usv1mXaMT5ZwczrB08f+Sfbj/MGzV
egZeZwxNEiFcPY9jb78JCd2S7cVi9RdtWS+/Dho+W7ffKV59hbbgahviwXnN07l0+19g+lGbVt2i
mxQa9pTmFuo+K7Jl7ZF0QWyF5XWwKgF+u0N5txgZECELQ/9ZWreKfbUlZ9nWSmcDIOrcrFiwU0NH
Al5mFqXCtLe5GJO3+7E2/Bgboy8enwXqoDjCV+OqVrkX0leTyYYTwrpeKDl5RVfYoWNz9RvMHcaE
txp7D+hzSBSeEWW06hUpztNaLVCurNpy1z5ygVaHmoYM/JEGOsNe82WBXsgjbqrEvOfthVXrT6cY
iVqyWS0lGmohrWW6NrXyk3PmSpxpz2Mp+9yTRmmmohOOcoiaK3av/UhVim6Ou+eQEHfXegFDaP6r
EjTtv4fXt3g843FPC2tAJmNx/MQAyUFx02qRfC3hX+AjRsqpMGUQC+AWXJMVce0ghwMHYkyBOxWh
mc5OQz1mx76V9RWFM5ATPLnhKeQqYfLTyP+QTFN5VsPzPB7NwanY/MxRYHP3+4X5yEkpyzZa76rL
/dCINon5PTmKdlX3VyHLjRa5ygAq0Hy1kjUcVluTGHYcnmY3sRPhi/Ar4FaNKcUS4qY7JHz3565o
AuIiKZgZACY+dofxSjOs8NSMXJq/orkabVhwo9+dtGD6NrodIhgErz39fesugNC5MbwDM+wX44yT
SjtCdcKlCaqCHeHhe6NKDmKD3T4XdYBjAUASo75gpK5hMPmRq5yVMcvTyVr5fXA2idYojC/9iDsM
xFVsWHtCGDMRXsfgHOhvWw6agEndcrfPPc/2I9ylT2d21ZqK75+jujNIvhBkOjhyfbG/HHZWj0qW
W2D+cpin4jVOdImvhn+ly+5dAaSmBi6KiGngYtPIaNQVDGqn8dpojBRH65a4Ggk7PjOqhy4F4yKg
FZD6dn6lZfeIFZH12QbXaFrcbk55wZx0UCSgqoykQ38eftTT7j1rrW70c/msU/uORGGk0eVMBYhI
KbadWnMuFlw2Vf2Fb2iPEMRihYzWJcLTTvQ5TrI1FdQI7NM8pGkhGyVR5vac1Btoe4lbFtehVoui
6bcDHnCScULBGoHjJd1UEFcVBrwju1RHGDrJiGmn0uUYCDT9EgdFu5aWTOp9dyTF8CVzmuCZq9Ey
OfmWk6i+hPlbSYgVOke8wd9CgTp3S6CXNqqxjDcGpQm7IBbu+A1lkdeF1YJVbK93BfLZWCPn0+aZ
VRlF/zYt4Xdo1/x/CjnhPb6nWEnw3uqvcTv5ObOPWyHbedyorPFpuOiDv3Joepjui5C3VZ2mK2wz
CtOxYu48qs5VmAMozdk099WH1HJ0PBEp+Np+/5eOP8j8ciUmsr07DKMnXQO+2ACk2jUcbWkryvA2
auafdoVWE1SLWDY8+IuBRuQMLH1+UbTBOYl2yTA973aR7ipOL9oTq7sZ0gR7PN8BLEHTNMzKL8Fc
BeiXl0x3zMFxzyY3vYRQrPppoVvwL5HtW7oysePVdZQiKTDtXdh6/i3G7psnQHj9z+mKGMrL6wLt
zwSFj/pKPKeAd3BB07Fk2DlWKdEoaQgk8fUfFjShBziN5zXtViM/kWIOpTGigLQBV0LmdhpxgJbv
xXcDdX48bGXD+bOVs/6wNApx9432TR84+ktfnEg7JKfbsOLGFAv3y1qyqzI4R1ERHghf40wt6N+Q
ln6C4ogbg0LQFXym8/PjVSD2hQYWzmdWAxcwYWLkrTYm01pb5vcy0bWtv64jH2UjK+SzGMwXZ+dQ
zjj2SSMnePyjlgYqBCulq+BRUjgV78MDgb98lILQPPAjppd481iG+94SqyhBUYXKYu2cGiWdgF7v
WlYYiCc20SvWiLzlGMdlxsgYIUacrN66wRFqm+x/7hA8S/x08HnL88i87mQEWAijmkS3Kbnuw13w
xncHXXsnNwfiJmD2Rt2OMA2h2zFO+fZ2JwVJnlMIVLBbahni0SQBvgtMNACX1nVBnjyDfvdhg1SF
WEdNj9la345Qa4XXpHzOfQLtFz/+0Kxcfpk49h0PHLwnf1f/6iMCyrfj879qRxSjAZ3bXCKzNRv9
Hxp9GJwVvUAnevDygbQMDaaDhV54130GENQF5ss3aDAKPa/mYYmbqZrCJUHGf/xCRjupjlrVnhbY
QhX0uiTt3f9F84/a8yt7xazezr3y8CKcAmDWqv+qMli4s8PFQxBlHnf7nkupqFfAG1Xh/iUzNlx5
GveHsim8VIRAHj+YQiv+3+Smtifc54K5qDZhPqqjcaJi52a6KDrMGVeCWyA3xV7VafBisLCd5UbB
Ls0mWJfwNsaIWC3KrMS/f3feR/stTDxAV0N8J7CVk9FE10dM2tyonWzjH0eeVpcjfrAwTGcyUL7g
k6HpOp6aWQeOBYLs/GRVutc1TaZViupjZ8sEZUTAkBLltPeMXmk09IJ64n+7WPBykCOjnF+sA3jL
SPZ5nYj+RDq8+wTsAxMAZbyF2S0sT7OH/bdWFba165VFnHSQNZbTZ2Ei/8raI6qwWH4XVkBgA6A0
gEf37zi9AR4Ixd7ATQNMo6hFVpUy52ugQQtwz0OV8GMB8u78381xfCocCkrHF1DDiSrB1XOb97Cv
07GpEHVB55p5jcWej1kTDmFAw3x1Wa6/yMWKbu9zVp6zq4GPP3KdWS/HxEGhesGotwKO282VnmIW
eZegOd2kreWKxtMq7IvqtC0cjrK/YGvy5TbGrrZxxzk/C5T+OV2ohNvEyQ4YFsqneDig8Dr6UW+u
L9f9I3fcvptDzAfwY61zM6o/cqQ8uWeOiWWQkcMfra33hG78qzbc37zKp5G1Vou89l/oBRFfcZzF
hXD05RFwnPnxJEkzXwKqZGYvXTBT/SMheG+0kt4Bbnlb8aXMHvED2WCWRBnejruqXRnK9UjK3/VB
ab7X9rI6TDAByYcrY79Bq7YpgXBH+BHqncAQiafO2SaOvaG80BGibxOORJtvf4Be5DzY5h/wyOx/
AGAmofoT4J6nFnEneHSDzT/hdTJExqIGMbkasm+iOabcGxOQ3t12qYCFhGgFS3CkRoOstyySv/IL
R8nKvJDNeJ85Tg9lESQ45zrp9n8a1qiLv2VOHardpmgUXQR8skXR838sVj1OCMacMxV92K9zAur0
70WEpYCyfcmeZhTcbRBrNbxFMTsNzY9DvV99zty975IKcu40pF3R6wh7ZB6ObbrRnyRQTpGno76I
bkyZ0XRH9KyFFpSBgRLnTwORzRVt/j/8Klud32smRsFEyUvWYpfDZewsEDcc7Fn9ZwhITxNVc50b
m0U24/vR4di5FJmiJDvj+2n8rY61TslL+pOcvzibEaITx6jS0+ia8yc/wWgarE8YeptzF7/NFYZM
kvcB26MS/dLiq8HQastgLnEiIePdpY9FtC/TwsgiheejIU5xS+/kt86ALP8wPIQrnpsWc1QkSX9b
Puht7URmOqDlbu8N+8985nwuINFwV36taLgSeiCcDRhtQkqr7Ictm4p2X/jWEDYCTPEU0Y0+imUo
/bdSmQHpCW1AU8ETF1KtKIpra9zuqyb5hSi0jD7RHMkRn7BS6/mrzHUagXYVSJvIw+6lj7rupL48
by5CNPS6o8lk3A/uaMc1a6uV6LlPczHuLHHrR1GvI4L+aboEC2GhNM1mEbC45FsnesPoFXqEX2KJ
fXhwfV0ozUdEUH1ZiccAC31gUYQf1Y9xMySyvkXOSzELA2a6uJgEz9K5cStqCrG/3CWHJzo+D/wu
7S+nGS6BWPI1s8Blly+WUK8GHiOyc/yYK+0yZe9Eo+dTCzzx9dzM3eFic3Bav8O5b/QZa0S4RRnN
1et6ujIghmN7ZI5PcatLxJnI/nrAuEGO9XwyJUSJunKTlrwOeScMVDBlxbwHLwJMTSJtcGgZp/i1
1ZjZssvsG7ge98tG/XEGiwSGvaWERA0+F4fWj/HjrAHxTlcGcmN/UPLe+CN5ZHrR/vL76zUvflM7
sNRKU5ZQ0kUd8SBhcXh5T2xVYryzUikl74t59PbO2FPBXrNThEJcEt6AFcZCLug2W5lELk7UglHN
bo32+TqV6PfsMCbatXc+irCiFqYUR833lvTY7ApJifFd0+BOqEKcOyVFPTBGs8L1NbdApH6uh4lN
t7adnB9+1a8HR1g4mSD0RJtlwVT73EcDQDzcBeGtMfC0VJcXSrwVsO5o7St0K0gYG3NGBnRNEqk6
X2y3Edx8nf/60WKSMqdRh1ojbLmC/SzlFrAgUBmeYkDnEuK0ztvlvuc1hm+oUwayT8qZnBCm5MrP
XrbyeM73b2xH1RwEfDInYLYNUBQTo6RlXi+mhcBhMRVcu5dKEsdyq4VkDtqJQmoAsZohN/VYty2A
sAd6aWJGAeXiE5DiD12gDSAJMOyf0IeF86ia4jVBLVdM5NIFcx346cgnUPmRamYaWQ6yMqjunfl2
emZyYYimBmiRqToG7m50DpqYw3R6ZXnsycYf1yyTnO6XEghORtcYWKuwxIr+nNOGsFkKc4y9/uS8
/O7OznBLSo+C/oMWVU22GANDsmTFvqeJgiGYPl8eYHptWBXra4YCd2j/ugFlUH3CJ6F0PWJ+y5l3
J9m4jONzuSrD+F+9JHzs2uSLyCUWZPhSZOKZ9AukbDE142YLe9UTQbeznUI9mUKeUI4GzvPtINbC
Ul7NDZkQAq+PsoOOtzWIEQWUoAN/MQ720rTV732pRtCoUW4xsGdTdV1Ws7NITCB79n+fIqq8Xfed
Q4wcwcUUq1aQ0Vt5dbopEYNbPWlpvgR9rXvOktYZAa3Fc70K6sIBtp7tMDBRNsHT5TgFbRwu/tDN
ZBuhxx2aUEQP1HNXVgqvgGgJzcKIgCG9oWKVz4DIca1JlrKZIMasiU9qRzEjQUgNO9NJ08bZfe+u
Hj/6KwO3jSyTIRsQN5tlQ3p8fFlhqILcPJNjQbtF3MroRI0XHUgx/K/IYlpkXpZUx+s8Z6wa4xcK
oSzfIUc4sgkUwBmFmncFspjffu5fl5dCEqsXEwaFyFsfJwZNGgs6ulL/Ou90+yaRAoxRygHLXIjK
tf124YVSSRs5d2zU9ptIDwV1R8747WH7lvPH9MYAtYxUqpijL81PPfB0JvCM7WZ+nynxq/Wu0ybB
R3EhXyXX8W22HTB9PcytuOEWYL4KAYTuXNH0meMlV60mvpIyzzMM7Swy8X/I7Av5oCftKghxnpcD
8aya/+poPq596qPOvQd4b/AJBNLDaTZIp3NT8DvtH3pAj0hGOxFPs5QzsZ7CncNkYHlZ2Jx1gArd
QRg6FRM7lze1zWJFOLpj2LQwL4JZBlLPqx4PyVX1xog1baCXYdYnA2p3iGGVIdxtaXeexsr4bzzW
pqGP5lxdfqerzIW4ucUFQK6XErHxgImhT20WZreqbaq54JRL/Ph3l9urapH1mbuSjuj3Mrl520qU
fu29PZhw+dh/5SNBjjwXco9PL2BTDHCwJ1nu9qE06Sp44PimJpS7qA5sEJzqAzn/J4rug8HVHba7
x840lU/AU1d3s2XTKrbbY5f+Nd0alZzKWuJ8hNpfvBSSr8/l/7qAqjSoiPnqVOVDuc1VeGe/HQrc
xecdMsmj5XtbdDadAUnV7ayNP3aV/CrGt+jsx7XCwhBqe5vcAYRXBjS45+cPWQdnCqJ1R0afuOvr
9FUyiN56Ym/ZwGTcxmL22qAy+L649UzgdDoJ+/vZDEIhYh8dRdoX3GezPrZhqyKkOABfSDMELbVf
0ss6JHVeLX77Dgl5EJIfABYf0avvpZRb5gMKaIF62WMLp0sSDDgIkQGnbJ2SXq2NJgoz9KOf1kdM
gX+9I7EqVgt7mmTIUaC6nXiSyPRkCG6aCkufGtJqRCWacnocL2aEFRPNcxLKldarGGuWPCPvLDFb
izatt5itsXC2LX7yK2bFUFPICoSe0HC5ZvHrjkAOJ6l9MUI3EqCRl31uY4bTEp3bJaJ8iOCuXYyi
AFxgNSN9K3AaoVWpG+R+MtZTgU/aTizKlbQ4ZWbqkFeb+HudzPIpjstyf6IK4dHIr7pV5zEtCYF/
2Sxwezts7fIGSxnK6iPDppQynSvh/6t5+kx44M0Nm69LCEGB4OlvDI0nYgUQ8kzcn0YwoYLewi1l
y5msOLUi6Qw3pNlxy/8o5hkMknMLHNHiWffadFsIOlCPu3eG8vVvjScRjkTNSQ6tLCW/N0Rm++SC
LJJRWp18Dq+G4qIXcuAcEdnOb/YghRBQkm5WqJl8CW7CJhxAZ5PIl5WODT9ADaiP3PyH0A95JlAj
WW+WGUHTl0CjBT94YbztgtgOyQ9xgviYVnrTao3nZfEoCwIa54NOnPsv9iRcOPtbNDt/LFB2QvrS
AIxiig8A4QV2Mmo8eLX5hUAevI2pTAGKiHOkbJa9mPwFSNpkPrXoykdr1FZHi1S628Jk3TZt3ETp
G5uRMC+z98X43rm1T6JxN2XxENpEaa4n9HcpZ1SsHRIzvCSM1ILOrg/fgGMrrMbDVeYeH8hXVvMH
mi49tliER6zVkcTMPLpz3ZqZlB60QdDpSu2e/TnpXsL3r+ssFjEOWfY44vbbTnx8bj/avW7f2II6
xPLm5pcglrw/bDSUo6Iaee/LNSG8FwVYYf7dt5POwmA7xRVvBVSOHADc6t4IlmQlkcX3OxI+lXdR
IB1WnoDM72sIMKlUbMHIUkoSUZuw2SPIDY+vFvjJBe7/LhuEQq8RhuFeNyCJwfTNjcdphma6uQar
RTAMFN3bFiFdBTnXSCsTDsGnWTOuuoJTISiQ4d07kV0jKPV5k6MxZ1Y/3IdMadqKdpamgIa+ZWyS
HLTkfATCHsbHQ5X36ngQr/9Hsp9rCUt1+6A6js9GMXFzRvxRIYujvl/qOD9Zn7u5pFSGBCnwZZCT
ELYdfb4z/gBx2wq8/wwmLbFdwgU8pnxYFUbqCaDUWNKSlRv1+cR5BALN0kMAL4BY8EcfxoDEofrQ
uqSrZeeHtFjK8QbKSiZXZo/Aa81qd35RCpa+RJ9mtsRRV1Wc9Hqbidyltvr6fEE1pC0C3SRZhC7B
yOhbGqi4OTa9iASv+WoAvZ4AxHOvmw7lDaASDKdRR5d4GKXboCgZlU84E37ZUMQxNgZw8PjDA6QV
tUf3vOajORRqoAvE/z8RPJ6bSpkftk7dfe+cL1JeXqZEjXQDFeIuJK6xOs7KBtrOEqlbutKK/Yk3
rgjzJi6oq4XgjIZJFqLkhnxmiIvkL4KowQKYqGjcuSpqs1tHB8Ot4z9yCSGstoUmfT9wfdoHCIKb
IJkinyRZUfSZK1aXij4c2V+3M9e5UJ0+oH+RCNeJGmdybe2SbSuwbcbxUkqr5sbUW+X7WoBt8jyz
0m7xsBCp1OTmXwcIkWAYALMQQ4Y3rHfTyxGJTdMfWVEDhibXtnCJjYLGZSHkJ6nLu2weDAMkLoeu
3ZmhvsurLMVmpFGuFKy3Khn23u3fQujoLCtzq1XoZwLCih7j27Gw6aZOLSjWA+qM8YsnIzkuO98A
TNGu1E9K3GZ7T5iqdyLsPT6n7aLUR5IC3LPZuT8LP8WsMbUXlDfg/ujVAgzYftqtI78ElAeBjA8p
7CakZxUo20jm/ertzEAWzGHnv6aIxeSY2ATn3BLRfIF+9TFA1lqnCApEG51hadKzlRAW2OmDiZu/
WehmK0NtuvafX9bdW5J36H782YcZQ8RgbcNbf4eBmkY9L9wXGdrTtzpufZRLqcbPcRYdoZ3TYwgX
8uQPWwO10SW9koD0Kpl4npFOvK94xgzdccr4DJIF+PQtQKkqcDt6BVopnsV3+cfStkr0t/ZNynS1
LRfslMcGkGZ61IbW/HoCJQaKlZBnMHWNfL+d4Cq2d3Hln5tC7O//D5LbCVBlBFLqbDHBQ4ZjKzbL
yP9/HfXNxuyxgbX2qvq2gKIriIeiWPyWo+aqRa9q4QIx3BXU5889PqxWPSJ9o05PsbsJ45p6Z3j3
Oupn/dwJL4HD8Gw9Yn56Yyp3iWROapLMA9MX15U4cUHXQ1ypnmyhyTN2JZKVDNDQ9IXh8TyyW1XW
rS4ZbaSxbmCrcC1OCB1TLjoR/7mphCiT+b1e/V8l+G+cBC8kadTTefuW4571HE4dZFNPMORQVupN
OhKnSFSdLwVutKrMndLO5ZzTVYeFdninYijOiQDgJ50AcOEluWqPP/yPdFR26uujx8S/5b+ik8UY
UK0baEC5D0n5c6o++ki6n+owdHqJGUx31Tti0za/qpTz1m2BMNE0+0GUmngjB6wKKDQEBjmyHKVE
Haww68IgCVfY8sp2jwCmrfEqcozfMhCPp1UvyeoxcPaCPTZ66r3IXupOhQ33TlrfDrl47ATw5c0B
/TzD0US7leCssRVGSMjz9BeHj+NegQBKBGN2p4cxbX824oc3EgBFTVk9Y/aMTVUlQ9oF6cduY+Ho
LX2oPvacOJoeITeJizRNTPNaG1K7z0dhFfhpEDFxNAXk6o2UPO1wE/Ufo5zrZ8bSFsDeA775EI39
fFVKn8V8WoWeYPK3CNIB8QrLJ1ymP3aI9REf6/cK6sWyl8zfDXZysL4rWYUvAmgOlzysiGT+HFgn
mBSn2Oj56lqSLTcH7Jx9djfYSsg88hUVB39vC9z0ezSMgIbkz4PgADTr6mZycmU2gYY/WYwmPNmr
mfVBff1OSjtwOrKjyXoQbrQCI8OJSAklT4isZoIGanBwyjuGxn0humIvQpHqGPbpOEBkxWkPym+x
d1WvIrfFjbwJcdUD3ES8Vf+Ifov3Iu3F3Ol9lDLl1yVHoDrcORY5jf+wCaPoa5+wMnA6HzuFlXdb
Et1mwRo1KO2iuQgq73rHj44A9rk5kOPSfszKfELaT8NN9cDJKkvuvNXdOnBrBuPHfME4pubHTaWN
by+EUZpAdz1/SEOuFCXlqSqobliJv39I7JXq1y+9oWb+pj6xGXROaAzaFYjjq+t0j2DqUSLsClKX
+xGiRRUWV7ugwHpB5DGt8rb0+N16PF+LxV/075p8CAgD7GFg5A7PB2DgqTjai/07b/UCAnPRARyq
ICG8mdZBgW7Qn7ptolzBdkBJ+EESCowySAJBcYk1Pwv141mosO4xcHPF5wTkBfnXmPfCjh3zA3JI
AxCC+lOxl7EJW+7/CueEDJy1ENH2cuCzqqWrnrJO/kiK//ra6yYZBOuEhTr5R1mokUjMDbRvJyPU
NGxLgM1a7lcFOxcvLWCoUcg5NPHo+WcZKpu4nhNMbm4X36oMSexZv9k7auVYU8AVDBLunIewNIKA
iGEOHjIWFpv+D+ja/a2RGAkum5OjxJqLdlGAhYJX85LZ1by1OjT2qMA2514O+vhzM0fdCRkfxCcU
bmf2X/WIso3cbESu08dWeZr3zCTFBfjirnlccwLFWsEXYOI48+M0E8XTp4sc1XMWGBIszaxJne+e
Iehbo/scv61yXXSNHmOj4NZXr3JXUps9L63e0v+icn9f6mHqwfDlazMem84AmXY1VzhNi9o3+k4X
OHgLW5PhYk/bqY3hZuZ75gZ2Z3H0/k68OdT90RM9lP7TTMkhxpj8HrWgXjb6k/cLVmlY2BMMOgcv
2Pg1ZX4ySeAp1r9v2VgUuoHIE706QhiTCnCy52I4gs7XQUsxW+IevtqXk+tNF37Q7b747h/LqNzM
ZXNet2oaKXWnMYhvyay/zWpxzgAdhyqPMHpoouqc3Fooc/8zWANdIv5SaXtf+LOzYm/xrKT9ckZ2
hPTZv1aMiSk1e1jOu7hi9Wcmh5UwLier0+U6J5tHdjygwS6QLOsP5fSd56HDX3wutFWud1zs9mBg
fOW4N2DaWZVdBiQgSTIAwK6chKemq6TJN3FEOAcukEqs7jKXuzMgQqEYKrqtSlQKP8cWO3WYxq4/
isg9BW0UgV4E7lVeL1W+Jq7CfZwz2QbPTSacrZ7YDmX3J+p77rAJlzbbinPTTY/e801aWwU5+q2E
WpH4uh7Igo9jz4VzzQ2zQupXryUecBAwZI/ZDbsvK1iO6CVVluGCddsRKI/80L8E5nTe9AnsRKwT
/p28OK9phrQxeovdHjtcBiaSh7X+mpRkRQTuE9DFfwXlRR+uU7F2qHr33x/zPhuVjCNhgQ6Gk9Yq
DgsozpX+uCc1FqvyIvT+Rs2aBlslaRJLvTbANxO1O7T0BA0n8ewDVaO5M38RCnSWBYXJeEh26rQg
p5Lm5tgb7/hY3PJWLLT4LnMGPFQCdmbQK53VZ7adBzs8NGl2B0ArE+vDCXYldUPrvEIYIFQPesvA
kJGI8pCv+X+MtMZcY18QcSFsVnUULTxXuNn7OvxNT06zT9FtQcDEZtNbJyRfW5ki7zqikh5yivoW
pjp6scz5t35yXOZH6uuszxdgpRjkhOZyunmsh6D5nMQAuzFTtAqBjJNaiIpTwjySQMpc9mUEGgtt
7rxrofwtKiAHrK7tm6DWSfgOXGpeeuASe7EtQnSBA601cOvJ4cnbtSqnycvh67lWt4ieEX8cm2PO
btvDxA8SEsJiow0Dz81C7Ch1oLdiSApaAMfLRyprDX6wNRhKTNYAwBnRIJj1iJucLDP7WpcU9m11
jkWtA4J9MYT4aQNaeEps5yYmGLL+gYfWlUOj+wj1GxULcgDtFX2dXv9mciz+7giX+YDd8P2OxVl1
KWeADknsV94mvhTdxxhHVYNRRdXTAAJRmQaOJzyRAxr8PVnZd6A1d8VvHMjo9dlPrOY3Pk0OETli
sUdi4VonLT49YZFrrEDj7Dl49NV2GCXaGAf0IiNOi1uLd2tiOSJnnVlGwXFnbKkXpT6wGb1HzKTx
n8x6PQTTyiVa+hvifTRnA4tpPLYdyTRoyqDQj07p2NK6By3DK4UclIFiffEA8DhrDGH9NsT354cJ
aNSNRvl3RIUi8T5Jpp4pa1a4/NUq18cTwHlQ8UKHvlJK/2Vw4QahvHKv2CxK2+1TcxbFT/wuZMpd
qu2GqtknaFRAiHwd4+EsWISaZSqItSAjl32DBc2dpNcAwWLYxCHXz5JsZXQ+vpDLWzlswJtqM2JC
qjR30r9LOFe4utc4NCV/k+VaDQAhhBqdx8gcnJymJrPYDso6oXyVpiA/ede3R86pvJGN2wEiIp93
MWt44lunLJjDOSv/KE2iJbKy98A0w0/BxTkIi0Af5fvgMl4UeaMTg6riwg41xeT5P2pEmDYL48qR
txkwXboio8ng02EvBSxrKOEsbhJMOw/WTi4dhsZoF9ND+toRfFrLYDGgfH1QVKctAKf8bPVdCeNE
zOlLrdoyrhKmJ3fr8FrMe/SC3ktvALHqxxj4+lGDbFoN6kKoFdufkeD55uk2dJfbU0Nln2HL1WRV
H6ZVkKCtg5ZY0n25iZMKRZwLlJvn6ZwZWs/RNQ5L3Kptx4TpRDH+tUxFtk7WbL1TDK/V68ydkadK
JDe7uuUUq8fR71Q2cwXh+u6HnyJs2XWXmRIt1MKOw0Lnq//bEkqmZiK/EvN17PwabdnuCgXkMVaA
idkCYPVMrUDUVr+SNcJ3op8hfFGGkjdcY6znGqvR88zHvUNc8O8QBAUolkM4+E0MPZ+4ZIPlG2eP
GTYukCYjPRGC7pof7VRBBGg6+T6qntEwxCIwBv3c1suBtg3x8k3/zp87TJGLIta7+dWIqb1RRf5c
Du/9Tfo6XCSdURadYU+lCobE7qev8hdqia7MWHxEnbNdCc2/3zoGA5Pf8fXmtJbQTkYHnvu5TMpH
uYo8AJeCchKqrOo4y1yPLdEHHoiVSj+SEkCzYkvtHFMPElRPg1oXDqfifeYvlieNE46A/sniJ4su
0cY/jgl4MCn4zSPapwhzDFzhdvJB8JlnsKSuski1lSuPfNyYSs/Dzl4hCHJxNY6znLeJIV0os35i
w1AidpFD0Uo9YPprA7/AGoc7XwZUexbte3LAmAjq89xrMhYDIZm6oOO249enxvOjmpnfUVuabd/W
2k6+bSKfXa+ftSbucEqM9FeZ6zA6apkj+DHfhAuhP3qoQg9EC7etCiqN5AhIqePJj4Ubq6Ha8HfE
cRsscprARbzAPMIC8sHNFjpQHaie9N8JVZ3l9FY5UvlnuwLF6WkcnuumcWnNXsxlzpF4fu9K11BB
5gQ71sOhSm+efdBp2YlawKzo2Ch0lVtupaOfmzaYGELkYHOwck9HQbzP3qfvUlKu3jUeqnkS0+n8
6JiPL/gbQnb96A6tHr0TxQ2y7heJV3CrW0xTh1YBTf2ReKfBYmHmee8giqRacLIqqsvE2MMy7cBp
Tzd15Qj7vCCHdP9bQBKU6FHrNI4pAAjnbEGQ33g60sAx3VGOz/qPACesI/pSWUJzilGOBV2QLIo8
YUhSgR1F9ia7UAjv+2t+ktNnuXSM1PaKJbA4LAOh2KYAtqJDFeNHeqeGGUgyIp7Wpk4OKJ8LjXYG
MsBXJ1TlsXWSvF4fb+lxDfQ8c2U/TJWH6R6k1W+aLf9em0rnivJMiC4z8/6TpQfYwbwovmMt2fqA
Acze2E9wC0j5nkitzwHvRgkBlhdWAr7yoE0/zyPS6mSRYOXW48CaJlD9GPsVzno3qmO5dPQJZTGn
Q/xqKJ/JUWn5TWNYOLIb/j0gqNikIFPvGN7KiHuFMU0TU3uwvaoR16e6o9cbLarxG/o2m7i0fSxa
N/FvrLbovnocOZMLpXSWVovyUnOBa5S3JtPUfhbeklNknhu6ltbHB/hRqJqd9135LwpxzXwsK+Yx
XcvgisZ6w0c6zCUO2EwHtY4y2WmqAvEetfjvT3WUk8lmp/PDAkSMaqFjJ2to5uZ13XNp9h3WOXeo
yvcCm6IFdxATxQjvlV5chh42xvbIZ5Z0y2bV0EqAfWJIPrS+cC74dBLnVIanMm9pyEwo3CiewSNz
GIHTe5yNAifmTn0XLaU5GdIRJMfzhjwhzaX3CdZVxM1iFejinDjHFwBZ8sGHf6mhMBLftS+3LC13
gNWaYiOIRfyC9VikDYTCxqeg6YPLmTj6bQDGXtNKh9eTAJOzoPCj7fG2DqMtCsQIU32IeX7FNPOA
kB/hllwk3EY2zoTTlCCZnPeUL4i9ZCN8vrnNIfIbsz4WfgALUYnHNymQY8/x5TtPvBgp1nRf0+Cz
S5iNMwamr669iSyrVr0hFpCQmIXO05s9ASklMmG82pmeHYxZgFOPDyeFOwY4CV0z1jwhZKnmnILX
YAUIbLSwo4WrCjyFmkr4gRfN6ktXMhbcBYzFssvJzorIYKDUyxl8/04qGDh11fWSvr23JwEi6JqF
d58L9waxMh2/KxqewHifaPlSvBSRRUMR4LbqX4owMW01PZsft+d544hBv26QdS32/APr9UThWEtv
+TjdgFDR2NSZq4uM+fK1DIH1/fPnYGneSr9YG3UMVn8Dcuvj11yEQvZWdverLsFDAMj47/1oB+uX
ROVHHqlX0BLghZcq584q2LFw0hGH74htWdtXtjBWn04foFfvtYlVuM5BkR+XZPUW4Epigj/ZeJST
u2X+wYEJnNsSVQAAgW+sytqhukCfRg9mQrw3v6xb7Te3qFU2QH45eYNWS5+luUVxXe+xzs9WACCE
AwKMXabj4o7LdUIAcxUtLEm86YGXI2sBt+gxJmKnEkpAvxB4YAHigmajHQqKMWPSA+Jg3X6Ak6At
kUuM12QqY9KdLBir+GmOr1+7/865+ZYdz9o2b6w1N7VvW1VyGP2U5lNHwBc5D1BSTRRMoHQndrx+
Jt/8J2uBEbPnQA6lFX4gkEqSVqSr1KiYwoafxtjpknYsSBOWxXDGhg+Y3jYhFETji+SUjQUp3+xf
XKEdhdAAuuPAUfN107oBbEw4X6x+dEoP8Pg9ILcUGeQ3IAkj0qE9s9CW7gZox1Mp9B7aBXB6x3cB
5Z2qwh5PWvD95gS7HKlKcp+PhSa+y4AI3G11ngL8kjKTq+YI5Crfulf5XFFKoNEnXSlHW/XEVo74
GNCIks0fzhCvsG1/hnOYqr+d28eHEMX1klCu91SF4W9/89FC4cFIj9uSHQa9kjTlkB6VSGI6swfF
5c/H40Ec4fRlF+Z6ws0h/E8Q0hFlV0uQJxmMI4nS/WDU+Cj3d5l6x9neGZwwZqbRiyeWtJ5k00BC
624qGl8AF6xYA1XzALWGnRocJdaVHvwjSsZc/JyGUPeKKZ/SCy4Ei42k6+lCVSOtdEzh/qSkIG1g
KjgsBg1Jx96MtfVZtXP0EHJFy9K5vCNUutDwL7DtKN5YZIvqrAZfXCvHy6AuBNtJGve4CcqQ9+z9
+VqDVYLe5Y17X4Qt9zW46SvQRK8nXvPnyoGx0goqtLuu/WqM0PkGbnxtctGNO1WiEnguFiJLliqX
2pBN6KTYDgi4GLnMA/B3Wl4jcNgFmbS1ECkcE9nH6JkcqQLTB0HdFKaVv9AUdIct1RWC011EmI+E
rySAWeihRi7G3+XfSMQu8b1RdhChHqw9/MAmf7A8Y2ZmPmNnyAiUmE+3IMzegy2ccUL6L4Snl8IY
d1WCRwsVzlHODDqll5amedqzB88/SJO3uItFvr/wc/Y6LanUJHik/bTK7RvRnznBfiOSZ+KwLLJt
cjh+IQLwElNVqCjMutcoP1B5/C2kZsBDlgrji0CGUDTnV9q9ez4z8PNUezO54VvNOf9gIQW+cwOJ
ld7JLzr/Lg2LhByN7lBdn4PIKXZ+rP4maXBN15wuM5XtJ9Rq9f6ULXgiBa+f8sn0C07fYgQBXZj9
AV7A8OY6Q4TAvjOw+daerZKsyLt4A6WsWW2/tX9auZyEFHWa1FkxDOTJEvYKitUKIjZrrslH3PSg
7rDqMkSQGRZSBn4+BrLziFyXf0ATBbfKZfHJDUtn62lc52wlUIe8aS0p6oh18ANMJfqiLAHehkrp
DS1ampXNqLAOflNMk84KlaZXSx20BncnQgKkd93I83yRTrNVu99ZV2lhcP2gq2Xq6ibmT1nyN7T/
dZWX9q/XNIovfTmR4nXGfQyk2dSAxTOvhMOnZdqokcqux1DLg4LTbliY8Fr1fCmWAyqbPQSP4iuW
n4D1yxatDuzjQ98s91eHNqWjjOsUHTuQV8zUEyds7nCzEUa33Q9O773JuJpNL50I4VNEm2wKHrtB
EGt16a1z1AOfd7b+KeMNvi+ilDCiP/W1s6jY1DfiK11xFRvIcNJskBsYimHIzRX3BRBwhc61cCO8
TGEBFvm74LAW2xciwAnu1IkDGZ/kJVzaB9hNakWvuG5Cy/pINfcyRTADLP/yhpn9ayyedblyg8DN
zWSLbUsBZKpyJd18ubEZhmJlXUK2c9bTa52w3/Kf91JL2RwWse67THcn13TuRn2uU9d886lGqt7H
tU2KieNe/eOzBanDNr3zuDqFTH/efnt/PvzXByIcL+ASkAOhqCld1ND9fz1AR9OevLfF2r/+FByZ
tEnoP7414K9F+PKefL1HwnOK0a1W5wdxmV23fh5+Zak39ERVZpV/2JO0E53BLvG1SCYFqBH+7OCQ
dn6QkUSYr5G/ISaECfRaPbg+YrJ/6It6Ti+OjFNeJ+g1lv97MEPP5okMqa6pLrdUKMK5bGqDTAPN
voqcWKYr7MH9s4TProX3WMXlklQgmCD0l4F83yTa9HEkEC2s5kVn572K4pmsyEMlHi876uMM9xoo
YyDVhQ/UI1Q2IQwnVnr0RbRcvdA9K+SRXsa2AORy7EpFgTA2dBIOPPLwzogtoFicOILeZKcnQFVz
N4KSgLOhEeoU0bDScUj4/mww3rFpqg0Km+8RF7pvuxUXJYVyrwhwc+OmCEXSiG8dDhCghqCjo9eh
QiYo0CBH2LZFcQu7s6w/C3x7ApRUD5cm6CsgRCI+J4AAFtAxYAsVt5qYlVJp/p5KdjcHj/oxcbAB
ZuOAZkg5NCsJCZGZYUwnDWYYppmQJRZfcj4LBTIljTgUmBCksDbnqc2e3bpfgj4opinn9I/T4kcf
zSz9xv8dc3XXvzrf/4/7mYJh5LverfHM7BsUGSlh28HW3SBgKO6gpFb+API7d7OR1ZGwd1abr9MR
TvdihwlXcZs2whPPU7mrP5tgF9fG7k+EsoZUyBOzUWHptoSEEp2YlM+IAF+m1CcxA4DZhRBYvJ8t
XfpkI0W8M/OIwiXrveTKJREb/+k/FOcJyuOhnkKwBhYAsHGwrNdRnwrm0i+oBxd0jl06FmmDWjD+
kOyeXu32sEqVTQdufk0n9LO1/titvtJu6ozycIwVDCPYnceUz2yjS2K2ugpa47jUIoH+AsS0kYXN
E9Mn0V5DCbdpCbMiKZ6VYP+taELUiRX8JM/ONHddEFffsBKpxBsnBTQmOUBpvmCGiIDNuPBUXcEH
3tbrnlBbq6ZTjwSOBHGYkQmR3lK2Kqq7T7kiq+BVwFy5nUl0J8/8RIYGishm9lhXkUgv0GQzKkBw
nS5f/MmsQ7m5UKe1+QOUpz8CpP+rJqFY7qCOg+DNbdUgFt+k+F8yMnzWt5gGN/U8WS1MIeceyt6b
FDF0wVSKi5BjZf4Qig5j6k5NJk3JvqmRazax+ntzORueQx9L1JWcvJ9Ud4Kf43L0EoXeQ8MiR9Xv
lGmJ9Z7a8wYB9u1nDu5Tf2PyzcFswYK+cHKuBseb9mPCEGfefcB4ei7MQ2V+YXmVQb32cQ6A1S+M
y5cbqubbS3bnfS+D9bN/rK7pXkaI9mdUsrgByy64962AT4XRQLEYGZMctx9P/UNHTQ9uzLdIb3hh
ss1e3J/yZhTi4uuRpCkFmaQWGki7FrKOdXXgPU29Ff2FQfnD0YGqrgb/4JI2MV1LAFAmlnpyuKXA
1fxk3T47nyynAeFxxjulsdeuH4k/v80rvsTSAWbjS0wdBuubm1/Jeqo99G7xH/IpsGSJxUycxh/p
dLXA+m97NtRHYd6xxPpDdQvhFgKLWPiddTcOVI8vAzyq5AmjT8shoFeGGEWcYVQ4QedaaA5ekaxW
FUMnLjNEtUk2H6xOEaL9O1WTRCbMe2160rPxXMk5POluapGL6uJ0IqqdvdkUuiQ2qVFkAv3EWksd
0nRH3nHuLzN4TEsIfetyTAjcllEvpJMdQPM3YAi9udnpJSZUB+TvsML5kRym7jSWPlPQsC0qvz15
IvfsRDPPNxrM+C3UAGeBIZWgywYXuI4KBbyZlX8X6qkb1n1pNIDB4fBRDqyEnEHAFZ3Wzm4n1qEN
mwdrjKyvk05SeXZptH2Fwe1vKpASkjIs4RvUcvd2sddw5fvh15rXcynn2lcpsI5llrmT8P+RZG8J
lwI+Ehgxvwxgu3IJdlRD77xuniKZ425wdtfTEJFHMY7WhHd+LoCNzONngv/lpHN7g8Y2mrCa3I2Q
ogBsOWtsLckJOeZqQtcBN1hU345ZDIwvxpENwkgrefT+Rehh8+qGDNwoe5uoLJcP3HAqVayptISX
U0EKaVXvD/UzLGqGa+NTty/ABSFu0zsa6T7IxD/3Dz8rkJTi9MzkLrkO2kNUJ3GLa4PObe0hiLrM
5YDWbk7gG44OCmlGaE/bNSolwcIYUCRlS5s2cFr1MijbMhzl5O7b6MpHzq3nfYloujY9OyckzORi
dVp6FDST32bK+fj4zZxs/XhRjGO5Xjy1maUV8sPvvE/+RCHKbqhV5GzTKIwn/JMIwpdlJU/tfm3H
0OShU1n6DaQNEow+rbEyriG+H0QWLwhg37qelWDNijLJ08+c4btAusfM8jaJbLi3GRbJtyClEaKM
sfk9qUknFtaG37VeYEDFNGnVtFw+lMtvRPqQ01tLq0/hwpfkAwJn3qYg2lg0b7dHFgZHVHH+bdLg
2Tvai6XKQoryyntEBFbzZPIfF/d2Yd/94Tuj0W51wxHmolAHgQ0QMZzn1yd1mxo5k/4mvxezgSul
Mf3r3/AuHNvaIPV/MIiCabvNXd9JlinWVs9/OymGpLNCfdAf0r2hT4DAirJIrChyiceg1kJR/7l7
D0f3lvSZzUn/rojoeAxJn4nIAFmqvuFQNm11ks5QZKTo3YyGuoQO7DQAAPKGEBJX1hKhJg31A6ia
I1N6mWtDqVk/O7ETb4g/JMyehSRAukdvuh9tao6HjAnSh66Ifz/Aaz4sBHJLfpB1fjwiG3CyZHKM
3UB4cNOL+vymuH6lHoUmYVBlGzjdWRxZLAOh2Izt3XejDVVwW/NFsBo7en7aWNxWd28kbEX//pdC
7TOOQHriCaZ62W88rdTEQR1uQRMXUs6gN9dnJyL2tZopGQG4OQOIUja2szO3JKazGLgFkE0PTLHq
9Zm6vC7L8S3d4FkBY3ADwSTUTTOXmhZ+MDD1/tClRCoceSlgMLFVzqmA4jEbqde4x/0QSct2+9OC
QBCjjoA7scD3Tzf7xuwVX7nJ1lUSeh/0iqlbKT9ngI2Z6GrjVIA1NmqINQObW+/23q2YLyii20e6
OMQ7ZdZ1M5Uf9KOALALCG7WzWBh/9z7ZNbwQsZEnU/owtGew3NFSh5tJ6rfmRNWRX3kc+4dyEc7m
exCafvmo5zwSOmkzGsG3WCMhOAhZxalm+O/O6L1H5w3i7e4Gq3Dt0nHQfIO+xyg1v++Kgo5yYxtv
nqL/6N0Ng6vR+pQF/6+EgLlo7HnS0v2lwrGzHU2eu2bAMOeuF3XyjYUM9pfoLhZcYJOmlyTfF7ql
FsYDeydRi1xQl7JKDosEP2VWV9lOO/yfdfysfKlfH3MnPhzwlyPrYy90NB3XwA4VdTaFL/xvJiuv
vJpWUozbO7zF8e9IYi4ukpMyfhooTIVcdXvps+4DW31zuPgoECvqWD8Te67sNkn04iLc9XN1DL7r
Dc2wbxnAqCUFwhUbRPo5uYOaAGk2lhsjXiTzbSwioWtHUduUvYwfESPpKEoszyDiyMZ+EGDOUAWH
SYgW9qfSbLFWhGb+IGFPBkUUjHsX5X0P5Lc7IcKYfqm4IJEtWY4G8SkRXo1vDBVaOVNGWqVtCHRS
5P7Jlx2V/m9hZ4qIhkPGjjxsjpHoL0E4FjCIn3irb2wu/OzxDhosfZI1TYiiS4Ap8FMy9JIGzP4m
ao1+mOFEigIyUoBiMmXd+9eqrftk3NYxtHf7fugpswjSQiTkL7az6Nxw/0P0inOjb2oXpcGj9LBd
x7KJru4tY7682bE29B80Qb4jesZjOW9zAH49VShPSCf1+WuJZjg3BVdSXuxvn+r6Cvc0VkYvOll1
MDCf+SdIiDv5qkrjmotUXy9wmzDOJrstMskruN9pAFslMpCtzq1LY5AJvBSI5FeJS4eeFXaPaiz6
d+us5OevVEblQTlf9NIcwDWi9OSRmOZvbwTDF2pZFSh0dCB2uI+vLPSR/cCwLca0JhzxJUJCL0ua
mqxWhfg/t8RLU1DEUwhFHYI5Pkb1wWeNK/uNEXDcLN3MMS4HO+yIU8c1Vhjm+dTgqtYeujB8hidV
AhGI6nt61ZaHNFuXMUasGjdpJsqBK4JhxNsJLyaHuw1EwPSAKZHrqWwNDgWwaWOSHr1rfyPfbe7t
3h2FYSiDXsyoVppNz+eutKh6yKgdGe8qGVe0JCH6sp/n13qq4LsuJMgeTS9KhOo5DmBtrV3aXnru
sjcOAg4WYx5XjGfI2GVNJhGF38rdFO/kaM30Uwtd4wBD6DUfhbAMHf6Uppq6vxKWgVzzTIk6pMlP
fWh3ADOSXdFDC9ddRzaY+Bd0JrAXGlIRNN+GkUhKrxwA8PG4VMlHXVS4gyID+OvH63QrO02TVW+Y
scks2wcSwaOtl6f1H5Pf5s9vi03jxcQ/SRPVLDagIPYbNEjhKnwKlvfnWnPIrgxAppQQJBN73xYh
WA89LzIWnK8/mq8TUSiqT4MjgBFRxUNtUdN0DNC0e6SsW4eWwYZDage+CebzW0S67s0iPh5ZHoyk
uxcwu1vkiFWYPARmW7IUozgy0L9vsXRfQYXZoelz2Simh+jy7gS29Jq4HBNNBMgsUvExtqMxW6cI
dvVjKEPO8v6Saoo6LWdaEfbnPiIdJLhSryxy6XY69dSg9fLmSHhq1p2jcb6Wn8kkWMDnVrNNwSqa
8iGKA0MknMHWVSGdwrS1eGaHGWtCxd5qBwXBoMaZ0ym8hd58A635Myk2v33SlLDx6Jrc4qEhSrsb
N+YbPlMYIY0TWBRPnHg7dopIPe1PhGKDrjrBcKOqVIKxUm5N18qtiSGTClYbGoLqaIsO0FECxzR5
DSwaNaiFGVkeXyrQOJlY35y0JFRRxDSfM+cpOIqyB552THsPQ27IaLN06h+OjHZNV79JRPESN0mp
wCObskxmMfhjtZjZ/7sjyW0RTfyCih3ST6n/hXXY4H9QHfpG+DARneMizicyaw2CXYUWmgGBUJVy
vjKQJXHdfiGT6J+eex+id51uS2tV6GXZihe/SEPrcH3Ai099SAMYd7WITk+u1RJpYjzpUpGNrUGL
e/Bori5kobgfdtsIkSJTWzRL90CyEK3rZvq44xefkOFI7mLPABMldBIUWANJ/ray6loJym0GuKBr
jtNHvWUqxZQ+faMuLj/Z7lDiQfFL/3QrdfX2Vs/Mld4/5YiGJho8OWC0NywmUN0Mlw8mwzP5fi7O
n/zGbTV4wIYjmeb6cqAb916bxubnkknsE5Wqx+sPVQwDTd8s4vY+FG4DcRXyWH8UUZ61wmX5SUiE
a9hM+yrgQeKuSI3nZ/FAVCI8CTa30HP/erlYsBgl0nmXZQ4P/2JEdbCsTH0wX9mOdUsv6gEZ91uW
WXWGmRY90ilNQFD3YsFwnyG3CuGnZ9JFsVqJZIRNabGlFqNiV19aU1FYPFFpF9IHlSQboHlTQaKz
Q+NYL1ZYLjV0Rdy5/NuV6bOh5xqbh+1obN1HJLTMA1nRxjMcyvxNrqvda1tO1JfrCe3OhxSV+Pzn
Xz5V0cqczd1vpT220jWBMESKTFm/HiC8wDSMLu1JHb7x+nFkQ0q7RR62VtL0iVgzxjfXdL9nsjM4
cNQTogJdaeap1b29LSpSy67dtLFgmI9OsEbYjiBv63WkXtMT61pQZOlvPZiVisue8fuSOtZuTz1C
rU+L9PX55ndmoS1EqE4PAgdzB1rfPee+yHGS4RsQmSelR3u/iMIKpUQp2BfRRr5nrH3+ubMcX1/r
upvO4B1dvyyMpQWFkr2MU20iUGhlZgVupbMrI0LQwRAEziGGj5WE+K+5Xchg6y9txAuTSNz+1/JP
JPyfgJsLdaGb6VOAvljY0TzIiewKBGzC0TyxthpgXWhzp/iQVYdqn24hfGAozz9LRR8lQxcwdRO3
zNshYTE0hg5wFHnZc6bdgdTWjutasbUptkDCqmeNSi6G8gzxLjRglyMLxGbnsl3nLK0bWdMqg6i2
or2VFfJof69g7epeEWyxagDhTW2PntAmluH2vnshbZNnJt+4WdVF4q/k1BAF2LfqojDjQZym9HZo
tDygW/iWI81qmevhK63wSgtuPV/BMG05rmce2mP04huLld8vyuxHeae7nOH9VBUULqOeyftDYWFy
4VDyqy1pdmvLmq7HwB5v/WtLV1+6p/ddAa8WjG7bpk3X6K+aVhScwsvwphrcAjLS2+5rH3W9beJ+
jTWTrNVIMtDutC27nxfrkWWuw0fSFjJXj9YgZS/LaLmDFWfheCFAeK4II6+StxciI31tX18652ch
iyVgr8n4zH+ktdBMHtVdYaLtYzaQRyWsUchbtM5bDx9vYKK7PBJ4byCfv8daz7ZW3407uCwfHQu4
Lh6WU8dPoprXoXHxMhcXoyxDB8U0vzK2K27PD7/tS/aKJ56ll4vV1FaiaLHN7oWgQ13Hb282Jwdd
oJzU94JVBCywJEWA1sV2iIm6qUFwkBQJvHhLKln2Ft3RHZk0Hp5NlAg0jnbqjTgrA/1axA6Q3SER
n70vT3G8EzOP4zdjLxXAo7qM8P3YYrufPzWIgxANLB+xeFPIaiyb/X0hwG9jnqu36cfoD2w65bGj
LrKJWpqeMKsao5E591IaOzbJLqYgnnK2h88zHIAEyHvH+FmgaTTG9jAqzL18JlqBKKqjXLvfby04
j6X4jDU+NvGWyi/Ke+swvCqnYQB006T7Ner7sVT4A6DtLVpz+pg2iNRU3/oJ3pIfvNjnyDPuyRld
yljO4gn5wCVzKcZKkb6RaQmufVCtps2NtA65j75b4sW9hDiUrUntQ7m4xtPI2GCzLRoggFpYj0Kq
9VAIAkNeJV+a6D5q7OqanN/FAqDVczRyYMxkCsY/jCOiGrI3f7uzDhfECq+e1zhYwBZnG88K7SWg
lO8Y/pMsu5dVJ97qA/BZ2LNWykSaq36YeP1Fe1rQKnbLS9ZM7ygFtzl9NZsfZQkWr4Kzs0yCu5PO
uT1VNOwm+yWkNOTNJlQ3vs6r/3Cm16O3+Tpr7lvi0dXac0pn//7IB3O8/vwxlntQfMDij9M5HXD/
7I0hHNFPPqxmXLXPmLjpP3rNz+3rjVdH/ss/irftjW0KDTZq8t5hv+7Llj/ztpuGTJ2aoHm/kDVo
Np9u9ld+ftI8qUzldSkwiFRqpvL/Q0j+1/kSzvsP4HrJ8GVggPD4jJkSAQddHLSK2QGo+Xj/WjfO
R9w8kF8QTYgeYAQdjaR4BsEMR19XZ5/wzKMgPKiZdQ535hg54MqyLefOdBjpv6DvtLRgSd5yfEB1
qQIfQjIaofuioBpr2/S1nJfFH9mHGCOTpEQvK15W/T5T0oISD5LGr41mf6kjY+B7Q+aQI9A3B4n4
UFyPSJDgNf8t3vyo8Lz2gJWIQ+JjJT3U85f+OQYdL01amMT88Q1ejtbmiN8Plh3c7eY9u4tNBTqL
jfKbfjjKoRkIOum6A0ZjHcaAIu6END2gBv5i9N0+A5Vj6GGR7SyQo0tZ2Yxe8Am3jt3QCfNdO1de
KgvrwQc93j4uXlopNHJdmhYyRBgZytX9yAGOJRoBUzj8Q7rX7QfprUa13la09N2JHRuWUbPXzlJX
JCdUev+Pfy99FPzwjQ+Wn3xuOr80gJnxvEPS2A5Uue2wp2hLFT+HLBF2JY+OyWPrxl1iOwksoC6W
hETjmxbXU6/ir5LdtBnM4U9kR3iPx/jjFuDOoKcEQdy6haNtC8nfnEJpu2jNjjrUgD7vY+3i/Z/B
w8D64dCxhICN39Anx6BHQEb5VPKog/MCxYUecvZWwjYWylNlWCAdMAu7ueCE2L/+wtYU4yuAqkGd
i6lu4xRGoN4RVXvuAylx11JaPlH2e6qSzJUXnc/6/ArVemvr6SKs1kjcvhW4FK0kGdYHGSMUeVYU
574mDv9S5e0jI+07YxNP8TD5KHvXwT7b44BfMEw7C7FoyuEz/3vhGwNjrIjfNEOpLKWN1L4aHrN7
35KP+BSCJkX/MoD7Z/rlc7eY/BPxGWTskCaz7x3btz38DL0Dtwae5y5T0RfMAEjLFKWql0uuyFaj
Db1IB1X5as0m4TMxBR4GSKa2q4seMUqqhncMRtVGMxh88pSfA7NmvRm4sj2VI5wQ2zMs9kdBuTAZ
FNyX1WGVONELw1yTPG+a6gH9yogjPFIQtqpbnGoaNrEA7sfiFftnwUeTQvbhqExtRh0+kfPDoFOA
LRazqV0zAvTZ+rt2H76XP6P0y0nOrw4qmYKjxyt/Xt9RbjUoBKl1Ey0IYaswjrxhYer+5kkARtls
j6Xlphdg2vVv5N1/TCEjQ0kkYenX6LSu/itSeKHnRLoVE7TiW7D1jwY1mp3hl5AIU3XH+nkE6Z3Y
qkgEduVQS/gSRmr7OzGAl9DZ38UlG+6PCzzVyz0GVp6wjzGpWVQWA/nd7k/HWt/f5UFHlnULl+H/
266aaUJskQjoyERxD/qZvxPvYLkoiWujODrPrtWJiDpdmcLUpk7n3gsx/0Cdbdk4XYS5P22t+GE8
a11aqXhUPgYaiNXRukVUg3Ug9T1DjvAHIC5SSh5x3Z/HkGIInW47L2+1pnRcLrvhVmaPJkHF/dmS
GvHotwBEZ1ZKsjI0oBZvmD7ZNEHl9LWrKuUn2wT1Hy/i7fzdovhCTef1JVJRDZQdndMpoZ7JgVFC
RcE4dM3yY8W5Iq4idGDFVE9t3+oNmPJSqfE6YMZO3tGUPVvX/dPfraPi6cjyvLwqXGf47ExwVTSA
x2BZXJYurFbb6xtXAWX1L0KvdiJaZaEVZ9mpZWqTFF1wX3mSUIpetL9EVITGH563KZzptozLXCOJ
cfMFZcTMjgEFV9YK7hhKbalo0QUHgKgs3LgLgxjr6wazWoO88kOuNOXG9Mybwem2oBBQhT/8uUdL
rWGJuQaRhNHCUU6CCxlvA16LI540SBjFM37Qv3dXWxfUx6kw2RXKnmdj4e0Jw8ccQ0JdSlsQaQyR
LKQgbbTURzPRRK+O8zSBjPjb8xpbTg8Xz3w2mrYwwF5+UFDbMQUGgyz05WmgxcGBzRam6hjw31Z8
yYd1exbCaof6IUnBRFGKf6fq9W5DfjVYSMJcH9QZlwUNqOl477GoQugQe5saRqZ8xW62OLclzTC8
PkohjXxWn7A3dlnYH9bdWXzz52KEndWt/wGwtL30Vmn3bqbgfAYg9i55wQTdJHQwXBaG8BNVWJJT
kDX3ePp1GsFiOASK4ifgNsh/uMwb9hJjoP03rdAwC7kCPcJtLR6Qj90m2RZhGtksX/kxZJ/H6swe
ikTlMpXAEzwrQKYUNFf7BXt49L090h0DMjMDxj7G0YNv8jvcROG0vC0ko0S0QhsSP9q9M7eqYliB
+8fZ8NibD9IcUU9kBqHExNoItMAlDHM8gKHd1UlqelXEkklMM+RJTuwSoLIm7/Ktp88pxrAXy5Q9
i7t7bj3Mk4OeSugyLHOO7s/pnoD523Mrh53ZTmNjMmxrqQis98SHNuYwQcLdR5nJNAD1QZbn5S6J
p+6Y4m6Bad4wS6P/+4oJ5Tuxy77m+e+8DLMEWK4KixzEKdT85RwgfxKRQhGFCm1AHCfRohY1jnSn
uMwWEmm87tJQdndXHNf7pO5P+AQxD1oOpqT96gEhH6+LNKMjQlO/tk+vdzg71EV8vLZ38kkI+fmQ
ZIbfdSBbj/g9rC1DGZxY2RRAdmZCsbQYoZWOx/zzvhTe1f3AJK3SOKHA0cGno9Hy2sPTA1UcmK3j
cAtypJ1XfOokhpcLwzDJTSy/lSZGRPlpTsK7uy8jN+LJ9FIZde2MqSTzxx6x7+uCls3jZX9kTinI
/hbE9PouBOtKNdFRUpPtL1tjuWmymBEu/mL0IaOYV2ffEl7XMjJMziwRLWJFnBQZ0UNDTrVVN/OF
+UtfUcqND2hQES8MgeKTKPrAfhqYkzUxZiUYTC+FSC7RnKpFikXepqP+8J2V5wPwpgW3bWJSYWQl
zIPhsZdL1zrAibUZ4MZAQSYQTUWvxxFVT1+Xpa4TeOOTZpl2XcZJH1Z9v2nWf079ZLuKX8+haOa8
g0HQyc5qG/qtNbLvs359AWpeaCM/DXNX+mYRIaNgsiVGWujjteuJutFXyYULf4O5auQ4OS7cb1Ru
G5635wbLlpb5wFchLqEroRKFSOVCzezJzPWtDiT1uY8Z1UEJvKqf1/1PiqtZPYn5qxx9nKZwqIgV
IzIqc6niE/k3Q8si4G+MU4mJ7ZbPisTKHy2RNd0T1mU02yf8owytIakwLgnlfe24qmHKXFdlQYYe
QIZ081APAnmh+AUsZA834Y0Buh9+cRGxaThAe3zejxRcJi7TCLZWnPJxpqMHCm43O1EBSg1kojmG
iXV4QcCdVTwvjDkXZpTUocTgVYk3DRSy8z/U1BoR7B4ynLUp29ty2NGdbjB0t3jqpaZ48AYp8u/U
/vvfpwJFSiZfug303G7F3JbSZCswpbKZvGQtCGq+5il9m9YUEQ7vJU2T1qfqs/iQTJ1xkg4Gj/50
p+lDaRN/70t4QQupNpuPTztLXyhUzoRKCSbUknEBEiLrAQBXmAbcQ6CBjcw9dobYHEUkRRgoh82w
wRwH8T7BdmrH6Vl/AHbwMvIagnJReGOlmnuBqXZMJFvI3nvqxL8MO+MLC+PHMyQLrmOpVDQCXX6w
YhIs72PcanoNemvdSg0Gx7X8d9fA5aWnf4n3kFNfFz/yC9Ua7Io+8LaqVm21Vl+1FRWPY4pwyQHo
F0cDmme/KFlETPB/m1IoD7oqDpXSaw+zOIHxrcagdITDNNEoJB+hBlrrrp3gt87uvWviBU6STNV7
BkIssCJkaO7SW1/i7DZM0s79rTW9+psDUVj8Iyv1/x4D8qewZQEhvVi1XysniTJGThLMuKH1Q4DW
HODQl57z1EDNWguTs9EBBOhBgK4YK0VsLXaNiLnwBCVr4qL3oEpBBW8/kbUMwcuS2piZwt1fMtd8
JEjOj3xLcUsOOdQgX6+b2bUtJ2vOY9cN7m58jLSCkyz95pCHGv1ZGbm+gNOk2ehnpaGMc4c9YOyo
VU+QQ0NmoQdnzuKiUE49m5aY9qK/78WHJxXISWM89rZSIodz7iIB/4BcoC76jog7lnop3LW2f98+
b2rI/y9Sk7UEQ/m4e7SkRoyz89XU0Ht7NPS0DxGXnSzgI45t9S5D+K0zWY1e8h0t2r55bYk7HYYY
L4mHva3jprAMiUeTbPAkHgpOvUV/b1klWCxe5lwtKGK/qFMC1bis3JzUXVPkSHL2oE6KB51VbEuW
rB5TkP7a7SlLknBSwDWp3Z9jdVQG/Uwg11uJDLN7PpE1k77C3kYlA+VKCOxxCMm+4nW4R16J+dx4
07oS3d+89mfD72/e4Yz+MlXd8DmVJXigVu61hx+nNL/6ohum8e4O9t4NIGviUtvk6CGPT0uuNQYQ
x0aoKNGY0aDC2+1nCxbFgjyoSLIX91apphEg/GayI6vM9u4Jq1e/K6yq/hN4v552SptCQEPPJUou
DjJrLt0KOtv2WN7wkVZ4XSOVXykkE7Kj21vmYLZzNKdsRbFcTOOy/QlJ5chjsMGK8bVWevugR8km
s8y8YJfUSqymDuWV5SnuHsYeYOfvxXF/Otxt9hSzsqQ3lGHLqvF4NSz4T5bra++BcGiPx8SxrSJS
sbZ4J2+2V5qxHW/MVucpOj6bpF+4Kct0GKJL6fodMOMg79afGO5vDrrG72np+K2eoPRztao2vT3H
jGPDWAMoIxZBguqKoi0euBVrwF5WPjQsIjYxArx8G2ar6Id5HTVngf+4MNsnlCmQ5u4MxLfbHyML
6m6bOflu0uYRfAAtd+B5XH0ruWOibLzi0GKkP4FQBdACb9Iq9ScwE8w3da9PpR6R/aXpc4lmqL1T
zm7auwLfLoZHGXBMJCJB0KOXPXq3phHvuBGvb/snC9pmI2whDFUL7s0dpUEdMXdJRebyfo4yun94
tIe3CZ0JQKl0K1P6LP5ZLrCdwqvxNjNlQuj8eiFEx8CH2j4V4OItSD0tFuqfgqpLCvA28fLZ8/xx
j6/TK+rFcssgbINFeTAnmS1MSpGianTESEn9YekzwwDeTxLMrVk3GgnVPkmJ8B/+iGrYCJnrtq/e
4y5jhDyHmbnWxrz3b9ddzoSpKZDZ8I7Gk6nlG91qgCM2lpfrDGfYf6uLCbQrDxvhXE6BtEfI5f5x
w/BeahIQbpVgAu0LYUcvb82dWSmXsk2cWog0nG4DHZ185ZQa0d3Ga/s6a1RvXqsIbjC4DuAAa2xY
BWmQuBphWNAiDFHhwiTFzruZElQ/2JFspLzMqix0lzPYu5sTeU/iBJdKPJEMcij/k2kGmOQvub8Z
epfutVJexCgREr4wf1hpjXQzPVQJ2H+pghQalz8hUBSS0bwxdhMZchkbyNv7cZc4qYbwJsfoyxxP
5YqZhEtpi99Yw/pNNM+gPfX+Ppcr7mhlllKXfX9obOlBXl3/dNfC2bF+hT4VdByQ2Uj+8jSVChpx
pk5jb3OF+DPFJqr6Wf3ZlMemRia0uneTgRB64mNwWkwgJ78BWhHd70WG2239kpw3gfPXOYkRxnNW
TspIsYntCSxBNepVBtPpK3XlZKZRCsUWe4asjtUzlGDBK15Hhkm8eLt1zceKp8GsPTWzRgzqK8SX
IfBahR4YmC3YeSwD/OfBpHaNiuYELLQbRcw0uk/vNwKfqsb99Xam62bWaPBo+EoahCOrSwdrQOa6
99PgYr3m4rSkzF7wOt9tdIezQauW4/2c8dStAl6HvN8TRB5oSgkJVRAO+NdJet2M67c7Ta5UgWxe
EljTCK7+hM5sQlg+UyNKxEsSQSli2XG4HDS2GylWBnOW5BeJE+Lai0erof8xAS0pOM+mQ0JOBefs
zTpCObZWV1pa6Z+0V2+6MkNyYYaizOAvNheHbHbvPEZ6mjG70A7uRXy7buHJPMC4Mqng/d0a3Rkr
kIf3jkhZo3XavNGO22JEFo3zsVeHG1HArzn65SFuTnHF0eXte0N+tAcoPz2yCiyfKenFCLt7wfEV
b5TQ1OYLYw21HkfBjBPukVMpkQ0nkYC53SY+2hPe05w80akCLQLrZnnIBTVVtjRPAm2L8/nasy0s
21BFSxgNpMv7eRrnnZRP/CfE8faKk4ZkDMgNJ8AlOqeNpk+dhxjMrNRDJ4JbGNCGn3gZc+MudfWw
oQGmyCkBBOB1rcWeZ20z2RdlqBLML9bVufwkLJibTmr48bOqyoSCD988qy4palXm4WWHgdvinbUn
ujx0ffYlW7Ae7CUoakl0SWormTFwKe6ZkNssdv+DLHszk7i90wx0u9REXGxcQYrxkzQeYKeZWwmM
U4qe5BzjVqXw9Xro84GP2+zLNr3V+l3kv9VK9Fq/xuINzgfpxRlr5cM38X7M+BfCDXIOtkgqAu9O
b6Thhh6GE03NdwCy3etyAFl4DRnVQAu3BmPdUqmupDanLl6XQEhmgEZj3JYe6mf9BbWAMhOBzARb
u+MbiRs9d+jzcBAMIyFLcRWRJtn1LU/IBxcKurxsSTseWKv9KKc0ercdUr70/pU1i165qm9/jRtL
w0f9Ys4oG7x93C+rYn2J0OPB+QCeepQp8r08qP3TvMm9zvQ6Q59aaZtq38AdRhr63oy/itzoWegu
NNKLRUhsuoCLShKx5R50EInk3FffGtTRI+dH5Y9ybkxY0P33RamX20vm9cUN23HUr2n8DUzm1JaD
gEGuF2o3H1TqvGZHB8oDhh4pqil4SsTUgI9sznoanzYPNdEnrugPqOXknCO4k1nOQQf4v3gSJgGh
vQfDHcw5ojgZb3cD5aJlEulmr1sMGWtNJ9ql764DK+DR0PtlAxlMoJzJhSGCo6CNGrr43rx+kWLZ
sG0yUX7DTpFhVTGUrn+fCc146Tk9QMtm5Jiek7miABOWr6EFLaxXEXmQbMoYJ7pLau/sm/uVOIoH
wFNa/la/V+3wU+33tlBCXiK/1gw4c1cZ8YtgDPsxGAKrh9Er/cCkmifuE3jHyogawMak1ETWYefP
C3GnAlQf30kDZLa6/aJ37d8KadKkmoDn187LbwzWAmOMEBkzp1Py9bV6LNxni7Jw6jLnv2S5O0QY
1dFH5r79Hguo1NpvFxTXVsYN6ADFA0tlFST2HGztGFrMn8JZnLJ/qBpUzY7gxPsM1fhTLz7pMEkr
yAgHvYCa3alFwG0Jru3dRovRGQYiBWpkBYkZBQtuPFGBypPsYxKSzuqRKupszZYZB5YwTQHcTHhQ
+ohSNJOEydtuKH1V5ydgevx6z59MWVEPefa2mBCshUN0WAVzBE/tcgVej3H+MTGFjbWoFb3cYbRN
FbUAHr/w6Bnc1Dd0wfDLA3cLBLIv6e1QPu3q9Yp02LZOj6X7fOfOolctnC3dURXFm+t4KxR1F3Jr
inHFASBEATt8bHKtVss/w7RThmY+Mxw9v/1ePQ0Lw8GoFERCSnHfn0ERSZgRUZymXftoh7Z45SeQ
PFlZi92vBYHEOqqnsF6GcVvXS1hphXJCCr8S6hZqXUrfX3oDKuYAE7tHJRMMxslxJL1ZsWxumKl8
hdS2PLVmbtFeJygcGS2swQib80YHV0UWtiBRue4sWuY+Q/4MJrsKzHXgVJFfDc9XI9+cSjLaMXxK
Y1OsSienoRkmdW+VDQkYy9lVRIrKgWFVgXCuJF/foYvB0SlYiWNMvo/jXG378zCvJ2+P0wvG5G61
ReXRSOqQ63Iuc/XZcWxEgZ+JyLVlXVnzpqKlVOBw5/YOTpuQgVs0L+EmSo+DmsiJH9tI904uT/50
o5ZR4el3gB3DVJDvvudUHiuZOQW/gg729moDTkczZMEli050REfQrewN53MKqmKOOCskAku++N9e
KHGhWVtL9n2N2R5kBEJ57zKKWyTJZbNbbvDQhUIe473ZOb5+g07rUJU8UeM/6ulXQ38EXnlAfbEc
pempGlFaFRiuBELT4gtInxgz5YqMyRB0WDYBYtEWjQfRLajZLxJdSl6vk4FkoPKcUGVFwgsF62ul
us3sxhkAsZFsPSvTBzYuEbO1T0bpzCfPmW1upM2P3owL4Pm6Uj1uD/NiaF83xUeZ1NFv4Tiqhvli
D+sJFFiP535YqyRYGT7kG1BHQ9dw9pNDzlRcEoBZZ0+sYEyewsnDOPvV4xFs6+lzHbuONXF15mYR
t+xcAlq889MeLzbqbHQgVQbU9jKozmMgW+ihfltDyV6AImISzqYw14P1DbD2AsJYMESjKYHHoWwe
hEFEVF9kTiMpdLjuR4/HiX1VOWgz3UZ7YBCxyFhxWsjTdjE474wHSBwS0bpqX15rB/UonGHs4Uz9
VT1r5mRPZ0jv3eLFrGnIbbBkrpMDMLObJ2ohqo5QqcDqqOkpfSdjEqdW7A+GoRc+vrPS0sjWYsfG
0XtzJz8GKzR6VmXsw+68bfYmR5EkCcG+0NykhiFl3LrB58y4AZm90Acg2d9w7BQsHHpoHyBfu4Fh
ME8mFT9tjxQU1Myd7wHeyL5IG4pC02zue/kRwoWccDNKH3lPxkD16h89laVA5ARKoU9MwIE+p75Y
HHbpLJFt7lrL6xjWQC48aWyN5Vrixo52cD2aFzf+LFB4PKfKIDmW3Y9/0Jl5VQkMo/ZVwyd14cPn
Mr9YwSWOJjvJ5bq+G4ux7u/40FAilmaTLR9GSR48WKvBS2MDhRoFvxpsSAkmJvtqWMgSXSvcVbHU
FPpxK8sxH1dhNjIjuP7QUPuC2fdSHvs6713gqzJJyEphDPe+4VjRQswOOfYT43sVofezFwkBKj25
qAbwXNhKs8jqn3iJ3sN872/ASEKpyFvV6+GG+lJQsipsqspe5mP4TbrRTuMt2pbKbO+GLbsDOmkk
SbmamyhDqu3Zl7yiCOFInj/uHs01BbKcnmGCA9fHfZ2BzPRuI/dqxLmYrddMA1j4Syoeh7B09YoF
numoakfxoKtMpEAjpOmCFlUqTFH/ve8KMuMj4HCAhdFVNruDDUpfA7OI+g5jfXvqLVnDhtx2bfjN
/y+zDUxKyZtiXcjsASFmQajtVYjhKZR5Tu4owOXjReN7lnF68cNx8gwKGAjvJsd0eyP6qg74Y0r6
TzTHL8wWnfZYk8qVA/kEtF1YGRHYKa10rZ2xdh88mlh/6xrWTMB82PJWqHZDypmWWYTM1W1dW+DU
Kz0IoiMYH5L5f5002sQKYJwwiwoCvWmgw5etXDnnvybStBJt8YAXYb48O8HS/mGstyWHVLYly6bi
u5tPQCQmQWbafiUPkv6mqfS+uQsbKD6PmPYGdhPu/b94fbIy8lV1Gx40yJhgdUmDxshzgeqQ+0Dv
g3lRQcWKoAX7tToBWRsA76GmjVOmvxEvTGUsVr+/uUZ62U2uLLJCYxHkBFUxPItz7ul7BzmR7UHv
QoFmbA5lOHp9KT21I1FU4pHhpZcZ0DypeluRr6IROurebWfIWNjyzpjuDFb6aUIccAEOsyHlv/jL
rr7rOPNqWG2DhxjdNcaRFZvLzVlI7hfJov1X6p3rlYJBJS1mQsAZWaW7Qzbmf3rbFJNpvUg6Jv5U
SSUTBiXr6Uf7xYWRyqsS0z0lD0uXv9BFT3AhX/0FXYTdmru4p7rgtH78AgNA51l00muLC7F89/+C
h6e/p8a3NstQYsZpCWSmvf919Z84gHLXLPvN3aZFxT/N4zlS9X2lxv74ruYnFtL8xJRPQcqgsvWS
M4ifREaleuBI7Npk8U23DUf+/mXKJ6dvH4z48xdB/py8D2V7En6WrqSjv8t/GgMmyNGysqSbUFsO
OStMsGKRWetVD/XQuJfX3L77whP1w5ziIwu5diZH+ykf7Ox+P4g2TAcFSB5u9toF0uq1gLdGvzpk
hpO/V4EjsjqfiCyj/g3YcqK06lGpiYCvheodWYPwB2z+B4J9vC2itAcXbYSU9NtcNPy77X1jAJoi
v+t0tw29z0zTnt9eFwZYdC/JHzP4f+vW1JWpIdgMHMsvxF97IFoIwpRPTa9bvynKReGPCZyTl5VE
nz4OY7SXlx/4DW+zxbnWLwaROAXlzOUsNFQQmLEE+QkY+H5z+j5kj+1jCUFcQwTVDJoalQtpx5Wl
IZMXi/GVuyhBl/gkpK8+V9gLcVlqEzXkds1PSzEZ0wJ+Xe2SIgdACu3BLD2lIzjBaS6isDwDfUwC
IvG4UN05h2SGv/n6wHHckvw0swon5v9/NS+/d3B4SZkm67cveqOeF95glM5zFBmGANfMu4EtNIJX
UjVEWiMB1hGPAU4Xm/BbtM/+lDf4S3bFWkwHxnY/OqQEecTWw8HRYwP33+VFEqlET5ZzDVKwlbzA
zTc0t/x30EYY1l+JI4ZxvJF/ROY0PiQAA/t5cGqmvwtCGosXTjFAqUKlHiI9jm0tyMuSJgjeJVxo
3731j0GoTIy2SF1nrROaqE9B6DlVFjO6yWRRvU4nrW9hxr81R4YVkLpc645I9moM4eA/v7aN5dtM
ORKCG99UVatQ7G/1Piww0OeCGqefI2FsdMnJ7RqowRUvCCIvKz/1S8NRIYFyn1/G1TXq7diKDl18
53EvuvgrAWSxTnUBVXXeKgbivomYz+dvRTZuYgfgU3Fn9tpquP5vHriZpFGNOqOv2b9NPMNZuyOP
yKOe4iH5T2ihxZ49BE+eEmMH/YxMSrDSPtxrdaGK4lD2mZh0I3fU+PEMUrJ5CCH7IVhIWzzHhyyW
4AYmOqtcX2dsV8pS8MvlVi8725y7SzC/hWdJehDmyh4Aqlqh3NMATCgYihjXL84Eo3w3ukmPRTGM
kDRyqVuiDw7jXG1g9GgqEEMidVZ018mBb7NNniI2BmQbiGDM0PM+hxpGc4kbVlYE77NWQMSNo6+u
01tg/BqfKOou+M3CyoWfdH03lI5aa7GSM3m6LHV3dJ/xhBaAnBMc7SCtqUbEQmC3tFzt33xleFbi
M9wegv6/3pUgU6Gp2npJrX4YB4swVXeoqWZ6LBj/6wzUZEauwlOgLLPsGWX84zYDpx74ebsNzN+o
Pe1JMRFCYEGqNvrC2CGD9K3RvMm//mctwIyyhfrshIYG/YrSB3I5z1hyOxIVtXqMFXVMjrnUDPIC
DwRzEFfPP+BsADPLx8CLTc7wW3F64ggtPyq5FQDQh+uoE303eNJUDLZaWJML+BRwF6W03GARtmd0
vtBar8Kf1d+yafsA4njOlL8x8kEEAGkQ0lq/+E078SE3ncslCmWIwo7qgnFB9Lr2kgQyJeVALIHx
/WHC9vtThwcymRp6fgNedYWhADxMWJ22akx8hmxrj9F24LZASNM/lnxNEveImTLHwlAzHrQRXfIv
4qHNwTiHqC1rk8qcbeDO2qlGh79WvHwemkc2txU0lQqVd7YJKSXvbNf3c9E0FZbVsLxUPxEMm22S
n+gLhm/zGfMIgIISeOnM9STeTLURvDipA10Hu2g4sBjE88S7CbHZX88YyJ2jJGiCptr0GuJhobYp
GGidL/aZemSjaUdybbYQW/dbH6wY7A/0oIx5R1WFyByMgPIwi2AsWH8NMpvbKT0baQinQGcdWcMr
WPuwshaQsk1C1mVmRqONu0gNCOnbIH6f2zSTWcNaE7km9DaIe5OTwK6Ktsqn+27LaIEUq3zfAqY/
5DpkX4/+5YgaVVEMSfxKfZtrfUwIwIaLPYACyHfpcs3hUpq9Off1+ew5EeILNs8uQ7gFZDp7akkK
WqbObNDagYE240PqyTlpANmseRwR4r1+J8nwsxovqvvWatSoDoOmLWC6j9Pi7sx95QglxMzOgJ9Q
lTDMV21i6lOHkDVcYopE2Yt7X/3PEq6j3byIzlB2DQvZoP4Ko7mzUjqujyLR6KRDdfJqJdkBGRnL
q3huSjdUkwZd8ZpiqaKhmiiy5FRbfl1WYfVV/o3r4/pAe3AGjKfrNQjZxl5dKhRo8/88O6/zOOq8
KrfXeXhnKorBnp2PJ5BddPlQk3gK7TuwDsPixSgLzBnv3og1xDSvCdA91nzWaR2e1G52T1Lpj/vL
Q3zJi1OPJ7lBSLA/00Fi6xlDA1a4jJzpbMIAIOrJUnwv3vH1aPXSjy52/D38ry83qT2g+gAYu3UH
14V2fbAkaJB/Ut8syGxnZvXqP9mhDeZlIVdGcrCMGqrtoPMaAMSjlHTKxmmZzm0HvzwVKrFLSQk0
WsUK9WNUNWWE8FNykIW9zUBgLXBeFLVxydGHV+BC3Mf/6JvfL10E2J689iwWUlppzo/XJIUhyUrT
rt+xs0k514hU5Z4PbL4kAWDW0i3WFhw87Tlnzs+ruQgMjqUZ47lwUZH4sH1WhOyE8AC33MjT6BF6
LtayybELf7bKlQ0asAKVgLPrYorWv/+2vMNZIQpvonB7e5exSELdv6X1xVuQpnOT2LjmCbm4O4If
YUC+YlvQLP8SS4so4cAEs5N+VCuv8U7ymZnW6uTNlWBgviPrAjnQOrgxgJQOAJpS7UwGndAr3dSH
yvgvQusM7z314Q2ZEBk9tx/O/XLkruKFeFlR5Cm/KpKJnT2LpvD8teuZAeesHkPXpCExI1r+q1k0
4edeeUEc9UVsAMiXhgql2ZE8ItnHvP5Wo+PZaX8biVDbOp3TgHMgY1gBkFWtBnVjkrSe0Y8yOEn9
yAB9wgnYcM7sZwSgEYn0Vwiq/s05DjeCOMsI1zICHKUnAYoF7+JZT3v+rrSkDyX3HZ4ExDEkmHZF
azBnSURjt1e7D5g4d++4ANCGV6aydtYj6jvieBwCPGa3L5coaX95FBMDJ4VUXhcsbtVYtAcBEKQU
DPnWz/RTkW+nJIT+SF5+PqcRyEef/TNxXX9fsWczPTHEZIYYt4mruTyJeDs5r1nMlxxm9mY1+QpW
ZkH0OyRJHr0qhiFQwLGW4X3sILUHqPbc20rxZ4LHoxTukWdmGBV6x06f1W8JZ4CvDbuVBc0jNc4y
X6ubjC/njedXr9xUVkGjqkcg3zTkJrpvWGQ6YNloZKAzgJrzNpjuyGE+oNTbng7l4M8trVi8SjSc
afp2UP9TBBk5Mu4V1pSQMQmDOwjFDSb1UlTn9QfmWDTVI2a23ETcQ22/q+jDoaUXBOYt8Jvy1QhL
J1m4PP4P8MAE5ajygIZFbVROpZX5aVUwesnHGXxBIYp9gjjYNF548ZC9rp204AgCd+6SwoE/yh/w
PA65szG0lA1RX9YmGH6AdNbqDQyBizOAYnxQHxHfCIk7FVVMkDRDAsY7ifCoONrJJjxi+CMhfS4s
CzoM1G3FL/e+vAIvlA42IJubXPiactsJcUZ892BJN3Z1TYt30x1a7t2uydquBIgNWZGXXVJpzE3y
kcgMiJBW4ItVuA2oKI5+KJYrlTBBwqBEpcT+m9p3AIesoNvgvojBhDzshOPdh0hLb5UqgpmeBb4K
zjiKU+kz0+Ce+Wqxp8X2Bckllb86hhi2qT4Obl35GNW1JqSNk6jK10LpC2nY/mFfdEOTcE6n9ryI
35QRuJ97lnik6xm82YDCi9cAGs8hdJ56fWV+1NHPY3sexPpQsO956FSL8mCJ+JSUIt3e6LmIBRP3
qxNL02YXHllhdRuf0NzthTvxvo/AlOfcSLRyW/Xe5tYyEojMOguLrOiV4YgaWnODL+KFzRYGqSvq
MVtvEcYQyItX/AeFln6tnD5LQCVB8y/hHKghub0zjgeK/cnENcE1rODXqg+mlLpvdGnum7Y7DMxT
Lu0G9scGBpSzSHoMOWOO7Xqzx20ykUMKBuUzIoivGNiFhBXJtjOXR8eENIXYBXtGXNHFS42XNkJ+
Vjp00Q9MckR5TuEjVymzirjGbWtMxc7VeRoaYW6NRw6x+FRXrgkMver0O+/vEKufzyM0vHwKjwSW
Q9Bh3n5JvbqchuX8qJBeocnS5fWqA2p/4u2cjg9zG1tgUqTzTPOLm6RMxZgT/Aa13f5TcGGWq+Xv
MlvkWr8380peF7i62qxOIn0X/GJlpuAFg5c6o8E9JkwKbez9xTdLh+t9RCXpnHGCHx98HTeN4aMA
krjKZvu9ucNtRs721I/tlK7OkTJRNN5lq+q7K/HJvm62g0pu+7l3zDHzIjns9tpUqxG/tlaM65CD
pjdBOrx/xxq0eOvNcOw4o/A4p53QZDM6gU0LbPg+SplykCGBMyAwWwGTuhaLTYTg+22skzK6hH3l
A0WvSc8KceemcU29eu8UEx6VgAUsbf0d+7dGbpF37rg5OLD+lgCae8kjaK2Mr5rlF8dhV5LF2jwH
1T0HV68dpRGrIDAtZgoE+/VvQCysVvXQlbaQ781ChR1MiInw761W2Dgu8F6HwVsSxrKG90xIpF2b
NgSBlG6IRnPdUGg35BnbFRTt03+5WjmmpR/rCkFOS8mu+NQAEuS+xz3MFwBGOChjgpXtQ/Hj1CQe
oTTdEKeiVldR+4JXdkAYvP0AJwut5UcP0bytFYg2DWMN0gAtG1Y+ci5ZsQCuGFOypzO4TNSGr6Vi
HCs8YSo509Lidk7WbHBhn37mUjlgmuXXE0MywJgTtypr+iJFlTTtSdXjkfy96WncbL3Zs3ZJhoc5
gmRKGXYcVneE/fQKWeVhWQQMR2XtxhcTk6jYVbo/v+OPgKrPvbDPUVlR5ElHJeXILzSUdIoX8VKD
vzPS4AN1fjJeKWIHa8TZxGxGhqmwtIiJbcZckF6JF7KfAdY1QZYUa3NHS6g+qspgboyis1Dqqxli
lH/qHewEOEpOCPL5ZQoWx9VgyLOKF3dHIiQCQ5Mve6i1ROUlZ1OvBVEP1/+XGUEh2tfBKFrrb51K
Ln2tgOQyeq7ppRpbaq4AKEuXpjE95ZMT9xQss8i/uHlcat6GtnUAc2Z/aSQveDhUVVrSlZ/OCZqH
MpX/i3k8UStWCW/jklGOFjR3A+apKuLcFsIptg3CT3ACkEVeYlnGKTP9GmIaw66tZlIY/5mda+eu
8DZoW+T87q8wy7AQTg9aaJ1PFVmnulZFhaJiWdmzfe7EcM0zD+Qj8C/xTr6P71OTEuOoypqLdgnB
Cd+F6JQ/kWXpKqIFEev8AD/iT2t/Kr5pVKPrkTi7BHNRSB6GAwgVxD7tx1UVKZkGPzN4redXBjuz
uDRIaW524n9V/DHZsECt75cQR1F5D41ApnZUUmluWrFLKl5Cn9s4r5U5wXuuYONMKtMLM1G4df14
/ezE4Fdatv4EZM4fZdR7aCfUvvIkJ1c9ed/kqC4Nj7NF6XtERGCSUsguir+kn7eKJ00F+P6U3XN9
NMNcku6l9AE3ttrPjvdbNhkoot3wpqUlu+E01gWieqHncrSbIrPXf7lQYLfnCnuutS4lItJW1Myv
EDqKiUE7EZSpVr5DeXyjV6aX2isiVO0hwOLH+D4qiuqGL0pUZFN6eZbRQymJsdrMUPDC3qmLeRrA
jP6HyZ6VCZNExDKTspHQwil3c1OurMjcyTsvIfvDNW2YJ8+/DJHfQnsDgUA0mpe0t8Spd+FjLqNq
Aa8H4Z2PUaf5HFz5JTd633iOZE5ybsnSyA+1kWZwl1HuachLJ2b31f7r/vNWMJKxq82RjpGyfBmN
HcECGQDkEIlLAIoZ6GvBWXlvMlne1N/I5NxATXQ111QWX8XNnrUclp+plpTXI1hsPiUUBaqNH25I
ftJIfvevTxSPCakkH+jcD5anuYYOsRHsZXiBnm6t2zN3ZeHfsVGsJYFuxKnVCKIFpeV+2bOC1tkC
nUHZcLy3r8O6XhPQVs1uQdWPxTRoCOT9UGYAKKXL25Qh2bLxskoHcMD5pz8NSeMVvASl0ABsPjNG
C+OdyCXsharvXrt1BJvkMjFgVArSqo5uhpAZHb4+CJxsZKwgaFwjpbRyarT/339k0FuWaC/JhyrJ
1+VQs7m3Vn1SDC5pdr39xrDDpaJFL6tmTvLNRNWFRmSF/AY5CaXkR/LA8+CNLkn7k9tBrgEgZM/m
DfCKPoAVrE2HPP4x/knerPrsu+upmDW1bebIjVHPk7GqbfevRGdQEpW9uOk9dFOJjBtuGhe5p65j
vz1arXOl/raTAPWewpe2CBEcZC7fHWeOeXHbDB/xPgcyh4ujHpCAcTSLz/PSZB75ai9HF5SwZvsY
zaT0hrgimH50P+Bv/yAyZUrkBvBF2vKhvecIr5bbFPr2CeQBeuAtsNYHtdnqgvm7uUQm9tEUx/P2
M9X/7E+hVuD0pslVV7uU9cqWwK48WKsLdLG/8RoRTTZC2fOk443fy/BnedIBLaax/z3HarUjjgcS
u2JJZfWRCy/WnJQdXp5NtnbHBUORDeV0sx9DgWvOIucz9sXkLHmZZ9Iu9nArw+3zrb2wApBEUwSn
g2EzIrHWvitcYYh/XoJ4yBHJjFcq69OMmj8zc1CuBb6kXfMj/5TfJNNgecBV6zdYtMM9YPo26nBH
6Kw5WAfMHyY9NqFwdQwaMh20i2VKb2js5XgnetOOR755TgB0GiKz5PNzv1pfcL0RGyj53rA9SXc6
kYd/OiLrC6abrPmWPGhOe8NCp46vhRBXlonAAjbpk/neLvs7z2Nn294mlLoQqPI3J0CXqqMkg3C4
2JjW1+47NVBuREHKbHPzpIliTYIv5Sk0U7ifEatBqnyzgZNKVgVftTjaA9TLJ3taOiYQBF8A8UmB
pX1N5yGA1t5TQlNxDU94c3AQj5v0Jfw5yRdJ/Gn7mAFBX3sS11ZjXIKiNKdvv5ZHqqax/veKemob
uElma5DMH+Fn6uSgAXCxRd2eyDlcXImXpip11u1A0RTm4uEgItYSgyN2y/JzQaCCKqCgiwFL9yNx
jTB3VZydssU/s4LbPCci33fBXsTNEIjouZtl0oyVGyAPNcUxQiBchn7PY0UN68xEoGKlsnCzrR63
pSzWrVl1Av8spT2G8jNxC0uPv7nV+4+KHPtHqC4V1LZwdQ/sMhyk7zqwaV+F2pb+JlTLUat6a3hP
FmnO9k07YZWNMvuVco9bfmkD1vYwTwrOhYnlgKHoytxcWKGP3aVWgSFxuEGdipnxTR7EYydRROob
fZa5g6bqt3/99WHI+rHj9dhDyHzfglspwqhCR1dsc7Q3Tdsgd1YnVMW9d0nKhs1NpI5CKqrfesJf
heFsVj2JzkpLg3xYlssFCJDnTCAfdSSQq5eHWe3EnrR6Il4C0qyg1ynObwDvAqXhpNTTiw7H2ZlW
xyxFtYLaV6EYK79OLVpUfAsLVckoRhptRQZBO03kKmDOc1bhEjOmhcnwB8ab5A1hXuRo+xQvgYou
BKb6QxZkW5snh2AlB60TnwV2CKzADqdtGfkpKhEu0kk3BsMPd9qcwvO6RCzvu3VqXY+8mxRUTneB
KfMsNLbUbhyI1TMsAFWQZbnKaeK2IzOBRxbLGy0xIZ8KFL2Auh4oxyMv3G0sb1pxOYOn6rdFu8Z9
vqxb/l8Jnd/Ws4xjMfRTV0cVpW+c4beUX9b5QqX9vktUxk6m/zPbo1aKgyrMlBH18adRl0F/sBx4
LuKYiwnLIhpIEImDN1/VMJybe1uiEuBsmibfqgdTO7Alo4UQokCqdUvDob7/dhQHDEfCTH4ZbB0E
S8FCO3RmCsyX5Xyrz/YDRUr43IS33YsZzhvjFOkf6WeqfsVBzxhlQnlxcEL4L40G44tm/FDf5xaN
WkVPxXysaHCTH9iuLKOruOMaf6Ad4HkpRSPLCX+PyDMWar+zM3ccqg0wg+es2oPpS3F45EJU8OGH
EZZlxWZR3eNVzw+bH0FiMyC3fiB+H8fl9oHQiG8d/UZ/GHcADMYeDmKuBKQGleTf7N7Y7yYSzGWJ
z5RPiAM0SOHyIQOJSkSWX8MxwOV0C+29eHboxaTr+ht1QSWB1cOiloeCgmIkpQbg8Q4dA5Ktk5so
eEPRHkiojXoyPHuW1vSkJICZqq3IEdnE5YXBxVd4/FcKR6EZaCHFC43b30sQuLmwL0DKdj029+go
2L6lOOQHrxoyXS8qNlly+v/Pgt5hAFs85/U/30+oo18N7PEgERj7Dt28enMvtVVIniPgdJQCpsuv
OI6WJNRleSkM/1Bp84+Pp0PBwVHvOG0hIOPnEIU1bFcwFlFwAGg72gQXEDicvlAvpIDmRYBrCUK+
z4pQe0rTlmvXCZZvbhuv/hle1tzii2hDwNFnArfCmxBGKmn/KH2xJvGMIJSdZB1O/XgMejEnoxHx
5i6zkt0UxAPh1nO8UFGU7q3eT9Zdsl4JJHXYbEADt5lY1+qaHfRPnsrqwfY83Zn8Q5RkeO//GPLo
VYDLKw+DyynMtXA4ZmfUrbm25IHa6HErPe+TEtV7mJvVhkMOn3C9TKpTi69huOVvDzj+QgBfTOcS
6pYU5OMzLHYj2LKpASY1BCqsodF0iHU/OaZ6j7WZKbGgB6FiQd7Hz5e2DGpP7yXbbanKtHAdfzrl
O2oAXpMG6Zd7jcfkQQC1GKvlXZN3iOkkzkIaleCWEEolC4OGkBGJPVjIT6dg1dp5z6S9aHzb1aGu
5clDsMNquJtf9zEidwrpIRKHAJUAynmjTFRJw/WfMxYDcbX3PuoZAjKWT9bvWoClPamnSNOF6ejB
1WdJTadq+uhhk8Eu9ZaEiWSiogbEaES0QEsGxL7TCk/5Kx1GpWQ0EOgYW9BtFfjhyI3xLvJRndY9
OFS53ZCkZATJsYcvTBHEv17ObGGiHlwztqvklZvSdMQhiB7ngGmSsD3BN9nLDJZr9TZ/+nqjNqr7
BC1iLLWmHP8tBFug3Z5UN3PPfDWE6ldcmE4wNBr0H+mdcahPQIeJu7F3cqObJgEbzpqFNRWduYuB
mejfvn39r+gXJTKAMBPtllqMAImCpfKyG29xstdjnRhC0GVDwWJ0HRbVxswrUz08p65A7LKRB1iF
avvost+Rth/rQOx6ooCi4NLsW882C5xeXByg09MlPyM4JTD52l8d1kCc858plWsRa+RlZBGZWFpG
XQwikz1ukdF94BFX8l1qtoI619zO7O78MNlHjTLEA69Dk1Etx1hX+FhJLH+veOIEVO2GflB2P/2K
ndFSWGNWMC4cijR7nMbppEo6OUF4dYNx8YGB00/ggbTFHthbTP7H5HPzb+APCms/d4qOO/I5kqR4
VGJnEIHC8+qafid1iubV1U9cvJS26ozcmV75CQ2U0675AMrXGYQbcwxZybgMUYB+921djVhHe2QB
WD4MtXfi7MaDvYcZ7WfKnjWe76SSovETCZKB5DHK837oh0+sMaAJHtBqMORvyyodZzJdAQSttnGD
h1Ivf7Xnf4qj8J9xo7iEA2V7hKFMm3RcdCrBzZlgAl5v33kPH+9aZgqlf6uDv3mPuJ8cMPWKe5Ij
ps9iVwwVZ/9Z+1EEr/zs17ptMORJ0vR5y+5BI47o6Uob/IUmgzFgmHSYY57GcaIk32XT2QafnmMT
/LigiLRQvvQIAzjss2bCUWmDF2NRJVN2/j/H5DKe3pSFVG7fZ8jzbrmVQE7Hsa9zM673al9Gwuna
XI3U2dhaEFj3DMJI246Is/pshQKWk3DpWsSvdaA8y/LdAd1Dsx1k7TThNgykuMhDtL6jq/FPwyqn
c71MTklhshNi+uUDgZfDUQOr5jDzNjqkQcd5QZlYIRivBbCflXPE1HwwxR9uCjyl1iXBCIg3GQO1
sgMG9y8ikY2bJRPGceBpr8Yky7NZZDkdm7pg/p56jVNKlXuBJr2yL/YqgzJH3KxzKSm1W/CQPzwY
j7781EbZn7WyXC0sgX/WRIKEK6IRsBln8rSO/Lkk2S/9Panu3WqXEgAn9tVkQ7ukkHZJ2myX19ev
vza6gybW0lLV859Q2r67OqQEUC66xkKJ6bryKja9gd6kyeJcAbohIQrwZDkTwGg9bPFXx01uhKyY
scASOJmi14m88dfU4g2SU4McyXWze1Hwj92NgHrUAg5SFHyOqbVs5ovuKuFR3HwhpvvVr9tsvtpv
FjXY4yTNdUiYjrwZOiQ9ZRBSdCTs/KxFBbsCDSdX1DILw6kg2zczJhdfYwDMcG/pfcGpnuK8KG4p
ty4p4DW9IXxZ5hzUQV0rqGz5HY7Zs3q+6x7xZuDPJf8SnjIxInuBRy0oX0p4pRkqbYNNODdua/IA
HYzb0SyyiNQ/yJ+M16gGQrYhuioRvzZm6GFk4DJQbsjZYMr48s3xH7b7IZD8fE73a0tpA1+s51DP
gAgeDukpRjlZmRLCkHTM91kaUQV2zhDkURI7b4IbdDQnD1v/JGZVLNwbWF77XFSkNV4iplnoxLzU
7RAUTBEkljIdlb9dDCKsRiWG/cy1enSe0tpXpIDfeAZWbDs5iP5npWRB0/oHXB+qblurGWwULcQh
XIc6vbbL0Ao2EWeV6V88L5m/AfT6Z2v/7440pHTxk+MUXeGPl7v8gMDSFU+qCoFoSkLQImoM24/8
71tFSbwjLG7wlxLnm8ht1fql7w6s0IYPZB28DCsfct0BN9mNxwnJTJQJKh2HBH77OWBtkiqSwFxG
5zXcoOFoLfQK4ggTKWHVzTp6Coaoz7ToQMqa9r2AmOtkwExJrz/VWTqnZPPt9q6+FB35GhqLKJk/
KmLAoYIaCujk0whhAraEiBLJsHay9pceDVHs0Pvf0xPe6QfjmqXQwteB2bp6bCQEJFSnaCicCZMM
LUClgNX6uPco526Wq5qw0iccUrgknx14AWaNrLqvNdhMVwzZOVIhQ21045yeYa8vX+TMdScqHnHQ
T5oorPDaY6x5JIXkoKaXShmILX/XUscj/PLO9jFHAHK52FS4OiRf7zbLCbezZYJD0Ru7tafndP/j
RkpCIUTrMln/AT2zmi1ohCPLI/lYEdNv3tWtb5Yw9dOii8xqtleoG7+XntrPm6oPJUjxLA1gmEeY
bq4jw6ozLVbnkm0YMYgKrHSt8s2WZAd6yEMSYzYP2KFDUT3Gg0XCIemDBXFMZwPl6ur8qN1YQu6d
JXVwMppOM7UbBmBZWpI7e2lFTh1maWC0ywRkvJkMWGBtWHcnL+a4sQNzl0huB8iVOJzrq+Aj4GTF
lmumB73DhhsER4kARjLnzEk64VCMPn4mIBJRv6qhdZSkvLJnN3K/draJBSYf4domIxW9ig8jNcWn
GpJQL8lPvG6v5I5qUS4MDYSVILkoxGRLumIREY/VUOJuTy9YiRayjJXC5OxX7gZGcEzuPMs28lKs
3jAyGALP7x/kGsQwrRe/3yRnvWELFKjoPl9XfHK3lIWWIHPdceEVzHWQ5AaKC/suIwKoRRJME3me
g8Q5UckG1N4JW1Lw5CZFJU4U/cRd67Q0nObSLugRl1bT2A9B5iAAXdbN7YvkONgRg18bv5uYnx4O
Xy1NVzT4VuYUCRI3fmpkjWBfq5E3qp2WDeyxnh81A0nBwfdvuEOtRXXiNhiJVMvq/wYRYoT1UR7W
Z/f2ozrAdChl2XR2lS6Zap3WZJmqsuJNF4fbgjww1XE27MEYGsYuChsO2M3gn7rTJXthQpCTwxqH
S0cxrzEXW0FMCK02XwzD/WbcOJTguzp0gpUBX2ysZ60kt8LWVu0gt6BpsVYYfkDjOuEeEogdyDyv
4pDotc/w+ufoaaKbbYakZdUzjxU8brsV7Ct63I5Ui7lRb2MBw8eAJoQMFCgai7x90uaBRej2qPUt
LeMg6PxLJLqyl9ICbbFA5hLGFxdL38uIF0UUiTcqsKgGB0++mawF0Epir3CJt3dtcrmZ4HVV1WWI
f0kesgk2/n1byrxxInwuYimp6VmHs8pRpxmVJY8kdGSWUObR6ZVNC40O5z8ySIzmVytolAX/TvFF
XoewF4OLFlu36nCeFPXJZjM6wwS032XQO6vADIEoaAj/ZVhVuLvKjTdAO9x6w3ITqdBH5f0ah9Qd
7O+0C+sKsZpOjfd/VWdUXzxNqGftOCHT32SypR0B7/sBmjEMvg7dySGhIc9w7u77Mg2jWVuL1h0F
t16ddUnT9cjpCtwxjPT2Tn4Q2NMjowK4omS+zpfLwwvvluSOFyhkZxg8XJ+n+qOlfslewug5OcBV
cvOpuD+Qtu+CDHoevEwDDzknynzjRGbml09Lvo8U26QRooQ1NdzklAV2X1YFBFDwIoBtwnDPCV+u
fSoX8oBnFPdPz8eg8W8D1gx9QiiAT5DmbFYbueFIsxB0ViDCaiNl0FDm6QtTWCdcJ7h5bwh844vL
2qDeoXs+ar7t4oMKq6wJB3mkGnztrt2nfrEO0Y3QiwR5KYd5EsB11uDU33r8ZSLQVNJ1lnBzVtGg
63NZRug4bgo9KtQiW4Qk3CJw01I/jkuczJVFykOMsXl2hCcP7BmBkejLmTgxYixgItq9QX3FSknR
3L5XwEYPEcddp0exF8bmCHNzDmddYCNlyeIHgAal/oI6dG5xquyKbw1y9sBwH6A/TfpA+sgXYgty
EYGH+lg6EFoKvTMwgzmxZP8Y3iOVw5Vc+v+yPhmpkxTw8AcPMQkk0Uv5c1EhdNzVhncTEa1WXUST
S6v4Bx83y1Mvhzh1KIAeIMBEoVDjP4+57QFt1xEE+khf3uMAX5G9nS7I8vmcgQZc4UzN23l8Youy
O4HxTP3jd5v77cHef7VZRQXxzLAxa9SH8vmS+XWK5f6X7J4OTHoehKxvJNfAAp+phWxRVMtmwI+t
xvMvZIrDZqN83ApgdPkuNijuClS8xAbresBfK4Cvmh1nYjQx0aSI4gIi1xBj5RNX5YzEhUTyVl1u
FH5hdAMLhHSXlD5JYJFGuVLymqmeGNxxSCRV8V0+Bw6VY+PHd/I8AJrwumGYoHSrd5Zgmm7b59Tv
juXdRbSnlHwmA90vHSvn0EJLuzwTWOHML3kQXgeY2Z1iK39/IXsZdjlf4ET0WhEaRdVylS8XG5Gf
yUscMs8nt21lW9vlKD2zaM1NrUAcviVjWe5lzKa6G6gZvNR1F62/kMyajsvZw+bUOIY7m1fg+MCM
ELwtT2cJWXOEI+wotK7mI/eJSEdqFpTxW561r8/67G31srca36FGd6aFaLy1VIJJ4nrkCaiuUKdV
KUun9uCgRiYkDqp4h4SDI4myRvrgaSNM9nWG0Vo+oXqWGCx2gFUhaUcSXfXH0H0301xaAwJxH6QS
e9WVELZ4fqRSz65OLeUE3xSN9pPZPPuEwvdoaLBxrh/DZza2ds2JaN7hfH4Q5l2kEF3SPfabSktj
j8oFzB2WQwCXdtCzr/XABqz/8qs5Hwq+vXj0au/VRmDoBcpRhYIKVGQTH9mho0qInS6LBZI1EceV
SP1eF3aR9Nc80i0OqAy9Oh34m4arA958eGtUgcYXXcoS67h6USuL7pYrLk4B/1B0NBzp+uKTmaLy
Kc5fTen++B+zHMEnoI7d0huUGJZWU06EIuAMVrUbUQ4mF3fHCmNqQrKBDgbfgM29At+upFPC4Hrq
2KRiIohOD5YwxHEGh2ntHArVF1H1mNW8zkbVlMNV+6gcibBMd+TrgFsCtrgU8BzaVB39S9URdZwr
lZkTv3JE0rX59kSseWtCAbH47I66X+TYHu8Ai24bY/0eX3lRwxLtHL50AQnsKSsIhN9jNXyV1TqE
4miSwdvxC0/RQmGaeZbcmtr28dGR/FWhOKfMgkPQgewgOMhX5lr58j5WQGkjsiwQ6xLv4yK9zdL1
ajZHBYNSRB3/hBZyMkPLekLNlCy2ixWu8xjv3x4Z824WGr/yfzHtJWcZNOC1zSPxG2jmfCBQNWzz
Jy9UDtmK4rNLtIfjTwrZxi+d3E6gYYdebfvTIfqcOwO1pB4ot9rSKoLAQGvEvljIbkFZwxIaA4kU
1ZFmuzDIG6IHSfucgsKxUu0ikQjAw24kjDyREJzSzosWdRHB1aTHKJWTF7Hl/Sdg9ziPTcAz20Hu
++bjWxl6sSIY0EB9yPkQq0dFQ27br+T/E+eGYJ4HD4tHRfod7hT7pDT49tCQA1OuIOGWc5qqYRHH
mmeTrCH08xSeZMfSSlK47tr3ZQOZrb244DDDuA+zBY+I0tU+k4ySHsp92u9WKyms5QUSmUpY9U4T
kkMmFFBT/UkgdKzhYOC06PJrynmzW8kpRbjfQNvWmlb/2lrbY7J7M/Fs2/Vo61vnjpN+vuAKQFRM
EzXFP9GGf8l2vnro2guN1Ch/tn0nYifH+ned+iiORE+j/o6dznYORA7tj/edWO45mv9fq9jbKBx9
97/yT4F69C9ISMoGi7HTnVj0Aa5MCNXaXVGG5YEdzY2CvlQNTZP+Ze0RqvxpJ6p+UpdIPZnmUxh/
ZJW7psUQMd8kNOcVj2PdyNSl6Ynum/3kvvA/Z2NRRcV/mb79uh4VZRpo96ZTwjsLvMie0up+/9Y9
QGkY46ki/qHro2nErK/BMnq7KZUW0gLTLhDveqB/zQi5SR/uewEtZuXXtgZze18udrUN3uclns4s
2bR1MbyjkI45hP5V4H0JLsg7KlNTRWLr5MjZSuLvrLklJqeY2/GwTZ3Po8GLfAqDm1f9nDuAL88x
h/4hgecLnHcZUaFFSQaEGLDlZROVjjxUiwJMZSWdGG6KcAyxYHMuajawNqRe7RuMKIAYwJ6n+7Ro
in3AOET3G9C1jJpTj8vuC0KPDYdvaFobw0+OlfV7IL2VomOlkzWfaAWINhRRQVJBEra2D37qIltU
y+odB4lMVmm4Dk9cR7ZcByM76rW5/eaR2cDE7LvjsTg8JE0NxKj0G5+mpkEm+ds+Ny/Ii610YrOH
gaTgelkj6CBO0L4nlPdfa9IWCumtpF9yw5+fzsSUT60Rk0824tKnA1+VFzpJZsbRxuYJHXk1RKeq
jgMBfzbNJDr0kNsVm3fTbS4QUMlcGU5+yghVvXa2hmqlrcQHg23Y9sHGhNG5+sYoV6ElOVV9AcQZ
gwjH6feL1le6TdsY0OnG8VFQDngLyCRn25fMCYip9ywfhiJM9jSbKaDSR4dqZf4z9Oq6LlgPGUNb
OksRIgsVoCd29MQUPjBl7/Qt9KDlMNUSHoCsZ8lLHzLVgCcQIuFVGyRz5AEMIKzhYSU0riqpPuRx
7XAxRIACH66fd3udzz0dksZW5SUgtLZ++oMaNzPd0ACvqaw8A8Le3Famsv1zDMt2/U/0JWcFCWed
INbFaO81Wr15U/Fs3gzPHCqT34JRuTLM5Pn+Gd+aHn4jNnYxPw1utP0qPQPWGGkO4eAUd7cfwnvG
mUsqjUZgztIb9ykA/4uoUN3cs6VtUpN6924gqjKPQb7OgMh9XoCjd96Dpg09Ycd9t7a474zpmSOO
rbrN149vxBDcmbo34qR0eiha55vLnpquK76tNGrujp/PwClo/KwtbKgn8BpDwK7rmSLcS1cOX6kr
lXW4bvNmmhTbYjn0yC0wByL+qAhN4CIVr+5hSmsi4uLPBPE6+FmrxKOlf0s5IkIFAWSlwBJIvAcw
nncIjAdjDPVFdjHQmcp6kxKfN8k3IGq9GEjKYYYb7I4J7VRbEyMxm2T/Eq4lzz2CY0CgsSKEODeS
B5A9XCm3VPbebF0TknqIhuC0WlzUPahY2UtfK1ETuTg6zGyvYD/AfOWyYyCz5y30Er7YjVR5NFXb
L9vdBEjCqGBZV/sP8pLSkIJFRTtnY32bu3X8wbGZZScoVLhTGMm2ZNS0ya3WCYeB14Sd9i0rYaTA
48mV7EaL74N2VfbIl4gQlUhrwnr4CRhs2Ur0pUlqjvkUpw+etOCl4f8IgkD3GL7qYAfqOqx8TyTU
yqolqB+B37q5TZk2vPH2JhoE8BrjlDarvocdD1h3gWQBharBYvYXFd8B9AQ3pdEpmWpesxNARaUB
0CxWDILRwAZpyjVTFQHwKnuRqgZHHizfc4/UQhqHALIHHQC8ThYK401PsVTiyAl0VeuIvhWSeiGc
9OJqC1G4F7j+2F0YtySDqNNMEoN9N8wfuiiZMV8rvCRU6ZKYOlQsQN6d/ZOEZglaS+LZ8KtTK/gm
6bLWRwyJzZ/mwOnzpBp4RM9vOPhEw12gC6gzckJpfL8/mnyI6pBRMQ3NqOLCeHbuXhEiNNWGuqXQ
/gfYguE2GdF7f7igRev3pFcZwehqdFkb+hv1tuCKG2SodVGBo5CvUBnU4apvmwD3OjYmiobPvcw/
ztO7x6ik6vBc6SyuDdnL1fRNlDDFCf6JRepLxx62wXAr64u/igs87EbrEQ80SoaRkEY4Inx3OB8D
Kah2Tz+QDp2EChIypHc5Sfy9ErcpDhm0iLt953xx8B1S8gul/QK//gCjkVtqlB6WoDvbMtVteSA3
/QLcS+9GsNSxERR7SPYy5S2Y14YKh4YIMXAgeprLNm8+XoqNdmgXQC0k8+zSXfHQZrDuImhXwUAS
6uesFd+QmSTgIkmiQSitEHHZgc/vw+IAENU7Zwg3N0lZvsLKqKXIEyiAhChZ5BvFtFonIrsmD59B
3fvuAT7M6GUWOHOIvwsL204DeFWaXbhMnoxdnwubybxjOsyQrL+O/Vto/nQ5flunE57Zadw76PY6
gmR+qnF/vaCPwhgWZ3BKgBncuu5nLgeXBhACDUg+pL5ZDyyTeMUy1hN4Pv/IDqsApq5tYgDvvXh6
mjP5u/ghxXsxGESy4gSWiqDMgqKfsjOncwXfIWy0QQ1u5kVgDA5TnU5QFOUjS6K3fw2NzwO1g51p
uzlQO1Z7R5B4O6QX0KFttVPXqut5Y0at5yqebRRTg5jhvEofoDv1o8sjPI51tcv4TnCOKpOUkKUg
ZZN6L2A5sSQkwUPX20HTgc5O0sQZnAa8vPbI+bMt17vgb6jLRsns0iYtYspfS2nyQ5fIu2Rpftzp
gX2LkCqVneXkXHfsLtL7qfPf3ho+Abqy9QDFJfSFtuyoBPZxCPYWJKqj3/EjTRr2PGDkDA3OzrDZ
onPuxHHvXt/Hv6tFOq6FdbB0FV/6vmlUugEQ+lv/N0JZs8f6/H7+QCPuTRf/h5+45RZ7KI4t7rzc
Ay6LifpGTfSRlbtlX1+oi/SqXsDEMxDxBz/WJpTr2GoVsNndJLX4SKavXTa/dbbQ3qOzWIdl74tB
obab7TiCK812WmfMMyiykKLJlb9zo7I7c+kTXyZKjPE23UmRvk8tEj4ozhf/vdC+fBqNPJJ7JlQv
OXeGdmZL0tmVsWkAw3lZQNeq1VHCOYBUNlDZOAF8qedt1zFZ98pysXDOZCHSwrzBZRvE9r2cnkLb
LvN3ETUmQ3nrAYYm9Dog2X5knJh6uvz44V0DJfddYqh9rdozeB5lZbgW7bA2tp4aewzEUbdyZKmx
w+xRCnphRpgW51FrfScsCh2sXmYgGGMIFUPhicEWvhJm2pP3qEqthrX4QysRfv9pnKf822f9u24A
rC0guY2kvO5AG5bh2PKMLwr/PDsikX8CaPN1d4Y5bwLawZNpqWPOAVl0B/64KqKX5RzjuyR77s7H
MwHAKD7yByjiCSS8rJ6XJ/1xJ+hUiwrLaYVrAyzPl1q2uUkvuTv6aMk49lpP/vpqms1Rgd3VXi1K
wznXs0YD0PqtwB0enLHYgqKNKoGTz/BWwO46zCvoC9ninwKmQjQrA94fpNSF+TOP5MoKp0z7n3Bi
FRjJqyBWRiR9zNa6lPeiT0jngqZ3E/YJpxTr/ZBtzPeh7UEBY9w6gfaNNU8SE1a0rzPS6JpvDH+E
oxFYVUtIY1uOl5t3L74p+izRm9DRrm03b7peX4bGBuUkP5oaMMkzvzzo2JK0iiaCEaiu1mtvhjOH
QZLwmCE4Nbzd3lv2JYnbNHu8nfznv1mCTvHrB0d8iNlt8QQxdKjZn0PBzreSbb/XvPzgGTx5XiY0
iBS6XckhOWjGdxAX3SlGbn4pcJor+tLyfmQnVGeSVrkdSx5wi22PLsCJhCWMCuAQd/gEJyMpbmP8
flBmZdwsIkiG4h0jRpkn6+dFh2v0+OIuUyHris6plGPr/CCRWcxo8uUOtoNDHq1ILzyLb44XlAu9
YlJ2Hh5eC137W7Mf9OjFczsAiVoq9P1s3ifb3LCr+QhX/d8296g0J1JHMpY04n1PAPm+itLcVfCa
RBBPIzw/y/pXkoZ8FFOAOcmBPBGpqTyb0PZN3ZSJz7a8ro1jpJrhiYTUlOMdWtlrL3ZBX7CEllZ4
xPlxr9C3T5Dxh+rDi9OYgD82vVI8q0jPNf7iEpL43/Ah0hXtMuwKctxidjm18CIqbWTEWDYCzzSd
+M/QqTkDSvLPzNNDA+GfAlOFU1ciHwwjS7jV/w6/krSRY8DrQatpDxV6psKqVZDUpSYVbVfRmiSL
yHS9PZYQhvQ5I+cKxQPy3spcaVrQTPo84LNTw78zfbejc+kPIUfhm4MznMsMwaatMBKurFPapvX6
f3R/FtnYgDcxWMuKp9BG6ToUq2DaJHZxkm5guNXHxkjj0773s/TcP/2Aq6m2e+9D4YS9XhTRGA0j
nKai2sixR95mOg7EU99BULp7uOfAObs+mtEJKztMIv2lDydWwOuCSZFEvXwrU4t8Ik8WFLH7F7W9
71XRh9vGYa/uh/osR1inru0SNJ7fQup+VsEvdbx9yHnLNtrwxTiljbD5uzwzmLy+ngPDWUyzx52B
pG0QgOAfu8tK5wfLGo+63BITkd4Ssqn4M/LN3LS7KsH7e6m3irIdST/Fw4rr2TXSaus1fAhOFxkk
OFtFV7XcJU6IXh8c40aLgRU/7fhMwXOH1IzmxxiDw4IM94Et47HV4J44YI0klCdSL0TYlIFfFXOv
v67+hf96VJ+uQf9bpHb7mGFFCQIxOd5TPhl/O+khPZLuQEaTtqe/T717u5e0dvZYgf5r4P4QWwn8
1Ggn+xp0ZxDkjlLSKmOJboPkokV/SjmjkGGNE1I+UIN9CpaTvwYt4krDxdbGmX79LqfMAr0aQdtR
HPR7YDdVWpMpAir5j0cVA5hg/+v/Gh6vWn3fKLkBD9u+nQN1r9pNgA1ldfOgNA5UEW5x25RePArT
ThVr0c7Sx1hNtv8f5o5+yiJt6Rl9EKOlSWCuUt6VKlEXKlU4YqlsGdEoceEsJ90mTbiPsZNRk5qf
fT9rGPDzzJbJHhxSLlYlZ60Tcm9EDAuxemwcUPehPormk5uXDoVVPW/T3ZGwEzsKT+vSvkR+sdFb
UglvxHe27w17/NtbyqYmJjrfLuPoDKOX5j85d23Y7h/dAikQ+TeH2405d6PmFCVftILjp4coL5e0
fEj5YeVavp5lLSwFEW1wUKPH5aFWmgGlf0izoG8LhUZ1PPnRKJcqVK1cljkPmT5UclqFlTdn1cZA
iw5F18QymeNzKpHGNt+P1eG/rHkaN5V1ifGFCN+1ONDLbQ7WxIvJhszGx3Rgr6av/+82G3InmKca
WuntqWJPqh25bQbz+1vemQepk0/VJmy6iuIbjh+33iFq70pMQ4ZCd8E02w5GJBARoKuOiSNeHFQ7
2SGze8Zwl3E7t75BdC79XkI03irg3hsNubOcRMzZs57YrRI8WaL52vX9GxRZEohe/Y7+EsabfezK
88dAdS1B9zyd1hLKNqiAq+d4CJjUcX3tPJBWqkmqtlkyMGngRw6+of9M9BZ/SPvo4P/b1/zwnLYV
TWVuDAbhKJV8JuWDvr2pZ9B4hZBYZoYO45pSGUfd+gpoIn5Mp95aP+Sh5xQMzq1qJufgPVcY2tZ0
5nT3bKpMTsy9yjCZmtlAvcnNEkTH/5MXmfc9pmVkvOaQQW3truQ1hGxKpbOQkpzjpKH5djZYYy3u
0LRE2EgeknU+m4AuEP3B/bY64VN06xvOh8ZKIwJoUora6AXc2zBsTlH6T0/IGZJXqLaVjeAAPEgM
KoXCipa7mBUI0vPbzXWxf79b7jF/UVBBaegFT7D9uFC3wkh4rYThCQcUqI/q8o0bWe2PPy42zwHL
WqxyZRnVlVh4nuHaDqKvY8dpbqEoncWmhD8oZmKb+x7Ey37BMCw41TwQreTz5mujCt1Jj4elffVl
goKOa4PHJx8mEn2LqWn2IInHxggyw1umCs/PvTxXKFjFwECim2lLwjZ5iOJYtjwRyZISupj1oQJG
QNQpheBNCZICx/c9KksyGHJ6ZeGTWUMLx/JhdNlcgJb6v5RsKbfO2pjbTJJnunnzaE9L4r6uhImX
iR8pklN+b/ckj6t+KHKfwDann8qAWymD+uloUBRw3jtCKlh9q6kiQpiCMeTWSFJiLT6uuS5AlqCK
cr7xABoIi1bkhQew/F26Cu7gD0o1HKw0ieNqlWAptH0bzQsRKMBjU3eg9E6LMETqPjPT/J5xeXnK
rrg3b2IXW+fwCqCecE882VevmZdUpOKCBskVdPsbEwoJjSWYl1HAdWeItkrLuEMnNSYu+TigwNQJ
7xR6iC6VYFkolVJkZnm6WKEwTB92qYMzD2ufMzWB2/OmporQePtYuGK1o8MM0uU7cTuY6xuZmkZg
65WzyNxjpmSZXtrvSQseJ3NoXEE84WUeQPzFr4aW4eyUnjQIGq3Zkw5SV503l2sIW+N6QcBVXyj6
FWKAEdDPuCz2AwQ1X+uT3joRD4Xwgvobrs1Qtb3Qo0vWGj6YErFR5A3Qymd+JH0/F+vLC9Aer+1k
jzLWe6rGPD1Wtoz+tJaPVctMY17ET+t725bLHMJ5IC96NUxLHtYz5gbv6yEcK2Nwn0apjpkabS91
bRUH12KyRvxG7kmkGIxrJEhXuHdM7qjFJ1p5YrC8Q/yfffr6LK/BiMyubMc2WXe4UrGEApPC2FE0
/YNtC7rYw5rw+uH4w2cSbkLXna72JYCggy+67Iijz5D6cQ2kGv9PKA7riSuAxUTVy2t/rLJ//FTy
/hxdjCdQlYhOsp6eZXvu5Diiu/RUOxfCJxvuvpwR29l7AiSfd0AqQMPXeA5+YAl39YfQFvDzr8ij
2z28FHTBW0UvKmi/zrreSSN7D/lqSfINnPg97UZpmgtgPOeNMgKXNIqJ/uP5mEX3iK9bkNkTq7JU
nCYN+5nPLVV0Ws7Ciywi8eO4iASDXsd5ZQCnPlLVFNoXkLQmOVOhZbemLs4AfLVB2TslMOUb1o/4
Y1/NivPN9vkitgXOPxqB2Ht6AaGgL0toRmsOlKqEAhZXYbTk//13+bl2QQ4+HGaswGZvVzPTl3yK
bklbR0qSH4ZYwmNd2T1Z75mYNurebRMc5k0RsbnYauAFLDLSZUmltJI3fIZD9l7tUIuegkfotc3V
0J0zdEslHBDKlVU2sc+YWOHIkVWgBGnx8Zz85dVwWXOnaJGWQPjbWPUL+ZwcB5QaA4C9r1Kva5ui
x4pngXE24kZY+YNJa6asZQYOPAxMHs/vGW11LRhHqWy3DNY2nx4tI/OYjbpfiIJ0stZ+ks4ts+0w
IrU+NjxKt587q4dYMrwzJfAPm+DX+5GlZ4YyHrvfJyiJvIinq/4pKp6nhy83RbWQvvTmstahInGd
iohi+VAjdTduhHhJC4YO+rmS7htATb5EUY9Uq6AxDkEITl17QPSiebrUic8Hj/QXuAp5DW77DYvm
uR+CrVrM5y7XH2eH8/XfKzYDHNXNnMLswGicm3EitdwlAHFXum9Gc2Avl07pE9xtvjb6PCCILbBI
kkQmZvYRJEqXTLe1hAkXklDkgDu3ZgDmqVgVB+bNdYDx9+AkGTJHz4RgN4juokabGshFNNBHh+3p
X4WJff/jawmX0gin8Z6aT7TRqS6EtqJY5qVGeyG1xT/UiBDLajMT3007uiMzLox86zNq5YeQXT7u
/JH+zWFaI2YselYzcznq4S3eN9SOSqAQtZH6uln27RH3kNOrgmktYtMIGC3BKlYCV83MdbtkRvan
SNadCnjEf4yopjSxeYrLgMAwDq416eK39jfJ/Wb56o0qoSfHhN2+iZDjIy2RoUCiANIJdhZBf5i1
fp57sEd/MbqaHAzciz9TCiiBu3xuDB7PRV1tcVjlrVaQTE4+HkCJRpkYaDwwBarMSz9LeGhv2DWb
Fm1skgvfOgMU074fgvVZF1omsnq6OwqiBHiMIn5A3R/g7CLeuSD9oOTrRei9GHdpP4UX4w56GXRV
HWicQi8/2zLuoO8lutNDYUwzLG7i0MJee3PS8evsNENbx6kgDFsyYNfUofqyxTorrWhA7PU32FC1
HO5owdqlpg+H3fVB2CK8BjkkVAX/+atkZxQ3duDWznW8E42AZbxiZGdBGySzMtZGPHleHS6EbX0u
vIPfSA6rJYjQJBfneLURFXTbGPchayYUy2sNpn42LxFF9KYMpPdy5grKI7HPn+/Lmiu7+2P1wmaR
wjZIrbJGItzBi87HUFmWbZIm2s+JtXynK1YSs2lJixgxGmALS+Od7CZWF6KB3EvzebeLXN8bmBe1
yZSnvg5iseLpsWdjAS3yuVTStprUcm+1HKwgvMFfGeTs08nIoPd7yt+u+vJAv/2RkMjyMCj5AnNG
5qoWPDl3KB+KFflT2hai1ewY5XmkbNlyvHEo63yoIAXXhMhZSke073ucb21H5RiA4mHho053Q3vO
IXCXj+uFG0gx26xqM2TVopG9I/R6Zyt+h94tf8m9UgcXDPIrrd1f5BEHK5hWhlRvgZz+jmGaxTFd
X/vh9sl990P9oJnSN8FcOg7OPMPNyGGRNzbuXRNEeobvAmb0zDaXsId7OXfcqfnFVoquveflBw8b
/5LbkBgSgmykY6aEzoUnDWjc2TWjYQBqE2pU5O/eR2mz43hpqXWsp3+kBubbloc6DOLTX6F8XmME
V5Crg0QlGIamZgX2map5UX3Ihzj5Rmsbup+iy0+gPUNHQesOg1AM3p7zonT7wASivRG6742IJfdT
VKhBidfkhr4YNBGPsBQm4iWFI3CQ60WYf4wvhKje6dlqI6eW2Z4HFagJ4+JJiwfYkcZ7EbFIduf8
ZrMKgR9x33aFca6cd1j/cf3N0uDrWM+qABAV5fm8w/s0M+152B91Ugv4FhoPouRWiOAaWi4SN3fI
Jrj4dIiYmcs6DxQnbXYhfAEYOVQvutYPXhIT1P6SS8NwsECvz0dT0sv0tPxuWz+hhiP7QFM6r2GD
vj/qRFuUJkEilQp6ukyvGWsAu/b1GKyCWL4S+/ntZtAxNK8Usb+XXoPQ3XjsgHfZ07Rj+0Ly0Kzm
vUWEE/0T6c5BP4zeMIihmmgcEPH/NersBZgGWwESguQyKOo4ZkfvYn/m6x8DvPTy2Wcb7m3UiYIl
4YYV4iNys9QIE6Qd+bmgpwNAIltzpiRjbekrI+V3iKXRQJAGgjoD3ZR1em5oEBJUdH6W1R1nk6uZ
luWzvUCi3bTwyoifsUr3kc46aLEmJQdQ/ymTEJF7eDweAUdRmwdRO2/ypVBnI/oIHNB3TP87LpXl
DcwRk57IeCZW803fm5S7J+zfuQHFp5Xx4wqkZgm5lmzMHkMuAg9FuAjaJkQsQIvKBOhlPvSR9yRk
dzfTMFe0QkJSz4bLKLXP8duAiRukC3FS/zbq7Iz1BqGghGMEhFYcg9bqYbquyK9mUdvMnT2G+Mbs
MzzMRwHYUkc234vFodEsxroVwkYpP88q966yeJ1BQaKi1m86CYXKWN+XNeDzJCCF911FkieIK6Z4
ILpvL7DReMa9mOiujmqo7GfYL1gwg35P2BxobD4XgI/YxjNLMpEhkmlMM7JbMW2NI52J0el3/Bax
ufGlHNMqpernJYVbPYkSk68gAcctFMDhYICmmYXpuWVrXWGGWKj67qww1WnKCGyWdQHODBHp61Tb
8CY2crYD8ZoUkxZUpEQIr5l2rjAMoz1C4LzRaS9JtIJA/BE/4CKisl/wJePqFLyNPiaqnZ6homg1
39EUs+X9L07hczLeEQf6GBp6mIPMGRCSqYX43PNzYW5OIMQjxBqUi/HtHD1sUMxKaYRvWOrz2ikc
6/fejXZtz57/Xt+GMnS2LCpKHdtTW4XjidwLtK7A0sVSvfnG//MSX6QzRO6y4cDGDgEt8ee7Jk6a
1P2D23L85kbEImprOsRWN10F3VpTCatlVeJ3wwVzSZc4Eu++m4l18dEMKSqUV84GOPBSHHrI9wa3
WxMEIgyHuaCNG1+T3seBvzTTvFD/wOPUTYLILNOutndDGyS+QpkWntwRbSftGuLawHvKkCgBrHld
Q9lESC24KYN4Agd5x3I9Jbrweq/EfutGQ0Qj2VGuk/b74rPz7lLzfrMoWxLT1X+hT8Gl1d1hooqZ
3m01+rxWpWaOTyoYCAUI3MTpBVnRPNyNCRFwQ4WbFCGTHfxd7fsCj+mrWCIXt2FrrHSzFzQCw8Yp
juGIsBpiA+yjkYY8yTvSpt90nI22rntPL4uITOl2GQpf5DvdIGh09EUWCXvUuESqiMd6JJKlR1pG
U4WmzpO61yrNBdBAs//it7Nv4l9quwy8NIO6iCPdsZFE4zhLLeJLHFOy3DYU861wBhV0Dr7bzRxo
FX2+PgOqrNjbZyGHvn3lo4f/KYip2VPrSAVGK//pAY6Btl7WSqFCgys2/xY/zRpzL8YR6EwE1mde
qPg52D0jRS+01OmfneKJ4dg7ejAiuEDoft7C9Sw0XAaFmzDESvuyxQMxyUmYfNNys2F/Qtu6U+DI
WoJyAY0uJpLY738UNOsQyFBngzZGqQ4KZPGkowyybyrQW7wfHwFa2lBzUJLfZEs51jPgXSUGxx6q
qZ45WlZHXWTI0VqKgurnQVTWao4/VurGKnwnUJdDj0nVfFh8SYdD64zlnQlw0eeFep2h7g1R2wtw
OGxBNOjgFLjLhT9fqRX7SRwKaaWB6Gqmc8qoE34bckXNyKi3rNQUyPA0oLwdO7zM9/3xJ9ct//FM
6PVRS72mUU439zbYie9wWvXaLKlnrjbdTZu97/uTXZryWVEB376x5SwVooZtcssiDVAgPY2UkwZT
47ATPeTXBRycnsIvJR6evP/lFD8g4dD+O9MMAMi+i0kj7sP4wQD1ifiQ6r/1mLIlO0SqU/E14B1e
D6jG4kz18soDjtCQZJFfn7+7LOnT9Zvi2TlJMYz94EpfM8VMcpY/7n/fBeIlzjzb1dtE8ZFL2P/L
juE/zEBV9pyrscJ/oHI1em3DSsmLq7tSQsdVmNHxb2OrwK2uB2XYdgu6Do47xc1mOR6OWnpbaVRM
vJU16FsgTIHdXXHtf/oefJzYZ+t79DEhvKynUvG0RCYpqO/CVolpqcY2WUOkkAybAnks43FOWjLu
UvPwVg8g89m8+uZYn5Qfw+DnM9fZx1+S9i8ETzbhWxbKpO1gjLranDdSy/INPzKyQUqqpAfKcbd0
x8gTZuhYPUpMCMpN14IRcSYPt4a6Uj6V1TUSDKB41mVgONE2C8KrnCfTDmQbGds95usgGdL7X3Hu
oIjt8gGLLwmEf5x2RerIjh7a4VjIIk4esVpog2N33iYZrYsBnL+obdBCDEY6dXiJn27itnlTXviT
Pu/J6lXILjX1sD2Atsj731mETItq7opElaSakUQJ4iDkDEuMQMcczhLhSDI7LO3w7b4xbOHXVVL/
dh2ECB+SY1uBz8Olw2eS7WJIcZDZyuX2F03JWAGEkh7H7YEFq5gaGeu1Gqr2bz8v4tKwWlFexHJi
x4KOSzBbu42vAYFal8hn5vNBAuvEArsvuL6taweoCb0aWJP2KfYfinx3JXEln/H+oGZoIRwpfia3
FLC4T1dkQxqHEaEAF6NHeN58e5MODo/z9LDlMyZBOb8iL+h/4+jeM04CEqBBD3PJyBmf2nxegUst
cXMG7vQpjXn66tyb/Pof4WHetaYvYX+FVDSMrtJ+a4CRQBEGXelRH0u6letXMzlaEf7sqjnMvBbr
OyVzeWK5kSJeF6urvjD/jHRvW5ZDRd91auMMg4+FwyJ3IMBuHcf6Vs1d5LQacntAI2W03wYXpQMx
yspdRtjdDoHj9ZvekUHxUcxyqfoQESZ59rJvl8b9KCQ31QveusnCfgOMpjEMZlKarsOk2HJsGuOR
DobwXkLcCXsZwJ5qr4RQRN5MJ5Js6L9tl5UgiVr2S/6tNmok02SLrEz1EDsLrrPDk+xZq/FfWnhp
WlSTrcumJBwi+WPuKb/wBedBZyXDOw5PXY3NHDbpv5HLzG3b1gPbLDZ3yOaqRr4c/G4jjkbQwnh8
zUEupfN1WvxScqMirXEEFsOtWezHXwrEehbKfJml0H2giAYi7KS+WxBXa1PjwWDbxG2OfiCUvLaR
FX6CLmtFPhQ+GxpqLjyShycvDvJJWAA/sCyySQRRJLXE5LOURl16cfltbpnd6gHow7D5ObNnnrq6
EQUe5y6Z2d3zrKlSOqghu5sWOXCNYKaGxqCMLuqvG+8vyzkw2t7XThVRJCQCdq660xzZ3mVdmj3E
O9KBPXthR+50OpMu3HHamarJH+GDSLKz2HDC6cnibAWN0gDjb6kXwigA3CVUBx9yTg5UM30GYA4h
mLNuIs9L9KeirpInZzDFEKezNQebCp9zg1v6y/TqkKwu6jU5l07SStwqx0MULxXPnWRI00+wcMYz
QIlS3amowKL2eQgkQ91Fa3luBXKPVWhfXYzev0C7kTpVuDZtkxJ5bApghdF/IqkMmFxGyNJASaXw
WVuwK/0BcOSSkgWZaMMO7vOIKj3sY4Wcu9khy0D8JjLZf9WyEU14p8bvnioDKa5gj9bG7trjQsuA
1ei5IogiFFvgGQMHJWwTcJKEKun7sgdO8nT9Tym4sEft1+Y9B0dI+RSxdzCLHVwwc0/+xtRAMtfM
7shm4/rpuiCKapZ/MYwx+B2SEJrPwz5anl3Rf4OEGhe1bB+noPX3ztNsYAB7pThECXBlF2lv9d2j
wHK1OKL+h2Mg0eS/GsU0CfrSehqr8TmuIu2qWEmhr+FDRC64YZaf1oLR+6cGWh/+1aeb11ChL2Lz
N3gF/2ioca4/QG5N0A9dFoX52AJ973BfLZ/wKKh7Cu70B1/BIY36BamE2/TuqhSA2NzGU5MP54Qt
S6s5AaB6jj7X1gF45PIZoRCsHx2W0Lxys7e4CULH+5kcygFb9fSuanLDHEDEt5U5jwE0mD3DH6JM
0vYodJNfBNv2jy3F36yC7R7ScOPbn9/XdgqOvDoGicDyS4dDKc8wV7WT68tCgrZm7iegqCTmZU5+
F49IHXqcT8Lyn17IYNqRvgxYtA/lYRVTgx2b3zyKJCv+5myBxns0MrHLiayA6qtfUXc15db/QonM
CEw+HJ6Jz3Alfi5ZoruD7/j/2dKw5UoQ1tFi7BX7I1LO247oOAJ+/9udIl5iPhHt+ueyBbA6tl/x
2OlHT/mPE6v0dfEDSqy/BpPAQkG2+sFmIgvmxV3dvkCRGkLAiYRB38rpHbFLLg6krwswD6W3NEzJ
REGJxB3I1vBMa35A0A4FXuDhK7qgXSB3ihC0ExDprkGl/SngOZO0eIQx/WlNs8abV1VvxMAzsIyg
2V4WWtFB3Pf1jtH8+qKBtqwhJS70t43f4bASbcznrHR6P/YzHJpGrnhuPuDHpTAnRizJ0L9zoajQ
Pzohg98Lp4/gQFZhkmtPz17WcH6401g3ar1+FtS5zifRgFDx0FCjNBjYuTNtfOL+0KTYSEqbgj1K
+mDB5aEAI2VHPdMlX8abvvHsz2Ft1DJkOVMLb/94TPkHVIuWk02k1lB5OJEsMdWXrV2cXnhs9jrw
NgzxjbXiW+19iPmGaNa+yuEgW2VDu6XVKHYs7K1XBu+Z7lNSybgtCDmNgiuiLJVD6rkmx775Zn/k
SDsZfNnmqXQ1iae7ZxCxIOn//rESAKUSZ0CeoWkguyfhx66e05tF6BUgdRMpaUEU4VmU6JnY6YoQ
t+LXHD+QlAy0393c2kmjipvMUjifE2ClFD+Cjlyaq37VIUaU01sfWE1inW/hhJkXX2VKRytjnZY5
glQNQaiMrNlBxo8xzn082VnDN3ipJcy7zxQkI+clLn9zIOs1MPrzg80wieT5pggXnaL8UiwXhGTv
XQMLnzGgNR9sxSTN8VXesbSE+UIxoYOaYZeMo+ufEVfC2lDazUwZhxXzDK5/80if5g8sXUv27zYp
FIzqh0rMGPryII4dZIuSdTYEDLyHxuoRfRzxQI8cw8tknOGZKJhn8Sndp0eoIY/2t55Ds+4n1A+u
qKzMqLXmteCTWnLD/fbfoP5QOa9L7bz0iOa31V0rjeigQb/f67rHnREl6O0e3he0Fd2HTKvKJ66R
bCIIKCRy2/7FO6YoIjRKNHtgTIL+WX4j/zDcPJFszYGzqGHKczbXJJ3QdRqaCLmUSCTSpM9pknRC
1a6izujePd3Suadwm48Q/ppl03WIDUBD4gr/8fxWNIJgheqqBrZC0d310mhurceqYLrVHVRI6U5s
CROM07prQpoqr2p/mL2yEPa+1FpskaQjwmSzoydJ6kCZsrmrrUJx3gHidkYg+LIggLL0QHcvHhwv
C/SxvQ73mjb6eernMsuwB3AYSW3m76gKlH1kxNPwVBnYlXuCK1UMj/TC5ZGN9sJE7RjNSkquy56X
I08AYM0rSveDeYE/gGmk1RIN7GpXeOBGhj3jmelE7MD8Kt0anPeFHa97DhtiwPUtecCenKU+mLcI
IkCgURuyPyFfvtcxcogmWdNCMX1otQwqFoimP0rm7g+hlUvYBWbt5TgOgwaPob5cGZg5CdHbRJgd
hcYqBkoypMo1eMykdAFhpzOtmbjktrh8JBa2vnyKFjJNWOYjoQVg925G/R259xvxvM1hkjeriley
TcJGhcR0+6Ymz6tbanibUcF48PET2gXde6Yb+KcLPM6VfhJ4gaq28lSglVKal2gK8/T8a+i7MAbN
nPkSm15UXYKZ9dj3ArIi6XHFtpkyRCnbl0NRjdRnGiv4NETIve4GpXKPqhmdFos4X2EmXSJ5axSK
VsOBRjyzNr3nvDjKpAeBj4jyOks7TNm79BZoA7Wrbrkyy3JR9RlSASxAM0/DTleaLa2s7a251adn
KR4lmiqkQxxWeJAY+82ZNklYeNDeXOz8dhJf4M6Q41JGKOua3HTRWQ01IKSCxIiRXRY4oOkq8Fxg
2vDpk2DabsIEMr+CnqF37akXY2YAu81tF917g+jQu91wxouKaElSDr2Ifidnfn7yhNqF5wQlDBBj
CGBWysd3aoueiyEiIb/XKZWlFD4k+O61fh8NqUdQ7W2g91COiZ7ZG+Js+eUtuhPva4tu6/TK0nWd
07Wo4NVnuCDyOK35QnGfC0EhvJaJdxdihQRU/aZh89eAnr5AdyJR1rxaKDQEOLv5XEk9c4UCH1I1
GrAmUdMpD1KkIktAPLQ+ixOsluWvHNGqmkwb6kjl4uCIscYEU0bwn+eVSq8ZEX1lrqVIL6dS7dvP
Y+24WxiIc6199C05BtLx6jaLvg3mbEHtXtVc2j3Mhey9e8+oTzQplsEVl5EQWYxcg5oYtkI06iaZ
Wtq+2+JHu5BRnlYKdi8xSv95HX9i8/MPqu2amBdSNrP/tM0iFGQvAU2/XNLokT9OpzLBRbERDDJI
29U11MZyPFHaYR92RgjWgDmJEAyQ5GKtgeAwnc0qiGOSD0ZOVY8Gnop3n6AmQdAWgtkEWfcoicX+
RKDsPOdnexF1bXWp8ClDKE2aKfh+Y5uuYEyxyJJ+UMPgvVQhg0l0I8Xo2yd5eQCJVyE/9UYlITtv
36evUApJg1hnYcSYtLbP6F0TPMAbeq2ZOlAVPyvgPKt1SotTWlGavr5bDcPjx7fgopfg2FgKYUqT
B6MlotbLrZ1oK/8UOlVJVUsBRWg5e7oXe61oKx/yxcRuA8QqgOlxL6HCBeFP18w+9PVz3xknHV9z
k7eM8NwbUiApIJWDD1gHhI4e+mOePfMaOWr3M7Jyy8u5Dp4clk1p6CGDRHY9wRe9B6xJF+gCd9d7
8+SYBi4qtncZX0aiJaP4SfvmZg5G3g/VU8cJKWw8hynHvGqOvLndHsFmp76RFl1bId3jZzU1kimi
GtmvTpG7y/LCqVoDuLhLXY8qq/yhUBHl6zF1j6wvAq6TvGyJxG7rMqTZvmbJoF8o8FoORtUNgHzh
MsNrkrA2J+hw1RdmDjKfbYUXA1EYF55t8ATeAhAmaO+uoker75fsol7qu6QNwBcUFQCaQhxADoj9
IaD+KdRYwn+n2CqgmOj0ZTUooFdB2bTHoP17BT+dRtqVudFxxSckpTkRFBzz8+zTnc6/CWVx+yaN
5njYUW0Mnt92etKNIS3HdfPAic1sztZJupOhd5lV7M2SG6ED32nD7VAPh7/t9QPGTgaDVGjl6UN7
rh5++XSECF/ppuNkXOb3Pa5j67ap+54Ji1xZmXK3lm+5NhjVEAo+cOdpdHL+VekObQ3a/PGVKX/n
b1PpdEAZGZG2z5SyGXJk/DJ+PWeBIsGDxmwTaQaiAM9ELRmbFw8Dq9QiNRBYm/EPTc2RqZjsd40M
PoN/VH0u/GZ5PZUKG6GZdwXAjVFb+s398HYlcCxNLMyDvh8Fnaz4HydvsGHltvHIrcZbw50AZCP4
WRnt/UQ3sb70LfoIYfrCbANMKBjHpyuSX6ntPmFOt5fuL57NiLHzpJweYrcLJblOMJeITRB+GdIw
PeJu7Y1pcHe0BAtl8/RmJzImtGZe9t1VoSuM1bkQDPiDxIgEXndOu90jyw8vo1YLyPXTgUAPoZjY
K9fc1Yy9/Cnvnqkstaqb+6Ep2EibQKm93jxGrZSx0olk3VlX5LQ6FH5Wcz9FqCKBhpslwq5CEmcr
F3hUeunkKppfpZ0HBMFHGXSsKDeNVXbgFxFiJvTepxvpCRwEEW1tNYJl0cZV6/tNcZvfxt7JLiAX
Vyynqo37xnMG5tFH8bHZKRjlm5g/ODDUfcwtIuk7x05aEtuVn4Z3kg3vFG7mW56ty78GHZzBFULr
R8NhxN83sJR40CEh2Slyxxl+y8YT4SI/g83DSvV+EQNJttfch2HDVEFuxKIqEj4X97arrVpjHGlK
DQb298yETT0L/BhKplZ6ug==
`protect end_protected
