`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5120)
`protect data_block
hTX64IeLyHzfa3tJyS5Dfu7W58OMH7owjA+xaI0LFp3qRK/Q/EN6ZnChCLudt63EHLlHyyjW7rtW
Slwjj3C7GbX4TV9Gpkyc04kq0hZL4Hb11/AvhZvJDGCURojEPovACFq8rIijg1OVHG1oCn9yCzAN
npntWoO+A0uOHcMB8KMOPj+KGuFVM9GSSTi4mNfRkSvlNbmKZNbplzshVUYVy5o3/7UofhqiBHp8
huSqQxte8qfRuIoIujVxc/7DrsuNSGF88itClD5hO7vBZIqlsF3ThpQFXCQBEik6sdEqXjYCX1Vh
ibz1Ua/n1C2gErEM6i4aTieusKa4C1i2ajvMcATFfv44bhylHSOHfLnrq5joug5GZmAlAdqRgYXX
Sl1C0ExrJdA1cqm2mi2C3oovWG9wW4rLZa2I2bkragxroKKM3Kng7GQZF2tZbBXzLF4aSX4O+Vg7
gAJZrdVmbMTtyRGyEN2CatfBM7UjBb3lXHZ6DiokFZYOD/+/u6kCE7QpiQ57ECHqMZ0dfUFqsiSP
KUVpxmSPecSl7vLZrMlN0oR1Wl0OtU+TFD95Evnu1aQGGjVOl/tSAdt0Eoqu/mj6BU8OT5OLuFq9
COg8oeu0C+sG4App9QBY8EhnNnd8DSHUKFnoxOaFpKX9vdjH6HVQH71rWhiKqpkdc9yVO1pf51eJ
gbtY5yMbh7IJNOvrViwSFzRc8KWwxh2hKHrzH7R9yUHVxTthc3UvZqn2cHc1OyLee5nYryZZkGpH
C4LK3oAcoh4tDjXTY86Rla1IxB0AMX4XZaeywoPCkswPRFM46/AbEAyR4xZNbicDp1Zd2TFHFGv/
BKwehTQEMw/K3/EtEIUMtqvDeBcXuHl0VhsKj7YkvhNUpoou9Fes9w0ETa8zsCWajMmVV14J+JFh
qTNe4w41KQAelfmVLLiP8mIOycxfkXmCPEXqh/yvoLbQY++IxSfL7wScHmb1VPGVbFgiLoIat/sE
qLqlf19cU2QoUUQIQIrexSVKR3l23g1sW7MEzcxZ/24mQAXPaD9NSQZ4tYn2wSC2j9v7xC8pWsOP
9rM++1yawSdm1K08empr3tpVchdv2LzeQ805G/RHdvVX2x0wcUhzjMfBoU2P+nT7DL7qWidaPZKg
iej9umvaOZNbQJ+oADBe9sSFq8d8/MT+MtwSsd2yWE5tKpLlyukH23jnhTqnHRJLV1RNLXxwFg/N
tcQPRMKvU2zc/1iBt3LBtLNk25AtkwRS/kCkExX74CuB8dcKS5O5T3cy6+DvbE8Jucjlcjozb1oJ
m2XQyxD1onI71IJoGmretvnpc+Z0aUnzBQbF3pjbNbEBhHsbLAALU5nYhe6Z0KVJwzkRRUK8EIjd
CGaZzrTTawxjm7vtegrTiyj1seGVRULVzH4wlUp2tZ3Xw83y+DpottrE+AwAuUNeRw1oMkzmMPc/
iZzHq196yh0+/+ghZ+ON0XehhggPlh94MIq0u4h2Kk0+N1KuxolnIkmUjuzuNpRkqcjeF4DFDocv
ErHFFqaxWyuilBYLdx2weT2QTVFfiTNLNmYRU4lufcuYvv4fF3BoW3BqssythPwb/hmIbVUygsB4
b9Y5d1x/dUJZiQ07fAKcTmf0rT0bxbrtrjKFc0CtAthAZobyUwKp7KVB5U7ZzjO061jZtlB5oj3M
quVAZGM+jsWr/rzAShg0fvriwWN8eNcLZMrufG2O99hxhAuz7OgDVo9gMdctmP38sx61urTlkQqn
WjQpHb3nqJ4ktqH24moSomtpPCHzdX1vRuo8JLfGefhQRdvQdJsFAOAoumSepQKPfH6YTCxeERaC
51HfcQ7Aku4Lun5dp9SVfj+GSr74dHrxkFgqZXa+JChoPEzEivamKtfpbjaZu8Usv9Nn7cIh6rTP
jHfXrC+fuc5SVlA3BT8QgKPHPbMfx8UIqoJ20Wfv9qbY3QNv1EkRUsmHcLqkaqpa0FnQP/o73B4h
K3uz2A7yqw2Zb8IVSBh5I3XMtpHIycriE8B07WT9Pw3CWAVnXzL2W5l8V/ijNlQxKlR7/EPQuMmP
ZzIvpKAHPobhyM6c1oakU0526JGPI7ZMa1WQRdk83OzGxblLzdRW7Of8rTW7vPc13yzD4RwewiSu
PLLmKtkm+Xyob3urTootVIawQ+uuxdjSbHMDmRsNB1t2XbNEwvN87NMBf0zNgw45oSGRZ9jg6J9J
qV9KlQQ1SXU3o9InaThLbaVOruNvb6iwamM1gzpmaR+Jyl2NUw7i86Ia8/HoaKbq9+EONmfyHDD1
/kXnmbV12bdAzWnRWTrJtoaSOz0RUwZM5zf1LkcXVtnzVl/xWNz6BQdBJstA2SpCLUZiFhphxv+t
o61L/Eg5gTlBVh9LRmFFXs3FXryAht3jDGOLymGDy15WFM5bmZPylVJyvdSP/g65jqoCc7JC4W4M
OZqen9o2JWy5alUW4SbiKRJEUDCMMjg8DVdn/mVqML+eD3Gsg4fiJSy1Kp842xdwF1SSGmhYjrrm
iJpbUk31HAIw4RhHbFnhN9zFiz4GtvhxXhjBHFcjZg7fAvx3kuuKPPjjmze3NqxbZj/p4q17CB9B
RHdyK16YzPT856Wm2NN8YKS7alBz2kIxsHTtJr9m6mwKEuxzcjDL8QGiKsaKkA9EtdIDwT71fkHR
+ydhzbJAHXbq0zixfzLhJ65LOgGoqMsj1vEGb8b9rC15I3bzzPc30+auFcP+KprJ2yjkkWbc477O
I+6OUVqdxim32iITVftJRzZHUR3kLbS1g8iszpPs0n6GKuil2AgCVyqGyHl2MUprBJHLNib/IRMw
l1Hd5+InXawchk+l41ZJOxG4h27b3Vzj2DWVM94gfACzRlGcCtPdtZVSa4ZvSMAmRBGwdysBgWo9
IDOQXH3/59vW4DuOxZKsxhXM55RgI3gquRyuUFrc6qDuzP+3XOaiGfE25YgPVLTLipuYREeg/ls/
8ImIUcmMW/kVlgyJO/m/GTWMDhxzroVkbXoeeDWzjvplbGHqyYFoHR+wfXCxqjRkrPH6sXS8ZB7W
FN9gsncB6s6XV2cPVMX0pCHKAezH1A/LMoY6YDHyJEbPy9a9TaRiffLq4hDdMbrhESOGpdtmmJne
PuV2AHxKo5bl8kWOjH68Lg3vsqPa9WTi/IWASRu8PHL1ZTObloDkOf4QJI0WQ6Kan982kRn5ww0X
uBZ0/XMkIvxM+Ucjk3J4FEc1JmRGBUqZvZmcsnyg376ljvXqeFr1ZyEPbQnfxfthvkRujmu0iRdh
/GybvRLR8BCAY+f5Dml9yQbKJJlYx5KbjmM6YE1r/UV9Uh8GEnHIqMxduiIa6VJ+3ysBi9vbP8Y0
j2Imwb43++qzfzIylodJndoNCgObC06UTm45vFvZlhX/O98obE2c2pCBi4AHTGkE/0yWshYMYHgp
XbKw3gYmMYYIAjJ+fjODXVeQtjBpSsMflHmu3NAQUGsOb1s0/+6nccctSpbet9KGDe8j/JFzkgqi
80sJqabWJryCfq6PoMJrEoYQgH5KKd/Q9/y8zfO8TlxV139X+UzQP58qJjYGbhVGPyQcGBk1eD+d
IO/b314XCVzgRJgOeQQYGrfZfj5kDE6W0AaR5C31fRbVE/M5/5seJkmnvQL5p8rQ8uIEe4dY1aRg
hyUKoEMcOP6uDKtpEx/maXMbMvm8BASn4s/BAs94djQBQNhQno3/0UuxfHlZNX671qMPXnNyke3T
R7u1a1/KKPYDWNXKzJ7+PbFKyn8VNgmJUK7WhmDKi3+aRN+1wgIA/kCJGhx9kR7gcE0+M42ykdFt
S4+lFe6s6+f68Z3Ol8bycy4SkLnuQm+zILQiF4Nxmnpz1Dci4/1yzy1znyI3uWAB0jyDQMFF0PaH
onxGOM1apZvaCPY6UBgVV8FjoQ5WovHHSiUCnVf4rxJFhf1t/VZmFIVyj61vbw16clfAeVcKBD1E
BcMyrQsQqHf2ivGOj/2EMGdktwgww9z4r+UOJKranBrArXcbvqIlNX694skKIbmTfgMQBZpgzrnM
rJbe4KtAcSSsqdT3DZXy+2ee0UFOUECAFaleuqiZnOiCJ9RSDWvNgqIy0ib28lutH+b51CoN/WEn
zBm9uonkBVsEltTUgH1ucbcSA5mIdxexYcu7ARVdY3jc6AuouoFY4krPE7Zei1qVf+uWuZlqNTcR
4kpaXyu/rAciWuH95oKiilsuQxyRSFYTMdx1qjvcPudDE5x5ReXY/fLPUy4bUCadfGtZnBaJtI2Q
uwbQrRaiCM+AdNPQxFm7rrFY5/LHtWmtS1ZR0ksGH2ngMO2anXKLfRFrUBynZxmJime51X0KvFVR
NzvZ5h8FXTHG5ABL9H9WOWaktVN6vCHzuGnaXxvc1YRF932MF/bbfOHp8VxMwHDV/Ix9LT1e962s
YZhPvW9x9IRY5xjpbyzVy1IZ6OT7NNxEcC+X7XII3SK8aDKeSl5C44dmQM0/tsjh18/9ud0cR8ZP
IkBpD4ITXNxCKqqbSS2DT1iC1JCUAovXFs/y9vtvIPS8eO4b6/u839sJWApd2p49pU6zRKgYNzxo
v96g8ihGdkqUAUc2qKD4L4RU3hN6YXpBpmrCKokwMP3qWvntGyPUlUcy8QnAzjjsN+N3oDoniRdi
a0TypL6s6wpKoWHBlwS/M2X3wpN/iI2i//j9dF436jqjO7sQfyDNXgeczaKgOEHGGLjkakcApF1H
I43E5GK5eqLsf3IYnufkNiNX26xXcXKipwQtD74XC94TbXq4PD9b/NFJSCsBTsd0fvp4NPPlEZ/l
IcdLKs9YWWsocXSIP5bV/9jp0nwUHaFxbHraRZF5k6Png5E1VbSg2QZCro12EFBWc9UJYJiHN4Tt
PyxSpTdn5kCHvHYzJQ/QrygPDSwGbBp/819d/h7XbfG6RP+Sh8ttl5BkAbjYcAK20BHDr5qHwtdN
meXySMxtRIpTHDR0fjgQRsOEuer5GOnojRYshCIB/DqP9A0VpYPqFOTOE9QZt4GK2AIt8x5vngv2
DRzW4od32hGCQ7+Ng5H4ABVdWV9aMfRP8nA0XEAm5qMzMpQIuJiiHhbVHUFCk7137uXpJMrcUPY3
ofjmEYgQeJZ4lMlUidNuTZL9Y+cgpCEF+DWXrjl9DF82jhXtwB52GWch8Vrez1eM0rSFyimfLn88
JL0JvXakRwtXwblwlQmZdPNk5dTX0Vsg0agucVDyO2R7W5mi9x8db3jmzn52JtP7rgDuemSbEUkh
2R6WH+HRfnj3Nzu1++KDzd2TLWRBLWwTen4MBAWOKuXlwrIO3Ao019TIrGI47V7pEBPK2Stnzhks
KAJNqJqYjdkrqkahGb55wW4mdDkwB6yxebEoSoBpI6fmT5moLJaw/G1hgELLnpVSZFXaXX87Au4W
YXpvSb6VSKZh9WwjgkF9jguPYXNPIKWOGXBxnKathQRVtM/d7tV34KpLnaZNNdkplJpU5MJkIBnn
pgWpzD4C50fLgcqW5aIV1lemxLSHGz03acdFnFO0YQufXGwIBXD6VyEAA9B2kiJegPwgsB/aWoY/
zuqTa3l84LT+Be+Ui/FNge528NsgU664Idy8X81XlXzaarddAY5UC+mxEef7o8rCCGMVBAvvMi76
8aT8DGOe5VB6sYzF2FxYh9/9jUKvSjVLv5SoRKps0eqBhx8fhVsYzlNiTrARtE7eV0CGGklfCHdC
mKceLjMOy0W5YdHWossaDlulfjr+yAIM140T8cG1VSnoJP7cV8HnlkglSFKDFf/Dw3TRmr5/15cA
8UtGMw5fV471502SsztCoQIGdpKay7N+JXaMbOrK8ZlQ6L+g6USTY4kRO8q2CeWl1GZPd0C1vLqn
CNLntlsxR3TL++Jjfnsypkbhauau6ppK5wY4oBM8n4fMfetbi14KMYrHirEZsJW64MzoofkclZLl
ikfJ/iK4t7WnBK4C3M8WUP14myCTp/nRjjoUAODDRVYP+4+gyvtWDqvcxnILNqZML65x1eKs4DHE
aLJDsyW8n27chBhnDlhbFQyKv+480K9Pa9X4VYbMFwLDtHAe1iCESvgrYVAH5mMRfTlnjHzOkYZW
bWBQzRIPhE8wy+Gj7QOJPSIdfGGZrQ01uh4AN+iZeG/PA6fPSk+P0qIpRDCawvHLulL8i/RM2a6p
pWcvmKQafMaq1nCDe5waA7cKUWlxdkb+Ytdgi3Dt0y9l3zh8eszK4j8QdAAe8dqVg8gd5O6G27jr
dqdj3rLvQXX0vriQcx9I7ZQDOKU42I8MzrH4qQAlYg1SvuW2G6yDwk3jr4J71Ii98fVu6NE547zf
r6XfGWSsZCJmcD7aX9NvxPxiiMc/Q/T4RzRUvvatrQC4XTFLGYGYJYpC3GBikNFtiFvQsOA+7HzS
qMa0njrUnwrE3in/ys9Dc9TTH+Ke3Cu04rlAWswjCAhAJuWK9VP1UIzHqsyxyAUKc+AKBCl1dQvu
VeHc6fMWfTMKipZUCk8kwSn41HHfIRlh1wOYtizGqi2ghprRd7gY9Yan/XOAxJzwTu7/fHLGLul6
RXZffVd6LwhzKYMa5VdzaJ5Qor30OTnYH9NGEgF71AWjUZj2en5VQrHYltuqTbWHvA1hsHEY+fls
iRm4qoM8EYu5gseB/y5r5BFumQDShQbYVdqeYN6cxP+7MiIgfslKV2eLDWs3V4LSh7z9/peGAvZZ
hCXPtvJksKUVd5VPjGGo+3LqjK6OxbClAekJFr/Xvbg4/fZjXnoXfmCsOO0ILfYiQwzkyjGaXKgm
0N5L6Dcde5gfgf9+2oskwyDdhx0/H1PFYX5wBtqCShybo9f6lxpCT+Tl3v5ecuk=
`protect end_protected
