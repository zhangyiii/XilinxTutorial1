`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11744)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAKBo39yeXSsyTf6n7wiP/+JPUw7WB4txgdDJWmR3+fxLf+XNw+OiU1jw
uyIiHt5MtOyBFrRSPyALUOIKsLO6g/amE/4QZ8BmkIeoBWRDcmzwOxZ5M70xU2HXkPyrpK77HKs2
p1EaQCiL3b2pl64R0sg8gFXMeVtv183eC4AH2R1rNz4psb5929Uin5NDfxc7L05BfOgRt7xtK/b4
brwgIBHTWgtmFgQ6gTmFKk22zl4yqcywnWzmhq57CK+YNuUh3H8kcqiM1JXhBIh7K9Yo/9goq/8C
//mqbpasLBwGzCsw5//P3TEyzMQV4br0n6xFi+oCEiyYfbEIERHkekiUZ951xzVjjI59O2b0J+t9
DD0zm0/xqtRMffLHALvkNMYDX5ws9pmQ9WxU/pMakHTdraqWhipoqtv6rCFVroHuSYMkSPkohyqE
iYw7liaL97+O1P5j4G1LbtBVqZLFEubPUaimvL2Dho1klepQl+p1VW/kCAXO5pVEEFgDq7kmiYm7
ty7Ke31rH4E4BZhKTl43lzjUKiIHoZwzG7Y0uR0piN208WiuBzOppMgAXR2bGRSVdkMaqxnbrPHv
dKOub7d5URF2cix8/zw+KZ+fh+lHAHLZiRROsyOfXtaGUVdaTI+R/OooJy29ljhSWd8JT64eaIVs
qUTJMMfyQE9gXevgS/r0BsA8x7lBU/c1SjtRiIzTiEOqO+pbgHHovrsf2jaaYn1LtXmpES5W0Znn
U03X44vKPMOMsD9rfiPgafdLdEqQhSWHOb63auwTFgcemjHbCOhHLwEETC817OKCsZXmOFy6fri1
FLLzkCnoslbgFK/ZInfp3n0jCqKsDc5k0ctzpecx4T8CaGLAO94jfliYZvNgci605cvb2bsLChTV
k5GhGDHlfCjNpYan2QDZ/V9t7xZPNTUXlYpvoTPSfLxLVXKdO4CyVjypGKMuhEq960dvqfJHglAk
44IvzTq6TCk16wmN6DG7tZRiAu3o1aUDA1O3UUQ/hpwNW5ldUZluCc0xxXfXoowO0WvYiMn7Ykjk
LzGOwSZK5qgtTxQRX2T+ea32+qfuEbtlCInxJVNyrUcj/d9mcLekx4j4WOrZvmez5+Ch7Vw33Zue
TBka3ukOz/mt2IV8DBCpfR/VjDx1rOGYN8gPuHNGfFeP+NtnS2Q+S8Fc6NpF2YPfzCRriw8MxLtD
MJR1Lk5l/6yRZiFeIt+4W98ALtjWgF83eqO5UGFVKidgGjMq47r/cs/9/F2QnE8TnDWCXZ0pIY56
MTlPi+d8CQv/jS0SajbEVJXvS7zZl/VoHzZl3YNX9GXRluDGS4nqZwMCgQl9HTAi61v/ooKM5z1r
YzUp3BalpBABI3z89MNoihg8GMrWADxqVVjHrUWsu4hRNnRCDImHzQVP8VUwLSop4szu/WvSjWNV
3JHABr+l/CL7kkR5MdUoMPHN8jAoJEe9aRbuifj/b85+l/A4BIo97BntjFfk+o3lJC1lisivXwLs
16z3PYnkauwRoSP0geTOoRfquJdj55A0x6/phiEm/FLSKwOufHsRIpVRWVh2Hfic5KLSzcXh8YMP
wdZvP+IV86YT+jm2h8XsWqk5ETaz2XyEqCAjAcqH74ZXaCldfCrazaTU+dUjVa696/4J8SU49PGB
5EpvKPd0Br1mT6FmD/xMeWQl//FfJiVakQSot1jqO20n3ibpxr2/trI+kBn3O2GbXi9EyHxrEcpg
Yac34dOkdGF/IL/6jXPVJ8/SipnFIiQq1FI74SqbTb9dd5m5LB/iZUltupOlN9IZGA8XP96/NVJd
zIRsDUPjGE5PtP+W3y0h5aw3/ym1w47t4lb985pBDzO5yT/Dsm7J8nGleBBsm1c5I7D/EAAAU1kz
8rDWCrhRj8Q/a78XkhvQH2FcS95weHmUfDyGrC3scGpnAUeYUP9oOwIFuAJyJeFZi9/ULRsP4zfs
GgsT8z/99V0I/YU2prmRdyDvXhVXHvIt1PBV53Ihbx0Lm3HMvjOh8qQ+g/ktZbPHflf00Zhs0fbB
XRa2PmMlOK0JX/TP+jU94nNt4geha0VJZbW3FWhG5WqWegbLTafpWhrmblPGaTAVn00pvPqY+hfq
UNo1ZynQN2rSJN4/jh3LpnAiqR2ZcNX4K+KEoRagjDOGbIfcUynesuMPidQ2yseW/ldvFg08ygxF
10gtliemih4zUWnmcHNBnUedfDpeezrYYnX+t8PkkcYyQpy9x3s1oqBv1l2gyoEQG8jqWQckHz0O
VqDG5dsOa2F/VHt1KXrkhFbrIntt17Cz+G07VDHpcbKbl/7Qu/v0WlWAa4sU9+9aT8o/HeqS3Ja/
zlagU0L/aEB/b2mcAhD8mxoOrgjqq0idGL/VMxdFfSt9YPhazrlCkkhS4g1AfNbVb9sukTmbvpQN
kVMSd2w26dVuuSJpr1YAnRdfHgeOkK4Zf8Uls1RhjiAsqkvPrdbPCFcb7mmnNRBPH0T7waTZUCP6
8MRiVby3yS0T++tHFbLVVhAu+bK0KfgrvLZ+3ha/PDZ6WAUB+OHFJmqExvegN0wbfB2Lj0zweOKI
ENtFckPXATzUGDbC4XtyHuCOPMfPNeCekoVzSuDTO4xKljXEJij8/URJILUMUdkHiYn064F5fVdo
xI2C81rFbc5fEmjrHT/gdkqn85qWe7DKNjzu+YV3pSfkF92by3iTE/kHiFqA4NqxFYnmd6jvwTNJ
c2NRXfrYOdWVOwaMsDG57XolaijGs0oo9E94IBICsH1SG6db28z+BSesNor5T9dz+CaMtJ3RxVds
NP0ALYrUtSBc+3S7Fx0lMjMZCsKYHfZ444AhdvXHkXIPCBpd1oZ46C2hI0114HVzRYThwXf+5mZp
rzCh1MeoT9Eqaf5fG9rDva+NcidjSnObb1M0xrFbnMkZIuk2YE3A9HhKmDBmxl0gqX+NbZNMj8b8
rdFgGxWcgJOORIyWytyXt1QLbPj5FTwsF8Cjl2uhTotoSpD0Y7synwvs8zTebitkdW8hnTyNNOEZ
tjWeedYRyxJNfQ1k54lWICYDpRSlQIsMdq6e3pKjYlegHPeRaBsyGSFE4FaX7v8Fbx1bCCFJE/rg
wd0LFWx5YTweNTuM59bpavuVd2a68oiQkZe/NfkaL+PJ3A5+KG7IpZL4OZpfj2h4n2MvoMVuxyo9
/h6gyak4+q1+6bCaUkWS/HiHwde6jYc24rq2DHRmg+I3YRo3RG4uXuWnkuZrF8Zb3m3jTKAx6cOC
3ByQkN31t81yX0nCvahB6jX3mEGd8d0XDJ5fvnI8Xzygtiy8p6lzHXRh4O9mKFjTkvPFWY3cwxy+
kn08iI5u6Dq8AUtidbrA5BqOLb8oH6PwwzSkF6UFLk2VlnYx1GxE1AEz2oHUgvdJxO4/0KDD2SHk
jPNgPFb6lKNs/oQ36QbYh3BPwkyr1BElzAvTMY9FALRMvimrRFKECYdPH/N00TWYklsab8MGPts7
L6BpaIYTOPFQEbBV1RCY0r43XZeib61fEaBgE9rQRLhztwptmH6SXcJGlSuaXnTzxQqRio83rjhc
fbUqztFewZWkYgnr851DLlNsi/3UkBjFNEF3tLanQq5GAtQCZTq6vLyQWUlZ8GcSI3pyk1hys7AH
TRZIh7IWFdz9lSJdDFzy1dVWEeDqDChvqKF+HqbbraeMWmjUUPX9BSMi8M6gM9H//3OCEaQgeioc
Nz/tReHItDytHCYgFn49UEvxLPkZJWknNuF/NVdvBnY0LxEFeSTT/Etf+Xqv778mv1uQQ4OpdWs0
rBXKsjThWvx6HtSIJsrmdKyb4UBPdT9b08iopT9onmmow7xJ4IVeXe+rT2VBsXWTcvVYg/1Ge62H
fX+IuBkCW6rf1bSQlseGL7pYWiDCXuNqg46Ug7Jq6St0OehkakIVR0cP9g+xk7o2F+UFeklYGpVN
VcYO9WkyL5wtrNiW90sQfK18hD6wNuajuPAGQj3E+s6+SrAI5CUrmGK9it3Dm197ypjb0ieSXuV9
z17RLu/yWspFDz8dnFI0h7n2QlVGF+FMl28j8Qq84mVzFgpzGXbVizUudZzJpyNNMALUxuqk9gru
QExA5R53bzn991ADC5OGW/lpRuj/JTm1tB5zYAekWfePabaiCgS/HCq4lCScr+x2O9ybbkRRAfLX
6cdQJOGglwfu+jrdJAW9c7v/S1ykYppv1Hm7thotYnKmrdy2FnGrCxQLljKNoHQI1/TCu/Hbz9fM
DonOsN4skwmfdN4Dl0jjc1RuoCCtJNa7+iStDLa1s7GcJ3fDPQKB0KWx5dDJHKQJEUOsrB1ZkMeJ
x7JE2O+ugjYrLQOuVkqb2azP2tKfI3vtTR+G0pYzuaZdkKYyiABkKqGbo0EmNnYB6MmZA/WCg/54
8KZdXj/3GEMO6VAW75Z6qEypK8O4UJWiPIIPwYPCo5wwXUGmqH14QWop29N/ENqh0sixAR/I68mz
3eckIFWegLW+l9WswqW9oV9F14d6SJHW66tKC28UGdZ/4tUacTSEZvLmop+DlDeeFZbuikmmCCCc
g9UXdP//zbmljyPmpwg2DtkPWTglBFsGSo4e8pNmfAL7QLKxEqTHYGoVtn07d/NXdrXh8iXlkNlN
+iP62JCQsbMmL66A2novAtWcRI1/UUpjKas2Ph7suZK8cBUd/p0xr2KbNbJAVX4KeVt9XPGm6X/9
ul8PXOZ/Hc5MxE6/2F0z4XqBPAOol7pRimiI8v3j3rf28/ma8lJfF1DLjvzAWjm7p+FlunljwXp3
2mTrTHrcTm/9mExcuU+9I4BJwm0KD3GHsCt72JNari0rR4b1ayvfFTNx7WnCWFs/TZPE0QpOlJ9A
8O0ZFRbrzicb9t70n9XPhtUlhaOE2bDOoguYpuuE/fP0/K2u0ILClvHyyLDwxKajxZ6SQhPB/H2k
3KMxnQeAZS05kcm0W4CezDHV5KbQjkxcQxMFkjmp5JdjXwK2jiAol+JnrpXn8kkDxNmstivEu7co
bu4d8dBrQ6aiIbmZ+8WGMPpvs/mKYZAVaulD4VBY68Of2dmwHEPZ+kuxMzVHnenTBfpwNMneB2aU
5Prw6bTchYHBbmCi8rqBYV74FDIJwz37F4ATRPfYBoMQarXe0Enx3C7Bxw9Yq4YEuxZJ0t58N8An
B3nD3UFRGlXT0qnVtcSM9oOuAvZmyDYxnazVs2vXH2lNI+tdEi0jnsPG0RMcGOSHWk2esNgEsROS
K+kzqag/D/xkkpHhCkUWM9u9oNWtdYmSPzZYZzb/J5eSjkdTqhaOQl69rkoTjbUnOkvIoDS1us2O
rQIzIAD/zK/c7Zr0JpX2+BloYGSWhkE9C8x9VMqdUE+hXcjUaurgIs+VNf5kuGXbz/6HRDkQPQDv
+8oTWZlUfDdjuqhQY+zIQj8+YlqYciKhEuDCirsRZT13Olgg76nubZYx0MrunKz+4m7z++N92EGL
h587tqRegzRAWlcWLyZW2ljAQ7kzvm/QuBUvTIQBxhxDuIvw740J4BZohGStGkYMWyMCVPLEfRIL
m5j15+UIgt7yl9O8DssB1qZBjx/jy5AdvH04i2PJN78rs2v/n4JZPWS691bzI7aUICxxA/v1dKVz
Jc+wXHz+OhluABw1fzbQBfrV19uGr/nQODzLpoLuWIyCK+TES7DSV+Vc9l7iCPO7/KxjfD4KTfVQ
UiFgYvJs3IggPlsz2CuBSvNeTrlPCWPWK808clrWdn01SyLGtuW3DmpTSvFXo90WZeFfeOXrkqkX
fKjV4S20DAQGLmHH7W0hekeclQdWOg+m15EWNbv09PDGiqaHTBxhS7iIUUDc1rHMCzSQEtYw72T5
ZEKcqkP4StpD5NiIfydT8KcJSrF6ajbWteuLEeQtgzlY6bI5+lxg9na2p3ePK+uZIIBs1xA3ZSQN
lyFO39JuFIDFnWg1fecuvywyEIAkLo+gxexvjE+MyMEZAeEQrBXw2+Rm93GvzVTr/qHIFni1WxBZ
lRyHdXDKJHq1K/jZ9Qg3NVbN+wmNeVJSe4phh3TqWtijT6N1wzqLm3XiqcF/b0zi9Tg5MTPN4Rw3
HKFzI1KCa8RIlWmR2lEoXhKNEcO9zpLwLqsNeGQ1uQ0xLdYikKv6KxHV+7Q/DYTPeH+kAYGAdxm2
AMAs0MoqSdh2t//8/e5D4HWf1SMuv2V/iMxUbTou7xIQ1sxgiguBXxWwsDieHHz7wiTbZmJdWh+S
obMizN+BeF6C5xbWL3e16LG9PzYOCUFH6tVxCJtUT9+hzBajAajDHlIoz3kob580XW065K2RuFLs
aLH06EvT+qcJ96X4VxH5w6b+EikXw0pNYJ9vn6uyXvDDpH1WaVQEA0Yj24kMqpxKH1Ieojlai53F
6uGLbTqsWAlQpJdOo0qjOzhXnbA3j9Je3VCiHz3qiuq8g29qQdZ1TuenwRbrQD1KuBblE3anYXsj
8W4xhsbvSbdZwbElq1ew2lxU8RQqvw3iYsuPGEFJBc+hmjsEQMySm2O2Km7fhhY2BoHbyz09TerO
KUyExysIg17oyMTY7XgtDixiJr60EF0HZS+ocZ/TaZ3Q4JRpaWSZKCIu6BtapqdNcperV2gCFfNN
95JAlqMUu44G74E4H0rbuL8Ys8aNNks+MAd6LhJKKAOd1uAoWvtGe0fh+2V37EwkTG81uB+FCla9
+63dlavnhdMu39PBPWpLn+TqRxGe26wm75QI9oc++Z1tdtJXg7SZh19R7QLhiwfL1qsGkOF8pVAR
77EeaOR1hTF+7dP2G4OaVTYo6UOJS+ZtyIHTF/qC0IRC7ZfpKntlBkLD5RUXKJU5NkanjuY9sCvq
gg8p2Kv83lriKx0PIOcJ3QRQNi/Ty+DrHcu4Mf39sXTbGbqDkMYiSfhUD6quKv2nr6bXcM/UCr4K
wACnz2MoGgg+g6i6ZZAzSaQi7y2JWCWFc8LZ1tgCN/QakhqYwDDJmWL0VRHgcECAzDS1djbFbxh/
sidytkU3mIE/2Mtk2WHBKsTNFtw1adAD3ZMYDboknKIhwqeICOpbkFRo9tGNi9n4T7D0eiz51qQN
Ff5pWzs5T8hnZI84fe111Yt95xw4mHinO2lL/kkWsOPnKspu1RBRsx0FfMQFNvALc5yPGphsr9oT
NVFgXeHn/wh3kW/r052DYhWpK9sI7XZVIta1wyJL12zlRx50DKsWvaATtAO2JeCAXv3GuyLSr3St
w87JXGd4qS1a1DsN3jxdvN+WfOJThMm2SMxJSLRRZxmg9HcORAewv9sSShi5rWb66PybyaRi7TE8
osQq3GgJU5ECFEW+nIKlGDDbu40QRdWxC6OeqTTlWIsVseo1NLWzph1xhAP4GwljDROyFHUK/sOz
nIlU0Yuhfaru88PSORBlRfb2CDA9idFjwYuUyF59sDeTh6FVwInXWOb54ml+LDXDgOx6arJuggUX
zHHkE/q2DiKJzgvzXtnoACB34crTi5FfwFKm1OR3dhSzAYFdkKMef5dzX66/DBbYebmWAD+HvTQe
q2ot0Okv1plPX3/Hcj4eo8LBsC17e5IedJETFUvo9oGlNxGYD+2mFw1AQab1wDgLaGPhldZhzQlu
lRVLWneXJWyVYr5Apm3mYbuEC5G6qXyxCEe2gyX+CvEHHBv3r1aE5sC9emnw60XQR5hb1H1UJ0mE
xh51a19rYbKyC8ktmBv9FzWigBO9tOHBaNrsYK0SirYTLLSkdt7gFXdjdSm6FymsvJ30JBLZWwbR
Kph/FGn1ZHmhb3cjQwQB3+QCXGrwePRl1pP/PmxJ24dpUJfdb3ZBT80WRO+PSLe1A5BADvtv9ex2
CnQDqQWN1yFtQ+6ekM4YPGYCDHPyIy3sAeXA2gfaSrxAgAdO+Jw/1nQbj+7wIYZts1Sfjjr21kPM
KTeNm4MEds0fb3tNGDWFwcgyh80sK3+D65HOqTUp+FXgG2F+DHEr+h7haenaxj0EwSXzu9VE76Hx
OEkDYF1ii1GDb4hfFKOEgrf0VzMemXqv5T5g6h0qqBZOnIqmyxM3vnjFKOk5vSnKajZjiFUC36/E
uAOyZZVoLvDh0U9de8NctWvg98mXdBxCYGw3VNUJJpPV894Vv1bJhb/fMYrUtuZwHbG0RrPYQacu
9CXzIXdQPD85KTnM1I0PsuJzt/VIe3p2RcXPwMFZ3YmqKCUgs3cPs3Kl6u1LXXbCUPaPdzb3KvoJ
JwhUQsWhaXYEqjMrgjX1K37T2ACZ7uM0fOZ8C5qYxIfHAPXZIY3ATIxXbz5xEsSfnIP2gIFKKUaT
J1qchkJp5TLUnMBJ3sgd0gKQNnEm02oK50ksvgKBRpFBzDS1776msAnEcRpNXAgnuCbX/gPfPzP7
xX9FAKjmuAO8ylv/jOmTYEsqIvsqlnlA/C4DulEFXJHXsLsKsDFUXvpGxALoz3gW/YH3ALajnQo7
SS2gV0T6NhRJvtuRS8EqAnVm3zxHGVombsEuCXacV4ecp5TMjMH/6DJokQfHElxzmv6m/CierJ/f
HzHCuib0IIu+LHLfHgWe4Yw+oBA1+dJNNtn/TJjHa9F6cjb1HDojifPgQV8cnsQcrCN/HQxGs4yX
IK7+wyuNLk4elmKrDtnr5VdgSapb0IZOusbgYZdn8JfAR6Ur/064ApgurifUDozGA+tgkh7BQNI0
tg7HyxouSp7+8SwOSBldElbA+Et0Xv3U9Pc1lvJDb4VKPpyd49FuTxeH9uDHBlV3cWU41rqa29z4
co7TU2EDVOSya9Egfj1ia9oTO0YB8Buazr5r4utgKT1o3KXpkzBG8YBWhcuxzFW9+BQ7Uy7rqPbb
rgieNqtDfOEj1QSJj2RCnXIZYIJvLIHXrI1HgVnMAbZpmaoyaXuCKVpC76im6kxYgHsv97nFUsO+
vrNFQCYjH77uShUbMXs3yAiHTKLwyr3cRuobFIXE819uqQ7xM6AftsUV+BL6qFBf4OdD8MW9DJp6
Ln4FV0EUIUn8lif+C+ZnUQXE6VXAld3ISvkU+CLB7kOxVFSZBvzLuqZ7Xc2GSNsC1C9yvKllWcQV
Xi8n7GfjTPQ4p1YF1GHY9u15NJAoSEuNeT7Bnb3CL2Xixaahf5TShLAfqWUASsqG/9wKgh+jCCSh
DEErjFi866Qr/EnkWCUchHez9th6D1q43o8zWG9cefADol2ReCdFCAq88rtufZsYIdNNnjDby7Yw
70+InzWOLum+HCatgU44Z5Kgo5JSbfhUDbmWxVTXrRUQCA9h57amxUWqqJ527aa2S9zS2z0rmZhK
qXOBn8lwUIbUbRpjhn9A7DVg7byHM6P+jpEwMsEUgqEOMqZMSfWueHH1bDbSUpB7mgciqwjGJzrZ
BU2Q0K+Msxlm00vhUx9xl3bMAf/TiHN8NUw6vL62e7V4CxpeZ5FHBhuNukwOomHuuZ86R9MmKqD3
bPUazzD+S1PNUPlePaoqufG0lmIoJsCMeniUlFnb+OsfqKcrtUxOPMrsVyGJNxcbjwkRyjwkwaDJ
0K00cbV7lCmT3RTx+Q3J57jfJP1gSs6Y06rE7P/hkF83ATzppqS/8tpnB+K4i6DMiaQnCXx5N5qQ
/5SXYJhJf3pWaeOQb/++iwDnmNHmYwujdZGp4oxE8/duurE1+FGDt+rwQszICnpvPCERWZV+NORX
Nfsvfb6bQkp8bFTCMhGspobLTJNe1AuRVLdTUk90lrLS3NSDX48eZL2wxbriQuBIaR88PVDxctcc
eMiKQhV5Q6im/rLShpu+H8ZY/9cGIIslQ9ma+kQwdrgSMGy7HuVU/PrII0nWhcgYH9pMrKMmekSd
40q4pwm3t5fTwUNpNYLMEMCfBPTy6/yUKC/uDKe4832d2K/xtitiikYmdYrKYNLBr2yAqZWadluT
YnNtB9/mAaaiRoiok+qdWMaIuXjuCyWGeVd0mapjJx6o5pFQCJiHKQdYT9UDTv3MTJ5KPWEkOnYF
EtdGi8+uzW/2wiE1Dj5/b6HXcff3sHqD7bR1rCswZ9Ay75V3CsFxoSgfPfzudZF4l9BLZh18VIAl
jyY0kxR0QJwTDao4NchA2o3srp9ZKeWB53qWl+WEPv7lXb/IwNfwqEKfs4RchITWwoFb9iO5Yn01
RVUDxR2v8zceoW3zl4su0Gi4jx0x7Oin5JDC/GSGRIoMpYDwuOomi2hPYQh02o+DtYU4P/S+3LbI
FexljNXk6tvE/X/GwZ4hUs3zgwxCGlMmcTsO6JOnqjS5Jfg7mZ2Nax3QWDtJ1SGCiq22K5eLYMHf
KwHKc2jEFDEgX0JY/iA01lPG4Y2Bplm+Hs5LpY43WyfEXSbSxykt9cN6ELE8WxsSmPsIMWtDIz7w
GapMfOuCu3JnnBDSiCUCadbOLC0GZpwHpAAhRdB1qm6x+PBRA5ovRatCGpRgPSf4Fg5vTCMLQyCf
rjs7uN6/hAtz69PVTxIMU/dlLb5T0cQNChzbneNIOEyscY4hjS93KGXlgDF6U6R+BSbJDN4MBRmr
ORPF33XIiE6vhNxq/jOPhpJXWv2EDi2WmGvPBBMLG+zia/bUO0zxpp035+Ykvgbk0mM0W3/DyR7v
Wy7jr7zQQWgGYtrxub3bxIQ2ITiXhpxEY4my91wWksCpGg7aSAT40ionU6PM9VVmQMiyKr7pKpYK
BiAgtb07LSbeOOxfYd4Oovz9ebJDCE7Z9j/rXn9f3veqxJ5eQmPsTkd1kWSCZYjBkmeqf5NoXpbq
IuGS2UZL+2LuGkKZz57Q0tD+cYYkHbJ8EA9JuX1aeiYyjVjwTWVEWCTgXYkWDFhW3bms6JWklds5
61vRRUo3oXBihQvkvGGvQE3zhW7pRQwUMkmcGWcr3Jii9Op9URvPII8rV5c8AeJPh4py8ViWxFzq
CQvbdyYUxdqjZGToVzaB4CK/9POye2D3aHB/Cz1RH59lD5ys7sNzVUNhQEGRjaA4nlBGtkhFYrTC
tlfKAiY5tzprph2jYWNyY1D6vNPKvNOERFRXsZb96YpI0iCW2sHeht3FvCZDAmqOsZYyqWlAEmuq
TBX6kKY3TaBbrIOylXNgjkBKXJeWSlPKLWqel5qysZzyqFwVbeG/NnrQxvwU+pQh4WntSFZTj2sz
85v0Rmk5vIZ7l+r6KfgEllqGJF6/b38OOespQ6NDWCmpPOg+vsULp9szvJK4Hvut1Mjh/73FUvDb
7c1zG5vDAOJzX4jedFZfn7bmmQJKXHds3b1c56bjGKZ9ZVOlYA3CKLsZIo4mo2xeUXK/ei5TPVUy
/idCpGl6Rqr1ytnIMGC9NsUCC/W5MnvEreXBIRk8UgY2sljFLctZH0F4kIYcNlE6c35OXkzxEhqZ
fxqI6p3sDQy48HTT/vTr2H/L4h683xBbQ/N6QUdF28wuDP39WChki9LbRQUW7hs65ZXR9ex3ln7C
ZeUl9CgSn5q1MjlZimXmI50BZxcNv1KpIqc5jxaWTwk8LzokIN++Ix+On9zFjiIqXtoeBr7QaiPn
J9/pINZd6GUZUGB5W864w51+nEu+4FZlDgj58NmKhy1TVZfbAGKgbd1y//zkiXDh60Po7FIwNtgi
+Gu/NAp5bFnm+OBOH+vgDhCQxY512lnYrrrXNpm5glRcG/yLmgtChUBg1eLSXSdnXT7OdCoFlIjH
Ka9IvUoyApAdiEi8+COHU3JHLlOH+prDE2GhtNPHqZ8s+nzSdJQ5xODXoZ5HW849eL+UHPy3ENoW
rSUuPQoBkplPvqaEO/23cU6nt1G3Ic1ObqX3fYADwEcv9RlGVNYylzAbRsHFfqJ363YCyxw1SPTM
Jc1R3OV6w1FAs6ZDmD9PLpAzKbr7b5znqAannDy2Y7RK+HFE1SI0hXULLaq/gODCE+/LnuH3GUwe
J5HR8PhavuO+j4qyDeRoSAO7HqmAE+OAzMxMP8seyCcbHbxofaay7L/zd281fgs3Wp1pYxRKkOj2
TBo6IT9U/c2Q3GtC+FITl9FbC3eLnTDVqPycbLdgy2bvb45cFdOU2RMpi2UWFTkLUPpl1PsE+lyg
7EhYkHiot3+0CWFVQdawnH8C/Xubmonr8Mm4KgPPBB3YRJmTljQU7qsbewOz/8n+Cu92mPJW4d0e
+VdlRY+riYrX+NlhPbYQUTV6w3LtyTd5d2YcGuXGIWCUDrEy6it2+YCLyQ65jBAvhFrxIgGcBAb7
SFh8/3TCMmjnvsyALgTBzWTWSWgl28jkXqUVVPA98uLSztwSHRBKlbpa28Q7JbmVfprtagkYdliV
kHPDkuWAWGj8Rq3JYAro83ACGIMLuUFHC+JdmYn+FXu7CUIOSqk04T1+Uo2kT4gdHkEPvHnAGTOs
DNtGFfC/E1DjD5wbFHQOiHGND18ixZFpcAvAMB37p3aQQ8grlCRmmo7zvY4NfKQDzDoc7iP4TT1H
C2t+wvPvsdXfrGwRSGQinPadyGb6lnBHwQ5hBd0m5qirYTwgSFim6O+JqnM8dWRRqWJc8kmNpy6v
2UovP61Ws40CTzI2DcZhoVbfYoCjZKk5NvEmNzswePbS620+gXgOnwQ1tNuOeHOU6gSvWap2dOK/
EWcssQYgDA3xOyD43ugmMG+9Ib4qs5EwfXCqyUw/UiyTludd1xWqDDb5yTzgrOs8JQtu9y5Y8tyX
tEG2h49WokyEXW9XDxj6MxDVWLFzNuOr4xurXgnGx42cxeLBIO1I5SAQgijXON+L6RAa406m1KsL
hqyeEeVDe36aS6o4eNYMj/wT6AlqRE3MAYhnmDcgwXIsomsDDBDf97ZCbOsdorzV+RsqJqIga+cm
eOAU/wsPVPOyiSttOO38Jr1tYHdSQUNNhdLYq5ooiPgK5ejaEpPWoAn0WN3BTY04RdG0HQ9aiMVB
rb1/ErTUY6FJIVwX4Si3/I9Gbv1oJS+YP/b3ATskzizggrb6WiWUHmVf9Sd9VvK4T5tgrydUpogb
7c6+QmWvWjJL3ulHenVybq9zeVe1edM/WHizdYp23ByNQegTc3rRjehY6QuLNrqEDL1JHm4YY1/9
Pw7+6Cb+fiZE5vX/swrI5PYW/745GwWIJ91gGtgjlZx88rQbrOZG2KiEa/5HNf+TdR3hW0dsdEWE
3j5hq3yTlY/WGgfcZYvuewmV0mT9oSWCIreBgB6lIL5phvV5mFznAT8eJH+qz80Lns4MQ7mLFIFb
XUwqSGsz5qNMehCNZsZo2q1KUhLSykyPrGSdBFPHDxVsqBVXjgEjjoY3T6nafO9msOXqsYp8iWcR
wL00SJ6Ds561vwJhXFpFewaB3olcoV2CA75eZ3RI8XbJm9KLcuSjZMLwJjxqY8wBOvsKYixE1wiA
Uy9yncKCOXCCQfeUIOp3oEap15mLMfTpnLYmtDwQp9h12FQjtCUcIT1jldQ6Lwocuoa55BLu0r7w
eeTZ9IC9AuewFZv7Ch8hSXkgxucIsvernaPsEEduKma5ljCB9/WEIExeluMdh8giPPH5e4PU0Z+l
9UyiRYPMcC7kvpy0e7KhEYM7yonqH35LvFz9TgfTrSuh8jj00VJFjBNoz1I2gxMDLvNNVAyAy7Cx
xfX77SQPhkIpE10biGOeLSz4Doude+A1XWvUc8kOaXE449e2kzHDFqLpu9ljwY/LYZCMtOq9Iegr
fqbwCIf/q8qo8Jd971wqfVhRngPLrlwAiC/eEIe6QzRsXcuyUzp7JRamMWVkrs6ChAamwojowXMB
GFXmwsw9yMhL/Yfm76L2dBpekdEeH/wAGJ0vTeM1UlsE5aATS3sPfGgl5kLqRCJnzkbeM4iOVZJU
0QL6D34fNw3w/rWJv7AzcAaGqvhrl2bcf4UbG172stLtbQypmS6o8gugRuUEXnBFAbpzoudGhdz4
+4Q7xHDzjZhLfY3mwgwm4v8SyOkl5aYHqV4WBIBIMoW7O03GCzxTArYIN7OSNZoGwDz8zFfZH3qQ
SNAG9H7opgRUmmWOZL9U83gOxbb/gtr7LgjmJQ+Go0Nm4318Sbhk4eWqI4z4vt90BXcn9KY8X/HC
hz223apoq3K3ltL5e6xYlxwy0o0KuEfUw7ULB/wOG1hDk72RfgyLngoOGvZsbHZmX1+9Bqb/bgpL
3NG86wkB9IMLGoDMYV2WEXj/vCeKH71ViCamMzjdzJMM2tbu1gmjirWQNSIlGsf+Bq14tmZe45Rm
1NvtUxiAruAzcis3OzaCBoLmBuuiIpIBz6093E8J2Veghnnodu2C8KqwwVsn2U+gykLRfpK+blg/
A6TeBxsMk0zzFYw6Uoup9p4R4vvMmFicquOeHI4nTOaukurqUOqnAA/vIfEfp2RMB6tlNL04HQ/7
R2kUNlru1qYJ/TpA+FJUd2MmopA79B9k318Cp8ivYDoJ7jI6TnF158ES9h7oNq40QhRL/DgJ58Xa
DUcZBKumlnUXSzFHvsXfFkzTdOjEEYyoakHO+j2Gb4rt8j92Ab2+KPHgTiQE2b2/V5xHKgNTjpDx
TVODJDEmirP8gICjDINSL87Z9YlVmYi57wFkxkbzMGzDI054X3yiweauGAKAITcr2yXyBOFz7vWW
zi+8vVQkqYG1AWPTQylyllMfOB9XhHRXi+216a58rpVeg5D0+whmQCWn6jyd08XrwT4VCxtxUdSn
zXK7pJPnb32WMduELYXoIlzMwaOOjyAz7lx47xBoKqcntabV0TwSdT9poANxAj5JLVcyc87z+Rtk
jQJd/e5Yv1srv1UW16qrS6eiBc7wRBEzOhqANQnAEikOFPJZcDpYp+6+7Ba0f5J8gLthpayr356k
0BgUSR5ez5/LjlLR+9Py48Sikf53MGs+vRnJwXKqyoE3eRHk3oi2eFJLf8eb4kW1Y0MX20a8x+XG
Df9qK424XX/btxcTPcg2o2ESkUBn/pKjN3So5TU51xYZ+NU5MpYKW6QJa70LC+wimBPlf4sf26G8
UVf6m680zmduT/ExjIlTLXS4quLp+VXH6AKILVPf9ShILmIx+L1sITb2AoBOe5/y82DWFxoA/3MN
mRlWRaU3G/vLmHMuvNJlDP2oZULAnH2qS1XZ3yt1kJWlPNQVaeggtPDc/VxpoJmtHDFi0DJbbxmF
550xX5TUWnBYat7BfK7SpwYYIVyy54aJlrwShoD9znZ/dkU5auR6q99DIZozO1oX+rVpWmVbwLhw
tuFWxJKJ+dE6r65OgoELx88+E5Aqz34mZ/uuKDzVYSliYw/2vmj++8IC+adu4N4RcdMbBvIKynvk
dz6nj6MkVrWdjM8bz1CbEKbOwuSnRj5PAjwWgpNlzjf1pyRbVFzPylyemmWDmDTl/ZD46Y8pLlqd
8lk7g1Md7tCglaPLZJZ60JDJL7erLydDzcgobmL3cp2UxXg4B9IFXX6ZCNPAO7KgZvYDc12RiXrh
q692ZoEMOrMe1Q0zl5pCrZjCf2VwEi0YHxUH77fgqByaMBSHn/BQmRkYbhPCqZpJHOKvAZupPQQQ
cIn4SsDDFMQzqTlEWU0ismwWNL1EfKAt5TmddqpNB4XmcF4a3sJ7JRa6lIfCjK6ctzwdiAOHPleP
7zGY5ivKvk3ptqbqmIYReCVhuh+1tB83RUXswZtD3pp580p5pZmYo1u8jUczLWWDrXqhCeR1+yWp
n5vEfh9zOwMcSBWnnMpH9e7T0WsfweOSmi312hwPH/gs9KByyqztpmI05Qs72ZRAPTg+5/9Lly50
G80=
`protect end_protected
