`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 92768)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMK/PgSU3QY91fBkoay9fSdIXCM
AO2YSxjwjCCa4kjZ6EGpHLsWaRutaBcN9VFBZUxkmYCPhW57uX4Kq35W4hcBtnnmjZ1E+QXh4TbO
qqfiB2PBRFfJhWOmoL452mEAieXBu0W77+B2mIjhJ+nUK6OZp8pgYLgZSHUn7+z3xWU9uhyJDvAh
trX2HYdrWoldQrGr3T3etfPn6g722IKiDaA4z6LkKhrMmn+m5EAk+uV4uxmhaJ7cr+C0zdAELSMu
LmcRTuW/0RmFS+OObRGDkp9qWKGuEhTyTb41MVJywU1fbUQmf/Neb0YhjE3JiQFm/tcjuqu8kJC2
XpSRTyv+8glzeI/Lk4ICUl12lC/aqC8g/HYEu8j/FF45uEaP0aPB3vZK5N5VaTgLhpqosNOH7Kkf
oO4d2MrNW7UimTmh8vf0gq6IWt9wT45aTQ4MqZurYfgi6aij5VsfE5GTUNtywW4XhsQ3stq0lBVC
XQLPdbOeUm+cImUFDG9GZJ+gS9nnmCT7hM0Lkjir8dzEdRoAV45DeuNKTOoFI4C7k0b6KCu1V86w
JkatLUn3XYhXRiFEJ3TBnhmvfFakt0MmEZWSNuNe2pYcNXeRr4UV7+Hu6CR6RBE6uQzR8qi7tju7
XL62uA91VXzm/g7SywvjV+GbHpo3PiNIw1ijU1v6P6sY20peGUkKJLAZodPQIiYW3Ek4cZ6np/49
F7hooHIX7brSWvvhabO7KEmRbnekO6dECrnVWmmKgcuf7wJx27RW+m6oXWC903TJ6ys4TCfQjJnT
BN8w0UAotkvAH58nFt+35BfmIfAQkj5mdDi7hvyQCxZk/Q1oH7L6TR/IgSzO5v4fZS8h+i8ZPVuA
ksgz6fRaNTPVc1MZrn0RB3bNB9ux/zNug99lPBGoPWJa8QV07ACzjtThArcAFDQUGB3RTqolPu8Z
3cMn3fVq/b9ATdwqaAoKYg+ttACxaj0flTaUwlB8fwq4NBALjn//JqgPzFiX13gbQcPuMh98XOkO
PhXK3OTJvTcpuM9a4XPOTOfasprfhvxqZdwJD7fbcC+PeiHAvdzW4MFpcIEIQKgfdT18GN7OJanW
f6YiA3m/2wNHIHPNfeVhC7LI/mwxrlxidJa9fflqcWBrdNT12Ky2gzpNZ0ef+99nTZuy/aazYXG7
mJq0aBpg+tnRpw9mm8+hPIXpIR0vCnT+sCVN7JexPnyzw9Hi0ts/wYz8QpLFsTezQ+czP6vKcwxo
9jgfyLeUtq87k5/+4/vPUZApR2WOmHLDbih+onh9v8wN2ut+5fdpaCJVlLl1JSR2Ax6fdRfnAEHm
NFeZ5CbPXP39EOYjnfw/OZE3jUiHt3/aB8lcv6jnAm5Br4Ekq1dnEvgpJZHJ+QyRte3F6d5yA3I1
jgDLN3TE1Mj2xufefX1I6LmeNKI9avG0fT7Ca0vUVaw0NbYEapd8wAH5IN3t1Z8t+j4iAnov7ySt
tBnBbX61JY3j1YBKDB2vE1KuCVSlM8bLVkwjRIUg29mto2Ej7ZGZEedc3tk4EidBV9uySg6p9JLc
4aEBvInMR5ANBbFLlqIde7+QRJ4PzeyYooVboN80E/FM3JU2gE+6OXQuWMgLvolH/Hue96Qvm8Ji
AbzCbm3+nxryqfGvwFohAc9x3bdAKjdQGMnxVX8rEHH2HD56ii9nB0aPhyDFmSfnQCdXWsTyL8aw
Fv/ZjblSXo/CyhIjwKDcPpeocJEclNZgQYUP50n0+aQ4raUpSYPYUyvjJZN8lSnX1gAz4j+q11pm
zNInuXpDzBdpl5YXz7KKzLVnCqjlnVLzb/Rs4gvoW3ZVVkDqHIOuG2r9dPWEDS7Z7hM2EeEFzie9
qROQZpxSlF7Hj8OvCpQK8vw22Doj/2lSxOc8a6odWLcs0rViAkh2ymHHeejqLvgksINcByeNaAdq
rr+507nRSYX+IvA8LVTLavT7N+bWiVJ677EockEWdgvaQXBJ0F6GrDj6kVTlm6+jAZokms6ItNZg
nw4IUug+/cqRmAWN361+udj2NQTMNToZmEqy8LNKHHEcaiIfEFX0ThCNS1iQ83Mr7aTkKsu4K78V
eyl2VJzy6i+uM6OhSg4MqQePXRhBFNRKV7HYC8oS7bTadoUE8woGvAo+PU6bkNuDwHtoUstVrdCg
/+M7vvV/z1aZyUiKmAKGwnO5stAthv+goF8OUaslShIQxNGJW2FzRFykdRZSqmAgvVbk+0X6odai
MBNInurfuivzzjaXqkBPd9w1Fp82I+vT7H4ASDLKeMal3O0I42kncAL1SZPnRMXFOXHDHkUnDj7W
Imb1QKzPSOBB1k9Wg5J7iYBgwdH2yOCoZUw+B8iJrmL/9ZHLda8zc6qUXWVByd8t8u6a1iKTmvKv
WRMpylqnWGLcjBhAALJIiM0y9je9ji+A1Mha7NDcSSe/vRjc7cjQ7gWzLlz21TViKHmfTPn32kVg
aLWaG8iUJZHjJTIicuy6FmcdhlV3k8idRHNrVLbRz64ylIhfr8mTyoxPmlTwUTC8nBO7zdi46QGy
YMgGMnwIPr2eDp/DGL/v64t+/cDUPgZpd1ktjPNeffFLEQ04UxZ9i9oFTQa3Jy5byY5kf42DxYh8
pwYzRul6+BVjp45i3VGzxOa94UtphvncFqRhKAIPn/qy1SLAj2TWUXEdIV3MCi3582LuZ9bSMaTi
dZofL9FWyiUOXX2vKZszSEdp3RattzhicTNVQmiPf8DupfbsRHo/NfCYSBW4bpdhIpRiKJ0DG6I9
/mTrz9uu+U6umK1YkDMtkkkG23elcA2dZDsK5qosFawFf8+v/Z1p/nIhMUX3vt2LsCGR+bQrUkMr
MvqvwmtMQLqy6em4mySlGZwt6t0BqyBMgV8QI3d1h7A7rWjg5M3jlsDYmmY06FfFu0QfxgL5+4VF
B2U9KIRuxJ6dwXnSSH0Qk+R5lu5Tbp13Pb7Pts6sk3RncxTp3zuJA9lKUp8Rsa/0VzY1GYuJakkR
fZ6vJ4ocqFuMGUzYAvX6Ga8cQnHcgxgvYu7BHjRDABykuEmTsM5FmBejC38o8houoGq2Ed7B+UII
a83TibIYBO3M0xAfo5/ahudgbWrXC6LjI/A8nJ9Ey4ma90JbSqm0o9/iWiot9kGwoxl1Iq91JtAQ
FCOB8kQS1tB0buhJtdIYjyQ8cjXV2i3Hco7bTaSFbc2CqX7jJwATTDIUyv9NCpAb2ijYIzTeHFIk
SUsyt0A9hlnTr//kmP/ht5ajvs6IlkVa4vBe5b6wL15yBrrZpj4p1h3LsVh9ju4TevXQMTWY3nlE
OUPGjdgkkna/iGfkUG+tCGTwsOPp5zbB4RQj6c+2sVK+8DD3BDV6D+nPcGOwq2YQpqVBFWWZKXX1
6AfmST4eXuwLkWU1Hw20yk+4n8n10zS374br+A1n3h4qebLISxStAcZE7eUxGPfswrqNKJjTlsYd
L75V/TJrvOPovCPi4ZKPGuM9dbhTnAUGafIWXYNpE9jVrq92eHLVLkJ7bZrhvmOv8BaLJVMkJDip
Y0sb8msIWexf4xXOvPNwZWIj3XxmA+z70XwHGZomEWnX9yewIc95meuDFWvrN7mmkMOReDV3BT/y
/ooRakCYnoXocCwTkpNMePmT2LQb00345nFDnJNaiWxxW6H5bs6kQVHe8GkwEj0CNXQ1Hm8nJAsK
t1KE5qZzZ9bzJNfd7566mM7ttscpUahzp75L0FDljyIus+B+rUqGRj42Ws5F+SrXZ8FqSpgrxG+M
Y+F9+hE0vdDEWvvjxt+5SV+y6Dm00zoxJVh834AVlE6LbcIa8zglu8fx5EO1z5ZvEP6qEitCMAC7
71XYIbVx/LOpNGQCN2pnHT2DDITxfOdsy8oY+Kk8ucXj2FdK8neLbrD3RhesVNVAJ7rOFDiiAuca
ITFhnMm4oM+0hX/hMgsIHCywnGTrd6oCTHR+0whDJcmod3zBA8heeYs54KSZUHNof+d7RNh56HfA
6HEzaolnLHZ4NO3PvbsoWf/jxY0DpJaxqKC2u0Kx0YALPwS6a+Nd48JYwey3gfC7ToGRh7llLX05
D0yBGJga2CGvg6bzMzQSXB5a+a5hJsQWWIt4kBiPjJjMsKmxZzA7wjjX6uxULV+FkF1/AAXGfmjI
34y/ej24SrBFvAmN5ptcsZbZoG2T2DRu23j7sjxEWok4RRC0C8uz2yWP8J2G4QzodaR3nETdRDjr
D14BhVCRvlB9vY+v9eAgNWZMB25k9EzYYZA72bfdIJQrXbFFlqy71StBOZJrxuuWLneImIrwFA+1
QwH706mu9ouFSD7dbP3SPNUMNbrbAlSmVAA0FHGtPU1ZZL5GLZlXnUklZL4JPRuMe90yyLm7e4a6
8FTwUfkl/6foYbfNGGkmzEEhb2MyrLwM3BN2APpnHJJvilLy6MIkzhE58h9ZVVED3K1JfjE/9bWC
qhDGBpaA2GZCXXO6ZdBdJkvs0MwU95NlLCAY0FW9/u1tV9CqKtddkydJsOYuULp9QsVU8NoX7gvh
wgBFRZ9uL31pda6dxbEsf220AaOtzN0nOrkebc7IrdYZWwnhnn5CDqbYdO1iFuhH21c+c7u5BQ7A
IbMn3ESq1fQxOxbgCvPPGMX6pgtaEBWT6BLpbmgdH/f8fyJFCV0yIwdPVyQHrGkpJIqClFbD8GJ5
+dA5vObChrZXOq4+h/SsRfHIlb2ynhouYWnAPHplY7uAQ0xpZTDpuWpn/nflMEdvtA7Lj+YXs/ip
ATr5Bmuszh/qTVYJwIdTo7prqVFu6QAkSIJ7M+v4yk+qqzPsL0kszmR6Vtb8TSLLpPJIwrl6EHFx
BRDuNfprtakxzV8F6BDHjfd3RuXC5PjZa84aVCiHYbOTkdaCXkOH5yvMyCmJlSXVKpDH7f8GGgwq
YnzmQJl+R/YQZB2wrHyEnlYKkD1oQE67qK4sIhlmIsrQjk1o5oenNIetNxd4jUO0AdkJC1VZqXXQ
jsbmSqfv9SF1hdSrMIifGSBgMqElfBagmOpTy34EQxzOCKzuPEbb4I9WEPkTroQJDEkub8Ns2pZ6
lUORC0uprVDheFfcCEi3Zlw0vkjC0iUT9DmHNe81T1u2U0oEVvJ+JfBsD2AB390ZiiUlKb8bGpXE
DpbjYiGG5LKVtjxNNrz6agmWyQpgqyos6U4HGn5l6+MWjr1UPqZrYGYO4tgfkh8kJuORkeTRL8kA
mEWgzJNw16EsoH3n26ixQQtIMTnYxlYVNG38BmVyaerjWMLlbSjG3754QmNVWItqJdkItEi/9A4k
Alw6dCdX6JLUW3XJr49LPASujoEe/Ugl6k0wW6zPzTL6GJ4QrYwQ4+IWH0v6d0WZ2Jwwrk5czbUQ
WBtqAvsXr/whzShaWi/Ts8HP43NWSyWA4m6n28JPbZ/ii/Xx90L4+miUxC4Cn76ktCCIC2wEWt6Z
WgStUp5HMOYmNFhbdXMZIonxuGG5YQ1UH9ZkGXmzlpicGg8efTtDivhKNuMUederERmRTYtDvReT
fUQXEo5NGzkvjF0OD3+zSIuc6zHfnrTchUpdTp8F7i4f2+A4Ay6FtpH8uwXojzY1nFGkilIntg+f
qtyrj/HothujbFYDgNPrG1VQzFj2tQunskToIl0GyKKxPMo8Lp66LL3uoDgK0OHCwANKmERJxcss
nOKfyUEtOVRkmqe8fjlGSjr238HjhmBbhayWECCraC4JgIev2yqLlaHTYfeImmL0xjPNB00BjumU
GwfDbAUZwqFyZPUu1oIeHhbu1ltKKKhlhDg49IcHIGoFCOonlXABFp2CnWYTgK9exYVb3Lpl19eG
5Tn6p3lxOUSn5ei7FQUMGPst82txIEU65eGHkRvF3OmST6WI+p+gWTrZch3QxIoK28c0vV9wc2sP
3yiaPIrMK4FXT9skSYKWQ88ob7ssE+jAAxaKx+s2veJEr+JsYsh6WyS9N1tnl2QIfcJurfwh565T
x1cSU6LlkeK3fNHlHpEkh5oxVXhnVRudsORy7r/RBmbTy+GVqv4zx4eDlcdAArONS70mBvzw89bB
bremhKITnZ8q0cdCTGiO6sKTHM+wRnj4LrRs5dPGSDliyM3Z++i9uNBLL2HZKRgVKw1YIMmaroIj
j2Qsx/ynnWKKs7ItfmRBdbFcBLYPUi2YEqzCdJtoHOm65a9VfRs4VIjGfk+fi22IQqTUzq4PmLQm
XM9mkVqE6GQk3Ju7PC171obxBBtzf0ODTWwvEqKV5gyf0Y8LZ0Mrah4nNK0vefEvTql/Qd5HxkfM
WnVnF+CUjD4rGKslIqH5gHqBeVXJajrRSnkVX8JBMzoC+C0FQciKbhaUfFJoFhvExI7JFTq03V1y
X0ZtIGb7tvHDIwXj2Ne0AvWTUYEb7X5P+nvTsmujdhyabjE8gqTRxSkJDcYMn99F8Sf7sR1CnCXh
7qVLc/Wy3s253IrJpdY5wD03VKt+PPG3vfjvWbGVULnXx7J06xdem14/TsiW51ZZsW8SVLy5P/SS
yFEqM0Z4QjgwPEQDb1lxdNEJS/73XxY7FMtof40V2PvrCgkqXIhKtRhmeHk6CGyvC9H0q797DjPf
8H3a3OAUZmqx+Q8cVvlYeLuPKH+Wu/Njj5oLulkG+q1Tc00PYokzSBcL3eaAh1DXAjHau8PnZuMI
JV9fjyRnLMDXhaYHQvINl1KiP4qP5rLl6GGybaK/1cGAXd9ICAoOEy7si1ZT/ZgbX0OlrD2Cj3Jq
RQ9x9flCfVG7lIz94q9xlDXAnR6P09Yv9Ss+v8XFQUa9QAgiygTs46BY2E9ra5d0a76+aJA4ZvEV
KeXXgolq+4C5dt6jpY0M/9F3vMYLq32NuVQOugyhStzpQbl5EpjPRPP2l8CDZnUH6ohUGIHmigr5
YDmOgUnUzvfwW2Wk9JCLTkMtUq/hB1wOLEupOLq5ikLgSGXxjKa2bNNnyYAbGBiG1Noy1EaCvTIQ
M01XJncopkJUdjE8jfi8vMQbQdIbN28Du4YTzX7sA1ZFUdKcUsXHdJXlw9YQQ9yROJhA2MPZHZrP
xhBZmnNjxe/t8NjgNYoGbIVlJ28/cev98eqIwIA8C+G2k3l4eMQcvb1P1JZaQ2pM7fUmzTymMXB/
WVyuosSx2auMVX27UZCub0y5Q8h03V08RlPsxk3h1Sa91/QZ0QhIUhSIvph/9jSqWXGgTDTuZDgM
xW13RQXpvTihXlkOaYCRjDJ4rTYf8Edb77OK4RAlbQ0AbAlwJxHksW634SeG4x01jvIl6MVs7lGi
5EDYBNd4C2VxMFMcqCCdOjguwsQ6XSd8jEvo9xNlfKXfM7qVQZp3aPk4308WdBYsULDK53D0j6sv
wOl3+wa9KFmsSfEjnlubYWgxXQu1EhqpEbsif17ldh8ESer878BPcqpCM0jXdNV7TdxC8bhvao/F
rCVrtsuW7G+OHnMYRN823p/n1FACBsWZLkvCn0/+HqIcFnFOIYa6wA1Wi1X/1PGP14QR5+d3emst
cOhnqidgEOvG+JmKjzznuRY8l0FkQ0FDnHDV3kkZsK6kS9O/TxMB/3AQU5KqPAwGRkm+QnCeX43H
u/bVgjaIcoz7EYRiU689T7dNyt4b0AQUBL4hg0p0vpe733u5x3HGWtlxY2JKtnHHE8Gw2CrHvhH1
cVacmO03byUV9zy63TwPPy+M9ittVRuBdHYocs3EWWn+u6saOSiCoUyMZ4jFlIg+z6HR+NBuvO/5
BMAZMwqbh87G9KzLUP96pNeOg/M53jZeGt5Ajg0CUqhuZetjNVkdKyJqFEqT3lNQVnz07FmC1D3e
QQe/7AL492H1/bK+8Hu4qPnK7Q+vVxKZ7rMiKFEZO0dkPmrPcec2hA7JMzJ8yTdADZWb+IXcK2i8
KmHkGksmH0KmgAlV1Xh8iSNvU/mBKX6Hr2bEVw6c4sdy02nzVITQmcyezTr1mUVrgg1b4KUxgN8c
vjeHZNB9Fcs6G4bu72WSDRBqpuFxSZ70hd3+2JYFznTa+l8ccWfDgyVWZEU5by4Nj98i4/OPKNa3
GFzWmjg43mlc5GGUQXL0S+5UFg3zC/Lbo/V/KAP7dBGXGJTFo6qQZPJfB7tO36neFngWUbUFilYK
/aU7hDkN21rIVwPKyxo7K0tZ6Q+4m48zyM2/51Husw8eXbyx/rRjfWWl58ma857CEevitqEd+dES
+fQNC8IEOLpj83KujEYZExc+8XreJc9nxvEGvbzywcCMMBxPwn5/KrB0JA1l6aHHKcAtn8p4tWFy
ESHJNVWVGg37Vks3rOfDu7ZqhCdXFFjqS+vgI8KxBxT+nSe1AovsgtbIab+O1Oob4gxIjFHaEGp2
d2I2KePTSTfKBDjUF8TvDimCyTPEFTPHkfahxCm1tZlbU+0gA4q9M4t7y6xjI1lPtVPYwaYBSQKi
kYjfMCjrcA/NIiOtyGe/4ZLpeJIxkq0OqM8Z+T08iEZkCk984wSHU0Pgk2NK31Tm/4xUHn/na8/Z
pRTgA+WPipeLam7aMQ0rpjE5NS98dvoZuYJ7SU5zKSD06hllikwXtahk9WWi7pi2/uhFuR1v1GRx
f1IM4SIUpsBMJtrmqLanBYfH4aKaZGd/boNdjviI6ck+pStBQ/Yh9j7sx1OVv8zR7mTqjl+sB6Sk
m195mbPMOIgrmS8F5m1x8pK0C1LWeJJ3J8tyVVEJ6nwnebBSGfRXm3vtWQEYw//xJPR1j/YBQOyx
LdLPJFvtAvcnYwrDKcgv4w6humf7INwJMlUVPpTx/UMwmsr6p5nRT0W/nYgon+ru6OtQS29OHqZM
6kTAUMmjEeVAOEkrPTWy4uXzQ7rW1vQfcK1++KvVR5L2DpDg/yAjsfw87LIbFT9aEbxoMmAUki8W
Of8DOmgOHzP7wOphj3QvORalrIQefUs2eIruEZkyVvp6ff/N9aZDQL6OiAvX6e7iTSGTzFSCZ6SQ
Q2yNJdUxX3sUpk/8dLnTGr8qTSQU2h0Gfq8VhjbGGTsxjWFJ3tNhNFBmYD8yXju92hsaV1GzFkH6
jaG31mKVWzv82F7ghvVdOQmZ9k8cZn1C21TFVZ9k5DDaSJephma71yessVMHAXxgeohXH4UQLuld
TP+dzLOeDO4bTVmvUDcxk08RSN1nZ43wCucP8tZgiSItfYDGVez5xuwoGRY6TGhDkPcQCpP7g0mV
wdJO8lDX7PSMYhYME3D7AshXDKPqsm2YMSQaud2eW9z9QDk++rPDQoMpJyfzKZm+bXX4XhICquqO
kGBVzzgEw7LRLaLaVtUsnDxC00VPLBl1HTbdQux7sm1eXsXrCNt1b9J+3zqZu7pq1mpMwnfol99i
yn7SsLL46gZpQIlGX8CtRP0iVUk/56JfIMWahcTS3+m70NXPWPoUtBajyavjoQlEu5/EWg9ZhmN4
jcZFFSDNmXCU1G0pmltZ2ay3F3lOFTZ0W/U+cjUf8bqaXtyD6t7fpIwoMwjP0P08hwJzdhI3AXsz
rjt7Db4mybdQKA2jTAngiQf90tgdzciEKvbSnQ4M1cGWH97PG4xfObjGcQNELiXT1xqwLiScDuLv
gLgMXKhjcreGU8WUqHoV06iQMo+5FVPK6wjaae2Oyw8YRCFeysaM9R5ciH73vPIo++BPNxYnN0C6
wTYUOT5FAS8vUdxL0TdrEn0ehcAEHVVFejv2e/EGZq0AlcwYVljyE1fn/AknZhypYqp2QrGW71BH
73/d1mmHF1hOwgctMAkUK7kbTd0RNnckyfXZITX/keP18Med2AaJMJ1wmAuuV6uOxiTVMYfOMMgs
B2mZdg5R4PK9wTLbBKWFpsPhJOJVdmmCqlGQK8ArjZxZBcEJnStsPf4Lc2x3L/DBN05atPPnwtqp
sXd2PqF25KWyAY+e05yngPLiazSLRwoZ8NbQTUc728zog0ObOciu6f5eDZgGX9JZarI/XPTfAVGr
uz3Oh3Avxan/OIIZIBWuE1DH6ZYC8TB40RQzQbKqmzEYt+3tH022x8ZbsKU2XyRkuuFIbSmbj+uL
IFfusEH1E2e9qBI6ePfMOwD4IPiweg3jP87GXmbDN5FBzAB7jYBZHEzS2EkjJgIbU9MPu1KBdmmI
4/u0tpjkfsPJLFMGevpY82vW2RALeVam7v2jlxP5nLD4M5WBrZuISUpwv8PfIVsaYsBrkofyLhh0
ElTCg5W46FlS/ak2OID1bglaigy60sMlrC1u/lbM8Y2WtsjOsXYMaavJaK00Mu7rpjkjuoZeIPsc
nWvzZkt1sG1fFQkeMdG/9D9qfCwRh77i52L0viUSA9kA4+ZLSneHWwxpHXY/BWdvT+tuAtppK733
6LI1Hxx166eigBiarxRc9rGiVu7sxqrLR6m2lBapty3m82OLPbLr94WGCmCq5+74j/z5EQy9K+CZ
AwYyMJN3QnX0UerlaIdN948hSOU29P6qu4p5sAZ4AZy0AP/3TjC3J1bmfqQ63BWZVWpwRCUNS0m1
oxqUZv+UZMVfN4I9foWFyrxFs+LcBmhM8GQ4X6grbagkPTP7I4pH5zxe3QTAqzTzD0f6GGyiKaRT
RxOAvl+CdVIEzQpeJFyM5uRtwhpY8IGAnR5pWoWvIqcsbj2uuoQkFgGTUrkLQ5+TJjO1FsZDVHTe
LcW3+HnkaObNj9Ny3NgKZ7Hbrpaz0jKovo+jiC9byjcl1tyxzVqRQdhjY7O/ll7kIC1+QU2xddUc
67HOPZJUTbPD4gBUbX9N3N3VBJTE7cYBbMcwFXwfiItPm15tfu+yFyBz0GZoE3cNEsoowfELoAgD
KjZ+Ep8KvVurMVo8L6GiolK36uK/RueWDV2HAcfzrhheHgvNviLcxRMKNz4LiFQssH5swPV+U/MT
JRYBdSc8Z3vvH0QLIKlXvuR2ExR+73rgAWrprcPun/WfjrVqtZN0BuZYwCpvmox7Q6AkVzgX4J+B
A9PktYr2YWuKvyFfyNQ7SKnfcpfIKqZhxKUip9Tfr734L4/fRRRF8I5pO9IhIpYrkFHFKBkaXJQV
auvOxVGEVNYIoE4A7NxidUh1ncCcNpu74MSoNTlUWDgoYLbCViYH0fry00CWSckToeCHuKAqcWCz
qab8oPorg5xIxGoDgKWOBXsDp0lIGYM+darnz8eUk5tpyu52N7Tz4eiY6rBCgSESbcVpGuaVLrQd
XhdaLgXfMjRhKbdntH0PcDYHvPZS2Q4CTAY95psWLDYoUk1ynbSfUvLGfDpIM9ddpz+xi9CzgVAe
PAHNQILQ/AkWM+FxOmvS4FWK8OJQT0ScjWI4XwMzVaw0fVjwRL5Wfa5xA2xVTcTLRB91bPTY/TUu
YmaHuG/dSIcuxY4UtmQ/CBaIl0bilFTP4edWARx80XiLfwOjAFFI8Pu7eqvj23psSGQp2UgyCjf3
uc7NWESReMhEcMeCqzQy1leLWeZhP8kwmIDUGtQ6g9pB85Y5rYDgoUof5jwPQ0Ul8kZReouFjCI0
/ZfN+q5i0ITQEByr2dB52vg6XvF239OGV/zoYe+4Wmff0J3HMSNs3yTigLrbRMwXE+azI7afKvHM
dsg63zgd8KYk7oIqFm3/ffYFMpOmA9C8P3p0fzmdN2nF76Vco0hMpKdcR4aEYyv+PlHRWzmAospG
HvJKmU+C9/IHenARWKvVVuHNYTuGJSwpwWjC4C7dIj1nMz6YI59MRfgaMTKzlVclfySANpBBIcZ0
1bQfSE9AKWpWxWmNMLUbDxPSzcJhMkweZppA8HD3hOmz004b+d6rZnleAvabKjrhR8RxPGhN8tRc
zkEBnGbxd02Uvf+qdmzfh58L09GeZkxh15mjFlXS/TGbcvf0ogtmIzBU4krOQgscmuLjAYqQ3pa2
SIrVy7BNewDIRoML4bgnwtsXsCVKaOHrywSrR3ubb/AQ5ZaclSDvdZM4XI9mDjjcl13R8ygUI94E
CAZlVhYhV0kQh+VY6+44HA8/zXlcuKNtXwfL0f9eNuVAUGtlvmUM3wOVV4HLR3epG+ETSiNWM8am
jXGoXiX6ANgvighXL9LtsTcOZDebdCZ4er7kMc+x8TLniEvOYL8O/6J16UzCoF6pegTGPRkkLyOE
uWaDuS1gmydfq7C0iGrYG20PNTpq+4qUnCQSOlQXZ2dwazojDb0FsgtRu1VlvIhKwy9qLJ7I0pu0
BUs5fOCvbNDEWKXM3nQ8xlWO+OH4ZZYABm2gfnLvodCejBi2YeMGyBzjjoD2BocaWHqp5ruAPicg
PmbU1qoSb6uWVH8LGbGvmGZEhRQtr6ySnkOqPi8pqAOHVQi7jHEmZgoNyJ1AZfgbm37eQCTYe2bW
CyijgUEBzVb+GIPJAYMdBUPfMAoRKkp4zYnPV6t+HObk5Oxjk9jrHlCNBFD7XFbLd+nm+beMQjhO
wBOsReEo8GEpetzh59AP/ztQzxSLcjfpeNZKzvVTgQvKqL0oLSAYVMv4hz9OuC4UnHbpVKV0+AhU
72m1olhMYTbPRXofMIi4ah3JAn030R/7yjC9jfXamGwfN1VrTn0W4AVU6d3aI6QrBWEFmnRT3Bx0
aoP7zUtwp+dUstTR4a7Q8p7OhSr9/hrhpo8/sv6eBA4DYsDuyLgkUtOnR8ltzuP0w2W63f3/y5/7
hFdYU9qC3+5ouECXY7ZFpfvQtBtWG0WOr9jk41w08t2UXtckiH/JXnEkTS+0j0CEBFtGU3dr78uI
Uh6GbEtYSuvEZdIsQwHPcLsw6CS7qh369c6RemtHXIzjibXUyh7r1NsYGPb/im80vUMgH0U3AgPE
D8YYx5WdwWVw+sbszmVYcKBVc9/h3d5Xd+ZhNTpQLN5I0LdCxFQgPIegjJnt8b3FkJJZciLzsFBk
I3QKs3fgrcEQGzWsD/z09e/8EHTkTy/o8cLTXWtbmemR3o0wPcBOSRkJATwbGCCg0q4wZO5SdiIn
ABbDet/syvDdYYgwsl/O9o/eqkfVtmIhm/MaLwOdpQJtpHXxQegO3Ie3GClbMH893SZ5Dp8fjm1p
7htYpnPuHqq+ltxFrAMy7nVntuefd2sxkiP5XjOFtFhNioXUviGTPpz022oLKs6YqFbYlLEmhAdq
XE9GQsbQtW0gP1tMhVDShpLJ35q8rqbW31U/vtl4fg1LBh69rSrJ286iiR9HZaP6CBHq/7tDK/+p
zZkr4aLRmdTut8I/YihEPCXw16irymhrimTdEkqFY3UKM0xQZ80kmUCIeM5Xz/p4B1J6qYU6mS3S
YyHn4hvnxupgo6Tx+iO4hMVmEXTsZLPQ81E4NBovj+hrQTipuiCFwiL9Oru+C19Aay/6HnBWBcG3
jw3ha5tuJRfH5zYZN4mNoVwmdj9P1MGkf+v1jun62EMx03PQnzgRe5Ya0WPuFM9mcCp9GccgU2Y5
7gzxQ2C4E/p41Sbu490PDzdoTiEPSA3GyfB6fWVvvx0p1ZayWHHoqBIem5FUw7yb3FA7sLs/bLWe
T1+kwkNi5wt4uXNZDVCaODOKxin1w7xgEj+kU4mMDjiSRygW3vy+5fp0SSCkN6FyT5wX1AOyrZ9U
MhRFRyKpa7Nq56/IDmwjieJjHKuwTAj/f+ZjlqFEwvrfdYgrZw/CD71kZy8pbCb5H4ksiMr9CWvu
2G7T6uoXouw9sJZoYwBId79tAmIWaB4gTMtdmVxiHnOYa8939DsM1qhQwq0/EAOdC3H/lEJP2Ng8
u+1Ye5R47SEsXKS87Wqi2ja2FpQADvDDEIodEYspI2UZuLnu0fyIPfIXlZ5QQ5ExmVO1/GdTPHRl
9UiSNFaqnZMEjKMmFlHX6Agswy9G+pElGcEkI8ybqW6do2o7ufyUrG25HXr5GaOD8tfy/NeUTltl
EkDtkMF7h7vHuOUdezsgMcKFl/gdwIWWwEGr+pRqqzRmDcbws1lz5zl7XbGyA5tVaJb1CR+02lhu
/uIODvIyQ66sm8546ccYvgmTaBKstf1YF6bXUi6JmDsggACa71orAN6U14zKf83sHYBGUEDOzSIl
5xXrsXpUbYm53xr4M6pMP00sdKW8Vt3JA7vyz/bweIuDCFJM4nR5FQaD7OOiJaQ+j4A7NTBljNvy
BvYpyE15DEzMKxYaGv0FXQf3QSWmy2kxYn22bDoYD+zlKuEl+OSx3aLQWG1Jki8x1XqXhluydKdv
UeXo6mE1KG9HCNTxxhv57PSR8w4t4pp4hAjEygjqv0/mPfZW6HL23So110bskRC2MqvUIp6KbPG5
k9YvSRcKEq4s3v5SCtCoibv8B44+OqAQnqm4ZKz1n9o/58xA869aKZtug75Le/1MgIyN6DOU3aKH
6sI2NCCApxWSDm8YrgHo+i6KXHoj2E0Tj2gbpuzaLc8NYuXUXnHvl3RqCCSCv51nmCRo+KkUKAza
aiNMhMeP06Xqw/v3ElJNJnY3GQ1CCnZs6oDpXQz6sHQGtv0XeOQ0b5FmigQjkqjtQKf4xHEVNxhv
dIsnphFYaWNnRBtByR22UXh1bg4Y5kY6Rt+md52+Nt4j9pngfllHyA4uXzov+PvqqZYONWmkMZJv
+kvpGLA93/sXVnExmtRP6f6MFfWW6JWldDtPqeGGx/RGdEX7CLqCWNXrVjJrE8DK6Y8w8ctsgXwP
k46HPskfB5W96d/WrrKLvVCWuiwXpp4YJPui/vwartTwpVVyrHVd4x5TghznTKxI1BB2rtN4EkwK
M+odO8eFDi/s0d2RWVQWbO1UG1GNoznrn+wwhPoznOjS0NvP74zapxSQHY5Xjfaas8fV2j3mjSMX
9N/xwPP4AwRZpGYHWKkC39q9A/WIPq0pXbq6nlBsxFH5DH2Ea4WyEkRlN8+/TfiZLys/xDlGIp4P
6tM4DSAu7AQncT4lQgBSHa08NLdM/eFpLkHUMkGvBOejN10dNwCRiyRmKzLKOdcXx8eAFPWloShw
VjyM7F3/NzYzLpW0Cai8+luAm2LR2WwossBYrygf+zpw9El2Sb7kPBYVxRAVt2KX9WZ7G9/tVhJ0
RIz3QJG2j5RCoZGwdkwBANJqVWu/LxquJXVsd+k1bLWdOuF+ZIxC9C37opq3NEWCzCoXzItxtUOE
cNF6VxYfz+wTZj0+Q41CbnA3CSL/tpVMlDmp2yF6mYpUmToy+rfAQhUagRup112bNMaJr6Evodkt
wk7BmJlHmEPWBVqdlt5XYcedWpUohqPAiuHuCw6LiauxABKhCwyjHU1k3z+dAjcEd4LIOm8Vb7F7
0voZ66neaKhP86jeNgCnCMcCKbmQjJkGeQnSRbRUdYRMkDIrxkTYvFwwSXMcwsLpaet8gKeyHkIk
UfDEdvTyf5oj61/pzz9goqtXsIabjIpo9cbowEcVCw4u1r/v8bPhP7bRqqiAzpFtvODaIUSyBF2s
b3+PUK58QzPfabd6Nf3i1r8cXITT2WYEgI5ThMjMR7J6sEQtpfQ9ht6mA90lF5lnc3necIQLhaPC
bJwMf0Iq4wt3bEiIzqnKsv2Y2ZaduKIq2CxfRtq6lYeOIpyytt80NWb6oiXBOAZvhE086fNYC3Rl
MXLXyM8DPimv/NRm4g6FuTH56BaWXGNISB9pPlUzcViQjW6j6JDkkaABaqPs+c9mvcWR8soMflwM
odGQZjeFqnN9WlDHhTAj4Ki2prJdR2rObLFTrwlLDtTOT8xY5CtUdCbYDnLH+l6g+Nv7zcYaVsEL
IAoTEpMTja4hU/HoIlTCHIfYRcrwCpZHt//cwQXMq0CRQuTK2VBYAp4GwvBJUemBiTxGEUjzLqWp
q9njVqPqp8blfVb6nN7kMy0u5sVb5ca+dDtDsZyQ0dIPpFL6b9wM7XV9X/vpWhllow/dFQzd0Fus
O3X5Cm4KAdj/GFJFMOKaLXa4kgYyi1tPW6FbuhhK1++hnsHjx8y1yJuieJZCd30VGuro9LB6pZwB
emndftJgnHeoDn7kenw1rKMGpiBjUWB24sAm+pla472CDBOsrVUnMBEAUn/mBQ/UtYi+TPsyc6IA
3EX+XM/mbHLKn2RqyK320SNsCqaxep1jg8hVtjOhXXmt2DwDIpyCCuOWs1R+267OmPu9SEMAsiJZ
upKnvwjbEf2ApgJf6Muizw+iMEPUyVr9sCT/4QRPDN1qtDFTiMH/lVtyCrtnhe7lYr0CY5bKiYtl
xstNrVFy5rwaUOBvjUFgXMwSGkhqTlyberfvL69LaSFYEvE2v6L5FNautf994Df/ZxPkeEXUD/ZG
Kf8M8WIRHqnXoWrZdmS8RGq45/ALPxvmPo/I/IwSXXXQ2sEl6zOROcz5DnamaI3LHkXio7Q3OpcR
4kgetJok/Z7cAo88CFDDi0mrgQizLhHrZMoq7XsAC8K+UkB70YXJbiTRDrei3uI1jWj/JsiK3ZEy
fMfdFpFKplUuuCtw+euo8IzdJ9gIEIkMGoaB3AgWTHlf5zl9/zgEwgGYvu7TYjVo98/t8cPx8aOl
IyeCoD0M3fEf1xPhwkeO1n4SGyKt3yt6/im65cfc16ucamPOSOLIOnfx5ODxbDwtqURhXI78KQV8
/r7Bh6HMOy7IHSk7rwfxRgFYPD4AClMOblx9GqdssY3Os8ouoweMQFBECd+EBkzTOEDr/7psG9Zg
8EYVE7f1Z45t6euOqOrKueZ8nm59IdjjAQh5kTznCcT1zwJvpmTX254QkSX0D8KsEsdFo910OxeL
kSdrGc3Xb5S6Pf33A5ECbH0GFPNTTtlihQYxOfgsZuhVXJS8C5QqoppDdP3kIGlkJgxhjEnhoO5P
uKLtJnQMg3D6RjRZF/CuWnYQeBABeJCc9jnntbhuk1jcQAAw4IfE7zoVwta6KfkM+c6QDX9qwpvN
zoUdSCWrtVJR1hUq5k1zKpQktmxrPtcXyfkSU9qJONmyEmYXfPaitdk64a8Qbq1Ge3CPHy61QLMw
+58v1tN0aDRWGrjk7HgDHpTBNMlm2bSu//SleRL4puPFcsnncBOPNNICxSK/cd0sam96jLx6VcYg
1AslfPHKzH/fBGKF0TubUlcBf9C7uK1alloPZUCekcnHcR5XDKj87//OwdlXHN/RSSquiO2WA1Ep
EO3OpUYn235PbnF1QfdYVm7v4C7wMZA71UoZTdH6DUUMS6a2U5BDA5lTSOyYD4mI5FVGesXMmHnb
QAXRDIgotfz6xsqhtH9wm7AJzHH6uH4o0c11/+icHM24Z8iG4re2JIp2gWYONNOJtNcwfHsYXyiY
ATfsLYiqwuHc8KSL+LY7l4iFLohL/WNA8zzOJNP+/yIojcwxdAG7AKp2x3YtIHMYju1Tyi13Zrtc
9zMItkc36JSp4zZyDBrUQgEF/9I50/FJj1wy+P7oYjWhJfOsj4+s+oH4eghjMYFPidF7pUcqOERn
cgJGVOa6yIjAIqOzariz+cBWdVX2MeetsXuoaAHTIQ5aza5p6PvqsvBT/PUkckKm+A0qbSGnS71Y
sPFD5fMnQkR77fU9iaw1KGtWchx3/Eaf1h56LLElfftdB1vu/ySAQUDomx5pf/YFF66nJT11xg7x
g2frXNu4DbcZZrmvTPz3cu0t2h6Hy4g6je8+1pynVwWJ89h71wstXxmosNpgkEZeSb5P2pqRAKzq
nkzrwz+pKmvr3UThxJlQJVQLePY+1iKTlAs4OEDUM7+7ATYsncwq3189IC/dtSt8l0H0HirN+v02
fYQk7P5Bj8zTUpJdIyOj3gKlncoX7CJiQosT1ByMTQRwSsn9IgfRCmam58fqdKVqZLv8UtkYo1RD
2bzud/WAVsfQW+k7QewpOm8hZ2p0c6ScfRCrW63Te4VhpGNNuUc3ojy4jMXKkJFfqply7DUQWj9X
edhzcyzYJnie3c+uX1saPqyEmzkXXziDXds4mfQtBtwSafPVL77CZ84kiXr7pEDcHfL7cPRGTpCU
WQoa/gvt2TpFgga5KtLwthW4Xj+0XYiESZ04BZf6xe78qZACv71JwTZTIkyjASdajlXxsJG/0SrY
db5dyrR+44VKIxWwzCJ9L2PGvsaKoBf7YxJHWUcnL+ewpMhFprtud/dQon7EcynlF9yo5flmjO3M
QYTzxwt6yJlFOi8NqGN01tK2L2+Z8HiJ+Up2dtwE/ryrNSICoCGM/CR/lc11xix6u7MFWLA2DplP
YBkRePtO6eeNkwVYhZnypoZuMzBjzU+RGFuXBJbNh445TXVT3wk51E0i6fyYFaH3LUSCU8dWUhq+
5EkcTVPJbAWivNTKhnRHBbAksskEZ5bI/sY0tZS8qLF5mEEqPOpD959B/i18XdkCwMM33ENTalBc
r95U+4cJwDeMoIQfIVjBrpZ5doGEUaFNXUAT9EhOicfHYKHrndQJ13EFbFcAKG9JCbnPAmdKprIC
08WU8hcICUl6q2LLis3DLlwqX2+K9J1yiVjKETpr3d6cxqrS1wsSjSRWKPVin0+D5JDT8W03XOz2
3wb+F6CFcovMjJzCPQVrS4+JxkK6V1HrPnp1JdK9jAT3M5jgS9YYI7KSBaM1e9WpRQwz3yUi5uep
/7l8MAyew5iJEumk0DnfxLsB0SUleGMabMkSjdR5skBzAzLrJ3KvobFoB6RqHLWyI1LDs1JnK0Li
YNjHuIbErv8Y/KLEh1SVPpFkESAlPHOtILacpek1nekInY5nd/W1a+Z1lQVRupIoQ1H0Kwp7o01d
PLgC0qKu1TCxxKuHmyeDycGy3dhMYhO90fllY15bWI78FiF/slvqQ9wcFzZsYcZ/2oQAMi7zH3Sr
zCDKaWcHg4bYK9tl4DNxXrqcJVzhnwmYCXHbiMFbcAArxQ0CJnd94vXBXDczEvow6abudIQiqGcY
G2Zh1RLotjbqOT6STuYoBQAPLl0Nl3ADlmuPQ4ec0Fup7mTGGKNsr6xKDR6Jr787OjTb48vXXo0+
t+90X26dUPj1j9gVp16y9SWjq4plR1Qh9BQnwUjeJNTqf5BlR/mq7kqs+43z5iA0+KPiLvYhImxK
mVQXJAxiAqJB05gofz8OUodEhtuwyHQSspZ50oRHbnQSyvZ089aF4LMnLh0hRstLUbaE+N+EMRqs
vQkzy0Z/jmpzIktHBIbz1oPWzUpUfG4s9bWXe4ZoOu5GTxqifPRt2I4V40mcXNTJr9tRVZYtcqkQ
gFNkdJLIn9JQSA0gKo+FTeRgdN0Z9AiF8Ya8ncYGDH15PyGaah9I++uyh/Z16cGq/vVemOitEw/Y
wFAdWgBxPyUwnFObD2L8dxCH4aNICvYfjHluukexKgp47pkyE+fhHX3bYveFuWrIzn8vnMvIL7Ta
vpMKYBNdFAnkzk/FE1vN4vmVVf+GaP2/hrwSjNrhcXjQja88eTD34qQTkE6fR5J6y4hNxvrKpCDc
+q6X/KCksmfq3GyEAFKRlcoYz+KOCfJh8EMJYdo/EWOXwqcgfZ6laSNx2cO+tdBLFZp0hlxM/Rkv
I87PkqhxlsRjeiOEZ2HaJ+yu2A/It7QhGzcjrY5Td6qKHbNLwFYdzsaleasRVWzBYyZXgHdyKuDU
NHbGn2z/ZwmjpcLtUtOasd4aEMIn9KsRqFHzms6JEokqP5PcYXSAiyZlpiSKpDpSzffkuJPlMAfU
G2a3pfhXi6YyVoAn6p6gjGgXKiYjXWE/18zdZccYmyKDhy39a/Ow5t20PCMWR19eWqEVuMNoUzmy
1GNt5rjy57niU+HJYahUxn4HWHjsNxaQbK4oY0ODher2POIKtBLDCScQbv/9AgDlXHVi7cduTBCe
Vk3RKDEXg4kob/S5lYfXUK2jCeF058bt4JQEfjiXHSkkfSpw2H0ZsDTxOA3484JuOHmywe9NicVg
BQHRAHl5V7RZAvnYadkP/2Qu5oF2sh6it2GTSuLRmR0RiLFGD44mATq602vrKudvoUk44hhvQenn
qS0SXQdl+8aKRn/v6tFEmtasDX1j5qXvnQVLcZl4rr8X0ZjJdTQOSVL3aKH1D43rfSEJPlkcmUWz
5W5SNJZKa3rN/RolnJo90BP90OPCMqiMUlDbB8TcJ4sh+QtI5p0FpVGsqNe7VbFzGMVL0/3aWwZo
9jyFBkMPeLpB9iZE57REO6VOn1aI1yVrUIkk8+QlXiHNqyC22teQif01eLCyW6fynDMZjhVyumKL
j90LxCeErlfkaBVlb7knU9XHLJhOIXKr6OjwtNGfBtQL4zxpfgb89BTUayuohWOUmzzCK3pElIhr
Uyws+gnZNXT9f4/SbDwJvw5WGFKgYictLMfv4Y4m4cP1BFQq/gFS6Qq2zUxDIh8fomRXtpd/9gHm
uIYS7fCzbBDMiLjDQBDY8w2UnE8glMx2iGgwgDz4uBXuIjA/ZX1m5TtcI51/1MRvOP8v1amMemLL
Z6kRPe46LwyB5+fcB0YHWEOYcU0KWiMsEWcLsd8VB8jrH/+QR7zWMRlGnt53FAZnBSMkidCPmEnB
HWQ23kGQ200njodfTgDmEJkAQ/87pooodN+8CdsaxKDfnGvsfqtXDifSBHZrQsxgSEg3P2q8wAXM
FMnZJmUnXKd9gNzU0r2JBjtetogrgoQwaPeBK2GFK9tcXKLH7NGO0vus/S+rsmizg71U/G5aFGYn
p6tXLBgeaL6LOkSiDIdRzdw71YLQk6LbCw1iITAUpZzzRXjVHSIzhwGSfskF11fMFfFq/PMhLw6w
WVCw9rSXNGJftxCRxC33GxegAiYLzibTMsCstcipKlJ2ZvQ3f+L2ezJrQoHD+LXY0FV6GdOCwBWf
V5rhU+yfMPGE4eq07/Y2rJzuVNURIRgrK4CjP8mFx84+GUkSTD1aOq3/i+Yy1lsm+Um/dj+jEOo2
DP3kYY8sVQCBPdRgyfdbwvLgAhgFntNJCTBz1AD0rYEWFwMmm9HuDyttjfmp18mN1ia5c4P6G6nE
lQjmezqVNG/S6aKD2XmCA0g5NrJsuZQa2VOxgqZU6qRPAAqdVEQId+SyZ+0rbEXB+vWIyFnm78nw
gA+4plxfV9820DfM95jBOUF7rlirlU+YqkU3DINcs8j4kfA5n+8PXk3+pFXqA2NWw4h0WCgDGUTq
SRhcuGVg2Xuv9OQWJY7NnksUTSSd3BciKYDoxv6+b/Jy7h9q4V1GXrZY1RyU+bUhQxzql7ohviQz
8i75+85SJiu5+Osa1N9fMogh4MyJIq2wY4ZO6iaiIeghAfa85o6C3ny4bDp9kOnBL6GrSpxLfYJX
Fj3zToKT+DgNNGp6IRUQfabowo7ZrNNL4HwRmwFCc8vQDgBUf6/WGomEbQiAIcVR7qMEWDqmGYqH
Wja56MR+NR9WBdiAEot0+UZj5hltMfgjV+Sz+Ye59QXDMIw3rzvMHBski12iuD3l49onSNZlPnYA
d4+oXvEVRIx41ycEP//SRDF94Sm9EY0rfCqJ40JJwc1gWIbk5Y+yDfhiQsIZq2Hw+lvTl/JzvKHs
Sao/0Hs7D8wdNjbQPWgwg0begWYw0x1lRVe7tz27zTGKeh/vrUDas4NxanmbpKaO4TOY3Dv1bbS/
+jr1JoBnb++I1YPnH1YwTdEGRkEFXFxWjqgPNpjpTF67SUt6xj6r7jsVT3kzUt3pa3cBiiRVko0E
tVpI8eV6ejEa62Oh5STtZubNS34e849hd2VIkK0pJzDm9IrzG8s83fBLl3awA0nxEXnbzS1VZM1c
l8C9+HOVZ5Ev5KI2Et3/xvnNz6vQUNG7/SUjVjaG5+7NyeYEZXhmoRm+TTRNhnKtUCEoR8+Rg2dg
yK6CgMCH4yBx1KHe+Cf7F4stdc7xwk0p5zSukzP1QwfaU5af7OFEZJOvHIykdHPqO6uZtYLn2oRr
Ib8PqR76Gon+Q8XFGRKFGVIt2gSOlMStzX2UO+6BdYOsmLAxdnvHSBU1UqkPxiEuISkEGD/6+x+/
2tFQYzIQlo5X8PRyw3i2rSU4RQfiwdy1o+4YbNvcr+Q5ZqKPWLI6Is1YMXiZNs8zoitMBcMV+Dlk
Q2zIqGgFM8Umu77vcFkkmMc+BBfry/etKsY5Q/FLAcQ15egVcRlkWEInt5hk61TolrA+96UIifpH
hPm1TeeO6vhE6pOUsHdtmJPm+AGqBBPSNdp49ZXE3KA1OWSj4Tvrs0JTQxpHzNmlEwNu8E8p9j7z
1P/oxfcsQ3pYDl4B8uKhi0hCQj1VHJ7AZtFHZcQAP6RQwvVhSQPMYN2svrgpopOgc2c38x2KkX/j
XRVqdCAWujigP/3xORhyzIWWP5D5Lbi5iLIo2LNG9A0W2OyjrJM8aDFM9x+nLOLLFjazygCvtnW6
YNSdv9qh2U6aCBAPuhUhIwHoYkvBrukWoqdKcOT06Rhs9B7v1Bh4JT2eD7p/WdO+/FjEr5GT4v8B
s8LPpiHcDqStLa8Qlp1O4REfCP+ni7clq1BYHHyQDkkXy7S9LX9aLATb2c+oMa8bYjZ6BxbbuvbP
NGjwkeUejXeg20OIEVnES7gFsPD/UxDKnVWMwboyDQdFPbE4n1uKeyuTFRKtBZdXZyDuC/EMvlHj
dEb/jsB04a/Enck9SU7zwbo+SdDvDPkgrrp24hkMPOEKJMas+t+4juECv3LTOl0Ebwc+3RoK66ko
X+X3bqKkR1zj1DrZQV4edDILqzw2BrM714hrDuXXaqddwsT6aA1lP8fVZlSwDKzd6ZMOIgRyZ07i
VhXi175S9GdkXmAvaRYj+4N05tt2lq1sswWCXFCdVLd0CZExGiHceZU/zpC8SjeAvQuk1EdhvE8F
KJfd1kUqqGUFFfWt3ceSC6UUak7Cga5rwau6AwSRybB2qeWh3gQNX4v2zFrQQ63PIG0iMw8hhVPq
XxDNoO+vh0mhZFaZbMYN+/JHfLSz1UTJQgAZ/JE+UpwTXlIxSFj8WyJCPrM8I39NKtj0Zu0RrMo0
GAw93UwJZxuvUuck1O/lIPVkt3CRlEp09tXvr8vvr08c9ag0TR07MxwuL3POAKs91K/onCYiZKuL
vD40p2lvv0wfXGOpWKGvniOQ+HfvYV23XH+KDnxwMwemR1rHxJmgsY7qkkzFwRJNVOQ0EYXRzE6P
ymomWbHgEK7QgU08BpCGXHVu17j8m0tvQeD6w/g4/mqtxacmgwIKoNT1OHTyScODpj2gClqtiHpr
TDjsec/nI/ls4i90JOF/4/Pgn9gwh6xnS2PYP/OnslfrQYbaN7xRx3l6mAvQ9dW2IeUUGlMbzzSq
jfwCFVmvPnde0PLS2FGrceBSvja0mvj8C412c3zpHefVjr5xYw1AscANXc6SDe/AN38rV/kuela3
ZkShtl09GlYsT4bT7gC7hTBRPYi6TPb0w8kPgUFnU1pceRWdP0GLq4wigViGMVqJg5REJhe4iqRs
YcJMcOoaGQWOqxhXKbF39umh3jqpON8QsGE8HB0aSQnf78nMSZls+UdKjQdNAbGJCnGAqL1v36Ny
nBr89HuWLKZdmuaqAcEF2wJzbSY9rA+jHXjr6hnEtmfI30vZf9VvWV3czAnep+M0ceBEiD2l+QqR
fJ5OE8e3aHX541UQOelKU2XrW29Gsky6AOoFNONe/OFX0odrt1lzcsNdEkF0w+j2gLP7t69XbUpy
3lfQxquIcjuaL5pqT86zGfMYUXgc2xIylxxdZbkSWWtkjob1gnFPBaiiQO/9s71UEvtNGdpkGe2t
4t4K9vxgeH82/DFr5lphczWZNzmB4LYe0EkOjR0/6a2V8PsAgMaQUT+M+Ofj7facGxx1oRUcTxMO
pqatACGDr/eQLDoUZfVi9PrCLVz9BzmYyqXolf2QNAEnxfC5rdQ4sZqPw4kNGhL5jWynlcnnanI+
n+ijVOEgGNpr/RThJ0x2RdKx6y0aheG3xCNLmg84qBXikHvf1wV/0PUh1ZVXt4Nk6YxBncoYdb9h
fMTIS8Of1CQMZDjGVKAMjHjoIy2yEv9mgLxtWxRZ4nkQ/0M7GsIqZ+xTj6dyfkBSNRhVIAvHrOnk
i51lv0Wwd8WSroaGj0re5o3JEHQDamva4/eqiQPQV0seXibQqmU87z+8Klasvt1h5xEl1Sjiy36m
cYQoy/nZW159eDtU5WpaT3N9B71vruG79EBrpKRoGOb/Qnarpd1943b8ldeBHbR9gX6bw3n5TVip
woUxiCMJGywqK/mYzAbm+l6rtnI9RZqYVO0y4IOwZJkNaS9OH+OXa6kOUvu5o11LfJ616fVbdavy
BRRRBBO76SRX2v6s4Zov/R7VyrvUy12HylKW/qFUrSna2J3TQVKvjVvoHdEuLoe6PJQQZUXOiGW2
ZLPqe0FaFChZiJNdU+cXgjizFsJw89N0pgJvItHVxrWg117g7re1spCCzxbnhFFRE0wa8us4be1D
7IGZOJN7wYAUSw0ntxSRHYl9pnh8sBwMQMmM1Hhb92iYR9wb/aTydzgxiyzMc93OkDC9MJ/ovRe3
4Om85qoWalgLovHoAaIQTICR6f0lrjxRxWKMHI5X5ooGPwGUjFAqopYLAG/q1DPmeSqEJ3H98+oL
5cOY932IyIHVBrrs+JT8lydX+ynK58PcWvZpCbjwY4P0tW21D0ukh99tz0JyGOUPNhKECHZiqFfv
CgaTpS8U6hkrpwgdxqcipuVUkQJMQpSJGj2LhQ62MZlDo49AB31hcqVcqZJ97xFKOR4jGQOeVdHp
LKAGQFhN1Bt1+yzIhXYdFtjNkThEx+sPcM4CdxNFdfSidWWB7+HRS1F9S/j9a0z/cKy5gcD/f0t1
WGjZYf2s+sR6uFsQqmyUYZbWKIt53ZG2pg0O98W6kxOSeVpEO1Ggm+llT+e6Bebbt7/IUdS4BIIT
kcwD9d6AKEar6s/Z140E9kvtMEm7XF4MArjvWpqI2iSX/9TRV+/Ks9i1P5EruA9Oc/khl5U6l75j
Ys5B+AGVJ21/9pAtj81jrvxCxMvsZLp6UgzPdHRuIHjg4xRZzO8YptOJif0GVSL8hlTMW7tihfJM
prwvgPNduFIq0H7Ocm15WaxOFwbH5tKarewCXtXFqxdYUxDufxBz3KVZd5K5kWiLLXeGSTy23Ggc
lVuZbAXxL+R20YmpiqK5KA4nbpLLuAqgGCudOQUfGvRI9a2mGVS+EJIGMuQe09H4IhPK0fPrJKQI
U7jj005UQbXcPxy5OicVQ3TFk7PpvqevDWbOiyQpcjIfHO3HmHulMwgqTV7fiBzR0RukGa3PvDtD
BmV00bqEMj+6fw1TmzEHdtBhq633pkCDzBbVqpyqrj+1iP/ajbZ5B9ppxdbwha3e4ds5WkyPLczj
EbGFMC4jjJxWjAcQogzO3C5BDJLvUjzfl1hqx+Qg2Dtq6sDMOC3HFwM5RyZzxNCsGv1NALuacLNe
MnaQxrMtNPHazs91FY2YAmuI9QE9/JPcJqo5fT9weMofRA+/jeJkrUikIL0HXpiGMk49wUc5L6qe
mvFD0jVYKCh953ZNUSEFE3+H7viETOOgpF7yQfWzfuBJYW4j03APlEfWodNlo3K3SspkEdnws7HY
zrJenmrlfNJc4I4G6wDYEkGFG+ZqlTH2Qi8uWKgSKduXc/6njw2prw0VEMdHAmQutW7ev/koC8vr
cb2bLGUB4V6LUuMIl+5tlvFJ4mT0JEnw9R2dfi2kmH4R7aZ+opfScc6wEn6i/eiRJ0Zjka26nMeh
jA2Hht4dRaQKICFHsB05qER+XlAgHVmUkOoKaI2yUjVryXmvn6HF0YuAooRXpaa+fOMOPzy9rFCe
rAWlLVMziCE5/KFKLUMU9I5N98gen+n1BEqlKnJs6Cy70O5dOxnPWETqxJGg4ANAT70mzmBD5Lcp
kWFSHKFafEqTtpPsltsffcAs+y9s0VecrgvL6jouznzOB+E3pYZONBHlKYteePoRl3a20Aon+Op4
QKDL/Td0xU/aYdRSpgS4xuZWEiq63TJv7ZB5D5iYERaryCwNTIiog8s8Zwtrnd6HQo3j3tkaJe5+
4Qnhp5XDqcYa5gRprVz3OsoTxHKdID1b2eYZWtSHJJRQa4Ew7Cy6jMqiXugvX3medfArW3ecC8ri
AU3Pq2JGTNtLujcaOZXUufMNuejmycVDnNa35TSGJhfSUbC09WV82P75+6+6dUjC+i9bT6ULg6Br
d8i4vJEOMeEMWk2YRY0e4IBJ4n40EozDZyY9yQeoV2z3C+8JwKidAXIPbybGQeFWJx3egJ6jVNfX
CcvEy9UOQLuqPdAnIK/XQxJ0s8eJZrUeqyhlxfraqo38BD/PtyEMtneZdWGHfgBd2AI8U+6Tz9Bk
UW3SN0DvWVeHMbxApU2pAeg8H020GYCdogJ9TVBHN8POEFIehNomUKABS1zLKTirih13fqj2TqtM
PmW/q4Fp5ZARisYzPy0RoG+c9VWpKTI39fDwOYl1NMZTu2D5jrJpN/0RE7ZtC9vDbnnwAv4nu8Yb
qPpZ9FNB3RwNLnNFIU9YZfULiYsd7tWeu6g0CWyFC6TI5as2cPiK7zsP4fGGJg8tcOVJqhZR5OCX
HTxvco7DAg4O/WkQfKR0uidbhCZNu2FZgPC2AHx3IzrOYzZq2jY1LRffo5LuzZg2iECW0M/WDTgk
tkY7/WmhWivksbIUEAQ9M5FxZa1ACyoh5/Mg4QN4XSysXRh7UwvfIfiUm+G3j8o0gbqsMEWg+MBl
jX1Ym911UFH+i/b7CQqDqjsHuzyt6EePaoXBM+KALgalK2qb4EXh2R9g7mOcObPdr9D7W1qK1211
Bhe+1U6A7HthzsQmuRScTrefcMvnfzXRhWIuOCLeIDcYp/7+7DCcJG8mIJgRKvLlIa6IhiR4RO4w
DaOOL/GaIzjvg7jFm4QQi747GxhUsRhulTWC6ogJ3gv3cfkZ3uHC7I4cReoDFLVEwaxcx2mkPgIp
0pz4BC5X5vXaXdrr14UqDnnRZw7SWCQ90nJKV7hM9/5474xDX+vGb7YJBhd7gDnA+hG0sWpXHZFB
e4KkhefgwZzF06ShIVpmYtKy2XM8boQuUqWO59gKfT5hceKJdnyaa9s1rVoY9PYv6pRwIpKSDiWq
/W8cadYls0obQT1ijB7yiJd4HVGKM67Rv/yWrbHFKRgp6z5aVwv5oV23ybW8rcpRZTg8dDxr06WU
sPDBQ61bvq77Vnhj7laicJ3Z1gsm5cbuPDzq1Wz9Q0HehxRRGMdgsM99ecuj0xgWs7KowqxmyHSy
Z9vUjUUzxWeYX8GjNBJQKWTuEmYSZ7J1chRHVX5Y1MPfJ6U9dsgRr4PIHJDPWtulx8w4723WTa/3
f6eJ8I0c2oi1fLuVqieXJ/F26SwzuG4ovwuQWu6PXlM9vJO1E8SUWPwdXwpTUDwPoLsiByS53Vq5
E1y03o8sB2VlIhEnW/W4kiAkenDHgmNNiqCAIfwbksIPlwr3SHGFq/YSccvyy1yBIUX6peUO6qpp
+WSFbksWGPTgIdgkjq2sTTen3v2F8hJVaAq8zyvkg5TcoPZiahH9qhQmPfqWtsxLnCx/sn6/eteH
Ly/BoXKypBY5/zhXIJa8WSLLOzk6nKOWf2NHqno7WZo/cNAw8saKbPtEjKq036+YJBIw2rUWD0vj
kS6Rg+6ppxeUcrKKOlua2/CWJyHbzQOwJyMYCOR5DWSr5frHeNoRkPRQNFT5p1+jRvMDeNkHoEkd
XACCREO5y1BvQehAxBgV3+X2LKDsCd5q7pzc8nw0GKg1KWy0ulANzpypaPQHwat8lsLAe0M4xMHb
ujCkZSe21krQ1lyE5L/tJaq3mJN7iexoAnJUoHH4QPHGg8qY0J6WwcaerdjOAHyLRwVtOq+hnJ5G
kXyKBJmatpWsi5rJndz5C5gQHJiRFg4JupIsMQmTyKG68e6TckBQxkpNCGZiJWXWlNmtQLPQRbua
JP5NB9DO3z0Kc2mVJiDf/QuHPEwOLeAhblM5ZVKssosf6gcNICmgnCct93q0UgCC7agn+z3/R/5t
JLrN7qSoej+jvrx7XHgrDsWuzOtp51HbtBxYBjz+Rfc9/53obR6sYDca6zLkSmQNvL9AhIQ6QEno
dj+HxkFy+TTHX0r7M4kcuwLTflLtEZcoT8fSUJtGHUIXioamH0Vs6xuYNwBc74WoncTiFgea4w54
xFBV9CWpyYK/0X7NUuT8PrNrcJg95OfZL48h2dbotHMi+e/JW0A8KEcyCJzA/x889FE7L8Dx8PfN
TdMGD/rbErT89UYnAovk4gT05xHbT1uw9NADjgWGze7K35taNF4KaoNAEHPMTi9+AolzfjBJVXdx
Nx35Xgy4rhVdTXOIwpH162pvlxX2MN+tdD0g17rswPXFrdp6uGMAwt90Q7fNKLPf4Sg9auTiryQR
I7Jl07easiz2il32ZaKwtB0c+/NtyvcNZRhABiwXqXYiBQk/tLqByEJ5NzXqCkKFIRK6mP9Am0Kw
QvFMuIwW35IwVEVUlhTDOZYjjRWGjaCoIfaebVntZq0tQvKRKm2g8DYlZ19vdziqMjLy6quqjiBa
3a2uARLpTMhe7vJaeULYWFWNqakdjAWY5n6PQNFZXKgJgi+gD0tI74PW7TeJB15YzzhYQCldqiKy
am/oJyJuWAIc3E/10l8a30rSIvbNzb4TWGxPJdNtWJ6XOmhf+IXrFKIFglFCkRyM5gmHbFRMljp8
M5VKvubA47/4BS8Ep8V1ylWcH1HSTV2DA3s7/dnmh2lPhnhdQdOqG4n8O63zFFw4tZHdTDaHPL1p
SmAmWEgzpeaVh2rY/ckRjLg9FgCc2xt7b5hJF2MgWP8YrQOtoWcRkPu9nxDWm4mkkV/fsy6Ue+xi
nrSjcjtw8Ehs3kc/nWVf71s9t+NRevXSvjaC5yRNbeSKesFVsr+ruzQlQrZRs8cPwxqo3RIFiELr
v/9zv1dVx7+iQhjerz8khCoIJ0R7lUWUCKWnVpKCgFy7ZeTwHgXdqWnvNNweOeveJmLkl5OXU1K/
t5rM8COgp6w1W1NJFh8jRGa+AVuZHwiX7AfoulPjSsFRJaN9W/N9DuJd5DBKxN4rikBj02pUM1Xg
WtfS1O7OekBwXIwF7YZueqho0Wnj59Dgvzz3W1N2OOSh3lyOPGXlMOXu2eBWaRtUy5471ZnUXYnE
LFyWNgaUT7oWCsnhVknSFivnxk++SUQxGkX6VJlajfzJa0I7l1kgpgE+tCy9Wv8W977UGtz2zHX3
VWOnjfWXul3Kz7KWI+PkOwhgBZrd+23kqQrBz2MTXyIJUIGQVru7JxOcassFUdkrCbhfNE7BvIps
zQtpNKFjyhS3HgROVmGe9md3gXSSnHQdnz1LJgk7KLL/cmvdfkVLJdjQfApzwwcshEZg87jAsNgN
vk8fQefXGGRm4kY8DooDKi8g4Up1Fq1C+V+9WzWh/snXTeCNMEIBoJ45LLcwMHUVNaQarxJfPVLz
bYpIiYpuRWSSJyfdzMCa56JEvufTvWFMFjXLJ3vlT9gcTlURMCXuEIzp6YY83waHtsP+WsDpcQag
gg1RGJBLZWD8bnnfoyeV/QXYH86aVFUxK/lStHVqT7HFF6rdyTVJTQ6ffjmsQXNibNMUP7SYLC1M
lKHUb3ADL24Olqfv6Uj8j16xmwBgFCphSjLYd7VESBL9O+T2xYeOfHsqH99qmgN7tuFj2wSmBPyf
o90arRBK8ka429BUIX/gsPT3q0DL4aZqXc/xYQcHuThDpPSmyq5OXBMlrnANorg1FMTRW3nm/AS5
vk+oW7GMJcb0xD+yu5VqWmevipfWCJWyLKZD5hpKVDyhfhwnwB+sLb7IeFBw14BHt43vHDd3kue0
WCSnlX1Ui/cXv7sw4VfLcsa6DTJbbNGij3YijIeik45FPHBcs472DtWpwgUe6YiydfI2Y+XcTGAC
uzThbKcwqxf2Uz6pczqkeiX9gHj5kV4vJI0je7nWpbUCPQI1LGASlpefKO0UrUuzYbxlSFfCnkU1
s1JQTHEMk73o4S5pRYN+kvyajtLYFrRCp2w1fnqjWG6KZnWXJw0a34OsmM3POje9CdsW5Iy6fjjE
Z+d9/Gjj/8yNDFXHJ1klNzdrP+PJdEe6/8AhaM8bInTymfp7day04EVVN3bBtcxW9Bo6w2dGLfmL
KSa4iDgNH+OUyI1Z80HVfHICCgqryrSk1hPDM5X079rFXy2k78ZyURXcwwlepYxb9aWlmazJJVqz
nZJy2lgCua+IlTAT6iNxS30eR/EI6m0p4Rz+2DCUVCaSDQUsLw3/TPLNe9yKK13XMEdtOSSnSU6p
h6og+wVrrDAZJKTTYDzTSV11b2GteWje9TgLwBn7TMhn4cQiR/1OmC8mZFgFIWlFMfjSXhFx5EV4
ifVTANbGfaNZvpillr6kXJ7BPOooDvuKxzxTWH9L54yvn8ppQgHaURXLkNC3RN7ftvxRhmkMQJIR
yKcAOSzsHDJA4hKvp5dVDqAE+N5fGh4KFi1WJms/2P7TjgwFLZ3uK0+gHBhhoHpt0Bu3kb0GcNmo
wUIcYWZJSDuAvHUP+pMg37v2E4F3ukHUq6ICJbHdK89HaWdiouPqjG0AsIOJfTlqOqMtshmINBt/
kuN2CspN1PN8cgIU17FoafAb1cCgo8kEihrtBmctPzMnC4fnhlAr3Fmf1bjZowVjSdvFCJfndJr/
QLFLk3SV2KvmSJO4gswLguX+hFrJWFMGQrHhIwiLqtFJLuEKFMcU1FYiY3Re8wmiNUE/2jWQFmAX
kNGOw+7yllbzDROIXr4bw7/CNtlWi29r4MvOHQ2KkUkL2CYkXlBwuSBE2KKUSi7FyKRsDc6JspJP
VVpcb/H+m/cyjHdyQcM7WBMlv1A4ucs7BY40KgHPO395fVcsdrE+8UGO3rPENKjlO7w8AaCvXR1Y
bQKBk3VAX/Sf9SBrfSbQs4UR9b3a/CTaFt2oW6wvB85gF6h86u9mB6Vo4wVMG+O/JrcdtRAv7yyX
Fi86dNTjF4VEgHnw/w43y7GZfUxAa8bxLCiDG2LNsnoFic4UJxyelNpr1P37ccqDRyu/0L2WAuQM
zW+qoMjszunGePpfWegEiP7JoCxHu2VIW/rKsF2yIl5LDjJFrpxB3l3uD9weQCSiWmjngiExG6o5
1jHiA7gFbWuYHxEUtioGDG+WwoR558HFHZwALpgd789hDPsrBgOrvjkjoShADjB3dtSOSf6h7hYF
eVeX/8A941mVEzunMTcMlEubMyRp189hw4sr4MzLAM/kbybPOybCGxLU1gE3FnUWvGOrpHYSA8Ts
0vxyQO/H7PNuEU4P++XInh99PhJkwQhSjz9Qr2MLSU52M7irqpejS3B84eXbu6oekT0cPlFv915u
C1hhiVqDrnqcK98ZQYP1wKF/H3BLK0A0oaleGKLg9LwDtIJ3S1gNUoPu1yE2enPr048nP8guV6wP
Xv2m386NwIlEhaCX9pV+aCg7E66oR885sbaN5xiVzghALwvnUnrvwAXPIShfQu4JSyCx9myk5SGj
0L7/Vji7o+Ycl5x+8PPoQvDpaherc5B62tUPg07J9AoNMC2PaYYEqO072ePjT4eEI/aSgJca58gO
pmQ5QX96rgKdb2MWVgonX/z/EimH3JGAvAxNPKnzV99NiNboBN+JZB3YiNILBzkec7ModqoTk8Sh
3s8rpZOKgOZXdRPJBfKuqpg62lJBl3hevWmk6wu7oXBEbRm7wT1p7SQdjGCaudZKdRyxnpQKRE6e
sVd0INeM79qCSRJew5tJTFwZbxPKncow5aAPsLxELQ7B7DwfK55M4jOqJ8LAFXPk9JNK3nAQGo6D
opDoaJ9wLOhe7bONGegjINXdFNoN9xXpfmMSFwiGsbmfCllqP6zGjcHccr7YtPJULVx9Mn5Cvs/A
mnUhYuuyTLZgZ1LsHuyW8OmJ7YT1I/kTty1lV7QhOHHERuIIvxYq7ejEY/dMB8F46L1yJ1TX/nCf
k6tC+u3YRnWTcymGzh3ZJYCVXNeCAw32MtNvbkco6y+H6FbdNiyYFBW//ZWub1Z5nJGNMCDr/nHW
CJC80LJxBCyL+nnk9oXoXV1FuJExyitdQW76fScct7F1tJuYSW23ZCuaz7BXH6T6uxdxgDopSE2S
FiYBPXB7e3tCxA708jja6amnNmOE66gu9ZLo2niT/GSjqkTbbI97djbQP0yT0srXxPcVcRm/N26D
Jh8tJ0L+0WYS/jXqPxCI3/rnHfPa4TBF0SMKnS29QFj4CRay8cRVyrpzuGrdwLIIu0BjWFM7h1e1
MXaH2GRCUXjhqeG0usOsV3iP5REbqiJt8rm2hQaTkgP5sRb2pH71Q7ErFkjNE5V/JHZ8K0dVDUkw
XFkJZhomWI1BTyeaGjBRtkCRy473qDfc2inZkeHenb6b3O3FofvFrdxpukczMbtFzWNBGXhuLvre
j3KSbW44AEIrawcVLG+HhJDArtB6pCA2d7BVne+TLQeN9oukyfY45cSiyvRLbeR1ML+1Pn7r72hY
V0ESRk5TtdFd7qby1UlcD1H4VkP/+1snLLpVbpLh/2Of+Ol6J5V1SL9cBzhPoCGYkwORegEzm0AF
CgqAXO4wB6DM9fQ9BZ5gQLoVwHvlz78F1l/fvJi6KX42MF3jGs/4g/FLcv9dwLlxmibXo9kkmnFR
NwTU/0t0xon58lL6HHjRm7AoT4od7vjvCIpND4vXcW1Jn1dWqTmMT/b2AtSDVj4KbJ8zAgHAoyMN
kmnj7OagPypbinDrA+0k475ZwlAVVmIO3mohfgrbDr0Zr2P9n/bXIIX8M+AxM+nKezCHMybEq0Su
FCfqP8HhMlH8TSTRGAxu0I5/qjf5QkTwnPYq/at58Rgq4dvMlkDDOPYe0TTh9ad1eH2R6O+UBnqo
osywiVDBIcUdqnqwi5sT0JqRhqwwvGtLoCjUeuGD54aWcTf2Iqhn1mDwfn0fV552z+rBDtkjmUXN
DLMR/X84ztlskhuvQxSXl5E0BqCneEDDUECyhjxOx1eld1vxCNzT5Mb6wtplKMne+smEzyYc7MdY
JkhjXPVMTzayGzEefWeck9gQB4el+nhV3YkCSwtbe3m05otRiBoU3X+2D1b8Tfq8DvAT58SxoqM5
jgPIIPj+jR2kh+HMcgTPogcxKPBlhH+bIstuoUJ8SYCdds2HjlkBnuH90/gzCqdjFb5bzDHmnnWu
3gF4az3Pkmm49fP40cEYciMNkhuY0811P9cJ0IMDXFs0h/ilXgRqPYeU5aaRAc1vWYu53A0/XZeQ
osDqZMt/N40p4uddv2UOJIMjx3GAu9/Lyln3FI7L7DyQ5iHOjwCrfInxY12TJNHyi3tEHeyHrsJ2
igvyCLalpD7+ZlgeQjWlfIR83HdBilAf0NaiFak5duiOXmNVBk8KgoFbkeMgKfruaEBDQCT8gI6b
Vea80rRBSrCnjPaXxhKbIJs1eT8tYCCOsVzOTLnXH5zDY9rPxoJ6ak21ySqHaSqLLBopjuViNeLK
qO6gp8g6qeoSgh1fp1vWr6L9Vca3E0DwdVXMuyJZpNwySzjDRG69lm7L7g/qTgsL1wAQO9QB95k+
L6RBRaRDqKN+5cf4mj33vQs8egxFVY+q8BtLLPK/THhUbp8ilNdkFOu9Nhx3DucE/VBG+yrznB5a
o5WFG9zO97E+vUDor2U72StGb5Knh4ntVdjJf2INpnWr1aiJfH/xPGPjCCtU8sCbccGxR0FYjkxG
N9gdPTOiSp8OiPuLjqvchlgmovyPR5pcBP43h+GbZDmF7Ca3PB21OXferWPo3kuzxQMIPv+ECT/u
gCYz2rATk5LDof+T2Vi72LB9BqwyJV86jNcToN/VouKHuB8qJrerrRYj39c2kgJmlrEaEvNLuiB3
87i5zUzvoX1saA8KLA+hpGtroX/up5onIMR//F19hnzMdStN8D8qUskkHj1PG9eNFuuF+GX5ziNv
m+4BsnGSJdgEurJNvXD6WES6CZH5KjMOaUzv5kBlRF9TxAGRICOkosvPb9me6TBD0eU1MIFAhysV
AwZ2lf1DAq00goNtj3O3LP3wzvM0nf1/kSUkj+wZb1fKWSMfORhIzd3Hq6ll3tbiK2EexNGiMwpo
qAi47u59w+VRVwGMj4Qv3suy5N8lXvvbogAiYmR1kPuDWp5Decb5Zb3IsAUw7WSvzkNtR/iquBzh
Aq6tCisqcT2KYl6u0+bZ43WDdXkEWZSahUJo8KLDBKQKhSJqcq3hInW/3RiYKx61ppr58vBgCoI6
4YRpFeBE66X8hqnkqkQEGiJDKzCMDxEfsMrzG1xhKqRDLSB7mvbnZPQn+G1FHpLNs+9pTrvzMyC4
Mj5paP0+N7Z2LDEObroqA2fqguD4psKbq5lYfNiAGX1LzxqCywlVlgndqxqeDVxvfYr/JxxGgtoz
FdWD1IKHoKAqBWEacai5BVHupMEner0z3kZYOmw+ftNFVbPn0Agw2y/PmTs59djUILu1vNnYFImr
HVffelPkW686TqJuRyTjr9DvK5oGcEDM7zSa11cbM7Ouv/UWHbyNhZLcz3pRSkqT4ULYGez8v3FO
PIqiEs8HHvAfnM1gk4GobzhRhBlnlpfq6ue6pG9h++XLYIgVGLD91lZGQJoea5usjEQdeuyuDVmO
4JlgA3SToHJNN91dASkIrgJGu4khaPxu6uGYkj9xTaT2L+Cs3n2uBnviYdAgXGLkCMIS7qaR30jc
lql8NBjOMykjazD0n9GlRK7i7kKRxCZFCPyoyDf2ZC9b/y7IHsXPd2x6trLjFv2gqXOqyh/mipZu
YtPxaLKYLXh9Ibe+iim63ab9kDEEY/jLWjvl4jnatiiWe+qQXxDR4sRFdG2kvHAtYyKPAcYOvznv
SIklyKeMk00+1nGgrPnx0OcSWWTLbnyqjrszdpdOfRSQuYirbOE6pVyhTkMaIPAr/6h+cDb9pkHG
dFoRnLP/aeHSVPTJFzm1Flj6Zlbtws6nLq5nkDcZ5cBdyiJVOb2D7kbS0b7sfDt6jObYUPC59UaN
HnjKqVY/p8hpyYLTyUwA5p+Mp6FHalXPVQs3yChcnST1Nw+L+8Ls5vWlyO1ZZ2fKJZyxH8Wso3mt
NLrcviGfFgyZXhywgiqaSej7DH2ZszE3ZTeJrsqMBWBKeaKrejY8CsqPoGjHI9NSah8Uiwk3NK4v
Hbgpmr9uapM62kJEiPda/fOgNTEapVpKcc7Mm+9iA/CS8Rj/5i9Fo09pxKiNZ1/YHTTmGQw261eJ
aNt8xf/h39YPHXlqSwQDBMHIhQOmfUmUxyn/U1WHw14hlZQjeqvjccwVyx+8Fi2robYSuMEz93gq
j03uEeqS5HRvYS17YPogsPbwtTJdzPRc8F+mG+KxZWC3H7iv783qhHSTM40Dh+Z0VZ95hCCshNXc
tI9fxV9Td47x4PvgeZQ3k4LgjVJaMulTU17JT30OejJx/fTjfmkcvOoS3OsbN8+zhqPqUYqvhzU+
VuSTyVPTrH1eyKqoZzwPMHrYPWlD7276kXhAvJflZYIKF/Aj5Yr+jGjKqUJDR87iiLascMfisiHY
pUkdT0TS/C490kgRGWFYDBygd5TP8VWy9wHgfd2cdXqgTaT46ACh7u/P2W83vlxY6n8MkO2S7F8o
X12/RGP/m1zJvgArO3tOsF6xfM2vbwxPNw4ucjyeG4mn8seYXEo2oYDIiD5CSAgjP5N1hyAxMCYd
HFGLiiR1YZ0AltizApDRQONxo8SLPt4aj791XPxcnoF1jnuBcnxLGJo1P+/BAXhZnyO/X7ZBnHJC
g64RyoqhLWQ09LnxK+u4sy7NFr1/mkz6Y3n80bIN3cAHPlYtgXzUDBbhpKhv/rjQr99OekXFhvWZ
+FaLGpYlPxrDbQJMRnQJBCYCOxkmGE7ZtIANh2OVXMQCKCskveTT+MSYVIP1q1b1mL1oUP+8PGUL
vVdcd//ndbvfcHS0ndxv/LcKtSKXt8MT9N9RM3nrKMmGxpNBWFpGkaY4Bc8A7U4mwTI2w5En3Zyu
FLQjRODKe8dbr+6Je/Zwi7brsMLcuSIlpmVlXhvtUW7ESYmIQ9OiM/65yHsLGlgYO7Q87X5bz5xB
eTmQqrCH87Ag3wsi3GjBXyilvKPYPNT45BdNiXzULTBanh5mRlaKgxIphLQRtOR/rHm4c9zjK4Jt
MRhsFumXWNyuEjH0io9gA9gMsrjfmnjNvM7z7etA/8iz0PXqnO0+0VXRqvzCESkrOnDUgnTYzHc7
2rz86FRjJXriIpeNk9XIr4oVE01ThvyYer9I0c3Lp4ryojxtxnf9HO9Ot+7wpTOcayZ/T9LYxb8h
KyA9t1e7KDgidbzfpPAVqNcuHzqRErxQBoCENHEdSFQjBQ3rOzmxFQ4dhTF5jW7Vfw+PtDONbE+8
icE68fE71xftCZajqsWWKtw5uqxya7sBYVyfG2iYVCdxNYQQiROpEYLD9gkPX6T3ZMZKl7sqB9hZ
PsO306H2nysP59U3v1fFrosikdSskm3T0RQiKFU/nyBzCJfrzTtYD2IH0AuVbw2j/loanIdzVgPv
dp6XbNT+/tCIC6iw9adwUPb9plVvbIvt5mVl3nX1bdU1t4+f8ixlxaAXFBdFgSH+5ApxO1hdvsgY
14LLpJgKtQLK+rVMK2qxcJfxqmNBd8SCkEUMUpCN8QqMREVQL7LPCRlxI1gGAEVkCwNry1xC3rf+
ofXQZrEyYtqhEvbskpc2dFJ5vQU7p/ZGMeh29CNUoUPLK6bSlz0BdYIXLg+Z4ZmCFofrXCYvKugo
hb5j3lE1Zmt0Xv/duMgawvzYOhw57/ClWW9dIQiAsBRDH6Zz5LJhaS1kNOvNJtjLbA2mOkGeceUO
wdPJN4zu9TZspVFrtxkP6bpA9PajA/7QuUdPW6DGXSZgpXiengfEUF+Rzhecg3FIAnERhPk4VxIO
hLQdfWFl27ilmhipdTa0V9ajmcNmFgWdvpiB5Opgt2yJBtuke6XVyZw9GTf6arquYM6xhTMMVxxJ
95GV5ONcYsyncI93yzd9i/2uCnD5VXJ9Yd+gx0Aryt6e1p0uKgOYHULZQkVLFZBDheynyQQK7AF4
U09ITMnpGmzRqEcBXwMvKHCcytpe/mXpdGppCGiItjaCZGnSV6PAHXAKyvr1K6Jy3L2azmhoG6jb
wxHtzn3NR9ENeGSr2xrf2Rdjtf7vcQzu2HWh+CHqqkAaUGUuKnls/yRa7dDyNz4jFL0IhK1Db9J+
pVWkLcoDFhvsZBykVoO4wXkU9HI2VdgimBHOJbjI9n32vsuh6haMcCfQDb9fYTauSJ7Bo2vWr+qR
eldry8lxqy44AFUKP6Pk5k+NjwRqAzl4EEYwlN9TYr30q3p+qEoAUKWJoLE1uW5wYx6YS4XKHfVu
I4DilBZF2nkU/XDXOX1JMG9Bz/AKVYbH/1VxisQQ5/ckGM3s3YMQwAfXmYgHVZxf05DN/XarYZg0
f1S0xlhoAdUaH4ovaCCz6hqoi97jc987oMjiA1H0tGIVVOJF8UP2rwPbvjvG10rEwaXdyOcZcJDn
0tCGdQTydw3VqMyKtXPDisxCIIi+JqPThNOjqq8YyJL320v30S/sI2bRZjM7mHsAwmmmfWkdbWHq
K/w+DtC9MXAmCK0myzTCFzW7ELMveA+TZfbO5v0BmU1nDV4PIEPmkr16rb3FJILe0gdzEF3ZlZBL
0jcV05+/TvR++/toh6GpW6X47ymtrjXXzVk/QOjDXk7zwRTl/fmk3OrD55bxRkWxyfUExwRNlsq9
0iaWfLpvXbgRKLfIrMJL8X1jECrSeYQGxZKGYE2Q4RhGNHNfGPUOZrzUwty3IIUWgggl1rtLnX8P
lgezywLogdn0FXwV1Fgw/qZyveGb4lAyPhrDRbCFGFw1L4mu3XyZpe8QL2wo/fyH+4V1qF93OMXU
uK4ofc+Cng8GiCxVgT7G5GdCN8GLSr4sMhGHG/dYViowTp3KJIkcakibFib8anhK70Gg5atGgdsJ
UJOfUlX//oAcPl20vTfqPr+901HbdYz/RjAd+VObK93SbW0PPOOwfeyJWCv/8k5SatT6AShLinXE
6d+4p189Uz+egd8bwPHkVT2oL8/90KH649I0o7G1QDvUC98DTJpRg6fn36qwwwPYMrKt/R5EnE06
wTiYvVDRHBlmIazo3O61hys9wEOBdU2qrpEHGjM32+DFkL78eyxZbmCeu8G1p5otTdhq/gmfGTRt
wu8osmoyD11g6dPNtFVTPF1MjFxJKo3G/SZ8/qVLQpDuDAR69rZJCxvHLiTss39U2DP+nN97Lksl
I53qwh78KdO2DhzRT2PpMLnamlDYl9Wdu2qANDi4E4B04JyyY1GQIXhUe2AJJKELfBmZawTl5j7w
seC/liD1hFY1sKcXTudtaPP0XzSezA5e88YEDTB8H1eq85WqZDdPhBp8rKn1K5iH5NEnpzefVHa0
Wh3KZQ3/QnZpS0Bz95vKzrNGLgYbcvJk/x8+zWTvwKiX8iXauePHKtqdaGfHZdIcJyD3/l8lNq+i
TALkLnkQGN2bupe0j1qIunrZjATU9FwJSdPuZoOEI9rKZgTuQSH+70v1tsyp43/7RMJtu9hsnoPv
ntZgGoviXKDsan7Hpduyv6PTHltsQVbHQrYjW8ZqBb9vEe0/jIn+BPegOEs0MGHqLcJ0rAlDnyCA
0LHOUA1QDYROCNwf2W9KgdImeTL12LQrxLYdbkh3+dpqv6FjZkUHv6mjOKcj4LlUm0HUFov2fuiA
mbrQCwdVHak0AbpMx+GeHlOwhua0Y5tUN2GT/rmsq/tqJaVmnpiB3dmNt4m2Kgvf7dJ0J+sIt+/g
S6ti0LX8dOJ+PprF36M8tEHWuHcU6fbWYjyuHJ+wQp8hD5aAQKa1ymVLlxK4+kc8gSC//4gYez9n
hn6i4Dr2KsSdp9xGpwAjaUT3GUFlBqVQddl6g5tKQL4UL3zHYwN7sOaR08Zcqjriwh5MTTpeVGPW
oB4/42VuSkNUHljFfDc4/wtfgp6gR695yebHutB92T/snyNM/JYCaeByp4y9wltunPMeiTDOtVNd
ZqTmWvurDJgxSidsOsWHrMUH2n+fbButHk1LPNYuVwO7fSmcp9ev2Esq+qp161nM5CGC2gBXEWyI
lKVO0oVtNm2McKRkhkoK02Oansf07Mzp1VRUS0Ps7wVYmTPaMq+k3LQyIFO7UU4eiC0PhBT8dAch
WqOez66/g6XdV+HfihAXWK5uxL02uEz0R2qjJqUJRdXD0C/PK5X6LGyvNx/JwJGOiUggR5qdCeQO
vJvO+AH45drEwDvuJxy0BZt/iEi7VVHPYdJG44vd11qehaZhsIUz3p9ijUoi+qrHtpCq8I6FyecL
AXkMyty+iXOTngfTbElJQA9UKznkKtH8kfoXhky8+C7mnzSgtFw41H9IX1coroYL9ekDJ0F0ugni
EvQqsBk95VxEnQ3f1/gNo9ajAxf+ysZ2G1vvyFBYwhiAJN30XEJGqXXgLusKtgze6Jm5xgOvoXGf
7eMKWO5ip61jzSwLzXni8dVZz5S6yt+MF0jUi9TM7c9+CfllNNUg8rGHJgs4QcfMOZXfQ1I5lzBj
mbSBm+bmny9h0tkRCmpLaF5CtGYTEL+3wU8E6K1q/n6Fuuh5M4FnTbZpeUtlt5B4N/4UX9j2uMHe
A53p7NiPkjTX1yYx1bA0A9cBKDemOb7X+zKWRejMhaFOsugMM/hc8KFZ3okNhDnQgRWVAHTR2AXk
sdye4HLH5BHGq+U9OPeMuJCjUNuOYucQAT3dmbKNsKTkFqA3ZcqJHMFjRKCrrToZcLxB6+YZ7LGi
skmY3OfzRx5ASvfIcWUwXtQC6uj7mM8kkA1u36qKgiToLyofsjkT3xZ81RlrNj63ZkdTucxUbFGa
q1vMAW66WQFE6W4xzIidYL+blMMo3sa2GoL4Xbc5kUCow/p0KFok9sIAm3lTc3KZFL09FkUyUj65
uvZ4izVQUCAANYxTNNU+8M0lTMn41Ex5RdKfUrgcKDE0LvIPcAEypjp5TXO5VwP8lQSzUR6tXG6E
5U1lIqmvQ74tW7Npd2WA+UyEZPKHkdR/fPHPuzMOfaxXjQDCPYk/1sHMKt4uGmsKiuF5OzJtuHQ1
SJOOfAt+hZqO6xwPe1ATwyuPWkUSAxhTJMinhazau/ZYxGjSyYhShXYhSb9zkovB9SXWgMdga3Di
Fuzx+iV10jAU2pbicPdIsblTVk08XMY7qEN3KPLMEkmcYfua2OTlNNrevuuNEnNU8iToXY5QhnQ/
UKVeB5lqEiIof5S2jwvk6lSeo5o0srHEqpMEzyAUul34xaCBDu1vhUQOk2wDNeaUb7ZQA/jJRrKi
YEAFnShv2iwkVAoYuU6Phc7z2QVqnCXmvH+xjglvWTYcsI//Q7UgtPrDBFqNOorQK0l4eZ6MdJ2H
ho04N0tq7+e/cXFcaQycJV9PYjs3H3kw9kJtOYtKST5XHeovpEziHxVBsW+yMzGpteK6flM3yKm3
qQu9j9LFcacIGzTfzd5rbQdsnSHGOHY1xWl9yOpQCOBPhJ+Y10iX4eO5rI8IochPm+fUVNUe/rK2
W2aBpF+BgZnf+tfdXeUVnveI2clUkKuHNMbH1aAsCKe1SsOnvapQv27KBs5YZXDCUeMiJxA2DVSw
R/JEUMAQnjs5QKKzZd6R6ZRsOrgf7Kez6QuK8AusCEqzoAbdXRV3hk6HEaabf87w/1keciEzylir
YkJndrrEn8k7hhPvmmBGftEP21WBygJlPuTWJVWSEJQnMVL13g3nhDtJpoFP/cbvkcC1ir8nXUJv
30RKm0MaLbJPYAo3K3vapxuL8NXr/W0q3mJiIJDdDmPXG++ojuKpWTED4VitoSPTD5hHSTed8oSF
ruGZrUY9d1mEIidxbPkq5G2nJYOHMPtbu+tv1numfZXc2t/FXmaYLe1cVj1ic+eI7elwog3y/YzR
hfx0DYhY1xK39Xd0qo4+LoKoOFQgJNLzmldcvXINyfbNdp5Anrwrcm+UgB3bdPQeEOBeOJ7HXcv4
OafhEUKOVmIT4iY7AfnOWC7Cs8C/C4XLuO6Y4YkUkCxUal/U1N1Cgygh+qzot3FRLKI85bCeZHa8
PpsCTCv52J+uU3V7VcF4NJwjAeli4c5AZTsK934WS/fiIgXQYF8Jw41m/51zidAHXexOzBbqwA6H
Y63o1jUdwJ81EzxhEe2e47RMkU2AifWQ9IE+ABfCRbqyGd1hyeOUZ2QX0YuOvxhKJyh23G4yPOP/
siK1WFEXJbTVlwTzG7h9D/irnnuZxwUIrxaPAJwRuuUUT/hRn3wi432WS+qq8ZIeazhWjsxGLBAA
Hg4krcHHpNVAx2S+c/bJupkKFHmZB0CwukzA+EzZ50TUgjJhYBNvpZlpb9sJ1ym8NYWAdHl5QMsU
PfW1eY4H2osiKkkDt+lUmARGh7ENhrNhhHksJy0KLLhWvYuDIMqC798ND7PR36jzY/+EBSifPg0F
lYHdbVeOrf9/cXv8D2v/+32s0amhbH1KXxu+kyZb+3+YHtUQwj9ML765V6wK0jHbcSSqlJ8zoxLf
ncOS5XvVK1zbRZfIWgy3MdWanB19pRUGDBBX511VqS6v4WsV45qsytxfoC2Zg6QjBENRjMXbysQ7
+wDVtVaSKRGavpoYDbnoEpMHPCVnP1n/om71ra2z0szrbqG1r+onUNf5Zf7k8L/kE981+PA1cFlq
BrqaPpq3zjsy02XYgr+u9cXDY30DxAE80GzKAXqCpOw1dEUWXqP6Whv55UVZClgUUAjwbqkXAvp9
FZucUHbPQ9Kq+xaqBE3ZcbKyGMzBEwWZMdVZ0tEd7QU9EZg4s0CFPj1Mr6k7ejOcQVAfk10QYDcN
0gGX+BhxKyugqWubxOIGdQ+jji47BCCyNOi8G1XL7P6GaiZyeMwx5Byc0xLPtSbW+BlS13HCuKuS
IJFwTIUNLYv0Ktiq+C631xg11LOwDgMA+J/C0l2vFvFRhQ6onaZn2RejUZhmCulZsIjFjcbf6DtV
jlR2Peyi4JPV5ZRZHET2j+OSmgCs3kIATTAe64Jq7m3DrsoLJjgnDFfYz1aDjmxcBIZQfZxzHOzp
NW624xKjcNfxYgR9LF9do+wE0Gg5Qx/10vsO5xBb6XyIFEHj1k6b8fKh3NU0s2sjOim8T0b2hjci
IrKpvQu4kJyDFRa4P28ImygLHJFT58zuy/ZLgT/ItDzVmu4d54xn88KVtJK0jrScW/wUZAC1o8uC
PczSUxcnnVxbsEjRbykAfdh14CrL4b0IokoMzgab3gzeKkpDZStlaY44ZB1kytFtLenNP1e47qiC
6KSoOORdEv/yjVXssn1Cs8ut3smiIhwkzE7tGIQD3U2Lprh6fMPrAfTl7gTOw8nwwRcFfKaFv2cd
CLiFjXOdVvOHhfsyyEahjchQnbAqy82UUkjBdsum58uHjMZUB4Q+Yn6itnBVEcCX8EnPOubarUcH
x9bIhADRJu5Ae8pIS5gqWpZWIvTwRo/8wL7KZjpKp4FFpSIEQ9Fdbj3RuyqgwdJFhLqxhPszmEqS
H+CpI3iY/fDISng2SCpodUh0FuXrxX3cbXbz/FQvPKMarMGi+YTWaXmIephhnamDvctUZwHVRAeU
H9oKfQFk36FEo8R9PLNo1ScxKGllkabS5n+YIPCG2hPq0FFLVxOC+p6wchFEtHxWyeppF63AgfXD
f+yuSwATmdkxn//fSJaNW/zqfBUQbUeS4oLaZiuVhsiwioeAqioeFHiBHeRNdqqV6xb4MDg+ppGL
b1x/bNr5LOnC+Zk0EEJWO2Tw0qCOgEuhOFoNqY6Oi8MZB18u4CRaTGtTPNkyLsxhRycUANZzY7kv
umnUyLy09iWO43I7zlvPtNMmoHfhNRUwjhlvXDhZpaGTH4KtKxSc6y0KVZe3iL2gRYZ9Z2lYJUj8
TdLM6gS4C9TkLR6gxbKFQyxcqZBLXqbdrgswHBE8+u31JzhGQpIkvpyYEK2EbB9ArwUjve5sQelQ
cdLKmqXnMYjQ9YI965lDwcRs5q0XoqUkDBYV59c37vw3aFh3vi7gKXZK8JOCrhDiKMd1YABwP629
+kkWn44ZPHo/7gy8miccXLEAffBByWTkgb/UdevNqtHboWeINUjj+gx5PWmHnaPlNXwOBFSO0rxS
xnSmfx4yw7R3JgVB7pDQB/Qxk+NLdzJj/swiuAirRW5bH14yTqN1RYlOe9KC9omYEDkpdMlX8L4b
TIr8EIva3LE6MGu3jyc6UriY7zhxMXyc09IIQwiU/acowoQFxKQUE4g43DWWzt2E4Qpx2joFCbb8
OC4h38BomEyXU/ZAi5+w4z9KvJ4388qydbGGhJwKgs2b3rqo9yBTMgNVouAdhVGAddyuVvapj8zl
rDW8G1PEPemPppKsFGwe4bBv3JmdMojS00IEav50fW23DTAD7Wa+L2qVP5OVhliOvzZp4I9IGnui
wEUCuLip968tvIGoZoOngs7wrAqRi9uPD9aLXOLTogboeRw1a459Zq68GQRp1LOCRtbM3JizFPRY
W7i2F4FJtv2AfqOsVdTMe+ZYefANc27EH5bk4LK75OGT91xwdsHu370qFs/RQgCf3DLx8jYF+bN7
/HbvJJ/zdb0x4fOD7qFu36+LwDkOYydfEyUGy34e639QDLf/M+AAQ43Lh5Ej8HKU/1D1Zkk0Fiq/
aN+bxKBUl+tbu+OKA7MzyP2QglmZrmtiBORB3fv3vNm7ciSnt3WWOhUHye/0YJcXFmFqqooBOIQm
vybqmSJDmzgLIWG/K1c9bijuzjVus/fdniorSEFdCJ+TsGzdk0bxDCwZ2KeIaiynkVAzAfnJ1gu8
Cu2Mk5zhI9V2udhm7t8jbRi6/aiudarAKAfme40ms/yqU/y362Ng6M5JHN9IiuSiE3AmhYAXACKu
Pfx0aQKhNogtwQ/ZPDOELY8f4VfRoKZrzrnq1hmKbqVPRdQSxUWQU+UW0AOCkxR3hl24JpdnvtWR
H1MzFqNkuqECjKyxv+paxeJFmqD8py3Yt7/EofBNSfPCh/4V3zXzLwSUsExx5LJbuXhX3f07EPs1
0a11F38A20K9M2/sqm7BTwcW06nu5bBmgbvWCtbCWNOQb1//j0ctH9LZ/mjR/lKPbldGvOyA8Obv
AAHahzvIujrGaW29PD8UKhrLh4x6eZO9aKKGHjeYM9ihyxGQ9lIaF0iKSbYLQH5+nV4Y/jPVL22w
AssdL+xHd5hJT0IogsxWiACw/gS0bZMAdwf4LXKWRtazi5t1QW2fuxEahkSDOAAK1L9OTrpjKVXT
QBJxF21Mdfx1hGdmpmgxcaGMmtNAU7MAOW8Xg/ouQiuxmpwjWH8TkFpS+o3JrrknCLdb8QVbu2+t
5FFVyoUT6GbWF3yY3w2CPj1yrGp2bvzhg8pUWa1gggvE9uecxkXB0cSe4yV2gb2+MWj4jDZGDbFq
okwjBBxM3CmOdobbR6m7OrDZ1O6b1q2AGj35r3gncHKl1YkOQIu0xmsX3hd12IVP2DvrvrUQnnp/
N/bto9B3b29TMfhu7bxslLEmC2ybo1Q9JaYCMFRwtfVsi6v3/Aq+jEIKlxNw76IdJO0Uf/+xRclv
+cKyJMRJ3OjKITVSKvy7T0E2o5ueSgDfLptEqyJyeZYR/0qxlY3+Da5MVCqLjCUOJ5G9AbJTu8Ie
k4Mu23ha7rSQD4zq73pUK4tfJKp5rzKCUrhVSjtyv4yq0dy4rUQelcD9JMKq91D02be2i+xN9S2l
8B4n7otPStOJL4st2gQtSTGHTENBp9P7i/2qOlWUiP+U31jlJ4nKfmRHbDMHxhAGI2AHXqeSaOBd
e430ycRynrh4cRTzEEpUYzZ6awhJPRATtv9MS3pDnqipKoDs5Egid1LFPMd5qVATzvG+LiyNs+Hr
qCZZGJeFMuwdoFPA3OjfYwmkX+TNhZoMNQQ+yVacSr+39PLKY+WaoOPmVUPjfsNkggCGrv0h2gsH
x2G1dtaDAtmuVUcGqDLdTLPKVy8I5c1yV3C+xZyyPTFKcqMCu9cVDxbmJruHrm4Hu+Keb8eEfr8e
Lzif/myKKg4Pj1WrU1wJFlghen7rll4XOGEncCDABj1whI8B5HCk4rufnimL58BfUEWxAmO11/hZ
HNwnQE1GM1iMag8NqUwpaLqergxZMSQMNoXxjGYDjzFRH3tqTuJ285SQyyBjvbSxBORwnf67m6EC
QnO1vzkPrK5M1kOagJwD0kx9zGqdx7Hr7erA3bZTWzw9/ETya5HtKzHAc5s1uLnLsa+9UdkwatPD
lZdJXo9lG0q98fNw+Gai8u6BjsgP9oiOM0+nhzm6174M47tHZ4DCfkopm6J79x4gA9xx2Ujsy0Jq
vj3c1IcF+LafIZPc8CnOvUJC026YwlUMhHeSG2sqQ50s+5g+/z/cR+JRg0CPV5t7NHA/T/aD+jA0
f+ghlDP+FtaxvV1mvKnRRziHsSLxDGW50yaFRY0AmhhUPkbthqvlsW8J+jVO3rZImUHNC2lqcLhf
aXW3XHKO9TahE3hQo4LbPqZeCO20cY0AqO2WaZy/QJCIsLKPSW6WVGBILSbr/FRLYYdEbrJ4ljk0
oaryG87TWO6psINQoVvCMbFHnb1W/whgP+RHYS2tDnmBPv7ZRUS22JuVeFxTbWDsCt4vw6NKUSjn
Ubi3a57VSKeapdBH3QuJIMfPl3Suwle3ivxOq6q9JRCWEf1sWLe+WvgiumYO5Lb9xNJvIk4TdlC3
cSssWTdqq0kqEBVJhkgiNK1QUwWxIRCMWL/6RqDrBWBMbm7dfl3hpKRL5uduB29srnEK+U9OsZcu
q/wB/MhhrM4uzol1B+fpvsDdf2IZiAs5zVauJLsHhq3ZuMowNGAb0BZdn+n9HatvB8mQJe7coQ+x
XQV54Cj8JFGuBVErPaRJaiAbvJj0LCPm7eyy2Kczg3Cwi4jI/gRB4NG54Zt/D4YrJwbk9cp96emz
brDRQH1crYdp0LpKZL9kVCHO7sS3+tWYdTEWg1TOKeV5KwRI1lDR0xNirELIp+lCycxoms2wUU2M
G/QuYYAge5snVs5AWZvqnNfv2QltvZWovxLu0IQOun02cVTFpgpXgRWGjSamgpH+RmoVjVRHKgld
X+nRcq8lWmKV54qHq6WRU2KpknXYtJRpmng95nUjLgQCesSXaOUjGOkTeupFgWcS/w4mGZSnxFj3
/9R2MUmxCVCPaBlWiIUKPkTpUklZMWOSp57uTCfA/EvNhCN4sxt/D7OQgQ5xlal2yPDHPc75Pn1U
wy0MbjgE88w8bXhj+0JQ69is4AYFFZa40U5uomhaAs4fwzAV2q7XjM3qP9yAo3O1mD38YttuKGrt
2fst2LF3h2CKpiN+b/u4LiZ+ZXU3OH3BT/joQ3kKQwrv59cWoTTWnqF2Cwe9P1Gs0kxpKEf4xiQB
D5pN7m+f+hg//D2WRLXY1ouXBBoRK3ElpFNocr3f/J+ykT1d4D+SRaoNxB9+43sXSttMdF+UbJd5
Ak73y69BGlqzvzDcDJU+b440vSQNei9zXqahlE+XUc48z/Joas25Bdhg5LJM/5DMdydZiC1O8Pj8
kXdd0nt2nulkBlLoq/3FCwJjnURMBQ6gRvUSWwmia8n8qbfieA6z3U6vy/6ZIjpJmzdswSfEYQTm
W9lWCBi1/lJ0sxnpJDRB0K6dPqSQKL671qYw+j3a4ojQhvWlXAQph43box1DXPVFacWJf5q9V47n
NQHV2FAVFd5TZahYn8n45FTn/47FpQ6NcHKBt/vVTNoSkl2ZkErLxW0lCf3MQL3feipdx348Uudz
aDcliv2HVB7if/SGzH2xnE9c5QhT0Fh3qlM4PXR79A4yoM3CPL8+WepXmyod3w+oeKqRsLYzfFJs
Q1dl28G3kqn9mK0ZgZEI3mDBeCVx6g7grlzwcilRQCBZaNKFvWQWwxPg9AI1gamE5FTWc3845+2v
S6BuPOes4bVHyrUFSJ4wBJttp8kMUdsFB8qoVv5ehOMvE+7dnkqYnxUKLtzpNaseB/br7MG6X+GS
FXXKWm8x50S4CKavwrVCWzjbAEw/N+I1t1H9KESybPpeqvS4Wyr8dRTogR+4F/xccyabZx5IABY5
Kq7G0A5AwerUvM4e+pACfhT9nlDW7HLtMDk5b+nPC/pZnD8iRFNQtRHZka6SBJjGNv+t5VpyXu1h
tYVzGMqgiDPxMj7BuWEQ0XncXDd0bu1aiMf4t34B9Zl8eNKMj++21PFgZsqlyWiDwxraFLTkFLWm
YI3+8xundsRSdA1jknr2LzSMJ9tydgLbT1w3Yo/EckyGlct4Bq/fHyyDxUuVh+0F3dMbHffGmlFB
Gg9vK49TDoiUyB+JEiDeD+5c1bNKwxEeW+FX8suQz15qJCBdTWgfoKMSXzVm8AESNqVgk/LVyKF8
ULSKymTuoLe3UuaFXBqG1tnG2qi6vU10erKNQZMxWyq3S98l+8sbQNqAGsZ3e/OOjmLK+blBZje2
80xv/kourHP2pNiPSqBFMqNQQvgKaf0Z0DBy9lqkKVH3wuXqil2y78VaRvVJ+H7JydH0H2/27dbE
KiyyuwQWcUb/0LrCrxpHv6Z2RHZ8P65MtteTVBPDBUm6J50vLNczzAYL6+8mXPPeGWp6eSPkjn8C
koa+xwJigpHuR5kHkNYF7HiVoyo+IhjJKoTaUcU3+oI5QKGatbIB/659DjXCQCRzR+yGAeK8y8vf
KAgmH5blkF5Pv3tmquvRXOITLM825dcBPZN8WJNtiJdwul6YOKMJeMEaLTEuWGlcLAkAa8qFU4D3
kNzG94GacbVtWmT0rwbvKsisMstY0WMQcSBGc03FgUha/00RLxEFmov0ejmWMj9nZp/dgfP7617z
oomOCe198VIGGfshEdXyPIuVpV+RHZXIJKJldTvAqpMnEW1jsLnrg6LPwx28Hn9hxiQtbTXe+hGI
w7NlWJ00xnNZg1ybq/rGevKU2kqGChSELn79ZmRoS6sLZ+dHI1ETvUNeI4Qa8gZg8pHeMLDbY9pR
FknhDH9/Ohi3thb5AsImwOVf+OXF40lP584s23+5hkyDknDKomts+Qo5wi9xlENvmQ49KePs1l+c
j8n7t+WE7RoqaQuv9x0SSO7UVRFpfk3/XE6lWfpBsuq+kUdWxF0EvhXQsZ1PDhAl5YURv6vWKOc3
WRhQjfv9LzttNoFu7Y6uAAxO4AyPpZrZGVtWSY9QoJjztKgfOLIhl3JXmlLNKDPvWTc90UyAchG8
NEK5JFpA5aGBL0aUPZIuxAbN5/AV95jX0xqeEPRHm/UpF3WYVIuIO9wx4hsgsnYicuDd1HlJCGTG
JC1EVBWbyMO/728KY6X0IqkQQDG0b7l/LXv6uSYAjwQ+CdGCKlsQpf8hb0ygDz6koh7TVCfcDuaq
wzr6Dlh6rryXqPoz9KIZ0WMBQT1UGI872BkQrBGi0w9EbQneuNpcqhncvmkvPk+v8+tSPc9PDXXO
AVzl+9yYT3T0XL8cX13L5Gvsi4aWHCYYfMMU2v4AtWxgGzUql66V+yAMM8UlVZRHkeIgNP/39lwf
G3u+Vu7GJlzJcr5e8tYvA0SjxeHyERH8bXTYN8jiDS0db58hWovmRxM/rO+PhvAUYTO431kA3U3N
2T64GoAMlhfo++Ov1RcXAqLLqvuhHa7/hAsh9oNpiiQZrxBroz6wwI7TCsluOj4LCDi1a0rqfL4b
KeT0hV43dRAV/B0thudHihZh7FywMoC0iYGFXMNnKuuq6X0x+1MHtNQNKf4soXcpGZelUrx2fykK
4QmeLJSQqgbcWibPvutEqJGCxFNsWszXWKnyov2rLzfmL+WmNWJXnY0ECMjbiEfXUKPS0+bj71ul
WMDF5oRHe5gsM4/oaWfThFJZpHWo2IZ3r/XPI88jGuR0XKn5RIonvgIrV6x84tOudqp1o9I6bHPa
a5ARwhs5fIj2zg525Mf4tQsdrf39DyG/UWi6sbPhP+BMTPzLaVIqzfP+lRH8wB/h/yrAHCRIREC/
K/K5VvMI8kgZfvuJriFUnAgPE2sdrtekqzyuaRSCW2qozThGDRaAoxH5rDL8Z8T/VZ/RrLHtTvmM
C4hO7Oq19h/0yyWXqnuSMV+tHSnu4/jZdIIXpGYff5BEbyJgXXsTqhtVm2HlEC1ret3UDRbTGxam
DBS3c/KvSoNHu7/fSjzRCDI0ag05B5uZlObJKmf5ePOziMbzvN/DsTOAfJN7gCj/P0UqZmhNdjqm
KLAx7V5NavtoMQGRvUD7wYAQK7bkl8EwWGQWw7sWPSkHlTu+n98KD85TDYVWS6BHzPr7g5R+dUmI
t8ckBaiaIzOQVHmkZgmcmamaM5QbDOZTbHmj1VrGk+0c5UNPVNJUs4ai6YWl4GRuRXrDA+3c0/jZ
A9SFu4sDMOAs0kOxEyFBXui8S2L1M4Q9HmMcps9saHdg9J2vA/gXebuZMaQtv4wVG1L2RRTOXm5E
i+x+fPKPt53V+a+RO5CxTapoAJL5RxuRQpL8Nx3Cse30+7+sVr4JJeevL3ag2aC2Ragln9rEbV5G
HCyfzkf8qNtyqo+kPdXnici6FBffUnqUXGTZEJ0Iwh/NLLMy+M4o/pX5iB+dcHDmyRo7WWRoAvYN
ho8Wgj1opEfCyPrlPPNqSJ1BiPkWGdSGNX5TN9X/EAV0FRTLjfqiOUxSG2xJkWhHmoPFWTbOT6K4
feYgCUVFhysn6t+/meL3pMtg/I7JvFl5oBeliW/xnwLbzAk1vSYwnO2fSl7kBydDbx5PHcbZALWv
cAwRU2cIhEvgw0xVF85aAOTAFL351xla7ou8lIBS6M0OyBwIu3ntByAOoBkDNPeOxkqOo7Wm1vAP
qbeIBvlUGfEiQFP529X/w9UbSP58pxTSrOX4+fxo649jkbDdetZQFIEi+MD/GH+JvBkAtBZ8Kk1Q
UPFiO4vxryE3fyL6ROh+YBxh4v5aDmh6SepUcJ9P+qQanndtJPUOIXl5JiEltcDirJTn+ASjT5lI
6MwQlKsza4EE/glY2S4n1J6I4seq+1uavl201evqMWfQ6fTnn0XFIqkgFf+NPJN0ZnI8IjuVdu08
lKcJLpKzDUadYPt/KK6IQXHBlIHqtADSrlE2leSHSyH6ONmxny7Q05Y/EZ4xtAOoFHrF+Sf347lQ
6QQgbcPOir9Wr3D8kePaSwkMQEHLcWLNK10u/FC70Obo1wBIC0WpT5cO5qwy6ZRxdB2q+gUQUWka
2+raUAd89jrrj2mVUNiyLQitcy9Xyr07NxvkaNXdDvZBcVMnmp/iEku8lTsEeji1Kx36UMAKY+RL
sAmNKV3AOSTBgf+2zlFbxAED8cFD9LuVzd86nAWGS3BT8DYWKYFU92rtB3CGc7VRYXnuUtFUOmLa
/DFRbfk/wA4OoPTeR7iBgS3wGAT8FX5RD2X111iR7EJcPBJkLWlhfibefaBAiQH5cEp2HpNdRcvz
kQrXwGYotEbNXHLTP3mVYHpTGZGgGE4OThoiZEYy+QfkNlqc46amWRGkLi3mOMFVX75xtz40tRa4
mkLQkv9X206ELZEDAY7HyfxIpOi6S1WMzX8YM8R3Nx0By3cppz/Oc35I+ETGLx7XJCIT2BtpBqfp
MD+gEAnEH2sXZjhYcIzJsy3EKy7TvYM264AbaPxnQzKGz/j7tbQHxwN/vP8fA1FCkbIAqVCnggMw
LJQ9tntA4OXnqLl/12uBUv/JUsVNNU3kGVH/4zE21BCnzXeQOAP1uJqoRUTH9ZgWqMcr5ZzzTAAT
Lx96iJu3MfPvlGufUXmPMlzOUg/SDtu6VjKA/U2LSUd4yTo1aoy4eZ9pNk1CkLlxT2+KR0iZYqJ9
UwTYm958/isiirMH9gcxsIoUdxlFNcdSAzvXSJy/ECnZoeZpV7ZibTx1GHOH2IzwZEI36EV/wYAX
LsZFcTCg478xGnsMPs+nu8SpnosZFr/MygHsfOfU4YDGSrYtpOx/gP+alJePl2vw0ejmeRwZg5t8
2QlVxn5+g2OGsIjpZmfsiRdnUUbzauh8GGNf0Jk95+GFZCXPY5NHAa0uY+ogy9+wiK/U1cER8IbE
cP2X0XKs2Jn4UjZeEheLpcvhcci9/RB0L8ZiZgonlD3ctUAYFD/zPzrySXf7/U2VP9361VTf7+AW
y1pgejgKOnHdaUJRVJ59qjjwkS94Y3DTy317FqVl8AOwhdpoMq+XyB00TKsqnkkO+3qzcHA5WY4d
yeN8H6EdBhDN2xEUGcPVrB6E2CDEG28zJ5opNglTdd9lWNH88Ie6yFnLmNXBeAOibSJQRS42R8fZ
VRkjlgXEuhD9NPODGMMDq+IxRsEJS8U5sUvKLOif90Up/dojDFfl4uE6yCPTQ+bhneDMN50OiJS8
PTDYsmtoBqIsJ4pqyhYjSnTUli8f9P5F4N/JTWp2zYTo56oPfRJrqjTp6HOU/xEtv7na92Rkfhgs
LVRZobtnMwWKRVsj6lU0ip+ledj+6cZZwQfpadY+Y3rl2hgXcvb7L6G2KF7DrYbIXDIgfNBz0I5F
mu93tCQFnowJXQwdVLP/+6H8M0gCRWN2e3gbIqD+5t59qX60kzjed7wsDEiB4H1HYMhbdnMuACPQ
wvQ1oJBRRfw8AAmxBS3efJvRUCALtKYzUQaLWB0BqtANSIk0vWlwz4CiskmpgeD3vXGvOy6iFLU7
cbk8mwNopo52IE8OZvlnqZiqRfatb7wo+sp389vfOecl7y4waBOLsVfPhGv6NxJT9xGsvs2qrFqw
fjlumNrv5A78DXh2vKxYxvfFcn5LftDX0X7muVOWAiXLCWKiqMEbXPltzrjx4ooqF3NminmmGkv0
jSLMXnbvVAxbH5k/agEGjqZgq9mKYCow9crXTCBz4CLjIXqhrfXVCBcpIEY9u9M3kAMVLTU6ZBz7
NxotYKuZqZdlzPmptBWz5VRyXGU3ZI1l5qPAdA9KkZeb9aMq/MAWd/DeMn4yvv6FnaiXsCavsklK
Xpfcd+k6HhrRfrP6QLnX7rT3QnTiFH1braN0UkQnuO3Aq8R5baHmzLrElO9mSsby1n3oHbbcrSf7
R9GH1/F0YWceUUsDa5F/3L3WM9Fei2K4iI4/GR3Ue5tzu4m1T9fL2px54T78JX4JNbJqownutjhK
DC/1Fll9RQBhyeeEX1Iv/TRfSmkIW4gLgRZXV29l4Rr0Qabt0bBk/UsuZGu9j1yHrhJSFfSvujJz
lSJYQzB3BfROZOds/LuZZ8C45Hn07f2X1rgxK13r0XYmwDH3hnZUMxncwKmyRXeMYOTKf6MInVar
U9z7fAq4/QZLZd8R/jjbnvo2k4gaYSVmqp6Y1iBJqjjRC+8dQ7IkTWfG36tNQbHC2qubsZWXGMMm
f0OnutZ/WoPhyyBmxnRn9IDfrw7DJNOMOpahWUwynYWttVZUYIjjovHNl09PjAzwdAM6gDiXtwJH
yxCUrG4TcxFnx+0x9NlXjaEU22FjOrQQF56Kpa1oMqX9F/qgdi9LUUjS9+JR3IGXtmzOOtbvxBcr
TtDBCwHJFsWtn+I00JGk8QSgA9mtEMwW7W6SvJH/cXHjEo4RXu36goqExdwZX02wjXRJJS029iU7
LoQaIOM51FQlxl0AXwytkGPQ9Xrqo3iHYFtaiSZikVNriC47m9agtRxUUzjFa8tbTR7JUKBZW7RG
lUfx4+f1iQuiDc6XJdsBE0+b5TYEH/w99kvAonMY5RT0SKmYZrX0hr4tZ6wMbAPARSfVS5bmIJ3L
P8rCDshCjo9Al3YhWorZ8GRH9mv4LkzjLeyx0BAaszhFrq5/yKllDIgvvcKtYBG5uJ4v4E3ovL2C
Gtd6E6YdS10Pl06SRv3Mg7rCJ500/sz+iocRnjWBtqQ2wr+dP5iRQR771BGGXlt0UDQ9SqE+6tAa
FctFne+OnsTv09lHYG2E72SQGyWhGlr3jiSLJaar8GaavR4Sqg4WDLJ5ZnIjslJwRn+SrR3sOwOF
f9AQ8NlHeVTCIGYzsBNScSJ8T2dteyIn/1fvFgjoEtdlOlXG4p+HyEOdVJdGTKhl9aeQkYoNxCre
Z8a4j3ti4DjdFU7Gx7sOH4cPZadNk9UkppXszUbaAU/F06FK4d+Gk9M36bj26TAC2yBU+Xx+1kgJ
67w/d6l87BsbevDQ+E+bf2rIHdrGTyn7hMCpJ6w0ZqDbbTwHabUOkVBljdT704jIhtCq9g0bJL+9
VqdwdD7oOsngz/0ktUj/g2VF4FnsKzuLmeGyFjkq162MCRO6oAmSm4hgwgdVdiHPlnfb0VxOxen6
2398KjJACqQL62Gu6qSgbk9sCQHJprx5b+/v+6qhi8k149SDm631gpzNf18AxThe5zNbpAdLyVBZ
PQnyGSn+/ZRftn5Y/duRZMCcAkUiO+GhKixRCBQRcfM2CbpQgWxPf4xjcUyFPQE8YS5Gg10qMf8O
mVNcAWOPcJ+rwpMln+3FqCy8wzrgvkeUOsIKhBft2hyaCdajqWqRho7FCfC+taIBkba6k7L0MDc3
MPNCLCUQCcUD9lFFaGnGOa7bNGrnk76GACok0L4Z/MrBYaZ16v64HpJWsfyHBXYdcWHWlkj6W/Ms
iHcgC7uNDN3vA+pqTU7t+EPe5NZLxtdu017Qu+ECpwRqgD+u3pf4QLyOQR95eDRVIFCRZdDJ/ewj
DNPbCd1gljtC5qA/fNWOt8iodnmnXrgxNHDdcjdlSd78k/BY9wZCa/nQooPeVAesVzCBf15QnTaQ
mi8s6ENTroCor921jfcjxjwspSrgNeb8t0w32CgDyUQSdXX3s2G9P+yxchJja2rOGK+fi7KPR+Is
0jjaaBl9eLWZOIEgnOfVa2RSy0JiixIT6NH78OJD7UzlDmHktRA6Y7N4e9s3UGV+gl5lLu8DPHzT
2/5wy/E2mjSoAC8p+kg5Z5FSfqauMwsffq92J5ES9AR7xUPROBl1e5V1fWpq0oMECFDkNBkwVbcQ
M5JPfltpHbQgdaC/H3SWmXrRAiV6TXq0wgvKWb1MNrOLvRv9F1mXiqSl0yOHW845F91d//uOFl1M
q+rnm6yjUk5kTTPYlPGfqMM7PfwdjmmxVT0mEzTZLaMj86y3BagDxSPXNrsD2187AqmhnbeSpceA
d5sWZ9z1RTaq5z/XYUGtbDRe9quvt3giTIuLk++pzhCKSltZiEe0LwYEK+Rus13WYbI+Ioo8OfHw
QI1GJxbM6EPV3yS1BXYoW11Y8zMTqgjBoVqRPtfbjHjnPZgAj+xx3Z+hlCuHJntSs9ybWBdO2oN6
VBBV4tGeS+OYpQUJT5hNuKiMnoDNbGP+Wn4r78Vc/lhMh1Jh8BHgGnpaeKyqZgJFUG22z3NG2wkI
Prz7qT//RObSJkOUCj19zz+fQbD5mfKaK2FevwDwsZnlCQ3+zMLM5naqyCmQFsS8GtruA/X4KjFY
esWac/5GrCS6nTgGY4K3pWzn2vGaV9w8JuZS4jZIV5eHN8zG8H2JhfNdAq2AnevFcAgWg8Y6Y9x5
n+Mr5CviTYRR/4/2KqMOXHF8RTerjmdon5IIm2jAFefmgiXK6m96PRlHri/fl63aXh1FjzusdRIh
wfYyoCPIkeVXnquxqw9bLz50Hxl4l7pb9Qc0W5wlvWlHXoRt452gJAj9teVzdt5EkHISBZI/jJA5
8pqLidV/Nv2aS7LRRNX/+lXIbzI5yjs+O01omovyLZ4BA9mh8Ovns0DgxhD6kNk7mxRVFdpoAGD2
k4fv/wJyk/tUTAziAE01KSkfrDMioJkFjBB7FgZW8jMTV8b7UWtOCn6atF9czOpwMG4kGdmsyRas
Na5bU/kjCtCk/lCjufkLsuQfZA5TCdGDMjXLdXxip9CY8jqJVXW1y4UAA/0KS59GV11x+8oRRGd/
LFV7vpxwrhgyHbExQmrZEZ67VmOC/mnAmhQ3HFRC+DneEAMUOe8nRs+hP9RowDq9TZ8t/1vqIbCd
RqD5aSxhuPG33bTEwp1jRsJAuUKpL8UzMv3K972NsQ1vCudmIe+nPIrODV+DAVwEmGsppmHNEOSw
6+OIQbTwNn1l0euIyLS6CeQOC7jAnAz9vxoUd54b/p7IKqja/M2QHsDtZU9StalEltaXKR0R0Pud
H97eNRCmUu52sR9XbDmO1j5hmirZNypRFM5Yn7fmlDj6zEfp5l1h78FzLN4h9Y9DRXMgQ4r8+fOv
WfZGpm3vgkzLuD7fxqE4xRg089izg1WlraLTnc2PqSoR3P1r5wUU6y08yMDgSiLbmYl9QIKYXyzK
YbEAKz9fzOwcyYRD1SLatNLhqhCcecJUvNmKhEqb01gzW9JYQ5iFwz7qJXbOelCZtHtQMpWUH3kj
qlmnyQJ3SwDwUAV6Ky8agO6X+IWZyQc8RZ/L+JnwhyB6d0nFIrCWuU3RdQrfJm6BuLP1B7OmIA2u
VEVQB0Ko0r1UV4KQ4hlHku/BCRkEWzYpuQPsysvzGK6YvpYSBeiF7FTT3dWiF2y/ZicRc1clIZsf
nCQlq2z+XTezv0Sq1aQ2llG9IuaSG238vE1uLhl7o2p+CMjPvqF2I1A6kteKXrs4I9BgMfd0KJNd
wwSrhA6wlDESWVKYO6my9Sq5l+fEx9Uze3ewtJyjHFs9fifcR3jyGIkAbAAP5nvMgGDeVRbWs3PI
53BOovJouxW6vb/CdKpjJbV0A+0Dc3aDGwF9Yk0iotdLMpL10ZvT/uN6xzvrHSsCirZFE47oVlYJ
Z+bMB2YS/PZVG5x4braJZEiQoQSJ+rjmnS4MRxOQ/Cv8Gi45shzelt1TgXAHjeWVhmMEJCK6nN8b
REPkObGZU+va8mbhNIWmBu4g/+tVTtH85lPtqUrumwSFBph+i+FzfasLWaCtb+bPUxGRJQIJiq4t
df64BOIKmItrlkCscuo5X8fpWYeuUa9XWO/T+8lhZS/rfxyZeqLBcQvh7+E9Lwdbzuyn0UxF56Ag
2uFgDeTSijYnM+8v+qJUxiCFH0x+5T+0SrgIK0pCDZE9fkj50eBIL1DDR+nAURuw2FvaFEzTZ2aW
whjmHxPiXPDcVKlo8beFjEOMOqTzAQcyoQXtvyqRGBx47mFQbxDAR+oVDiN+2v1JAaHkLOIKkjXm
VAzidW5a1Pi0u2Te3qHE19Pt1QHDcN3v1jPMV7CXVwH1rs++WlM9q0FTeVUVgPZe7Vybo/t8sWBo
sEiovBAPFUtQSDQ6LqmqKSn2tnWF8/sDdjAz5vp3vgmUWcguN51lzYL33yEVixv6BIjZdxkHbUzU
Uv9+IhAFQ3muGS9r/VMSwG2+7X/tnHL7f4Ia7XJlA2L07PVPe3jxvi7GkPJ7PuQosqD6FltxM4c8
oyx8wsNcFOfAJIzHv2EiX+590w3vyRmL8LQ8ACY6+mlskEWFMgqN6eqtxxmjFX926OP9EhqqJXe4
S2CuGoAdMccqH/ytfdlCjBzjG1O8br83J0a58UgN4G/Qz4+I8+jx4XhyIP0TPGMLf4hk94+/LgsB
T4BeyHR+v7pWYVHtd1pB9BVJQqxguThce4MVwcpZXiUT3Jjmwbo4tdBcYN9Kh+uwMTVryKBRQ+Zl
uuXNKFw2i4htJ8kSXpj/bElXafAc+rUQgUdpQhe0mJugepSj8iEEeVF8F0y4e3P20i4Z2HgX4uqs
uuwR5Oa5biZVvPPZtl+z6AHmt+GNdETWjQUym0w7Lo73p9RZ6FPYJ2OfAm8pd5BKcvKZyzXKbGdD
Gm5pfgE/uyiQWd5S/qjm0q6wvCVqD0YkyAyBErDFge5gVArfb1cghZBFPCaoRP3z7s5R9ElElx3h
vol2ZEalvnbY3fSbnuG/jyZ0NI2gWIesV/rR25G3Lv7z0NFUn54GV2Zzxab09AMj05lAnZIX4LC3
0wgcJhQCK5yLFV0i0JZfHQlf+EHYn1/oygkDxR/1ZgD3Aj+bbqGFQI64av5kYb3Gm8OyhOsVM/MM
kBgMC/cKOqKcWov5BH2+6hI7zQ9PJyi43sSviuHSBbKtrrfHFgYEKJcAYOueVC3OwopyH9a3T5My
OgPPwasFh3rzDuUPgkSyjXxVP/+E0yvp1q4+110/CEFXn8OigriWeVNkAajpIhrNnrmNuKx8ihAq
0RdCNAVJ5CsHnIIxAmoxOq956ceLHLNjXA+WG9THZHVRdGC6QF3IJhQe5o/S2IQbJNZm1fkl7/IJ
8TMhcteU64tosvH3k8H67cjjR/kabeMj3i4scg6P98YiQV4osDcmYt3X+PkRObP4hKYANnNfw3Xw
CUQvcvtndnGZ9Odeu+KD55bv+VAOs7+QA4fjkTFNtaGdopBd3VSU3wueGiAfSX4Nj0J9yLDXExZx
QdnxkycHHbe/qkzBhjxQJ40EjhatJTS1cxOGVrbxbinzC2IZakQO42VZjEAvtRCWVZBXu9P7kxMk
tQdPojmpJVo0WPlNGbzCf4PXlZLBUQrjIy0adcQ7l7TtuA+gRBQ1UidDx0bVFxL2QRMh2bMwMyAU
/Cm1Cef5AxSWcfWJ3jds1IYdoISd7ynWdjwL77DoAiNrXj0DXE1o0sYEFPb/kdgabEfsRuQcYwsI
uqeUyFpMhr+0SBXQNELkudNqkqiQ5SzTIEM5ztergcVyFSROS9awXIx7GpUgPZak7gNgl3HyJ2R0
Q0LiEbij4wOFJJRQddTJedxDNfRjz0Nu3/TVzGYLd1jlluHLrv4yupw9lk3IGHkJ7P7qw3/cu0yM
ybraVNzt/r9GZ4BgYXuMRD6HnC+3ngN2og0ITF5qXXuEoru0XI1xTASlHuLuF/QXhUPPmFw3odBt
PvxfHtER+OqyrHEFePinELVNRPqOm85nS2U8aNWd32aKXVR30iwbVt64EyYwPXrzGudhnxnIXKp1
mWoTu/hrkdWVTmwkwDSpiMPZ1uWDw5QRIf+5CrziNfH7B3TBf4UjtHBVGvPPOg5G5UoA60mAAocA
GGPowc/lbmxTcgzrqF33CLBHxHON2H6X3WkdiLcKi1VZtBLv8KXPK79Q/xS1DYdtL9E5ThxepRjZ
U+/bbAnQvQ38j8OSEgsFS47mOdaPbX4MP4t31isq5/ThuEoHJBAab7rPVRkTp32Y2lxySQdqUzMA
SYQdkot1meu0pnJdBou80MqYbcivvtUoD4OcqfLqPN1F/RvXNaNMRySZGPzUVicvSP9iQJzbrSux
ALYgKkRfumgjAqCFYCtdo+GKgM58v7STs8xWvJb2XL8aDy+8y49LedSgSMpJjg6pNNc/8GzzS6J1
pbCYkHF3dBdqVFk67uXq+PmKOTetazjZCBpL3xU39o72yWBTd/Q1NIFWdDOaqPfkSMjPs+9IHMY0
lwIZx0m9m9b6uf236AaQJfFTYDah9lgUsPDoeLGyEzBIx4ZX/WOeT0YsOK5otg42Of+fcZ5Hlddj
Cj+RUZJMUSZX9ZyeYeCs66xjQ10abO3HezYLAtkag7MT22ZCHjDuSKcfGHLhHgKZ3o+ovgPl3v3j
NY+2Au/vO3yBDS2miSb1cpC3PnvutCj9FUimebCevs/qCyPMlJSMGSKFvE2sIdvmVHifpAnJw6pS
zXXVKDadgDPNeKkKK3DFeyghdrmoU/qSihQqLDvYIrCXiIK0luIqwsvs+dauyXttZWwh7d6lXmxf
d35oBSOmhZx22rrsHU6nP/hjVXS+MMocp2ZMkVk6enF6WLhK57UoSXCyQGzK+qaerJn+7wnpdkvZ
OcmstfTf5B/lOq0W8CbkEX96W+5r3J38+zLRykz4HRruMORPFpzZKmt0vCrG8c2Npd64ADMb8RM6
WP9pQKWdoKLajuyeHXk4LVgfFvQFrxPq6fDoxWab99C2/xu577q06ttyG43IyLniweJnX27YXZjY
2clZRSI+ZTrqKtryamEQwWSphV/KrMDL8F4s5miuN02FOd6f7nU448LIKo7rSH9/vJCUofi8EM1M
QmbRwD7oypUMPG3axbwb+G+Ah6OHrfceZ17JyHBFrQF+EyLW7N+Lwvr9AJx57H1Ow9imrGrxchZD
dWBcCJOBzzvjtVLwuaheSKatYC2SqBzvPVE8fNWTLX/ronke5yXdWwb9XvX50Hz56RyjwCjY48L/
yVh0XYy8kJ7SQ3gSIGknDAYBSmGWW4m351VRBJuu+I59aDqfNtmVlx9VAfrdB89qx7uLKRUBRduV
GHiOG+Fl97EcZ2jAZMLyLF0wb9u264og3TWY1KURzHXQT+Z28TDP+9Ko0jtWF+fPZD00pHWcCrge
nVVvQATaWeCwx6H6GbXbByok1ZyjSLbzMwwGgszlZhxAcAOj2bNghgi2aFRV3UlLYH3+xk/Z0hsE
nKMI2DunpdZfaCREJSRa31woPiJqUYcfXhu0wP0MKFsTZic4yoVshD2uQUIAwmQ4kGsgji9/JR4w
B6YRLvSptOktcTlzgedw8rGELSG2DgqBQDd9BFUVleLAwlGFbesjmeVbZX4+BEAcW6OxH7Htep6a
oZU4J5pcC88IGvEjc/hmH9DWo7aneOHi6lbLvKVH4MOGaMTXEHdRACnEodYKpiBP7SogG5hOBwF2
2qX25EYTvMMnIhcmsLBilYQYILPXOWmvwgVOGpf65/Ti0q26baFzIjXqqtg9yVF86EhWCrmZiZQy
QEDCMZZKA0lvQ+ROD1YeBzv/YnW9N6EBKBqaxyE4S2IM8JsMVFnxD/VGed1smahj99hbbzwqt1TZ
DMuNB1yja2cSkklG6BYbFOx9W/GKWkp1NZQSj+C9ZmMTdyzQ8AfNC6btZatXl3/Kw44xGjwYXqk4
BPWNIYecvPc4iTE6EknXiYeY6oiiZPvAS2WVZczTY4tmQqNx2EQbdg6gOf1RBzZVUQUtVesrlYVv
pBuuRHWbcTfvHoVsrABrz1iWrzQji1x/FFLxeOvlDOjcbkDtn0kB8gs/b/x7gqWBwVzV7JqBBjuq
xQbL8TUO1As/WHuu2DYFsktdrpNKSnTU3jRiGTYE8A2z8Xgrh1RBelxwwVMZGTso/cKVdR7D8M3V
SqX/lembbnmvnOlc0hY2TgcFunVpjLQiC/1r3VudwHpayB8zObl7Ut6vi76SK9eWNDs577RxzzPi
raWHZF8xVhBajkkU6fgM4xw7bWAVHEio0j8L+I1lSjU5hSN9dX8mTTbnxJnp9nnjfr4j3NZXzvXf
h5tAl+7iGcV8D4IpcU5Lv9B8vdcBR5BV6/w8RNQ4uxGkboxGETjO964KLLDhnhFQbl1xQMpRFvU/
u5Ss9OtL8d+2HpfhUfCISuv6M8JRfLVvpQ5DgsMviGw8L0LN5qcEoanHsPdTu0GqhjgjToFRfRVR
zhyzAmgezWjGX+abnAqOscvQ9ss4zcHLjFgkvtlDRcuRqsXVezvnvX57bbTzEqHz4p7/zBOP+uQ0
qSPayoGhXC6b0yewdnhwzyuD0yosj0Abdp0YjCoM/yP06wdLd4IZbkLOdZSUuiv8cqeTXLVIuaOz
gZHKX4XOExEhl/YQCskQYWv73F2UScE58gw1Qe0tE5g06ZInCbRx7KWC4dX6m1VxD7mfg2hUG918
AGGkVerd9Hr2XG0yD2itZaUgqv+WY1KwejZTrot1u2wi65O1/jPKxrco32K8A2RAFo7qBHuz6cNc
SmRanEQKiYtYPIflP7E+7ckpBfPKlzUbiL2sIZgNaY966+0wwbFUe4V9soxNHan87+a9rwVFygJf
gDLP+AZaVh/Q11BD+nto91IsQ4kGnFZwH2JvrLLqDdTKEbx5zFT1SDd//9ehOU6uTTfbmvYolVHo
7bNCzcOBzXtW0ux500rZQSio8bNmWIV9VH/R3jPK0LEvekozGrIw24Btve1GoJNizmXR7yEDd03A
VfCH4kLZwJAJ3ILOXsIvMv/oysOrb/Jc+zBPlHEBby1D6uf+YBvcLyuRTjJspWSBeHLZ6XuTFUnV
DpnErEgoTO1g10sW3aLdRWdvqzoOHtbTCWck20dhG+bFanBJOHbfQke2FV8k9GRs0uhwoAVX/hrk
oHJ5mvObtnTGYj/64HCuVjnH/O2iZrTkbZfDdXynoLMjKL+6vuNJyqtMLoFNu9OFwMgEH1hDH30p
MrSRYw0yT87mVAxAlFTWJ6xOMMWDv6VejinKUv49fKNI7O4JCzJYGQTf4805NR2LWmcgzpa8Fpo/
U8cYcIbf2xWVKClF5fd24coqQT278wEqzCvm+6zr6Ffg37Y84srKmVKMHS69oIlNtaGUELbH6pV4
EGVdJ99o/B05a1WKUuzXUiZovqeiXPftOoY8+RSb9dZFnJDFAsyTtktKzs+pFzPaO+gwRekJoHBj
jIM78fLXZvILfxXe2DG1PnQjakTwXxsDl1zr3+bXb1Xa82UUtwN6Sqfe6opxlbL90HN/fCCAzvyL
EzQkLQ15ig+MfAMPOVQVivVGTkZC9fnI3WOIUGR04VbNaiaQ7fSvRlNz6HgpHIyPQ9Er3JOSVaZu
3m0YpAB4nl8iUBH9OlGNVUQa8VpVcfafZb5lWplwk1ZHx27tHzd1u1KzZHlsXQo9kc3wcixC5k/B
wa70473yNMNRuYtUcIgqZC2zDlkGP2rxmm8pNDqn3ZTiMVG+CLZq9S57AeF4ifc+Yvex4npWJx3E
bTYtCoqv/N7ca/hOC0klnuavbngLDe4G9yTtrIlonS69KwWe+8rOe8rEkHx3dBOGCTeeF8BNUNLz
IgZdrmkiMNj2duiv34a2/jaweGbQNPYv61YpsQ/KLrMR1O1dDZ0TL2cuyGpWV986ZwmUjtlcSUGY
XWYSXOiNYcX403O4bphkGx5trVAY/rrglByDf1GD7PhDTyN/iKkpzmXP20ydYpIqvDi3WURxX8bJ
ODypyY9pznCXmFCtykPTZfKL/krkiWIDpLlPZke8Wlfd/hKX1UEVEtsNsGS1+VwMqy70+LYZfHw3
XQZuV17DnAIAQ23JzcVeaf8wOdaVpjN9+2UA3fjT6XDn6LV6XcHTKSRYMnilhLWg4BS5WBfkeUxM
ExnCML1zNwK85wgaATuxedugA0CnemfTBgwWKVpSkvRoy1zBVnxl9Km7uPwbkPihbLVPZL9RrTC5
//g6fclP6ixGweAzzKIE8rQ4dpkj40DbOhrZnf4TpqKq59r6i+7B5eiPlRRXq5twGi+m+QYSzeiL
hjixVEFvvI9zOVLTMVEmDL1BCWt8ukV40v7MC8+4MDfOV42z1eYVwvg126asO0T3dzm0KwZL/9j+
KUYtxZGlj8eqHG5Q+IP6SU40pg+9na7aoRHmBRhrtDHXl6I4wZBSi0nvsQ47XtyyOse9wj1p1psK
7YBS2IoND/Mn/gAJXw7hPoUqhCGLw2XiEVWHg5umYR/OhLGsyeovHCKEuA4H4LIIvYnQXwh9TPIa
dHkEtq3aLjDEqZWwXaP/S4fFMXQj48EATzEVXkJ5ckCu9KWqN2Ob9qLuJhJ82HWTUitVpgREWCJr
I8lBNGQpg5SQbBDfdzB/a53DSXFu6DkjOQACQodLEnOlgraPiiekWRoX2yr7lGrGVq44OcnwLhCO
hvtsXeFYjwIXcPcRA09IuA7ymfP67Y16z4Uh9Lnvc7S+Piq3cyjAR7mHx9jvZwlrJJ9zs30i43tZ
LfrA8zNQLVP/dXKacFvuQqFCRLSNu2UEnEaqVKbqd6f/SLCcaNoHc/b8a9TBNRAugRS9whAIHdhz
tJNCMBFB0XwpbhT69VeJub+quos9gNFREwcpa0TZy1DKFFLK11+qfmMU2wlsXJLK+Z2AeJpYRsJi
0JpyWQ8WiKJWS4qJwiIbiSdBkAEg1Rurp0sqFE2wP8IFqj2cESNlxh8d8stNpOVt48ZFwanwKje3
PJLvOQcrbQp/aqxmNvAhyW4vZ7lRqAdjndyg0T7CIfWPRdXjq2J5ZTcpOAI7XHGQWRZj/PJ7Q/Se
QaVjmd9ade0nKLO39nDPCb97kbCU7gIVL6G+D4uhNEFJngDcPJOlo4Pvf5oJtGCXig9xRLILi8z/
tWX9V6ZYOFtkOe9A0gJsA8JBAZZJk3NajrcOMDIBa1j/ycHxdRu3VKJwGqDJM2RdXCooPS50fmxL
DbjAipmo/ihqUepDlmmwWjb8hLJlPKPORmzqOJTe+VZ5fsEPSkUtUKohe3PzgInOjoMN1oG7seGY
QofzCfH3dwtwGu7XbTSG2YfOBajSYkwkkb4vkPVi70QR07XZpg+WrBK6ad8n1FS9YQymbLDBt8Ta
Mb08OLKsoDbidNy/UqsxXBJPL2V7syeE/pAQA6vZ2Afno39FqiIj5KPPRqj5v8w3KcXYJYk+OUX8
qQWawJyejefAGV9+qXk5/XWV2DSI5s/U5A+FbdFcM+56/V5yfTIu85pLRnHJUsUeUPdzQbol8aJZ
/6QsfIH8Zn0szPaTAVXhTS6gN3nPEsz/2XoBVREpC2radey8uPFQFU4Awt/BZkHoXN6+Sdo3i4BD
qbJvSBBxMmiRghUCf076ujnCze4NMGXX7LDeMTyVg2Y8nt3s3Ro2WIUp4BIWWjaEVv1cKm2GgCxs
qm+74sJG6Tt4j0AZAbXRukVQW4MQe9L+ogMXO6lyzSO+Z6Xhs52hO8/OOSsi2eD6EPqIWtvcaulv
901Ot3r3tGF0maV+Nh5jiBFPTJTDK+qd4s0cu+KNUNw2pyWj97AM3LsClRe47vPLyvd+/2VoG4hn
zpwd7zKjkTvUyxrGR2WsmtZjRwHaJ9CiqOex3Drp4nP37I9xWfJ66RcIunb/fx3qwMM3MUo35T3C
/wpet8eN0u3AKJD1nMIidjCfaf2Wy8CpFhrKvMwqMQfnIZ24Gvi9CBa0RT5X2K2+Gj7BtjnpAN4E
KS9I5psFKt6VA4Xg2AqX5HvT3zGrCz2a/dOApTeaTwdkrpa4VUYLAOMaaq+p5T8KU4YymYXyEl9F
JIdErSt0wXefZo9EdvHHU2MNblCKISB23OCvcAtafGKEvMnRCCQri4RCS2UkKMo5jExGVyVY2qws
vU8L8sqFpssHkVPJvJ6s/YIyHPtTrYktt4R/vaG5qXOEF4j1bZY9KV8cONZQ5LdOW/bGe+G7T1nP
gYiCGVWBpzlAIMCJ2f/+huNGS71X5VzNE3hMgwousBgY7hu0VuyRyWB6xqM7LWCgnSxt5PkVWYwV
gWNNPQcLYbY0uzXF4ui7hIa3KqdKl/EM13AB+NoD+DoDptfu4874zg6J89V1BZugzhu5XLvWApJ6
M3BoJq3E+AJOyofjg+h3GH1tK7+MH6jt86a2j7NZgI9CbOQzPMma1vD9ZwbVqQk7r8Zie13qrg5O
XFHDR9cgHJ0GlHqxCDAeV41fdnZu/EmsN0LdsMS6DYf37uWL0/xVvToAxoqEp+u76vZYvQaqgVS+
YmsqnKPYAY8KCg84nz/i2UsMCmPBD2PdkDGxf7GGTFKi7WorF9YRLbeedpUdLP9WuqxCOUGUZDH0
eom4hGkJQQaAbz8o0Zpww3Ziq0K0JfJOFnH1LM2bhi/zUnt9YL5rZ6xtLEeON26EZ0d6aZ56ooEQ
mIlpBCwipblt3tkdmtQ/y4DD9ACKjs6J68Jfw9M8vBgDvtFf4nedV7IHJdnT5Fbe6kxIwmaav1Uv
i7iEP/whUC/M9Ac12dBl05XOLozVrQZFk+AapX3IRAkzxxfSINECXShmFRbXreFMtQeZSIOPOCGb
tcOR4PtSvLQJ58tFP/KnT49tub6Peg29+TpwQUdPnvVdrZ3PHKmUQQK/1gd60kOa+t1TkSfWqbhQ
mcKuQV9IE0LHQONs7yCWyNBL8xrUKvPgGTD0RiRoScclRE67f4o04ohXFqZqvwQVE2zXqf9ni1LZ
QOfxmZsm/aNws2/RgOVAy4JYUwV+Wje4J/GIpTYp1/SQFibOShjp5j0VdiQ4R9wvD/Om/EWVp2jw
GDhAJr7xYCItWajXsmC6vi9L+wM1vQcJO2MOYNJQocjNRVfGaLA8U0HJmcC5a5P6HNDv7qfrbQmh
tYIXWVBVdUUdUyjJ00jT3l5dcrHHBIbFTfRfbt/HlMI0a8NZ7dKKfS7sAlQrn/+cORWKg1oqugc8
HgcXDEBKiEag7hGzpqXWdkI+kNy4W9TO8BIbj9Dy/rEuq6t7AJqd5rw4jOw7RmaR+AV6c+tqykpd
o/TevkqWszmAnwzhNXZddVOUt44r7d5nPIsX/IGBJzicgrCx20gpdFfypV1uDjykuLtPttNMvmUb
X3EmKklYP50UM7KTN0w7DqcfZQUKBsynrWLYeH0bvVjAgoiPOlYV5UFewMwoIJHct3NO+hkG4TyM
pGE1azRj4NsRL+0FOXpDfJ0YSRNQ5SzvyfZuVsnled4Bo5gBh6cBmw+AcHvEr/om3ottuxDjEOpJ
LrvHkK6ZXQmk6vAk3tbURnVtMUPhxBREuhTkjIhfq5SiPKFtOObkoKvfDZDSH/2iJbZvZNCAUkmA
jv7wZXwxKkev6a0a04N0N81SVOhgeqIy6OamWODdKHXR0JoudNInxDb7KrhO/uBohEfcakDp4ocr
6NIuvltsH1u7/fD1rGqDfTQF6+dTZOSCWaWM2v3xrC3eI702fQVllcvQ1EnYeBDg7R9xypz4hQhT
1eshPz9St/4pHNGcXQQIXmNMhKVpAUxww9HffnbkqR+kgrwql4Qya20VGRYegOgKXHOptUMDS+C4
TPBlySdPyk+7dzYbiIsO+fYeTtGDGNOBOUH+M/AIxlSwFdktT7P2/4ClsIGGZUaEgruDuhqWnyxc
H830IxQ+RbfsYb5KGVBEFn+cO1E7cssY8MOQOS1qFVR3Gdpcqh6RHi9wgXIW61EQKQrFKcAsuYrY
6+FKvU9zTNIzN463SxRqlNVJaQhPPhC8HlsR1dYX7PJ+EO+sinMrqusx0yt53TB+bF4Qw2Kiayx8
OR9iXi6OLsnVUeRMTH+eYs6IQFDFrh1Eg75GASfPbtkgJnjua3YpHS6AG2OSOI1RC9vYlWcMCu1e
ys5CGuoCwaoWSVALS81j+44tzfo03vwhZd61Tm1aJWGCwxH90eK8XHZBHR1QLVHE7GqZ/Xw/K3/S
VmUD5p/SlzvseQozD7z5OdKrelocgda6gCbfdFq3FL+s/fMmKLWrdhiqW03dE2WnSRyA6L/KV8lk
8qPkdSZLfjx8SkZFolam7boCZ8DWlvOHkEocsiGrI3kXRT1eAC9fmQg1l0DZ0LdopkMrAB+hOEjK
0lSY+fuhS5LNL4UnGGi2jQSRTLqY2PaIXfpy+V9uHUWvidGwHJJXVRt/K2X21BgH0COJcHSCouTx
2TgjKOBBOCVaMoGDcT7xRzrEAUm8H2277NRyMHE6EQ7kPE8G5araJatTrZU1AEHoVpX7O53yuDnQ
hw6WQrqgtTDPY15vViUbCYvMzJ8Mi/SD64ntOqM7MpEf9Yl2HsNuhY4yw4jsRep86k2mYyA1mTH3
BOvrkypBJXG5wxUsV5bBOASuwoILPRAZJpWjYJEKo24TmW77goRYDAIHnNZ7CBVmz0KGBoPiP4Kp
Wo/Y7T0EKkSuDh5fgTZJwai5kw+Bp/H0bxtzGkio4fJgn61HmznfhiUPNpnnN6vETUyWZH/zeWAy
8Q82aVV76pkX5HJX0+Q4k40GKZtGLVLxEbL2kQhfG7rla5tK7d5NP7Fo158v3jYJC9AR3va7Pwe+
sZdtxo2fvj3gtdaMoQFLnpiGklKFyiQNi54lBanhD4RB4TZvSZdZji43UffRTaCe9A/eUotGYN+E
a2/Qr4yGqPTeWF18fTfSQIQTJslH0WPSNTWi41NxB7He2NHooHfKyQslFuF9a1ye4pKrXClqBo6o
zfVmG4+X3o6kDDfhby236UtOBh4t5oRxEJpjZfozKq2hv0GgLicJLTu72Ti32K5OauEjE/Qg0pL1
6j+0iRgZ5HaOlmbTqNz0H1iGTc/pj8lRcbYD/bKHvArp/wIGhVV9jGcqzBQ4v0NXn6lAAzbldeP1
B5q8QFb0jpNhwmvv1JI9Ev4Gk3Wqour5hOw7OfkUIIifqCd3pSAxESPbseAsL+d+gl1vVIG2KYUd
mSUYC/fJTUe4Sv6PEscB4muXQYYksAmxl1WJ8xtT9q4yP1UgaxK8dUBhKqYR353wV5ZlsOenUAMG
120sUNfb6FwUS21D4JY3NHuqU832ElAHvvZ0GMxU1sC9gk660dv9oaesUDsBWSAcHCNqhOEF+Tg+
nXwF865EQpt2FY7VTKO7KoxIJZlmbSQ3lixOSPbOe89KSAZQo5LKZxJbSb7gAJdd9cWXzo7Tue7n
OS9XeAO5QbdDUVd13ZkYCVjG3ShDFZAHTwUddar+r3qMXpzF4XM0juGdLGyUui6IPQoXm4pxtHGt
c5hBvWMGzOQwpaNMjRDH4N+piYIUkOr8LLIKneLXLs/DvARGsNRmNwUvWvcwsKw7FUJ3EmAlmbjd
QyjSBnQpT3GJ41xt9kd24HjHplIZfez0ulnoq6U8joivguFnqWJc1Q/WzouwpDz82BHWFaZqR8rc
a8PFtSdz6oRHs2drNo48n7WAN/im5E0zZuslmLM+z++hwXdCBMo+xVnq1GRucOJ2U6bs346wZL7x
GMltsCybUWKBaeIOvee/prIuKONfyqXeaudtTWpHv8TAV00u24Ux1363zGmj+2wWw1l1gPqf9QfR
SuFrTB9+6gN9QK+I03s06C4SjOSEp6nocGmpJpFPANstAOaNN8IUe7WamPVGdGGLSuXobf62Md4t
DgbevimAAPT042je8qHst+A9Spc/Up5D+tL5+jPI+4XeJZmW4hGbsAK6zc7BRNwjVv7ZNWqwW35F
408TqDnHPDjzpZxl4tmMilIDOvkAuF41ng5yYPsivWPsVePIcHVdiX1i59bR71hPebIdLMxqePv1
jRyYC+4WLdKiUPECcn3YAN/noH52ApP/oRAHvm8xKN27Vw6aNBBbMrucHdojPv8iKozUL7DinKj7
IUIOwBhnpDKkPpecMYRj4IccK4o1fGT93RzI8S9LGXlYnTmuA8RjlhqCnda6JMB7qHAdW4Z26SlT
QiQEeLstwnSNQab6ndi2EKRSbfcxnUknQP/87q9jeeYjRoTdp0Xz/OnWvDUxERvUrTNeNA/eB3xQ
4/7Lvpt9kA+sMq++R89YG+WUQWq64OxiTkyoFCeWYUjlLyS7970sjCMaLITCMCM8uyQJjgSuytc0
mN+D9HNApGvAPG5NI1mwLdzVDnsXyw2YRqHV/JDqt2ptaf8lg6CJl8YoDDRvj0XG2kfng3QtCgjc
/PI1k39m4MvsaWIXFNfMRxtq1WRsqN5Rhgy+jSlgc7A8BCa3ksBvIZ3csQo8xEzwKS13E+hkUsPJ
Na7sagjlMEB125hM6CrY7jm/CDLnr2OXDdW511gMZ+h6VBr76aJcQQVw4xjY53B9t2kDuypvAoaD
+QOkikCfZXPfecsv5+Eof4ZvlJxH3Q4II24g1Yzx3QskBPKb2h1lwULGElvs0BUm2WJfBHK/l55Q
7zIY+yuIVsOi5eaNmRA0K3lqhYns9ay8QCzLUsJjIt/AljMRkkwPKa/cpUsU1CroORbJDfXwQbha
a3IDIXHsZGcS43pN4h6z+baUi4FzbF9dlPDnzTFru5qfj48/ZE0UOHq3rJHAD4jjtob8IyVGYsTq
KFZJkTencfnp2+Gw4N8xnozAGY+/BFEEYzfJdCENbRNw+2ordk3tWmIo2ARsEt6rOc411A6qQ6SZ
WjQw5sVFuvxk/6pD1+N5W5Rs8Lz/40eCWmjoBuN/XC/vVFLAK9IGOikgrbh+YJnIPcdz0PCZ5Ufu
Iljc7v5fTVntqiJ+65I7qzxtD+oL/coi9pBeW5Pr9edRYYe16IBCRH58pQQbsWPk/mzwWhwWMF/X
yuGWKp8hro58xqOSYOunB+6tC/2faCThBaHkZhKMZA1OoA2F28zBI66u/BrbACmfcg8byKROpnfh
wFBmavMskIAdZb4f2Xyj30GbvhkojvhR8qXY6rhZJ0GtHOPmyWkg3j7UuFC9z1eK6Z/MunY2nqhO
pAtNOzDudN/g/zOrvvOgi2XpM0XFNLgE6T3oACvNXNfAmFFh/lsgjTP6sFqxnVUVXczGg3CIqDm8
5wDby35F6a2d3//GQfhDEXcrdK0j7mOlx2rGFh3VVjVPL3WdhzrvgRrH0ge9amWWquFNsLRs2DlF
Zcn/Nj4+t2cxFK1fXJD4yKkUFqjE/IiWgScgxM1NLCLLDCU6D6niiGBw8YFhqGUt6vJE9Jjoouu1
L9rDaJYDmB2rvWUuHxGtyipeci3leFUAN1xxPM93bmY4VXWvedDlumtssglL/3K2ZDeOEUZHdvAa
SXopbkH8JQVpzJUm6arvdvJErMx+Do1gEt+nEgk9kpDREN7mWHBXdnZBT7m6B4kat2BwTq0DV3qJ
L3j0trrV6CWF9er7y0Rv1PbnIdVWhz2yovwIeh451t7K4jygpGuZwSde7JyTu5b1CLRNey3kdhbz
Am5MM2M+uTeJaj/bc6b9LIEHhJcansrQAEUlk+NpIjsKFFiM8Dhv5YLlBalv10bfWtwMdAlV77PL
e7sN3ja6dX7jCbaH18EPy4liNAZvhtQcy5jgmIZ9mWa4V3zk1TBR319PfuE6+GJNDzHK5X+CL+yT
iGJ5kxsLZxM7Mn6cEiciBeBVScaUnJMCU3F6RJVtll4xb2ULAU8wv9Eyr6qJJ/wrvh8aCiA+czqm
ch3S3kPizjL+kfqnG+VQ4EFEvvjFkzr9oJJ2up20SLT2vL/npa4fLCQWhUN5VJ60ig7AYP4/uB+P
NW2gXFIClXwyY4TUrT/sOM2VVyKZcUH7NQ91k4A+p0oOcxNVLg49whxvsq0jSW+PpOAta6bfb4Ig
aLKu9XBuEJuzvmJaPGwDm7d29xgroSABDPyJh3UeCohYrkIzlpDRS8jhDfPJXovwe9bPyVDgZi24
e5MjWsEg8gIv33Odm4+CCX0TzlarkqxuA0cZ5r9iIo7V2GQlpQ3C4T99nsiKHJ2Abpu2TQ12uZLl
li/9sf2dRoM8xiZEc7vParhTxmvu0l7UdiD+yJWxqd2ZYhynyHN0XheggrtXw2935CvsQ998mc+w
/+eUHogqeLHWJ/4lRuq/A1t4z8lh1cM7fRl8L9/1Y2iSifJ8KwvN2bFFWoapRv7eD2tlut+XMrMe
LZpe7azi1i8zXrwBjLbR5e9izTI8zcdJ82VGSP73XyY+nxT9LCdJuhkE/GXZISnGu5/aWcRppHcU
R+viGUENOtgkeGj3hepc4mpW2dLUZgWM3NX0L2UUq/Hcqt4Vw71XHI/9GpoxlxRGTdEKph4MgNAT
vp9dL3sEyKxlY8la8b4bWJGePDiHe0hVpHk11MnSJjsgvOKloSONdaoXwlppmz9gnF9dYMuqfBrS
9GJqZ9KuVDnmSnWORYjPXuyL54FKvplA4bLAbmjz0Zk9BeUoXM9+yhedjjzoVdCDM8bnt72JlGTo
UD9xGivDTCFoCD81NM3tIJGSysl4c6cpfnH6i9ijQhsMyXCjQctJ9UFVvjV43F/52S4XoEh9xsor
2++++E7K6aCJNysfspgGBVgAJcwQWUUHw2nWmgxjZY3bMbti6tbQX2cc+gYxmhoJIHdVaRMSO4Kj
NoeAccuxUhLIczjCe65UcQgmxLtxpmPyOFU/U2t8UzOjWeoSMYmnk7EWOJnOSfJLoAu159mIWIwL
cpMmw2Sv5xhgkncUSt8VmhKrp4pVhHs/5qqDXJiBExJHdxTGwSCkAyrHRDkABdon6B3BjDbN9k0C
I7nlyV+7UnhFAqXTfv9hQM+0ibOVqXa0V53WYwtbZRhwZn5xGeJH+2TXpvJqm1er+2aRZ2x5U+t3
0yex9QmL73JNbBTRuv34ck70etLS0SFn0T1ZSmUCXeCJQCYWdGDJg+ujUL5FDayIS6dyQXXeJa13
9GWKm3rXDSMrQKflCtjr6MUGjhbpFkF+Shwdl2XJal4nqlF7ESBfiAKnXVqS1wd4QHbyAtiC7vgx
y/EjIxx7kEBqxfWthHmPRY9pdppiFdWZVz7dQ0IuKayMI7kf3O+7qebOv3MWhZPbP+76iR/MuL8N
mU3wbvnpj9xivwkMZpRx4C0cPCnMIlyBsY2X4DfTgGEtF84scTzVgtWn1rFzGF7NoQwrcwUkccWr
E32n4mDFLBA1CX4TY0/k0WVcE9cDdcxzzm4SXNWZh1u6xchKdfPxMq073TtpggyH8s/kCW30+xnh
+2YzqAubeUk5eq8ihUOH2yTW1uDkaUeAvYSUXuf1OP8BePl89dzF8jQpXxrz9TiSIJQX2Sm75iM5
qvoPqS/bZutuHpSOoUiHK4Q5kSICQW2h8aUOpfgvYSJP02B+YpSlXe9UyUfvAIKU8hTZpxnl8yvW
tPu2bOm+S7uPAKKgy0oH2yKr3sskfizFfk7dr4YaGVKYvf+ZUOvmNW54pzhUoesqqgSPM1NJB5j7
KItyTGf+DmeLEaxMFRKHqbxq64cN5jcFawHwVPQ0xo+FYSKg28o7WBIBYOyxOD7uMqpX0Va8krWr
VgwZ6KLBAYePH2WlDqBW9AS7RlrdxOoj+7lID+SdvBUJbJP74Wv5ksRSLQzFXWQU8HS6vJK6jhYZ
PrVay/T8HfhkCCCZROTHDDqQCMDgb1sBI78r1AosEgP48ACzhHWL2OTfRCcIBZZ2Wto3oieH+7Tw
03KXduhyVBgji0s2V/ZziVUr6pytHGti966zLefg0EBUL3imsHuv60sRZlncBAA2Ftq1mLYyXE22
ZsJ4kpQ4C7ARh2P8g9kF/uz9LkkblYDONEIzhAnc3R21q155FH2o7cQ1dRV9exBqG/D2Zw11v6Tv
N7jf23n7oThsEdnB4PsAZX9dqUZB118thiFrlBtgABzumvHeU0V4kvAB3YMQBw1QtprYq3hDcDR/
YP8wIIgR6f4zRkgcIbK/pQ7X83s2ZSRszcnHoTq+4NDBECmi1kQphkGWLvWn3j4jucsFGlAlyOsR
IlEfFeBx+jAcqh77wRtPO1oKd6Br1UYcLiXihu6m84U6ugU8V/gCZjflBv5H32qQen8rwL/+BaSF
IBQw3G09JQUm9W94XQB4RdbawXCs87RWqsV4tPI+NJ5s460sltkYk1HwSZRBbpznVdRpds5dN/LH
cDqXtaM0kCkB+OA2bfy/6taDAPeuiSMwJN0yVguNCTt7B8aq0TmdMve9TA8pMLo1pW1anmu8Kg6V
knzpIEJXGfrgxiHpW+ZAWpmcyHwGmIq5Zg9n8wWODruZfgMTeR9wfqUA/8LVTaI9vvY9nbbmfONt
7LP3W4BUPa1ICrdWDz+eDOb8+2URNH3IUb6r8Qr3M3DQ7sdokQ7SWq+GMtcGbfyRcHPP2YkdLENb
GbNXQCHV8+FF/WXBvmNQJzNOo9529nFVpIZU4H9X4/E4v3BKurwaQoEPQWGbgtN0X928R/y9IWzO
1eeZiirO3biTUtqst3K9U4Zcs79jK7nI8bqMihg5jRW+63x34u/DyiIIwfslnjbPe0TFj0kC+Aw7
eTEDS6D9Pblc4unwflW4nfiAa1MX/CWOaRl5G/94X2L+0KKFCEY4f3ccQT2qPrccRP3ofCrU0MS2
AiQc/GPLaVUJFtpY5fC8cQTPGxyO25+3lghNAFsbmEOoGTwa9952d2Wz87YPKsHygfCo/2rYTUdd
J59deuGCOQPcmnP/UklD8dISW4tbRQfIIJUvIfZsoCibQqagtf/fgCrfYDtNLob11ITMRNUVJah7
n6ie7gMJUxtSneI/duICXczDRyF3Mgp43NtA2MN9H3Ofn4bvby/MdWn23xa5HVDonqBcHgDx8iB3
t/M9TeXYvJxcunEN4sW/c5jlPY31XtOE4HLnnCjS9jtMPxh/6eKRixPA9pkmfPDn91GxVq6aILQi
YRGDt2RpqnQF6rClCsafxoOSiIm1fm8acrLNRL7+9mrtyUb93OFY1j1V1ZF2rtd6Vj2L2j4+uZC7
gxcWDC+RiUu/x6ShIQuuPan4Fh2BFeaFJw6RDiPqo85dNCrcxUeYeTvSzS9wv97/TpT9NDLM0EAx
ZSdwcEO/jJuhdtJaQPRP5K2RPV/RQE7MBQ6pKVkfH6uku8DnxXF0IPRkEfvhO8N32T5YtVi2fz20
k1u25kWqYhsGoV4jcq6VtweEh5Bek1pQZ4cQbXr2oSM5uM8/w8hBDL4YWnqSOKHOlWoTODIEdCy3
0+WxJkPcPZNXuCWlgpWVKiDrAN5pCbmc+cLs+ntTSSpgn1hb/TdqGaHUjtb+L98nZ4qaumGc1nFR
J0fTjoJJpzt2QDVPBCE+Uq8RO4g2fYMjLCjTR9WMf8qzF1YsMh+BtCHUYsZuqZYvLcWzlzFf0Ua3
8e7UOcfxSkMwNi+TdCYZyo9PBO0bCXWGiUTbrxUZOm5HeWbI1mcMYRUyu8XdHntwPBC4qQVh7wQ9
Bu1mEJlWi9z/HUg7ji6H51KaKOOAIuQ93LyMZCi18tvq+CZbLbKY+W15bSnBNV4m4saLSxAH7TZQ
Ntb09sOnFFttsgMplknyWtHjTqEQ26YEy0fqeKaj8JLrX3emSoQtZoP2m8K10L8OFi7umfTexR9i
LYo+YtC5zhq7aPIe6cqJyXIYy1HbH+UjMVMLmIhjjNeQjcsACSMfBdplFY89+UHL2Yu4DerCIoOo
p4L7+MC1zx5hVu0wbViRYUUNZQa5uHyQJKNP4hpDume3q+lz1jYXgFjchcMVurf9wYlzoob8S6vd
AfDHlb5QfVrb9yhk5UUqFKAFsqCN3OEXZcZyxXEKh+n5gZ0gUO/i5+CUMcK6BiczeDuoQuHATJVX
vMkNXNbTplsiemYCtm79+Dhf2LKeGVc9JXYanUwkk9oNH+89kaan3euI+fyWvfS45PYCxqMmUl6Z
rHnWRaAqLNHRDTIgLFUPzUD72XBfJEIJFlVG+PrkfDrYqNCzT8DNh2+Y4uyERZw6elmyNHvoeOW5
FXeV1XEZmXN6mHHdp1EH4BLaRnJDNDa5sLBXlmDtSwjsVxWGTBX8IDk8jl8Vf55nCYHa079MTdtC
g7YuZ1x1uEHYNvdvn+KfGa3fwaie6xpWX46yLYcnebrNcfnT7LCW9CvSG0qTkTitrsUF7GAoBxIj
JTonPMUH2CwxN/h/OlgoX6UC2T5q7kJ5aPRpEZWWIa1KxquML0Mj70fQgz8IbwUyLOIWfRYGAQIK
evOs2aSiiN25BWOt3sCd9ZJKsSHN2Z4rww7GyQZYkWe9v4afJMQHuzDG114anDBUytDVn6ABi4xr
Jf82DPYS7jMVkq+KYSz8wlN5EFOcXG/1anVTku7mTaARvjhrL/TXZXDCW3Y3F87Z3eOzokOOp+Fj
Fe4nGh2dMQdF+PSjeOPMph0RxiIxAcJroE/mE2KWygGMrjb1qiFpbNKk/DZSjU17vfV9o6XF3T0Q
s4z381xbJNbh0wew1PV71fQfUZc4L7riyqiB2eP+S2r4IAvuxN1fVwVPKYz9mjRvsPrBTrDq3wuy
Qp1ghPjXQewmCZDWEbEdOvaMGgbusm4mgpo5i6bG42xJ2WM/FzFTCv8jUtoex+N9r6wPSlLYCrzN
GY+vMV94bBtK0pkdJvF4cIPgeiaTBuDsXWIF79y03KC7mxYAO2dQHOOIslc3sObEN7KoU/IvLvXm
BR4ReZKdLB+0xDLtT+sfvk8Sqi+FDneMp/dmJvZACM1r19WG7GI3G+QpkdnNCRalbWj9s0Kz9LOC
J44JZ1jJmwspdjkYfQYOqQwu3s2k1vR49Y+ogleU5PLKOWzJd0SEv8tJRcuKcQoB2lhyu0MU5BHj
PpUV2SaVv0BPnh+2zDF46V4SXQBteZ9F4E9/1E7z0oUV3djAjdBLfF4QF2B87vaUatBclsGHxNkl
vSj6np+DCiwkCVJEYm8SW7VapHtf2SOnaXuzD49CMhqqMoKEqRtWREl4y8jWbl0cLCNmrlCkrRMb
MHjRE5HDiJ7PYefm8x8aW1YBalv+qYg14amO8p3zTTR2uqR9grfq9xOGZh0s/EJZlXJd3uFGQcY1
MyPqW4KBiP1lzs2HjDu6+jTQlW3yDa+tRshO/tQvJkRRbf2+LNvmhQpglYHCnShu4hh8E+JQHSLg
b95pPn5NNjrPWKw2zD+ktOWRXramjGU8XVb/HW7wM7MWs+cqA14OfdS3fXA4X5jnbRk2CxIB9ZKB
ZmTiw8YijQfnN771Tw9JSylYOMHsNGo2KfqrsyiDglpKXqMllYtYLQ6xHziung6bTVpqATNrI3/t
btabWx9SFV+fUAP/wBtxBo+sT/Z8GIlr9erUj3j1sjzoxCeLFnI22XUy8H2C0PUcoA4I0TL3/CFy
b/ccxnylXgNDYiz+o0EGJQz7xV8RTWrjyDtLfYnHtCeGSzFSqTywB2ql8h6k5dRE7XTJTad5KYBm
/9T46yu/4bSuexp2BGQRdcyN9XaE0jEtjlWPAdEgNlq0zAmC/vNy15XfHg3R8MdUw4ENOy1q7S/B
qPiLd5mVyeYSi84rgvY8CPhsnl9rhEQLORc44L3zxZ3Te3qkBXHyO56IZ1dxgzHaoTY4syBb/YGr
oI3/OTGH1HhMfHR8m7MhWUmSg7Xknuv1k6h2YEZSjWpYiyt0PWw3xfMhiQrJz5cCxYVqkWrdjJch
OeibGZnA1xBpwoE2efPRx+bH7DhVk3KdzLAGL5h4oczH9/w2XthonKmcJFkwpVKaOKVEzLTrchaK
wqihSYgdEeDC27q6lKDnM86I4n+mzFSz/8JP2KjlAI3gbd2qn9cVaCK7q2hv+U5LJWTYHqWn+Nfi
NcGnPJHkOSngcQ2ZWzI+NPJiIXBO/mjUKj1hpqMR6tmb/UiObqMky+GAuBWvH5AUU9pkhVzJ+hMm
b03ePl0AGvNpf8t/h+tmnt6IlLLcndb4FcqzdBaCeHmQZOgFq4+huHhgzDWyZxkC7EeZzkkipsYK
0oNYShlOurZrA7RP+mipB0KWV6NNEdSeVyAcbrEf1r3uGz9Jno/CBtukYGaoCGVQRHJY5izgXPkA
3PyqM3Wt1DPbC0dXnvB/Choj6/Xqwngaoye+k09Iiwt5yuVnSsGwEcfzd3NVvzf+El1SRbueXh79
AMZFfsYxpyRfE4PIhVhLgmImhH33QEIjabydNtkYAP7eTvAU86R93AC2G2Znr8oemBCmgLSDtU9i
YSypBqDh3M+chSFjGhn0J6OvTp+3in5sdyih2qzh7PTBrtyMhZUfyJgYAMoSB5wQtZK+Cgg1PQjv
BlO3oPc3vx0/8bzVk+jT9Xvd82yVKkvrf7JX/FSLVhGXxIaq+I4SE0LkXh14U2NFnB0w0Qo9hBcu
BC8mDeV326QuFddtRRu3V2sfqhmEhQ0YrHRdCb0UxgkSrrPZf86v7EdswQqtmFiVuXGCN03Lb/OE
kAm1JWkO9Hw2Gme2aFQkp29YEmBf2KvmtvCAKYYRR7z/isPmsO6dloiSNa/+DQIJXuSYBmUD8vcv
kO0/CLmAXCVx6DHWj3XfS+UhhXpNU2qbmsT3gUXxfGhdWLz4r3emSa/bbCma1PTL+o7f/ClwZoCX
9Iuzz/cRoxWcxyyBfnRL9yzFbkC9nsZgg6TeSYS7Ye1qJT4n3PDuYXYE10MUkV886UGNiaA16YDR
A97yUyhbDAH07TBPUfBk2jYJKl3rIXVkh8BQVL6WJxWWKNNJBwxvWIW+5/RQjRr+iMKiDfn04hcR
mPLdUof5Sc+TgbT/XOkEJStKR2j7v32hBKmaRHYIN1Miz1wlpCn5IHWYX6oYWPVMZFJN0zDYiduj
IX7JFPwznQu25vuUIlKGg+MkiB1GCv+78uPtTwUfI0649h37FnIxX4/Wb2Z2ZvytBwGNoyuVLfDV
bdbN9APrf40a8MKV0nSpohe4ZaYoFOECb2//JIAMsjj0xCdFtgg/CC2NF81bby9FNs9Lzxl8J1Ku
qLoD3FP5X5dQOO8GmPsQyCJppZg7n99ZxyjBCN128PGZYX6rPQCxdQjRc33rAOd4YqS0KtBluYmo
ZaVjiEf9kunsOFBvGxbW4g58phMZ6qNcvvL9uPLHzXVdfvTrhN8kBKm5YxK5yvJEJRRvSsfglrku
VgYYYaV6iEh7DzsEv+MagzYlOvyKI/JDgYEjVpYFoWb3v2teMynEsKC5+GpHd6lEBRAjGMyVLlIV
KnW7nuWUOPfv89XNgrzDGEk/6i56XT+x7B1r2vkYczpLQlvgTdtmcCV7iF6yXk/oAwjc2J/HyGUV
nkOHMPkYGJt+FhUuqOYjqSdt6XlSJWN0McAqyiMPx5E8nUMxphJrlxhYQ7yALwMgJ50reuruOzCG
cRGrXgwdeMwPWoRUKx6zUKgx0kDUHcO8aHhzcw8yE0kftEPfkGaUTwqwPBEXXP4sj5cEE2JEbwp2
VgY02n653pbZ7OzOpz3MvHCNKjgn30uKekuCumjDHNMrq6Y0HJpHRQaOM1tfSdgX9LMdsAN1sGI8
w8cAXm2lzeTgFgrCUXje9Ip+/zsfbS808CfHeW48MQdT1RJLko7EX+mmUXqgB1HU+aG5gwp8jpEn
64pT3QsbX5YX1646WDh7MbYs5G+T2pMUckCjmRnlzA6AvZvG6gFTWpEjnx/Df7B5/+C6QZs9M6xd
rhId+D8X24T34DzPFRXcFECBMS0vS8AoCMIvsZFdgOf648sx06mJtZJg2TZTAlIEdkEuPS7Orjj9
k/omkRu9ZNKVX0QwhKi2PYiRDrvyLhSc1AU50GrI+CtjPgIvDARRS3Eji0MLbGV4lKMHQgvG/+1v
6euC++PO07YcIGdynI5E3q0gPLUlVOsK6t6JoEeZTRNY5LrPo4zetGP/hTFNe8fBfhc6BogXMVmJ
tuxaLbTKhlFNHalYvJgw2ICRuwS5CCNuFYExElpzT5ui0bblqdc9IXyv5JTFdJUx2mhC/qn4kSwn
XHGvrSeZBbzRa5dw8czrzQmY2/QunAA7fxxIEduduGvtj04yXoYgytnlB2AeBmu6XHfnAHf/UV3C
7c77tpQxRTDa3T1CQLRm+YzYdSrU9n2FvmToaUv9yCc+/ugEziumTIjOFY1wGbyjWKXlPzUM5GmA
FZqJJwG2efMcSYC/soGGZntJB+nsOp8LCGq+PNwsSWDD8HUJvvsQK3e2szNL/pBl32kCtmq2EcS7
+eksIJ2PBZrvLJTPFFCspw2mIUfEBLRS1ISQD+YzRFMtSa8aqsLb97q+9qrfgSWPA4Tpp2wROLa3
FKK8RiZpMSsCZXi0zlgEGzSxiwXIIk3OdI4cUw7RfW6/ejFDE+c4NLX2ULO2sQxSkD6HsWpUjIvP
T99VE+seGZjCVuxpgvhtr9VpWdryDuQvrt4tGDvJ/DOi/2lDIb/sEGOpNt+GCwVqgLEMdbT+S143
ol5xkgGUYEBM150bMQLF5S3P4RGNluXZSxZGt9aunJKga+tT7XYdetDodS1db4duQiPWXqoFl9XL
YuuRlz4X0IrUoG1mXn5GrnlERvnPe8I/pRhIvGS6004x3XpATmc4aAexih7BdpmKwgsEVS3Pzfbw
3+b11pMhvGW0+Q8Xzcss8Vc7jYD6NgzSjpyWhybXt2P+RxrlOJvHzGYQewpR1azDcgHyDp0Vc0u9
ymnqeZJISIrm/5KH/Hv326/qW+7nmTva7cm6zHiuUbO5axijuxpnfbfkkiu0CkO/QALVvzsCsfzi
YMkFtIsTD6H1ft3WXEMxNaLeVaq1nGINuV9rUFmwFakMW3q6VA4YCzGeZ6WjwyPQEeqZJFPBo9M1
uepn+EJOLytmCDBS1u/hL1qau2MKbPXDkiFTtdjs/un2yElZ/3QvXV3nYNGr8PYG1hc5dJqDWtbr
FFSjOdE+EAt/6V65/l3BpGBeAl+Jaz4k8mzkErG5sOslEhv74sTlYx4brtqigL84eNpjl+dnC8Zf
m8tcd6j22BuX6Cl154zRQ3U2W5HULpLyoGGrr/DqjedZnK0yi0Mn3FtHyQiztIe3RL4eO64bLIB1
G7rOQDRGnu4PY4TGgBzzJepqyr0X0AHi2UhbRFMwzRNS4ioRAyBMonYTkzb/fg04hThO4SeUdBtY
izqkW2swW7CdnYKRRTLQ2wQLRvKFxuR+JfL14nozBWFUD+xF2BtDurl0np07ntcC90hSLK1w9EOZ
d1t5krJYEP7wlPCl9j6mG87IB1aYAq0KI0vSL7G6FpX2sSbjrR/7edGnTs+aF5bi/sMug8KO/zbX
XShymMFgxbiQrB6fJu36oKPqW8rOmaQwu0i5SbB0R0N5s5JrYz137niQozbPHDuIgz3xdz9M9/YO
+f72V97rdBGg5I0Ko16Xy0tBICG1XfRugK/chbanQq8KjOZgcRY8uLcJsBdONq0rNO/tOpSIuCag
YahsG+JmG9d0AS4bVn48eHgKlSY/FOm5mFWWfWYxrUevSVnNyyd4H3p1CxqTDkb95x6VjO5x3W9B
0g/2zURxypprFWcuF8XBlMRJXTyYfw9RRW8UOmf0+bdZ2z98KzhT20CJjoKXBlkJ/TtfubC0nxtQ
noiQJaPNtMmIfzLxMqwr4bR3Ad2sEEQ283Qha/vlIQyAlCChdrVhNWJmmnU1+RzIJEZjRphCIEV6
sEFY7y/w7tcsJZ+8NR/i7AXVXl24f8K3AiQbLLSTWUZ3x/q6f4F+iHJbyF8cygEZV+Iego38LDFJ
H/bpPcc40XdHgOtKLKFQe6UJqoc0fACvj770ZugocLYW8d/773lfPuOTolg5+Xsuum75bvxFJwyZ
eA842yUmRNGngelG/CU276bu6E90Y+NCv5/hK6YwtXqDbHMnHeDvv4QzV6j/AnJcZL79Vre1SUlN
LNbw87lT9IrYUMTsr90HJUKYxSnFWF72t+7BAcK5n1uD627j0PVSA6KwrRf0o5tf0WQkq3lQrNWv
QIfix7wtmjVfpxbbqJrBsfHVaBKKP68+ePZp9REki3CtW9iHyDLFG49nLNvHF/THScUaNCItVA5t
a+NBYLkERh9Rhk8I48QzPdbdxwM+3HkkEZp2T/7WrTd7L+OpUs/pJNEGhH3UhFZEE8oC4Vt1opif
yfdszMBWUahXlcuo0igNDUIjK1p+KUV8QLLTu9tXMMr5kwHPVupRvFLeBjoO6dOAMVMIOGHHcoc/
gxbMn+O9ZKMTrq4n7HQtHvDue7ky1nUP9H9/2B8BKTlsYQRBgFGRJyPa5ebcLbyMGq8OPJtV4moB
6PZpz7IejT7jbDBZS3JaJeU1UHfSI+XJ49o7MnaY1kkJWbMLyj+/PgL6ixAY2asBKIt7abU1Fk4E
HgNZEA+IwqqlgC8Kua54kUJcXbNNtm59niPzPuidE0tIU9t7cnVjxG48weq1MD9byvTJUEcvQyKJ
m7OEsc83W/tUnuE5KIJwmYUO40MR1MeWPiSoFsT/7NDCvmuGeNXWsGtDasFfgqQ/rVGuyuyjA4ml
67d2fLNq4y2EWUDqd04rR8pjesCttUDwgvqw0bRogFWG9Br7pjm6Y3KzfsOx7gF9ovqu+frwBcRR
wG/wx0YpinF1iXqkDMVLaQH7EsVxNB9J5oOUd/KMDSU2QiXrqsa7lTTzz4y3r0HipHdvbsqFCy4J
uVPJbfwslKIkskSmCv7VeU8lcVqqdOA0K1bmV+L+CHqY7ifnEEeBGbs6yuPxR2xV3xvT6ChI18l2
jspGxKq2wSv0TKeAfZYfF8EGfxHiAiCH6a2thZbEgPLvGFUctXKRfMi4CKsL2zMLtLt53JS8D97K
vEF5ttUjcKPIO+BcgMRiPUWRWKu63DFy7I7eRDNFGolPRP28pDNOUp7eeN8A1YpSlSCGLBiJmKxt
Mejt3BnOFEiIuFgd28+Xjr4JRQbSJOGHc5I843qMW/Hapc0O7HAUN0mWM0w0ZkbOyjf7ByszC/zJ
trGMdf9ldfh9Kz3XEcKegCW817wMj+7VnG3wZv5yBiF0D5bxCfTapNvUB95aQu5/ddayJ3DjdF3z
P5DdmmmkYAvxBjmZs1/a6oMPKrCN7BnQ+y3f/ocOV98bpwGc0u/4F76lw4AmfkN/2J9YnHRhw5w2
4jxbnKaBWF4z3TGdJ+wD3ynzpdn3Z2wLie+ZosetJlhZ5OI94xiUyiLVz+SwLzILtDq6HNdcXaPS
+6cein9RxdZmUGn8yjnQl4OPTNx9XMXtyYp/0fc9c9l594UzvjsSx1k7nll+8DZaOBzekRij5u5m
+1JVutDgXS21QK1xqoh/nkvjoU+J6vx7PV1jNX9KVsnGqPrpCJUjRpITfV9HIpb1Oz8rPbdwGVyy
d9pYC1zcokUTFpWjb+z9hdfWh3Q95WbPXWLPikV26V+rx4KHpCCVqDPICpTwNdhAkflURtxojz4F
vDrxNKXP97lGXecOXYjMiWh4TQ+K+MSdDHJMoosEJpKS1jvB9/6ruWwSmM+naLoK0QvrOsCBoUH4
inicE02M1l2G8hRqovg0KSaa1c2sXXyi0vHqgGtONqE4Eq6CyjOP4qO1utcBF//Zmz9NDY5VkS4+
36kFjeHkk4fusN64pQr9HXeDmrvXvA3hEWIe6I77/V3GXrd8JlZGeJpMD3XBWBCCqiHzfK22INcF
XuWMeoJ2rI1yMkrx8k958gjzhotmFP4HubSqBnvJdQPg2Wb6Q8ADTCwDycTVDwDlLsHMxtlqyOVm
Qq0tosVIh5mEGZlwjhcGkZelVU8ofnOkt4ZKCOC4J1ODvEC07xForZFEhra/6SySdrAB25aqEU38
g6hPa+Mm4tCmX42RjdfxzodYj9TWt3r08E26KiLkkaQazMPVkr0R0LJVGTh7Yvj/opAlxPQ87hQo
1HG5v5Rt87JXDqUjuPFq18ZElun2N+cGcTBt9tEsQVco/REn7YsNw2GwCwrXUGYGtdLQYoj46LQr
9rlprfuUH/9W3rJRRvho+9poy8dF06DZsntdN48cvXKotAKp9VhH7WTCh6pgaiWmDNnvxC5+Cgfd
Cju8MJZ/vGXUP+zspnAbIJArLrDd5he1JSxy/YAAcKk9gbg+8JpFmEt2dk+SeQ0tuf4bN6+OQSW5
sIxuDXrzT4VHH5+dYfeaMqRQLNp9qKb9qD4KCAlc1FgAS3u+42NBpkahywx6hvhIpin8w4tJSkBV
zS9iD3Xj5/Peg8BgYWJ01L00YxmRr1kgQ1K+vJnqYpf9I3YK4INQOrfzYGhGOElp/+VYxEvtAMad
wwNvxkd2estkT/cQhGAt5SjXrN1WdTKsTAgn7P2k9G0kuMrBwG5r7SdGvbLhCJk33aOpDYHNnqN/
uBercvxyhmenuSjgzcHsIDLGPvbGkm59ABJWgqrzNGbrfI6iMUjbSzZtz5YF/rfx2dcprtoXFHBi
HSELQZUdReViKz3tRSZxMwKFt/42E0aGZVjtWSRpi2XrgG2iZRGOH8wXuQCyMrq0W6eii0V0Dh/V
Dayosg2/cL/fy92ESyt6AiCosVggrgwainvfUxRcSGh/PHYBcgmejPmCUNdJsH6oN5E60HQ9CBdR
6Yhh3qYy1GxQuOsW/hhmktV3ixCQ1yjFTHNaAd3jX5lWJk2c1MUrA8JQcgzX/8uzmEC7kXEoCQuh
aoNi9hXiVdapqRj7fe3hXPOpPUzlPS/oCw8PavyA/n/5G9Nohj0PMCs3f4ZcEUB7h8M3KEvuoa47
YI0lJ7JmguCdZzu4FI960dH4VCpCxSJqpclLbC/ayy969kMlXdExift7mKL6HwkxXHzH7H00GgRE
X5t1QazEJe1+SMbnG+cGAhwXxmm6a2r74IZ7KLfgv25Iu2Si1n4h1ff0fso/6fNBkJ5Jc3N9335e
oTmwC8mB2xO2gpsyPYayPURVVZCoOMI/erCMiM/WzM9p0RK2WhBxxOGurnxaW9n6NKbo5VK7do6O
WNBYVdFsWve8DiBPezrk9ZKwCm9zfW0QmJl2u9/iG0IqNodMkVYkodizzKuVDKI+jXtOoM0gErc9
0lodmTdCYZ8yTsISg9i0tn5hv1BdCRop9UQEHRizwN6iWVc8qEqOEVOMlTHzgIvSCFWzwlH2vo8O
74DRQtNJ8DMdOWgDCpvO2u9on6agTio3DwpVMdIVfuUrOWcSPRm2TJIS3sNMyVZe/a+dzuRSAJTW
Va+JAkfcXqXPYFYQlwBmUaDEPVIqeFOBh3WJESA3ZclZRML0XUMxDm5AB+v5NTXjOcyHC4ZTW/cy
bCXA2OYRRiTQH75B0TQWdhaw3ekYvLk88wXuGxPiEnXoabjlDDCd9EFcQxg9s5/rZ/EY0hX1xPyR
1rav86egcWIYAPI7DRMJnGYRUWjto/cQvS/uvDLNUKweVEMCZPFYwUORM5VKgM1ZyfIN6Ux2Ezgh
TB5pSkTe1Q3gCuE9HdN/+pufAH+4+HqdHYNwPlaLQLAsm1c7AlVwhhlKLDQnfN+36u2fs8dLMy2J
f2zDOJTgsQ7mtYiKoLQih93FYsesJrYHxhHT1gWIEvKnGSHTd4t7u+vZKaoSGZcGS/lp3c/aUevh
8+mwxcxB3C5vZft8TFz2buSb2hs86sMrQxZwDAlLy3peny0b/PTv1HuO1uTmnNXr93zP9hN9qxMq
fvA0a/3Q4Nw94f1oY0HBU3rQWgOhoIqyH5oMcgLbGB8bN+NX/nVfHcAOqXroTesb6H8nrYO8S2xj
ABqfB4f7DieSMjYfRIYGH4F6VJ8+j9Iv+NegJRGbC3SVHOsM1zUbwVcUAbOuW+GEvywBIyNiO3fp
L5reFPlAV93OaIW1EPRwfd+KEc2MMgOhpANGJOdVvBV0C13AqMiT9spT6sWz9fJtDdWuxlDUP11m
r1Z0usCQZCB8iyVyYQUgNajv6dI4dgTtppctjexHNNHDF1iVP+i/19eRmfX337OAiV8KvRU3L+c8
Y4aC6z5C6L5Rbe4PKgKeeT7V3rLR5Zga0qDcde7avE6OR5M/+Pdmt62YIEm7M3hviinjNNJsqkIX
9qBHs2k1nLd9C0X8O06K16WEGRoYN0WhfXvk1C4I4E59NkdYyOnLj3Tt16kGGVSiwQTpe8+6u86n
JVXhOZly6sajku9p0HNbuL/5R7wydN6pGMAzQoC43S68FGBKy6V4S6gulitaBn7BlcbS4ReDM+S+
IyYmfVaceV0SD2DxGFMTUZTRBMY2QIkZrJRm0gNy34vhwnufmL0xQmDlzb73TY9/0HvwHiQMsvYi
f8hMQyBgQM9DSy6qU/6GCbbJdLwB+NTWcItE1pzsUErLt1LUscGjeKExxZ8TWTbEM/JqutohSGPV
gFeY94PdVJd+SX5pPf0RD3gZWzJRQl5EdziQqLMHpFVe+B3eNcr7M00iOqaGb6tlDHYoFcu4fMhN
qgqxm60/w+MTowwxNMjzeZiJHz22JLjbdhrcmgrgiyVHZ2eZeTpeRsrPytfOaeYUSQfH8SrQJGNk
09V6D1x9/TWdiXdE9gXoFdQ4OqzjILJyxqqhnncmXzvyJSp5bVxMtgbj2WV3e3MXvhO5A+WXZhM/
tICywvhSA97gUZPoEGcyuLqmAMqFJ7CbRd4VzGlRfIbXoL1Nh8FRz8Ghum+XM240rGiEZwddVdyI
+O98eX64vGk5x5d/9ij0nkQmu9FeTbTGkafT76J3Epez5TIQmZ84cd/UQWt5bHRxs+OpBCXVQBL6
+AYtQ1xF2vmMmFoZT5sK3GacpLLLsL+9XKeXJpj8SWe6f+BRHh41tSazqAsAW28DXMOopTAV6nIh
fI9uBh4q94eSFtAFpYODfKENKPGDfilSDJ9BIMFqDjo1G+98oLp/c+X+d/popP0jTJaTIsSVtzIQ
/cPwybyajofa//PjPb0M/SmMgES8t3IG1A8gl1tNsjgszcHvkJIME+A/OVPPHWcun2wlOpwWqmDD
XSbqNobjtMrXQoN2aVQMdABeENEQXhSLxe0vUwoGlUCk8rUtiw5bS/DyzuQ/T9Ownmbd6FyBwPQo
pMwXKObMbQ6GnK+DxBJX7foMEU/kpuM5RIoUSZemeblubu/mBjBMKK1udzfhdWg7ug//UskaCUwF
vWWCDMT0vBFYZOoj+JatTpJltipxSRBR3wd7u6YR6kajE3UuIXs0WCZDsmObW35YodFgcOg6NXiy
4g05oJAkJpgBnkMTjU3tk9vkO2II4PWWJbcPznkYVX2cYAUCUVWdfz9V6J4mjcEtf6U5L8kYBy8k
Govz4ld/ebrbTzImCE8Y7zghxfoFAGcaqlhJ6Rfirxs6VNcNyW7/RJN6O3uzQt/UbawHvAH4EL6a
e/j2LAbHXmoJKqLqfbuHfsKIc57AOJnvk46Pb+szIZxVhk2x+gpZ3tHH/Fuj/UtFdkuzLcYStlEu
8dRyrhi7Uvoqhr7frOMW8WTDC+RMmkKGvUaUQ+6jLlWxeNO2YGwcdUXIJ0foGe4uNkazKQJmkpGr
ehnojRnAZ67XB2i/CTUZukgRcVxqTOeMHJk8MTkG4eFDCn3EvOeIHiMdhOxNBo47nF6BnXulLAr0
s/TZ5+g4Yhs2Yb5GtVK8H65Al6IdSQ/wkFteTNA3+6GgHPM2vhXlc3QUju+rLmZcL36AMg5SCT88
B3JUvmNRBleWDOnJtCyphqWvG7EO8iKE+H4QedYqJsfg4cbaEdxYn1b3R0faRsNUkPrvqONiIPw1
zsTA0DoOWM2HF55wJlC/cuSF3y+lZlfGeCAvBTgPVCi5TxbJ0W+bw6LJDIVAt8p3fqbk3nUcJJLq
rcgsAqY38U+dMFTtMGPERaoLXloAFPxbEUm+QpZ6FYIeFW4v26+phM+am4M9WKA1PMo9eoMLFsfi
y5mSMOaPJ+HkSmayf//2FQ1PhcrlDuTMkWArb2aBzcpx+tGDZ/mGPhPlYF+j+8DZ+/0S3tbJtEYi
Q3xocMfeB5fkiGTpXtctleExRV5eVivKH+Dgu8mueXTXO7I4+Q/mJRIjXlMQ0ZXfFrblDtmOmsQZ
k6NXkMEB+zF4N3ENaa35Zcq17SIUtFlwqZjzqeWRlp7Vcxt5T7WNsWuq3CGQJxclbjHT8htR5mVH
zVm1UH3woeijnR1yVAHS6U6u+wT9BiztoK5+IywiCNotdhywv7+UKnGW6QSn6qG//FIS+TT9rrWs
JXuDViEX7D//sQvDACr+IdEH2SCbRSJbUy69uenduH026+MnRy4OGYIpWWVdDU8pgWd7rdP7zVmO
OUyuMj54DBJdUP0RzmjxZmqRcyYqeJWwE7nLpM+6zwL2Rb0yAIwEC8L+8ghn1GW+O+ukgP4umJHi
KV4GdSPk7DA531xBZgLoy56YHWJUHQuUjqRZfrNhn5SqGOh+4fn7fTerqk7BbOBlvsNuZMQIul0F
/OIodVFmzRi4FVIJxoR+7OSPa/G9dBsBScHez7WD7YnnFx2amvXYulz/KrvYfB/OblftHYg5mbpa
Y2erjr3fEjtIPUOFuSzJQofMdR1YRs5NOWN7LCXNOR1FgSaKS8s1oDqsHX81OMaebrtl6pztZXb9
DaYFXZ+anN6QY9+eg6Qo1V305yhn5Azb0HuvHwP8i/R0LrhrTPk3cciuMo7S7UQBv1HI1GxkQWJk
U6UxCAL5ABh2aXkNt/ijZHzFESHbQGxAhzu+pf+4nkPV+xqSl5Fc3wtMN0eiR7afFgDM6dsR+Jg9
Y8FcGwpMcWUGr9+Hz3+S6i8XKWBUA8txmL/FJEQJxc+OCF6IAF9aIUluOJXMdN4kICd9bISFbVVE
w+jiGcem4YQm3g1r+uLBaHrKJPB1+5MLd8aPHz8xKtA6T/a3GrEjTydqTW5akFr1qHirTnxYug4d
+R7fFXS389qlR2Nh2VxH7X2+MS6C3a4L0/7wouQ4vkFJIJtsy3PdlpU6BIoNWtlewTB775FsIxpk
jkKG9QKBUzUP1oieKeBwZWa6uaAEngDKCI+U/hzrpzv3wiGmU2Sa/QecwWsqEw9HCMxpc8mavUix
C4XrT/bpZXXTKpwKZIqQZZoWU4ClCY+F4CxnzyDVJLPa5We5rGEBhbwS1JX9Q4dbUnTfb9/AQKdk
4mfbMvhfQq3cnSmHi38/rby+B3+siciRa3UfIuTy3go+4NpjuWcdfIZZ64gJaZSFbt6r2zdPJvlZ
ZiUTLsvJTwCtUwUS3r4dsXnSzrb1iD0pjYpX10yswMMqxxEEBdL4Bzu3an9l+7ThLRD4UFHDPbkN
VWiG4KrUHeltB0BnCTzS+HJPgxnLI35ErEljy52W5j3wK4siFXhokMEklGQatKKVZiLxwq7aEUgG
U3PaKqsafv0aWEMJ/KrPDmUk2Q8LNlPMYBEIAtBiNZ45+YklB7hfO7OaH4HUygzaOmWzDqwf4IBG
DuF1NNWUocxjfx0SFZL0A0k7TwFnL7x3Q+hdevcKldS90Yt9S0U4uO2uVH2l8/UDeE3QcBKxiGVI
JvbcGzKr1yMZTM+3f6SHyzcrzNeRXvffz9KulIPZOPOG2IwRZldZ2xxXrEkGH7BZF7svJw7/DIsE
ksTpryTQT0z8tbnvw7dX33qDamjwwi2Tj4AhL9paFpZcH5tnjH1F4TE9JZwrIKBqxq0JiXKrusu5
2YtNCqh/WY+rT+KSyxKo+Yx5ZVzAULSWtoeAX2Y/mHnreNtEg410s6iT6Zo6YQxmq0PjBGMXEAXk
mM1xSiu2b6xvcznp3p5vqmkHNCCc4PTHYIrTvSZYHfD0PEYcoTBANxBD/S9R8C7NMc3rQ4od3dWc
g8KjexyGDWhrgMA3jua66vWSMmsvn7w3dyBfim/a0c7ikZoOcQQe1jvUmyzkJcGjyy+TSZ6q6Xd+
N81dv3xvWAKLGrJIAzepQZMxYdbQHYv4vDlZpNVlsaIxhNrdVBdDh+4YofvAH3MYeXlRHKIki6HR
T9PfpI6QUng78eem6gvsuCSMdlLTwfF126pQK5L/bEwSNP83X3aL2N1xBCtmfa7eGcmHY+iUDhCJ
zlrhVxsj4kChWRY8FrFeJVQTn3tCSXNMMxj9hkdU52uY1AM3a4OqGer30sIUnkBZKQ6XMC+dk+v2
QBXM1n/tuKlsPu2/7YSEpXtRs1T4120jnYesUZZQbTWFZan40WeUFAch2PfoDDRLuvKhVlIXOK+G
/NaiRh14fpXDPFA35LDPInWEkfq4PBdAUWBMw7cJ8/ygbHkML5cZ7c7E/tH7QO0qb8zE+enH1jc1
29d2T6Yr9YVwI/k93Rsh+BSB+00I9pC3wpT39gmpDttmcFGdVBVbTgopms44Zdp6sauvvHSMY1LF
4wePj0+uxFmet3fw/TJurQNDPWlgMkK82VgN9lik+O0qdayZaWmn7NiJnkpqkkjpEO8hYGofVm3+
6HZKGy0edGwc8scWUXUvGlfNG8cWeBd+Oe5E/eytLhxYKLC6F/QXybOdQC3v2TawD7FFD7BIGnQq
0HqtoDzBZ7GvrjU53JXceQRjl54bgx6osBQNrxAIBcKqWITJNfTroVvH9wez9uZ6PEXyBl7RCHHS
1bQjKkkRmYRz09MRMrXQCLpCY6tNhO67O3L8a6VjFSS6oyLMhPtFBRhgg7nIZInzKH6W4546N0NF
PDaaI/Hg0KLeMdTF+3yBqZl+bbQiXROGFPyJY0gyHr8oCPIRjgo/wMR2dGOsa9wMyLKox8QYYgl9
sWknFY3giFZkLoRsf4bN/7p5PxpJj6wNfUXnisvuF3GqyJeKnD/lljd/a7wmOubnlePMvxf3Cwyk
6mo1pvI0qx2xG6mRp20OwF2sRJKUKn8lXKqxAuRmADAV51RsF8GVHQf1lyd5fZnqzNBlyLr7bEYp
B0AVSuRyYK4G6PQ1Irj2VqFkHe97wu6mKJpvfNFb7r+uTTOjJaRW7qqrl8Z9Eh3LhHwemR+1Uks7
omGxp5X2VkklEzM81Nf0uDwffEN4wSiFZ8C8sIRF2O0Gtu+DidNvkyU+96R9KTwfQY+RX8DLyEp1
kTS4nlolvT1Z8OUzNKcbdoXMVchtM/zy/aTWqXfgQVTXF6Yb/F7M9aIMv+YK4p78vPe9iXqP+H20
d//q1xW8cQZc3g6vRa12BbVUlfQLHWKGOFQLlnSQLP6KzLDhkbO/uM39ClFwnVvOOxEcDjPfJ14t
3gMEe2g8JA5fRm/Hsp5cZ+hm5MJ2VCylnK8KU4VE1eFYG1eS4HaaR27xI+4K7eXAuQ4SFDfoHI4D
DQ7ONusK0wO7k1zeQO6E6KRO2DhTDj5flhNjyAY/yij6d66wJhhYs8N04DyXPGVKVxbUVaeHdAJA
8iNRbusy+TrQIYQ39tKzQV5rlSdkQt3K3X6664mzX47VQ8HqfKP5YKd6RHhifRfHaa2psE6ahzqz
mS3UDYQ/byj624lHGykLwuj16SvG+B2apIB66N3aTOTgqFkd3/lRSSF5CGSKkrDyfytZT0RN1SCH
admXAyTcBSbsYp0oCsyk4gKeYyCCADXkHVIppugsRWDWF6t1B9nLG9aSn9X4yvRrhwCnUC4ZXTqH
zkv4ytVW6zD4CCEr+WDudYoBXAljj0NVJ4cDPwsU4K2EaSzx29mRYqDWVjD+B0KeWRW3kcsDbnMr
T3MPvtX19ACNTHpOkjDcMk/QcE+awD/TGgjek5OaYZZrTptWRjmuPRJXPWDFj+apKOHl33ybILgz
k/MLsEwrzyYrLq/Ri6L/SsecLecNosKG/OE9cEPOyxD7Z6nOLE0X5HLiXhU6QmaityuLYykLVAUt
zrd/S8uOKBysUQZUhrfo11Xm/7DXl881wSvLAdISzuOYb1NNXlnvsoHAu/sw2266guI85/JKr3H4
9RAGapPKkJLW3dw5WJFtLal3JDE16cZaisB4iQXdfe9wS7wB/Ls+RxkbIpjCsLaFNeqj8jUnPsc8
tYj+HKF0WaxqLav94J1aNvLEps29i6w9EAGDN5fiF7fLJfwcT1XRNK65yOO6KrzolLNVPVAWpadF
g1QxfClOU0CE8p+5MQzhxdi2bmIAhqqr5gnyv3bV6ijX2aBUz9Gs7xQ36TWaqF9KnVEae0/P0U7n
KPWa3NkikRuF6aUNdNoUthj7j2Orv+cvGvR+RxqZ4f0vAm+oT53ggQS2GjH/uYuw/gsVP0ekrnc7
L/kesdkU0DMVVrauMUJioirPSwkohyvCKaYgEidmpR6Lt9fMEQV1FbxH99qKE8hE2O/tsslVx6Lh
C1NH0oAaP6nbKyb/1GyVYFAQntjMl8oBnpwcOjUYa5+1erV+0kVJDhw/QjSpsklZiRVgyvuDUtPK
nMK1P6RKEE/Fkg2NXqFhIlxule8Ppfv1OPDsbUWPReSKaLdvEvhW5DO+u7R6iQrdh4LS4+3x5zoc
sTpzW6Qipr0mLiqiIEmHUEvQjoTC6SAQFSogcBHPUK3vgRzqQaJ6uhy6vZ8jWFSxHGstwcDxNRXH
CVcnAxNIVOQgcar8ZT7Rxl+A8bq1ZVUxu1Ah3K84p7/LOk1tudciOlv/R20SZ2hDRjH0nRQD1iWd
+cCC0GsBYD5sA/tw4FVYsLUHBhquIC9F9p8cLEfe9V5wPPVTgmECuVy0e5JZLhfpexbjVYkEmWft
SfsFhBwA9c/Wo/L1QZA7SOW8ld+GvQLN8lYR85BURDn2AhePkXTEBDFaGEqiQ+WTh2SPDU20+IZe
CuCrICzovjQ3zdhSnknYrGzWa7czd/zGz7AmYkNcs/dYDLlJh89APCvzF45HUlnSpmioO9hMWzE3
e5cmgfxproJEVK/pI6yK27IhOb9GxfpImLIPGHA9q7XsFPSeJtxgHNfvt+WJshhZb+ToUsBV0d9L
0pF5NusmoRykOXhB7LOmdRvE7FCNxQkpeXLcj85jyF0alSqv8FyZmAtA7PG624feuafB5HnusqnH
D267ivsytdMjgsZ5mKf3xi236mMJqaXJYFV0x963NXHhtZi1mcIydTzxa5G7k1YDfWQ1PnD2kkCR
sIRaVXGqAzYjHm0BmrG0Gd57NPPXOWLycP0KQRAYAqR448QouAI68TLH1BIajTPZHTGVkX0P5wgb
csGc3rdSyQbUtkDjs+YnAQiadVd4C9wWEN6dBpSyO5qxuIwporv/kExk1zyOV8bJsyuumfpj5MiJ
ZBmoTpSgk/usfU4i1mi3Vl3hTE4eXiPbqzNCTKh3kima2DIVsi9UMWFHip+/C2jFRH4R8VgRct+2
+/QpE5Uza2fmZhC3ePSHPk0MW5TVF5DWKs/imAr4sGs1nmIzhH1Gmercb6tduFviUmGXSnjB1Yo6
lWiWVfcMT61piOJsXELwJbacU192/3Vdk3kFM0Lu1ej9dBEMPyk3EeMUNs6Cg+yerPD+YQgMK4eI
UpHq9EUl6pDsvVe604l64YUDYvsFo0RZKRsmj4qw5uZjr+ZFNsax//x1gRsklA0pALK+iyJxOaYf
11NNKlSUabmfCsgEVG8yxTrVnJczz64coUODs1V/G1c5RqlfZKs/puymM4l+i8vP0/9fzggbWFig
jR11oq6kxJvZITVFuhNJl+vwMET+lZLlu7G8i6AkJ135065+dDaEpQGNCp70EOLqxbjaVJB0hdEv
0pKqZ1WUmVvBoDDZnF+Akm3/yos6KZvxbn8in6Hp3G6xTIpbGjN8Qp2Tmm6HkvtNhOlnAfPeUR9C
LBiaRk/zqVtnt2fhnwAtd+W03LWDAcd28ykiIGPCMol7KwxhRmGv7jeH9WSOQoPNOT0jWQFK2xbm
mhjYF5Jnv+4L/p8wIwr3IWKTzmoVBIw1lbADkFE5UIDiNcPeHMnBDPbMIE8x4cSYddFoG/IB1gw4
IsZfMIfCo+NKl7h/+daejbQYfDRBgWGQel7w0KkUDwubICnSXQCipyTjtoVrDjDjSr8ONQEGaU6s
lgYxX9Kx+7mhDWJmxQpyxxKfZ7fuWLyKFjcNNASjCLfwKOi2B8p1v5KD3qxWSyEOGwlUiuByI69k
Nkl83laKWkwS9kGAzNeqTTmY1c1/F1QLnTXHacjlmVaJJ3csqso9gtz9rarPt59m6RbFDAujK6lO
1rize96ENZGO4RkkN/Nl+v6JooyqrY2ymB1zxXvDkTYM3l7i0ygfg7pj6xpgQmy+Lyo6VRlrD0N8
fqzj7H1DI0nDgrQzPWsKlSeM3HSZfD/INjWKR0kLfg1RqE+lHtjgzscjhb4KY/5GA2q2QXEPCb/N
1nVzGJOPH4TLlVgAm7k0MKwpHsqLku8CpjYGhO/dbd7ughjT9/BSzzYLlfrfRUty2IKPeA+18wMq
7v5yojeVPNqvKOcxpHT0K7GESpaUhMESo7C8yCaYD9HT26blWZbA5Uf9s4RuvuBpUEdw3PlCSUZC
7oFSPiJeAUVcNCimo7Av1l39YuO/fdKfii3JCr9MZygjJZ0TblQx3o14WltUakNUn8NerbXIefFW
fUVo0VD0UxpOYMxNEBWo/ZEoiRbKSG4VcuzHx6rKpJriGjYNUSORkM6+PjD13keC5f8FhpHdyH18
m4/riWubjIJVjKayvFuvRC8nFKTi7viJtIyHJ3AmZ6CyixurFanzDBnuZdzdc0se1EF0THLWq42R
xhTVSUROnq6sCvBUlru/ijMHAkyLIxi1Ae8GQzptyomXpHw9VK8pRYgKvy0jLzLRKRuE5Ddqedwr
n14pLMaTcVOb9d26zUvoqpv0pnY9t5qxoVX9POZb2jDS/IUJhr6FFUIKszT6jX5tjwmeweBRHFdc
/2TTANN+DkRY4b3VSeMiP4ZyWjufkNesLsZPqtBP2fLcCQgal7w4NwyS7FvAeC9x3WeafOMw5Zrx
GRPlFhsrA/0Xg/u7Q0hqG6re/H1M76Xh3gdwL+/F97B/yBKKtnjEPcN3dyul7p9jYM7qo292EZFH
5JBnWn61lEdY4qSFg6flwrt9b7s3X77vGW9NxG4l7G6GMG1H2dHy+5aBNY8Xh5aKm+gf/QgIx4bu
nKoW6KGw3aE9Yp6XEdsDOcoKrrz4pRy61T284et2hxzwxTpb3He9njMyemd0Aq1O2ZEwlvv7Dpq1
3RWfzAYA8atO2iZqlXuSLSmxKvSGj4tmeV++pgPrBQ2vFsIgDYsG/71g6ikgPKz/z4P+QKuCuPEm
PPytWwoHQv18dXpoa2LX7udOoe2qs6A1TPmia6uINzPq71hhVtwFs4M+XjxML1gfUdGKii0teRiq
X2eySEchtcrU7k6ZPa6INtFcaqwXTyP4Z78slKZISPXbql6mb3F/U09d9g+9BSP81lbQrEB+agBd
SUfjdb8vu5JoSMx2/YlXry2O1FtjpR79XrHuhZLQuofRDGGkaA/ZMCkSrPVpl+1Z7nJY92nQ/xvA
EDrG8eU26PCL21fH2gn5RXCju6wstKTQihHnwN6XKLe1ziyHNPU0Ux4FGWLIO8o+bRtszQU0Rx5k
69oTnebANyiNrSiPiWY8fBiJw36SRZ6/DnK798itRyWvWnRokvSZNM+08cSRG4a+78Z6h9H6FQXe
9+KPz3IPTI5m3KwsA9MuSKdMCHcXhKJWweQBAOZjhPphZKjjhHC/ty2aH0EZet4lqiY3OdRcH94L
MSw76+IoyYm+L+uhZdtj2myZoWyil7O2PGkI0qDNueimt84OUOsiBacKuNFGUQYourPS7Ul4bZeF
tHIUdFG/bW6PcvqrZcVq2Ja+SuRKkVrmJeevpZieEM4URHIuOWpqZ3g14bX6qG04oPWnQJsN8Iyq
fFheUUeMLdcqR649e/Xx7eYhoG0sOWbxxYMYalq+XdQDLeUGIHp6/aeMqx8Clzcg1+JrhC3v9IjT
Lj9bXP+ZdtOVOeBHf4YQiEYJ4QphSOKx05RjxweFE9wnFwwLRhmh/Z4ypCErNbUn0428qUJDLTNn
8gp3Z+PUF8SG1vKbOjXo0bzOgm6fDVcfDUJywJIclbSYvc9HAa2CpLtbDr//yxN7TkojdAATYwp5
6ZUMa2COo6cpPGmdSxFH9jbyvLE5fMyGzFt2w9hFDzS+uGgoJMLNpecKEBOAYqW7b29ytxpAY1rg
gb3VHto2Cdz44avnC76bMktLA3PKqJGjqA19gxWJVtfk/fKT3qTTsQjXn+AaDoOMjtMyLJe0hDB/
tsnYBlZapiZURf7QnNNECxdksv+IixjEZA8AUKAhPj/ekRjP37vziQfQpWtr1BbAty5DLz0dgeuQ
NeUM0zTEHI8fXBi8orlTtJLyiJ7cacOP9S5CyPBW2h6mfhrj8j5bUHA6DBz16ZP5ILAwQAAix95i
SJ+WKEkk7zno5eNyT9q2PojtSI/E73b5S29xZyswx3+ROIk9uT0oN/mG3qwuX5F9gd4GDSj0Dk69
bOWNeXQHMH2T5iAMVXrOIC6KiwAxcbxOgMPWaw/d1wzP0SHfIUujcHasOnci6UngMtTzjgpd+/qQ
9Ai8XwcXxpdJ52F4/shREIPB4wpoA3a92BISAMXjGQmirJ1gxFlODJkPUwvduEBjWMciCvDopdH9
7htLKWtkrLA+jGDeHO+uTwLzMD2LA+5eAAGs7KiXXy6jiaOZdgwidM1WQatj6ZrKvwhjmqb9mUR7
Gn4hYHfjGlL1iPSZE3Nr3zFUjCieuySBQbywH2PSeHrZWOB1BN+U6lKl4VpWRGETKpqTZeNuqsSc
jjNJvMp447Pz7T8tzG26dIRO2zuKKHi61JCOjCz3GOSwaPlCG/1XH7lCO71+sKIA0hgVfpyC+zaz
e/PTAP5zkcf1jvgpjEf623CIaq02/4/c/GTnTEWJ/wFSxLAUkQuE5td3TvANfnaIkpe0NUuruaU0
Z9hCrx/Kwqjiy24h2DVAIegw5Jhqn7E4tKM9EbCIDvOtZa7EdWEyAAMnFjTc+aw0I2yTSCoDtb6g
9GK85ykk5D65Hf+4qUSZH8eHkHePxRW6nciTL4pvij60gaY2paaZ3muRiBHLTKCqyzzDXH5v+1xg
l2Gd5bucp5qH4aqTRlyk5qHgbU2jkuUA/sr2VtaU7hovuz5NzL88siEl4eAT87llAMdFj3Jaq4Eu
fTUG6oeDhVTLczAUAJMy805dg2PHG+KSf6Mb/wN3cHFVdOc7P7+YLTflyK2NYWsZ1uVh0eRZzfgj
W3EKwoW9URpabn2V0AZYeJpQ/q0qUkJfFPJN5++WuqC9wZw+vo6hLVxGD/FvOUZqqdgPn1phTHoQ
MYtYyEByntV/bMIFWgXkWdMN1yjPzrBaB8VxjyD+Hv0otma5pCutveIgQi7YPGRz9+l2fUjBG0iX
EfM63PT+REcNFiZ9S3Z1bMJYD/PQK6GZMKpOWeRWkzqaHXnwmDi9hOqmLfcRDnZ8OlAMpSVOTZWH
kCa3pM5lfp0m9Ui4uNLoIYoyNb7WNretdUaBSJd0KjWgiZKddF9wX9b6Ll3vfHr3tNfzapsQ/XAi
yuEueJwVesRuBYy4LzcRO1N05lbXxsTAIPkwFJFzrjYmHq0ljwD4GQ8nnHyA5nUKqE2fuEG0uuM/
HmdS/5QAgUHoEELsDqYIKcZ5CQT0tzQY2Xtdd2/OfFCks0TVUacxAshgt84JSvgHjM/xuoUCv7U4
tCVUlPmsm5A6gBVP10YRc/W5LTJUZdKcWxSJ9fBTy/ubu0ZwMCXgjrqF3szAH0UIaiv6bMHisyM6
LZov4WcQ51jj6XJAmCd9JYbz2f7GAAZlS62dWjGcBoLOB+iE2b16zrnwmf3F0NCA90mAkJM6KV9s
/3h1gJkw/Wi8R+YOxaRW8IDgxJPTljeM+1fdpwXPyUODdUmwNBYGoXgFZzLdkpqtkz0vYY8aQ86q
9GRViD3+uTrL/LgHiuEoPWo5lmSc410n5nFgvzLIuht+RN91YznkKe53RmZLs3JLuGmkBlsspd3V
XtMZIztuSWPDg5/DAFHk3pSzs/0tMgbzv4vM3NKn043fzZAmtJMBq9SyQG/itKkEx6PSEoe1ILjh
ov7dGrvYM2VLGFUf9pkHuKMMQA8rmWg7aCBn5dqbATiReWKKMPpYFTuyMUu8HoQAb4cefY+Ho7HC
XRVtzvYYRHQ6gx4GMS+tYPepBnp2SI/IpeonQfMB8EnFbRVkFOa/nvKH4LVRRiAPIWZX2Ko1OOz3
NHZeZX9Q7sPG0jLFvfBXJdmOZ0MjYgekPSlIl5tyelWuIAx0b6pLfRDgzRY0NgItXTnnBicxCdoM
PLtA7fsY6ljwJpCkFJPVnrADCkWpePqqR0QpT/DFD3AT3fRAbXCjYIMGUm3paNSXkFHuTxRSZEE8
GOjuVeeEHWW9t47ctqPl0wjePgLIt0vuRRflcQkgnW4LQuFDkqUwmMiwJdk/Ri4FMeHiCI3BPN4v
RVwL3V0xHfzhAa2k0Vl8e5NrLdrBj1Pd27FW4rWonAJ3alweE7Ibyco+uD0EnjpC4Yh8PT83WSej
XT5yP8gr62+RBvYc0ZxMfLlufL36GGRR+ySphoayOG+UTQQ8THXtAKFTDn8AWNHR7tlnXJBTfmxm
wSOMBnFI7BIqj2lPkKUzWKQNoQBjIRY/OxoVO67eoCAv/NvUpHQZShULQzi8BsHYU7lGUNBNxJ2Y
Fk8xxr/5NDfOU+CRv8tUm99glqpCzktGs7gWLwQBl9BG/HulCm4mrKKMV9MZOEfe/5QaU9uriA5P
KKCCU6/bsidC3kHReUVTzVrSrzIrlKFJbxuu93UmMyPe2+vI24T1ljcMkrLmQAm/JBu0dbkM/Kvg
SgHsHp2c5u/ZkgPZIx3Ciw+dZRRRvIn2p0XYWs2Z3q4N7eK92kQNZ+X6hquavqi/CXiF3+mwpMtp
gbI+B7ucJ8TcdtYkXdj5n54bkjJsQNZ4CrbNxLwqXmEjN8vFVFIAbryT7j/Z+maoDoGjHVNbT/lU
Dq2oVg7X80y4KkNcKNhkbxX5S9yM5XuIgk3JTknS5S6TWmgQ2Ghv7omuRSUnYzzAif70SKoSWsRq
a6uFtwVh+iOOks8b1rWvXVoZzNNQvBudWuDG3GG8YpgA1JArm0TxCksw2pcBPh7HSbSDbKx67tzy
j94dd5MWWWFjvGAeoKfb2ULoFdDaEObyvRMyvqVA+cvMQVJLeK+xZFZQ+ADGR0G8nS92pjgbwE4s
fRbUourSHxZaidJCS781EhBf6v+SNxYHwpxDJSTQzVKpPr4LsO4FNxp+QP5IJXAa/1zkLxis+r/h
L0LFsZybsougAUfDyGqIhk4C+rE2OMk9q8ivU1Y6e7p5kzvwVnMO3u4jKHoH+HHsj7yqVi4cxHji
C/3AyOeaAXqLw7IH0li4MRQt5s/fdIPNK7qyH5TN7glgisYSduvLPv16laPXiISXFoxKXJMtLql1
Lxkh/eBoMrMDeNxRu/QGjgJaUOhHua50dbzbB+y6Q01oeUv36yQZzfzzI4ZThJF60MtVlQuWq8Ol
aSI9xgCxAQzsMp4wbQIkwKqckVMLq3CyfIy2tD885LyDkFN79MalfWDzUHKsoc8JAscfWViAwucN
v/mRD/jgYcStv6jJC/udvqWUiLw29iEGM5RIRj0SZNooc3tkbM9mHz++ZxcDkDamXugQkQ33xXzl
UKYl+sLrMy0nPVIGCbTQkEJVoseaDUqyBJOauWiVQyhPv+/V2zHU6OLj/pVVlrzDSzysyIkRWSJt
ucf8dhpx0KFHNFzN3IqLZdlGX9FmDj7DcjY+fgqGkcyddo9+YOVS0r/3MC59s9QM0KaQG1Tl35ce
HXgOq5Fc0V5hw8/Pgi4NyunY0ZuE+hFhEgA7DgmKpqdw0mwP+05KqaBYm104o8CltwkJnsRvq200
86WzFb6eh4XugGdKTXEnNm+N0o67/LWTzUkNfJ9SkxGu/Sv3W8TMSgsCd1gecsdTgoSIFB0yVA3M
2k8zDDJg+Kisxhebb4KFCUV/QXmPWNZ3ISbq9nHCj1lTCJIt/HKPKr/EX+iah50NZS+yY7C6rd/y
hWrEiZZ5K9ExF7hq7852vJ/9FcuaIhxstSTSuLXxzAeZkZoBinQYx92K9oOXwYwTPxMGgU3UH08V
D8w3zhEdU/zI23QWscBcCU1vUoZdPsRr13YO3N0AgL3bLYNo23FHePzRSwmU7NlqxX+I3xK9RqpE
hop7qgqEP0CuV0hnNhY++kDLc7qNeH/WUmLo33fVTdtWiVRubrIwS3SMUwRuqkaFxphj7R21bUI5
Ic6SNtKnECzYti2EapbL7QpTKueVjkQ5HgM/lIyg3C/AqUG0hUoVkN3ZKGEBU30kqNDLqi0EeNKi
EKk4rRM8aLDGY9kAhWU9d2omzUjzKdSL8r1KIXq5e9Tq8l9fjDOfq2eGNVyKfZmc/RTuYkCWNYzI
RxwbdQ1Dp2eeuU+hE9y6xiy1oRvu3EeX509mgy/lqFTmDSayy6g8IUL40KT3vgQwsb4Vuwb3sUeC
h7OdsLcZPPqpErI2lIzWW1N9p0e95B+kR2KWzlQxbnQtydwD8MDqwGJba+21UghcwI2b5U/k1uRu
tjbED09O0GgRRESGrA/ejqHQlZQX6j5pZtMfZL+yjiDWGtyMsHWpRgPA0iVBdFzJTZ5K9bhDeqIo
tuOrC1XeDvq6Uy6tMJD8y0vPwxC5VjrPbP8G8smR2xNEwOcidK5ULZPxRRLVyUh5QMRyUlN32qCi
MAtDkklz3v+hZ0JeB9TslWHXUKvNKWS40LAHae6Lo/Pgaf5nZC2KFfOwBta8TzbDWeLLc7uEG0r/
a1mZ0FJqXZKhSpZTqyItUtVcegoFJ2xmnx1+NTe3d1xPjgzwNQMpvke1CcCGChNvLbJ8gNG9IyO4
v7RPho1YYkzhbbEDvol1PLn4SOQZMvGEUthYBozcS2dokUuiesyiwykS6lbpX/hvB3OOJZn5w52W
EpAyaeFQ4Suz8unfKknz6/W3DVubrX7WO+XjEIfnfACb9lYfDnpK1nMvU5hbLQ0uSrD+UCkhL6lf
4r1WWRjwHcvbUKMntGwjMwtRe7HsaqQ7XkIOWsF3AUtnScBYe19vPNT4g1FH/Vl1J2+izWNkIcs6
6+ThHPpkOkBCZZSoce72agCLW8ydjEH5S/UaJJfKiMcKGGewnf5Rxrk5CuedNmViBfNV8EizrqEg
QsxwzPfxXD9gn5h4CqNIkidOiYfEM5MisGqgthCiIFLhff7fcGT6Gcmk0fhctbtl9y3fwHQA81FZ
eTanOW79KGKZFEQEdYZC3LBbfYxrCa0HWBgly2IbLa7r/hTcu87zpS5Ug2zw9h5E9u80vQ/p551l
JHEJ6xxwepj+HwusYkFC+/OhCv2Le77mUylYBPfP1ZQ74Tf/ChTYOHGfjIPiUyCRdkfBGjJPKLSQ
uVJIa3ai2KCLDJa97eOlHwfmVqdZAkM/eqyE0oiCppHKskX7ycSzSsWigtVfDkSc0QVygfGlhmfV
OP841fZKwel5nzK2+fTbcGCR1BJ8dsI5QSR9uX0338G6wKjwP/QVZxUnGKUVU229zatPzTXAok7n
LbEB9fm4uwnDdI/jHJsj+Qo5E2wB+0FfYQDEZ9NQOAk+zKQNUN5xO99BASxk2WALohtueF3DVdRe
0s5vT1rBEAJpzqPFJ4UpONnzCM0TD52Rb7Tm/0p3nEnmwV7m10KaO+fawU4VSBv51Npk14smIQPX
u0TaNr7ABT08JZOpe5AfvGhAbHqu7w1xez2sM7P98h0FbJ4Cs5U1v6GWGVkieU2DDybjQIDOrp5a
m1yH4e1Jy2lNSUbIvMWr2vkCxPAm6zvmbuvIxNc46KB1njLoTtQE7PJnyQAwxQ8/inOCHO3m2KgC
5wnarGeyUOF6O1T1gCmOYPajkZOqKmpz+8KG5MHW7SaXYV3nhyV3v36qTR90i6qeZ1TROq1kw+mU
X6vRhdLACK7SUxfPKnPEB6ex3gUbvBllHW9hqWdTSi/O29glg89mFyX1QhOBFSDk1AQxFWu2nESf
0NEi+Yn0cqCDl86o002W2vKNtp1xafFxL5l3K8P3oV5c65EAz2E4/FVg957ESzo4HWopN99r1vlC
Kq3vvt+8UgQZ7SDQE8zp6t0BZVZ+sIXJB+xBeok4hkuY4GOVkCtmSbgvxetgrLXRFStNzWYi3eLK
/tj7/71HdgVGuG+KUiZSH8e+0ETZ5n1Eg9PWdzcjN9YItzrL1Hr6/AFDcamtYCfJ6xrZYwCTMAOr
LF0iU0cWLolrvMLBOwiChZp7UqYTa4b4pfj2PxkaMEiMLZ4PGPxgkzTu8mFjbl3uspX0wnlNafVu
01TUtKS7Oh8aNlq6GHa6zrIF43bydapFHe31MR4rTXXngnQOZOookyTL8K5pmEFzsi4ZCioGl/E6
hMztXNcVNvMeAbpd20zEye9Nciv2UbuknHxOWetIAvIWU+clR57XgRy+M4vifkIXNfzHAZ5AtoNp
T1rvzVlnMwF1sMH2+Qr1/inT6SH5Y9fSxfs4TYPsSd+TxCWP2i5VQbrXS2D8+i6njshnl7nxrIy+
13WuNTWtNAIZvm1xbOo5QucegIkJiilSTMboWR8lfKbAOZJGDVvjB5SAsQh+d19zjPiAlDbe1NH3
nAEg8DFlR6J4yIMl/wk9fmika4Y+dV8McPSq0ve0/tBpYjew/9Yj2/jhGiax+4VGZP9hn0Xo5Ee4
qipr12+Z9V4mG6UUXhB6RrKVt1ebYehWvhsImR0kjCSLzWIlqmF3ho+EoTlrOXQGXLpAjRnm4Y3m
oa0ePYNcBQnjPGNkbzeFrJzPbgY/RvZRFUFgYH+9aPQq4ga9ME7Uve1Lm2pZwqQ1e+c/nBcsISIT
Dwi+5vUxuLbZ5+fswOGONtxQpR2JwrW9IIa7AbMUQRhK/QjZrZYxZSrW02gu5wJtzRv7vKwfxfVl
oYOUp6zm1IS/sLeK3+ZRcfnAvJHy5t8UO4+CpxpMszP6vVC5rSDH/LSItDGMHDco7mY8eKb/Yvgi
1XtUAS2afnWOzcjGP4ZttIhW86IKhwH0/aocE67AHJ9hmeF12rtEBcGSSdHxJCC99ZJBCbwOSFbN
d+luZxmXzr1YKpLmLy0fxqRc2EcFdkeKvZDR2nANqKI1KZ4TN/0LUlglLIzYYJrdq56g5fZ+kW96
mOz6z3MysUhQe2wZ6uaSDw3zOqs+YSCyLRvz+HG7yif7DI44cukihoLUMKu+ZO0kyTkbdM7qhPlP
6gEO/Q/x1TCENYFg+HnESxRJB6a5OqvSRaQEouHn8g5IOC6o+90o1EnDVkJoJLOQBv48ML8JHRvk
xpdDkGnawiTH2Ii10kOyuQxyImVKiFRHwHrAlKtUQRHxf1IuH0aQWCkGmjT1nZcZ1CJvW4eAL7lH
WvMyIxVdj8zn0hn7+9W9+ocNayNxRLIu2TtO+rqYyncDuntMKCmnFONYcfUcRI/mdmQtFukmPq9j
zS2zI5cd7pwD3bJmME1uQLITZcPG9sluCrR2SIB7PD4rpPEhin5JGTu064UsKn1MigtVMPiV1haM
Vh8PBj4+TQDvgk21ru7OAvlyQ6x2XF2b1kiDAGahPi/cht+lQtACkG+rEw2Cka0bdK0mQK4RPKbr
aiHrQBljhv+XWLhQdWNC+Lld1cl8gagK7n8Eyio8mcVMwtSYliC9/d44DnHtO4/hMifbBitrVQvH
2zNH+uafnOn4lGvjcp5ddc7l1sXUa0hMKnMSxxZxpZV6w7r1+83Q/iHRXNCyziGhQUgcM+l6YjxF
2MN/6vQMywyGPMwAa0dG/J3JtAh2A00v8sZdB3wxs4drvg1PllTRXTi1HvA49BWfWwoBQ8ilZ0mu
ECjRfZYGTu/Q+KJvfbnMGSQx2OL4qaCWiTrlNr/AMsjJEq2ldwSOlJchTLt4acj6tsyhkLkdImb+
I8ufx+FqamKcb8ysT+VqW/2EtEQIeegAlFvHiH5Di6zZv0oBrXp6Uu0F/ZKlRUlbim/kdyjKHRld
z2ZJYtgLvhCDDok2GeRZ+A+XWu29dMWcfqXOctEzn0sN7TcN20OUNRcjUnJLecX9RuCxLbgWqmv5
0W0mO/aIIDypydL1t55/ajwD5tqp86yVkKqpE5rRovJm1bGZ85Y/zPjlxh1aG9hqqI2u7Ee8uMBb
B160LCO5y1JVhNumMEPU6B6Jeh7EbbWch3l/BfN46l+U4iCEDKdePEPAA2WfbbOjVc2ZZHFbW1l6
nGgiVMaknjNLqrPRWJOUVGmRq1ikoe4e2q1PlnVU+m0mqE5HPlpIEua3p7txandIin0D+aF2QYJE
SSwndAaAVHWvkzF/oTUgVaorv15Bw47H0fqC5kqgDuEE156Oi3gtEq2aKNf/zE+peQJVDuyBQW14
0gHRcOz+cExrFI7mJFl05RS3AQ9MJZ+ZMGjMKCIy8Iz6fLU2g1zJLc42dwygaDT0Anyk0Heqp1H/
l/yaRmOEdcCXM54LbCxuYOwwzwPVXCIYnBMbLXLuIk3yb5KHkWH/s7A32UdZWDrqIENSS+f9tU/j
t6Mw66WkN6yOUvrnQ+V4E5PSGMzxkfxW8bbBC8a9JLpY+ENhH7SSqcR+gvDdAuTdHwifjSqIFmFP
xcVUxo08uKtuKLhYtVjEmyAsdzvO7GWvy40UVHmu+mZPQRmtH/JlVv0eUu1l7M52F3S6K+6DNehY
k00Op7VnLT5k3BLkJdVZIIKv/vh6uquP7ytSnaX1g9svx/7zhfMZPZKKgrsMlHdlXvE0oP5dP3U9
Kr8Mr57EJqkq2TDg8Lt7aMch8q4tQLlKIIYPL9m+ZLZfx8PLjcJtSYLtL8k9891tTz15+MRy4mRJ
Rm4vdAQ7UGrxibVdZnH1/b6MDOdtN4NoU9JDlZJOVAlCjHqcWSrLfb1L/xt80qVUdFpN7w8adSmL
cJcyA46h99l1hDfXz7+G7XMzOgxoz9Y7zCr4KS6qn14+MgO+tmGB9RWhmed45swRm9/KnPW/Rp1I
V+gNYxggoDSC0G0ucutOXbScrwZuWYKQlYjDu5ZMjAQGeQ6PA1SXE4w8bLRWCYOLzbkaCCzRZGE9
0Gg4uHEmUx+a0+2xJUaTNythZw0I+7t83mP7sl9iYOXVn1UYBG8xoYmqFESs0SdY+a8B+LXXdWsp
ATlJR8BLxQR67CxNwpBFX59uMTcSQdtLU4VnQ/eonhuxN2vsWaVHeEHqVmqvadjxvud8ElQxW1jc
68JwFN6Wr3CSYwVtxPRsbB5EPz1VsY364QcpCmqvIXZu3bZm8nVBytkLstnKUvoHbOTbAEGH0ZrH
ClxlGxtJrWmmadbqL2O9tRuPlPZOrrx/iEjF4umXcciNCxGu9yUiq1MaECKbPH7Mn9VTPels3cjs
oc3p4vXEHJYvObvfc+/+5KfoVW3UYv77NZ2Tu8FR8aovLm258H/hwae2FwdfB2R/XlaVdqsVUTEy
KQyJTRnvjcp4YC10rrviwOyvyLn+B4rODyBFK4PUp4pyEopT9bB91BWiqYfJDP53OxpoWfjnVc6w
WowpKyNVtw+sDKu5lkATaFtkNnpwwDWkaQNONhco5h+BR+0/WUCcMuCzghiV3MWFEkd3llMpE5tJ
u5c7pibayRM6XZeNXLNFI16RI7n8eRYeaLVt3H/OPvMQQQvhD8x6nFQm5UxowN36QrWq8oUKwaOz
iamJ0K2UwTWsmeNVY/WO5dTWNoOOe+rQ1Xzz6YiFZIk1Nl2PxLxTEHEzmWhqS5C0JXx37/zsVIQd
Wppo/nJI0rsbNfo2ik7MOOPBjUfQH7vjvEjo1BDamzct/gCrBntzO6SgdNvmKH60baDkEhtJ0Urj
ZJ03AFwoeLndFkAxUlcD5lFD+/dkgMJB3p/JSUJopLK51h4izbaxAwN8H8s3C+/QDtGcC6hgCRbs
L2kk1gN23YtRoAYbBHGt1Q8JYmp1AHquiKQK1x7Dm4Se4T7YL8JZSQZFzHrWp3qyxtDqecovrY96
CCcp0puflLU2NE4uSArAkQzOun6t+dI3d9cCoLjZCLxBtz9vwRDuQBjYXMDVotgk6TkgYWSZiiZA
otCVITie3h+1sPwrhoHGAI7aAhTCb2HrdUZhYkNJgK3FG/v0bt+oaLbq8zOcD8fHuHmN0cc6lbYR
am97nrH4UJnohinAtU+7l6BuS02B5fZPNYmZ9GTwVvxANcHmiGcJ0oroMXxnH1YtxkjP4CJ5t39A
A506b6hgMp81UaC8XUvBCMoeF7xd0QpbtQLkIGaoE6MkPK2t6Y/fvdSztgePhiPYQ3TKtHRcCURe
HofdHFeSh+Az/AucgdyAVrz7YYWVE3VNp1lvi5YCA447qQG/19gi9s7tFZFTOXMcVarAqnHieRIn
N2AMQ1ltjOjeDsCWgS+11NYT1FD/kTq2g7fPxGFpGMnxno8dKt0MyuRMiUYHYer77VQngj7Kws/7
TW+7cn8Bfg51Qnbeb/DVr8jX/PqpF1ZfnpMEiOEy5xliINvg8IyEoJI/M/qqjX4gOR5dhghGDy0T
3+1OGs6K8gcYGfMIv+ML1IYoI/UkRBxKcndVIuSDkI4wk/CJy2GcJ6rJlyf4JY3erwawEt8MQrv6
9350dxzHuAuN+oMNxLQEAjFS5LFWf5TvyyRQJAEfqJap4Eyg2D8G1Qg8iv5D9TcRGjrT8hiF1e0F
V4rRzhnBNT9X4jiC4k/OC3naHWNRv81VHT2l8CFttNEczocTT9J9/cWiXeF3xW490bX8jWqbc5C7
LYul1o3P5lQjMDa+LTm677jOOy9DQyTXS0twCiTAYg1bcWjsGhvzGjEZ0hAKhmlHm8FfiiC+KwY9
xwNrH3QMW9CnXzhgh1Zvw40IhK4wpjpmjpHLvOe5AF3b+jFbEfPlybJfeg6GfuX78VtRrHllDmUC
Yt85gKraDytUq6JPCCCuqdgrCqZz9iV7GWmKPfxWmMKz4Lzj19qXwOCBboB6QQlcq1cIMKEcWmDv
JyLTg06gKr4f5kCQw8AAM6fmljpOlU5pRbjMrh/KWzAA/18uX8TimEg9DTZ9wRiv1lMAe3mjH/lx
gxN1kSPt8rEo41grHmzdGDyZ2mIdYBfyCk0v7LH29qROWpHpYYF8NhI+wME3uUnfeR1f6C5Up/e2
MYp7C3Fns0vQWO2ug5lR2oKHizsJ8gYzTgq8IZKdAFSHLKeeViJ0E0LGsBv4q7n9VBWCfIHDZWON
eGLM++grMLFTOwwc4SR+ujksyEt9DBLWjMHuTZpMxlY/o5SXjjbkuu8fqrb51kettjLSmNDmALjZ
349InjQSf3RMdfwK/6F+XreLrO5+PdMoFT6gsgyjY1tazic00nInOvdXp/PJtGIPvF0KHZCYHcJW
uVeVNHL6vIiN7ROloF9wIZ4HNuyKTp6/Gh+E/2lyB8DqbbR0Q3GV7Xl+WlAfP68n7LqpRJICTmY0
k9tJeySZ1VQMahx7M36cJ3Tq8uSQoSUjpvHZJHXM5cijrvCCw6Xmlw2eGouMHlglvrgsp2WCu8UP
1/qX1kvzxDR21Fs5RoTJlww5Tif6u7Fc36rJgZ9Wauukadxn3U9ys/Uv1u5rL2InIjJIOEtnw/mG
Qy1YRb1W8iR8Eele05UX+Y0wPYN/O/iLv86CboSdRREHfL5qH7t7RzVXMx8jNuCy8FVeECI3AXlk
0XvcSl1H5Ofoi3lu8nftvpwsu3wFtv40DrrvGsKagNk6BHc5+P8eYYO7uo37Hk6BXNhz8zBQKMPw
W/Ynvsnf8NpmKPr+EYC91NCDMoG1n3RWzxkAfGQonhegs2EA0ZQEuPLIbmezGfcAi1VO7P7+PnW7
8qPstTBDhGekQ6eoNf76A5hqWI525lYTkXenDppsJnWVFGtnKS1bqxYtIPUwWc+XGBzvAMWRhST2
yIbgZOHDitiXoaSD/xDF/CZ9DUb8hNG1OsyJr7Iurz26nB+yXQB8vPplbrcosEcMi+f5vVIdM4q8
A5yVhLHaf1fz5Ww7NqTtzNwHcTHYQMlB+BrEK3RF3OrFtmNCPEK/1Qw118/Zx2xUtij3RLC1EkJ5
vWzR28X3LP+8gIWQJJiXYVRxkTCs7lN/D8Bmll+NKxWLB0iFf4kdiihqaVoq+SIrKMXBwes8Bjmo
4yXRphhEoTYcHzI+srjf32SE442Z0ys6TJPWOQFm15QJkfd4DqDWsEcKgSggzsQB1JAQFoPnELWH
2KhsIjaHHOeo6on6l4/q/nFiN4h/OLs98cVoL7j39rJVyjWIbD3Q1xt6yivkJSJOhNBf8VOv60AA
lk2kuD8s5xNlyZFq3nCieweYv4bHHFROgqtYk44wj0m1SSUWn0sQS8/Q0gQAG0MELPrOZjWr3UZ6
5EhuTlVpwl0M2Y0yiNSkoKMV3R1AuF5HZmGMEcmUylwC6HgwEGEzlCIpnxMPXJpfu/mvUNc7tA63
NzpizQhBq79WLR2i8cDLbXsZmnRKbzxQwN4Of+XPL7NtA+eW2dNPsNcqpST4tslrwgR1+C/bHB3k
h9+MqwVmYhAAmlLClmVOW4gB3GVEu8PUHob5O5PtGf9K8YT9u/aUtKRL1Zyti5fdcL57hAuvtT1G
1RjHXZ589ZYEjkimblTXKtI87qyBPdfty59w85fLvC35+/aEg1OHud/3Os84HQHdyp3X7R1nmpS+
FpfhkQG7juuy0EPeEzdPK9M+g24q49Py6VUCw2VWa9j+gSOFAuaMJRhKT66c0cMlg8T63qq9EhHw
k8ppGOoHyv8ATjZLmLBIOX2J8CjWjlSDCvdc+oNgL1JJ/KL3nOZqv0gPqNwkWrkk0rbxhls9EWPH
Pv2vJerVGAoiOFxr0wwImNBmgfQ+UzFkC34GWh1K1K+ENFlXCHJg8OOiVyTW2bbouEsPaM0nJVb7
60QhkFmvoyUhVxuvAh+QGEfu6sQ3mruxJ47pYnvkWIjD0f33tY36LOuOOEfiu1yV4iJxHl1jxb1z
iuetb1EoDZgu3Y6VQavQ1TXTg4H0+fYS27AvyAUkyIvESGlDr8Rv1OK/kWJ9QBlNSDgTa96AG2UV
B/3yxZ+rWHgu3gNdKqkP+XA6vtU1ydP081SFUpKr76hGwlIimtyq6ODM6p0kNfejsJmbNQ8WHZ5f
siAHzuW+6VuxDMeu3sE5mD0uw1HRBokG1lTjZBucBh5C/zbFR9cYAtXkU6dyNj6LQsOlJfY/j8CY
Bhh0vGyztnrbUp3FmX818S0iM27RksVUsZSWAhgU1akC5mPW/Q2RG7Dh9OfIx2anl6GPfwRr2iiA
qH12S2xVEQ9DrfGsVTGG3y205Iopj490uhiqsnp1pdAEeF1UiZSACECisX1a1EqOTG98ul/8kP2F
7AbbnjyexauMNfSuzsl1oDaYv5fd/hNu+6BFgmI4jCBoqxxCPpEr9CjQ81VF59GlXqqsWAsWgT4q
TJscVl08I58yb1hQyGe4XvIEYSZcViVjsryBZYQGLOVDrZLqjmjcnpDfNNDiV85nmRlvea1LXqfK
rG5hnsI09OdGt4E1+F42f5zLObY8L10EBB2b9UlL4Fc2NlGKIYL9VAxIcA2g7P+hI9z4+72omWAz
A7iJktmXNrE1SocKrNT1NjvQMOqyC8vZUiz4bpdDiszkADYJH6VGoShwQMpOGWuUTd+WHxEifOca
/KN0MJ3d5FjFTRYxXE1Iv0SBXBqJ6swBtfFxA/AdfaQsiLUxYVhBR6xjkfbTuFO2o/W26PU+a8Co
ZWs+Oxo/GpPUwEmPdktsA8VhRwgFxPqfDN9AKBJ16L56zKixmf+d4PksISisFUzzWM+jTpGbq2b2
15zqLRSvdr1KeP171+d8FAfTu1M4A6QHzwTX0B13obmBvhuTNIKdiUUUby3pK7PNFPt987+hmt8e
U0sWFmHwBSecQaZvmlvrbo5+js00tkeOYe+hhCb7yjNOgTpGCBC6MJy0F2jh2GIS+7I39GXaB1S2
oo9S67nMniDMvJGPGeQHHbFtzc9jJwWHUqASoduplOTZyBwhZhYl6Puw92YA63armOyT9t8l7j1D
b2xIsxvMnbMlYYHBj1S7wNyFVW5tCBURxO1drklAarhjhIiOr14M4zxdYauT6brHiGG6QHw18EL3
lmzF6sHbbyjcfU3msmbeznaqVpw3VILsYBmKps6jXHdcmY+cLucmVIuhDoVx29+jWmfiCPmM4bxy
aazhFMJohv/yv2JkK6SLZy9Fzy2zeNiSK7ZgY4UnI1CWSxgUGp1IBGnNKYcZgXRADXk/U0ojJTtW
AxoP6sFsspzO8Wp/fEK+v7DEva74SAqQK6vCYlBWJ0P0U9cZblPStXReqFROP+mJFhDnDmdCohr6
hoaL2zxy0amGVlwukmDWZVNM7cK/3+kVwh3m/M50j5ZAukhcuQtA4FvmJ5wkY8deMvGe+XfC1lIn
uSd+1Q0XY2HfXsJQBXzm7pqNvWm+XiwwoztUEJ6p7gW3alNgHOYjYh3qDaJyKNTMoiHlc3EhUN6Z
pGpBCHzgqdf/1xVKbe+AD6eUVSYO7TZsnbJljim54EXPFFWpO8f8RBHOkgETeW+28V9JD++5OCCs
esfuDY1gn0hM6veOtlMvd2f2+uojt0hGHHMtcDKQO5rU+B8dj0WGtAPDrdfg5leDK4K69ByloKgm
Zv1GWMGzXsprYyTp1j4bp+K5VWd6BKNa27a0/Nvo5MS4IuMa2JulZKk1C9lLF5T72f6h5GR+DbMI
Q2dghvHeyithMg5BUhAEUCb+jfFTVO6XAYauAqa+E/qtvXhWekedmNp24/7UllOL3vwd9m8iLrqv
Z3j0fdJo0dJAmH/AdlY0qcAk1LwyAl6VOtqIGXiDQCXxUj4bkzTrMJ1EHJSrGpHq//bOey0Ngszk
kvnXrIvvUOW7kxP63gIZ4hfwffWugOrgdLBniOGjKbaXBOhnOtshdXerygrjqZtZOevCvk8+zal2
/iMyklx8HCI5B16ZGXwKr9SMgQwTfrlhzlL1WXqj9xaGCckaPG2V+7WTbrcEEFGpT3k6cLNJ3KuX
MoBqsmLgdCjosb04Vr1jdUaYyVVr1FSSyt9YycarPejMXt5I04Q7vjiCCX902670bh8OHhGOPpVy
uvWWk1sLoj25K5s+1wIwxPYZFqLoXp6hdCSJOUk5/yvzdqXNsvblbw4LgX66SvTZErz2lCoRzwTn
7OIs+KtXqxACitc3nmsZzBhskWtVnpyXexWJpfpwak7L7pLnxJuESg7mngagcBSVMafATsCoYjlr
XOqBzA7OMHj/qFzcR20pBs8gJ/LwSjKxEdTrhBb+O7MvvGTN5lL6Xvi25rSCrlahEHuRxWGVj2SS
6DIFD5Z5FT5d9wjmruUFnDaf6LoGMr4q0souJJzDfJDiOiAdBXPxcoaEIlSp35bjWfS/GVJ+YYKF
vwtym3b85py9sJyMtYuL/7IHesosx+RW887cr2amB2onc3U7OmlSFfR3L4RR/q6Jr9pA8EIfJGkW
InPOneV6+cOIRetWGlGwuuLMcdXngxf8+V6LTnhNradqJ54VIObKqe9hWwb/vt3IOueYeuOzxPEh
PJScPmlN0vnnAhLqPqDAKTy6WL91ZRtEHv1+7Vd3OmKYVBAuzyrarW+AMu3C2DDYhiaMaZ3OQjhg
2sDXLVAaLY09kKnLf7R829aHxwXSe/th1PWStK9fRkDMinW4TjJvooQgLmq2WU170vXKYS6wLAXv
dy4BVcMJnbimSn+nEJquylhhRpcjG1/mn0k/968pW5VDzDf+FjSFsEYIXPpwi/2prfwDyFSxtZnD
/bYIv9L5TmNS0gZ126nPuerLK+ch/VCqqzAgLfsTWlTnxfTWBH5EmfQWn23uXtELb+CkFWHrZRq3
iET4pTL9iIiB41/chaBnYruojgf1wWf710hC14rtgQfuUBnBW0ktDtPnaEJc6uu58EK+aGuKDyP5
ax1lPZ91LVwDeexCMct8KDNR/T6DRCb8bFj0Cg3rhL4wXxQ1GChsEFEKzN2tom7c5ZR3owx+8PE1
lYVnqcRvS/9MY8eisq95dzLMjcTRrrn3qSIxcI8ktk+6f3DVNeiT9HjMpwzYjwmuN9VqkNbUKoNH
eKcwC3vkVHdMD1A9aIGgh+VDtInNPsAMvZGEpQ5vVkRLeZoaiijn/HMcc/e9XesPByBStt2YY3Oe
mZYX5WQludsQKz9Nj2LOAhticHUJz5zkAURZzpV/u3WvXNYfYXBrFJduf2KnQfTcaoQuxB/b8BXc
/HSYShOK4McGTPH0QI0OHt/N81wf4xXHeq9cN3zb7QxaLxqCDKaw6tZiMH63n0tpSU8atBm/DXKg
oO/xgrn9qbiLf4d5folqpCBZQe1bRUGEjLOo72O68zb8k593y8gA25Po5D5fRkGysMnJN1HHlZcd
iAYvj69nXP5/+6lmr+TZ7Exwj9Z/t1BupLy2TM+htRdZwNcKL0zHCTT6qHgBYKzp85PFIlD8Enf1
KsLAhHu0d1XgbCh4ha3ZPv/e/v+3Jo8nTlhTe5BelPcmQD6VSnGOk/WkEppuHC7GzdJ58D0bZiIU
2YrTzMNn45ByhClGhXtxEPO4OPINFhpzYfqZzpLLWgPfvPUhsMJzVR86dnvHhxszSWR24J3wPCmg
Gu0uR9bifGud/+hVtvgXEJ7p3H3WGzfH8dWkOyb0jwt2NipKYxAQ+DFNkdPQwERrZo/egnwjGHHT
0KR9wcmEg2ZEjbd3FMTw1d0N36j/s0Eu9jSpR8jWUL3fYBRlEGd7O272k/9i5PORp/F/AjknYihY
CF5JURckHNhxRcN6fH1VG+yXckffuegx8J1DoaFiFF8rmVNN4vvcPfU1AMAhaXRc0Qzr8m+nQQGs
aZx7jYkQlD70VCjEpsYUwRSLSpVrzkwnRQDJfpQ3InzuUxR6XAqWlCpNEF8bzWRaSEXahR9b5aqu
tuksKMMn1gJRIgiZPUU8jXVn426wX+A3bvm4EYmpBi7146lkLJZID9HYsD5Bf+H4SvZdeK7gPLgP
w48XtI55sCULHrAJgPgolxzwui6Z9HX0T0DV72J3TtjZ8SG1kVkq0sl1wB+0LylU/x9WOZNM560X
Xihx3785YYU7QyJoWCIoQtm3OTPCMS/b3X6ZgLWO43Mi+E2IxZamLn5+j+s6pYuIL1qYJue8mf3M
wVY+Su5MV0zW+swyJkiWg/joiLOggltI6vCCKIFB6WvC1aQNxDQG4ekfhaoppt44QD9APhbA9lkJ
wkzBCe/R/jDbnpEQ9wPGnrkY5w4G2WyoHx8x/q7mP7ijUbGUUA6alUhz7Ykbnvc9OohmE0tb8/dq
VBpJZJd9XQNN/2LXVT+L67nN+mwfSkP0h5jckiP5R9/rGzWPWZ8Dv3hDddDLBUmTnnirvlIWmwIE
lES6oEFr3eajXR3naiygJ+C6eBwRP6m/WNvstVNNnWyCe5it3kX7zQKGPCNMmFY/1QSk+kKFTIgA
EWNxEwlnM8xWT7qC6DlQ3GXkGV175DvIHhCAatJC8f7Q3noFkEbFrJkOqOigTb6Cv8kp8uJrRekl
2tkU41MTIt+u21eRSWCEfnfkYJ81uRfAx3Fvj7qRxvlfx0hpv2tM6h4d1Ow6YIpDODA11iM3gNqp
YVvsXN28tiGtyq1/2gXxXlnk+MGEm+XXYqgCustcZKIIoZCKpQZ+Q64COyp8DS3n7zqfxzD7vF9d
f3XEKM84n2y89bdjJAsIP7MeM9QciEkkWYKQPwM1AAjaHTD/xwNz0reGh4KS80rm95c4maKjdrbd
/Gzx+4+aOk2ShIdZaN3FhUn9zoUYGCK9lxcbFSFV77sFOQklDoVhsG2ZMZsJXqKktD7VfUG5vrFV
os8YCNP/90v5R1gvKSABdHFVGvYgLDYjKZv0SG4jcRtPglsd/DP9uOISEmZj8hYzXYSeh4iuaOGN
R+U6BzxGq9nLTMHGRVESa9DyUBHovSBJXY0HcASChcklqFji4tVNqhc4j77+vsxSJTT7wB3hPE00
sRF4N7wQ9uy3jUbzx5B6iMGfTKXqyzH9oU5DhLllAk5VEPF2Qs5QAT+ROglG9VtQmIsfth+6OItR
zB48SVCT4aaiGjdjMLhybNV6LEYbDzFMeHcPQ6AnfebSKTcUqWcoTj8L8SpXTta1MRj+jsO4XWyp
Cl8+rtzRWYviG6DnGg5/IRBTO0unBJYe60KfEF0onXD6zGQQT5eJy2TdcxZr2xwQ3tULOD2+5jaG
CzDU8EQqOitXiYSbm/Kr4haWpQQ9XixmCMDjHKiFNMussfKQdobM0B9SPgbf/14gAAoAmfruevKd
G5qoMFSwtC+9ZmFznp1RSqxSlYX+j/LzwtqpvFoliSdf20mVI86fYpYrZvNJkQNduVUiUwmx1L73
JiiVwfmRAZTLytaASxnlms8mNrLvCWST1GSg1YkZKk5gANTULsNtHH9sl62EMm9b5eWRRlzKCcj4
uW7II669Ol26huGNt9sjFlfQcGMk1TSRYi99aNKg//cOF+DaRSe4nOZsdAVx0akFzJHqRQoLJwJ8
8EYzzPLam3IceYn2tFLL27x6CyNOu2lPexC8MeVOJJ4dxO2uz/jI/SSuB4ZZY+JlZcSpRldhSiHB
4N49wo42O+Y8SFdC1Ch+R4klJmlF4dyDV/WBolDAJt4bMsnPelUw6UEhxluo+pABy+vDDSnc4Cy3
r2RnFw5JkpO2GUaDZ7WsISwd9YG2dKYNtvP8gWOZmzL3tG9JPrKe72NkQaG3DtxVHa1ystOWTrC0
Y0gEs/1O9OKYA7ur27MybJORnzAs6sZCIKL3lRqnpuqxb+Opcqa/oPOCB8Se5pdgOEulrSyUcdMR
BEBi3m6WsEzgYITUTdUt+2VV5Pq8+ttF3nT6iR6zCDPcYC4GB533fB0e8K7DNsQTGh6gO1jCzVDn
BELK1Rf+Q9YcQWelV9XdeZ8nY4NkDv/ymHj2BjIWcFWla60xVfRBD4yJ1QzNiLfIEydBgjL8QbE+
DpqYZR6uWoM1Rk3ekY1FaB6O8+RTj8hQPAc1xoYF7yPL4r+GRJH8yl6lzxg8LVYs8AgqeyvMRgDO
j0yKNalBti+MgpgbYTSPGjDbIzluhVt6InhEArYLC0e2HCiQ64G0MdTUuGgxNOTsGn7H5X72dFl0
dkp/M1S50p1drXErN9I9J5WpgbyG9eY++J4Hqc77DInUIpO2bhJKUS1DIOOhum+lkyodLDTDfd8e
/rt7DvqqDkIpiNaRqH8IzwQQYcduZhKF85zOrmrOKaAHVnDDFPuKg86xp/fJ+umenm0lPpbd4rym
ztDWa+qms+EgidvCzhc9rduZAPT8Ye7UCp+9UUxfln9aqEMNpAUJXSDLYTUhGvg8tmbdi6kJ5tKT
hMrCDydXfj/e28KtqQ6hkHM4j3WC1tzDR9ho00g3vNljChx119Gjdpwlx6J6iGylHbP2hWB9ieNb
LZ90x5O0IQc2h4t2Nt2UyF4N6o0Y+G6lS61o/Qf9N/gA+Iu/Rc7aHxqBzC12btRK6xOiftRIO3Bq
iRmqr8fWtqOigsZhAGRwlvemUhn7U8zC6Fl3ivBOajtBdJtLyhZEl0VveQhrByOkM/BHiTidQ3Yu
MY0H6Uu3IjEVSEkS0Qazwg1FQpBnLfB+f9abqKnt6GX8hmChzugRt1mLNMAECeapgEqTsGU9EJaz
4Ce9aeYdVTz8SoKg/g5P+mQdnWPDlnYosiAEfDgCFuS8I45MfDCiOUE0IAPkC1hS/Mis6du9IsZR
aXT6scRCA4nrWy/JvO/OFAn38USGEyj6ok4FFCvXT62i6Snz1cO79UQHuI/586SG3IHAK/wOIB7D
p38G6do8MkA88hc+jr9KDJsv/V+5OTv44PbXgQ+bwt1YYa2rj6jxK3VPja6axbVxHx6A6YQJWHeN
hv1E5B6VGtGis9+L8uMbwhqQr1pB3nTtzgBTqNiIg+4uziYP7bhNo5fx9gdtzJ5C+FrmW2o3bCG8
tSjSh4qIb11m0SJjNzXkLf6K54MLBulENp9OWvjer+CLkweEh19+9pUzKeuwK9fYSaCz+3901bfu
zhTKnFhmtl/qfEVHbCK1CUa/yR4ABSlF5IMDBeZvDJ7cZiBvefmAPo06Vi9qj9pTo8tSGzIgzanO
b9Pg7QIkwUwZKqS8w7OPOQ/P+WcXovoTpKCWz93UF9BVCTYAHxdXbv4OGac89PXLlXUSdtuNhmyl
Ax1MblTG8f9nJV4XfaJervbJeLvKyVIMHFbqE/kwgsb20lFl7YFnPyJlNMC04qcQRrJxcfXBFLAJ
OC5fkB7ua7NH67EtFhgpNYwRoNvLnAt9lHUe+hqhc+KdcYm7dG4H0M1JQe9QvP2Mwsl8WIdshVFA
kRiZb4RMuNrFG23l6NLalXRoR7IVNGnjIKyx2S9jvjfjIiBigvLWyKIbzI+1/2qLBoE7+WMPmCEI
nm2bstB94KxMRkTiqQvqZlctrrrcClgTshA5tkKHrkQBK2Fsr1IM3Fbjrd6huWzb+8/Lgks3JIdm
uqaQe9U06oOQE9sc0W/ot0CnzpIYwu94WL9FAeuidcscDrstwVUfVtgWYHvt6o1DFH6DVjlCe3PY
XeAAxlUtAh5lSm/GtaOgjiDyPaE2u4Pdp3WNVEO062EJmtSr1uhA5fgUCf5aCkFeG+haG0L1W8uY
9AAppGtMImJhY7uE8s+3zpX80EdS70Dvud2zrF7gMSsEvscDXNECScWVuyFSnA67nqPzi4r8gPU3
Tg1xygjV+cV+d1qCbgutBXbvoU/yielTa7oFXbJhm5FfIkTjUEDKfxzMOiSBqkD9qgnvlbeFie0R
KRbaUmNwRmiBitiFh9t5cWkSXNxcq5Bqf4GFf/ReP4A8cyiWujbePbnoRXLBadY0S0nxrBL+ANLE
PsEmjZPXD3kUznjkw7h/pIu59ptuqKIR7qXO8T0aoyUAwa77od6mp11V6x7GB4/5a/73lyqCVTtl
wR1CVPDi9cMCvU5JQk754uoS2eEKvAAECNUrnArUkarhPvmtHYSSKQa1Da17x+mgva0pZ4dFUZBh
WIaWNQeAhIwlg72PdUWs6x3Z/MGx4D2SOEhBTBwZR7ovTyhe2wk4OcG8JttJVzFT+3bzzB6X6ynP
qMP5b2NhY3/+PiTMf/8GX1E8Gw11T3a3gawJ5+fR/s4PM8hygmMA3y7R0+x4up/hcCiWHGDD7l08
RBJAiSN+/7ShIufHc4t7GTovabtSycHvKSQINYor1zcm1LhWSHg+3Ykjcp0ZLkpXO55gTXxaTSiP
R7RMxNqE8UYMQT1H5GPLpUauAMRhYb61CfLKT5OTL8FJBUe41mmmDtqWTbPM8p/hHF08wbZwSpmo
e5quMl/uFXQJXNx93cJUCc2n3roLbWvW14hH2rJ8meCyUEn3jw/28SimxYbdcrkmZlLdeYpuFz5K
y09AJeDJxgrQYVx0hni//5sBobLdIJEBVBCTPqE4J+C6RKyBuqzNTbA57TB0+mYb3HdQ8oIsUziw
kIBZY9YBZMjS7KaOmzzNLA0sYDzZfPq7tvnzVWQP4sbWmcOODye5Sm2ZF1awquAh3H/KB31HvgNF
ECTVgKD72A8YuNEJaaaM89Sw6qyrLHJ1hdc/4x9ETQg+T32ZVLvdcEesEqD6xpjJ4hZmdgIskL9q
ZBF6AvYUTMUd7GeI7fvlPKzOURhA0kLra3WnKq+7GS8tzrdZDK0TSxwAw3y//O6h4sfUpdCKb7UE
l/7q+zOFxzo48yYrwkOewzjGxT3pBBwET1Bph5kN1nC6E53j6Updvuk+4rTU2H3eJz69qbZU2U8G
sfeoHPQH+RBsXaO1kZBQPr2pgE44G/7x8igxAm7D/XWRqZekIwmB3y12wF+lyWZ5JdAyY64DPurq
06+0u1MR+alox1P6v2BgsFZENn6Z+Ggt72WMBFjoOaZbjWo1FexIiob1Bq9TBRA/fiIe9w8hl085
P7p4nW/JFH4GYneegB71WS8auMpnjIT7PDJyJ88KsZ0w6ubVHTLXS9EU0447YNYpku3rUXRSDY2K
c6zJ8MXNJruXEnSNr8SXeNLpOS07MCH607exfT4KaAQ0dxI4XHAiRyPCVjlIPG9Y0EOkOXSsfqsQ
hFf2ZBEZF2v9SBvVBLN3sJSwq6mvYvBMaSNBelDBbxFv1eC4I4wvgycddXb+atIigSmORK6excuw
BNcGS2sMy9ijYqUCiK03+FdTfbjSP0hk6sdB/fmldyXXEx8Xr/v9yLKQ5dWghf08HaKBLYKjcLF8
Zpw4EwWDaJGCjvWZXZwHo85H22JFouFRgrg9dOsGzXKwUg4s0P9xiUSLm9PXLvNasp6SSgoDY18I
EnVdZxQY77K+i9/1uP6JPZLqYVQPlRT9XltYphvT4WHk6zJeBZX6rdc2OKVdyJr0avArSaUc5RFh
br6A1ZTus0sbiW4FCBXCml6pmuiDMSqmvq8G6aZBiBnM3D6nr0jystOhWOOk+Q/CLJPhejRuJayt
B+ESy5wNiyf9zIn0GIEdugGfJctaqAJkbo1pzXpLaJrxZESTvNS63tcVzLYqfJXtKfL65GCUXMtE
K21umZeZI0JHZU6Nqil9vNW8Fxq+SyPpMoVuAbcbOl7X9JSwZuEdGbB8Yd3Or5tPMfG/pb6cWSCd
/pXWMLrCAF5swhQZy2FaLrXgxINPlIa4BSqoXDHn51TCG7Q37mdN4CIw7lIob8JjhNVWctmtLDV6
sMT9ZGp2Zz60LLlBmiwiQMloaowP07s0ZlGY5DH2EtupPQ/udpIu5iiubnj2oHaYb+uKpkuJ7q75
iH2/UI1c0w8TCVQpRvcySzUbYJaa0GPb3M7rU+su2WWtxy/eTojcgiUQfjTwkk/B8or4S0cDyUaa
e7nIPEZMNIjQyc47ujmv21j4s+Nn5Vls6fiwpQFzIAxhG6Kz/nupDZK6WxR9BQMtSOPfRgvLS66P
YfwFb/6U1vm6AqizrubNgVbnEC13Nr3nV3ARgchbkk14yOw8EfIUi2ijeJvGFwEOUG9JNfrtRDWd
p1P3seP9AafZl70sKGSDYG/jVddiZfYldWZFW5/DzwRUzcj7iCJZ288IxP3UghRXxpVP9kYQAnvb
Gdf2QJY2hsbd/GPIz4zNS5WsF6ZJsEyPOgx82+PyJKsjWt3oOmbPeKpKkXMAOVY94D/Fe6pxA6D2
lUikyi7QfDoLo9pYBBocKaqA6F81ryowtoPq5g1DHz1NsDT7N2EzvnIrx0pw/77Q60f43ZiwHnvt
KhhXZz0a3qg+JvyyBcpDIjMBW329VOd7iiqAN8FaZWMxks1c4V3Y4ExhdzgNaCYYLVuRQwCCXoqo
bYDRKxkZZxrGj2Q56aKnkGkwvRopbfEMFPmBOz3Ljo2G/koIAGfM5tDa4BsGEkiwy131yZq7I0e4
ZvIRIA+bfOgHXigWq9l2jabTLzMdly2Se2LxOZAqAh4kM/8wHpoBzRFn0pRQQ5UhpX3ew4p3aaQe
GthGaTHtvTuSSstA5hF1K1iAVmBOB6jCfoqmdiwq1S7BcIk8jvawXz02xjvAkf+quBjcQCHjFooo
2tOoQMB54CjIfxVdo6TWkE/qZKmIH6TxjPVrPrhHgnJBEWhHcC+GOkiVPaNvRwTSuGBei1wiw9qo
aN7AE8FaTdoP6PC1eBM/kIdoGvzMoHUIdqrwajnTQOQcWUB9NkIYUWikOK27/yF4w70X8hBzJ6iF
K3CUBroBgMl5KVbJNm6vBKvKj+HITFLrDbxVH10X++V0SA9Sv8d7kY4yiWWR48vk1R/3Ep6rImJ8
xoV8GUMXaM+vwnPP8P7MyxCItFyZ7EDl0wlYyfMsSgosb9L9QGTE/LCs7UF4800FOiTeSmHmqNnK
SZOWdJpKtpB8T755eQtLavOtLWeXrNpkmnr2ASRWJlG2QHr69u/JNbRIoPG7TNRCRzXVsBcIOKzO
MLMUfl7f+u6bZswda2iJpMqmCeflPeOjZ9equUEbq9VQuaM41mRTRgvDiT92eZLxk2l8q7LI2dHC
jybyqpt3OndASBOtrNZ9/IktaRhwkOHI7y51PTdLkVHm00siZVxen9CXbajEP7Efxr0qkG1oPblH
GeoRJuCqNYVrj9ahDTatKbFk7//65g2eQpgEvpNVqXPf20RSU0OZiXy+aMijWWIG/Ty0w4ABPIb4
jpQll7RnmMlfM7U2ZuBddbCLSnsJvW5JnbPlQW26LqgL4hF2h7NQRnM1QVqDApie7XFkdrEbtcB3
Mw05kTPICKIKkas7bbxTp/z8nFWSfyv4HOoiKaBdz9ecIgW7n7gpBqEeUDsdkhFjAFMUKzbZPCST
Da8MFAB8hduhd7jixahB3S0AMaZRBGrjTXVeAzB22zgFZVW5U+83Pv3XLTAJ5McgQ2Va9I8Acw8W
4k/NDSG9P06WJdHVQFb0RxMkTWcuTkIFxtnAEZQBSAcmCmGBlinr2NZUChh/evZuC3goSJZWr5/U
WFpWWgyMqijvp867C+PBN9Bia5L5Dj2ewUvXEmYyzZqQogO67+yGHHoPn0iNHBOGWTHCyoqCqCIs
8PiXT9F+5mCF+j5Lq8/RrjBrhIigVTWFT6yDmah0/dUmnF+mCufHo+3CAJMbVhHZxxRMX3R475jd
D9ZQWfyVa7ah6MV6y8r6T8CO25d9JkHAPxXpmq08loNzw+VCN7qZBrbB/FmSWh8ms29nWY93+P8t
6xpjITQ83akr2RPyoQ+gCOclmDkUZKSTVbqUW/zt/STM3IG4C9rHKR0FJ26fMSG4u2y5j7nAu5Sp
Wr6W7mIoDstJ7E3ySjbin4RbopBjWnsWur5jqcERgrZqNmQdfanq0I4evkCdbFbWtxp1+sABcU4a
aSK+PAKmbUyE6FfWM+rYaWCPEA73NaSbZvgzD694K69hp6kGb40l87ij9lTJr/wG8XqY+Q8H6GDu
8+H86h1rv21mDOlUjNwaPUzv044/wYCRFHFK/TZPUDGkBKNe3aNtcjMgnAhk0zsIQGXTomJwPZqO
ZJfqcclW/hH8XHxXbHuJYtY5n6co9UEKpor0bKUz0XaJbzpKDs1O3jOmfyd52e5wfBvQKAjTBwEv
TfYKS6wOOuWt6oQdWcUulnBYeVXJb0pAG333MpuiAWz7PE7GDDuy8N35Q6POZeiXeHL4uuMMa1dd
ib3yWx4zk5MriQFu93kbydCoWr9PRUNeoim77cX2fV6SmNLUI6XHey6bv4njjtzvwgXLX8YTbOr+
COgFBGtJTv/hTU0o5Fzn9nchbnvaSbAOR2riZrhPmiHyJ23MHp+Eto30qJnSmz1iiCMGTejpmg2a
l18RRwbmBH3CorVbs29OAY5MKAb2P7vtbLFnJrE0gJNKoEmYxGHIyVmpAHLMuFrJRMV3E9eZB3kU
I5vWwQN6hB0d1mzYNqoWtodm+HuENAbYZmCEXfgNEc/0ffmDU76hDbt/70KyBjuHDexELLiFtKSm
m9F7n//BGpp2NwGp/xluTsqMg45XjEAvciZ0mtPHQfx9JzROXKlBc2JWGIDW1RFe+5qlpJAxPjep
tnrDyKIU3hO6kTHVL6P0MxohEUwRjiW0Nyi9wgM+s+fAM0+Qu6MT1W2QqcnuTIPLSL6xkUijDT5s
nUr4wBPUqjJILxB/RxzC5KB6s0YHH9nl+fLz55cKZray3YAQAFn3EaP5S9eYe/VrL5a59FU+hU1L
ieXGDByzbtIm3E8HNvukmKNv0i27nhZthprQeCsegjUcNzmnTy+EXXibuuaYwkv3Ulki+C+rOut6
2TX8S7lp8aywkT3MKG3ZnNfx771mEZgIy60d7Bmoe8l9hWBunFfsdcpiTOE8fNjt4EeqAKGybrHq
uYfjxusrypzbq+QpADa3gzv7qa2YFP+6g1ls4PphXqGu7SMriVlEi3Mx6o0B6Z1ltW6q3htsNtV7
8Vcvceo4Jrn74qKVMLtZlwY2jWFh3stFd5jnc9DtSvQmPD0dJo6DPDsVj4UzGLBUC5KK24xuOdz7
2y9q2sgj2W252AJL01gH/DBWiHDTnNVhpW3ZCIR3Wn73n0IWbvkKMhyfb5I5x39XYToyxizqf51u
NeJSRCw9znyBQshVlBXKhLK3dZ/QmpLIzANrku1Xaf0A9ALVTmfw21TW/zEu1ZIy+V7Jfyv4nFXu
+KJlQuPpu9OqQzUeCkjGYcE57XPomYNtZs8yoNmO/4yiAQRLeri9B89TYjp89j3X1CgALpMixmtj
6xbmdCQt28djEugFO7wMPHAB69JYN2WvhfvUW3F0TUVuGMy4Z5/dOHc8XAfqrFqjDys7NTmnQXXk
xyTfFNEFXOj5ZY16NZbR5oADu/HPZdwmhWhJs81lZBVSECoRmyoyTso4HlOTFViOrYQ0vxLt+6U6
86Ncg14sLFj9hOFgjH6QOa5QLNVwfT9+ZvLRfssRfnzX7cMBb0+Krmb/lXwt4ZxQy7V1YzTaXcOB
vfzuendZQx5nVI+7XH941S9yrCkxIjrXGgNOY/nOB6bVUapzJGTdpR0rEIEkWAf9my/JFhQK55vi
Oc92/Mzsaa/PUDPJUnVFXlP6JA36GNu7IQIrm5uQJdEkfc/OaYwVk/qiJ95cxmgXe5cSBZ0vdSka
DCw7v5oX387t1tMv8HwUGVigZcRZGBzkj4iXsyf7Swlp/mxC4EjHabJyBjBMnGhItaXmbbQPhUcw
DTHcy7td0qRFLQY6/i8jTAjbMMGSy2Uu8c6mH5LIXxHMb3/du5qr1/C2fHdzImu8s6GMio2V/zHd
dtf/6qlpKXxyxGabu7yl/MWDBSWA1yPIxnzTHOK31lcOzlt6Qc6aivE1Q1SdwB19e8homjSIiBx/
UWEV9TNRd4Qsy1+NSCAWSI8qaQt0ZOFtvUzE9RH5pOeQjBcU+ai53avHKCx4KuYy502NQN1saiOP
r1ja2Y7e5UUK7I0wQfZcB1N939ewMQkp2GOJsHJFXi+yKr9STPdHJN24U77H82yy83pAYXfNR9Nc
NtypXTAbqjskKVgjjxUL6kZdpYvOFtzWFZaTAyedTgaYif6jCeqGwc4PYuMmj3MLBW1OTQsM12JI
BDvogz39izLFFUCFjmS99LqiXZYOonAvC6alaPLN1RkPguIznEcu7cZB/jvto/3gpB/48Tc35Xbl
Kscv4UdGkzUR7Jp87eHRRJ7guB0cEyabCZlZlmmnJn8rOe6B1ZsIiyApomV6DpAEdow98tkPPgnT
Dm7c6QiNQAO6qwMM31TSmMTjA2IvX6jQdyUEvl/5zCvy2diiz9nz1C0slV56QuEVn2IlZxOEqsis
hHa/6Wy69CAIiXoMNRShti2u3tPtJvsla5W/8ywRkMNOqc6Q3scdn3EhDeYf72DfHgJRR0AocO/3
PGywBGv2IPFk2XkJ0K1+7dvwT6YsxuY+DJgfI4LlvX5UrzIoT6gXQy6d7xuQuP9x/HwrCjGFMzDw
kPrvbbnsgecSp0ujpAqLSk1q+H3LrmUaTFeGm32A+a5JU1W51XiJbHU13LUn5ub12eTvJb56wDqw
o1ATa3AfS9ParQxmq/5rHNzaOdq/oQ3wsMLeMeF8GAoXxO49Ga9WAW8iGW5pPS8+cvnVqNu7UTx0
VQGQnnR8wS5MDekBMcYgkP3nqKPlC3eWmtaTVaMCWdS/EZq3GFmWv4A2Co7LKx07z1JL/+2lqS3o
RNeOYxj6zoS9Edt8q+pj6KlhpNC3ctw9PEkQaKlwnuadHxteeeJYYLFGv9i7h2TKEgRm9Bf79d/L
p2HI7GhOeHYQpEfQE2X3Z94uvwtCl5QFx9XVCt6vF0R9jwBQGQ9Vo7vAeo0z3YysZTO8KmS6zc6r
95HKqNqCiv5q3ZC0jgspuL/DacLPuxKiFFQVu2zTrMjMs5XI5VZwSXz5zee1fG668gfljf+NV0AW
BLKM+YNx5JUd7yXC1SdITAnLZn7OOJS2vKS6t5TgADT28TRpjtH1E0oTdijooVFM4wuFUX4P5LyV
PpbSZAzHe8f6kpx+6Pp2ZV8tyy8QfMkTlmyABe9vleMP9dPvACu/aK9GiB4dEmwg6wQKrZvw8n2n
1PtHQyV1PT7c8ELGb5rRAUnYySHivMK2r8pDIjABKeLxcH6YPhDODRtemnHLYcKUwp5pZyBvgHD+
I6eXKArn7YDY+mYe5+S11FZPYnFsRBs7vlCZO1Y8823C772Mw6gV7GmyWY9AQzdSg7CKLKb60FgG
7vxh3jYoa5mCkGzWL+wBSM1h72OkhxE5QWYdzUEiXRhpSOPPXUjf3yEb0DAlHUelruXN2ZRxosD8
5BVU8q93vOkTzDaZgkGDV/V0ETd5J9KscC2Y0zTWmby4W0MLzEB0aK8QMTgG3ze6lKUHqXR7z/hC
d35VFb5ebMJljo+7FjhySUdrfXpmzFqpxfUOolykqSJzTEkzYqqVtYab8XmeFG+BoZ4oK2g4I0I4
ZDm08XN2REiNUg/mFRGXITfYtSfu/LLFXTntG3DFqdsnpVxzAR9txActD2ft218fmlc08mpi7Y8M
nNboxx1LQnRLY3UquRdJ1WjqPYuq+D9EvnjQQ3aSJ/zBgFORJ5WdMctCzbfvhdXG6W5tnl22UTHq
vFNoYNGNFbzFFyRrWfs4Ei5h6BM5ZxKQhnU+MAhYc50MsJXWhp1lOJYMCLtuZ1E9+uunDiUkA3n+
sBdZEMOe8zNEmp6Tr9HWwFjN25H5rb+dzD6NBkul27lC8rEv+cDBbE0lDerQDVlg4fKgm3SFh4FK
73IIgEb6Lyy1va3jlP88IZr1MLWfJV8k/D6LkOdt3cyCYKgwe5KfVudZ2bRy4jG1NlRjvm9SOOWG
THwzwxTlGj+pz0VdGJiYb8m6uqC6uO1wUO6VauT90jnIwBrZuqcYlQGc2uWiZre1Jg/VTSanEhP/
Ewl4w2UUneD868ychtOt34O+XWaCdnI1RZQnQLjMdyS6aRDSQN9Z5GjYPyIXLNb7nOTbPPi7OgLj
xsxOmP7i/6jB6p1RMhCramA46J2dCPgmrW56pBgfBrcWUtFucGbCpFyTS5Rnto5/ifL0kM24Bap+
1NXmtIWjk/WqUMPGyoBe/ZiOOtG49/jsLGhlTIE3CVHAHigYlAavl+9Ct0TGBxP3S8BEhPZAm8gk
txi3rEMtUx9/uUp5f6c23d9OiKa4K8ll+O8Rr4BqRPMhVZ7BKBgDLjSls2IFsSGVu7o38/W/e8dU
/s9qNXhY2d3N/UbdFk7P50rgsa48Gw8RgwlLFwOzdAqNsp43CviIe23YcZcaV4G2GdHrLhnCjB7Z
9jQDHY7q5hkmy0HaRJH0tpn06eAn1k3orrVlYhhhdArhPA9dcgHxSFnRV8P+RQB5sMbX8x8YYC9F
ZoeyL3Fl6hq6AvIao7K27vFJUShc0YsEPkR4Jazf2hgBEKrm4aL6A/kr8m9pQu52xgZWWwgJAMb0
3Bf0sBrbncfu6ZxetpRiWKUpa1277vLOaoDKwRoABIbfHQiecxLhlLsfJIeakGBwxZG74ZjJgIuU
S+fFr2VEkJRu+5V5BNGMzgsg365Q3eTVQpOeVVdsU1biexKPN7Ecfrf3ktDcmPPoFp2oMvP9/hDs
m/iFZ2+GvMo6mband+hCLTx28cOG35et+xGcL/z+VQ4ij34JycH82wC+omJz1b5dgGtjvGaYAj0E
cebvMlczxbYMHVH918bJr1ZNphxo51/RrH7c04C6GOBXmuhPnRfLo/nvTPWf+yLQxBRgl90rQlJQ
qET45DjrjpiwobZGO2Ha6Ct7bNPAUv+ZXDJRolZLSXPsemR0kNPCVfrEqceNGwhpoEgnYOw1AAVJ
gEHRezAlShOUAFmrWAGUMtgFIMdSthZ2jUBAfiJTb0zASoG/SL7I8qi2mbYidYowxXFTBy+oMSon
/XX46oii/AC5Hd26iOAhsmr0FOTsNFmY3tLb38Sj8l6KZRpz5znYpUhv29jwyiKe5ZGvUL8HxYE8
2AADUwhWQyrY+4Jsy1GTm8UfCJAjxe7gYI+cvdDtqNJnh95F3te323HQzI+BhTEOoe1Aswf+5XHo
YoGSGdBFVi8pvXDtO4OsVdozW5xiP412eDBFYQ+IaadgNR7Se1WQxSStjOtBGIpPTj/kZoUkhsS2
Xeh+B/2pLm8gJzl4VsIJQ6ixMTsQQrGm51ifGNL4l8nNeShPLCx4PMGPhqoSxAViQWTGw+Bm4aZa
BJ38jaaHdLMs0dco1okgbjQP9xYEfIZ5161z4vury5ihmwMGDOavPOrgAjeVCiFQFbAtCyrQ+QwK
J0HC2gU0NAZuwJs74LlPYnAfS55f4kKOaYCsS+A=
`protect end_protected
