`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
crsuNbGKr2+HGjsnrWAO3ApjaENLE5lmTkmDpqy6wXOqFQIJnrktoh4R9l/TVlY/BEwSOhFtvEbq
RKvf5np1ZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfoL36fNI5DjzIQX15YYPTK98uQI+Z0aMjl+hiAVWq0lzClrfpDjXWaPyQGiPvnYkkUnnCNmSyGP
qGrNm7GOsjezCGzMgQVr0792OKktWuV2kt0zVP1RUZuHk/37eznwh8N2o5rw+1YzW4dGzl1QbJom
tmB1UpBcp868gDBGaIo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nZKDyxkYA9uy2Xb3FwpEri9edMFM6SqsP4Aed0tRsVeeX445M1QANBu8GOl8sJ4QNxr6T3VU33/s
FK93SNbe96iXZq7rd0ZTftDGFn/wlb+m7r0WSjfp5pkNrLXaYMROFr5Y+cSF68dabG3s3COIhufS
z6LjxtxffkVZFl10/p5NYIyhVlCgj28/qTLowb5EYe1tZ0WPUAxBFuTyFKtX6X8Ha+x+nETiYK6i
PAhbV564AhzWOG1ohxDJJcn/sq1JfdeuDFdYSbNKycH1TqhYGY4rODz7EB10q4+UCVziUOr4Tv4R
NCotWnw5vu+fF2mIxu+vVyyYTSX+rhEfPs2iXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZ2XWhB75BM0Dt/9VMCHTjvBqUtECoyfIkFt8UyDN1IrerieLUkQavGMJnAyOgfgB2F9GkPnzVQV
7H9tsdZ87Y+A3ybRmsawN7gt2tqx/GGsvZlikuuSepi3sHN1vWxch8VpcI/SFn7CnlCh0jupM6VR
707+yLDj5AJkQVyH1LA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S4eCKuneguafnmn96ntdnponlGVTmyJu6zrxyF34ICbqsowM9Vhvgm6poU8XDQ/BrjS+RNPc37Fg
G4CZX64FNy0IB8M93ARmuOVvrGN2bYMf3jNRnVO/z1hOqr23u4iXXLcNjJcX+q+ntygTqDn+dkJa
tNf5JDJd7KcZbafDC5iOu1RcjafQnwlpqyaxuvNRdQkJM7f5tDyB/fmqWMaeSiYSf6cbwC2Jk6x0
7wUP2rAkEzcYQjkJqSGT74QQ9ZxpJuO1xNUbfsJDlmWbSmEyg55J46Q3XRBw9O4UV1TNB2XnSxvt
0rRnDIzS8sn75CDPR31VCmG8K+PwSCayofA3ZA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17232)
`protect data_block
HGwVbJA7sypyD5yh/+WUmYczAUp9Ilw63ul2foAahIAqxWWNlG860q1IJCvcDi+ST5/TvxcuzPir
qt27wGW80Ur84JcU1ohvXeBLj7wUxE4SSH0YZIS2OeLGptmd6Woii1yPHSWWyQ1+Ft89TS1widIq
H1t42s9uzhJY1plY6gOnouoeVY/HgJ0sHwZ1i2numW+xMch6UwmDiXp8dwMiFGXeLkpf+aUcxl/0
aHi8WAt/n7fsTWRxTjLjE51dpURKKgH5KBYzwqhNIMBUM1wF3Rsseod5Q0mhbJbXnP67R0Jkif34
PZ2eMroK4H3XhZVpvMW0ltOeCzoqMLX3av1oKi1yZyuuqfsRv1Myvl36c6keRzMrkSdMfXjqu+ah
9jYFMvijOoa4kA3J7zOzWOo3J/HG8sFjlPRxopCRckWlkuSjC+tP31TxU2jhtpFNoQ/aZxtE0WOn
FFevCk5vzh+69ZpgjFS8XEaJo87wUh4Zz+pDgkfQSmiiKp2YT7HvupydZHlCZocqvqESJ0lKD4Zv
r061ZrD0YijeEAaLwM3Q/8xQiZaxd2uE7254dGGnyDbxlI3RZHEyjaIYavC+IJC+26YcGfwma2o2
cGY3nsnghDQky3eF5HRZhI2sAvVagkBu5sfPvyaC+/qQzE8gm7BPn/4OnAzRxPkAuI342UobN2Cz
xtTVkIiYGnxtaPKrdrJ4eNIjC62nIhZrieeJLt8T/l3sa5mjAa5fmO1rc5tvaWWE+LfKmq9DN/1w
RbnhzHiwhm0E6coOBzsbDQNEeM18PHcUrBVVrm0XgdhT2KqLxqoefcn+FtkTqozQt5WaBTsYDp1q
7BGnz8tMJsH1q4t4ehOjLaZ2+vhHXlcIHqA+9lYJPRHFKDJPZHQaSuex8KrWpGO0F32Z0N6EqjJt
46H6JuinwMFEu5moKqAL9KV606NLLDkql1x0yjHCmaWvcd+CiHqJ95ncL/mryXnyjjeM7Ofexi0/
YXUFdv2EZarhTgkPMC2xXrroPVQLh8zGZyt6VBkGeMg3UGHlx/tdR77q+28IskfB5G/MTF2LTmqq
P7SBn3HNc2lL7gKxaFGvHdrePTFRwBow2A1FMbcDp6NzEWaqMdw5mAaUC8r7NoFvi5+QLhUKUVyx
UoSo0KZwMe3Th3b4293ETo9pLMGQJx6R9pscGbWwNsnuBz2yKFWvYH8Z558NaE0uyLygbcneZ7WV
rbtSGm80bNoT7jRvtiL1X1O0YY61IJd+h0e7/ChknpCD4wCL+ZIzodkJZS9KO8sWWMeidwm7ULqU
3IYE9/3yd6gQmYvj4im9mWe2RsG3oUHcRyUGfugeArALMuaETSJCgUGbwFA9q3AR42qW0K1xNfdr
qVZt8SDxpe46vaiuG0fiLYMWGZsWBRzbGBMPDpntXXP0mwK4hwdkr5+5XWLHYNR4exFPWyow/jq6
REOhi/JmxF9cDscqRc3RbfkprOUxTSMxePeyw/fUS2Wm1fFEq1Dn7vkZUFFYLPxhTnlxN2R7jpdR
oFO06xy72qS7Sv+X/HqXaoTZJD6HUBxnvUVOF1sEI0STtpSh/n/Bm3II0x2ppyO7ZAM5zFxUEvqr
OI5R6koGV/N+Wolgzzs6zICQCsT8rUbnHvQGH+5tiHJeLblhFWJiSWnzquBEhJMLTMhbE1NdwfVT
nXgmbG/lNVSZOzuMIvLJbXnFZVjy6bObJOgra6wwSQaUEkJZ+DcVN6GOS4snnW5AVnoqb0HzP9uu
bFkX7AyZX5ce/nBbT3qCXDfniHSFQWD+TjIDeFqk8UMbeZFEzJG5eQY30IFQCZjWlzPrqkQhJRZo
psV5UOQW7J+1jhp4H6AopDkT9VCo1IttsXWm75kzyw4ebAiC/2yeK/23ZZnzanl+/CHfh7T7Hd57
o2OgMlKBL1ZA+KSi3yIZEp1DqvsLLn42gjs4bJjM/dc/eLEUSFmJa1LCoEHSUwYF2acLrmhctvUR
mO60RQoZD7W3a5vdCZ5We6kZSpilslqhhjq2KThgc+UzJnokYP2cDMWKDmDpXDpa10XIbEng4NiG
WdWggj82bDjJY+bO78DCUU68zQXRal/XHRn2Wj3PxNVHV2ibrBUXJXb1TXAd3hHdPBqH5o/2FWEJ
pdC0QAJPnPIFTVrsmwQslYC4WoPyDZeGx8hebuXDKAFznGhxEmQ6UlJ6Aal6qq0Ixh40s3MYFtls
xCNWbGJZijqoMEphlSgTlYOgpHvsBOmuhYw2l85Xa56sTDJvBiPuOSYL4vPQ5uJ49ddEllfPk6EC
+VUWDdXlUYmXEAZDf0ACVRodvOQgn564gqs/MQmB+vJP3uyhHSAatjnMZlpuD7t0AVxQIMvlOFBU
k9DQ6I2VW6WEkf2qIe64kyvz1iW2IuFd6bnPNIH30lNTzp8hSxXkawMswffeQ8Z7wZGENxtKdbRo
FPD7vIyuZUdUiEb4BmA2Rz2yYQVVZHRWX+/eLYHZ6z7Szes+p/HLq/JLjNi0j5PwIusPsfmX4Jbn
MWjf6AJVp5fpST3Aa2undfoODYjeda+3EThWRuSipyIaf6xd5tUbwGbr3r5dXmf3J6ppWVzgTlny
M4uVxm/ztRHrfROQzsssm06EOtDIXiG4wPkf3Tl/+6VAaKNZrrbwE67KC2KKrv4sXHUeC38RbHgM
tAB7OLecPbXLY2OIbrCqGK57nW70fVV4Q8m+PgAAi8yOYLGvSHjzLEs2SIfwWY6UQxgne3KHkDW2
dKcIPIdWlq/SU2IdYmfOeVTk+x5JsoNFz9cO5eJ8J7CUILrUT/59Kcl2gxA12pmfqldt0wTjvJBu
0TGCAWSd9H6YdyU/8frjDbhZXgNK54U6mUcA0imxTmtqAj8GA0hBv7UuGjGUt/yBDhZHr2MeGR4g
kuI0pyYmefOxMwjkbhyHRm4aWDMXhMhUlRfkL4SouxDVdqwAfa/n9HGJV4dnqqTTc41cETNl7M9W
huOrz2hjGupaxsko8XGeyZnNg0VIbG/OcetHnDGsPIXjlvRJ9is00TBWkEzDdMVvlCD6lDdsW5JC
bvrsfJ3FV6POPqf4sCmGpxI1zcxcQbUEWbYItTPcxHsMibQKwGNbBJhQeg0H8AJ/2UAvPuVIUn0T
ZMhsi4rdy5wI+ahnRfrq2rA+g7UudcfeUoNYR8oxMm6M2YlyRxYIHd4AuBYhd/Fa1p6OBVC4wKrc
tmZVRFNrqOwHZpkEWx8GKVxk+EyvbBA3Eu+0s1hZxmEqQV+t/m6KNKuxwRFGSFjqiZPkyxEDIoIi
9HSIOPKazJD6aTDh9LuFcE70jJu5C0kwU3NvoSMHRREm8VbtKn8augjObpcvUgmktyX1GVxEAZTU
7qBjad1Yqj/MEQjDJz09JROz4ypyvsPmyCGz7KlDOwJ5Xw0IaugQN3ZQgSoeVNBeSIPiQLsf4cPq
F/oDHTWRtFg+ITDiAOP1x8iXP0riJRzYn3rQFXn/NXO8HC9iP3PuReGq+bSI6KxHIgIyzBp/v8m0
RExdpPlU1Dteqd/ZvMc09+ye+1MJkPBZe+QI3YZlZW8qmWVetaGENmgxxOGDzUBP8HAjy9kXHMzL
T/MzS8mQlUsfQ4qqUkYYlVlbDEuOROS6A94Nsanuv4qbs8PLk0EFMQP4Br1/WCahUE/19hITJliJ
nmGbTJLRA/3T/ovIA2Fe+ec4EWFHIPMqqVLixcspwqHY9GVRLQosKwbkv0eRQ9bzfJEpKFHGKt3U
ao8+cXCiQDlRG5CyvAdJPom3AVyTnuBt3SfX3aC9PDyqo2tD74gdE5Wk+inEc6foFJZRBugLH7Z/
oNWG8j45grXL2md+ByTocmuqt2ycKAKV1Pn6gsZdcGyilSBGo5bMTSOFOScAs1yBtF0qHNzC4dlg
8bDG7CWtmZrs+IipTar3IF6hO2wAKT2WpGOmlRSfBP6uxliMYd+tkK9xadW1LjDfoFrMMEXSMRrO
r8wl3evlL3DNLcBnYEW08kEFp0OHdEYZEdMgfQF9tD4JIzVk57mJ260iSHrWd+uGyk91qExVg5+R
1TXR/mtJw/NWKELRlNbrQnLxWCSF+vHQ6SaDgLuFDExHNz7mmWg+66kTgjet49+sLp7aGKMnk1Tt
04yIa8B5URy/UFK+ck7Lb81lGfrVtbLEtjEvusoEEIYD4JTiQt4w7uqNllg6NMlf6U0N+rXcjQuS
2Wt4pZ8ADi/9LVfB8mJMJDKhXauiuC4HTDVSQbQDAeiqRDxsXr49hxCh8TWskXn6REFtVqZSRdsw
ScMyXLUYPDES0E80ClCvd5eMZGmsKMbAXWWXy2AwvAJtLzWTLdA1p5UnRi4aLf7SphE3RfeHyDHe
4TzYw6NVN7vHQ5APyl2yNpzaxHkLevetwX0d22mDDr80pMhpwyG/J2PHCmtzQYBoMqYhPY3Kvixn
Rjnfc0XhfIddcn/MO5mri+tVWwG1i+AC8T1FwZgOXMdlvc4wd476OnT9Sct67/CrLW0BreVCGGWt
VvZe75PhaAdeMTymMr1GFGoeYLhHtDspqEOZPF/7BFirmGm+hzHSMPUrqYIrsdX+reXQ+AOoHJTU
qxFetK9oGtEW8cSpT85rF9Z2AfYjRyLyiOlJwkapGPfwkkSer3aYFuaJcGOwcuFN/OxfdmabAFiM
PSTin9lXojvB0RGWiTnwwTn/9pOR/0Qs7/VSXLiCvpvo0eabddWgKz55iDcjgVNlAbs15YBfcwvc
use4V9d1gcs+1g+3+vNswSRaCmH0mG5QF7kZfsArQqH5wPqC4bBX68ee1IVggvd5YZ0G1ML4Rtnx
wSvK+UlLiBNoSU3jKna48Ah69ru8rA+3/vfatsNXFa/enTCPuS/RxEZqxbY21L6noA4rxlK4+gR2
m+Ru9+s7xYPkKdqsLAYSybzt78JRKRmvbScsSbcq2vf+dlYSxmy2NJKi6pa6dKikWTGZ194oFY29
HdNb2r8N/YaRI+sPGmuGaoTWxxhwV1K0Ty/gaSjrKR0hq16coxdnUVo4LpsfXUlMlX9Z6VjcG+vN
5uv7lzPgqaYKNtPzKh2/U6laRx5gz/Hf7KzzZDkMX6wGT890Dl7t9H30qQeXekFomxYZr3i+Y3XS
ZV6wRjI3OA3gNWuJjP+1KXi+ETF1t4Zp3dlHiI3wnJDzZKyT9qavcwpcNGoYfAJJUMjOErtZpHp9
yZnTPUJG3KMXRZUq8aolF720RrxZYCLmatk1c6WF2P2EG0BTDnKcPZmrWl+E0URHd4YUGftNorl/
mTLUxPazgwkLdGQ5XDWq9X1eoQqZJgmsZUSrzsc4DD6ch8YaeZ5uOwIX6ScPLgTisLTV0w2dPfXp
LqNmTxqEl9s46ItsdC6U9FHC/nPhuwE9xI1Ulj5hamgNIO6TmnhZkz5wpgE9OwuaCjFWBndb81tV
ubjE5GNMBsDjjFJaormerSfe+4vSzHgVWLu98HxFlmW3FAlDU6HWUa1EEe0VS4rnDv9hT+AIb2+K
ffju5IWhUUF+CT8ekUjPZ121L3VekTI+kK5u/ZMDgRPvZUOfRQvFj/a7UPkQUs0+VpsBDjVCjwfV
bZyEhJ5RucGDmHHwAu/Wvkf8YhX7qAxPm5r8dcdSCDZnjoNMpCbzkLUCOzODEqIYgcqwnc9q3+yL
qxBbxrPdjQSbsZgETMnQOZaf0lx8NK6JGcM8vxX0eKXA8hFanI7TA661LLKb+hh4VD+s4+a2c7C1
ZVfnSeKPQ3EqY+qBit6MjN9MFyT6X/WXfFLqhvy9PCI9+myMcImdd5nwoKQbk4aK3JRd7KKUE3aq
tSUXSQxVhOc3m62MMeJSmZU4KiaY9FyHeMOP97I4Ms/09xQMqGYiZjjze35D2EqUZE85ktAfWcaT
KXzGeAPqi57EU7Y02rqqkUzHM9y66xCPPGRFo1NOz0mMMKEqAIEjgyuuPNt1To0u+2/LcmcrVSzs
S4P4Tp2yTaHO43UuY8PDd5wzJxX5rTEKW2s+LXvr5QzLF/aumsEGzi4+FXnIOijmI24y2kCCYW0h
WScleAHmcjdnDrY0zIqTDn87klMgFzY1L7XsThxi5Qogb5lonpRrr9NxpjiMUpNvYQbJb28qIXYv
jmNxnIUj5h5xxsvMXrL9FYuTPqVF3fuHtEw2qp+/+B4TBopzVvzyUmDFtUYAjnmASJEO60uKmeIF
lboOMWpMLqb+PvKslxJbiWxWEoFAdGNfHf+jMnfsiYPcAiz7ByXul5HXbAafGL0R0twQfxxV9uDO
kQH5AOzYz4gITng0JllQ7hNm9b6XB1DHdXslUzjqS0XN8F33Yx8zmOPnfy+HN0uU6AyQwGQPUIO1
XCkrHmUmQtBui37vXCUk2vs0ZHuCCUtwtcB7/lvlM10lOpGZI3BuEoIeeHGyJjpWktqxHUSuG66R
4iJxA6qbxi1LkKIelYIqXQX60RFrvqftHuKZlSzpOlv6OzIyH6w/KnCgqwEfIXpibvhfP7QmWC+P
tBTptfJnStbSN2nbF7yBQDjQZKAszk3yT5Rb3VEOBbKAGvX07nzJmO1cNIdUpp281rYJHtxxJ6/U
iib82cDc1Q1JfFQnZBXvv12KUWZML82nJU+Kmj7G82HOtvxdR7UyF7aWq4krFYr4m/cdmxQ/YEbZ
pEjYy7TNSU1+npg5y4HtZ3SMGd2d+mOMlkX4I5YK28eCaWnGl7zl0aKsa1nHIMuFP4leAq7VmYJB
ZRH5d6FIRW9HSO2gUkuxMBqHBQ2ipBQHXzy8rNC+FBamoeyIa0UWnGkmXNVgik6Shr+NGl6FoD7e
v5KSFZkB/j/uwg+rBlGLOJvNHLSJKwAqlF6coKCtIfs741nV2/C/D7wASnexWhGjwst3uad4sIo9
4dSCgL5zgeKjNYRCJ3dCoSGMRRTfNx5FJcZS7cS3vSxjqVBzbu9FnOVVCB0/SfcRfr88Ftcb2VFG
aJbfiWrxPyhIxchWC9gZRw7cjMw7Vuq2i0HamZS1HNn6r4TWWqSWgjzz4EgwKBSfw6CAvsbmrI6T
/Twgc8LD5p4ncQMge6wt51UqWIn1eOvzQ+74Y6UZCx/tWIIci1HI/ATsNk9BTGeKHxY73ZaBit+J
68zp74Aahd5dNb5+N+xJo3GQqtm3AQLsCFiDs4VPy4UfUE5tx49O009DiUB5j950Mq3K69yW3Kc6
xd39e0eyk9IGyn9stXtbjeukDAEyxoKGCuIMKDRAtCnUzAvQ2gh34Xdf+LjL3CG5QU6LrOB1tkXE
+eg4r+KOrDFQJIHqMJ0tdyR4m3wZIcmoJK+rt93Imv8XhrA+wwGwcGJHFcxp07jUjaPSxpv4LLPi
xgRVWTgI7uK86vx0LgyFgAbSt0vM15qE1qOf6MQbxfPVIhoVcpo/neyHw7v4VE2jrK3gUupzC5WU
Z22aXwush7tkn5x1rH5Y8xdUV7iSAO0XVmqpVe3beDt/jv1xazENe+Rng1aadGKSdCoh6LoPSlNq
s2CROD7c2RH32g64bPHl7UqWmC7YrMQmdulrUrFuUqVdCxqXiFjViIkWx1ArL9gBMsaI2U+2zrwZ
JhOyzXB0uCA8D7k7r84aQLaGpyUPowGpt407q6KYsII3W8m+m6l7EWDRCTvfypbFv5FVfX3XEkTP
27kmr4wzlHEyl6hwr3nfJnqgTmGAkvY7dlnO4xny83ckoCgpCLX7gatTBzLBK0CpWnYwnk8ArejJ
Ks200Qh7RVu6u5eNnrOycRfIvJq7DINGylkPC/f3A06TtLj/1CEvaxbOhWqm5CTFJcSZyxHJQdUo
E7SsNWbMyTjYnxkojOBVANMS7VFtLBQnN/ZAM8IPjexyDQLMWAdvSbT19SgKXGY+CqVIS1fEqpEf
7KWAWUT9IYAU+hY8Q/JNbF8QSJw+ImnPDilyeBOR43/xncwoQ61lGRFhi3apD501h2plNlu0KIte
a1qITFWZTZAraPT/k/gX9r1jv4uGCsm5wn6FE0FokZcgnyowJ/hdCqxWQUrSRl9loiYg7eHlvv6d
djd0pdCYwxrKPfb+KImqL5UOSRpFVG26AtF8yO+fael+aah9WPtyXqzbwVkkXM6Afr2uw/3kxyAF
Q6sOerxre2aOPTVbzk4vjL10MB3oBfB2z+0umO2LGnxHcBqSydXXjr516HA38IDZ8FnUguudv6dT
LRJnoUl/Z16Jd/N4b8MT0K7oGNodOAeH7t0cZfOWJ06faLxpZRIDmTTyFtEHbUs+aPqYDi9uiLJ5
OPh4ZtYh66eW/7GJAHM0sZdHBCpDep+clZv8Hl5ITMIECvh+LzIIJTuFrOQUag5k4s1gtf71ZZyt
U0bQSjuTQGV65C94rwtPLcGFkBG3BKgJjj/NeSbqz4vsYn72/HIOIZTYMaCSu/wv5ggyAN6k7cZo
fEfWXtInjGYAIampksF5HokSZ6n6iie9BK9IF/2OSyBaPD6WlIaBJeLvkdUdZVIi381NbvW25cAJ
LhdOmcEZiEFA7eWNnLQGanjAyCxwguvwQqJLBHSBMgCwZDmEcPMGsGKHrbvq1aMisZF9CWo6H6Fw
A4cNQwgaladpE9E2ir5/Pm/x0eNTybYIruPYwdmVe8zL6WrsKPCzddkJsh2B73AexwJkjeYgyz9g
kfcylkBZxJDcfzGVotKwzsOe/e5TLigRkbZv4YPIEaAni6cn9jGdJXHPXnGVvw0uzi9cSw2yQ7KY
R7YRRIks8F9cFK6bE2/cYQh7L/LZjPkuus3KjhhoQ+cFaINrL+el2QbP0dvCrdT+p1Azu4BP9/NS
HQN5cBp+xpZFnwDiDnyAC+qMQOnM4F29X69CAu3ooQzDKVAKtfMSmDjVRVFMx/eJc65P22MOz/hB
ohZ4PZzBEXhn1m88x+nDYhPmfnGy4aM34yIMvA1NewlPeGyFT1dZSP1VG9eG/JvjjJi7PcBJ2D+H
lbZkwOOJY2cbdd7GtY0GEMuY16EK7aLh9c3qTbbfcuQP2TC7gIB8JXWCVCr19wxMPzG5UXvOWT7z
U92wCxfU1cl2egVITDy1NlRD0+5lqyOncB+EzvK3CGGrrO4cm+F9rTV2j2ObZ3YizrA2Ttc/JAIU
50VjjcKQ04Lgdvbx4ippaZXdo2d6ptmQHHzqR7YR9FV+F8WiH3dxyc5b/zixKTkJKSo6+mc7mwdH
GJHv5VcWnFD4ZDDI0SsasOy/l5GVhmEeZuU45AI1Ux4hMm2q+gynJ7JpiJl6bp49T8cJmaUdNrRC
9EN44MAYgnFADu7P12KsDGF3mgeq4cidghJOkFqMPcwmw9llP0iqmum5bWVWn0RMPid7arQKPMaq
PIyPRz42QcNM5OFphQ0aYdiZCtZL58HwZ+Dz+h2WJQJwOlNOxyr1SdI7x1E3YMJSPlaLJeGjo+Cc
omyC2VI0Y07tYObIIqaq2hOZyfq+z3LwlRKNEut7TPNQBuNAOhQlonre/M9QheTtavcQPwYkIHdO
yBe29HZ7436rilifcM9ghvQXq2C1l15rFGg40c2bNNKdbzWu/Or94yM/eyp5AiFdw03u7+MDPCGA
2mjClGtbmBhLsiogAHG1xW0icehw+lSKEVajgsvW72AcVPBWBDr6teyrf8E9cC/MAcgqclOF1tbH
jEeo/3KDW6W+odIZUe1yF1YBBwniqFkoe8fWv8/9kKj9mIkqu8+K3lHPhsusWrHBR0js42eH68Bq
f//vcHvOB1WQLT3oozE9MMGfcH5YC29EZT+ODOqszFa0f3E17JTCGEGyHOuRVppkfZjdZj0dUivI
nMh35BRDEM5xQmDqpylUa6zz1MPqPNO2p3z1nC2zTs05sTYAuOk64MVqKowFWBX5W/+CRS/MzZtk
S5omdk9Fy5WHv2AZ9Ua4W7qDWFKEYen1VkcXmlQXU0Z5Z1yU4gTFReeklzuvC6lodiVPY06X5HAG
bKc6QO/sZFNiD41PmaYjAd/4ka8pYhRQVSHbJ1DLqzapaExaG3pI37IpE6kq42N+s2q6NZBDE4i4
7SYmPKAz4uN8qaAWtPxq8GdkUxUWOBMmSh1Vv0Q5gRrdYwH6TFSdyTkP+6Przq/bd6VB4AIVU3eC
VtWNCSA0Mq6l6FwDUWPr+de6Gj/DX/JTy5RVj+zrClKHT4L6VwiNSc5hXlJxpppUyhZozgd3qY6V
LTNHRZ4sAsK6kkRCnPlstL8MmpCRsmyM73Mw7JEuuGb3OeY3Sn0qqas1OpM/I8L+3r9vLZNcER+a
lAVbJfFMep4KpiXWEgXbl0MLbPtjgH4Z4eDCtWKsj+xGyamK/d/MA3SfQxNcBb8OXIOQVoySf+Q8
voHYyEYPdhN5mJsa49sWmECqpIUPgofnOf0OpM9bulgOXMprtIzy54SeblAtumCYm6tRFyZeLwbh
QtozROC/hJ0WE8MoOhFLMh22nHWVK4oecdwYG8ovnw5f0dReoZgMWLKvtNxjpKYzgj5Y8UFaQokh
OpXdn51yIjBwFI3eZhFmeCX37O2p436FFIwo7MF40tIWXsr/R0Gft8qie+1TYYu0DVmmcEFgaPfg
u9YLPAdh/rY6U8n3QSHaGikGQzIqxH/XpSPlkdVwMRhNrPd0SICNvyLO0TbALXb+8u4fIJsWrDnN
B8jCHTFR+EaIQf0F2l0LtXNKhyQuHNxBgPSaChqUW3GI4uuwqeWywYpbsyo3lvT9N0N9PEk/2nSr
U2jOI+49ZtKeXsICxnQuKz1ZxPn1HjSBpRA5mPHObtTpuLYgoHWT8hW7XTjEG07s6iRzeZPEK58G
m3QxA3QMfilqrjc6vCEKTgL+oPTSVmyeAVfI7uJlgPz/jPvJ7SvIfx26/wOvMPvMMq5AxfWO5Os1
9wZUAh/aOQXrHiG+PZY6BIFzurF69G+qDeSNzZ+5WIAtVG2OCh/4JMyNjR6ti9NeAAqhVD2avKl/
tsBsffX9EloMvdS4r8A/CwM6ayCijvllSmvRBtGIE99Vk09JTE9J28FQRIfbbhJsvuBLFJ5CYj+W
oMwAs0KpEXELok75tDu08wVORDEIyRCgUyGgFW8kM46DwlaqXhdC1l0V7qZo//R+C7mhSKIizCmN
uwcHJYIC1O9S9xAGrOvTTJFRG6emvwKKAgdT6E/2oFWM7QyEU57MdNPitPX/t4wUdSrtVmd8jhrU
FAzxWTpPAOYtA8qUUxgJ82QBXLz7/ndRlJDipa2SnWbg5kqP6/pykVA7ootPdjnszStXpJC4mjgk
6C7Wg/dCX+tPEJRLvc/0zmcCsAYZUccSr7wasCGrDcS8tVgDjZzcrg8K9DrX633fATY0ezSzJ7YJ
0Ax9218sHK+fZmHVSJxBiBN5Bv8Lg/KGzgCGhRjtjallaNVyJVCQyVUzCrcXLUuo6bzlLcFN6PBg
QoBaE/u+C0MlXmi0W1/0yAL7ehJKzfyrWeArFZ/4qEiFz/u3lujGS9KRFb6VlyzMtnZxRQzzF+fJ
v0kWDWSkOVWWAeZWOVT9A4rHmhyWQ8J5ZFCLP7Y4criTHbB+tgg0Z2sL22+XCIAPNgPPS4Ac4Hpi
6l8cp+g7WOUAzz6CAkSkM9d4dUXpXS/ycDVY59LtURSPS8Cqq4+azyDp/3dLSGslnvD9rvRw0oJZ
+kJtRRhRYNa0ULGC3FiJZZ1UmUGL4MCIc31ZL34Hyn+bUsO4CLvb2Mj/dxYhWE2lbNi/LvotNTbm
8cBROX7L7vY7Fzpd1Mum3jxcmkzdxqNVhFcke5HjI/tSZN2wSQb5zF2kAFJCclRJIV9/ExuJ6bXA
6h10/GaBhW+zhVwhtJSNI7uMa/pW/1/MnRj61WvesW9CWYga/cPYhwAfHgNVnvBc6swPT9iU+Rfu
EgB1CUQZsf4ZOO1Zlwpaow4H8qG5mQ2JYimON5dmkyDVY9vO5tk+iW34vZAdUptnqnpu68IS2KTu
OZ4aiRnF6pknwl5YEr2cOz3cU/XV7c932G+2K4cejrBb+TxFauj+biwnyH9rTL/rTZsf/j/YPINW
bh01G/Z74gluIpahUq5RCfiFoVdP4quGcGuqRo8JHsnJGEsfhGpEABJhet5X0SybjyZzL1IOC1Mu
yC3z2hFUHyXy49Qao3TMOtRX0JFWyCC3umxabH5G1Fm5Lpdt+h4n87UgaNLQgKIQMZ81Vokqono0
HxDR3jJd3uUiNS+bB4XbSqSCu7qqeStButK+gxM8aTtXfiMgwPZU0vROlpmOWx24UivLf8gZ8FtB
+ZW7RQCYbD7B6F7ZiUEB5dbHATYkp7UmxjGkjgXxb/GyKxlG1/EZRR0Y3wKrssxF3DuJuL33kCpa
IgAIPmny4MliOG6wlUiPWrRyzIgxqOf3qkWMSMx/224GhjZ1U0gZBwB9lE1QvQjlzUzpkH/gHm+9
9JMvj+t8iG315bLHus2sO7M97DW6umZZ8apyJGlebH81DeU0NRYwWbxvJCDIRisKDUINgKenCWCC
P9ooX68kV/oiPpOBRmboS8S7zUMXKq15SOsEPyRdSmdjQyQ3prFWHlnA2PKTMTtrR8htMqZhWeU3
sGczjT4KQNWyTORqWaoR4B1Zsg9jqf0kMPFDMD5/Zfey8KE67Roquia7GCImspILV1cVvaKZeUTN
5N1fQVJYfpwpdU6aP6eRnMu5B5Edjr77O6gutDu5UsgSidHAg3OneNmDUXxXIimXZKTIEOjAxWaD
YCjHHT5Mk+Bnqr23+RkFRyksZUIGqogeNIlwdJU+si/VCLBEHA3zvyKd2EE3byTYOX69qLZOLCgN
k6nijfYDXOMpZIn7xkwYUwY5LyKdF3Gz666BP4TVq2m8bbJ/2fV4+MCdFcXcbiF55stmeZTwfSqz
qw7vcuttlQ4Cuh9DQY/I4c+X4ODC3fsRSUPuxxywL5j5tWwHUJHHIYovxL0R1M6SWnm28cOtQxUY
15Mrg+zOkPB5EB2PTiocaWvXbNQRp0KaftMfikx0j2oPWYAA0G9Do4jR0VhKDUdzyzj3qdDHZLyq
RvPioxEnJHHSoBOPhl8QxL2/62FMyKhl1OTXTjTuH0+CSKIdd1u+/PpbnoW7dJlGr3ttuylKPxjW
00LSr3K10mpIFMkkVqZteuzdzTaO0mvdPxM8oxHqgMWG0+S4zBUmovfHWZYjja9YerEnvIEYWCTx
tCqHpHkDA0meB+zE5sKAwxqKle8taTmMLyWEm2JGGthK8f23bqQbwQw62WCRV+AlqnWYT3fWlBn1
lUktuOtaJYxG9TC1H6CCbwcINBl8TrmJ6nSkJcud3ZQ8viVgt1sywUXEacNY8+5Iau3Rib2pKKob
/C3tKwOwrpZxeQEt2hJYHKADYkfvTVJawFQAz/alQqCrJMOEOHq4HS8w6XUSzkWAzION+Asx0VUE
3FAw7odu27yr7PC6C8lKWZFxlliJgRI8GAJ4OTHqaKTub766eAfL9CDyS7zI9tGVmOG3cEH9zc3S
YMhynOvLXabcHNZvR1rGkIwtpCxmAKhxpihniXqqWPdTmENB38etaIBEo/qpeTZxV4NnsYOUnMmu
e9pMaWj8c7eyXlWrrf/BVvxJevAKtAbNgxgvKwqoDk587vBoLMUxsPvALMh0H9R4KHMftXqWenZx
m1x3nARRqOXTTNS9atVtlh4CxcJAjWnyNO6104SgRm/DfkEeur8J4cHaiRKX4I/xkU1O37vGMAGN
LqU9Fm/DiQ5u869qvjWEMwwgtdkPT7Q98BErmIjZWNsTA0snwyvqPBHSs5lJ8jyBz4dmUcbM6QcZ
LFe0Vku/vkG+p4QtS0ULgmkQbWGrp/PXpx31peAofq22bVKEht7DCcDy2oZWqjOBmPVaJ6d9BYXD
9cNoXOYbnhaSvJ3It9gJt2CGKlKg0LrFTxsgH8AaMHY6QHI1tZuK/Pq5I1UzgjZhhWIj0zGAmJap
kfBW6MaQZAQaK6lARvtglpxTTF7HBLQsirtdORPw/mlEcBae4DCgtXTW4o+SJSfSR+U5fF40b88Y
iN+ESljMt2lcHIEtwqPqnzADqd5ZFsrJyOvE1qVID2EOgQoFujdvDP9Ya95OX4CAWGxUKWd8MeeY
N+5UYc6sslqSkLEKPPPW8LrHTBH9GxKT/F6EcyM1jH+y66ReTFhNmi3iJ+bm2be8ZBTAjbpnHbOX
dagSL96BfaekhFmJouIyRZPkWfhhIFoEKNiQVVbnrNh0PrpLeyQut9vjGUbxUuPeMEdWWRz/BeYx
o6oatJ6bZakUai3AB3JW5aCOwd60Tr4qVxeXZC0qVhuYtTuaWWtjd+cOrLEo9fxwym4EOBVBkN4J
S13HH22lXLRaDF6CFC5phRt1ktJ1iQ4/yneFL6EkgEvrSocFc/BBpi7I7Ewt0DfOxrPFb3boHDtu
4jUwBC1Klv/zprkXc1PjNo6bkBqgGL90EUGO1FtePXk01LgCsVRbJIRbKgVGJtctRmIKrHDX7w4H
RyBNIHP8p5SmPh1Io0t3O9q9LZIfmqh+e68ICGZsBp5N+xfVdu95GY7V5mpnxx57Nxo2p8AUl/pT
CilzvUVyo0gS0pE65aBWTPKhatcQIS7/QqLU2VouK+WkRwUeR6Z9WAd6ZH+jmTfguYp8F7Fzj4st
4xhn3N9d+w/5SejYc7OQCdhn8pEiVZCxRRcTriICw9iTing7aYVIY23L35p4HJQ7j5qDH8X48Wjy
c0j8NYgVApDissK9Hzk2gD1jHjnaWsA+cjvxVO/+yxANPuzW9zDTdXYm8t0QCgtDFm9dmvEbrXqa
npqI2TeiT3vTwrjlk+JZYkOv9vg515SwOB/au92ucVx15eh+y/hZMUw176D7e8MaQoAdJt2WNtHX
tlra3teth5xhhb+y6bhrZsf0W829RnH7QztOYeWiNsgt/ogveijq2TS3cvhv/iajMIbEQbXNEg1y
c4x7drT8gz5gGo9y5hEwndc3VwLWSfPLb847/RluvToxCCLb+bVd2fZ5HHRQ+5FF6C2kNfdQ81eL
QZ1d2ZI606kDxIGxTe27maVFWjJx956cpeo+R6k9JyJp2qWuqVBlgwfAw/iwVRBIa5U4CqbxTgBB
poJJEUtf5OK6unUEx3o6y63+Ni7+XZ7KyXqwQzACxA7F+7625AbkpNgjc5axHTd9jy/yyq7gEhU7
dmMIt/h3mD7lMHwjhb9ccfYPgZLBlotNkQdZOXTfy615n89+dj0eN4coMdNqmKqIkb1ZBoNzEmVs
F4Q+JHH7PVDfuxwNUIXvXL3UV4LOBbBaHXGWYPpbJoiS/bawBghcuuVT5ej3Q5++brInC2XPUThA
7elpC21v0fQIGBl+h3Wi/H8ZRpPUjDIn5C1jnJKM3Lie/VzKADW8j8m6/8w+lHvvQRbW5a0p+9tx
xBTolLFKs6C+K7XzR+JazWOJSyn7mr5c7suG1pZ+6ekWQcWjVfKkZZwg9q9CjBbY0p2A06QP9PUb
qNlk9UFr0EeZ/XpYr/tskSrFce6LjqEVySxE7W5uRFWiHw3PPNNnHz1wv7cDC3SOKE6/K4m/UV7+
IyrnR4nLlxFXO8uIqJsRCB12iocEYLWFFRqPhbw/oK+MhgNSFBETfTxun7+gGq+AssaM8HDaOTMs
ebVIS1FeSIGwathEUDUqxS4SmHoihu88ZHsVZ7u4vRTBxrKHn+t43MlhJfDTxeRgigWJFnuS44To
rmMofrv5mMAY8Hbb4VjWRkWg4Aanare4nBJZxB9sP41w97oyKQ69sEXYbutm6KXydy6/ZpuSsNE7
PpoTeE+2TlTWrgP81WFcsl4DebMaKUUmekVU5H2zJtG+LwmuJyAkGD6QUisrPDeddpdcHyttQgam
NR6JKgf3JUAAD9MjIk/rGlZgboAcHNzxy8UiYUznzqCvYbRuCXb9n1ke1L2QuhqScoTlAV/TZzV1
3Eu8karm3bUZxaj6FjWGUOMJfAJXo3HknA+vu4vqz+R/cXfMxARVliB93iFsTD42HfvtQVzmBQWF
v8DL+NEJW82fo94uDYDNWeTRzdw45GXOGCaznIedzVSNLxjN7IONFFekS0bpIXxsDwEG5vTApx+e
AQ5VadAg4znl3FPp8e/v6TxW49EHAIEeTyB7LxiyCE6WNnfv7akjBYTDQwtW8Z2ySEkoaZcKClsq
JmumQqZxpEdPcXfsce100U9Ivf7cGrLmiSL79PP7SzFTZ7WViye8Pf6fuVe2IeFTD5L+OMFEm/WT
UhX4xx/SMVoNw7HPHRSLfKZebbjBhUCDS+EWOIdGnd8yNmvPT3ChRjIBVJrWwfQ+qxjZCABWvEcs
ApyrAphP/ScQa3WWmJXz7OWrZzwK7NVUIBvsXhMGbqtBJ2RDPrC3VOtyuEWVUve4ftAB1Gk2ZHKi
6kGXCXZ1QFB5v7cH1uq5AnnD300Zshe2Z2N8VN/QIj926+LOa0OzSZ2S6mN+gJ2kcDnlX2OcXE+J
WVYUrPRA3RUB7cLmo5TSPpOpxKCmOwFMQrRwS8oZ4Qx3rN1fqGh84CFaXPT2XAUh0nQ450O5x+rL
SGAOr5iefGvLsDK1QOV78SebjBCB/xfVzwgO0qwrWB1X6J0dOeDVmX+dkTlXJdcrbi8kObREhOe/
a68OTBHV+m/G0NmWPaSNFIgxOO213i1y1WZwiY8S5egH9Tf1AgB+/aCdYeIFxlh+bIv46ikdsynf
PJHcM98AgwYIyeReJ1CLtwRyyKMPlXQT1AQAspJglmhq1/UHrr6f5F/hflgqpH51JKbTemzDN+17
bPzjVd/GlcshjlNNEm8ya9flnIVBZ5zYYl0Z6ddXv7xzVR38CZPwV+4ngqJg4OxvJj+wiqND3nkg
TFUbtvrm2aJYQLW7AqLl4ZJE8Zag/NeRonDULUjGZGUrdJrttHGZRE/2lPpmhltQ0yICnvUM/rbB
nzeZiijV/DfJZq94i6hFgGqKGHRd32v4EOSFhZMhzPpDP4ojQ3QZFrH7rSo9VM815NlvGH9c72KM
KAXV/8e0w9EZYdx9LzQKroNpFcYqUlzSKAuUXnFFNONVzxGYhsUC27dNUZc0q5W9Qe1fLwSFDOsD
8g+g5YIcQWOx9w9cqBpL+5F0WSLq1Kc1JzYIx+M4Pmhh11v1s42bRZAg7xxYcaqkXcd711LEEzfg
ZWo1WvXeK7bWGzy8JBE+VTu46A3sslbi0hJpCstVeCg9QrUyTtiMs6RWpzyxqcUOVjf8Na53ke6n
ko9c93RMv6qRa3yAKXV7T05E6mwKhG1bCkx/74uN7OFIjaG/yAdwq8xSwSyrCoTxgFoTK7dsJCrr
Ixo22IMoAXeyk4KvW4lGySn78HBsI0K6hopDs0uAVu71B9pD9pYPg8bCAFOwrFlXl3frAPwggXOb
6O4J0FOqevm37uudpGE7cfYAVY+lx/iOxeGwLXfQNpRg4tvz+AtBFsOi90FqFoFDaOG+57nPRIis
+iUVvcv10QGK8hYe9WlzeEXevo43ufyvE/bQ/K/pTomub007LIf97CMO7nlf9jGgDByS20y9nXOU
U45B6sZ7cJ3zgSLAUDFIwMRYBy/RgRPGADqb1RxErmYcyWZYKZGwB5+aki+tUWpGEf83gFKU+drG
C7wtptBxt3Mq/Yr0/485V3fwgwrbDTdhCfy/LRtVBl0UuEZrd+TH4b6IUGMQMBULSkmBu1NZ+YvQ
yDZ/UewNwcAn/rxhh3ZTvr8v+ZJKag1PVRBPNBKzYpMKS5EqWFoz46aBK+TGlJ3g2QGaZqxG5oVC
vSL3yrkY1tDhAwxS8mW9NX/GAPrp7oCcB+BaQpnsyA1sp1lIqEi+jqtahJIznrXnx9cRSVOerixW
hSDHnE4Lcfy6F/FZMfa/QVeZImOw7tC5gmH549kCRiw74NN6SAy8BztKu+7M5JWOeOZSVA6ESiSj
vLjuFB5hp3g987rYMfz2q9kc4VF3dMXhBB8hwemqLmDbOxaqBOxsBLB8a+Ti5tMOHcp/fWZ6Y0uv
+WWGbWEoBR2Q2YaeHJtDfkE0qXGzaM+/wF4nJ+mYNpwgyrKugFcI7GGlKBJf5AHss5r5y/Y4rC8k
U1KtkixdZmzfI0kyGgZjEfPL5VuWXXhjFpj6EM4pPYcTCsJ2fZJUBexvuFisUfudYWHnPdNfqQ6y
oBOAz+TsKH07BfxYeD0/gMmOWGpsDOm3fJJM8IQs9C0R8Vlf2XsSc7+1A3Xo6bUMMcw/d4UoCMH2
Gu8zlx+jldP3EslZGh8dPrAxHu9yAruvGNm33vYWPpVdaRVGiRaBdYt4mxGTyJsUO81U7ycn5kfW
8FERFBGChysTZI6OGgIjG9D44B3ofMeIil9++QPbsgeL1NPFzTth3XJdKH5rbfSFyi4ypU7E8a6N
DIMNgkvNQEKp7dSJKpINOUIAzzcOM3Wka0yibQiUAPQ8GjtIVVxuv/TaQSLyqDsKTBbOCXYCsQ+R
iZ1KZUBS4jVzROPo/g3K/CIKvGEUfTA6H894ENntwXhjtrPWgemH3EwVIfCO9Yr2lfcSdRir2dhK
AtsBOnxUfU4OOSXls8jGFMDrteB6Z1dQ0+35ZaExJP5s8kVjSgKnw4XCW8guJNu6phVOWTdg34rW
xR5EJ3xG2WZBnaM5Wa952TNokEFLYQtZ/JPfk21qsZfDMufdmK2V8rlmY4f83dnH952mOmr/oTKN
iSVRk/H9CbyJCqZw4lUHgD7ZK1/pn1zlA++Bq1F/AQcXufDvtmTXMv2aRvKqpRmdxtwFLpX4nL7G
fQt9GbrtMQ/3Q0vH87eRFQd7EQxaETmt4K0+O5IksfJ5VeiRPjAGeMEhV66J8oCzK4vhjUuTicv8
ZDlQcNfPBxSyk7r4l23AVCcXxqrpqsNAkp4Q+4EDqe+EPRG4bk166bjJ0h4YmghuJ/VswVMEg0PL
sNCW13px0yshi6sdU9oWzXvosOkC4xNWutuSkoljrUOdOoOdjLa3mXA5UE6Mnf71JKjBlbZ5/jW9
OVt78iUcDMl3TQyoz8ejzqW0bM9q5jV3j5jXJbtLfsazlqEcDhdFc5ZZL+4HjtkGtQ0hbD/fL7L1
3QlpvHaRE6tGONK7EF4FHfH33t1f2C2PTvCGVAB0rsTItVoKl4wDZNBUj5ZewMvKpf/jws7/noPn
DV+rKzohdLaallBC/Wn+jDOUqADs3nQSh6vbXKZNntwjMBP7183abq7HzE+e7zETEpxTkMU9mNkK
glass/kGgUWCdPosdZ/LaD7SsizhDu0K9SJDgNAax5Fn8XGkWGzoZnmBpDaogj7Qakq2Lbt671xZ
fmozDt8FdCyWhVaHZY4nk07Ka0O54BDGxbrf0XA92mG3LjQGZ+hGzfzPv/zDz+71T7cpc5V/M+gd
9FvLZSC+uKjAxmNNoea6TiFqSVduO44psSN4Rr5W9wqCmVqqzw+Dn7pgda4oWBy0JDDmfOUh7xgV
Zys/TyqWSF55M0aVRL0MqLcbTfX8FoP3oQmEuZYwSxzeOaxjI0eDkUVrNo99pTMqg3f6+fA2BCX+
ipbPMBnAuMuOSENF1xzW4My+rVahrh3zMO9S13g8xbPy9kHijdBef+b6fkI+UYPgSqKcyrBLR93T
L94jfM8lVksvJPj1o4cXMPnPvhTN+s1RH21wikKTGgohGwcpWoauws8MmuN66hVhWHEzctSgYp8e
P0KsxUJ9Hf1KhYccj9dCcLCePthzOlG0FibtXuJZ9xhDLC6uiERdEVqKdTB1pJOZxK32vsmtI7j8
1PmVHNEPWZNAYR87udjYWrMuqaX+uGOXfoK/5lJpn4MjAFM2Gtq/zgTgxk5CkriTwZMRzBjr3Bsi
8DkbZVGKLhq5Rdv5qEcnUykC1LNwtWF5iqAVLteumaFkw4FXmwQAofH93eECnAvDPpMekvWpuAyh
ZzbrVIzsPrG63ubtl4Qk1i7DoxdFwg0AuUIq/EU1C6YrA1gCDFjLHAMtuP2EBfP9aWfU7ggoF4eL
Kfx2gu9iK9sVvpSiA5dcYXefc6NkuVPmFTXMBR0VanBX8LWUGCUKCndGgFdNEyhwnOABpyj+7q1n
r6Jtm6JiqE0L+1WR51O4SGrEQjlUOa43YRzcjndJi0O+Iaqm9rJdwEqePIEcoLFptpqmQcsHKGDw
Ak3ry2MSnyFrNfRtpkCRpd+Y9lY7jMnOB5RnWkzDoErHN2IwBrDNuAN7YT1llqmgwwAEsCsx6+1V
TgDvr1Zans/AtFA+t7MqWqxpUdz0U/jK7dCUhjYLHUpPv9O8BJxZPXUGlRAs7+e6XdErAnkRKSyK
hwZRE1iD0NxkaVYpEsrlbsaRqgm/zzZNCLVMWVRI8XV0lCWDT44+Zq9L2EpForpSnqwNNAPpOlx4
A9mXk/sIT/EPWwD8w8iBeojbezRV7loK5WrveAgUJPQrs4iNvylkcmXTQQMNVRS5bb86YMpCovE0
hLU0dNhojtWdTbwt/dJvoTUVufqJnhJrmlAElODGmT4PgJeX7LnTtELGJW+bn6TM1O/Qlz1Jk5DE
BStCKRzxhA+Lwl7ceGsuyGvGEjJkeViI8bwJhHaTKKZRhbPnIYhYRGFmSx/zdiXYkf/FTbLGhrQ6
AKgJGcWbJ4ehNT+dE5+dqTSC6BdpsgyuAf9R3QvblIecFeo6efkigJCElnvRXEjb1izW/ygRupmr
rUE74OHHZnsIi21dafpkk1xomzTpsplv8/JNgaJ3LdyfQIw9V/IFHC6+UZ3HARVIDqfv2ZbqwSCx
IqpJ4c1ZFwSTVs/zw0Eltj/EOm/3ZVDGxbkTOkVUJVp03a7qYmupqruTh4sBoVt6AOL/Dvbmmr/S
kyIEdV6YnFRlqZKFNt5nzFsWZpFdy7VHgURhY8E20bjB/yltsSsw3bcSTMJKaRrBV5jyInAxzssS
Vqs5X4Pb3K+UVdm6wQ7XA5uxK9icRCuMd5TSuqB2ftY3L6A3zd4zEAfOL9FI+Le2TaBG1QylIwwT
DcjL6+hXlLI0RdimLYAa299odMqojBNk/6PIZYd9Fj/1N+DS6+MzzTdvSA14hUECvEllOVea/E5A
laNqdWpOsYDpZXErOFHabvXviz/wS8zun9cl1zjKtGJ+B1t7W8CEqMfpOPAyFKGcnOdiIr4JMDMf
JYdWBqIMKyJcJpisHH4et8QXaj8zOU470Zp/LrOORmCM1hOwtn9Zx5MT/n2PmgOx9IFNXWRVInh/
IOG8AAGdJJT5VILTloeBHdubTHhjlqJ5eSCUFLiRkt9JQyE5PEkUF48Z+UYLKkGSXK4Hg+/9qvoz
AI4Fcv8f81m3zEbNmexhXwBjK0xFQh/g7pHszxoueHZQujtgvNNnfCfUlJfmI5YuC5wgQoLsHHWv
pdzlNmW8FHyCYApknpSFfhpt3iBv6NDvUGABbVm76vnjSbKpkzjGjXtcNhl3ksZwl3VAkdRk8gxk
WKc/52IgEP2W/yk1QhvO5CRkrm6J1xJUnjeI04Yf6M4mSUjD2pb/UR7ewOncWQuw86K7QcLFH1+z
PmrZlZ9tB5AySW/6xRAEDUkF+tOaj4YSi+o9eR1MvteeuwkvCwOOJCi+ZuN6AoZEk7xAWIpG6hov
ZPF87lho+NjNSVrrQGrRrO6QuYJOoE9Xfk1r7PMp7pu9ZunLhV1L1SnwFEDe7nC6tsc72xYk04dF
vP1eyQjcupcbGQ7Hm9+xaW2K8djxpvjaNbczt4aFZn0oEzqBbcPpFbC+7chNDLNfvPlnzGQj3oio
UDwEQMUj2xWd3dszumT87pGk26CssHCg/HZgsCu1GcEEwr5WCgZ48oi8xjP47wUj2ehKpvyqEsxy
qLdkW1w0Ng0uMmtoMUS+0zP3BeotjObOTq9RgVLhRbDBlkBp/QrpbiiiDFlApvyYgXl6EJaX1jjR
x3+zk9yWlSNo1UPUmaRSM91usRJQiVwAMAN2L6BK9i3HzMx+fjvyOn2wtw7kgy8jrGSuiZEsRyZU
ssdrrNoXXRvHIDLj2FjyGAGQ9HaU612F4Ma2OvS2OkBn7LE31VJsU0DoHlTEkG91znMFmUzChfHU
ZEeQlR48v5d49gmfVwoe6a1dxh/RKMQ8CkgHFzHSHPUqFEtmjsbClqYQFsBds0k9xmKRoIWZ41KD
kx+fTflrCWuXDP4+1fqZ00Le+M4TjSCYi4rvwoj006jwuz1RA3mMJKypmDADyZTTLX4nEUupXEZV
92+52orR/NhQGIR6D87Ug76Lkj1Y8BchOPebm0mhVQzRBFcQ2v8oYeEIbS6qH7Acoa/YeAb/m5V+
l6ZrCEWuIrpghT+IdG/1dKxl5kk0DfgQUtL/G1hmGCe3PrSbOPpLzvJhrgJa0SCOLaufwOtc+yp1
Gh0ybu56/yi81sTjf4To5FrkkAVTmNQSg0S62wTaHmH1EpeRhlU3HErkXDD7WCYu8Oxv6hWs4ncK
q3DSnAClCBQJGprrs/YGP/D6uXsdZcSK6TEhcyD5ylGy3V780eDSydeXRSK9vQhHfCqdPlNkm66U
l1k51XundM08tMb7eZ1fwopxnYkuagm9L51JvWjOvWyEIeBu5SANhfGvN1yV5yP85aSaOqhs3Jhp
17u2K+oT/EA1czIy9EOL7i5w1M+SrkzZ8AHMRfmMZFj8WnpJUcfsYLAugg75asT6NpPjmf7dTrGp
8qI08epXTM0LeDjqdgDFtx8WMlHdtH1Rww7SCZtOphpld48aLEi7bemqJVVpaVklSYTslGFVWuGX
vkxKhfPXrRVD0PLjD7kT3Qd4TPWpxGB75mlIFa3EzecLvhR2zTzMPIFR8pNu81mmFTXCAOnwHkjX
/oQ2CQxGkETdlrsSriIROkbJyPTnCXexcLHlrIKOSnLOpwFcs70D74s1TAnl8iD+FVY/cET6vutK
FUTSXVOFw63mIv9pJz8nx+Mf+dz4cLIYjR4q7EjixwKmQHL/jDKBYMVJFQi271ejmsLgQseJVHyT
WlXm4w8cCfCXpiPz6232xqRbC+e6AkMmnpwtXYyut8nWKzASH2jm463v95Ho6/ARTtpyZ/YDSP2P
kDBBiME7InYDa9gbtuLItJF8nxZDfpmIXBSPVmxmgVSndZ5V5e9vooUtiqouxU/0svGjTW5uESP5
6vUro66p3w9cpqHNCXLNugLl
`protect end_protected
