`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
crsuNbGKr2+HGjsnrWAO3ApjaENLE5lmTkmDpqy6wXOqFQIJnrktoh4R9l/TVlY/BEwSOhFtvEbq
RKvf5np1ZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfoL36fNI5DjzIQX15YYPTK98uQI+Z0aMjl+hiAVWq0lzClrfpDjXWaPyQGiPvnYkkUnnCNmSyGP
qGrNm7GOsjezCGzMgQVr0792OKktWuV2kt0zVP1RUZuHk/37eznwh8N2o5rw+1YzW4dGzl1QbJom
tmB1UpBcp868gDBGaIo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nZKDyxkYA9uy2Xb3FwpEri9edMFM6SqsP4Aed0tRsVeeX445M1QANBu8GOl8sJ4QNxr6T3VU33/s
FK93SNbe96iXZq7rd0ZTftDGFn/wlb+m7r0WSjfp5pkNrLXaYMROFr5Y+cSF68dabG3s3COIhufS
z6LjxtxffkVZFl10/p5NYIyhVlCgj28/qTLowb5EYe1tZ0WPUAxBFuTyFKtX6X8Ha+x+nETiYK6i
PAhbV564AhzWOG1ohxDJJcn/sq1JfdeuDFdYSbNKycH1TqhYGY4rODz7EB10q4+UCVziUOr4Tv4R
NCotWnw5vu+fF2mIxu+vVyyYTSX+rhEfPs2iXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZ2XWhB75BM0Dt/9VMCHTjvBqUtECoyfIkFt8UyDN1IrerieLUkQavGMJnAyOgfgB2F9GkPnzVQV
7H9tsdZ87Y+A3ybRmsawN7gt2tqx/GGsvZlikuuSepi3sHN1vWxch8VpcI/SFn7CnlCh0jupM6VR
707+yLDj5AJkQVyH1LA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S4eCKuneguafnmn96ntdnponlGVTmyJu6zrxyF34ICbqsowM9Vhvgm6poU8XDQ/BrjS+RNPc37Fg
G4CZX64FNy0IB8M93ARmuOVvrGN2bYMf3jNRnVO/z1hOqr23u4iXXLcNjJcX+q+ntygTqDn+dkJa
tNf5JDJd7KcZbafDC5iOu1RcjafQnwlpqyaxuvNRdQkJM7f5tDyB/fmqWMaeSiYSf6cbwC2Jk6x0
7wUP2rAkEzcYQjkJqSGT74QQ9ZxpJuO1xNUbfsJDlmWbSmEyg55J46Q3XRBw9O4UV1TNB2XnSxvt
0rRnDIzS8sn75CDPR31VCmG8K+PwSCayofA3ZA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16704)
`protect data_block
HGwVbJA7sypyD5yh/+WUmYczAUp9Ilw63ul2foAahIAqxWWNlG860q1IJCvcDi+ST5/TvxcuzPir
qt27wGW80Ur84JcU1ohvXeBLj7wUxE5VLxV1phQs3c0mTb3oMLfKw1HyXAHZ0yl5xQ4h/F48khg8
PLSnPazC/6wIz4P/WoBZnWEF5ujNmFELOxP79CWZc8NOeyPVDjMv/REG1c7TWeyRUwS8rDvGpbru
yP2yQTGjbH0r7U/bgCVEvkq0UdJ2HFDL0jpj9l69g1rjc7eBZ1JBfhx+OKICLZnsgfplycjJ4V0P
+YWpokDIuIU9BwjNDOU5AjlQmpxDonl8EIbnyQ2X9X6XljlL++37lSnR1rF/qzeivZOdG1pEHV4A
/wGPNW33uMHw6vcLRLvQKLQ+FhMHvlw2rbI03kICmbIr3UwpXw0Po4M6G2VOv27mXnhuSSNtve8E
VZH5mC8mm/VnWYlObhxijNC91SRc47XUr5+odH0FxU14p9lpqKlV1W61IkWIUnIZUNU+J0EJv29S
3vZ8oTyhJZj9DDJRYDVibx8uTbWSRP8ZxhnuDDmg48oa0lAMjX+88gebjkl4gm+wIMw16LfaHMkG
k8f9lzxK1in+1+QTamG8zEBfV2anfvbgIFNwrG0mqstFgfQis3o0paxPNaEpfsg5uz6rDH+exExD
+28PFMVf38AdmMVyZSVNXwKgVZZdUs6mIBmdErkV24tb1qtou0TMRntKMEM1hAGh0i8tRrLEZdfq
DeDXSHWYbuU0+CxS8aUWiQ6cUFd7wTHtycvF+l4xrp+2SfkIHh+VoXKOTSEp/H8aik1EUgaNOhyR
ScdnGw1slfJpQrLeCBI0B6fPx+Dyh3JSmIn2gX/vCy9OySx8qz8QWCwhZQc/WMKraNsNIU+gmaaq
AlWMn93agg5VP2BG+YP8+Hy5WwY4QkvNld3hgHOgLdtjpLjN6oig0HBxhOgvgYclXMGm18YeDv+G
rf9L2YKjOUW9UzKS1cCqOAjCyvlR7Oh/Xxqj92SFqVhVJvizG26oAGWO49dXmYNGxWtQRJ5idMRI
5F7lSnWzMVb9/lg0hNysuA3ASdIo8ciMHv6mZ4k9j7Rfds1tpdPtmrw9bi8GH0PmgOUGYMTz4I0b
0qsGzUDWG5kmzMzzZU61YjWWXnd+UJF8Do0X0xtJ7PvVgjCPNqpuL9pdjmjFRlkVW/slWvJ/lPm/
N8i/hjAZqu7v/NonpihmatCUHNkyeH4e4RCvm7CsRDj69CmgFWGp20MYDKnGoIcFAoi8PlTETtmM
z7obj5xQSk1+eBgmDcxJOItsEXZv8gLA6lJEmAL5W+VX+YYNQWvgQ30y4hCZs3fEiIIBtlrgGIed
l1mMLH73yyf12LDiaL7xu7bUN+P12nxclx+9bIGY6mIlnSuqQdTM2Yg0EwunHqb8GIFI277P7grx
mNeW6QkjopOyVbFZYlWRNdfwtC/8ZswAkGAvs7aepm1K5uxv3l9Pgpud5biXAP6IbEET5wLQmyRi
323Vqn1acQ6aB/1/p9HMjDcmzlFVozSW+iqg5X29CrhsmFjpR+BAKJi2T4xQBctjNen1FP8wIudx
Miqz/u+pKlZXi6eS65M9VFTv1GvKn94v+bskz3UY/7U6l1heypHe9NQMdqQj0sGJ/CWfCsXhm3zY
S5KAQeTYMUUx2OWPb3YlegIz4bZKDJ8LE4feszIuha3IjVPgCAXiebXS9rofx8/ewZ6T0eL/rNxU
mEhk1bOhcjO9JmvwKPFvb1Oie4b8c/ro2EoVYwCXNsWmrho7AE70vnhFMVICw1L0fydp6aSgS0Wh
ZZhldCtCIwenmvgnVLZlG2XwwpY80xzVCDPjsNFmmZfAjDyV36jCgH2ndxj2CCWQbUeBOCXLHKg3
9MI2B1v3uyGRlGd6/faWgBw/hGClPk02xILwghzXfru0MQY+QltI1SqLNDtul8FOWalm4SD89WS+
C8rBq9hDRdaEbmtyOB4kTVqi/s/cN2o+wtRLjQrx6j8fFn2bokLSX8U6EyqsbHqR1DhiUfEs4meH
XemJmKR93YSJNY+2vv1ZKVrjrv0QkufNzukQ5afP/IjfH+GiqvHLw7pHaCNJSKCWyKGUCOyaxBCJ
dPXyqyKZ6wc2sfM0YFRBRfdTfoGPIlr1xKi+W5PFeUwQNO/p9Cu3L+YeGrWTRQNpZL99JEjV66cL
BtB/FXtnGQtUwGI/W1AN8qXFGF3RD80IRLT7V0UH6a6z4WymHonFVAir7fGT1vnsQbLPsoOD3Pzh
3R/o0K6Vtr2D0Z/qKdGmznVWeOC1WxJeWeKIFuBlxoUOuOEdMnz5yMGBMsx4K3AALa97v7V1NsNF
eUjL7UhuzmZ0R6lSDOkXfI24eFaC4E2DVvKcwFQbCgrX66Pb75saSJoSMrQpZDaB1Tw6lWpvNS4H
xxdj65QD2WtFz5+IKAdF2TqY7Tji4gqo83cK0J5rVXaMEBt7fXQb7JPIe6bWMluSLyhVTjF5XHzM
tvWylJfzrpc6z3RI6O5TfKDF4+HghE+XCy+BLUAIkhZmmMp6/iNAyno/hFiHbPIxZ5NNCT6UoLf6
MFq0mIk+vemuaQFcKJfLvSWx9QE1+gOrq8o8q4vN3SnbBZ8cmSY4950FQjrFi62ab51P6JGgVptD
Dt7SuAQF4q4cSlSe/fd8+i5ciXdtubJqSlQXZk/6AqkLVJI5e7zaihzuRtq1ZoNXQwgXEHPtq+7r
A9d9l1v2EHy7qAV4wgaKCkvDxeiqerY6lkLxRbjsJfaCtQFiBBeZsgfSaIEzHlKSUxG63HIV7xbY
dAZNeSykQeSu2vq5XgLsXfmSYfM7A5zoLz1WmIPOVBzLMbme2EQ3R8ovakYbHZ1oh8sxPdYZUCsN
oE1NU1tySZLccmGIgL+QHFK0U0yM1nSk81ZzUi724YkdHGQ/umF/7JvQvr3xU9J74L59y4KvrYVR
Vd1CQFCgq4O9liDqueKOROVn630zxWzY97tjuTkxXsu3tIrQUnORwRkR1+w1lAwz4AXzBe+vsf3K
Dzyi7tJPH1T3X5Y5QU6sg0B4qEQ5X8Sp3xgXqaPjVyyf+3ul1WCaa1Y8OiLxMxRvwJ5qBnGgVcYk
mRcnrPcPhqgNgB2eSUGRpIMBSaItmymfSMQM5iLfdrL/w55YQsXrwCQXtsc6D6a8ImxTGo98oR25
mpp0FvprOo6YK3B8HyQN/x1Wy3Fwp9m4I82CXYdHyYRfhoAD7Dz+0MCHWSNeP/Z8airuCJEpQD6m
2fmobSRVxx3OIkupuzpZVcEOHQSY9F0WPHtnNAsU4YWIg4VwLJva27L0Ja+zvR6EYRT87WWClHUw
U/AoIdiS7UKP1OCJjeFqybqDauhGcdgI2ygxIgq1xG4jxt/dthlCNeZnOOk6Yqh8Li5eGRfYOaBB
rkvjhw8Ca7zl61GG0dqkI1OP+Bkn871hHGi0PvVWRj2DgLrh2kxQ0iHVl91ie1cZiy5EoEJEKdqb
HmWKoZdAMvFh00pL9kvX3NXEqv5Ff33i/vN6fmEnFa93YNZ/vTQoEcqFjHskf0TUa8bTcBBTy3dX
vQSyUo3xsyfVIF5ax6omh5CGcIZcTGAN2kIi/J1aeXoNboAjV8Qt/d8PvrMKDHH1V8kLghANnc/V
a7spZUUrh3XWaDRslmMcX3FQq6XEabdHmknW6TWs9OBTOXPFMQjx6XEB2QJShwRV+i3lOPuZBgew
7PIXjSn93aFYcR/9W+IbgYwetB9qcCVjB+GVXmBebghSirTdSxI3x7nebdTS9wvhbDRH02Zh0F49
uX6/tf7Jbb2XCcNQYIj2w5QyQsYJpQie98AHT+F8i0F2mK6ZoqSvpRKK4apiFu0l3tf21zmBC+JC
9PX3HyvGfQgv/Azy2MDPo+XVcNiu4NFGZcX4pQb9BT6dVfhI2c6OEwj/hiqmZIQ4dK+XToUeNtLW
bXT+meq5jG1sKuJW6LobTniSXbzPdsmbKrNFQZWgUAM1Qq+HCHy0Cke64hQDbNEisglLi3V3snbL
GoN4y9OftKc281enhdtl+ubNc7PDWqLWTk7LpaW18ouaWQnP+iQvwFDSluTqmFtzz0j8BRm9spGM
OI7ncwfxXGPAVVZyeI2GjWT1Y7Y/hm9aYj4JXRHVeGAR+AU26k7GYuM8D0nyGpU4Qc+JbcFD9SbH
c0XLooJl23A70SozGrJLndcgatkHJcNFX0TprQ+PO9ak65bqGqHYFGTGP0z4KDl2+bK1hnt1Trcu
3qLWMuK2R7meEaH3pdANaTNrU8mImlZnbuXvZrsl5ztUr+I4NxBzDgz6C0LR01Yu+Cy0dGBJ/aaw
g2y9N0MZetUb1wT6g5T1PT8WIYxzgj2uE6AKV8f2f2yC5IedtL1Zx5lsMjAjmLnR6Wqle1DeiJUE
A5zAUjiJ/wZGV78HraZbqRp7VN4v+ZLxMnjlTiLmW+6FvYDAwWgzLOTdKHJXQQuEIDK2Y1B0sepn
q2CU/98lafv7QfbG+DClejbgieESwKfpjVyF/yUrDPc7cWZu7Sf1j+Od2xOxo55mIY25Xit9QaJi
7bFnIDb6wUcwh/+qzfy/2+ZtFKKlsrEkEy3fov48WpDRczGsbzyj1lJtvhnhPfEOgVYdmDGb9uK1
ht4ywRz/JfbXfvGmBAEBF24Uztih30ASwpWE10N/unOwOILGquBwxPAu2YbTLwfcHSUeuzEfbCzJ
PJ48XFn+XfSt6jNffaj88fYZhgLkJi/VTqv5PimpmKtrKvt3D6FRyZ5+1Slsrol8UTq8Esvye8+7
5448qd6sb4hS1MM54KfQ4sgE25E7JhgaHUnD8DFhcurCST1Lc9jX50OVJUEWskiGCm76GGDjvCI3
WfGx16Sh/cR4ywygUMZTm+iYsbbV7yYapIJZus79msOiLnmh69nWBwrYgihD2Ew1aI+sFqN74rEQ
HPzi/g/dgW1Ft1TVzbUshmbj4B+eNBWs35D+g/t2mFQQGphn5p6DTijcNFDVH0VtgDqlV8SqH5AQ
o8jzQRnouSG3jOPgG0esb5863hpqY/d/teY7/z5MxLQwBsJIv+U4C+bg7bvxRB8yl5LQOc9D8os9
CCSgk07KvSzg5+KdXMGs1PEF4VTQUDDMvOJLmGQ1xU2AcUnbD/bBD/dzJZigXecIhOrlsp5HDGi4
AghdYY5FliBBpHwN/bW2sqn2T5So8BkRdMkavHev1tlvGS4gl9JIzLE5g+ZIfEp7yApRF2ybye/i
XlwTtfzEzGZvThizGzzNflztIG3Dt6TU7PGAm13rXL2ER2MV8En2O1a7EwzIYy1F6dKkcGR1Vc0L
1QqwXyn/4ff3HIZfa8h9myqtfaRXvmHn5VcO2Ayhy+CY2lVJjzp1J+hGaY8b/rmVCvhvS5zLT3/9
Ji/pD7pB15grR1va6MhwZrrdzqKVouMp2dRahuDH+avpO7T771FTO0P/WeJ6wunZl8E05jLklqHU
gymkManMqJsbhGkRma3U5Zu+ZNpyp9ax3iy2wRkOlENxCB7J1DmiKsoDX05NQRAiiFJk+HN375GB
yYPn0GpnLKxOZXVtztSYgqJPRaS1QDSNaU7XhPRj6S9wZF7QRWuwQVTKc2ndQSBXOqvqZ9G1dork
pgTwAsBL7LOgsygywbHuGn3zcm2NcDUHklfEGSkY7tVSKAClJnHm2Fsr19smEVWZ2Krc0Nq64OHA
zrjQQgWCZs2Cgn4tzBM0JbSTSZ6/jVmMqpF8SohrDFOICaz3yuaEUp/Wi3LOVTysRvewsag53xRJ
ziwkB9qWE61nB052QJKbB+/xqONctbrVPViyWEVg1kkjnvc2Mun6mzuAiYpBxnflc0YPY44iEsQV
zhyyjgt1D/OVjT6ZYat7/p10nHXfIZPx1EinR6X0vJ2mS+HObTxRlYlkVAmyWX1/TiF62b/Bchm5
/XOq+L88kyLtIjWZIWTaziSpDHaoc6vp90hn5YgBLBop64pvjRtGzDZ3ROaJzTCD6Q+udFPDI0GJ
UMP+BG30j3UuuHkmsq+FJ7O/7SbJCv3N166Saq/QYPN0V1frMBbqCiR3b07KkljOfy0S7g53iOGx
/CuI6SO+k0B5FSG6gupCjSTTsntuYvT5Y58kxkbifjuFszQZVwcmgZ5qnVt8TuPTLF+peIAXS7VB
aRhvMgyT8MkPIoNeP2c5VR86qL1sEyfCh869288+auYXCVpWN1yxU+4OwigjJN8UK+HYC+y5Bbny
KgoBJmhjKMcuZUqHRr99DU6rHUOsFHxNo1ErVlkHp4Gqy5nFXVFCoqX7Bv9kaI2roXf2vgAzbzUN
atVv6gA8OteMyMAwTW5Wk7brIPae+1K1ODCODgmwGsbz8ynebcjqhc3Ja8zcoaInAFPRCOlxtQPC
HGMzS371phl1Ipv8NL4SbJ7JZpT/KuofPUF90wdMd1yvn5irra+0yLrfTidW/4F2yLInuQI9qVbG
h6ZVPGYZydlSGF9Cs9RSt8rr5JfDQrsFuDURetKDN9vVJgwO18FmC2SSUHJY59aCpc/Q3hG+xX9N
UiE0rvpmVIHgiyt3qG0CkWb/w3bQQNRLbnSVF3ssCZYGyOOG+uSR6xjO/roOaQYSTEwucm+4EXWS
GvIxoCc4GwS9TDTG9KqZqOALbDC3gjP46fo4L/o3VC/keB+0rHK4euyHORzAapyP1nHcdBAoz3Z7
sTTbNl5jM3JeLaZts7zMHaq2FA93/Cx4jjId4Zu7EEmG251NCPeBKEIHr6cA6/oB+jRanx5QqFe/
+XFXShfMnXrtG0U1ADXE+zpqSdOsPBcP5BWnElJ+YPZ4C4+HrLADgigMzQuUOVs3huTqVkaBtL1P
jIcsAIFBq++VfWmdgfQhfl1Ica27e1n5Oz1uz11FLpCNTxapfvpnY+xDJZS/pE7/HX8auQDs6Tub
remQ1khIsFjadAyGOjTk0NIeyZ6fiP4FGQ++QN9ylnCsGMZPgQ52V3DN4y5NWHy+IYagtJv+k7zG
TP0dy4lKFMofCkoA9r/LfJinSE+qUt8OGFm1m7BSgDVmhqrK5OxShyq8pCKKwJSNkWzNjmV6WZ/A
bASbwADjOnqdUOHxNC9qGqDqlVEibXFiYXgQvCN0Wrx3OyjeqAoG8RJ9IK9908/cxwM8ZAp2ls/i
vsO3PaLeyGven/WKN5u61LQLig00HkZOjbeQPOLcc9wndv3dMwCgLj+rHDFbv4lf6W6DCr3v3TUs
g3X7R9fJ1QXb01PAjRN3mRpu96UMsLNrmlRVJ+P+9+6Q2pVo1Ci6qtbZEBoxu4h3eP/v0IAuUIs7
XFu8B7ZjCSyVlWSJDhOI7xweKWOpkfJl9bDpjX7CzsBsEbuLFF319nXbGQcGOhLB19hypqoF0mCm
CO591/1NKRZFXpj2t2oDEZPul0TO1qa3EZwupuImEZwsPg3GRliNqQeWoU/I0hE2r7dcSgQuPydd
r4m92l0De2oHAgTKXIkHWn5CYGp0OpivFPWtQSaIRJJEZaKHW654knA4G/QrAATuSgjXulHpQr4Y
KUCkmUCWqkNL1llSwud5iakiERU2HyOgPAZacbf01nZexxaKAcdAYIgMjfsGeD31+VVpX/A0eke7
MmNt+qeLQ10Wl6jw9WhcxIbj4YURGr9aDcFUZl8XHn/sGYUno0FtlTJHlfWJ3TggJf6c7EJVMM1Z
EN9T+S+DFy/jGwAz21u12146U7gABjyXCJ8QJd2q81vHeoNsNNeS9n3PEmTBHcnyAhuVE/YLn0lG
9oBTttyXToDhbYDEk/eTsjorvhpXx3LiZWUlRRDwkhS+d8Ql6FsfPGHiYlw3QL2KhLH23j8hTdIq
GhPHoIg59kvzLRyqXeOoyK46Co6fcQqRhx5l+bFywsqctorf2p6bMHvT5g1rMlx8UJEuW5zj6UK2
rBcoq3JuP5vGOX12K8qcVZZFENtkbks/jyzEewcofWa6DkRS8Eru9//Og2IaQwE6nVotzzap5SzP
ha0PVOg+e8soIoQY27S7bfKLaPdF9cQJ3RYL6cPY/GdU0FW3p+TnmvJu27XDgCVIvwZosqy7N6i6
A++jXq1NYcoB7Nam/SQb7tc9PeAEenmkVgejzON7oWSjSHAdVgf0nL9K/a8SH+ucqGDXssHEnUiA
n8x1SoVE2DIOZIFCkUcNh8Zdr/Q35dAdMrzZXxVlC5vHNT40P+bhNAuTjfiSsVifKBQf7WBYyW1n
XX5mKScHKALCU8hIKXSJ01GWLx0phjrox16JhZhJY/oezWzH6z4yom8XS9+i8UrxrCELlWBydv2k
XBzsy2kMpm9L2QlQGb2XxDy9Nd1kX43qYCu4bFQ1ZTeW6zZ8x6UoLPS7Hvdo4kWYUxAWKtV6Uf7a
ifWRbGcroUnbYdSxlPGt7brHFB6NdnMRKG5/nDtNb4R0i9h7pvZUT4omWDbJSsEg+hJE7Wpyk2jV
E2mEDxHdsTHr6veWYir3ups6dlXpZhhm0GASH7hd13/KnEgb7COYY7mt7XVcd00fsY7fkS+utyqm
xYJu4J+YKqmi3HUC+I19LmM4PvwY2SFDETFx5HKHVepY0ugKd2SFPSEfAWBUBpEMSHdHwBy7sotA
YAqUzgmzSiOnGwaWs5ir2cmpIvdNnNFRl3N7eRuvatJMOzMi9Qu57R/yZDOQZd2O8Tc4D+RNA/qC
ldy9XTu4KSSv+CHEZYs5wl7fz2QAiqbk9wfxmY+GHinI7WXxcfaOdU5hQpoeqe9qmvQSI4ygniB2
w1rIXgotIA+G1pzDb8YM8bmj+d08Q26ieg386KqN4TvMIP/4O0zuG0l5YI2O2Ns/ZaKU9y8jsk1h
/ZhGyk/7OymlGRbQPqTPLh3hIQpNZ5Upy11g2Z3IyGK+BBZ1JBjjxjApLVR9IB6zGSM70KBvmk2K
ES9PVER+6RaewAhaS8zK5GDCRDtr8d+0cqbf5+GvpLcG5QrL3M42rF3tKKYuWip4//xk2nwJ6FV4
rEztPH6nEipQRwMB6ZtW0mVY0XjlqaVxC0fNFqdfan3bGbpsHLO2bvns9aHZIeZR47VuXRRfLmBq
bUzwwm/zaPqcKqaWGPaLog7Swqqf9atVlwV3Shpx4wsIw/kI7/HP03HDv8kYJyLdii1ALH/Sws11
zB7wuSwPFVYHmVsFu6bpm1w6p0OJQwoIm9PVw7NLH6e2LU28LIyGuRsQRBMqKPGMBOdnHWBASiXO
O8SK3Q0G74BP64/78y9exuFTZiFU4216D5ALKn2n2bGVGv6oIYSS1yvru/rdFycoaNg+z3in9sdU
WpYhnYGc0LQjwNe4pWQqQJZjhYP7giIyz+6fWGOdNtiGyhS0OsE97/Q0joy1CxgJJt/abwTV5QY2
a6T7xknBm0VY0kV5ClCgpM8FopnNC0MSJ26Dcs6jgGAhkjon7uqwvYzWesKbsWqZ9Go96yHmvZvY
zFCvjer1Wi/gNOMmwiQPyXuQ09lZYbj0qfDEaFQtGpxwbyGFNR0uj2XDYznzoIc+GMLzS20U+Wht
PrPjuZVlgsGKPRBx4tah+FgUsibUUPI6gkneIrdLJmob/zmqaOJjqdy/YnI1muROPGLHQE7F9jIg
yziynCggZUgQgD6jUrHXgMCDWRjm3dljX/sfu7ReDQa0ZwTlv5p2fjfd2VIM0dK1aFxAXwVLybL1
k3b1fjZkUnOdHu754k6VnX09F8QihPGq0MppSptb7SxfmbYhjDBNpkjSq4t6wkt7JyYi7B4cNgKi
IKnpT/XswwJgY8YlOxw4ULnMCEzdRbVoXWlWdJHf7DKNH2jbK5zIGcoTCvZTvhuIZpv8QEIy8EMs
8OqYhw3+RTHjtCxeP8IA/t1O2Pw5ZbQqgDNvUpGIyHnCs3W87ADWwc8cngZE9WOjz9Fyv7B62Bck
4FsCYlDpiyFKTB4NCsfmiag6+fzhDMKACxx4uZMxxBZwFZnG/D4qVtAshWXP0z3pMQcv2wNAZqFM
V9oZmI4A1UaU2A2yrckvnH9dYIsMtybdxJwIRMAj9BxHXGHRBGRurRTX9zq9n4nNQ85s3s4YSBT5
GVc+tVUdo1/XQqf7aVVX2qnlKomuOFtvmpL/g2zGKBRj4V8z+QwkQyUaGBsRVO79JyEVYG68qG8U
0K3BNUSgqPatGgV/F01v0kG0Rn+PkW1XQuPwNsAX1kADnJsWrVmrz45KgtAc7JgxT15thx9hc8sG
/pjT8QVILat18/kd0PuPjgTl9wN/opOAqyB0u+pCHODaKE65t5jn9879GSb6ZwhguioqrhHh0erk
aEz9be/TlVOgDvZ2mYMD1lBbdZ2oJb0B7g/np2wHhwdrX6guQJxPdDnnRlSdxiq4GNncLL9cThpY
Goi8DL8/gUsObSwOJXio3fyuGhTkxkIwnYYQ19XuRxK5mZXW0BsWwKjwLdzgXJ+/J30YpO5eWije
NXYWSiN8ysjEiy08I35LShBSfkwJXSknDhBuJAOdOKITAdTxdkWVRt/B43Prh3HuF9PC3ykgSqPD
gzkC8QUad8+JH3kFNW3IULoD/5aBDTCIPzQe9iyk/GDn3P7ZOYB+5CQ1HkLA7kmKQXC7oAbVYWgu
Izqojp8LaBFekabVui+WWABMKrZOEc0ocj7eSYBuKaQAR6wj0D45XbKCOk6+hzPzoRDjcjNSork/
zETTIFGlgW8Fc87iNP8srstmPFZ+tlkc9xMJLpwtAdy7kfT93hkHWr5bjXB5xxD1xzh1+ZaVddLk
CYA68KgrQT4qQqHohTSMW+nUjdssYBBvhMTj3ViqX5/olgVnkJE2YX5R+kgpguNylPKUkNLE9miw
DzsL78w8lUOXMSP4LjUFZxnLmO7dWxpju3hwX97aBFkIXJ/R8VUDr01/UnXyY+at+NCzTVi6z7bf
V0KWjh3S//02FSmKsKViBfr0ckBray8k+Pkxc9n0YrdB8L6F1ZcykN75osdww4STefBB72iKTfJ4
3U6IJQV8NLRY1+SiC6RQewfRMfvScr3QkbyzVbPP5gq8e1/yBPdd6hdmmUPJC8aNo9S+yoru7m4i
KNCG/y5px72YEGng/XC1BjEWed/iEUh9qnQhRQvFYLrzI2V4z0q6rwRSV4bxO7IAFJFv6NbxAj6i
IHJKRtclKB3MUehiYij1SPsB0K1EsTl/7EI1MCxQVZ+4xyz0zjiYC45Bv9JLQUgaAPpfY7woqrWQ
xl45QgP0OgDzpNoCa7UX+cPXFITDW5FeQiN8llVBh+W014/xmGWFs6XVzbyLPvrrhuvNsZrTWVnI
LBpoLrqsrp/tlHZD2aNGtVe42FkNt4XQ9qR1QTEKcKPAf3KSxToH0HC+CMFCa90/goW+m67uzn1S
CiC3Y6wMHzhbASgbIUokPLnFXcxLQ/zkQ83WP0dbKPs4KggsnRvhEUa/myDZX5u7MZQgPJl2jSUO
WzTkPwWkT4jNQ4jK7z6GQE2rTnVT/S4eYaj0OO//OTFGQDzKQcHSkveWkr7Y7/f7HhBbTRL6fYFO
7W5C8xO3Ox31Xxuvxmw2JDhOECWMzprNnAOS4Eb253VHeSkvxotj8ANnV0reW7M+Kz6UCvc5g/kJ
T4iAc70pQcpnIRzTVAHlpbdUAvyMSBEBtvLxXrnN7v9KRIij5rauJmH/QLCaYSDaHS6m/FWRlgU8
wyDoZSX7MP/wj8LSObHbC6+36b/+ecx+hRrF5XvN2H6VuezI7YsWkI1E2pqKPz9+4M4hSh4xn+hB
z7tijfjBvDfX5HDjU0OUpWnEvzfNqWPR3E+KQokXgo6vwULyoyWYhDjaIMh8+7LIGLo/enZUdVYj
pbnE71U29ANwPIe5RZXuAZGsX1GxTIRcAsZRdbCuE0KI+85o7oouhrtTWK4r6O4udXyCPDvLA5Bm
KjiNu9vDmAJ0Bd8VTZsyONFI6BFk5mDEnK8Pfnj0PpD/Hwdo9nKxYcHzGRR5zANwrkytTpe4Wia0
69IYlB5FmB1EIRuLoKvIhV5tfC2xdEtHov6Q66RsqrudbTdqej56i8ZOhTuNn2FWKHh/7A81bvo5
81K701y9CsmfyeZfQBac+dW3bokBcK5mEbutYw5wVb0DNRhg6UwzVF5lcEGUqx9UpYuucXCOJeBO
UjJBPmzn9K5/njEACPx4sCh3A6FjaE9p8qsda3ugaU3obSil9jfajzYUcGKzB+TEtMA5DOIL5kga
cp5u/4wHmylNQCtjd4k38msaTqs9hPRoD73HJMMmWReuNdptd5U8fAJV9AUYUxuIhoryacIyabE5
M7ETRxG/CYZGCK/1rbBeNZSGFdu4441BZtn8r9/accdHADOBHdQ7ejTnULNKIiXBReG22RDg3SjW
nusTq7zKBN7Vf74KaC7P47xgIWtJsK336rjn4XhazDJjFyuTH7Cpf4lTCXfpASz8Bji3QVFh/q9H
Q6ysTS5Jx1oS5xQuFLs7F84+njl8y0tOoiIUU4uALDcNwfviY19pxk5RrF+Qch2hut0Rpr/AS+nE
Vf1hweu9YmW1/bu1pmYoIDkbemFj2YVH/fNAXMGBFoVJOUlxVAKa1jcEpD2UPt5wFcmIi6TJauA4
tykS+qqEvwL9ayirUViCwjRJGVvEsqiRHf/wEXjzgSPCMnYDCG9OnSw5mlnyp9fAcUUu7DXvMsbg
DbdoTaAaB9sLIp56h1OF06DlnZSq5u3yzyAkQQdRRD9XG/mtH/nZfYVhiJfcUVrSXKkqK4L875OQ
2P9XHvS+tIEW7y9H/8pVIgeicKyUk4KS7w7MS0bidPP2mJhlKOjcz4rFjOmpR67yZ64+p5NsPjjB
tQrPofTwL1f+sShEbs0EVsZYlkdkEKkYNrJqj4zcgiErXrIfIPeTaZ3UIJyiqRwqH8l10pujZPI3
3YuEfzIEFtELOjUcfr1BlCZErtrsd/Bj1qbB0s5FqZTlKo+fRV+mObXuZ4Km0QltJu6ObqGTzM6A
ByGIhovWvNs4137s0iGklWWgDsBYuFi9MS7LsrcuCOJArbklVZ4c2FAyK/w4Q3aUE21/Ebde8KSq
brpsiHNzq117SeviidH+2jcYKfr6Z9T5d56OWv0Fs/+qxxNUNbwXDEwqoOaBXqX5aHpaLXF9Lq62
xnRZeqyf0Te9PlQU1RbUR04g4ZWW0HYgHiBu5tTB0X6RX7itUeN52PH+nhzz9mT2+Dtd95cE/249
ZYakJhes+RR7v79p29vkcNauEen7OBYXlxuYzyIvDbc2v6bbxC4nfa1xgNvNMxASbpH9T4WbB/7n
GuXuVauiZZOthelMrJWbgfyKpNEwvVFvlQ/lUEF/pNN0zgEbb6F1Jbl10bYeYdVGfWyBNIWkVDQF
7hUHxvn8hLweVM2KsHLk9DdR9RHPbrSXeAstrNn1X+vwkXpyO63WdWOFycpzc4AFer7+P5hkueze
WDQI7q3TvgFsq9i7XPHwUJIQLuhkKGNjegfqlTVyi6TuNwcJlgEHo+cep6anATpay7IhiaPsuEKv
alKkI8JWiJL0UM2ii9tOQXf6DTnIOQIe/QoGWPUoXCD8t4mVYwqkaZLkZbaJfdqel6hSt7gOvQ0C
pxa2FGQHQucfWOgYzG86zqES6Ncpas2pKIkWZkJk1rS2HBNHumvobjIE6eyQx05kIqPxXlfNaW8r
GDm8X6KRIvwP0ROFL4zQscWmtRlJV+idDw0StNcUFGiowtn31TNKm65DvYQ8XYz5dDgj8xcay6QA
VDQuKXkKhD5jtOt6Ja6q2HjSbcwEQjTRrnVy8jBwtlSR65ObceNooc9+6l3njxZ8bXbIRlkekFre
k6kx95a6D7yv0p6X/Ah0kTbFQS75qj62UA471omZrg8IGM7FYLTeBuREnCUQofX2gIT8clmey+mt
YNBM+vJFn5BXXg2eYBUhZgckUxmNRguHf9ZuCkU59vDtuMusP9QpFRxkJnYmhXK8/3dmR7KPhPh+
5SeTApsipCC+nJbx7msVX3dK8qVN7T8i1+yckeUQfllCym2Y0HXubYjKdXn3nGuCbOnHrkFrTOS+
JeiBj/JluX3M5GCaNc6PrV0hzmyOkRsN1glZL7EeIZwT4SlPJ8VFK7V8t8y6TPZHuvnLMnxZVNGX
cpHbR7J0Ajf/JsEAkJanmPndYFzlvWki9SHPy3RDxrvUrXMkzn96rwlSfbG0YWSb/sT91hhcw016
HiFRAOyHrWmHlcZ9/IDv5QG41xDYX+oDJd5DElClMUCsazB8WbjvVX5jXHBcCGPXgiGjV0qOnwRq
PXR/wvmPeeNY8Pabx08HZCsrf4AVe3mJZlfU0wlPlxeG3knVkkDw9JF7qKw9n1VBc36rMZSZdTqw
qbBxbEaaXaNoyLSJwq2qW/UMejPknDAZ3qM/jvcHvbx5iJeCCkdAf8U5JtgAOX59xq9cs0FqlrKU
ew5cDIPMedjUYMyS8Bef0LMBtdtZZeDnDCWI929Fiozm8WdO15mIcxMlMhrAn46cvBPs0OCxFekX
4z84DpkZvmhTKm/94Lkc82B3lDNtAQSoQbwFx0yV4QqSgDJvIR6vF1SkElwPhzixsFMieMExdKWI
svAJrHHksz5msGg7EZh4/a62fK+1ZvLr8SxNqydUdZGnfrRMwPs3n1Eg5ux2NllVSu4op7zdAuuv
/tNlVBF7LKTtrx3GkRQoAyXHMikISCD7zhb4MMrsJb4W2Aj+Q9dpKDrlv4x9vSFHUoUBDv3nUPaG
i3KOGuR9o5TpnDHmJsDzNpYT4x6B2dI4TuyhCmAOQ61c1veOuagYUg5ebMDRQ6thYJjFqB0XX1kA
PRQYKYyGN09urc61G9SIswoDCx5Xzk5rGzO3fl/ZZA5RxvzbYzCdEKHw69BRdawydM84BnrvGcPS
k4kSzkrN7pjoazbD9Dk1vUHOGujNMfO9SBoUVGwugdtAn2IUVpeT0AsUpzcsg7DDj4qakd2usbgM
4p2QQac4PbQn8qPc5UaxGo7xxW5VMSohOdiD/ru9asl+RDW7F+Z1wmmcejg4Yq++ASLrSru728iP
V7jVk2MxEUmqWdiDS5IKW8ehdToT8rFSE5i0RT4i18JrYCjpasAKwASk0vPxbNeeBQFlBVPCwNAp
YmGEHn2FufVthUAdWqIpeiurF3clO4Wva/DYkrAkSAMJNP7UgxFuzgpNrFK8UQgxEJzeqrbYBjWC
mxwZfMOZLMM8X+45joKLYmvocLZCYp+5MDQs7qaeUoBw8Gdu2f2cGnILwMuU2WcW6hPf2t89MHWa
ba8vXF3W2CZdZgyBfbJIm6frMTTASrsU37BuHQ8vH0SANguezWvpR5UEU/3dtBMoUU/5unsok5AJ
1vNLDLuXUL+EWGR6yHTjZ1+Gzcpp3jGthunL+DBq9w2aiAW5H5aH5W9kH3lJ94D0sgZLYHkWAMno
715kc/LkcmtMxAmSlKwTjy9ek23IZVZ7qJqyTtMUt9/ZgFy8XnsF6Jfi4Dvihw+/6tvMnIa7nWdH
70/s1rj5wXyD/e0+aY/tv6i6INbpkSt2w/M0gR4HSdogjKVXjHh+LwESZaEDa8ZdGewguw2m/9sL
uH0v9mmYBLlqKOuQzNl1K+xteAP/XgJX8AmRC8DPKVGipyAPDJRKi4yX0q/YnP6AKPQ0sqYmaGy6
5M4+DkUD0fY9Ihevi4AMCiZVdJ2/mjD0GCNCPGkMDpK4Oqg0/c0UKaVR4F6duImHKCED5MhV9tl/
3qfoktmUiJQfGHYwOjGn6SKEdilji/Au4wlIkSUXa4HcApn/EdH1g2hXYKXYyk1gbNn/XIbqiNrI
Zk2u7f5ADoq/wvcRuSxyfnlGt2jsy+g6gNTdUV+i0lvi0KgIAb52x1fEA9v7TzUpFZNO1qOLWHjV
oqSuKMKejLeLlX3qPrNBxoG4XYgmBhrrUvzX0zuDIsYIrOk/W0TTeKlbVL1K5ymiSQ6VbhzPT1f2
hktKKNKp2ELcK7K6GQusuTFuLJL40D6isMwOkExozmJOPkl2wZLhCOLhpM+u3qeptTgvhoKGcHtQ
Q9LHxVUe+snPctYY/0x6JNpJbXJ8t1MqGZVddtv7BnF6z8/gLJUvrUkUD3GjBJs3eujDEm+bTXCq
EvQIs6jvkOXHWF3YJsvOzBGGoPgXpW14Gj8b6yOx+cgpvmBSiEysmxJqpwV7/YFb6RtcNxwSSYYU
LpJGeK7zfKB42/U5jJn25W4xRyosWaLF/oXASu/vGCN3KNKtXtAoaX0a4025AmTF1z4O0u2FbsKg
AThSzLlCuQj+POq26+huOQK8LDwkusyiGvWXrpON5UMZucFbHvK1EC6iWEJfKKfFff+L314WvYyK
3H1WVonM5vzVVZZdiG6vG6FCW7pbf51yYNxgr87dWzHZ6wpL/XaBN/UQSPUYlDbKH5RUi20P8i0g
pnjAulY01E/GQxhJyFOvfVTV8TRbxh1u72igooV7pj7kcYw1e+DM4HRikVKNQ7G/ybqgT0vJ0VqC
qSpicsy9m4UUaxBGLcW7x5zoI8pM3qxtKEBIqn7mK+zvEBds9yI/1PSzaw3s9N51mu+9tPM557zt
I2DSk4Pk3nTRLI9YOKb1dZvmLeZaq9S19s+TnfygdWqHBPU5QX9aZ4jA8ZTDWXrBkyCoLvG280Kr
XekpGYBGzmvD+A9yXBbsPRZE3Qhb26A0DO/uoh4DuTK7GeK/Vkwp4IGsYOUYg26L3wsYYNqzNPC7
yGjHV6EGNyGBldCpJmI2tWE7DdYENMJizsAlW74GlKbE/RThjddtGC82KRdacYB79rV+HJKckgD4
+ljjDispOpRVjNr9tTK3WlcmI1wzdbucL2cmrmyImVvXDuV2R53yNr4/ex3ReKZgFZqZv6NYQjhG
U055IldA5xbNVzUte3iTwN/f3TJFQdMd9h8G959TA1SzpIK8YkYwFdrmHeCYyOPiWYhL6U4ZDLFM
xLOY61btITqTWwU3SODDZ2ivmPted8NdaYcz1/R+4CsORjVFqGaBHDlfoawPNgXn4H3Vf/R58gfX
V/oj+zgXf6U0DogHXk9HVWWmowsKFNBMxraj9nUzYdFebq14rZvM7lab7Ym1GhxgECiy5/CGeeoY
+KzXjADkS9+eX17pzMMG0I5pBx+0W4Hi0zSr8dMCv8TlEkpOT1t/OLqy+NErrLkgL5ypbf0aubwK
nQakzM/Y9agE7gZukXVuug66l86A/au675amTykQ9cmSvQiciJqkIz96+IYuAEwDCiF639YnIVSF
GPwI3evvB3+wIzQd8/yieX4EUFg0Xlq4JWm3tpFBqNAtVG5mnYFqxbOu7d0PExp/suKTSA96Q3yg
az+Xup2vfFnJ0kZWx3QsSGt7T6lM3u3TNJOUom6tghFSSJxBvvHhhOtMnxmGbfEqKH2DG//3DPu5
xlAIkE9PKgQ5Foj1NMTJGIoRJyCLMiIx0q1d17W+BD8wvVH65VOZUU3azUilXbr4gwbcZd4aqgw3
rBvhQAbcw7JvVcKYfUjuLQwiveoQez3NjmEq4gSGbgtMZ7E9toz7OONObFFnVPufVhD7nJAZVe9B
MF5LAgUsvYn3tsV1RistBCyiu5z4alGyQNqSPYjggtk9xBl0FhyaAFui1Zc7qHEL6imEU3Q/MdEp
y2/Gm3LyPQ+MC6D1oyD2Prr2hfA6Mr1nkMdB3RFtTMHZzGDwwsWm6thdUmNY7Ypel4V4ysarw9G9
0fhmZ7lI2lnl7tZHNqXVrjx5yhQT0qE64zS/TBYRpi1fXtVJ1EaIIa2zI3+lJEZy3AUIKo+uz54y
jK/4VcF81LtMYiNx1TMAFcwbgKHQq72Dv76smea4yKSIJ2rv+Kcvjw+p3fHTZ5H4ltrHibEuTxSY
gvkboCqOyGD0XLRyH6EVR0Vq9Ksvrk6KVmaIVuyBlUb1nFvf3d3MeOhPPkeHFdDiAnNGtuczbt59
yDlaXIhnZujOKhGhtgHMHRhWXCdlKifV9v2/tXhbtnaZYZ7pT5iSpHPgcORjBxjRBJweKJDjuqE/
cK7njpM5CRfuDFuKV+05wwa/YlNSpS4SzSPGbwa2k80oYGM/8r19bG3SMInoUIMBUnZL/hLlA131
c+4KJ6shW4LZW1kqtIebtvD9JDwJtZCVQpGhW4CCtrrxIMW0Wqjsgm26eaYZzjrIOEdokxujJI8U
sSjxY+UMUyJe34oGClerM2O6wAhwv0MPss/4UGudO/4+8YInvtgQT8/kKe7Ner40czesgnn9Yc57
JNIwm+Yeb13YgzMj8nujetO6ouhxoVVjtiXzuY87VFOM/Pw5RDPQQa6vTl2hgveWYSwUqSWtX3H/
EAx7dHhuxe2bLJ+EEphwOy7IysF6ZxPQE1eQJcD/8vAoLf9D+UHjf2gOUOqXtgw/SnJdDp9TXzU2
HcjoiC1yp8LrtH5dJ6cIiBVopKSPOW344rw7H2PwShptG00qddt7I9MxvmZgBNs9VnSLKXukr1wT
/FesAxbQENkGKfnOqMMBsSLr3vcy76mUg8KmOj8rdpeZT/PwtFql4iItOkh+8l3lwl8eKoQa6DJ8
YBI2rZJYqgAxpwqIhf1eTUIR3Xo0ITlTPKB7N56hDnE+P0RC5yL7uHoRsjSSxmjOMkgtpBq5N7En
VmcoKXrKm4+zcXDPAYnzZ74LACx1Q1vEw1InyxAvbC63SoJ4i0CHbh6+siR/d/q52qQ/PUVpsi9Q
rW1YvHsfjcy+OXnB3eJZOO14wQhXflOtfpjDNFbEunbw41K566kQos8NBy3Iu9tjPbIkurZh5vwr
fhinGVeuWIdXxxgqYNVkdVEEvo4iZ4D1YfPcWCtvNaExlpvsFrQDL/ROwT+b5Zxo5Fcd7e6aHLQn
Jds4hZchLEXRLOZcSODmX9IcghPWRxxpV+HKjz2pgAnFgjsnGTJgi/LCFUAQ5N2lh0ub3K4WNX42
8aYFFUTiYCzetQwkLJyOa/WOxytCeMAz21Kzy/HoHp6Ln05b0eNlKI5nXZHh78QFujOcfLlRCKS0
/OIwVCZmO+RLzdAkmcIE3uMv5o18QISsKnXqmx7OztDrpJCYeONUYdvbC6RKC/noLNIP93SIAHcx
pWHFkxT9r0rtkVQIM+pctTIkfhtF5oXNZGvT4AhcSG7d5ngB4Lr/eA6irsmfwmpkAqs2eJWkTZc9
bvutHd6B6AvWfAN2wlVmfQFjA31cwjJnfRFH2nfPIwa6jnSWfmMRUhjYHQYe/4Cb5eMJh8OmvrZp
VgpiWVdfKcw+EL8E5gCucnlt7FX0aT7dMzXO36Oh5SrYvuYOgs5pAo0BR7JH8KUGJ5CGBMtFYqX0
KK/GFAkoL2hBvgbVw5g3zX/5K4Ai4eKWfIcg1l2frVM8Fq3Idkp6W05+mbMMvs4IQbI3K3w7LK7B
93Jpyxz3+GOw65MQTlHsYKjwmFH1gCPq4tUMMwzTn+UhpPohUJjbBoS628aS3FaxJ3N0JgEjE24P
AeoRP9LgZCTFMmYi4eKotbAD+ZNiGWRtyHEvfd8swtLMNcf1WqS/WcwS5j0Kc6aBfs7QlYE63BrW
I/H5GKUTqSd2+yINBaWRjUIlNYWP5OMFVklY3oW7It1DCzkm416Y+lvVB62lFcP6nLnodXUHqjiE
1j5YyaDXDCa9rSS71SsmNZKt9cKU9wMD/p47MvR5/6s7NCTC0sli6YxoyjClwWU4VFrVTak3c5no
5VxM84C7zU7kanhyoI/teYjDsGghg4BcB9HtXmOKqLmx9hn+qGaIGUf7hjLnwPS/XW7kqkH0oS2x
i17638X7heidXJtgVqSf46eVBVfvopV0gVspgacVGugkkYdHl73Vo5p076mMR6xN73bsOqhiY2TB
pE636CZqtbJKwcBlZeFxTsRHoLIKrw1nTaBH+sIUFGevOenl8SyieWURCQ8s7u7+r5gKJdeokHhK
sFG887uykrW4ia1geknMC7fLrqiV7hAnsoCFL4gHACRG+geR6FWHooTc+JnK//z48oYNgiY0vNZM
0YWhs43I6Cny0nmrXcg2iX+iexSybTDTfLpFbpmWd61cHd8q5xl30Z3kuNNbRJEjQHN9wj6dVwY3
uY5mBDsBEOAn3ncJZu0p+99mS9EEwGcBO+1q7KxXeQaoAIy+3K2YkYj+uB+6ATp6LhELGwY2Ty8+
1lQnCU4nAyFSJimp09tP3WBARU3flq/3dlehsKHcrpcByadEj6ao9x6VZtdII3c/OhETcsp3Rl+D
KShz5/JWqhY0beyY4k9OyASJQWteM+mS8gHlUrCY2g0jZgTOwOh2sszCQNZkW6VTbY9EPSK5DC+H
ag8YvC/j/wBSfPXatHPhTjHsq+9mM3ySX10JcYrG+C0QmF+zN/WlnG+p/6HZOQ7NQ8x8+GyKvk1D
TPP6e1QzLuXBL4a6x/K/tTR6o5XusSEyhJFocmHB6b8Yd02Unfeej8g4+K0RiTsvIF+2lE+jCtKm
Htf1dqRGo1nmqsHho8HilF7DnruUqedAqkXPaxJw+6YBTNqVXcTCDmJZmQ5fuLxemt76zWxR6btK
I5/32/wKuVJ+TL8h+RlLQqr7pu0KetpMFpbGFYCw3rOGfsIkZHnlXoGn7KumJP1BNdNDS0m5N62Z
6XCBXUbd6CC+9jodpAMV8DF87WVxJbtuvebdtcI6J89aWWA0KGG9uJEp2CEVe/d/cNEglTBlu6J/
U6KYz7dFUeFaFUdSYKXWM3rIFmiIw2YL1l8N5U9kzIpyzNmHyty8rc2MH2cdU6In18YyRMvrt4Ks
F3GZs0QTt2XfaVUS+35Yv5rNC2A1LMjcUBtU7b7ij82uHII04ntierHZujQ/SD093FhyGDMG8mvd
QJTBRGqzI6PEZUkGoX64ImHRbF/ooabgFaBRXTjYZHxASdCKx+aNuWSnAHW5I48lbRdVK/g1f6U/
gCeo/VjXOnDRPMhRJx1ZFz6a9fXstPu0amr0h1yfArmlelpgK7scdtnl75WRnO9mzBjSMjY3NMXL
G1hLfKBB1531NG//6w5JIycjowBurLZUBqdjoFq4H8tdT03Bix6wwCHd5JbSKwscyHKxFo3V7NOy
BrKIrJXjlIeuaNhedggiGdAbmdMEkp2qoLWkf1GhLhDw5T+xxQ48xTWOyldZ+DzssGiDASFbnlZ5
BCqYlPzlpzAm59l0/21MBO7G3AXZNyeyspGCtfkpgLjteAKU3TJ8ADBBWceOBXJFwTihZExcTKDr
3gXbU5l8EVquDcwdSxsErtcTFVkGstxW6zh0a1OB4uGxLYGSLqk74/orvnioowKojf104FhjfGJG
FmrYGS4HjQLRPkZdiYrg3e8kMIBfBzVbdMfXrYPpJsYPJMxqkCIaLhdA6oTSBQ5cPR0+0zoZK9zC
NOlsWW8FDUwr9zXhu5Gc11UeDVBU0xulkJ1A2VRC2joohvPYr4Fd42a3KZSLsE4nf5un8pqvyFyk
iGyh6s7sZ6sXU8OONWnt2FV/s1+QYxWYvr3EMj7rc1Lw6YWU3hIkLk6ea1ug8CSUViVulUPs3I6D
X+dkbSikLxNe6plP2nD41qICDkH/2JSlC4Ay4PcmUDFNABELocGgEus+Mi1kqOlAx6s61YVzd0ZS
ucViNe1KeVX8vJYkxUoyVEVKR6QB4RYGqfmQ0P/cUQYVNsKu2nwMdegQSHDHxQavWXLEIvzkyBHr
EhcdpuWEUkT/K2U91wlOqA0h69tbQVvan93AG/MYBYAANn6DdYbNwQtNExIuClc07nvbFPWUG1Fa
dniy+qAdTaGC0MgMusFkaiWTaa6fFcpXqWsWUjPd+R8R0EO/KB2q3vbd2mfkp0QEMIYcB6c63V80
iAZ9Ak0UUYTsUWtMljPMStyFA7PLrwFlrRYs9Y8l9OfD5BiiNPuDSPSn+XQ7+8BsLkmr3cTu+Y9I
AkRaPEfOU8wyBtn18dNBOZxiUev2/0LUH4dvR7Lkz6nY/8YxxIZ7RB0uKiEsowBB2XAWHQnMYq0w
1N7400rBvZpQmwc8RG2QmWgMSSnv/s7BmWRC2jPD8/4Lt+BskDuebJZjoJ0nsPy832ZXMakGGKR+
I1bK7hyRTGGka1dbXoRMIV6yNAdka7WL7cV41+wRAMQpVDaJ4i5LSp9s56ZrDnRo/5VDSasiLBR6
rdGmoSgT6ShtjGj2BFdBGvyzA4wFbooqKuoim7niygP3IuxbGpYAU/evHXnpppq2Vb4809+chrI+
mfPl8tVIxLX134pw82pZvAFqLhauy2ANB96YhcD7JhDe9UXrFhWemS5yip+QTsHQFvOtlRgleBzw
Y7LqX9s7kRQMWiE63g/WNkCZoaJKc288XDnHPitGwrZKYa4M3dBdNTOon5WyUSBTpB46XDyX3H8J
Dkmf
`protect end_protected
