`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5328)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMKRcNvzOG7grs/8lZMh3KNjoyD
IXsq0a+K7fwBVl18ZhYb0eThA2KxtLNiji0jN3XiOCqv2M226W5135b+dnU8HQzG3ACuxZltZ+Rj
Sz+ZUvcGCLD/Ltxk6F4DUw0UJ81qQRtqdd4Ums7PQsOCXzqVeUUmg+r2vCOiscDJjQRUqrTYwFy+
YiiQiU3XWY7+othSNggVs7Z8iSWgIXTwLUrz064Fi9oEeo7s0aUB//b5V/KbMb9wwzZ66Ieu4YNQ
aLkzVulnMVmlpZajeQ2G8blt62lzlzJ+zjIzb4Qz48BAsKAIYkNPGWnd/w0gwBu42Xi59CgK6vzH
G5BAeOnMnj2f/aeM5nibJ2JU21bJSAbucHkcdtlGrPxlvN82ezdHTOgbEBdEat/MzeB/EUjO5gzt
bVJv5TDXEcMC/UKchDL8uAanRABV3LmfL4ZIET9NSehYfiht7YEnlrFpeXsWzyRG1C5bPy9S8qKR
FEXx0UiDfyd+1Baj0vCWEfcpvgrt6sDMhL+7RfL3N3mlDH+P0GqULsmO/qwiwW95LTjdICD5ZFJE
N2eBvqz9KhpeRwBjrccWtcdfxi5l4PqCh4BtsGh66ljQQ0vaR78aTW96ii8A+iU0d3H6arT1D3sX
p7hl0YAoY5RxwE/Dbh6jtPiftp75CCvZDVvo+DAeSJJ50iq+aorG/l4aMX3rsxXDKywvo1Q7JlGA
Oprr3n/DAIRjs4Tb9qtjILbf1o6fN1/GFhYAv3xYJIFBGi3iY6cqgjc5t5JpCLWy5e9klmpqv1j2
7JAfseRf/4t+B1QkoKFHJL7HcqKM6RduJJ8mAdHFaHNiwPsSNxpFTfOT10YQzg3zW25DuQQO7nge
sRUNzr/Wd8RYYwcFjHcZPkp4reOGrMt8CinY6GcJwKYf2J0fDtFzgNXKmbplYJB+zKNWlQQVwmrK
3RtFAe4oH7bv6w0jMErUS9dc6X2pvswmcufd5PiYWgSWWvhO7A8WrgezO8aKu8ykR6hGna0V3+zM
EkBjAME2vqrPSxdnQ9b3ngjai3drIW3iYJHljL5Fs/1csXqPbJxgNBA2e++B24KArhcF1eJqMK4V
q8wM+pqOMRvuQi5+UxIVg8+/jZr5eOMU1WeoSgC4QnLPwkLEFzOdiGVG/M54QKY7DPM47tmb7iOp
Xe1q8P51CpTgTDubIby3Fzw0vgo218ox/FgUYQIpK+1mq+4QpDX9kYWpcrbUOAd2iO0RBEIBNNPq
Y48n0UWqHCBhy0Djmul0FB5Qxy+bPnvCFzdiChqpBpUIAVPk3yNlE4AIfSeC6NYKPGyMnVDtAxYo
NQB6SqPoGEOwbdLIB+adF+bPqcjbFieS7Q74ioehLEhhEuMzbjmSGzumkpuSGdMvipijjsw31NZO
c11c0FwGp4dqs4o0aPZGlfKjlDdqFF7IF2jOT3Z4ll9nzUKVox1IH//L4fyWTM+AgdxcLauwSejP
QemOn2qXIfxzcyUMi0lB7jdwPA+1OEutIQjbrijiGFw6fINRlIqP3iCmshDY7ncKIouuvfLkZxDp
et0ihxUoQHNZZx9lnDa8xfgnYMlO1Ow4WkJDWKiIyPHrAt/wdTVzxvF5X1oEfSf0stuY6nEq/gEe
/5vkXXD6E5aAAioLC3WJ4PNVkMrfWwN7qkC2xOrIJPNy0ifbh5l31aZP049maSnVSqXcD6tMthPa
C7aCxcsG0/naKi57mKCTWWYHRAHqI46TtCLYz3F0ZLPezJ/mUTuc2Qtir2oLe6jXLYD97NG8K6Lw
iI4EsPkVgsImxf76RBoPCr4Yo4wBU67zs5G1eMLy5XDb5rleldONminBHj4XmPGnGFfm3+e+JL8t
gxg82DN4UbbyQUj40lOSri8ADhukvV4sd1hLbcrwvdqqXH7Q/C8B1+RxGdndb5ZROb8mTnkgRJr9
g/E6tQD9fQu17L71w1JMiFhJ96936KnHTXHKyOVrHR+E4zBVe4Llh4N4ZvsEDgMFjYiuP70sDOlw
OsNJ6orw5u7xpx3ihsE1OT1qyvDtG1qrI0IQrlbvuBSeqYiePtu3fcXLdTziK5pN9Mp7LgM9knIJ
QgA7zLlOgrh92cENGgzK7z52BzFRdELgEDVI67USu9ZEmPKB+uDJ8ln8pP3KPTQKMEghOeIsrcag
e/0DixggtATQoRODQiod7EbZGKDZvUkoZEkWdr4SoGFwejBszwKWpupNg/6VtNhhz4rWPKoTynbx
M+mK2LaUKfD5bEZAA7c+livRdCojvJMaVwGByYzGd2/I0HKG1ZjNPIiYnbEmyZmE/ksuIdI4bkkv
3aFBcqvs5JkzTrAOSUILMEQbxEtRhzP2C2QdySJZDFx68gf0ohkLLpt7rIg0qkpTfAVy/yrj7eEZ
Y4onWMh/B5QkdEJWmYwvHOhYB0RI2m3+gzbwqBvbOrr915WXIHHKQAj9deUDL9WNbHfDNlKX8HU0
HAMXwX4vdRokXqPuUCSS5bD/ixwDB5C98cHeBow7xl03wx8EH/ohJe0lvPzGpltA7k0OmdoVvmy5
i1eWO5aB334OCafiAgy0CEHUJ0Adq+CUW+xxtyCD9CwOhYwlMtmlx4RdfmIHVt5rFTFhbYwCVNXd
OwdGq1eJl+JTp9DGNNcegYuF/3rsmwmeiV2x0zyLvDw8iw+ePUEHmUfwyenLBiU5Y33Tc42J/Ams
RM9PACivcMkDJtx8o9LB6+FK9dmTSv5USDPH6Fu6dY+dINKne9koyBqFWjfq1AoTCCb6viC5EMG9
q9aE5ITDoYFnI0zttys6doAQTz+hc8Y2D5O07h+YIlNV9hhJdQ4fps2Xy4QlCCUyK2HrD1DQpfUD
fug7/odSgbVdr+7NVRwBcdBhnVXOFnca5vYgfznRjh5IPYi+JbpIutgqTtK1mZSmo2ax8308x6WD
I2/IzhujFj5c7DJGBygk8ws9EtpxZxAIalNFP4PX8Gw28/N31d4S6DwM0f8wz8/ri1047xnjNJfV
Nm+b/Cn0Qv1X7NtftapKsXaPyrw5p6qG7qnuaihr4kKFka5rKElPGXP5UDWWxXiDk/5nXdRJo4Cd
/x6vCQ9h+rG6KEN5dnab4iH+CIztDEEh+tv9jPVuqIP/LRMto0ay88pnxjEbA2ynbBJDT/eUaPnO
kbxxIzXod/mAeB7EqLvEkFn5ExfTavxu6dWUBDvg+E2/MUXCJ5Tyzjx/LZSUDqrRvTbg0EtDSSKO
Q6WxoW1LnMuQfqMblS3D5t+aK1jaPO8XEcqbsYjQL8kd1VG9aKuBH2hRgwqIXyebfen/cHI/hbE6
n3Y/9uiX41zwYqbC7Efjyax7mRAW6DXMfM9omWldt8WmjbTWogEdoxJIBze82RGxFGy5BLqGKrmz
oQIF3qPWJ5QhhEhkBhSSby9E9/8dKUBCeAn2BsGuZx0Ao+9NPthgNn0vqQ9I4hAm8EeshpLTTxJM
2zrNERzT55UTRVNpOXp2ejjWZfm9falUFbhdcgf8wJ+nV2dRwPxVo0Ll5E7bie9DT82CsXjjKGGj
AjKxtPHjEt5PwLomiguOwWLPF1YMaMuTyFpuBJxZkBsPRD0mOCHSFYgIQKSW15P+fv3ijiqhgJkf
NYJSluayNmlKbX/+3oKsN6JOk4RZnX4ydxSmP1qqnRbYAoJ4ING4xb0r3f59BU7CYGKppbDjsgaU
1/JgqCYsGFcKX96IY0lOrr6mdpJgFm///84M/VKussoGgRqRe5cx79URpP8it75qSzu5YYMWDd+D
sh0mfTkVyNyX21hJdcQ1+MOVFAx9kGWm1tZQ3392xMLGQEXG9bXWXTx/IbWJ5V5YZBD0g7H09DT8
++3COpBQQoxFQxfHaIwwZSTm2DeqrVz3E3UvtpO+ttB773kofkL/VPOHXujjDbW4pmn2djd9t6zH
9J7Sgvuz0AbIQfa0stksUfnnFvlKxx797jtAC5Qcb6hmr0ohfsQLA46cQOSo26fj9ojG0548fndC
P62vDep8W6hufoGHJnIBpu6HomsbruMvVSaJFvZgDZxbkZjZDNZXzvpV+Dff02bwLrdYCYF0Y8xr
UupUrZAZGpqKJTTOJIZQAeXmeuYK2I2UqmfFOtY1svhcUhjUz8/uXpooI5NFefZeo18ZJIgCQ3kD
lIk6z21fF6YBq0FeAsNnqbN5n+yRVAZ36KH73jv8Uky9RfG5hWHIMW+DDt065/M03froFmZNFI54
yqVHoZOel+ixahQXz0qgXusTtTu6tEtYRsmTggcx6z4VmUafct6ezt30tN3qLCKwDgSYFBmfa9VI
Mpw6jbbsrEgP2/H99GC10MLQyAGPZEeJVzyyD8KBuyaoZy40YCQWos/25JeSg4S4dLUuJ475u12S
dltmGIHWYy8nlKDwRzPl8K5Rz5cltA2DnVMP768zW/cl569MqW9z5AX7waboiPB0j2xN2luYXca2
RkQKB3T/BSJ4FGsgLu2WJsvFgCgp0qA3xUJIODUGWURxnHT55ijbz2KxIkT6dB39JwM+EnXsN05d
PX80zhpxf0vCHQqognlGT211jwJRrJYHe5ljr56R/zQnp/Umq9CYBww3SEjUQO1Rs7SNGlCojWyv
89KfDoRJ9JErCixN9cKdfAxrqEO5DGwTRfPESgTIAgOAEw7dawFl08ZcQrpx6KMjM3ZalrXm2CCl
nXn+Mhz4+ja3AYH9sy4nL9e4IgBa8knMpike5mL9Osj68QxyGOybK//qbbOlBWeVg2Ae5Ms8AC38
nv+eqyCbqsTIampP8/6Qy/POWs8uKDHGEspAKXvkrlUIYauTiHXxNM0y/6I8yHsuHyM5dtcgmf5A
nTzP0QEQ1Xe2vkSIaojS0xq2g+Q4G0o5ofhADP5ttzb7GYpqVHoKf/Sq3iQFkwZfvFLGxG/Xs2+1
zuR8rxnIqe4e6iH91TjuXgVQNqlKUoGX9jDhOwlPdHe0sht5Le5JbybvxkB4/ODGxmINO8QoAILG
cVUg+oZ016UH301HDrUm7OCIrsPjk5GU9IvISEWTLUucQl0JyqRbyv9IGQJ7FgBshnsoK79mTWFD
c35VwET6H5d2297a+LuSHnn9SH62kI2NrlUysm+iPRIUv3x+lIs0Gy2jCPM8h+GoL3s3ugFWgAzf
QJ8DwXKKWlhuVm5+2WgzCA/SK1juV46QpOVJLkL6cyalBXTUJxaXfLQ/odGO+2aAkTVf7dGwdp4g
seRqRaTc2z8cLpV0DbnBr6eoU77ueVtCGj+Klsq7BW5fbRKzzcfyEREuLCrMNkl1iQWK9V7471D9
JF7r05P8wVzo7rMNA6d3c4GhNmNlYj1fimai5b/U/00VHQzf3MvyjLiD4x+xiRqyjrKffx2+N/Sg
gcBibBTrkGNxFWD5M86fEtTva5tYdYjPmRsGdScAQqmVY8Lv9eO88A+yCu39vyumpwQ4TPKck8vq
8nrI4Xo3uihnQGSq1WDxQzgoXqy1O0x/Rh5+djRssmHRMjDViKQJ2gKoqogpZ0doAN7a705AZXbB
RytpUCl8/amgXjxDezrzcKf48IVzsBdRXRLu2FQtBtavU4GQoS07Ec3plHLTBzkwkouN42Y2vKFZ
LbRZneT4JqgD1hAnVUlPrM3kYOhMDjn9uo/wnceqAH8tEQ07E0NwT3yGVKdoT4P2SvYB6iHH5o7R
V9LEiTB4YUKpNbmChuzlWbcuEsyTRC0ihZXIaBl0Koov2ymqOdZV5vzqHuMy0wdVBUCKaok3Nvh7
B+GFBvydJ6HRW90RDPQ3yYqxbOKY5dh94RHoID0Q+lD3PFH7Wj4MV5bSP9y48/B5OxKaDnJqtFH5
SLyhjhZoPwXFT+tgoY6Z952+fHnnupshwK3j8tdb3J2h5Xh6Twg7m8BKKLcrVEV+83m1MP1ZL56r
slqsd4vCVsTfb5Q8Mio3mB9L+P73OzL2+FkzSeg+mZqv0NtYdrmRfl0oG9Z/kW2Bdeg5/LPiIjDp
aTIXX+cK/u8D7NXIMM+ZRamwqCY4KtzJW4J5tXS8nqVTsCyZyweVbVrUQivrFEfEf1ixnfiAzilg
E3jtijyJ6D9GHwPa4mmro3AXzTcZfwPwLzMTPVxw9Az1dCSZCwdxfhRZBmfny8l9NkOuJiO0HuxO
bKcxLD67yTbZBsBvX2R4bSpqeMquPjerNW81WUntkjYTmBF12flOgpC4hmAmMOXDLxq+ipOVfTXw
0yCuszMgVd69ZMvXcwRutq8pgINPt6til2AM3/tSqCoQbgv5OQxWLIUZayRvF2ZBzxjBXcmzRpSR
bsS1bcZagPYNeNLl0ZRbuA6C+MGGE3Xj4WvvVz+E2YjCvw5+Q/E76mMSS4dZXnaTnm9cq1Q+T7tr
u92ljN7HlLZirxAUCaxsAv8PAW+40czuAlEWkynBQDHxTXDG/dMnA2pzJFgoNY3q+KdnALheSq7e
quTuoPO9Pc94IxxRig1D4myGm8XH8hvWgicwZ6b6WDBJrjbGcfXXEkaegJAtrTqPLqeVPHaQb/xo
yG2JYo62/NFukwAE3IonSSfBRY2dueIgMe0VaJjuIFlZhFGXJuKaj8nXnluDKXxiP1pfwAeMt751
ZNrv1Rdjs4urJ2Bapnag9rp9cQGKvvnFH5G7IJH6xEKdv7b+Ql+2bYukSXt4UaGzRtfjbFsegFAT
6tsdHnkJb37xxbkOv9WrjGhM4gVQaWE5ntFMAEu/iUvrtoXgkhdunUweVhPmdPpA7c3fRPLcplHN
+mKBbpSSVruU952fVQJ0+256o4iIhO+Qc9fTUxTB2CZqoNicMZleXvWt7rU1q9K9OPWeKmfRW2jg
F8FjaEGfKBuT8dz6OKMwXbBBcEQ0UbAsZyd7zNW2CdAsa+2GgWvlOs6f/0yPXxHtfXNasEodSsLt
LzG4mKJx3Y2TbAtkf0evnYGDXQEY5RgS59+MtS1VKxr4ueR+pRZFOPjgozA3MQgwo1tOOJdnFqv3
R6fRbyLttxWgE5H2SgZmj/4aTXhwDaHEYD/b
`protect end_protected
