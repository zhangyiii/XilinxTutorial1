`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12608)
`protect data_block
0eB40Voek3XE4QOCP93RnZMokpuoA4yK6p4m2ISYcReSB9ICFfoz+B1ZalafF8mOCyPYN7n7vhGO
NizHpIO4c1JhyZLpWkne/hE4+YRP742feVYVqkU/PyvVKAKKkcfQfdIDxzek6HS7QF8WqqrLLh4s
I/L0Wjd/JstujCf+q4K0hLbWoDOtGwffRE3ieEJaFdQ1veDgvN2WbIai15bVWxBaezCKP/hCt05r
fN1y8MdMnUQWPt0HI3zFjjiweV/AEHzXD1Gwd6qJ07UwSXsS9iKksARGZdGwOsHy3/F6zHjaWexC
Yj//FdhD8EFY1ELG990NBqOiVJXAoxJh8CwfaT7J3Nc9vXVxz43eUzMUOhE55wg7c8qGijM8YCR5
uq1QPZxF/VDP0r5us8KjWp/Kf9ECQKb8iwIqLoHzVuz3nZlg5waZumYvbKlTWUU0Qa6nZIbg0e4W
JBnKr/aUjCDJ7FPL0ABhgAMUrZmwtYmZIuilrp1bP1oolryN96yz463soj3DTP2diJaTq2duU46L
0qJhQk/LQLiXIYoa4eDTQiwrZRc6l4PE2v1J5c5doDwuKsrxNg2aKquZ8g6JqDNpWnl+Zx1ksxeB
A5gieWW7g18BuRuM5nHpobRn8bfGtxtrydgmGjjnl0dhqM637xji83f2nESLaqeF7KI3+ws/diPj
rfEVJvp09QAJvX+wtqPU1GleU0/ZoKUcC/syJRPf7euqW8qtOvDM2W7c4iLWEsZfmzDWSVjrHUCJ
oeJInL7vSs1fqfI5nHynTwY5wpNheOzNUXvfeU60HiTbsxfcy9/BQE7TP1LZcYblXKwx5AJx7yRA
ky6JAknYJlLr1cQgBJCVA+7J+CBRZcJhCNKhao1iCzVkAjo4/ARGT43mEcDg02qsObMtWJupEWAp
0xcljQbjFrFjk21+C9dxuxFbd9Z92KxjUNa+rhgjBu74GJphTNd2vD5PaMTmG7sTi91NZE7sYigY
Qig6d+3o2CYp7lFvbrhalIS3btuE+D0UKsSr6afXgeourYMwubjmitSZZLiOTT4Vza29UbbTjXsX
aL+nrzVVxB4AhkF7Aji5fE4edxyO7LPlDXwdioKR2fNzknV6HrhAw7UQSx1r8CEeGx/XKR9ujvLk
QpxfegKnf4CAxhPbBgbmErBrU3rb6ZHlaFPYa2EJqJwNeBxaHoUptd2llIVEXe1PP/y26AWaZxHi
T8IKbZE0xnldmeKxi+LYgm1p37HBr0Pe/PoKmAlTsc167CFNwU5Dz6hfgHfIEGUVw5N8jxfN7nCf
t42RUxJVqOs8PqJ6fT4AQKuOWMeMr1CYT9tPvqGnFMS/PC3momB63x6gzm2J3eXT6ywvYWd4cJ8b
ONjCMHxowl83hKDPi7Q1hC9PQBl9Z2FG6dqq7YoUmvD9NzAP4IxTXfFWiXNEKUv3W/cnJSPGt6+F
zzn0dwM970Dg5VYjC8KkbC0z3TFR3fp+V21RMNgsR6gtFmEZUPBbFd7uBUBX6hCbiZ7m+pyeBt4+
LmH7drH6kNft6y93wTTXqdvaWk7ZsgedaAJFgFtNkd0gP2wr4HUYCJDnYNGmc43UyviP6v+vhPVT
wSZtta3YJ9rQGQpUgl9YT5x6Bqy3H5TW+6lv8l/mcktPfaskVi1hA3zvbYA5omwbL/IxsvbB0eOx
XGIcu6kyyjId+ldkPhL7CZDT2wQIEOXyQjYDG+yjPpfXn75ExdZWn6wdBPsR5+LkCkJe40d3xg/e
kZhTfvaQf4l96MS9d5+IgvPchlLYkML+3gPyM7nUTys7ORmacO+SeaMdjfBs5UYxE2jZJuv3RhMj
Qqb2jnZz0EsfYdqoGVwmiRlMswFnxaGYeoRZOWNp4MrExdHGCxw08oNKQ0/eui6ha7prl6Qufm2I
il68THNtOl7kOJ5/GNCZtLponis80zuxLEK7PnD88ec6CWkUf+yAHR0OFWQKxn3TbxNtdeMnWufu
m31kmgBpeJ9KctymEA75VQLLtW6nLWWjiy4uh4C7SwRopbk3TlvKYXIXvxnEJ+KEIaNwQGRK+DJM
46S0HH9mIEJRxf1QMNGn9TgBPZ1WYRZd9V2+pj6DpblVLXR7fzlF0uB4D4JpaSFBkLjvAplGZedj
zhqzx2rs04wsggp3KadkBRT9HqrG0V8PB7vTGZorDNwmsHe0JBySQf23fkKe9uHzueiuKJ92/eQF
4uyGGfAffGhvwgjJJmTj+wphIWULpDK/RmS7u/wgOiOX5A0ZzdQwevaKHegeaOBpfR6FmH4xw6OD
XZvgC+HrWozcdiZpxfLqvFYYUupAVqYk2Fk5cG4w1GhQB+ewB/Xo6OfnUHNBVwe7Q+bS5cfmJDQU
+pUtQBIN6wJjRWO0cOn/degd8aYu+ddn0DCtCbnpCT5bTn48iH0HFs5WcFB+hjx9VtPratXUrirm
2sl1ikTzIccPCiuZ5FRBvNVGB06kmGnbAN/kPgV6UPfSEOOkZjsqTvdXauUISE7JrmclftGetx1z
a+FpfmkW45OMbfeXd811+WaZUY6RBzzda0fapcsyuorsbePCSdtiyeNYJr0emoVrZrVrozNPguzz
O9oQ/OUIh9YRp8Q9D6Z3JzRT0Bpl9dsNCzydkf8cZOYNiCzvFqPxRdJ+gt9kFddVXWa3EjLLWwHd
DwXC6eDd8myokJiyhplDGI1i9q5vQBpGHsMsgFkz9DzB5ogVYuPSQakWVY73fUd2ede7c3j224h/
fkx3e8lPF6KI+6pKubKF1vTy/BlL/1UdTXhElHSUeMURJLTOL24K80SRU9S28bBBqf42YxdGMCIH
v3W8UbPShNap9d1t3OWITKTvSryh+l4t9X+mRQWb8tG+nT9FpzgYbVgIaHcIoA1/fXUxZWoC1K8v
Tic2vHcEE7aglP07/Hb7OmWgorhl1aXOt+0EdO6e7EDQddXcn8Zf3q+o97wcetXEanYD3J4JmUaC
HbvaMoWJ5RgDBh7zW2PemSsIAFTTnvJ37UkXp7TqhKQCbtxUZ3DFIbF5ZkjUWeqGaVywvuYpSi79
TUIZKZV7sSCGsAm0D43uOiT7TEWQZGCJelbx/fIPiQESkJOr4lQvIGV0ANtgEX1uL0VhovxLuEqT
8JBrAiqp0LEigxakGQfdRWlYtGJRRMoR0mLfEQYHQe8ZYrAbuRcK8lNzdOTK3tA03SRep93FW/L4
Lc+E+Q/P0i1z/A06mVlbHN0EvhjqQBNgil9389ipj7ps9vjS8vKfJGbpXNjgg0B3p2ygZP6/DHN3
BVcEa8ZTMVb32iqKW94mUFAwbszcw640EXxkPkEdmQmC2WzTZPOMOpYMBy60FPkaVWCIsFeR5Wcn
OIKPCp6JuLlyZeC1Mcazy8updb2+M/YEeC2O4aSlAMUfti3tOP7sqL4ii8ORgqjaI+oDiL67lqYH
/CDBOplNDAvRt1wUsKZt3uLUn5xyDXVLNkNVfqy9FHNxuTIiZxrgpkK+I9ABH04/We6ArMQdEJL9
/Odv4O6xFnf4Iapwgf+IprAl0PUpFwDE8bEQYS4HQLx2zfmHDWQB51o2wl6t1xdO8hkPRynROr/v
kGQ2xv+IPqXimXPD8nKvjz5RFvjLJ2C15eJZh0ftKCY/lP7reLl1z+KGesuAC6RpxUcfBj8nwjd9
xniyD/Yf7QxZIhJBInpq/mviBh+GkY2eJWD0AkWGIAHuwYMYLJhv7jX0yZFJNXWlzXHONNsEDyQ4
UsUYseEHlntaPhq1I3X2yvcBqqAdK4aeGC2kCl1BQhZHw6RbKZrdrEIhnhzGG+3GzRWzXLg9tzAt
Wq2PdQkaJQdbeY2HKC04qC52dHe6C08mWtWUUu3kNIe2NdSpFM8bt+KrQ4AxCNe3bt340IaNf0hd
DJD7IM4ovWbZgy0mCwyEXZP8WKs7JwuOH3eSNmqhq3E54zBLV/dSLEBPdKx1MGzDd1V+/AYhiU+B
Hpv6amNxeMG9ZMyBp4lThbLaTmaJhjCBPiqGd0GJJRXMZsNeI4kZ9RQ8QlD4LO4J7w4E9MG+f9W8
49bctFU6JilPEAM+KgO3eMBAbUp3QGp1szriD+sYzpyhii8TOTQRmgBbSOKJacvgCKQRVRz78g0A
aRPnCMgXcFWfJO7ciWs4wz0bmKCA1UUrCRfQYEhAeEBIvE8bPynUv6EHtcQQpq2Et1m1rCVaIw+Q
Lk3h4xvg8Dpf6psR7U3stpa7TS8bD+OYv4cts8tu8xXnL7lUcGr+kR8UE2vhnScuaxlE5aBD09yz
CLuKVGQFgUxQx2HaRSvY9FSZ0S4o+ZPaLpNKHUvv+Wqk8MCmW1ntWQxCLTt3R/nrCqse6XnQnRwm
tZJxLduG4BtpDmXI22agtg18njvR0EpgExebQ/W6qwsKvielHrcvue/+E9BX3e3/OqjLuzc5oCbK
89UmcZGOLGJ7aNxA7FoD6Ruqf4K2E4KgB5HQq4h9pZhWfWRJxs3P5jYc1M7UKEMdj03lItsNgiaK
eia3nAm0gm5CO52KEk5v0ngFEHnUs/fXbfuics0mmGRfGtczAggmpSLsEixBW4xShnjs6rJ1JZb3
9G3HCmMbqjKA97c9V51Vz6lWZsPMkZ55ELJoEUsSutyUoi6uJg0xa4QdkQ7HbD2D4poxHeERtg5Q
w518hytnS3NJUVPLMJzoUkhB0UrdnGhpO7eiH51KL/sEZemjjKEAtZOANtkTqUl8EWmIbXopsLym
L6ZbjzzgLsb9zOIFe4O4mWhSir4h12sSsvWmEqNII0LRRFQpVZBv13Ho55IOrnHehzIQ5Rl6mIkD
mYatw+PvxeO03+hg0qU2H7EC2aJhNCixmrawSip8ZgxhBIrITCKj4EneidPY1RvNYrv8ZmcHEN37
ZSlYTJDBlwvg69OPloIBRAElz57u2IMLNFHw0W36FE8/ov09vTGBKI6ksjUeOCbAGspZPtrcxnAT
CuyEftZ6pmPp59nlXX0CcLO9IfID3Fw99qQuC7TcdypRfIvzV4fxyxa2wHUGiWj02btWuEk2clKi
GifIZafythWHGJkIIGoJ7UfKbzu6GlRRxv+cCRcjCyAL5+Cwcl46KoAbXA/tBcXdqpxYGlIhxHFF
AehL9cVomrr8sTl/iWMEDz0TJSKVFmEfU1AgGBNqvOG9BOkoc+rnsLijQW2W2XP3rzXYke6IehFU
QHLJ2hlBE3163hkVUaQWIGB3VB3VfEYv7NPm/WZHbIVo+qWfGIPbSKbazZNKGBX5zYTLhqzMcpPi
Bw0JFXIhesJzWYmBIfBVAfSrCt4QPj9jc0I/h50Ca6JLCN3VTXePq36TYRBrDfQvXln9VgO1Z1Ve
2PSSHPaZpvs39Cwe6CF6dcQrnKdvAXUF03vC51VdEU47yQgGcxbsYe/Qs9BqkCWv0gInCci9YgHQ
MX3nWJYhLZEV1yw+1Kvmesn1QJISm4wIf0XFiqu89Nci+iISs901gOKS9QjSUQoI4F0ngl4gVdfe
jtvR46UqaKS3UwV2hv+2NCq1+5PGCbhkN2NRLSt1TYBszkeRkbO2fVtQ7xZPT5XnB/thoFk80T++
0D/ir/Tx660ZQ4bB4Oj4pBaUp6cXCnjZbBLaeL3nrDEePVy8bHvJ8XXV8ruve9fTPkfXFoS2plUb
GumBM1bwDMHNR+9ga/R0115zA9QiSaFWZNDgHL2pm+B72ciuYLLWAkbqmvBjhAV6vdJc+snXT9ru
YGShr4WtqMnK1RjNz0Bn33qdRqzBXMBaMQ9TiA1vZdPwSZUsUoRj3TV/z2bFna6i04THd65qTXxv
neztEK7Ch22Y47yoTDMTo54Nu0KwPRcbK4RMOq9XVEhZsCXWz79yYPY77RIrhgOi5V9CXOAREX6d
MbAk1P6dDlJ0tsS/QzyemzEeJKFFboFBGMW/OK8s05pNjo0Gjy+xVGUoXEtGrEVgifGW0mNQwyMq
9DA6qm7N7CEHCitcjJyslV+nS1BgKIq052Glbz+p74x3EMxbe7kiI3/R7dqVoyDM3nBY4gwa6k4j
dH86SuO7SpSQYqh37YRjXQjtZ22HlbTuHhfcLkE9vF1d4sag9SdZC4+ycdZ7p2LdwWue0Py+Gyzj
eLjaBGtW1tQ42IZ8p6LuV8tblHHUhNj6FDU6aEFb9byfe0MeyaLBut1/+AHbRhG1UAWYxP6NFyLh
MtZ1z1zSUeGlx8bTbgvJdqcfRqwq/JfGEgdbYeg5HzkaQnEEynswQl31QkLe2OkYYvYDrEivHtrV
hjjxqpljQ1TVJnNmsP5ft80BOX8Q3ixB8jXjvi7VoEiRF/D8m4/kSXtPEWdQTOiTSsZCy5Mx0rIj
OJPl6jJ3nTFkdCz58TJIS9CQljhfMh7BFoIcGJWNe8tdJHCRbxq1uGXCy93qAs+ISzhQgCH9BcpT
uk/k1cfznUuoNRjDjtmstCZIKpX6aZ3cZArE8tC72/ugyZmkcdSeonOsNC68Pz/h56ArzVsxc3iK
bJTh/84wB2xNs2LSqiIG+ZaaQ/nY2/G9Vlb2YTjNB/IFJKzl+3uh2wmtD1HTAf+whXDC1mhsj3AU
YpAa+Kf9rRU7z8SfLBDvhF96yzt37c6+7h88j5XyupgppnjYuwrXfqjKjwsx1iEgpoaidIWz/NnH
vm/5Is/NL1XtHshKZtYpU2aMxCB4ud9kKy7Hj5GsHS94cNwMQWUybK8Oh0DfP2ho0M+jN06H9Lp7
WENM8214G9Qoja4u2zU5tEA13gVGn21jXDiEE+aDCFkNzO/zDvNeB9PB0wyqYceBikXeEmg/cIRS
tNslHNam98xQMtcrU4bO/bi0F74qvMUl/+BQj7jF06FEnbiqykn7nmZnKF8U7LroYMmqsf81/P2N
+AsWXQzoQTEHcJj39VXsog36aCjLdpBUjjRa8UJkv3XnPNxr/4FUgOHYZr6tO0Z0geoyusCSTa/H
DuqtRnE3s50hfY8ma1LiHKNXpniHgZyXjXKSEPa7bb+PCNrfKRn1fGaLnuyOGgzpppYVKcvSE/AN
1dwC3bNYNhmWANej9Aj6yRCXWkxb/uxCjSSo/jVv/7/gX1n8dYMndEUq0P97TCZuv+ijSvRdJHgN
x8OPqW+KSBag1+Ids+eYVKmMzB88JCVmTKZvfmvr9VNkCVau2bjoCXylFV4Vg+FsD9MkD3O6+N2F
W4fMutM9FNeNFAHYyg9JoFHD0E5G30zhg4gYGitibvKlEKMOmYll7vHpwjeUzjEqTUJ2OhRsz9iV
5Sqy9w9wcq0Qw90ooRqQmAYvzMq6z8zA5fqbJ9JDoQ8XsFDimaVHswZK4NNwmQHZhmc+lnb/Heha
sOF25LdPE1l4oRJmhJpqPfVHLHcUG3UVEZ2iCtYZbfm4pniBRQbZ98YiHFphVIddUfT4I+r0IhTF
vvgnuYQ2TsNbY1RVVD/+o4atPq3Ta6JHh86EU0htK8f9n+xz6WQ4OdfW92ohiFGAaItyu5IZ19I/
+5TfneTnl+yW9nOOtpH80V/olG6QpS/mjxSsazdxVh66QYwOpZHl/193Mu932IyNrg4X3DoM+BJp
Veb6U+fGl8BPxzzxZKDX55aCFEn3SwBio/rTYTLdVpXwSMrYS4WnSZGV6eE4Nkh7joyVuVbAm8y6
MVdSdKDKGiK3jsk1FefDMo2bo4tfAic2wUG2T0Jy3MDQkIvvxRNe32mpHjuKJSSO+FgC597Qu4JU
Vjzg5T3oGrA8M4H6nnMMbq/BUgq/0owhTsEbWF2NZjHD6lF8i9TDKbYVJ5MTpZC001PnVEoXqUVV
ETW6ebaqbhkat3tuoK6yAi0JQAkL2kEKdBgdHLouSqIkdIQtl21ebm04dE41d7qw+MUKKBxbMe0l
xwRP8YpIkYShTseCWYLNmsDKoLvbB9VraMbh6w0iG7vxGIatNMsjSTYrIZpOTdtc4ZFuziqobNG5
xJiZ4KcWWcHwzSOIoWJV1fZABVVXc6663aLY5MswaPI5TEI+5R39DcmMDBi8HNuInG/k5+FWPis2
PY3x7UMnX8A8IgJhxN5kv5SwiIu4oSl0S8zehBdiX8lju+cDNUbjYL6AqDCXaJgcHk3zJPsANzKo
WWJhfl2pk4iNb2w2MTwB+B8V+yt7f9dPjuMWyxsbdQYGvfbr5H1ewjtEyUDl1JC8EF8RFrQlYd87
ey1ltE6WVIlfrOj0D7Tzf6rZkY4PIGAFehBVTqZo1i47nvyGBlDtCK89cH4LkHvj5TL8ekeLFlpc
YE7xDpG/VENBR+ztF9zXPFq724LuWR0fyHIWrzvGHgA1EuExiCAH5ISwmslomvXYqK41UPIK9XNr
enXijR6mP9qNf5wZYQ04PK7k4Lbfr2Awsi7lv1lMWm//Sdh75fjenEoUhAOuhc1V362j5CvmlJ9/
VvjQ0CFf5hIk67SG6ZdrtiReayLXj3HgaeT+asGTMhKWIxuB5+BbLWUIYnGp8UfVAS86+U+j/UHX
LqMwLCt83wJYiu0tIjD6KY7kk3aS0Rn4rXtpmLYX56ybZcGg+JaWt10pju/WwCg00iMOBU1Tv8G/
B+N3cwcdBpGKQUfO/+lfaaQ0SbuYjA4CLREqr1aJK//AtZF0kX63qQ95g5g4+9R6arETPhS6US5v
xtz92LZhCma13w20LUf5k/LzkgdBWPPF5UvzqqEF48AYyvfns8bOCQ0d579MLHQZR6snZxtmzeUv
GIcMxO5R/wFg7nZoqpaPvOx4QmY/YaGF8INkaWvWOgcO/YAmMLw2mkhPjSM0TdC3ApuyNe93XcPe
9IZ+ZZofrCaA22PrA6A2WfL9ZG/kpYfCdhkhyNZli2MvXw6hl1fqHnfRk9ER1B4wV6NFI8qTET9e
cQSydF9bHuC6/6X+esUcTmGVeQ2E8qxt05HHEUjXKAfWEGg9CVf63Nyg4A3/oz/EbmyehkoAbQ2e
wMhnf85KCnf7su9UzlsQKQyQujiIytFDH9XY9QODGMd5NeSqt7idaJlpFV950YgsJxkJiOLGImkK
jGIhD3WCetqdE33OlJnE7WS7yJXBvGx5xxQIgb/HwulCjjnkr1jJYvnn2xk/h4xcZ1w5GVeST5gk
dXJMWO53t6eLlAIkvcdcGEfLbyW00cKR+BeQ0lxjwVtPS93Gay1gOwRmXz6M0xaIV+C3eaz1RrcP
85ClqFdexvwz81pbmzFwfUTO/6fATSOsrfHz9S7H35b79rypGNeRynn5OIou89+29fuCatXcaPQW
MyAZYNk5KZhUe4ZmAKqZCBSQvUC+ewpNAeAXIoOTv+ioqmVpxcXdYSTAv32XTyN5e+kXB2zXI30m
HV6JVb4XNWmpDzIUYq6QhCWTzEPeOo/3FDq0DeA+7VRz/G9bRPyWVnmlTLgqkpJlEYfc4ulJibBj
YXJ2n/sygj+9rZ72mrYxG+nLCv4SHTndjVxwbVUYQlo/VKRI8FIC6lEqjq4f41Poi1DPd76TFxa4
WnLsnJ7h1KfQa6s8ZzptOME1ltlGwIU2SI8r7fD66XQcTVZrOcHYFkoJQxuIXszZEqPI0778E4xK
vzYjj8OTFVdGP3RrTDJXiTTcdXlBKlZJZERYp1FvvBZAWomIql8ZF4RMoA5x9RJBKXngooylJCN+
QthwelQXIZNhytd1hLpVVpd0Fh3xL0QG5uP85OHSvfkGTlg8OCcrX5nkOj+iZPjIzZRAIiPLxhFu
lSEVACdsJ3xPq+FzwUBL99AcUukX8KoIxKnZWd2QY08zuVtyyL/izNp6a3Kmbs4kEQwPyIh9TdK/
ozX1IEX+Kmae1LCp7MymeOW/iF8YvYNtbJPLw9pb7TfTbpMHbdRKtHgRj9OjzVt0jThLcvZekajh
ouuF1qgfjPwdsPHKpToSTQ4ZyHXaifr7sUZIvkTYDaf0XYs87Rw6+6Xe/cvl9BmDEbvWfT3Vr6Uh
QJDz+7ulDaGh+gt4CvWfN+iru5JLRBda9Iyokm9Po0VLvKzQ+WjLuHRE6Vk44pOYTppxrPcZwqMU
Qnv0Q07uTNOdGAvd7ei1fNJewvx7jjj5+g8R2WQT9iUj06CDzhLAFAuz6pH7bpJjAHCiUM1XvnrG
wG8xMUTqJNjsGCxRAxjSpR7fWzaH5xqsMfSHhE9g+Y5cxo1cvDRK3cdv3WWVCy/u0IBtbJ0wntOI
qqXq9bhsFGsP/qLIGbD81bp/YA5/kggCOHU5aJpDi9fJhIRsf7rORlfXE0jxrmf1Lh5CdE/DwZZT
u0zDGumJBzIFaFAXafsIziHOZA+TailQImj76ThUv7k9hFPJ+uGxkh4V3hLE4G/pxcW3cOdgTUh7
sdhFO2i3XtBY46nTvxVL0z+74s5lgt7J1VZiy7VhCqMxnSIn7xh05UpsIdOuD5diwhyvAdqR1Jba
cdntnRZvjOV4fZ2fZRmWf2+7bmdWH6bOlJkk2yJ1FJiGHO6SMTpV5pDJVx0DESA/Si6vi+JLnReL
ftsD8VE7ORLE/WjNuqzHO+gCtpGQiLSTa8CGo1OG7nH7cEFvuRCDOA9bnf0Cqqk2Z/pduvIAqj/S
Xhr3sC4MLAE6s78Ag71R5r96xhoJ8s9mGmFkoV5LP0Zwo5uvjgc68FW2Bro8k8l4Y8Tcs+/ZFlyn
uxo9qchCAYeyco42rOSSN1dqDKRAsiNhmrU0klDAddcvj+IIl/8R+C/5RKE5Zs2hGWBLw6J7TuJs
tjkW18mA6mw0XdGs1RS6sR+bN5UMpx8TtAXepYXMTNRxmZexaYC9m8L9pSiNIiZui/JYF1ACrX0m
9zQop077GA7qWrpGDMkMvaU4BdhODwEoMH0B/JiIlsLTV965HP8IUUo3Y8oy10XM8N1A3PxCC71R
iNr2NKVlosmbdCseTqea6WpyrTXC8OzDq2/4xvus07WHS612m8mPptCi9VpoE+90hpF3F0Nbc6De
1DPb6f4wJzSBJHO4EmxBdqleq/lywRT2X2juDNAVUI9R3Ma4kmaIXSaN1bsOlNuFTxMRAC593vP0
rlIJNqGu6HJmuwiWg6NiL4VYYqW7/kbUTugP7jmwyJpn0sKIXkdpKCWB3hSMAE1euc6NWvhAKpHN
QEBWTycCSwn74banNYprqGE9TPZNtRrzrzXIeq6b4elPUfpZ/rGYGgUC32Ipp9QjRgFqk8k8+ydz
VQ1YOGJB5wpfbxJHn4gN/cGtEoLn0ZIZnQzgIMvWAYz9emmxPqRfT4lfsH9ohgSPkT7G3J/P/Kge
8dl4psCDN6nNAcpWSOJbUggIC7xYYHDIPddW+v2v5mOzYY7QCSCZMO+2cd6/WDTrCk2QD/OQ5v65
+T35kdhzIjfWR6AC349U+KluuKdfgisMSVax7gUsc6dNVxZ2h1hSASdIwsa40qO8zp11cA3IqC6k
BGd+FeGFv0oA5Rd+iuKROpmIg3XEFUjljhs1EXgfzzpxPpOwoULLOhabb8+wDu4LF7pg0Nirjlj1
M90p9WJhEnW6JhLAuwtl1GgStBvQFQn1iT9yc02GjRmE8xZAovd5wHfr7jQq8DtOhBuwvwThLsJ0
E4fRdqQkYH80/HAgs1M2lWyV5do18MBgQkkz0UGw0xJnUYyTkvxxCDJm/lKabca+shElCJQidiPR
quqCLKfntIM/oSZP4M+baRoo5khstBTjsdv3e3/e2LNrLLEo3ITigrNwdB8bfo0KzniUhzIPbyCG
SBykeRWXjmmu7FoGZzClwRuyiNvzuc1CEnu0mH598zFzzJeMzHG5zi34nmz9X+kOUilWGflRYcD/
/FZTCuex903uaptEF7e+Em0sVGRfUPJ/dLYnOaUaKFysfIp4UJI7Bcfi/fhXOBfqf8pViCAy6K/i
4/zr3q0DY+kU4XP/RaAfsVhAtVPe0YRau/H8e5I3nqtKfS7li75O4ALAAYxLSzK39aJMchtfgZb9
Y9P2+BTRquh3EtjGhNQCf7hZ3ifL/zgV/txJiD/RBLSnx9VphDURNjaFN8zuRc5tRT/sR6zhrbhz
Qx/hle19ieXdXvz4T2F7hYtIe+Om57bU/aoxaXoquOejE7ugp+OvdU1wl5yufeeEjqZ80+RfbB9u
CvuWFy6DOoVdzGr01eK//7TKSvPuB9sG728/420urZlo1ZD66Yf45r5+s+uqGF4czNuz+P/EZawk
E0zNm9n9yeBPQDMvUFx/zgdZPVLe7N4AF0Wema+vCsc39X3xcpWtyrRAcJipDyToEwsMMg3h1lhn
/WMZhAncmyddDpm/SKtNZrrjLx4Em2vnA3XF3y20zx/bwGqQe0m6oNmzQpnjQAOaUxjvBeU+TGhW
anI9cBl4nJj1M19pFDnzm2J+gzP+OgOl/WAqpQbVQAwCDbDqYf31/dJzIsRV2DxvViBeYi9ACgq7
OncfV6PDuCi4E2fpQ5MDY6Ws5Dypk/EcPA2N13RA6S4ONCcXZBJsq0MUQQ1gCJYJY28MsGnV3TRW
lKkBzYxD0R0L82SWt8WepWm2AzZKjX1XLKOCadxne3ZyNcEyg5BSA+YL001bBBf7eJ7eWlXnpgXN
yE72OYFv4dMEUI/vS+iy0qL6u/nJMke4cyMf6AkbSsCQfOMJ7npVCZsLaNJWzqKwtA879GGSR32r
RPwJIC4wo7fdI7KOguXUX4eYwShszaj4XHKIRArOn9A9+WQDpMX5drklfa2N/Wmf3Uu8Dt2BUL0Z
R+yNPNP8Uv5GHpCGH/9EC3T3ay2fQ/usSal3K7L9xErXPGtC8ofrfk0JoVUZEdhS5b1qigKP2sgY
iyRuSGphOZfg8Gp3wZL+zea9HVBBkr2wqZyAwx9SFwMJ6m8RavwCRuTdtRnLmKrmFzCkCLxNwP+I
XoxnxTvIRoTiG9X2EBlc99MvImvqa3Z5tE6YfvoPdiwerZUGYbjp/IqP4ZGiSmr3muUFTSjPg/LQ
iuwIP8oaOHt18kbTbRvZl6MN2QJlXsPXvubEesBWYBJ+Pl3zEIRKbqejw1GtcBlt/5kEsRTySRoN
ZS30nC9Dlae3WoFNYcaXFS77y4FD6tjWDe1DUVpJzYiNUJqILcsq/6Nk8+a19mxbewyblBVIPbnQ
EXd2nnzukCWvhjdpbKd7gpU/+FrvdWdWBXSyQssfFawoPprSaJTy93BVNNpGcjVuzVbXyyA5xii9
BcGM3I7kd8rl/Fw7PXoSFf9uoteQwBfsMobpiYuKVDE3UMf27PUihoa8GupuqI9hsvu9xc0z+BGE
DpQ9TyuBArypuf/tMAOCK/dUPV43owvZ50iJ7mReu8XD2oDN+MT5mI9Hi8ajZ4mgKAcBHCfxfocr
oHh4S0zXW3HT98BJfuoSkbJ59ASZEhL+nyQbYbiGSO8e8WhzxaiEEyBU9PkGfw2fG6ZqjIeepUps
GZTU3q31/+PhdU00QLPflKPRj5MI6wl4aoXwAPOy/aG3+vQ6GAP7x1PAHaIogATnmxgjC3LFMBY1
+/GZzhvd0XrLtrEd6noMYH3S01vgAYLTIUgG5lBgci7IoCOfzpXitOKwqJMUKFVGlALfmekUoZdH
AXGPZerVIK4Ullin0wV39yoIKIlx+6W9Pi6K4hAKdI2deMZx3BIPHoFm1t7RiLkCqQK9xqowh8OJ
RyQa/OHYBF1QNtZD/afCxJSoG5RGUUg/KClAq6i1bJ+1uN0phP+OFaUs1aMNS7ySpFLtPGEjSCse
vxLexWDEUvv/SRMR33K2yicGdwa7RZHDmfzxhAjyh9yjvr+OIAhR+EhNX6bZGIYbyxkfYPhP7Wq8
yJlVWquK7AwuDQhuHDXqfQQlbA4cnJ9fCkOM0Cb+aAJzaQZ/YanX3KprzwOVZaEQ+Js36C/xKeS1
1TW9gU3VYWEMOehNSQAQIbMQlJrOO3eOlDBoFX7xUdKqUi61798W0L4nBYZ/WGnGKc2mgB9d6I3U
m6q4rSel/UDyWFIWp0UEWhEqRUImVWNG9XXCGfVt2yAOXJI1n/yxpDIhwrpXh152UdLNMVWugKpP
4YdYPokn+Dt6u03EqVwySylXel1R+36nnJMShJFvETehXWNoF6MQUvih6zdg+CL+GiiZj7D1Kgto
AdI0LgGFfjrCxYh/ngPICcx6Wn4esjM3RruCM1cv0BYE/48v232t2Sri4DAVY7HdBlyB6xbObzpm
IgGNHbU5ISZxp6KOQ8mFWPS9rDVRLPnlSox5wJNlj3I0gPX0PEtL9sn0XClPxMwOxi1suEHI28Bd
m2ltOtt3WdAgfDlwAiWiwyja8IbV1/2QuUn1OTY56C9yhg2eGcDKm+RoHqZpAZ1Xmoznc24+Bbnm
/mwtzF7uWknCR7yjja+EyGHdF84p+xIekMajsRJVNfJf7vTkjFRSLxeY1q0dVMNIRNIyt/HYuVFl
uMq434VisGgbHF8HnCrbscFffMT5OJTiARjQmuzbugajgF/1WO769+qQocPdwXq7y7aXU8XE2fah
KQOytRjMFMGCwZfkdJCxoRhpJwAw6rta0iH8GPLHZ1qSvKCLFcUU4faxpv+y6O7wXBPB0k4EdBYq
E/eFELMNjxv+u0yOrRv2xWCvH7n6ZMl3Rplg0Y4VTF1z0iFJTewTCsVxJVGjLIFUkdEkHY2LAyOL
G3Om6RPMRmkKvZmtzY920g0wW2SxEEqMNIzbAQ4ucrxnfIsixshxhjkHH6AGrutqgpKEB0ofZM8l
Ub8fDqxhkBmFHxLhfblNAM70Q64semT9vsLMMkLe4x1lYBh+89m9dp0Al2TupyjPS7EpijX4PcfG
bDAgcNI8Iwf6bHqarrIetj9dRebQtKIMCwS0J41wrpO0i8TsPCZJHwj91cvQckWJ2nIuimMqk2kn
ROYjaXwZGJRyRmAhhz4V8xWACF1ClfpPUE/RKVe79hHAxkkm93oOZuEfO2P+HO8VMgMSvcK80Q96
wSeGKEiXJSkxvp3YN579/aE/0UazY+9f3ZnK6RiwirepwSaJidn1FDBx4BMzwD3rybBEofQEm+nJ
4ar3EdI9Ketzmfj9s6DcGnMzMNOIuQI0wJ1+jeGCZC9QWX580rP0zS83WjeYOhODJcNtTJpOJcbX
cVYRgLO7RZ35CXPkgpFRDz2BkB2Dk8G0Wlsv7ero10QinnNpKdeECcOVUFAfXq4oG+g+vVDXvNV4
AjzY3xabfQe82KOQ7L3HdmWth0avFYDReU+HgSDM01iK/XP8ACYAWqWViXSiBWShSP0+izqxet+a
1gdhBsCM4kFoP/+d6K2gtKfPz1FnH16H9VeMWPfmIQYD9IAceCma+6R8L7E20espr/0Zo96e0+D/
PaHDtIWJUQn38JnV3txwEAYaRWaib5VQ+fzG+k2y0xc7Kz8h8n8b/geLu8nc2A5W0HNYPfFV2uOp
heb8YnNPfvXX/J19xi5aR1M0d+SXx2Uxh1QB5yrn8w3Oygmn/iOBiSVs2SjnyC9aut8Ocx8Ediy7
q1uhfSwaVi7nun7sNfjAfHLVJ7ZunbszYL14FYqGMKss+DSGXiRIskbDSPaBwlfrAEgeBU9igLON
ByF8zrUgORhuw/FqsYlkCkvx47x9dYXMN9bT7qte5wPrHCi/mmRaUi7TYkU29hpE4HSMjf3FSpot
uctr7vAY/5ghQejKYuczupI1LjxhrcW9E90lhmsCqStbEsQD6FW8TH4ilUQ0vwPZEEGSbVYoG5XR
s5qSmQhuQaXMlkDGyNgV/mELTOZPCgy60aVEgOmOsrG2wGKmhH5/aFRLBJsh3iXg6jVWb+aM5QKV
xJGqJh/pB4a3VOTBIXEGQCiX0NeeXQ2iMuRrARu5m7XGb5e6jV4HQc4mySCzptSYCFIjRi6GOw/o
e0rieJXGcdPBISegRShu3hELvFytEJFCiNuNUzfIxFFgTL+P81ZqlNtCSXc7y5//WVhxFrX975ue
5zFFaFErQc6YqrGZO/+hWbWwkEha0c2nQgofwHH99ETIK7FpiGQFBwi93FfiEx8tMTmvUBHTY+Ne
lyTM9JACqFZvpHzboZfJ5U+MoKPrOyhGSW30kSKLW4xUdUoRKKvVE72xdy1yXPTmKT5aTe+jPCqz
SHYTKenarTmiAXOCtpv0UKxMlLnNgSdo0iyBvjnpUI0n3CKnDFKGK6FUriB+jqI0PMX0kK62HuIT
xY2IXtU8tsoq+S6RDP84sp21Rbx88qu9P/JRxdgcZdcg2c/ZR9OY7qys1jNiyrNXN1cWV7dZfhyQ
MK0SkRoFutzATvyG/imSn+Y9tjCRBkcODXxHMT0zjxVxV/bHII/MNONW+p1mVNJRp1d5Fs+NB/jZ
+vKLqztTcaznEjGqjARm7SaTGINqCiA+2p3LETEp5zEFJ900WB/hJwOUMfd0iZ3ltWAwIr7GqqFJ
tqoRKYYIfTtGQ3Q15CHOOlCdsCMHmwBDDy8Ai42klzWm44aXsEwI+XqzASwH355Amwxq2Zfl3Y0c
SjFeWq+Scf8tM+Wajeh7zXXc6V+oNh6c9Uryk5NITW9E8WcztE6e70jCPZowvRK6KAgUrexisCdY
oDOqyEODdQKLKZBOFuOQ3cYOj3NQFKckqjQ4VS+BgdZQiyG6r7MiNCKioN9dBoJARzd9IknkEbCT
C/hTZsT0cycxSFIuNTDDaouJq0WvX1EZ6sRyO8P5cPmnBk7I/Sq9fjVS0baYxlDR76yEe6/zytKW
r60CyiY74QPRjPhsQB8GyukZnD/xPMR6KoKOAa4M4vcee0v2x//XWhG6KzSghjpe0Z1MejL591mI
74JH2/cYcUX9xW/4lawSUhZLBheWN8iMyquDoZsYjfYl4ni1DjdqKuUjwcCEaJLrNd3ve6azaqVV
Ri87sq3oiOzhBmn8M9ibE3LT0MUtbSorJa5JZXyyXdU+DkVirMyCtuGzxR7CJxlWvmFoegoR8Jft
V5KgLXDUrVj74JY=
`protect end_protected
