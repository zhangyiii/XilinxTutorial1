`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57376)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMKRcNvzOG7grs/8lZMh3KNjoyD
IXsq0a+K7fwBVl18ZhaMVq+k2ZTg9lhurb4D+qNsORECx/TlShuAyJHIKPUj6Iho7/rBcVYF436t
BschO2PF87X14abVNYjpL91CiDTpOKrPtBKfg5+Lz2hIe1Bs1ooLtS/NXyKxPz4PTeOkvvb2+74b
GsrYMuFBhVRsbnXBpEGFyn7o0gnbYwPvI+rs0wWAsqkkHHqpkhXdpInN/2GIauHcpPLmykQ4mM3C
x0yc5+wqQ6/cuTkYmjZURAigJqYtVXEKWvz/LPBmTPDR/OkYrvY/1f7n0/8gOraj2rk4em1R0LL+
x5rliebLsBLJYQdZpnCMXYggUI3mNuW/Q5Td5tLBBMmT3q06AkVyVpqOBheQL+8Rxy2LdG5nvAzD
LgvMnIwcrhRg6452etuv2mxO1GXJweL+5yQvW/XvQVhDvPMVD2AFH4PGw1erpeoZGNZu2IJw/0Ab
L2aK0mi0gbc2s8O1WIzFpDWmWiFnQjnRnHClxcz+jjQcKggJuybEuHMInHtcfRWczsF/0Dnum9kP
8m8vHCPUZrgnBaO2Jz+BT7irdL5jW4U6vdgteMFHdttrUcbZInQO557zxl+G8rKCndK+ngB1lzC9
SDsCN0HyerjxrPx7d0pIpVIOopVC6h8MnjXapr7bkgkgWZkvQnjPBwhcv7KZGuNrHrfZG0ZOXC0T
5EH0nPwErBXNQurSKPrxbcJOXK+QrcGRH8IfyYs2cSgs8xNgPdDXlUaygEfudUHaiuyQNiiRCBgZ
81yqAxR3kBNsCQXRwJT9jNb4ST80OOzek8l/JQQRDyKTha5ZWvMxdGiKw5ZST3ZiNJCfPSSIBNs4
Xpg4qnEaK2YU6BsPq7w62Bz2hSR2VQAYXJiD8RXxCavS+Rrv3tabJoEC4gNmZ55ovLZoeCbm6DmQ
zAKIUrJvqAt9DYE5wlGK4TbaFFsmrEh8uMBCAO1GiZgu647deCmwJ1BPEQ1e6iysY1xMxjT+3BD7
hYvQGk43lyuuMly1vfhgWUcmU5ZL39xkeSbSPVK6p/H1H2Bp3asOQXBzsSUSEFbCpgGlCfdBfTEF
KLfWVTyLv1i814jVvAW+mAgCySeL8klTZnwNMYXH8aC9zoksL3rFiDTJeG8ugCXR3u67yVZpLtcy
2dl/MBnlJGTBIpi19Z6XcAD8T6k48/BOUvt1xX8hfKxIKHNqTS9gzMH3QKLmPZN3pdxfIYoRtvnp
gIFYNPkL0yEtMBXn2d6G9rEV9OepAye9j1CtGL58QAvDWfYY3d/a+0BPSGo8fgfbtV/9fRmpb46d
2rrmThX/V0GVAUX+UJpUi3yt2B8JIYGQirB7GyHa91yGNYATWBJeomRdoPtaSwWpNnFV3b9YHsEa
KJFKc2DBaPt2sxNVWRHtnfUzzK0YFwvk1lJTJjLRLwxbdVKevkfOreWHrKxK1foENQe8eQz7bMdn
tJaEL88DSlw0YyLrDF2vX4m1YYreZBSlz3LQElz37LE4AMx1YHYpaVPLdL7hkM09p1WUrllmdnzI
vS/reugN++q6m2KU9msKCyo4phpLvh7eLj+Js+IqX2OPae8TlAXt+VfpkPGJHtqkfD/Qn0fsZjuE
a7fs4+mbedGuBo2bU4Qy4gAH6dgViRxedPJySyQXl7QG+o9BvE3WJS5maP5l0Ru6MyiZ7iU4RU8H
1IWQjnavr8JZjMHYGOHLGk4J9uCBigB32sCX4TaaIBdyh9qTymZpFrTfAPqf+u2lOHLi0yXAwc7n
cr/c/iM92AU5ke2DuGqvi75WrwbSVabo7aW3UD8O/M2F0EdnGv/IXOHqgKp4cR2WBKalvKjQ39nF
xckRCm2ZHreb2nM8/s9niJH2ZDHnJ/y/xX2vLrXP+h1YkQfk7x0BjJ3Ty0jmdSVW0/mVuWNJZEI5
o7aOqExdpxGg8nE1HWL6CZ0a2E5X7TuM1RYJDePLnCMrUGUKRvTAIZp5P9/2OlWZsedghyhPC0K3
VreCmsWRWFclvcAF+F7sDvgBwrFDWpWSLOxPIK1XZhjvel2bNEsO24uvq6GOBV3m1RCattlf9the
0QcDlaAzEMeHiwnpnlTYZAx6YJ6maxpgPc1ndgqlwYaacq6dxSintAhZ97yYYL99jDxeyGKtr4gc
ghCj9iVCtv+MwVEq4uciNYQZu0xSbKJXW7PnSpWyv+fvkSgYEJKKcBo9bzbtpd4m8KESaxSsHJrh
g1WNSjhPZLctN1htXRd7+QVGp2sSt01bVUeG2Lha4aze1cUDNA6SSyfAcEbis8bQYIxhGkpjFO31
OQADFW+208ostfKgpeR0luKMPxpvdZJOoFhvjb5PkXTHmIuLY90EMPNVGtmyJ0GZf8lbokCZoO1U
a2KldDcNXKH/0BltyBFvik9Uj3Ze6rbmRozqoy/FEKXJHYR6+eMLo0NssrhE6uWHzdG6YHgTB9G0
WNe1PLqrNMIQJWlYMMo/+UtFszCsAGPF9v9E6w8C7zrlywH94SGMdP/RBbD2nFy55zVSyi2NujSX
T//jt/1+pOMhA97VyEjkXiKIIHmrPsQoSO6TckgPmLqGRGzyYr7KzUjZ65ol0uj9gcV07nsEK8i+
ZgwOIeCgok2RBJsnlhlPPZFZeK84+A03RMLAM/PxDBWYK6BoBeh8RHu9HmKZoremz76f1hp6ZF+t
tO3t2FKC2p2nmuSzsK2ZWbU8aAlqzhzzUkn91CnvG+bOwdmbwfWPdrmgx1gp8CVWzaZ+g4kN3YMD
4v+OGiguABqC7u2qRMgFXAsSlIcgQaGl/l0NRbGg73Nk0EWHCzxNQi9ED4r4qTsSwEsj9ki8QYDF
joQGUPizHz9F/vvwVT4Xk1fo+ohUD8eXcsHq+nQd3oM89lbmgkddACGlv4NfrnI5Z7UaZTnHOLtX
DO+QvGMDM6HiesFVX/sttNuHxzO/Fm5/0hMXZ5Os06XCdmAq8tpXb8/lJk0kOYwHjI+kotblabWb
oH1Ibfa2l0OrxLankgYydQ00RKFqo0RDmehKG1YyDvIMIMN8EAaQRwCI1K37AyxV3YyRnRjFV9d7
fdu1/2IWbnnpNh4lhq/5pOLSPe2iJe3gw7kPlL3l9wj+8yVzseqqZJWDcohzMadUz0/qZNSt7hV/
Jb/krODjsq81SB/aYWv9rXC3Q4JIyYrctfrpz4alNyRN5GZ5m95EXQL2OjKt+MT5fsXgQwmC1Fk2
AZsO1TaGo7qTpoEAgit6wipl3Wx3UO5jZZaNfm/Mez2VquVxgdLHWdVnRqVQgDGikGi2fXjUQxY8
XkjAAd7NZZjim+Nycwg7m3BdNB5TvpDzC9BHggiBeN29XD5joheP92C8PXfl6DmORibj6dG0kJh1
q/Sxyog21rdI22cCQIGrsS/L2K4m6ebdIaeuf+WhGYk4sfciYfV7LR92bgLtu55dAwaaY9rXWR9P
rN7+HqNDtbuPPEg8SkI7tSJrj2yX15sixa6eku1xm4xVLsGFndD4+j+I2GGx1vG0nD5kwaglqGQB
iA86rlrgPnAaDjg3kIaHBlMXEfmDbh63254zvbUWVdYaPSLDw7fBW6hQbTWnQcUe6q/Cyv58DkIf
hjp3jirWdui6PsT+2CS5BS71P0kO0Hv7a8xdRD7r/OV8SNPHq6Cz5GHk2wcI3EETXrSRebNbERR1
iNpi2+j36uCYmjo4jlM+ZfsqQEDGnkIQRPSsb/kont37EDK7pPlzUnPwU+h0v7QOKXSC5fggbqrx
eAfA37O+3+ONAHDzTW83WnmA4UjkZokL6JYLViGE9Nw9ZQPz3JGsgp47nMWq9LeXMFmHPZNqjVKf
d807A5L0/EOP4O1kQpODK8G/kpFzUzW4sPzyvdb28HVh1kJPPuuUkbC9yamtjFteKPSE5J+BW6Yq
by9quVP/YlezB9zg5i0VtoDA1DihIH430v5/849lX2RSe0gP9XTQbGHAgtgju/B012aRHMYoItX5
1UWEFVdTbrL286LxYUn9ajSc0D85RY2porGwOrgo8I4rgE64L6ntTppzBKSPt3zNjTADO5TwhEpp
FfG7lta41RW62+x7ulP+e5sMuKYcgKLAysAvrao4z3yLnZmsJF8rB9JHV8HglX1vp6DS2XW6vD72
fm+zIYYWcFrYKSFbSCZ+otTVBV/mkDfkzwZPbzvkfVTOomgRTsD+yaRgp+w2rtt9cUQn8ufYdSVG
p3ZjUtCYpLqKh+yS69e+BsD6VxahhHRcF1SPpMekBnMa8cZc/dOy2I0AycEgG8ZptSQNjmh+LrdY
J4VkZDOdn0WdTWqHmXZADwCNx28rexYM65b/ZN1QEdXimtF8NlvR1Ht/2eGLneBvHyxTsnwjbbG9
qM+QmlgRFm/4T5j7dCfLR/cyW2i09eo/+LGFmgZQ4JHhUgQUauWwKFj8rzVnbADZsrPe0BiP1Tg3
IsLszOKY92WXqMcwFE1J3K6tQGUfIcUcR0rIZyVzofXTVn+zmyxJO1vBgDbYho28ZMt/19MPkl+D
s6plVGWiASkh+ueJX+Uqhj24FkB0D/Owur5ITky+2SJEMqFX5AJdKkkfLujHxItNNHYvdt9OH47s
mhSnY1C1VbPE761EspLjqOxjpsilYHhe4Z4DNJu8H9TG5dMsXtZOWXy9XrU9S/ZM+PnIC4VwxJ0n
Da2ZC4YwgVNOnuXAE9cAj/q9B+OlIBvK5fMq3fdx84zMY3a3NqRzbXwXyXAg36ZVpkyNkejFUdRg
eCPt45+vJFPGH8rnq2Kfh+ll0BjE2riLHGw1EM+NxtH95apvztnZwsBqA1F47fDucPI90aobMxnY
C6AEWff5URnrbdadiyIMgFZiawo1yYRpIbZSEvboR/URlF605cq8lXEWClidRTRg7Qle/IqZknVB
mzviCxuKBrrjlQZIHhRayEEwztAeDY3+l46iRQCWAWFC+BaZiWH6GshQpj/0eOb3p+psjzbUdBVN
oaUyyPJO+6YkyhS8mE0tJdHIKgFwX8Rgis/fzjdoZysPu/ssUtFjkc/8qwf4J+tVeqsDBactJPtM
Yo0Rs84d243608zw4l8+GbPmTvm2FYfvx13XSDQlf8O3CEhBpbzrviQPRP1S9WQp9GrWKL2f2haN
9f2m4I2vfhDxups9rjKaLiYD3aHuCse1Z0Pg+D1hgKQx0Gi24xAfAVTLuNM4y9YUh21gSzzRVA/H
nj4CClgeBKtWCD9Pqbz7yuQyP7oxpKUwkqgDU7mzDq+fFivFH+NR6WZQziFoQDksKPtD+HvMqvkW
Ww+C/PM0V0TaYtMi+j1atr0bC06O6hTia2PJlywLfmaU8dl4SgzNArUbk3zxf1mcarIpivU+W+q6
VJGR9t8+aDDPXaLQTXjGkmXyesjY+GxoKKcf5Kn+o4M4zfdsp/TcOLzLhSsfKQ0byJL9bFu3Y/9/
KvIgPGRk4zUy+F297vOvBW6wZAhYhEbqRrb5A5rkRTSxYT8j5dzJI1S2JNX7wk3OOxGYLNuizKWj
KiLFS+PrHqCEa+p5HrL7HNu22B1j+WomeoIaBwaQB2hvK8vnWlRKQen1E7JezNnRV6ZKxhVjZOkK
uKFVj91MX+/90Q6AI8zOLJ+qvA1cRV89vZrkEmMrN7Rk4CVW1JDYuhuJ5pCywe+3W8IKg3G04s+P
ctrNfg7FKwbxJ/2a8wsTXy2GZQBsUpE5FnbTzbTURhw0Uzd/pybEPeSkbRpNgi378aLhdchPBZws
csj9gOVrzcDlAWmmOI1iRx5443Bv3SM2NeaDCt6d19Fujgh1r2RHCVt5gHCL8zw8Eq3EugmFQ789
N9c5D4clXFKawsdxVDto4FX1tX6ZoB1DkztATU2so0CGTtLzCsGtYwdayMk04mdcjDQKOqPWSSYz
vdreruZVLwLOnYElHQOrIf2RhFR9ARRk1+HAR8LwRkjn3HXs4Rq6fWR0M+G4MZAIgyuxFM6ybigk
wc2F28bSsKA+kT0Wvb5sf2aaDxpCCLS0aaMnzlh/GamhPn0IkxWgOJ2vW4MTy8SCBh5SmKGwbptH
ssXM6HiGrTUKhUDAHQfRrWIxgsY3f4z2dGWrj81b7dKuDmpYmHRdYL7oT8eztqIJlVjspnJI7bCf
dm7Xr5XOSFiXyDWcnusmUV/0YAK2Y0SI73LI6n3BhTi07dxINriPPhPxkUushihFUXueX+YaIAJw
F8CWi5DWjII81XYqLixEWNOECSCeMxZSy7d4X/2NlJgIlMyJfYXNciLLHsZnBDS2wlK9cZJdjkGJ
ta7LKB6HHLaskJMsyLAm9dsZ+C1FqwcuhFQ/TpfIMzZZUSPu8WnWu2Jwk02Y999vS5Y/lwzjPilF
6xUmR0pJq0pYxqcuFWebVSLGinzssEL6Atw37arYLAugl5pX7i0AF52coqHf2Fmc55Yhh9uVoWnr
BdcuwQTsHNuIKluceHL4LqkWREh6Rq2pjSz56wd+B0oZgBFIKOvhs/UB4Tw590nc9rZyRMgj76jK
sUVkoWg3QL7xBgBQL/cKt8x9El36Hy1f4SKc+8JC5Equ1qxnh55+1vcyKNkdNAABut2U3tVdwmao
4pXPwY1sC62PUVqrylRlyNAlw7+Rz5b4XMZk1mgA/Lyp1eYLsJGoOwk5FQXSlFUtij/EYHqPbxDe
mcrTFirejEhKolQmW74C2/9Sbgguh89zAehJkOnJ2zfBNidcErJYarEQd7lV9Unf3vT7QEpgT/mh
GSgZJ/oMt8y+uVXPeoN68A2FZltMkOGuQM2D6q0DfwWYSk8HSJ9/DYE+xN0bXwC8IlleFJgZGRJQ
zSVKukxAb8dPhT9lLyFECg4dPxFWHaI4G89nwaZg0oS75rLqsdrJFaG0To1gwu4RrUmFyhQY8lba
wvJ9MU5sqCT5ylFTbnRd2KLvJkM+iFZiFyqLNV7crySK0O9/xn75Yf3eDNxA80R7Pe3KE2ARzAzP
32waUZX2GaX9FCJAnUC5fvar5VK2AbXNg/01DmvU12ZdBrWHQoMScRDUXa57svpbzDUcqeYv8NUR
SjjnnRpkhnMjgjB8Eu3YhhEQQK+8X3g1h71ufN1zKqJiPL8oJHnF564hO2Pe4pWP6FEa4nRN7j2m
/WgjrjeJO+qhnTLC3Z42LJmBi9Z+LHR+AAcMk9ScxvQVvNpoABunQbLIxjP4TwsiXW2FjXcQz3Ve
+yBOyej7GSK1R/XD9c96YXlb3QqHC4eqSsaij7knrxkYP1XLJTCDHTsds9O+AtKxTe4Wb4B/y2rU
Amy0Bvn11uxI4ZqXKdhFkAscqZt1EqkMoBsEueGn38uEw6roLFVTYMwkIodzMHI4rOFESRW9vzCx
T6XOJJ2GVLDe1TATu0bzNNsyNfxngpaK3SF3rQkB4kMdd92Ep0Ofqz5clYACiFMnBbIjs1NTAtd3
hu48qG8V7DyLiPZYtgecIXmMxzqrlI4KB6iUaY0/F9cwaKLHO2L0rpgaZxQPmmfPXvXObQdFALb6
tuylW4V5rFgks94Cavn49GPamOYkgOxfY9OJ//oTx+PJ3gev1rnEkLN4VSCV56G3kXKXHlZvJHAV
MCWm9rRUr3lXa9CZ4TOnyIjtNAMslZu6BmmsJHiQFDVE0fS/0q1sCiSRAQ1QNT+4sznDdSozEKTO
yBe1kqzJkD81GTzVUZsrxf57UGFAsy4g/1FrToEV/Yk8eX6aIobNnlTW00YX4mYJZp6bGX+ByflC
ouLScYYLFs2nCAzJr1JkIpWjY+0Na5toRaCb7Bcb76nm6FeHfK6nBxygGBLK9eBaeNWZVIzX5J1N
JYKmdNtDepABVVetKj6RQJzoPhFVaewU3UMr6WavO56uNMBKrc/KhsMCRvhj4zRrxQs1yOmSk4vu
UIVqTxQQ0myuEgMhD0VwxmZMNu70ArGsXFhKlSadvjjci2j0MReT3bOSPynl+rLKDc4MHLT3eBXf
Yw721OitnhguPU4BJBR414JJg1J2Nni1W3I3YQg6fps+KF5t9wtzbteSDYRCF+q2zqH7aFjQTl5y
oPyJ6QJGKAOFseqHKZ7tMAYz3fT2aU0Bxhp/rEQ4GsgaOOx79reUYhK4pjpp5nZA9b8EoVWwigMD
Pbq1o0D4b/hDnlpKYabkjQAaeDp8gLOy2sIkQ6c9L4n1MmfKuPPUZQhHrtMeD/Ryjo7CrO2WA2rW
QvZ/osr8RtiCXP0tvejWVV4YjnlVSx26x6ElO37RH3CPgvy/8LFM7FLRvvNkAWQIrY/qC3JJdl3M
Vq8Ara3T7DAXRJ8cU2bgX194sXMszepZzySMtySLnf9aFVYwceGJV02lRNqs0gS0XAb0KUWzDjOD
cD915EdTlmcKtc8SDOS7p0hKuQMFIJxHhoRfwttT5mRXAMNV2OJrwjk/9WDPowUjdN4yrAApYB/E
3EAbNZmdEJoL01ohuW0vWn2DuffYRaZnBPbWqZyzKWgabRreRzNxUBUmHYinCGxPMwZBgqzvfNDR
CS5wENo3IBpZfIXNj9CBkhIV1fw8e/Adxu0+HySMnH+ftkYwHN4mnFFsbHHMU8/JEcrN8IT4eYoe
qEpM9GQQo0FcxVU1hm8P/hIofxS0DrUGKBU3VJnd1tOLtjRJ2mRu8/PGef6zrFG6y3ngvgZ27CHo
Iiy56Qr5BfnT8n9B0i0dV+yuERQDLwi2m35gOOFSqYGNhmLiNwx9OxVNFZJVsRxPJOuKcTQwCCI2
tB90OIzHbw8AWudtJQMqp/MqJsgZXOC08qYECx9q8nrGn+eT5wzmORHbX8ElCI7xuZ3fqsXq3AhB
fdvZ3z0pPiloLILVPi8HtewcIeEfn2HQH8biMR00zPcZ0mTUj6zR/kzL76ctbInYl4h/YKYIhcvv
d8TEpD1R4V/z7C/5LBAA/5AeD6vpEq6cRewhy7h1fyJBx7Vr4i9IbP0pVzwzpvJGtTMH7YMV482d
/OROh6snNVR7MDhnj3m2xdVPNXmEQ9A17WSmZgB7tuft6gviqpV3qRno89/T4AlVFsWskbOebVgy
HRIniXYpwykJRDyiMmSIcHyioeCA0ULUsuywGOREi5+lxMMeijv96z6t2tfF0G7kUWp0Jg1bKjNe
hBvJAs/YCjEDsgIWhdTSw4FyScW7nLQHp9XdQnE9aUnpVh1mpwrjvdiuG8bq7GbQoWF4pObNqyWe
TwSBk5BOI+VpCmTraoQQN5Dlrfjkh9wgJ3urk7UTupNuGiXbANXhUUsF0ezM8WDvZMvTiD+1Dk2Y
STDcDmwZ6KgUQt1gzz8OZ/JIqYSd+V53dkiDAQeJKAoirtv3gHhWgq1pgtPj7yDf3GGV0mdk/BbS
Rw4iFyaHfzx2yumVdO8UiOnGcW8Tsel36IV2kjnzft5KJPym2iIfSlVlf0Qs4sVzskHqpLiJG2wX
AG8ZE5QLCc7UUbfX3lFQXmEDwjm3Uzm3/rMtQBc04q0MW9xxRj48S3QHY7wYETnpzNs4xeI7ztV5
ime1yFzdncXnAwzryshydqMGfhHOeZChIcbXG1NYhtVlXBI3zg9lpp+gjnFYmmaoLLYMcSNfLQl/
xxvzT8POYvSSwzZWhYOpwG/Zyz5gD3ygtlsAG1slE+0BlZo+94GmSX5xUC6MNsr2GGPr4tqAX7v5
Uag8Fx+1KwuNhWPUlX1SCRYySzLxAM/Gv0bGrHQZb1KzmLDtqfMR0yEm373HWB+kBjfCkS3M2fLD
RhcLWCEutKj26GEDl8ShCagWsnTuI/15hASaJVUUDy2m0hlq2YU2xEfJoqxEN/9MIkVTg6wvM5KS
wcB46kYz3C0QhdAwqpiwwzefGonMket+avhv/QcimU2GnOkLLpA1WSCrkNHec9mO8p3qCtlFzy22
5oN2Z76zc9ixVvoJJX+UeDqmJfUNcE5YyA8u52+WESjYWODoMxXVQANUO2jS/zdvuScyn0MWu+dI
OrzFCt//TiizZrQK7SWIdhyGBQgGu6QfpVwm6Mq8Kr3NAR06QX+y+ix6XHOO23/hybxBr88KgfDl
tb4Hbw8oxocER4X6SwLirWGVlqBWHaP+1DNgjw255wK4w1YkV5u3/4lUcEIB6QRz27jWj3ZtEMKA
Rr/0AlD6d8hXCj2VlX9jNKvG66nkwkZTJSO5+cThlvYZQQmvnUXn+ixeaW10W/O5yIC3XgoDUetz
72FLfXKl/+9C9IqmD9PmeOT8O9z4rILflNOq69BhfgvhifxVoHzjFXOfi5jC7wJQc8AzzvBtHlYr
vbePJ+wbJNgvGIY+qsBGwRE9lt8rgDadGhtcoKm709ehZ8lVxk7H/tajAVEMMR0pgDzCaPvBdluk
w+JHffig9CWnABytZgldWLjDrYDHsrzgfrV79gM4SETXjjt7IisPHAclktfV4zmlwjAKVEgoyQUJ
CEnzcx5rrfWEWbh5N0REj1nQXDMN2Lkx6LNrJQZ8/COZmO0xdTS4Oesoeijny+qOxgqiAywd4Z3v
zS0fQ9ep1NbCgzNPNG8ec/YcVCaZSePHYCMiSqkq821/PUskaU1jHsa90/RRHuPxqWnZgcfk6IFt
IcxiG73bZR0wVVQLStvurMyjPTDnhes7rD5ItkKgUOYKXVbGFhjVo5HMSY6/Ix0TS8lmKedDIYZd
4yZjis8jgi60+GwObGJG2gbTiL8aTpA2wmJzNz4YpKlDi6PpB57xgkgzC70UiBZCDWnnN2/yKW2l
xE+wDE6baqJrJ+NnAO5lGlOursBFH1YJ48i7vUO0ua91SjNIwq6xahcmPGuMP19VbSjJ93/Q4Qhl
Dm93a6oKtC8FjPiaJtrzbm5SpGeWCf/rY6Wn0GWskhob10FNlK72F2eZXRWXztqkOu/NZmA8T49K
FiEJu3yuT7GolTdqwgXNxAaXuIUuFHQpFlbdcIAhfnaTvsIPDRu4IETeieKwqp4Q7da5/TLbfOEC
i3n3W2ZiPNPB0uTdPSb7WYQckT0fxXMCd70wHTF25p5kI7wD5AUtAOREoUkGVGJl0f65j398uC20
3gb2S6Da3iWNXX4p359P2fcuDyvrCZCcLoXviW9FjNvN/jounTkrDj/Kl0gD03Kbft+g/vthNsGI
PnDPw8NUVRdIXz8Dge2LF/5YyPqr7HS1d01hwukJ2IWYm70L96FGdU+ZC/7DxlIty/kKaXg1Qvh5
uv2O5E9RYffO/WBL4pGAO4Mfu4QJPOI8d1kgNvrn0eprfXCsTXPx2a4vDMSP60zcYs7Jm82FBffS
QIR5k6rn3agIws9NKHQqKlmmDrB9RKIkJr68OxBkWj02csPjxGDdylnt9MOWhUUGyWiB0CZMQWXZ
74D6CNebxtphhXT0CAneLBEE5iHm5OU/TbElgyKj3KIpJeBEfvB6WQb5OVo50xdsYxmp6FCcWnUg
6cVnl9SpJqib77ylKS9QnRj2dm5bo/Il3/0zNxcRt/onqyYoUZAmxC2oAwmwFcKQ05sX1/r/cz3W
55bdBSxiqnfN0zCGckZtB1W9ApOsv/yGtnropYyBgN3hGZPGHOYSNB0wQzK5G8NjRIisw5pN/8r4
Z6LN/dD51eM2fhI1VrHNsUiVLZkV/Tk1LGlCNV0Hj77Q3ggo5YmYiX3jvBXEKNI6NopYJ744V26S
s/61if+/IXgkx37kg5h+IOAeD4D41hWkDJ8FJMVldgGhcLdFIUwaeJGAmQyBvTLzWynhNlqAEDCe
PZQ+W/pFjjsiXBdE7i8mCqp0Xyfi0auMYczfl4yLoRWq8lyO/Cbtp6E165sOcR9kdoowcAiWaxA2
jYOHfJXTDyevd7EDcLF+lhOL86EmrCcjyAWJ176kOOwoVfZedpinpvus9pYyPg229P640G5U72iR
gyAHlcOn6hjOU2tbppQUqpn5ZJahNwXUIVuPXzmByoHerYuxQxQMLuCo0rT4Zq26twDFptozkp/9
ixBzJFFy2Uws6S5LPyleCFx/sxcdav4D/OPmITwQU7GOVFTOhArqbjHAtZTUgjtm13UM36TJJ8qy
GMr/TwodiYyZW0G8NcbNNImcMs7rjB5geGOR61AP6xW3EtAWPJfIiyeLOSKeyzhi3iskNJ8wLdm9
4vZ8rV9G6DOGsa2Gqz0IJVxXPnd+YbSDxfT6EFMymfLMZShRc/qbDGeiepyWIAMwrhZ0lsfdjfYM
CzZil9faVv2BGBxA/RkGltUv/y56ovA3rrVxLV4fgF5ORpAG61AVMsZpTTNfILiWHRSdUCdSH7ak
rxlKzOsVdFPeDtThTNG+A/GDRGmJYK+F/d0sAt1htv28ka3mvQdGfBiZAIGQQwCHWNMwyLEfdMCX
gUdkJ+q+r3rKHuvUcUxPwvMgFOBNeXEEPwRs3UA+pHbE8Bv9p7+JU9mW62a8Vq2qM9DUGPl60JCa
yokr52c0NbWZvlvwtLqZBxm/qgLBReX0bPyVjuXYX/vjcAxlOma0sryCVmhUh32TIOs/BOq1Sygd
ojlxQesZDWO22pFBy2zu10o86U27N3B18EtxkCmDvOuHbQwzgDlfAcwC2lrK+cbJh0+QXp7md8wp
r6Fau7Nr0bJkgHbR8ajyMvVycxd3dAqQbi9e95SJSqeOb5DF6J9rTNF4U1DKBvGR8E9pUcDPk0Ox
xxqwLcCUhTTeRGix3Bs6IVsUWflvd5jWScPOqMTOwPLxfEM/acsHVzSJ2aLyI4bnLuqPymdwkOUo
wm91qTgTzfoHOE6a6FzC9V/k3Qc0BEBpCTGbVUaDwDlDv/X5Dg/6j3l7r1EEp0Zc9m+Ewjp0U8vu
Tqn09NXAOpFh6XX0ioYLv2eQiJUJfsW36iW4zlZf1jw4zWd/jp4/ITqjK2Qoc2Cy15+c1r4+cLOa
jRTDwy0B+21HcfAq7Lthi8mBYUudZn0vd96gIGqU3C7iNWHYW0fCP8ubjYN+WdIV7QUfvkIQb45F
ATr/dysDzAZ1ryr1/Q3jw2Ut12DQVeJMpu72jGbUR4Z1zWV5Be3P4Ca9iOCqaZ7GDnJu+jqv/++B
slGj0HHOX+Ylet+YmmaYNjrZ6ZkGu3mVi58bWFnx4RsGKl38AVuysw8CN2GPReiZA+0g9A8P/k05
mp/gWhk3y0ni52eaoylpCzSAQ+8gSOfcKXJQyFoTVBXjZwLaXHcINJmyCZpvwGnp36LcGdGAOyH3
v6DhUnHv2RvRku3J3pw+wqyKujHtDKXliki5t9Uk8Rk3bQzzo96N9wSGYO5Z7JPAY2TjQRnkZdD6
ZDNJETRr+bOAoslaHsktsmzdY/RayAREee2OtU0GI8EF9l34boXsE3YJK+xHIXLLzPDOAifRAhPb
fPKlPzFBH61DdU0cNj6vvO6A7iuWlaiM7Pnfl5JPN1SCMhPQxdcOCsveifYfi823gKWWcEjIeTuV
m2JgigjEtmKPlX566qtGcGkUu+g3Mn/MuOf+4SnRp0w/Et9ocl7YPlT8B99p9ZjJT8VyA3t9nPmO
g9T54esC4GkuqyLpIEskatIcjScrPe94uaMXBaHxYiK6YIpJkWR88RC0tn19HzMX4f9kh3d1AHPY
HmxSe4r7k7Gpt5tO9TvdApyJw7CJzxRCgiUF8ftprdf0el5lmMZjz8oTriFTV0AON31jgnaYFaHg
cpxtx/mOW/oLa3W5IB71rRVty+uD9qQdWkQXD2rnf5tpdtakknALRNvI2zUuU6yRF6QzuwPohbUo
YCgdskUPAmXw33hOEUbtU+mqh5PH6nhaRWpYiXZMKvAZURRNhWvVpFoUov8xP36a2RMF8D8M/vqr
grnsxrBqvWsaOl+dYbqOhy+6QQQSMDF/jO0L9VBGHZHFehh2h3E65ZI+jq2vogAyzVvCWT2nNH8O
Kb/TQcTHyOVso7Rt6VHrLIlbGUONphEV9ESZtmO3UIdL6x2vQhJPtrVUL8MeeNnnvt6FS9DLKk6b
LqsYl8eKCty18T+FIyr8HCaAloVBSJcTK6xzHcEI6epaYupvxlDWv7kgVwIDJJS+QSGjgJsf0CCR
sJAUrkv2T/vcx19z+/0QkRpb1Ira/wUofOHSu5yX67a7uc9dBCkXOFPJUl2R/AdCbYhYligkXhtf
zcosTbJ6pJFePbRyKTi6NijJnjmk9Q1VIKAgFZFWmlpN9cCDkxoR8noCPOLCbBT0JGYd2yhsQ76t
zRA6sdclhSaO9jZWgtChiLJW/XtZ2WQOc8MYbG1Kwt0dk9wgDkGQ4i5mxSPmIhTt+9rT8w1mNMbP
3t1UrrdGFEJzlT5es8odc2fxJ7VeVbKihanFFCqhDkBFLi2YcFanf0QF0lMsY2OQJejLT9XzVPjd
6Z8diwdnF8NJlwqptMg/qDZwtG1FeLyKArjia10BRsL6SXJbEhEmeppuUB0zbeS6SA6zHx+kIiix
4Pz5jyPFZQUr+eyjLj7kG5TuJ3Izv7zZ3elpT131Ez52PwhHEzhONozMODYxS1OGnAqklr2djri7
pGFVihtIMkb+ckt5IGFiE7g9AK2U1AYiv81Rukd8w8sYnaiD2BoAHic/+AtZGPrplz9ZFy2ssrB1
a/y9hKXS0+fZQyC6xWh9yNzrp94wq1Ngellt0etwQf1S2tqybLFr4GtZbLTREXvcB/8on2+j0y9m
W9McXseuWRtVVFkNMmvSJHSp2J/yIsjPCyCGtLeamu+9YYVGOO6AksltEVeXG8DGs1X0rOxGJiN4
zpxvQ/jF6IvbK0xic4Eq+g0BPm0l4TvEtNd+HY76clQ8r16vUt9BCAWTVjG21NNqHpeQWGak6gGS
l60pH43BUtbPLJvN+ChXBMTz+H21cwkaDax/PMeu2wZusP+7UAkb2cMkUm8dIO0CJsy3JJzolLCG
GKvoFkF/F3IvtfjniNs5mZ6kZrlwWF93oqqZ2/fI4XEo8/cRpGBxgeg91/5JGump824nIC4F9PrL
2zB+Y5hdPxKttzXcnBU0r0N2uRMbx/OIJujCu6sRfteoMd8OmvrZ/quf4Qrw1V510sgpjohlYGrD
T3sysdfmj2dE/b/hJLBaaHuNqepkI2KfXZteeC64mxnjPSp94UPO2yVAXDhymPqBWAnmRXqWUsf3
RywQTpJ/k+TjIpuEhUWxxMHgWyKHB0DMnwJhnSaJkWFbvxLqBve4MqTBlfjx5Ugr6lV6LyVW4F5G
SrtJ0CSHg1zxItwjsU8frm3GA2DSdTuQRrhxMIsS4/7O2n3vwubZ+ciPHauqK21enP+CSBKXA5wk
8KVmjFIsVZN4sdg7KySyK45s+OIqBfgUkZRMCMh53W+y/mHSLrLfM/22wTuSzHxzrtOr9kH3JUYV
MH89jSwOnACMMj3tpAPaqjTeflMCmQ2RvkiXImfZmKeBoXUuI+JCBEQxlOZwUn62LTiRsPSrQKG/
GFN2V6P59sikkciMJYNvVOWNy9HH2PExDO37ziYdUgfTrK9iPq0/7n3fCytJsB+F4h0/v5W0tUSN
4PCwqLbvy7sILxbG45A6sPUlqED83FWxGscV6HXXv+rCsiANhr6iCzgcPZC5wODVL6MRziozGyIJ
P9FPI+81ukXsuFwjvDmRHeBdfiZN2GciS4y5EnqJRsEnPf4p3UUqa5t7g7MDqMZ4TNXlNfHm3hNk
wHrMqSN4B4xZzSAaoi8D1mFvTtoJMvk/mUIaZaXC8XKZqk9tU7u1bTJQ50jmv5le9JUFggQH+cOO
0y+7MRGBULWVMtfavh2HiDg6gGXfEfS7KuiuQ+M5I+1sZzyNMDRLBbNnoznAt6XbXehrNu48xq56
bP65dUYLOqubaHiAVCFUR7OEiVJlXhEWZ6q3w+b30NutMkb/7ckn8g2K2U2+kOIKTLRnsIKwXnYy
uYuFne1mwhjIPURhUezrRzS1IZH2Y95jEXqDoFIefdr3FecyurWJcEqREUfqtBLI1hpBftOYI94X
EMrnC7jbsQusclECaPgelgIn2ySblAUn8DIYzAPK48uJVtwT1Vpcc/2+TGbcBG5jdqGKyL7a12dC
LjV+bBtUMBxFGfMByVt1XGiXCoHRhm0DGInugQ7aK5CMeS3wtpoQ87kb+BbqDtr9b/yuehkJK76O
uwiy7t3Y2E9ab+ngX1S6zqEhPyyF57CChV+MItzzu4wpzw4RMkw6Dr6+C2SrXjFDfJ7LN4Eo3QDp
ILeqDj/qtVSW0PsMgq3kyJ0Bt4RLqrU8ZQ65C7wgOMmwDJdVd3lgQfmHX+ctaCHcurUgZ5Fa3Dvs
oxbb4PJF7DrVKk6K7z9QpDQeqz6RGaj1lJGFPobjl1LeAlIbSwWk07mwmliyKf+kt92yy4YNTkeK
C7nh9BcbMHOSbl8IFfzm/NWCm3c7X4g+09l4Pmwwbt2SsPpSA80qMssANxc8jj2gR6lJcJ929OAY
fyeMlKqZfn+sJzKi/TI8y3YiCA0zQi6Uyp/fCywzq+KR9mutwysFCSSTKS1WizfrSKPu19dCwqUx
xj9ispBpz3oFQ1Z1FHbHhG+vLG0zPfr9kVOGuAK30KhqwMggWJZq5GhLg2XO1dWzDsFafYR6tSG3
X3rhMSOcfN6yE2uZjxFhrtTVTmbj6DtbOwlcFWN8rykiTI3NAV3QzSfZfL07xcnCvfPg9bU22hDK
LKw7iF5NnjWd11R/MZeT4bQlgxtV5Yoqx3hgLf89i7CWU/VjYj5vvQGGnTawHpsNJhIOf9yFci3k
kKVG/MMUced2cerx1qGjRRczIDGF9lINBtDvim8yaSOGyOxyTyPp0eXjTuU4VaHotounaDUfNtlu
oc4An+6qA24ZVpmHlL2wjpVvWnbmgDz5ULDCluc20bne+qg3BGOjf0ZGNnApPfCehqpnDIzhYNws
kO1MdI4S2dz6j8AfK1ismhhE/H8dO+SNAQonToAGVMdfqyat8GIPIzUILWbgitsboc7OJQCev5Ao
Oxuv/ohCpYshHS07U+5EgPTVqzCzJqQAwtVlWmIcq9VPJ5b0mBBiVMp3d4PeMjuACPOy6sBWoqqu
d5/Oraf51uY0qpZXkKjmgAvqOBEncB1AvxcX1UaQf/0+UVsh3UeoZCpoPH7+XISsEFN+4wRI4QWX
DyHtbdTfO9s2VhiT23OqfCtmEewPIW/jwnll6nyVv+QqtjqI99j7jntWxf0k5VTJlbU7eKP/Tbgh
UEJlLUH4gzhWS5lJHkIznA3wSmVo1lAQZWs9kHwgKhbJQ1UM9JqRg+P/fBYN5LBwPyvAVyu6X4rA
YoweVhJWyvt7BqUwlaXmQx6b+8yovTWH7fdukXF6LdqvLZ/z4ocYUrtVGuckYqjwqhZoo0YhLHWo
YyA8RUGofOygAO6jFAT5wyWaDkbDXtyFSecP7C4fpCia8S8aevM7/W2xd3SAcG4Jy9p8zrArcWCE
KnAOLve/24vNWsX6lcAiU+q6n8tCGa4/Smvz672yT+B04m6Q6TKRP1xB/4ri7ujj+Si7X6KGEtVL
RQ4SOv3VFzFJFJyD+9keZzvRFlWygc8cXINzCat5txD6ENEBjk1zpzEI7FHnCRhAUs+bsvjjswI0
YCcM0HIC3dvaDknt3dQnjZ8obYqGF/ZaXq/kiYu0tW+3Z0f4pnsdhHi5bR7AqUeo056U91vU26wp
WRx18I4SKfVpiG33PBWe3nmQWRiOmWS21f6qJ8qFheUdaRUX29xgrbmy8Vuc1SAvVX4EQ6DvsiNd
/gun2xRAWAkg9TD32FiBP5cM89Kg1LVDKPWks//AXCYkbiFs4f9Aq9WxEyvS2yrPlwH1cY/T7RLg
ghA4mo9oMZrQlble94ZrHU0x7BDuQqWM7oJcqbyve+mkraQu30LE5LKbKFiQsLkBNq4fc1L4++gm
QKK2r8zC5Ho6xbVJ4RyAFc0FQ0QaX6oiA36epuIUSLFBVExGU6LR2gAfI1Z2U/+qlX9txowf9Y53
LMEBd/RhzidcI2BadfNNnjOrVg0a3spcIciRUf1OdowkPXqeMF1wnsOP8PMkM7kkD8zaoK7xZxai
GVCmQzFpGKf5Zmu6xEm3j77FRlzt/GP24tkI4QSLibX6Hg6DQo2VD91UD8txhzJWlaS01ixq+57b
pkaS+779UHSLqDFGX9fsW65JOfAnfwedHhLsWJeGKkyB8qSktmsIT4f3tux0zJlEZaJrZke65b65
exet97G0wpYE9O5dHN7Dk2B6+PcgJERdHHWkyOW1p6WwdkZee+cDMGq7zB2aiqEitjndjl1z5cr1
0RMI4m0GNtfpfXgNXefTVVMfv1KQPg7S+5WP6Oq8EhEOOwMSwvVnuh3V005fBO8jONzLqnAl2qJo
+9KUvMcqQLXRkRriSMRBVr8LmWEVHixI63aaVMeLrbvBx3FHYHqrXYXspELlLnFBdLV+SH7SXphw
MduNZnYnLALgo9/9sPggBfC9/lr4E73YfHUG88x3iyA14Z8t31jnkw5nk8cuy964WenEPBqzcRqK
zCXp34NjILnN3lXurqcOU1Ym3JpMXvqwjghBJL+Nurlvr8cqvCk+NiCYDCFhDxQqnw4S78IEWodO
7QLZrBkWjsyslBn9tt7UbN7CAr74UeBxFADdybe5hqGLEDGzkXl7oANI2l8qYpIWTESNoFi56O/E
UgeuKxsFHfN37Ef5RItULS5JdofcIEBkfHAXbPo5qvUQ5UaT1xJ8g1MHuWmj1nOJZbV6bfvYB0HM
MG7Eu5q/sXUW5FfuGa7F0xzSQ3hqgGVkSt+wQKwKqNrGcT5LShunJllFCu7kbmymQsQOoRltG0P6
hDOr2bCbxtFHS/oV+yXjbJuRi7Hn70uMcpcS6uyryC4QVX/Lr+sQM1sHHtfyxWO82AH0vg+kn8I7
HR4oaiY4Kz+r90Rf04h/y9xbsp6jrlXjmwCotFaBEfIeQ/BpJXcjgINpkeQ0V/2WPfd7NJjfZkXt
6Ppr44PggDoQyvahMbIdHhzA02CXJ0KVugW96kSVhp95UP6R5ETSouU0HX/S1XvL5vkyHbJBeXRZ
hc1GnuP90YbuSCbVSP5y4F5mOX3Hr/u2sYt6P32eSEKdXA/X/KXY//RtM3TDoyJUKAep1UjtaNzB
IeRp04hLPIjvM2RjbVjQ15SydeEwOuI3imu05OrTgETUuvHGB8FbiE6TOelJhi1JIT1pTPrDvNRR
+oIGPy1EhEEyX/Z8GtYeFcv9JDzxDIvFQfkM1dfz/9YQ985HBBlG4NTp4U5q3dGHbUXw7Eq44xp3
+PAcGLTY5vV7L6Y4zmEA3tTjZX2K3dBXlEJeFKoiN27u8pWy3vyf6qxKwRqoiWceXx43UrClJlLj
hT/7KHfolWWZ4nsJSOf5mMYQMM2eDwEE5i4yLlC6cSZugWcYfwepJDOHQwJADqu6lcLDNkzWQ0bH
wafRFfcFzM2hnr08oAuKKXeFrsnAAWg6PN8TMJQRfldh54HUSwz2XhC5KTj6eQufvV6td0NqvEun
bULB0jjjXV0Z2PFSsj0wUWP7eqi+1QgkwDVNZWpwPe+CJUzEcBDS1Dih4xqY0AT0wbYfzyis4cTV
4NdLMNEtuLU9K+/sWyvsilA0HKrB84kfpuhGRfCcm11+00IBihhnMoWEpFr+ZoMBvPw3bv9M9ueF
fzSTNVfJY2SwlkNhXU4KLoRNx5EOl17cCTAQnQAamX3W//MmquUI2YVeccwRzaIRMP2ZB0BYtxpt
2yX2r4wPrj04plzBCZvTyxhf/qxEpCZv2xzaYkSZ6guozgLJTVqFaOkA3PvszcZ1uLE9FogZO8U3
L9CfkupoANUvYIhZKocKVcFx3rIEON18FtsOBskizpAD0i/Wh+AKXLCWDmKwxnz2y/pso0TSCcUX
VsWMmuTQ5tirqe6V8PWbTP7jkmovS+tcU4FbgddM0e5KzKmKkD8UopbUxhVB6SH4iEI/onWZnKfM
eYD3TPTjC8gjMHYvG/QmWJ7mXkQNmQA8ouWnK0O3E0YUxuMqn/RXiuUCbW7r8PeVQ++eKES8BvIl
3sIRJqtjxMW7M/52rHFIdfqnrZplByMSy1zsjU8KNHqvBryVTgK4F9vmAorbr2GgQ9PUCE0UFK6A
gn3tPIYU5gMsi4F1iYnHyEiop/yStE+y5HBKT0PJsKoved6gD0tzBehwFpy8znAScmxrvjdrRDG9
3YWRkkwVinaRqHZwmhJY94GL46G2rGycEPx48zjpsm/4bjuwWkHPvXoFjfQim+G6aBaBLVos/zJ2
9e9Df3iUdPo779CyScbuIMt7iRhmOlyP+sCxZbU9Wlw19T11upcZ0spTwnDwbXQdWum807KsY1Fd
q1ifI8crJltt1QQ7U3XVMl7rIAFp9AqPl+2d/MqwT3HtVSRHrnhS9HCUVjjy19u+d1znExiM4UcX
nfOE0LOUQrdicx1Ecs0i2M6T9wYX2autXGkZ+Ue3r6SmeSBJugdEWkVapXzV/f4mBusIjT5+hKjY
MKhek34ALlr1ZoVD40Bj06s4iaCBbfUdW4m1j6E+YJxTixe4qClZDVN8Du8yruYFfsFc9OcPt/ux
0O2e+HJrj25m2GG/Dz15jMskuS9T86jRCE0KXuPAgV4qxvO6TjNYHGhATyOU6ZffTkvz3blIsijW
RWm99H/we1jIysl2wqvVVIZgmH6E1UuMNXXJL53YZ/sk7DuBhs+q70OHd/OaZ+9KUA/AA0B69SpY
/T2YJtmK2fzs3Wemqggx6YuzYZhFNHDYl4WTVBAe+DvXivUWEEG3MvFsGh7w04N6a52zHeSNieRZ
1f4cUsNpwmCU/icABQvvUvM2duwzSoDeLE6cjY/aViK9jn44JFs5qwe5Wg05bxeo3ktloaGxF/Ae
CRB2S4TysjiqXMtLoi3DzPzPCocSPWVTyQ5Yi5IdOnv2QVhGKUGgzVkUGBOLtjCPTApxCchQzXs/
6xyGOYhlj14jWnL8j5meIHXqZLRlrSteeL/PcLuImxVZR9rWCsC9Dk9CzvAmehkskJVuDxs4M+bD
QjBVw5bmeB1T6aQPhVT4lJx5kevMj7tczrrMr4Go1aWRd8/QhoJqg+bMWD9mQ3SZjIiKi0crQT9p
hEsa59KFDHKEHVx+zqVSN+KxEtM8btUY1pDaHkvKT0pI9Mm8vmw714H3JvKsTwnrDilFbo6HPm30
AJw3xIDuCBOiDGPKnJR1WIHS+g+9qtbulYp+QFLBKgcqdIaQboPolKfr2dI0X/WCRmj+2yUcPyDm
c30QKUiitVmJliCJa1g3ZHIvP4kZbQO6DYUvPoAQ+Ah+ViVzpvUdJtjgSUmvuURVrnN5UFcD4ieT
pPf16X5C7Goc9iGQNnKQ+R9XVj3WC0aFldOinyf+m2Lc+Wfc9vJmcz60RyCa4OSsVKeVC0esD9Ea
kQJwn3OZ5/asHogfrIze3avQDf9QY074qvAnNpIV+Kjb+Ci3dd388RkfH1sulKFe8WHEGWMG6qa2
qQpfkoySgUFghQ4V79M3CmmNkpR+VZWLAYfFLOQypBPI/DF4EleycRgreWtrl2g/jFiFiZMT8dX/
YjG7obP8UXcrfyzcwww5QqgOjHlZaUiv540wT6GNdYjfIhODfNhsJv/ylqN75rOdb4d5Un2ZwbYy
kTmsU59WyFOomz1oIPf7FApYX3HYdrf9lxE8wadkO7dfoBTzyi4s403Vww5iM/bzLL8T3v2d5Jqd
iNZItGN1Jv0DkUr7lW8MWehlr6oNeZ1sPPfSnZ5rnfEnxmtI383X9QwnIX2jYyzsXn+RfOcBZsxS
S/yGQjSyO8CM0o/lpKCItHp6wghh//MurISTUU23bEfFtK50JfruKz8svddIqmQWaJ9atmF0K8B7
7mYQZUVCq3vG9WnUSRts+5IkxlSqbNnWtYR4puDL2MQlZ+2iETtlBwKIGCXjt23Vk5gLMJQ6WRY8
vVoRwPE38ogmK8hM2gv+0zJ3B4Ys+sJjM/JSkMhXZqBQALun5vNgZRMbLhrbaxR9b89uu/Hhg9Hx
0yDbm2WqOoWjNLK0Dp8Li0bOsLBA8iSzOOYn/+CWa/trQW6QmjrzDf1KrUJUGSdbgc45Ryhcfb99
JZmQEbj5jJqIr9ph5TVt9t7GZ4IkpO1OUO5VRqlKDUNjKhqLPkRI3m3abcyi4pnuRUS21Te96OFY
RAB+WLBqbuddq6IK170SuN6qZiF6wUFQnFM5H46MMaZO6H++oZFjBhKdlTvJZLIumWIIC//lQ46A
9n9lcQOun3hAxswJtQotINTKqKDt/qbVRmmrL8UlSdzEMLZr7//iemdeOTnegjgiwqMxmvNXT16q
0cEg1uxKkO7Z1ItmsHWGZEvTuokypY/tjeq1ofi5CprH305rD8dXYKx/XA/rjqe4PNSVomT99voC
rteWjgAiSvD92Nj8PalCeUizJ04AwjUdondYQjwkyG3UNFAGaChiEnTPTfCnCLTecUFAQihtucsG
6PQJ1o4iO7w4FvBVXuVnr/xhBgG02UYyMnu8Bhozluk9vLTNgxkPGB05/ZyXqpf7JzI2+CYHjQoA
yxmKzK2R2WKAbZTlCnog8x68NUJtkG9qlHx0g3jblbWKZvH8aHa0uNiPnY/dStTMGYPF7HOcQylI
kfuqrlLOifjyj8zO0Yl/B1QaTov8C97FJjywIqgG4l19bCw5rBlyNVXn/DMsFhRx8Oe7DyCWhOl4
T67OD27XSjIKUgqpAPa9OZucSbV49SCJzG+cP/xZ0vgnER4QQPegFYeAXVLDSYJRGaiQfVUO1lfT
PmFNpRW1oNy2Xjq/HQfdgp/vqffz6cIUSY2MbfWkT5a5hwzzDYyVjDCq5Dsa2H0cYPt+6VDcyWe7
gKnKCqMSChxN/805WPNqaqc2XB8tcLCnXLGhoATylh4R0zPc7F95V6lzsq8BJl6J74uo2ck8/5a/
pSuJLz64k0gOr4VOUdEJ8s7iViyJTcwR43HK04KuwTeLMu0RNsXX5ehX5OgWJ2B2qTDUVrBCgGtD
23itOhoa3xBj6E5o1acSTeuY5ZsqVKDjwj8151v2TvRXJz83cwcFMNQjk83GpSA23SbR4xyQ7euX
Mmuy4bNpH9D6wzEgzRA1FeOd5BkPitafz/sQG0MyRV99b1PXODcJMisP0BojZazSFjxRtHZbVFEq
HPx7KuXpU+1CGMqT88Cd4JYIb5HromihrU0ECouv2wo1Lqew6vOasw5oc7aPhndEoxkX8aSpEc3M
BpAum+gLvWLK374Yw42114TEW/s4Vq/agVzROwv0V6X2mDuLwKjTL5efmRPMbzlov6vunQ4YpTUq
EMoo8wPNw4RM+ubzn2PwzEBNogNL4kyljj2Gjxc3GKN2ZbX2wRqOHoEYUGhnavOEIhGRbkj8Nd8W
6Q0eE3aDF14Nl7llK3+oXA1MI8Vy1QG1MuSlGEjhHNU+wBTxX6jrU1D/MsQdA4Mtc0sM2IY14EF6
ur8kTK771a7cNg5Oh1/X6AkGwLLeU0lEf2uIpmFWKykHiYx78M0Iufk18qRIjlasHnxJlhY8Wzhi
PdUALQ1QH5JSZs4/ZNV62uuSc/GY87jefzH4re0Lf/m1iDRI9tX7x4AzHUEKblctIzQVwoKCrpdQ
2VkfwJO0y6OVdeKQC0YQ3N/6BB7pGVZl/XwFdJmyH/a4FKWQLeTw38Y4HQWLd5ddGsr4+2fFY0vR
PeG/KTbdKtYqCdStGljNt5LmzlbD/l9uExPMmGUEktRTbYTcoxZsEz1dD9q81GlkbTglAdO0azTa
y23KA4LCkp8YoRswf55/Yij53wcw8GHTcr35OONw3Fc4147dLt6ucgkJnwGWh0KeD+FKTXdmF7Bc
2Ul9FkvCHnf4Lm/RO9SIBztfqJYrdii3agKaAPK2PPl/D/j/LkDKC3mDqXb747dXkLG/qqKUA1Iu
+cP9uKPo9AdD2xj71bwl5nLUH1y6BK0o4UNN7djhDfWXRQeZgM6XMtr1L6y/iiLKxJ9dX8eOqyRY
lRERpu3XmfsB16E6QAOOZu8FsX/5aswEsYQQgPtChRdPgIvsoOD7pAvjlR3SOj2DtPCPfrHkmom+
mJWXybxpYiLT0I6phCcbsLahUBGgiUAYasaeLahgJIf2CUCrucEXli7HK92XWgWnAaVy84iAMJM7
rlJa0EzFS4K0Wn4bEXGdxwXKF1YDWXKlAP2lfwQypxDVuTttHKLYR/WMACkkukWG1hnCosPA/F9H
Xas4W82VEJ4KVdCW8+7dLDCpXe6+3ycTKWJKvBSlkOYORYtrp/WoCZbLbOl+IYr5K3RjazLoYN5G
ym5TqNARi5IbplCMmm8O1ONOM9PvjSwyhz0Dd/U1ZHxQHeThSxMgWV56FoN8HQH4MKAXDecVncgQ
Wg4XA34BXECfzLqO0RbGJKX8w8+x+K0rgnwPlMPKbfSrdCgfCIPrrzj+S7/8M+S8TZEQ9Bww2DmV
E/QvcUaD/zdDwrEejiepZeNmu0fvD2zck1nYVkOIDmD6UKoV1JW/URNjZj4gqGmIRQ1EuP9UUn2v
ituUbSfpBPTPIwVrsuoJHb+4n4bMmT44cArKPqpYYewnAObgyd/+jPMOxb0f6Tc4LF05SkkKFXj0
RNmrMQBL/a16wkPJf1vtlzPh4epcdlETXn1+jO0Hbd9lwcPEpUkqh2pdV9FNgyf/gW5mPIgHJ3wI
UA8qykiNaQEmBX/47FChdN/cjdpOuEiYZilLJUQ+G/vhBDXc23K4nEN/h70zZDBIuBhT8iXpGus4
ePa03don30sxLUBkc7KHxEK4woXWDj822a+jzYpWoUQd0cvzZjZtdYYHWX3W1cS8+PS/47SvFwpF
lCgLqn3qxMXwN2GSKaz+hPvPA0dG+31rC04jihMI1MxtHnUx+kjTbneVK4yfVmk9lmcN19p/q3AB
6i8pbYkeWTdzropuSUoL8xqcsJ2oG1RCj1tP+JUkKs2zOFTaQvWv6jbyzI6sgdZCHaAM8utmvweS
q3aaaDANoIceBWRjI4HXw8RnL87KlEFybMdHSvvzEAePDKyTgaQjVt4YhbId6egJ73pEUsbQyter
4r0QE5g42xDXj8D/8dXaQ5zAz7RB0VrRFz8Omyniz7CBCFu1wpO0JrKAMHFpgoAU4HJdoTjrcAOC
LHt8MUXARFnQf6rAMkn68k1e5MGWPqX+oMLTObk5u1SOuAje5IfMPVCEpW1yCrvIqD+z6jWq/sF7
uKYpZQ3TfV2dpF+h5XAmJW005aLpKet+q46jol4vi/V9oIkWhTFOTnw4ivh7HiqqNPYaHTc9m/5B
9UPCuHoFXU8aKxVUVMlhiLtU918CbM4XmLCAWPowAtOV/P9aeAH85wKfSCSQ1wVfTF6w88Lja6+a
DiQijsTWLrjUr2tcNxm/jmkNlQYpM/hFSEgDQe/76Ny967xKa2jLRpV+ECxaq88JYqeA+LZNsjlx
G7rTX/mAufxi1SsRq7JINLbxFrP0Kxt1dn/JiMC6KLyXo5SZSA4Tjlh3qHIZ/FIxcwLOpHFnZvAf
y/7IS2A4t/30LWAXp9KJ8jld45PKb9GG9mAvAk9B+PV3wl8IcEMWAoR9enIIzxykGF3/LOgGo6BF
50cR/bx95vSrMrdhDV4igaQmn/oSxsDa9N+dzsE1tk6Y1rFQyt70nZnpFu/s3Xay3Y0RcWIaL/VE
1a8l0eD7NFZCcJl2C4iS5zvHnT7Ip6rHQ9tMlMY/OgFbYERiGz2PEXfg8kK1qUlRBD/yo8DDamfW
dAGDgnecs8B+QTXZzvIiWPZU49aF9cPBmqDh23+xszWfyHUCtpCRFzDEpnyWQgjg32GCgHzkHnL8
JI/trtKWETL8oHKw6A4BU4O9wXmylsN/r9JITAV59ssG1UpfQ/lK4f74UnDrffwDR2PFZ8B2WNNj
cTH7zERiC3XeIuofiYkKt04lPI7E3xn7J1zl/urHI4LG9oNI0nQntwGllIznXCvrk0Gk9j0GtBNc
X/HlKYNmkOCOwPIq3o2m1TVmlhmI9flf70c5UGp5NQ+ypfBgGFVVuPZBgRZ1d9gHHpH89mL7FUjf
6rUq9g1FQYwsNEBOzVVa38sC2sLMppZSLFrgoR6ercQrU93Zuuo3pS2DMus7nfKNRZYdyL+dXADW
xzgnxXOKvbvJKHNC4s0i/Za+Khvj4S5RJdkMKt1PO4eF9dRoammGsnutkS92YaG7w5nIPlYLHn1X
mC+URoS58L3/1L5XbgqnlObOIiheuvqQsZ9BCgB6pHUu9/5GMyzIN0Xshn2hMZsjKr4Jh12Xu7wV
K7oVuZ5QbZetGMx+4vH+GcdYDT4YkB+A/4QsaIbhcAoPaiV3hLD/vz7r6LoXUMScwTenAQjLelXJ
EZ/n2+JjHyUk8Xq4TqUvFYzlFByp0BqT5XLB3l849qOwfEWEUjNIhwvwsnFo9pO0Pg+znyFkQDdG
CR6rPaxSairKHZxpgV5mimQiyY0lEZ6EPsWjdE66c1S6gv1S0OrUnpIrPYUaigMRhwWibmZk+zb8
NnMcEFWDLtsI2qlL5t4nZQOIRvWdIA1Ew0w0nvtnRrMGn6V1IT0iAKF1irqaArC03V2HHuLo42QJ
Lxlw5rsKhNYFacMw241FdtuviG9UEVIc/6NgjGovJrAz2+9oC8Wg2y8pBfhYphXsNhmHEA5WE6CR
+6y3Zx91kSuTq66FB2iDu01Q/wb9lAcT1E/Ja61gUOYryCNtRZbNDLUiMxSP99SkKUBJPm25krso
Ns2fW5waGTWrHu7Zbs4tkjqJtifTZtC/3oRbmKuCmRyf8ryx4Rf4amvATv7WVgnphbBeIphSdM6Z
yL2ngEgRMCrZIVs6mIi6kW89xcbUfrFxbR5pjrdffhs45VZfjT1hVVr5PQw3F2Dv7jXFOrd5ruUB
mUMtLTA5rg4098Zu40dSYSOxeQLdMG6JhQwoHuYSDnNYrt2Z9mc22TY7kGgUGdiW92n3/4yVKX4b
TPOmouGUBsk8E0lzIJtMvgZSXGY/K6nK3SM7av0dAVahg2zp7fMaQ6sw6zc6Fk21lOEnBHgrwZHJ
fJoJuTg5D4uop7NQFxHL9M8/7pC2OyITzwJKR44OYaRjEEj7PLv9RARhuUufE3q4LUMhI8QPAGA1
+LTc2MTTQYu3zv74kAJEyaMg8SZcgz/GtYdgLGFFwuyPx6635RW35d5KaohboT5SVAJj/oh/vW+o
LItmbr+XcIzjrU8qd+85s626xXFrmwfrW3dfzCMjFr0YnyU/Q/PIp91Nc1n69CVYiOr8EFM93tky
i3WJX20fl0Uc4DdTZtx7uQAniLVpudV6OGqdS4/ztLumf7pAOV6vK6HVHG6KChfSjiXgnJ2hbGmO
Ui+7qTC1qlZ3UyonDYMuy6GUEX3zYPPl0YdFx7jhmRu6m5btf5l4c4xmncxYJV+MBT39AmYoLu7G
5r18BSvlID9cSXareiT09SUqyIlwFTjbiZgxF2fSRizjAYlo6oVG+cyR5F0TCQs0od2f0eGBVUCx
swX7QFoaYfXWAI5kQPlkUg0Kw0a6QyZmeGlGGLvJolh/j5qJQOg23lqIO9m16VwOmz7h0gXTQZ17
3NS2FOk4glaGouj3O+pgIkm8boszVoT9QPDXR0kSwVS+fLvKkJnU//FFksWoJ+8n19ARSIYeVGtl
kUNrQ24Nq/W3EFZ2BISdiYTsMfapTtNIFHnDFiDnhX8zcj9lr6nX9eo9XMnzaeL7EeqwaFL0kl8H
lOnicm3WZ8dN1UdYJfMMRCC+3ePpd3tnBrzLV1v0olMn3WtLAKzDlpkN0gF7z/7zJI38bbDMLt74
JMdbby6fVcqgydK4fh4ttAcUOFWF68+ArzQG/yWhXjGVvyR6qFEK1MECahy3vZmWUUOmjmn3deot
MC58Z5+/2wnafJnyIkb8AWs7CN1+XyYjXIEyfLi1ik6pg8iqoLuIJ/wMPjd2BYAMHnvweoEcoeyj
WG+P+F3n7Fnt6zvQ+sPsBVzv1HquNv2oLLFo66tf5G5YsWE1QgM8Jmt+lpTPlnMFgu0BMTo59Lh5
QQJhOhv3FO1V3WsOtdM1K8Ux5WabAkmq1vQNgX86yH3Hvfbu6AEWr8SmdvKh1kzDK55bQC0v+Ggi
wJy7NPLQnoOGnta7zHIYg9B46oMgNdfhwm6sdnib1OY0KDxg9wifBexPbFx6OulGiYXoBoIITu6w
K4OopSf+o9kP0ws/5ey7YH9+R0000IRgYifoXxOA3KkpDy8yIOJBCgXaiinZTkkN/RmE8uOmlGY0
C+Wr1gLjyDD9XCQe/62bDACBhiZa0+9Ak7i7hhU40Y1Qog69UCC5Ut9lN5xb+gR96mAJ9uxe3Tc0
L0qxyh106SusLBNM+8o3ZsWdDq/qHmRleCT19PuvbOe/ejl/eZmSnbK+mVuYSbx/ITChaZSXsif0
eD3zubQBcAtZrPAyDEYsTck+9c+XdojMHkSOkpQ7BmH88qb8LU/D9FMrlzjlN9P7RMYLe0ICdvMF
wzjBrWXMlJeZZms+gW8ZjZ3VhMnALcmac9A7LJSrwr/CCDO813Qtp0bcMhAgHOX7+R6CLqdHNd2y
aaeL5hN/Kv/OZYIesEpw0JSoocp5I+dAZRqMah9QSqL7g9fC9qquRXp6Q0E3TJnjbQZjY2EuZps9
DrpHcmoK90qxuVzKbz922ZDNCXLBo3am++bv96SWWGVpC7NJSG0LLmrUGZ74KK0LONM6kqHS5MUX
3zPXkps3Lcs0dpHRL+bUD5ny93lDMqDZSy7P08VLxR1y2yBQwkxzJyS5bA4AJwPrqPNnzmMQhX+O
8jgIA8HRHfCSOUJK+rEWkCzgl1AVxLm5A8GKhFGOwcOTRVkW2eHBhPb22vpHrolKeK1/jOj9DmFs
jt79UJldtSS3FNML4LkyYyvedX193jbnc69juEVzwac6iUGs7G4x/HUX1z8DLJTFvhuU5wAqaZi2
BknEi+JEJYuLvsMy889OmQ06gLDEoJe0K5V1XhdPP3bwPqyfyMBuZcjV++PWfYGwMgakdXkHEMuK
WWBkefEwbOvFMj9nDdNVJVjzfBwBG+1YarKABtX+FEENf9LpRm0q1ICOE4IuoSX6+4MvI1vlbdJK
bchpgh01oJc2I/8o+W37XCMBZSGTKmtWxoWXgLvU5fwoNDfjgtqYbtBtflp6MF1p90UoQb9EzaB6
NV6OeAC3txvY5tMykFJvZsxCc7RA2Pvy7wYNREkI3N1t1JX6yVDjMOf/e/+Zx7edXeu0bVB+HO0w
SX5BbiAAJTlihHvBGOBZK+zLBgj22Z12Hd0SMNoqJOlDN/7N/rHwUBAJEzwr7qv0JvbT/cRmjylu
UrPyc9rP9sL3/8da7kdpYX7wQWuuSVeAhu+Dxyy5C4Smmq8/NVR/Y51Am42oDhp7EPKJCnmRzdQW
rVos05Lj1du3m8P8Hb3fX0qwiiYF7gxDWpjQcxXL2Solsl2E/Bb0CYiXlQaHepi/Sim4w/0Ea/Ny
4DuqbsHvmJCn25ScFRmNo3naxzxJeGP0/+j1S5tTx2DWMtpJYcn9te7cRvfnqgCIByrlhE2BVGh9
YuZARWk5MbIFKCp1ASFdIOa9csfjYdmD8HQlERRNw7A1kEEiPEZPBV1porZl4RoN9K4cZDk6Y2GL
4bjudBzFh1drfEhrxHGJ0j/e/UPD0kGuQbIRIye1o9cQdNOjblt8Ij2zr7qrUhAteLsTyLECIKZ4
VPE7mkqk+9/vClftsXXL8AlAZf/vcu+W5mo9TBcjp5qsGYG0rIxGou5xTqqouo8at80yGu5tpP3z
4vLdARCppFlJznS+ZZ9XSyY2sqcinkPXwqGgBRRrT4P7KAPVgP6oQfkey0EyLJGsuhgtmMhXgxhC
f+z8kdgHQk+eMJZCIj5sUqtELQ5l1flwTHQMB9LZORFQ2a4y8VcwLlPx0AMwt4V9s3LT55fMEu+j
uZksqzA0zk3Yv3K9f0Kg/J6ckBq6Ru+qqNotfFsZb1k8GhtIhrM8khhPqQuBdiGPZnqU01C+rEDl
zUOEYBZDwovLi6KUMPvNXiHg/vjwhC0NoVeLxRejOxtXemhpDUuURG40GhX+Tm7qF6GGVQYXyczM
TePZuO/uex0mHUJkBX+U20pRANtl4M+LgZyL8NqIVv1TK/MiD53zKqWhO5ZDX2t1MSycwn989VSw
ZIzKUw+7Biqg51Y4hdbesryUZ2X1eqq2uvR9wOanRztt3dMRa4WXtlRgK5SWhiKOO3i79c+UP0Yb
lUniYopVRpvGHpMS2fBvtVnU8lyzIcZWppqVROFjeZZVG+nORWQbNoUfE56tiVrt3mqV5l67JMSI
mfnCjQIAZUri+IP1DkhGii/ERsJio4SDIyuaoQxZgJUUEuNeh2GKhEcw384U60cDjolI6Bv4tLT6
Dg5NsV7DV7BO4EJkEPbm5eLKenygwTanAEmd9uk2hnUo9GtnwoGBiL15TdiBaIpBiJ2i9illRmH0
1uaukiLH+nkKqKp4ZW8udquVi0vzWy3BmWWeMt7MxfsHwqJ5Bbh+HcwR2vFr4XjU4GLX5kHR+0P8
B69cCRtC9ZK9ioY7FWz4jyBrnwaSLf7AUL14Xcyyvi5nxE7qntGYg6kNljpy9lee2WcOaEcK2ctk
mP+Ll7sPLUcM4zMSNmmU5uacHPZJe+7CkLHMfHxTbPlmPIINOYBi42uv//1GCmsc3LG1HhB4NWHl
0h7BleK9uY9wOPTUCp3jALdjnqVqus+LVPz04fP9ORqcEnTMTVlZBSVkIXyhTJrE/8W/sI8d6nX8
kaf/OfH+y6sHMgvMMX4dSx1Nw41EkWAFqO/X987ZUkqfRb5WtJqp5jeSxnObkPnjZWLj7GUyGIQ+
o5R8JZ+G8oQrU9bd1u8dpIEsv7JHMKUv9VtjnO0Z8RJf3DK1cVBjFw00wNQA7ZRnI236ZVmxLWsz
vrWItWWh0NzL1KV0jPP8rba9fgxPdiFAqH0sUXweb/EgFzZ2oZ5NiuIXEuC6OzMfROnK7fqgrFmZ
9HXQJeN8D5RfgwN8U8u+hlMvZo13chrYkKW1hBpWLVLfnOxxboih0gnJRntRUknQGZnYgprmXaBo
IvdR0QVmUtR/xkxVxhtsDuNMnGHI7lVoL8eMTCYboEDmOzvaOF096RLubDLBgLlig7PTcTmvaqT6
2A9jPw9D1zZhgcdhodSlKcCQiVolvnHh0PkYP3aZfY+Vn6SgLlAnP3ca9O2wSSi6PPd1tlOgAOsc
4J0nvxNld8T2CQ+MHZLl5tMDGQlsLzQ+4en1AN21k26k7332gmPjMGl9QA/bQk4/NOKmiDU2MFrS
hMK14NcrV7jrIvwyAkKi/yFUfx3rgmN/oUTCiVWvwUQ8IbH3rxKnPJ0R6Pwf5CSVW8VxWt1Tevd1
z1xlzzMpkCdKpPRPW93nOLq68NwSh0jaS/uD0p0xvGiSjEtUqNWKYfv3oJ3OFD94zJcNZFoZ8Jrm
1uZuhDsYP7c49sIYYJl3WGXLJr5qMfWNCd+q7OO9BjJEfDIF3GSLkH3E3JRfA10CHQYvb4ol920W
OzXgQEjOSgnOQJqF7AHFmduQt3qxLjXQqUV1G5zGO7ZZ9EBhnRe9LyaP2EsCKR82m1lPB6Nk+Iyo
ec8Ri9N8Lv7hDeJbwYWWGhUuISKwuw8uxJiH+swdWkktHlQWTTmffxvID3sJ0llfPVrC4I/pl3vr
5lZatcej2EqQK5dH7qXKQZYl3yMAP9Q4o1Ux8YpAg6IPqvUwZTFARwYL4mb68GGqgnT5eaLU5+Xk
i/neVXkp2gKAVQQmekzM0pWjsm3SVJS8VHIoir59GL+Di4hvunVow7nFzGBbzK9QG3Q+sXJiZJPr
yT0/AxjBdqB7Vekzfb/IB9/MzwOIGbHzPlRZNTRgay47TfX687D86NMqB7rYCq+Ft8m24RacFMKo
6QbDDqv5aLueShI6hdVnisLhYmgLbkogPdOD/NbPgl7TR2X3ZOEfqClHDxMWI/WeDULS12Dp6lxn
uiO+TTr2WxSRQwpbjzpcHzLZ2pPecYAemt2ce7/yJZIR5tuUHNuc4R6tr53zf0+AIJIO328NU0w1
2hEkkImoPOUDqmJXNQpBvol6p860ycBWVTtxhimk2285YLqNUy4FPso6rBYaO7UhofbCx8NWo1e4
8K/8aU+DM/lTfwcNPuZf/nwr2R8TrD81uCKM2OkUMmf96n9uOxtp2mfUJ+vU3TQG4NbwQrgsY2ZK
j44Em6elMrq8N3alCwNMNh1xlZdlrYkP9akISn3FWUkDZP/edJrCwSZ6/II4xADT7WFvrFR9CcRN
M63MoGqfZ+cfEYrOlY+KjhkRUcKc5QP4M9ztP9dgqAnK64kk02bUizElhMo4aP2/Qvf23a3eVKKX
3NFtC0u5s7kzC+JnLBEYovcNZ/ro4S0fiWX7/sHPJ+vXTQfbI1oTGgr0a/LMn4pdIGcVRb/vRwa0
sHbHX6AnVGKa0fwIWuYBrMOJ/DM/0w8LlviK4sH3wMM6oKQSxbZIURPkUrUli49mCxSJ8k/RDDTN
EZSdTDe76erBVYjpY32gobWs3bwP/3219ImJx3moZa8pfnuFGLN3p91ixEFW2rmNOZ22voR7Vr99
1HB0f0X1SjE3FXyepzSESaEHoSh4oyBsRR8TTagD9sE+6pRnuqMs6cnkl+tQDwQxDxPMPlYw+9fK
Cze8G/9r9kUcqLwmYw7En8AHtow4t8k2bEp+86C8BbBUjMXyViwyy9yslk5R+EzKQ5V8RSFKH9Zk
w35nVj/Ogq+UmrqeHTieLWcwlPRzttf/TaW6X6eAmXBAnRPQDqCtTmv566iQEcNnQtIlMiKAXXfS
y+Veqd/e+xm2iMrr6JjVfLUeXVqAPWpXMdy6mYTDzsevtavbCavC1xtn58tBq1kJKbuO+UyNYBwZ
znpFCZfRcottmcuIa5ZDc5YN8nbylVAwRJkjdI5tSmJleupsecxCAI7EDmitZAEguOx3hDK+vhrP
ZkoZIFpwBNcC+mkc0r8ATKhI2c/2ae30ivnlixsNuWpNwWqXdwYgf4A1PV9fPMnReoDnmq+sKwGL
0WkP/HHIopiy+775WfQZUFWEo4FaUOHS9rc+Go+p/ylTDGlbOatEdrQU9+ic+Oo1Cp8aGi3xDuLv
+JGRQrivGHzpNyp6CcZX8/f286umVmwLICzSvRYkxCHKWuQA+aaD5/t4Q5hR6u3FSQWmNi2/rCc+
06omiSuF3JpGO8BVjqikGFufYjzTB4GJubgdhjK8yb0CXVvd/upFqdYVZBLw9rIdR03kvZ8ibFCp
/ikysIjXyeZZ2vtn2hoceGKCtAaWS2lphwW79+WPR3YMitzfjOY9HGRLxI4U7ThR9/dc5E+Vv95F
5hFMGT05marnaZlGcpt5IQPL/NTLJZaulKJcvFGWDUUIQ0HddM94p6TIGMszJf3578JeLQ/gDBkC
fBw2nUB5SIt0RQfy+KAlswTtE7LFD/+Q/1td6fx42FrVzqGaSzV2RO+SKZq7ASZHyIkREgMQWXhA
THBApf5tTJ90LBC6wnKu+wDF2VB77PB7NwUzP5Iq6tYgTbImqsSw0DBE5BemIfFvGaNdV386fU/X
VKrRqYHPoD2cJTXSG/0o/R+j8wNs5D4q9x66xUyltsGhj5uWZ/Sc+yjzXthGBwPIvbrfuw08auyr
fUrpaQvLaVTuw6MvClRP13EZ+L+uzF8gz0CBMej+5v9+acdtiskf0wz0TnulfDaAV8Hzc+8rydCG
f0GT2pnLZC3DrqnUB/9a/GQ7LVfHhRUBpnAkJRtNRxhO3QyDYd1ISFqWY8DAEiZqjEzqkSlpUAOb
LnuKBak8yGW2JQ0+fc04WopsqYIxFQPhn8ft232Isz1xqM+H5/XyAMoCD1BHyVqEHSR2szKp99JD
p6BixmfkhPavDy+PAEr5L0kEHkNaAhQBXFaJZGS1lPa0wKpMH+ngihfXW2CbzVITnjf/bFPAQRa9
dWRcv9Gu05jKhlYhHNrM5dLgfg3yUfYVIDT/tfwfv2WpsnRY9CFDa22WNcS0wPBKNAvrOtLoE3R+
ar42erWzMWDmGH9wAH0sU7Z+iVblyI9g9BXA1HjP96e1Kzk2lsR+GQTsjoOoAdulQtXyPsoWmuLF
V5g0ID8Mmi/XYmQhCltQRfMVGzJDTgStEFzRQrjAKRsis9MChHp59pZS09d2OBjhsDDdhkK8PIZp
bbjA1upZpuJ+d+6m7LrSCHH/P0YS5wNNp2M4nfwKLoiT6whOEgScgcEQRIH5xnglTM5RODMKXxYB
XCjNsXSuygexr6/8iRWL44Bx5B60PLVauNuiGNV4b6HUxtOxpVXw0Ld7OioM1EQpscfAAIVZ38VF
3Fmu8AF0tRR5Us3Cx38P1txaNr9mdb9WQvC5T3EozVcE88xNN7bJR2AL4wdjPASbYEG2Y+YLCj4O
m6jMMM7nj+XbVXubY6u/AZDL4uwzMYxbcjVataUnk9/uyvZHIA4VWOg/ZliXlF/a5xzJlZHqC8ws
73I2A/DbC+T+w2VeRdU8nOnzFmvbK/XiTEnEEs2RFvC4MDlfD8HK7maXwdgZixMlJrL2nrxVTiYu
y8KNwdRsHGg6pvGVUXkwGi3XTaE0xCTIywXol+xzX1tfBGKNQ+EOaN0vFUFrR16SGjA/fYcWzZ5V
3cXmgeqiWUzYFemlAOyfqVYQsRujd8kEl85VN7yaKG17gLJPB8frALtTxjLlkufTFVe/ULv3QreP
Ba1/bUc5hNcD3j4hFdUgqZ5ramu/4dQvDt20DvDaWfFvRAOCrXO3O/bFx/ZXnvhBsvJ9YkpU0qUL
8OJpAPnWPefAacRZOTH6UI/nyqPuj3xkUFsuOWVH/ZQlT3TRJHgehNFoXYCnYPHOIKJpglY0Koe4
AmbOlcg0jIrLLQRzTOpJd3OrbsBCGycfCSWSbdwZmB84QesIH1ObAMkPPAYQhgY7AN5aXc1ayUdX
Y73GxqYH8zteHXOeP+CK0e4p2upZXGwGO2phbmvsTpdfXJI4WbKB3BvnzAGoDnVPLMnGiTPETk63
rav3c6cksuKNlJCyK+XKZjBIw2NnH7StzXrrop1qnwYGUNImZeoL5JzrLkV4vzHHhj6S4ysAg1wt
auS0790OvbWXhSzEpQVbcQ8oyiJ239GOhXmMFn0+oEtQQXSvGujec5kpsQKR5cbjwr7P2Szv5zJ9
YVxlOsTAZH2KHm220YBBx+PFn3ZFaJUGmv+zHBpZEipfnCPKf9lDAd+wvU4dtiF7S4ssnouHmCGp
WKLa+MGDIFi0P77mNJM3pUj8sBTeseDpAKd9MvhQhZwEV0hbB0yd8/zOYhUzEBrMG81r4RDZvCXl
ls/1RN0g7JiUD2xWN+HKvPNzNqi27s94ub6jxILvzu3VCFADTbCt5L6j59pDJIAQGkgdodJmWO4X
Gu+/ry1fVu3FAkYnWOAYhkHuD8ek1JaZMZeVUXj2hvBKTuB/ICxDXvGmMCu4Rc7W8Z/EZCyK20eK
BDqqo20wNbdGbFffav3IB80TYNBm9jfuD1uFkdqrbVztndgFtgi7vO0NL0lfvFDKjMNwutT/MydS
JbVbknh1hEjacB5r8GVkp+DFl5lPnjmvdfp7aP9sm7scFaz5pRSAU6EAM51/mMr/DWfiPHsIOm0p
m1L/V/mZB4SxveD/wDUr7Hf8hvVoY58rtkT0g1MeDjECYGWou2+JqeneyBEUG8UwJvz8lZVR8MTR
qDZ6pMMH63u3BAePWhvcPa6fB1ia2PYTnIl943b1BsnZSVD01youR8M7pc04BXDGpjyFaWpAxGCu
yYErro9hiJbUcI4YGwa472zApF22OCbEO/wA08VT4PFpGjhzRtkXI5q+7edxPqFOAgkzoyyXbgtV
DHXgH2JizaNLizodbzgfXKkLKurd/FLY+vy6C0XI6oq+mL1RiIcv5sfQB40/TUBB/Zkf60pLzN9E
gc828eVCQomaFzu5Pm2DQEuKlTot8yei602YoRfzX6OcLzIqSwO4vaYg/tcHKY3XxC+1TjHIDfky
iUOFsV7fBQrc/0OHE1vkqGX1j4ZeNC/nAB7LQ+rT9KNFsiV70NKGQBmi6Vu8boxQ0H2zubNo0vJ+
pMR0xMok3Lt0zFalu8mJnTtYmSPMgG4DoWdZjhiSrOJQttRcMYZu6WccMumAtuysLGSOS0BYIUAU
KimjPepxqgM4zed/J8IZft3BB4uBZNazMOqj66ZWDP+gajJR5i+JQxa5wqBXBlw5UKla1FbJOMlK
D15Zy+aO39vLuTyuM8/aHQOom9UB7TdMwGQT8HhM9a/PTYDc+ae/pm3LrJ9Ws6NMp3c1Hl3VKj1A
SjuECMtwWUv4Nkv9zalpoqbXGhpcQcbzbaENJaFctDEq1A0OVEoN9LhShNl2FE0QldqJ3LobZELW
S5BqQdBi7+RbFZmQfYu6NzCL5L6dVn7zn/+45gcLrtjXKS2KQ8bGSNhdNEKW0udl+hHr+8BrbAJ2
Rc5UBa+r6bQ06bnRyDZCXFRl7F3UqmmcCPMbnjfpjj2LXxTPUuQXZWxolkOUE780AVYC4avnSn7i
nk/VGgWlNdAe9lQLXQr3QoibwlalnDlM9L2z/rVh6/et6eTzyAbYUFMioQkgtz2jL/i2cvpABbdj
nifEltYjFTBp949KNMOTH9OojA6eQeksP4BeQP0k4CmCMtVYdOqwzd7cigY9c8hOLvoNVW0o83tr
v1gvnSz+LDT1s8OQDk/HCyyDE+WQqgfEiMo4IpLYZ0fJTyIJ9+FDNFMo8Yy0PVpdN05jVYboAaYN
7JczVQS6NGghMY//OTbrC26fizZmfWs6gE4VAIDiSArcCHuGqc8ECYs9Yi0xFVXSHHmxqT229WcS
dcDwp1xebQ7ZxTO7xoYmefrn2gFEv4FSnl5wNw842gNIXloTMr0dQqZfa8vpUmbSOCjchmE1LVNL
YgGXPYLaUCZ7a+ynzrJQsMUvpCBt9RkAfinR4fQjCGftad6AndRfNA3n8fhMR9O3kPGfSmyR1DFM
67UrzqBDcNcfshJtcYxXOyuaTtW7X2FrKM74T3saYUGSc3+0qp0BE87zJ12iHnslCcYizb+DQP1E
Saqht9NGP0FIk7oXnt26uazJsw9uLtCYuoybDsrM5Lvad6eLOakIZDMPqL7IP+R4D38q3LxexWEb
rikQqxLaUQObWsz7tsEWImlQfaLRMPvXuemMOTIFZPPZlpb26Z+n9BVRdrSRfGgP63i72fniOrrn
oHelD8sf5Iex91e2RmFozWVB5cif6h0G/tRx/ul62HEGS9GQ8h/E+DxEotd1f+1qAodrNGAsyaYN
wgYUUUlhvVbZ7c5r1PZJ0qhIyi74wux76OeBCViFbqq2XNiv7LZVmP4bVLWLbd0jYOGjGV34mDjY
QYpcdd84Wpf+gpKjZXIQMOgRMrtRe7FK3EAZ3oLAqK4vSbhaGsTm26WPMHGzSiNXm3LkFRsy15t/
33d+bBo79rrjoBdDWCmbOllvRLMX4jW0ixKAS9ZSA4Br32GnvDPxQT10paGbQ6dS2FpSoueb2dFp
TA2fwzkMokvyK9WRmF+Wu9Hg/3ZCRSSHQ5JQ738tSRNTeSfF2zEI01ZfkEK5rcw3Ic/oFap37Z2v
zLb+b/4P8WtKvrUETr6h3Xb4uh0cZPpsfW+A5eiH52ZNsAQzBVn5BNHVnyBxzlAltk0k4fN/hegS
N6AIK/e0/PN2GtM3blc9B+N61CnbTLzTbSOGE/2cZWRtDQ2tLKWnAtlQN+bzEcKtODuQTAKJtJl2
N8rPW1UejBAuwW/Vwj8p9mt/gR+0W/XCkMmLbpeZMXLTq9OrltxG6jzcqqLQGgFUJFqS+yjjyXyJ
dXOOesOTWiD6+Z03Cj20jyO7dFqqSA0X/olk/M4mMXWvrkvVxAkihJnznZY81MlJ0vL7ux7HSo4U
370p3GtRvvQEfhkcfWyNAIihVYPMFVxB0ThAIhEPmkBNW4axAviqcbMT9JLunoGFwgoJdbguk07X
+8xrbbTh4nNJAGEymXcLESZdTIItBcsUFt4PjEgFaQDYCBBFIyo7O2//L7shMU2gJl8fz8FjSELF
ObctTsjn/7+ZMRcVJb/O98bukFUDV8tX5wyYHfJBTHXk8XIJnqDCZbIvzxJXUEwBC8XpwqC0h2A8
/a2oldUYyqieifn7LbMq4XJcQefWr3N62sqVfV3UDmIo/5O2ZBYdKwBQTEFKsShoORe8J10bxY8c
TL2nojPmqmQDssX3srcysrgxJXkPY94BKyfu6ATHnU97jW2ft8O0INP2wGqpAwAMiGnw9sNuklJJ
ODTWbEjy8Dun5BZlzsfd48NyMcVRJE0k7v/GVcn4TsXlhBpB53qFDxWsxPHc90fn+aS1uIEuEpiJ
kj11GXrflcgr6hxwkh9SZ7DnlsbgHaLZ68U1yWCU8PXch3o2e2OU62Z0igt8H8JvWwjjB9Be4v8j
N2y5hQEuAKHxrUmgmy90GstEFqlLys0hJyJ9FwvQ9ZgNQDnig46AIl6jsp5eYfyLiyrKHhHA1c+k
Osaj0yy/xxli23PIiSvQB7CCVmznif9tmT6K5pUSHk49tXd6xHoG3NO+oN/uvfGwy3F8LW1OxH8O
KYpgZoifdUt7IrOZKL/pMuaWi7D34Qiq3tyuXRLUAmM/DcQ1iz69wSpvsJuaQBat3I8+VRVSkNag
pThprU4I9KpNNio88TcJ1sokAYtimiMaZaZsIZTVFqKSelMfl9m7NAoZNkgyJsEhTRx7X9gfXqqv
MtHrc/IIhOUKI2e89tsR1CLG7fxXUkve58XcxbajYEPn8MmHyj9V8MjnYxyxjmd1eJvdac04Muj1
65KqiSovM5s7oCgrm3k8weVCAzL6mTHCL5HqQq+GP28oqWqTQB8TxkWkThKUM3jCrzV6gXzBp4l6
r+um0uvlbBCYOS+6/xCzqH7pTYojABURPre4gtfp7FgVbPt7BDlgZWM1Tw9PF7p+XQNblK2Hc3HA
6jXLmFK11cAWyvTnMXu3M+bjSVDQd+htADZ/5b2Gku49RQg+P3e6OKgzhL+6rRSo46PV49Z9Qo3H
W89RIxQNnpn8ekkst2cLxASQiQtEZGlrt62748A6sbkhUA6UylEZ4hxAMBRMRJ48N7W/1JCibhBJ
ajVX4Tcy+sEtZX5WJ6i9eCtTYx4bA0h3gfa6qpue17FSCX5z+WTXcPL7Bmxb+5R0eeeX0KkRkjXQ
eTMnoWMCJwVLC4EYBLp4vRuyrpcAn9JraF8mnSpD3CWjI7CbEP5epX4caIh28mmg5dCnO7C1B4ix
Gou5MRAE/Z0S2J8dGEV+m+HPG+FKAsPRYvYrYmf29LNbbEARHHxB2IEtMbO4KUTg7gAF84rGJewj
a8QrjOm96AOPCqEQ9ujza7Cja/fktXh496hEG6J/Jy+UwqbSVyWYQNdNvV//ncdvlfdR+RvqUmck
v9wZPvWxu7F4WDLBg8sYYY+cH93Nl7DiHpyqTBBElkd92FLffLPwNnBpQn72AFLDyptNb0ee8Yu3
zsbFyqnogSnyTgcOFgYty9coz1lCg6YzWbbK80yNPk5f/ZQ0T+HKRnwt6IMnireOpPnkdfXZSMFV
WdOaZsF9Z+rPrYys1NjT+nt84vK2TBFAKKKeEQEOjM9RcaVv3SCa5j9n5TSfPLmtROOt0hEuqevz
SLOP5CQ1hC6zYTXKW5i95Begv/gE8VOhvy7wAGn6UGhzQ6MCZK2aT7aDlj86J+if/OSqtjfWGuGL
xwyNZN5ooWX7noJvMy4q+ZXomlLdQxnfPvbYOZ4IITPhr6UN57KaNqbqYfLHejH56LHHZjuFeNFP
ZZyvBJ0JAOdV6s5qNTbTVEWd4cp5leJ42T1z/bnIXCdymeaV5yB0z6YLeuhvstLghpZEfM0AR0FG
11pQLIXCGB+pe67K4PhPHY2AuDyW87WUfQp9ZjKEefGqw/f3rJDxWgotULo42WLNimVkmlNTkLdy
shHE1yjAaDHg6wZNob5HbhzcHYwJwkFU0aChzs3z89Cgz61D2coUyLe4CdUtK0RXT1OoYPO6tNy5
f2jx02yte8tV6LDnmkOmr/ENtQe8WAqxZbcv+p6oOPAOlABMkuFmbxS946M+cKSQVOUCSEISYV3e
feLgqADi/emm1NHTpZbLoK/ilLZJsrJbUqHQ5ePYVJMtfc+I0VBlewD7TyKwJ0a1EXG5RpeeaChC
orgbMgdnjJqmA9s2DfsgFI9pVPOsftNtackDH/O31SzQRkoCJWde6iFNXVTqI9PAXvT2V/H31Ceu
GB7uEeQbvclFDBfofrXjewqfgaSY8KpgnnbkRLHAc4jqE4Bg6ImjKpp5UQZPVjtQyP80W3ZSuVhi
tlEsAb5Sb2p/2W9C7UZF77A5jNNyWa84haSJws+c4R8X++6sbcZ+kZRhNkRXy2uZe9PRHEmGmf9Q
WiWxVzd0zZZxxmtpoK0XiEIzWoF/55R+6EYQB5f+pXgjndanCHOu4hlPv35GnvxBK/pj+L+Fjx/n
xaBD30aHrwtbuoRsISTwAyvDAS+JcbZVSvIWfUQaZP3JcTLKwv0cYxvDUmr9RPmxa6MhHebIhpb8
4CaBseiARyY7XNRDj3kAYrezeoLidcocFAomgE7hAQdisLgNrQEuzhehE0ZaYqlSqDKV/Gl/jeqd
egTVC8BxHY2V4D79f+li7Uc24Zm8yzr19POuIP3SNRYmTSHocwUu4rNSq+aMZzdN0b0+ne6GpMp6
Ah3Ovkm3YDDKgS++utlJ6OnfENHZFYsTIiRyDPeuqSXbrEfsL/9kOA4rm7n8i8mFdmDOpp3h2561
FrtOkSCK7ZAAcAMka/FRGMe8JhgwcpB8lTLVOUM6MUoqzPQUsxmi/lxuXE8fszddRrS8kVwg2saM
3BcoUlLj2xmLrCXeXGtClGJrOu43j0vZeLLIA3IrxVgmmuToR7QVZrpHNeJdevA6UMS3quNyfRQj
NOurYVyZWbGAsDEfigXztMX5Ghlyj2ppjWcgZCFQErOaOdIYLldFEgnTDLvjkHYdVQ42sqc5QN3d
obZQeK1IpLroBzKZNkT+w/vPe9xPfi7vtOXJa9SyVPYurn0hJS5Y+DD15fTvFeZD9hcZPWfsjLwA
lQfp2fZvsNARcwZ5yjKthOgf7gnhd3yGxJNeXYNGRaWhpuOJMihXm/s+MwudqQo6olQjP7lpolCl
+nIVZXAkmcuaa/pmP1L22sxxfN9gi+X6y4WgBuEFaGN551e2ddWxGjbcEXLhpLH1tgp82AteUSNW
xq7R+ti6ZNp1Vy42MnlNEl/jOQTtSWZk6W9MR99MzIYKvidkWGVxaWBJFOI7kxi0xoDCs09KbFwc
U9QRRletmfFJF13sHDnMG/iiJGovmK/Aa4vID6qHD2PcnvYbqzQXdHiPmpK1v1g0IOOzjCnhV5At
vbcU+u+qeB4p7fwYy47f172660WG1k1FHDx1o5FV/9XMslFGZT/Zj0KhRtKEahdrW2DL8KZF81sz
aeCQxOt0VOBuO+hGKhF9RS7rQLvgP5WePyyUYo/HKAr8QxiJybhhUBpAXmCfHh3lQcx9uDw+Cp6M
DabKOQ9bm9AotY1AhHxtf64qxe+J3jVmZ6SSFGPb2Hnn2wtr73Nha+DGtCpiEygoe394DTP5TObM
uhNY3NxQEZUATTTfK9MR/kBKcp80eKmpmEvbaGB4eIRSLH5B11AzOFMuyljLvRn0+wTwZHvD4Bjr
5X41JrQJCqCTy/TTEB4bUy3Zpp6bS3DfS7K3ThNehE1ZP1zaUxK2Lkew6q/P/rYZ+8zEvc+OPxVY
X8xb1nreJ/1BpjRcBoR8mX32T/z96haVJmRDRvY5LApL8Nmw5fVHwDlaamaDfzW8bcB4u685q5Qs
CFy8XnjJC6/nRxErHVQfg+zJTu/KJTcEZfhb7Vm38JHmeRgobVF9vXG2UmzXWy6HVveC2H/wcoyD
AJ/iholpbklAOeVY0moE0pl6a/nNVSl7xJBJ+7Xe1z2oVlQrszjYh9j6aoz2S5a1jYOJ80d/dPg/
fpGIX4ggTitEfpZhmKY7nY+3F1Y6noq9yGv0Ik8vq2GSTRP0AZLnk5DALkAGq+mBSR9Q1adviSSI
5vwN+EOStzMAispha+QeNJMtrhfDFhmH8+lvUuTWVqGI7GRVhleUaeY2EROr8zG1giATFf36eO6/
O2XZ3wX+vGHXh225P0oceSZm7jIxKpNJuRQFMJEM5dW0SCK550p6ZZctpLMLeWyrzZ3dAsWPuYuL
evBWX6HVJbcyI/aWqeRDL+6HjQLJQONqXalLgolxhRvLhHp7b6YCf/ILPyd7tssRFcvhWILSkdrX
PIhgGbXgIaSITFGbRkRHVklwxYltuRgw4q+aLQvtWLcK0DHQ1JAr85KDwphIqUb0GFuRyBSmyP+K
F+D6/xKRFRw6LbbezbH47Mbml4zj17sUGXVYBmQxMjqTDzJRqCKhCMi1ycWXFys96JabqJ6Li/k4
83QCpDS0T2KNi9UN95mK/raAvUGRTuDkeraMSAPoYsIkZ1E3auppyrbYvbu05Efo6QeThBmt2qVI
9Mb2iEVNK/OKqoisXZ3fU7P6TuXmUT2HJ/GHsNItGcshMP8I46I80zpi0D17q4XiDTInjRQnF6bK
/8rQ3lPbd4GYheHbuYCMQct1LTtXPK/1xrbH+1TV59Kayrbu51stHcQ5Tibnn+/45ieOoET9vcxV
XdUUw+xWO4EcLV1wt88YfnpBQxm2MloRQdnZIZ+wnY/KglhWDfGkbopIh/alTL8+jGOKyDdojhAi
F7B92b7uRavTidfsYn8+QZHVMT4mCyTg9BJp64kXmi6mBDtHhgetgpW9eTVg/pvrAR9qK7P2kgyk
eLCvRPn8+fooEK9hMZlk8f8Ob+0KlElRWzjOIIjMeX0gdl2vAdXWCFOjEBi8gGfzA7Gp5/k+99eS
LvuwfzlxlXbFPtu7xxXOaT/Ze7++cw0OFzDyXbNbxmfU4i+Fjm4obR17lX6qFhuSm+nmHifrh0df
/g3QzOUHw3/UGfGC7PufY9+GEf4o4qYP6EECqoSGt0NWc8v4gAFfrxREBG0EMPhRwsFVFlD4Bnst
2ZbiinlY9RG/fJUdUR50DrRRwd8yHFH1+vDHHiEzycshkqT9YRyFFTHSG+YmU1Z+44e3wg/+Z0+q
4Bs2Xsu5dd3l9oWlV0wPId7dLW5wpzu0jOttZzMucDjyCDl3uhs/Y+Sm8HpDFTLpwYzDB+GDN7YQ
YRM8m5amFKkREtbBf7GdILkua7F7oDHu4Sd5He8BtCEpcSJTtSVOSRy3pY/s07RI4rTYwKeFcGtm
L/wnYmMjLaOwN23JeN5ZjLyOcFyLHzxv63UL8MtulFkOOQ+B/8T9TXeEQ6AWvERnsDKNf64oPKdd
dnjXHMBcn6WmfPLbXTErkTkT2DVqWxMcklQ3tFUUsZNr75QZvpnMPB6C8/p9moS5703sHrrW3ITZ
BUEnO5quWsqNCI/RBOyO+Jfp4h08zS3X7zef/28thq6t0alvtee6FeD/cJ4sIjlXiKjy2guzjcsj
n4J6m74CkJ5h3nx8VUIdNYhluV859SjGydYiwDhCg8SsWDX4wkFJUiFx0+GTs3kxby+Q3Gxs+53m
ugp2gSFTWboiW2zmb//HyXtJhkb39IGE0lfcuzwSWy71ScGpnY3AC8TrPEojT3PJxMprHO6fPL5x
V1FFE7qmC2XH62VEH7KuTt/CRfIm75t2sIbB3UHP8SDxB4p2/slwTQyNhGwZ485oFTV2D5yZw89i
d8byJzGz5r/aOBFBHFJ28HYMlFFftzvZqfrfGFlKBPq+wkO1fua9JxzKm0NR969mTx1W0RpJmF2t
exa1ZCH+ZbAFoLWwoqUwfj53I5RhK+kT83cmN89ESbsxupkpS4aMw+Hy97duzv1O5d6OE/V0BlDg
mO+LG0f00+iyyP2YFZhbh+I2KxreuYNjgzV4tlkYm0odR9vmC4mp1AJ/l5DjE2ZraDjnj2YPMt8l
cF9xClgiOLtBCnE5ru6jREhSl6J4pnvs/0J9CY5ccjLwvsZ5+Ig9hguqwc7yxZUS5xme+l90ssEs
VY7k24fFhuAyVFIK8thoLaopjqq+qoaqAQvKpeH94+7HkkOPtyCEUIUuDATbFNrZ6EuHFp0NLVgk
ruHbWQr+OVXCobjiUivrMwHAaSuB7GxqNqfa3m9lkbO0PM7PtY3heqMZaNJraEa98Ljil7NRxOOW
psqc1Bn0BjSwIJUQJyqDzlv9qTP6TXTKtKrLXc0fBAn8B5isupXqLbzTP54AnkzMMlacV2WXPPyX
bIKOkutI7i68isWelMaT6fSmsIrj/61fCyZXrCJtWHavXLX8FqXC2QcMisJ02SM8sqZ+1ajn0faC
ZMXt6olM7tdWx882pI1RvuJpSEKwBGHxskZCWaEwPfZtmEzvJ9S7AXU1IBeZfEvC+h3j8PSxwafK
2Bhldf/a3Efoktg3HndmwG7BhfXDmv4es0+yQaMq5dpZ3uUq0wgb6jD5QAv8e7GOhMx2AFXVDbQS
QldAQdIp7KU8UpPVOWQb96SeYrNsZmOP5Btoi4mkasGTwrb8bEtYCSClDAY6coHW5h4/oxpZnpO4
P6x1Y6msWmAJxvk39UJlXLFwTGmOKgWk5RStHMrc6Z6tZMwko6xTRIQEBGMU6KOYP7ol7KqVBA2k
f5zWbJtmxnsWtm8Pzoax06IGBa/vLSDNrk8yECB9lDf6ntxAqLePMhF355XKSxialhZcfHQ7+xAj
mSowXvl7kwvk1u+BM9/yjtI9hbJ7ef7JEe0LUHBrhxrnA/laE4T3P9g1+/rCL1wyeMbhZm6jrGBv
SY4pE4mtC/7YN4IANqsB9ml5Ik5IgA9BOjdgHDi1HS6l6Qt0mC/kjlm037op+1TgFWl9tpIEnQJ2
5RpTA6o0U2jsK7T1V5C0LYQ3thjxkCAzEYGtHPG3QCHo+KVrISfWv9g6As1eAviOAXT7U/iMQV7d
8Rsps7Ve/UVsnJTodbSAB4Ru+I1BobwuCg7sroHldW0jgMKfPkGGDJRwsH0D8fB/+H7h1cJZGCR0
MxQmopHGMS+fzgQULbJ77eVPxsOfkjM7EI4ip+yat1UVw6cJxpQzb9Odqhi9Uer4gzLktE9CXVZ2
G4/ybDETYlnBcrJfLyum6m1geacm5vmJXoKmzZZyln+q2QFDq06hO8fjCvcjeP+s1LXngAPPcXQv
aR9r/OAq0YAqScDieA/0BQvUro2qFJ26rgSFI+xBQjO9C8on9+xG+g3xvTrUucrs2H8zcPQ/NYy9
T61QWHRqwXg4gNMhPXOHITrbgh3ivxSidODjT05zCyl4dc/KKgjM1YsnuDVtPqgAIXyvd6JHb9r1
dw904ciM/8CdYsAONTWiXegxTDaZJ4vBtMa1E1IySO7tw7f2aqEJJTy+TAOmqbzM2D3wYA/MdQ83
ypDqeKtS+8IyQnaBA7eFJaK+OmmnutLpyM5akTS9PaQM1z9IV8iNm5oSOyxi8B5Q9FWBqECiOhX4
J1WLE6mxluZP6FxhnswnXfR8gS4EDKzlueNq4S9lo2p6H6HvvqFsUmiEqDGkM6oMdAJLdKErDrbf
4goel0NzW47psR3dzri6ZOFgeK3FlZBe0A4cFLiJr3174kdEEIhZcJ5ySc1/PszliplesWRqMS5c
7OsqCZM7rIOpxq1jz79rGTWZAsUunWDR8SNGZJ/JS0lrBpXVuettOoOioNRYhhv5AHvPsO9wVQV1
uM7Wc3A5nELWgAYjYcXFDSdq5n2Bv7aBZl2VerFtkIgxP7VxcQckXRjxbWu6YB6uKdO9OAamWYLk
fIYMxt4wDvELKa0hx06C6dTb2WveprLY9+OooDpv5otXqC4pmyk6zfEvrFRvq2LcaWB0yUbOasgR
6dEc5KNik3w++4GjhSE/HMwaTouzCOqoxTG6oUdj2xo1pPzCOv/u5lGWlaUxdaWQkGhmMn8vwTiF
nR3hCY1dE+4r9M9urmDP636rw0OdmjW8P1nTdorIkyRPao+3K36ppIW75rcliz4NZhwWwyUKPmxU
SnkuEu24hlwnukdKRBFW5Us+4PRe0PP8BQUtjLF9ePEnrzFqAw5dgS73vg5CTGMwaIlvEn7ZHMaE
cq5OXxHW+9n2XKncBxvcnqUVVo4OBp64ZWlHfFdhmurxYVtIy9bNP/dYFbhNnOPtvjPV6IuSIjjI
FCHj2izrNgHgbefzEZkLGHWx3fmzEMAqcIX9KkL46fSsuniN8BZphXsgpyTdiDgmJhQDX6y4EJCW
N7gP0oPXoUK+AEUnexKiBr2KPh1+0P7o6qED1R3SBhV5yh4q7NX555xt+7WtZ6bn1lclkCWet7d2
2tTEIJ025/6Te1x4mC6q8rOM8eRdD0o6uwwW2KO2AMHqXfcJ5mxKa7/0l9Avo7A9bgITxqGL8yDA
cDeO46J81o46djcCaHa30Hcj+Ktzs8COnxkaBIhmWRBjsGXk1P/fZxALxFnfhSa+JyFbdFK62LD2
9qHQ5Qd0CXH8pV9J83SkfCzgSWy2/794XpOtVb1bxLR9fdqiUfgEjlRZrvs7XXcNtf9ckGvW+OgU
4AFX//ieHEQaEJuMtZOKbS00XRcql7cq9IUs1u/BSbuPeCdara61JRHZSmtK3YsQ6ajMguufpfsp
v43GdpLgaVC5JLL/ZMe8ji4oEQXW3IM3xD1pQunVbeXBS98FLYyn46HyDm5edjdVAGDFAfq2uPdu
iSTy71TwvcRq/Yb5vHAPyuORcdwsb18rz0xD/IAepgvlwGaR3SkZWb1xX14ILNz46tdjXSW0xZPW
TqWfnF+dD7HDP2Ui+k+G5YAewp5osD6GpI3U7W46+W19qPBeICo5AMhHXiGatkJ+VZicIgT+Ln+B
jTxbltGX0QyaO50FJkCqo+79iHkgCPmnxPP9E3WFCFmS5B8wLVBUuhc9+3c7JYp3R4uz+d64PT8h
rx8msetsGUgVGeQkD7GXlmKxbbZaSmqpl957NHFz/TsBgEnsmqHu4ksUyJ0V/eBKfMjaari+pSOK
csehHSDoBTv98DnwhPanoKv9mR/GhjfVBih8qt4DYB+9oGiKSGwA+waQippS0qR+m/63exGgpzK5
rt1NsGbGRAso/LunGZ8+8i4UXlnW5Df+Lto1Q+QB5V7E/15UHK4Eamywidnf7krBn5PlPhTi8KKg
arTiRVtEmxFYfPhpe/cQ750/YvFgKT3ynmKAOKfKYm11SJMyozMMzMoR5Dow0Cq6qvDYwQqPzwHW
FGuSrHquL4u7fKKxdJfBby5UZ/9ygMMMiIhwGqcdbJArVbW1uXNtcMFhGTmjf2QsAMRv3pTdSeg/
9oqaqFK47zME00+Ydx/515/xXCJaioI0Dhg0wi+RpxQuK8TwGb9CWmkuTNyAaApoEOXTl6M0HVbG
h3Qh23UiE0fgcDOVLFk/sOFiZoMxu16dMW4GoOA7FVacno/AVdOUrjQ5G7fk814ZqUs1gbJz+qjg
LsrKk7hY38C1iKDtyjWJoWmSk8IiGEtxczFFJxjuq2NPX/PcjGRQxsD7KWgTdjmOwvOvuLdC7Q02
fLjzk0grfwJvd3UuRspkwa3UA7dxBvluVtsDXPSKee2webVRVlk0C+N3Xv9Nef7dvVa1Y6CdLphf
IonLcrs6dX3860r6lGizzRw8YJSPt/lf5uRj2Q5IwSP5HHU6AYFRHwnBCkR9c2C557+j9vPxAstF
5WilIMosQBPXzu70ztGoGEy6tupzVbeWh6yrSVCmk9+JXNCnh1RIUyZdBvjFK1LLGjn1BqSmZa+v
+sIdCCw4nm0kDDzLIiP41oGevzfUfxZZki24wzxu8aysxjR0iWq5y24tT5tD4i6j2c7Yy31cXd6G
qZ+BGV9NpXEUq8vkr2uIKxrtMtI/zPniz/VfkS4OPidnQE/agDy98KsTouwvYAmpb2zXzPGEPqhd
NGgBmOjQrY6YsoRkLSFMEwIUX1bhsGp5oIUTF5Lgh8ySKVEsbMpKe/UkmEzi3HiDVYcNgOmrJgZb
BWbrfX+v7n2GRVznVWIvHHAfsv7r5Ne/F5uUF4XZdysjvI7KZ5a0UxXs5mgK/xg5Ma6CNR2UuXT3
kNpTMmavBKQrHd5Cp05ukGyjSzvZHzuv+lLJvsQ9KKH2hJYetQwNKWwuS+moNXd5uvtAuZhb4E1Q
TScFejNBBg1Il5Hp6tQxRz4lnUHUZJJrQgIyUCF18j/RI+h8svnfBOHd1VJaJIqiXq5cVaB5/U6g
4/hCFJNiZq+2VrIYYoYMhVfsGEXwIBNgp3+RxkDcMfAMP8UTPPOEW3YDpp6mxO/hvcei3qqrPaJk
kPBhbmxE4JdnLmyFm71f87sXs3scU/QFdmE/LpK/yV3ODYciZBpVxKDPFkWPY4QK3kxeEwNNNxnr
Y8ikT8sdhlcFfh89oTdF9YSjqTYpJUCyBpS0Av6t3wyOUdl/TlNtAoWpeUc/rtDbhGMH/rzjMZI/
SCRK4l2dlvYgjYj3LXIHnoR2qhw4BAUUW8APVmTo1ZR+5WsEgTKw12ezhE0va37z4dQoQcPpivIh
YCkFLnJmEb+m8K8DqwJ4SCR8SwrMoGBrLTLJmiBgFrCj5Y2ze1kdl3Qrfy5jTcfg5y2LtsoCtvq4
XDNfqifaktls1E5OdEupx+CK9hurEVTVx12Ky7RKapOetiTLpQmkHGADeZGsyno//QAkxnqxJNq0
rrJOBay/hoAMJ41lpolwGJGMVDZkn9JCLcMyYqDsolQfKAtjEDWnUXVjvlsN5jFkO510qkjMY+dZ
2olmYe6ex1u014372tIL/GlrZaTkUtMZXQFJZ2BBRRZ9lMXbB9f+9+fMBothzR1sz7FHto3HmTlU
hK4upg8lHT1iGYcmVB7q6G1BaHRyjzVOudjGv0Xtvi62Arx5dde9ytpp7gz3pJG2lkb0rTV9cQvX
hGV7oZ2Lg5sjVIC4/liffMA/btiG1SQrWO/pdMbc/3L07Hg+cIiWONpYTG6CGymhgINUBDBKMOW7
0u8+JuLEIl4Mem9DL6PLpwPVcKgHcDJYAqt1t2zq1eu4CLlmiYOKh7Zjvy20bOWFMNaoDIzv2AQA
T/O3xcKo8xgbAclANXce86oJ3eD4zdNt8qQDcDSb8UhDBEUToI6zG1aMOpGsyJHFNGXD2yFqENQ0
D7QGBhHgO441piHo086EkUrAyQhBtvqcNRr5o6gJMHZsexhy0Q9qmcLNiWZ9ZhzGQsbn6kKkD6nb
CVYO2RrQLIETNkyHToeh9rv927puyWaWj5hmEzRci5CL37TKDScsLRk20CxAlpgKRBtHchMrLNYc
4AiIWxeRCb55lUslfrzKI/2teOG4P2hBlRH6RX1y6k1RH2d73CmYjsyGh9/S4snyp2vCEwcXxmae
bNz93dB8fAdvbOHN5c1Ank6CbHE1hnEgFOJQ2YtGbuxjAAExxNj20lPUWIG7BIIYd07dK+5yGBVI
osQag+dN/mGSC8/nyYJct974btzBak6tpQv5H5Wu2bpfpTqalZWbbDPH7a282IqcXENTLFrF4je0
D+il2+5fvVd/ogubn/s+yQWG7pc8G1X1b8J+YP+9F0mayef5oCoG0GuoP/X7HrgoMlT8u5ZCcqpY
JastEPygEdHwj/JM5T5A/w900IJxRE7kfliaNCYkXPYOTTr6BqdrjrYK6TQrB6Pzn25/I2lPlvym
J/aZK4wlXbJrcCJUXwHz8Umf2bM0Aqe8j4hX2Nhskn9IEfZ4miK/Vx/aeXs6bzFmmJDjk3wfJ0L7
8VZDfNdyGoRt81jBskywjpXBDODTZmhVJPQnizAQuOmIoi5iqQ9F6qH5G0Vk2QfbXv4G+2z/lcn8
rdenA6pxM2q6MyoXeCie6SRrYCdVTUReEvzO2cSrSpXEahWwnb2+5/Viv0OF3OMW850gMrlP4y8e
pPJoQBQm9SxlKXzLgm9hjVx9rGKF+n1uvnEgN7tWeXN4XtlLKrZ3eLfDV6mU7rE1F2lVvKGMg+w/
V0/ULJjKgcaIselKZVeuVSamzERs/VI083h2wUz433P+EIg4GtcKyfuZ0ULzSe1oVmXRfFbqH2Lr
476+2sP3Cu4MKH5uHElxbDTh/F0vQ/FxN0g1zA0gKa3O2RhEfZD0JhpTL2MlYC2eTHRvRFttjtXq
Kpttlsh5ts4dWv3CISjNbnXITi9sBP/cyGb39p67ds3xlq/8QtMQoXPpDGaAodRsj1u0HyTXrl0c
ZmwmF+uI737lZvVqJi3sbhznjwoX3SuKQmNnCRGgFxy1QjxfogbzSZrzA/mH8SZe1xpnpL/TrYLq
icKHdlEJP5jb0PaIgZLhhl/adJgS5qBIKSicS7ptXBBtkzXaLmfrElbq7hk+3oNgGUamBFhNZ6lY
dhn+s4ZjGXsraQttfc1BIaa4Asr4CjxO+80x8Hd1GfKiSgC9c4mnI4xrAyQCQHEVKhXZCg1Q2oxv
U2Av6Xial/+7nY6jdqZyvvTwRXfJ6V//xjj72lPzuZ85nrt/qBN+pFW9Jz+lvQmWuxpFTXX+vHHB
xnySW4xGcrJiYs2HR61RE5tSAIenWzWcQcMnwMASmz2to+TjOzlyPyVuOhTpbZGFZPAx43fhn5NA
ZVV5mg1xvnFleIF3H8MFz7yXxSaw6RVUARPMcLkcrV2r1u0UGCo+ImFo7oBm1ABacQbI4Pf5fHK+
f5scsPZvtSfQzSz3FNJldlcYdC2K0PVmjJl3fP5TWyCas1YqFqipWfnqO/ATUCepqsCKPZyfI2UZ
s6LwbQrZHaBAhyHDKwfgFbF8nTCxzDFz7P3Y8kfoxRpfZxhDAnHWnVgo+sYVAy5I9cSAnk2M1mav
an/BmGstV2XabNLhsq1C+dUsU1deV2VsIrnDQ52bSijcozTLgmnq/eDi2tqb9dSnW3gBLsS7lO4L
4bvw1EsFVbSUSpXo4/WQBnnHZlwAJuHY0CuMyreUKJX5DwgtWYZMdnFATxwNuy8k3n6QROT36d/c
AJjK5HGXQFZPBLuGXOgxPFQVcQRIkBZzSbgug96qylP/wDvJsE49GuHNvNO/9sJ7Hrb8yScupF2r
J820N4An4IjXIzcPXdNwgO5lC1WtwjBGhOMvll931glUIPvldguWJJHDFWlq7AORqBGb/0hacuZX
oJyThQ+94C8TfG4G/oEN+ktG1hI83o0bkmBputNAUQWiBUIZdZriPLwp/HSlqvzyARO7VHoEiksT
fPgX1fNWKOKDEii9b50xHRH/6UBB70jKyBWaQJ4l+0+arsJGjhlSsHP5GrfpmNBCmK11QeDAhFq/
YY7w72C3HMgbeVcSxSvEQEsteEJmg3P282IimOAoUS6lk2DGQ+gMO7IM5dol/UPVKjwdYjFe4S3l
CTl/anJ0XJXukNK62PokG3BV+3YguLvfeAwvdtiEKNy3Zm8HUkN3lIZV7fbaHNMLmj4kqMzylfdU
HxP/8dNEzUnRrSW8MNN030f9DcCIQTYUMC3Ry0gcyBpplMflJ1j1zfGWmfpEKF/oDeBcstJzF8t7
emE55cyr7hjhP9IPTPJpb8AUzfOTONNcordB4zP5a5vLlvnEetwhUhTDjKTdMyJngrVgBgQq1TL7
S6C7RENZUX/hFMvvjuWEH9Em0gfBBDwlc2BmsniVTgMVIH90s2tY6WMNfmuLR1e8s5TWeBrRzMSg
NWS9Bohj3ABaEjS8Ja5dAh3OQnDqIsAEj8I7F+Om1AFQB6Z50OKYYot+OlGbOu+RlmgGFAIz6Y6d
iRsLkBmFh2DQq6tGvn08OPR9pbthA+I1AIeuOkvgG1IJNj7cnyBGBhGyRTqIAdhrc9QWKLC8SPDM
z2S9W3U1eSSVAxk8f+EyomMRlNI5+1noRosRs5MOYQWENHHqmLAvzu4LjuzSmkJFZ1Hoj1MMDt9p
C5MG1XN8hortAl8cuzBwDuA3wtvAo5PK8FB3OKwKiYhX3/hO0RF1oDnZ60/pCFbXmibjb5HwAk2I
XcrwuQA6xj+ZdLYnE+Y/uCRPPfDnQz5GGm3Z/lw/JciY45W9ig76IKJFI9moalhrwJJTfsDvuTzJ
ujO3JV+XrK5FlNTy7jt09xw9b1llCll3V9K238oYRar6PjGBNoZGYqRI6OBie+ULM+0wQqQDiVdL
IFDBHPsAJZQxFgPvMVE4h5qaA97gSX6ZfelV+lKhLCLD8QFiVG1Q/lfzB6XPvagqRYTwpFsumiYa
JVbHfNeUiZC+0QWmSnnTeWzuJEZspX6xyAgwgWLJZIy1lpSSWEjd48msd/kUESc6DNCJmuTZ4dCv
NTAGYW/M9kQzSwNNWl/opUjQCu1BEQ3TDlPrxGQAL3qw8KpV/ErPZvFcckFT6Np78Kn3LMt8Bf4v
SvcN7ek35XxfTSNpGxgE3iK8uddjCP8B/EC9dEb0eL6HhAB4pJXpufeyo1ZXTcIFbhJAdDxQ8q6R
gFH+380fRoNPCGGAmhhAK/jEDNJT+zkqb+CLpNnltlLnL4JCp8iUkFC2EoH0BNT7hxT5fcg6Wjs1
4nUZ12/jem+nIQALlvv88zOnoQrhDKhtq0oA8LQ5dNilSsZMWA0sE5yUereg0m0XnpO6eLIZ5q65
9eOhoinH4inHCarBDFThZM8C36O16kMUxD8M+K/XVEZsr6xOOKeYgHMgXQieEF/vKX3fLYJL6mg1
8UDlq8VxpsYXRYQcam6yNPao+57x1wet5+Nn+0YtLIMVzbcg0wgbeTPLetnpgRK27mFsmFYcsT2/
RlYb8UBkUI2ldvO/5YxpoqRC1mWxHHo/XzGOBtuDAf3TfgcyEHYFz+pM882uodsw3Eoa5Y/xirjt
nWymqfBw9Q57pDwZos6BInfX2ShMTABFmqGH3MBAW6UmNiPcV4cigcUGDskHi8euQwwz/Et7rlzz
QNopwSmHZ6xQ6CEJUzHGflSv7KE4NGYYxMVQrjlco3jr2xdqZ2EcU1YT4dpcwwcQb9fqoU0+umXq
qOAn+yRpM4krpkDKEABbUNwjfbhdjaWed55P8imQC4zUk4NVHICovRJHx6euwgZqKj35QmrYZdLz
GCahtG7BEP6yO5vRqNFQ+iQjnZlCdBDzoPfQVSJqUFRFQpDcndufb6kbsH63m30Fv1VESEo7ms+S
qgX1WfrVQ/EW5nxlco4kt1LGcPpOaasmv5FduD18FKtI7n4aANkUKdSH8TqhZHNr5BtsKj8XxduB
qH6OrhHgHm0TNWu4B3aj94YB79jwnod4ZFctNsateXWqyvjMquUPTr/F6bYXDltgsOvFfG87x01G
ztW009OB4D/4vMieuBJsp8QOVyzaBcA6ZswHSsV+45AF9wTw5D9fgq3tm6uXl/aS1hOBZxZZc4C9
2X77RIqCf95jK+gwElBKkDAwfelDN9LWKWJubwB3NTBO6Tynj6PVDdf1vik1g2dy657rXslzqzxR
LtcRbaDaZ61RU0k4Qxvf9K9RIIvvROLglC2vjIHTXv2n+J3rihzfjFeBEwkWs5E/A8z12U1B5Okg
aQ93ReH34eqHhilVVlsEpbxBbLzDTfQnkt/Gm82KZCQsZIm8MwBjCusmPCIfRtdJSb9BqpXGqvBV
xunF7ASD0+1WG+jDyIG0mLcbEauhxE862hLvzKi0CNG+nusOGHh+a3ATsdl92jsqT7D0mE/2wemn
TLcy7D1EeBHhqwv+bkEreOQeEVrz9G500MZypdAxb/IaC51wdjXsNpxRX60cTvsAiwN28yiNHTss
bQAvcqDIof4I6xmwXhrXZPNILl/kYJUl6WMfJocq5pRyAWvV5rWjfhDAriwp14eQ+6tlI/5febF5
ALVu6+mfAEuk6iviC5461gwbmjR2YlSnR2EFHTf8Tj1O0jGb7siMu+PbmS99BAQi0MGCiOZKGhe6
vJ75y57xqf+j/60PIdhoCn9zVmxoS/hAuv7xlJGG6K9jqVgmx5T8/G23Lx/UEthDnOlils9Wzqhg
KrnhEZbzVCnQJp373fbZbmAlKAxA6/AvvUQPi6vE3yVyFcsy3qrXmZ2eyT2JNbyaTWXOjkOXhEJs
F4Fz+/VqWd3QkIIqUsTlnz+XyGBkYcRhNuQyPs4zyV8iC9frYff5I9V1D/6nA/bdPA3qAsnGfF7a
rTCxaGsGhZEj/DUToBXr/rwS83Dl2y+E7gmWnpUP16cw3BZ/XF6wbXnLDMYNmC5fbT0HMJQBZLAX
iyGD+MvNnhWMdvlPzvSMOaZyQ8tSsqyZKwWe7CizK3ofYfvTsCA/82gh1daPx3xNTtZaq3OipmoC
xKKA6uGuRMvUp8gD7zrEf8xEBG6CEoYoL4RxWoLKBQx48P5+LxF5xtiPhtSTtYXNwfBb+YIlNBhr
1Aa2TEDHP4fwvS6t23kevXtFgF1OIgVchZa3j++Lj/LXhbxccc/TSlNzCqvlsHLywFudEo7xbb4l
yuhqC3plH3wHxdUn4OMMiJKtjE4wUrz4fo5Mxcgeu9bBQT8X+ZmkQ+ytgxxyvKkuFOgR4hfgfgiG
Vsqok1e5Hwygw3kV6P+9/QTN0i27L07SjE5yx2HEbR40sZ63pN0qzPDseCfXu1UqJayHQvXWK//8
Qy+FghNdB9+/wBKwswI8Xw0HZIIGOGBLnsRvr8dZf+LafCdtHOErXTN+dw7RdJEAJvtoZJeavYWr
NCNugq0ork4mbshAgXxHhgyYNExBv5s3+7BgQ4BswJe4AHKNMA+8koJ2UHMXFcaPIkDQjxKz1loB
EgSt4gy5K3QFegdXx76E8gWFFsl1ruWz9XChqoYuQBDyx1s/m/YNMod/p6VMh7CCY/pwhURKzJB8
lEfWlnnh1MLUpDQLtWr3EVVEWcJV91F/DAKxLnUf9OT8CYpVD3H5ichhYlxaO1+PqywGvFmmIrVl
rcFN0823g0tYzWf7IxlgLJuMfoYuD1WP5GXqJFWRhBpdox5GgGVp04GPyWJetz64Qvi9ziCDSoHJ
11Nv9l+JXQBe5dne1k0bl5A5vQBexX3vtI3Qv7wdQegs/62kWyTym3ahHIhkBf6oP+9PHNCfLd5b
QaFq07fVQegQ9m6lEbA5VDUa/rw3csM1aSs04l0YWw6UkKj1Aj5JAt92+BgW8Y5dfTW3+CNh+dqf
mxa67ddV9H1XIpk1RWkH07rAdz/AFKytW4FIsPbMVGiELc9FBLuuz54LAUGVvtWPlhdyCgrCykV0
zgV07k8Ix8GKZG36UP5OMmUVoHbprGLDN9MoSUt0dw907I9bkAxX14sO6iJFvhLeCnmKP3pFvheh
MDR9LGQ9rOHSr1vjY6QPK+z2LfxEicS8gf5sCcaE2X7OdAz4qLOO8VLsGPv32EbFbUNrd+AOUZg4
OQnfkb31AIn6eL915tKHTf0nlWtu4PEL2tsI1FRXduPgCgJNcsPViRXwlDfLxJmQ59uDDnbnAmmE
M3PmB7fmPBCId/NykGkHONU+KZkSqMLzECqWBwvbdxBzfyL1cI9WkOXCaEYp0uEUQ76ChcvMOmo1
UuLJNDHF39wlZXhlMKKIsdZni9v6mRJwjNV+8dPahsu+0OpYeicKL0qkLsK5koEze40R06TzcG/E
zoC2Xe7DxEU+xegH/QX+YRllXjwxidx8FNqmHPtjVtaEFoseTRkAZVS05rsT+H9kF0xUF+Icgj0r
hiWQS1Abf1GYT/Xe4p+AtiIfgz4aOzSb5miFZH2V+eRZLMqX89ABgXAFTtV3kRUZD1ozFhFKyM6J
VTw3XCJdDPftoE4L5cxIaBsuCtgiWJ48O/chutr2Eyg2d9tVuCi5JI2XdXMR/EXsGAxNI2ujtWk8
hcjvAXRTkljTK3C5BqARJutuFwG+ek4iBoHy+c5d11UWf+DY0Ievw63XffMcCJVbr9FH7s0gcNy+
MWEWJM6RSY1yPT/djDWJtxck8EyooWFxT43MsXLLOC2F7a3hbyn/8v1nwHsb8GoTR6DKXRCfP/NW
4/+vv340zx9PQ6R8t0pc776Sd4C+2y6+gqoD/etfiuNifwSUbFKI9IHd2RAsyOG0HBh4WFMGzHRs
/sTwV7xYIfTPbN/91yqKgIrYF6xbMqxan/hBFxv9w1vxKGFFLOpNgOYccqMKTSCLiEeTj5FoQnZK
Icj5fspi3vj4OJWzVSPZJZWkHj+Yl25vlMd7Cwy4dPkzrzM7A8ouKj4BvqLoyJ+aPe3lC35ZHpVO
CIJ3tB00avV6/XKB6CgIvM/8/gysT1gLWyJPnmlLBBIrClM9WVT7Ez+dg3cdBnALluYqYEF+MPI6
je3RpZEwEkhx+5RbhnjSAiLiwLoZ9HM5l88HdZ5HXeY4QfpEC3k6KKt3nWKvvWca9NeiNrlBg8C6
rvpR1OJqU368XyLtOAEUjgtqJwPhm1i3IdUZ/FlshWc/1Pcot/KS7PKgdvWu4WAZqbGUGDsXY3ce
U36uPmgfQsQUvxOkSyPU4cfwfWV4q1juZZYFyy5i9J1WVhNVBkXor1juATNLXt5wREPL4HoQlKRC
MSXHwypN1MhTVTvpAdTQgk6rs3Ni9MgNfY+QQU7iuknksBTlOxPh0AYG9LQGhRC3E4EA2K/0c4Kw
E/HFVCw0G5mTO4T0Iid0mofjo20QzAusGHOfVaWx2IkQCXckQNl02jpp/9n9MLy7xJgaP3bAAS4V
tEuiJF3G0Uj8M3sZaNGLkQvYhMvZ8nuzhp4tNrXnvLX9Rh504I9vvp638WtTaQwKaGhVgvgbMUCj
tna9r+x5/rAh/5TDC6iQnCiV/FmnYf0nykmyHnPkN/MkGI3/xW2evJbzOZaJ8F8agyR6M062aGB0
HQ/pAq9cPaaHlrgbXIqUjopHKMOIvT7L69fJxmdSqgtOuuW3vq8Hr4vaYUBmWrmFqrTQp7pXFItR
6WL/UKfdgYEadxbe/HTu5lv0jdy2gdjsz5Ca07UFvk5w2aHYjEcOWIMGi4LSE0oGRd829PAE8QU3
s2Ry+0IiAeEblYMW1jmzINibrzw67qekh3BNEuU7vcZoTBnUcmi/pxe615CKGHUEBiLPg/v0znhW
g/CF4v0VIDg1vqYiwWr3+whVOodV71+xYgsK55Gii96fTHEbtNsDRH7NSFl+s+4x37lRN4WS+AS9
Dr1utWxckWv2o769VX9ZrYoYGbSF4Q592a+ckmxOYm4cD4HNwL4hph5LspxmDPkViKPSeLHbD6gK
+f+RP3dlUPjVY3TwkSSdGB6VaGMGH2pw7bJDy+V26pxtNDODNeD2YDtPEtThQ5ZrqUFGfMlypwCZ
ACFDDITW1ArpLGEfqDi4W7vlX4HdRAsokEravIef9hXhoFJiQR8j9K3n/cmqVBkQ1YZkiq7PD//K
KNulbUaz2SLCc+731v3KARvRTvu5UIBK1z52ZvYZ9iA7c9KuVG5VKQ1IxNmkTeDdEzz3PZrHW4Cf
og9939ikmKH4iEk7VCuFSsh+RLsYsr4FfEPHu+oPv4Qx5/iswogAWCQdZe82uZXlplieqH3QzHYA
FZv4RuY3CVf/l9hO1GA0sfwx3SjZMR/MskjkeoIgyGgy61gYBdFZQ0sKADkQDNt7p6RgDVc2hK8+
YBBuD2zSvO63ScaP7EjI0uw06/7aYbqR38Et2Vnfb9n1gz8JUr4t+NOt4jN+q5XZcZUXY5Yogdmc
NO9tB27Q9apwfJgfZqPTr9fjupM7YAo7IrpUNIHMwfkDKseYY0vSJwMpYn3XObZYjpXvS9Q/4PZf
+rgWwK7XLM0Z1TsrLE5oAEwezkx3HtLZMqBGMtI3NEB/2sA5hfO616eBDfN2MqBbN9Xn0q6guCP+
p40r+H1BYrOFThUDQiLfbd/vW6C5bSDwM1ZrUHk5VkLRPJkjDekqS0478IT55296gPIFPJzAR6u1
3GaqLqfiiDInLFdOxqJZoym2RYT8K8TKfrW06AY9LJ+BmG9XHNPf4zmdqh+rndqi0T0RiXJ2jvYf
edlJ9bX+0gf0b72vMc6KM4rKQ8lf7+5Xa4aQXfbYFOkqpEkIb4qbUHka8zmRQCJjYUKVKJ0SF6aV
Blyxlh6BJBw/5PsSKuxyvDd+G/5FJFROLwVvE9R6Q9Ljb6m15B+OZ4rbe/l1vAEoKpkppa8bAJbx
Iy5qr+j8FyNz4jd5O22oo0JnCMcCAUsr/sVXun0Dna1OWq5v5aRa7zKItm7osrOQoTlUw4oMOvug
n/u0TzCPonvMWmeFlaGcK+C9LPBpZmF7+3KE1l03YwcOlEuPXD8xu7n/ItCj37aMV/U92tbyYMq8
ZoFmsZSbOY9+A6ReNZ7CEWndKZxm45Span1x4VSAmZ/lqFlwsOrTsElP5BndgFpgz1mfid1Nc5qw
n+6wgsqCvG34WNCZ/AdOx8hHN+PtvubhfbGPa4LMauDkDamuy43c4isaFHLKvN5psIg+HoJd1Im2
sf30wMEqSKCd+vJO4VLY9ix/LJ0HmQPsCrx4EDnuuBbj9Qbb5cOA8IVW+R2JBTBDOFaWoqXW80cY
/CxtlAGZIxM9FP8BllKH8l4IAc/nl9mZWoBytAcQf68WyM1bUSbQSszKE26Z2u1SO48X/Yan4qMG
CpMCbD46DWT1NTyOQdDO0NBdV62oUcHnNY7TfgpifbJ2rN2xclLR0pdT4R6i3KvR6HHV87miOQyU
1JpQlYWiwUYaaIdN8ipC2cf/Sjtr6rw4b/tN9MIOeC9nLlY9kmbXYdZu8lybKa41n42Bjuw+Mrus
8wWnOqFUrY82gJzNtvuyHr/EXMEa8JNHcXL3oMBhL4j68/yaHKBb/H0ipNt6tXk1pEZ6r1aDq3On
92AAS9K23h44Tc7yYr0GqBHFA8NO/RjiOXmbcfvQI4QL/nWojfFu0Up7tFxCPGNCG5+kwneQqI0U
Sde/cDwyNnvEscBDfC0GGm9HAhZR6ZvnOlECivak4YVYBlMtH7eF+syArI8TXN3kMH5jo7+Us7Kz
NQZ0+olXYSBzQSod1qi80fhWHqwblVRQIhcK58MdXfHIskm05Ekow+EtwbX17ZDfjhPFPNyczQQK
hJYSGFs04+N45ZrTnZjtaEshgWtBXCWvYKT+bObCf5tZXv8KYMQsfGYAN2PgR+nw4VFU42/ssYaE
F/7+5Q3pJQVZZDAnNtHL9TBGhCHUmt0gZrXVKRmrdt820zwb7yz1mFAT9Y7sjEqFUMyPiy/mmUJi
EuGm8W8kQntVQfa6T84qOq0HYRkVHuW10PFsC8N72Vn/VRopTU+cCwz921uDYXWFYTwulqTKKbVZ
R9AYcpPyVCcNA9wolKg+u0iDdS7JzzZ1S+eHX5mi+5LbKOxcPHtYmO93+EXgIVXrWOENbrEbKDRy
HEIZbc+EFkhV3krowh84Tyt8MNk+5hQ8FI8KvF/BYHQNQ+pm9zOkX7GpEwK4vzQNXSuJ9+uGkewZ
EnRbW+WgowrT0S0uWQU25+udSOJpt2yPiq6hCCvEL3M5Gr35TtAPOvQCsjMm1YfqCgCvgo5ZHXnQ
jer+HYTBjAZXbO884HcJ+pXop83WQcpDnGhAmS2khw/M64idF+o1Cy3YrfOsvL1OnRzRPY8l6jmP
PGz+vl3bUylocR2Al//rqI4Y5eoC0Xy7NiQNN0hK2GZZkrG0cKlKdfOlMvEQKJFezoLr++WSME6z
aLrjNVMzKxO77383rfc6egEy+cnH1urZIJm6rpjDxnp1kQvWO5/afB5CYRGUZFZGRHqU/4+MDGdT
32mJE1T2P9BdID+ZaOnHaXSKxrDXcVXLfrPsxObJKrXb5nOVdA3Pk4OjNRTbIMILOxKm6LvAWivX
l9rBvlF9WPq6Sb/b89tjxDHll2HKqjz52ggM8XZOnfmUHxdMzYGlJtgWVyFhzh80JJFZJ7nmzvWs
VF+NuiVR4ejqAr3kh448+rSAn/gD5sgwQLK3UXGrI0C9xql6Xk74KeLCyHPzm2Im+7Dy8JyldUSI
87vdDF7qc6YPYFrNCUldnxZHKx51mhCegbxYLDa5SzOgR4rcXgpOnV8pRhnrIQ6bav8QIcjPmyI4
6r/JwiofVC9Ni4Tl9JTBHhUBqlqS1ZSKk8SyCJRyjjrVNlLvSMLyNwzjImAC4matNMxw5ZH/wCN8
zOgNu7vOy8KsxBF59rZ1cr1yHWTmlqIL1ay25ZxLCgiz3JunaOok98iTJiwjJTdgPUpFvDgxnDz4
LRr1eQeZgybevbDqsvBW26tfhaCJDupsQjvoymyOsyhkPcU0dnMZH0tehauQvjpGWbiPJPLRAqxx
/pFD6ugbRDaEaPRi3lXLlWxvgR2zKXPx/ZkBqJlOV1Hva/AeF7uvUQl2PIm5sdj/aZFOlMk8Wby7
rVOJUUkh3VX7ie2J2XptjhfFFIYW5o5ZTfZ79RS8x8LqIbGvtQYoJ2lkggcxHGoJlV9XyCXjqfHs
Uck1k7ch9bb/hWT/lVSmv1AtSJLtq4TwN/kdaAEnxTF8Ex76MYYmzrJHwfWrzFOcKwFfDKrfg8bf
LLxgq22rnVe48AC81K2/8onaUUD0PqvUObOwQHUqwSxZ62/y6r2KVAIK4ZKGz+DzlbIyEwZ9cw23
EfUWAu+0OkqswiqVAvx+TQdXPslfnEh/SAwjif9bdYdMi+lUl1dDeN3NMX5XEFDYbuucdAsKkE1A
Aj+JJ/VfC3PZI62t51ofc1+FWm49ddtvciSBFotVq599NTLKEPL9p/XVy72IBpilSyVkqHbm/Vgk
3tawCUSPgBxjimCigFaOTfQI3vsjj/NZNfQiF/Ygr3HtB+uCMBoAiKgxr9yEzRiU+KGeX53SHjQn
5TAUrmzYAbOcZmpZwuWbtzcQyg2jN2nDFdGeKw0tfIuNksHX5Y3uKYK10XbN6zkL1awlOBv4kAee
TQGpOnVkJOMLyu4vzIV438mBI5un7MlA/MMSK6pGuQgaTMKzaeAuUYNndM7jgPuntby1Hb5biOK6
DcIiYUebM9I9lqaFipnH+Rs4pOjH46fqeZ2cXX9CQqGi782jJpOCebwNw+V/2ASdKaBj8aZHGxjD
xlTZNrKSewlfunAeJmgjIGKNrE8isiP0GS93bVuqkwNTfabCJ3KZZHt2IMbRAWrco5TZufHHgla3
6BelMwvPbxRkagLRqi///ba+OfmrUuOZObA61NuQqVFHGEIXy5A3pESZrJj+mBJo8IN8rNb9e/My
nsE08VB3KIl28SQbAP5iQtCrlGyhh2SJOlFGYO3q+Njj+/rBZ+YLkGL5rqjPhwOOvq6HAYAutosA
P3PlrKXWQThgcR4EVMbjNlCUjkpivu+hxt9rVrF3stPRJrINWwgpIuSN13pJcQU0bNh75Eexfrqa
ejuH+zJzfkExrP25YPhAx/08o2ZopqVhKsFgpiCl/COCIx8NoQ6wLTrtBjKjPIfh3uXgnaPTD50Z
osDjT8IMb6Ws+0ASilQ1Il5oLHQTJEMRgu96CC5al7envQxEJFQYK8UDWvEKtbz5sSpqFNVLhPe3
B3zvPxZC6H/ycJ9uuOAUyUtIYtPvNftatrRQT+RRqDP4QoaRyfeAE6L2tKVtfqflLZvxite80IaO
byrwWYatUyN+4bp7a0UY5nzyZiuKc0AItzBKpFHS2IIuAlz/vHqLgp9neXRohQoIVKbsp4w3pIES
6/LesgqRlbi/gn8cYT7FuCSjJTRvdq7plMALhMNJqXdjDL61VWvrMJWsUMXMrf+JkUH+M8Gpa4tz
jtfDNjU8KJlMEB43Ce6CuKGOYj3lpZhoYsMGra7puOHO+HWBI90DyzJm9eTVDqE/UOObBneU5HRa
uexc8ob349F343zAVY9Du2Lb8vNHvfPA9qEJ6QEv7oUjhc9Khu7mCWM47r1/fSwLhbljZAS4lb/1
V+E/3SU+AKtE8YgCWFmNlWQY0EPvz5jVInCg3XlkIBOKy9Ihi9qMvu0T/Dwu5fFTcPwyggflcySo
4AoL3V2Sv9+7wco1h+th0YQXaDOTmgsXiwXqaTI/vAJ+117P/9ZKxPXxsdKy4oW5CcoDP2FmSfDU
+dAhCfraIOUcQVaVivOQZeWlCPcqQLu8vG1UrCiX4PRlvgRLJfqGRVO0GAUG2vgKnXQRR5KrA/9U
jw9LVjurMXUM+4h7VEVsWEXMIhlHeqzD5/llV0MZSwuHWb2ylahXYrLClBM01bNLwi5Gq0I8WHtH
XB5b+LwXW4YJRNPAnRkLZlq08qpuGTCOfkaI7XddgWmbtRYWJuHx2u5lxqR5+hBl5r1CltQNyPNp
LdScHfimFqedVyEaRR4Ns1HBaqaLxJgUMM/z6oH7+dt5x/Vcf6xiuUpmXkvqv/Ept7ks/cpq4j4g
1Ku6n9XeOoQbmTBvg/IPHuRd4bFJXStfe5olryR/WENwIHS2aX0Nmx5YjT55+ZoP66Qj4n9fhYf/
fgD3GrfUzrB2lQrDZCBdPDwwAy86YDCSm0LZWCiWc/RA25YY5BZHlsbsZU66wB5LqjvoxMUtfBVR
12ozn6DMK+zntMD8HFv8kuiKd0jcHrLqFzNl6IJyOYUonNSLg0zUX6lM/LL3/DLD+LF4qiQ2djhq
1LBrmf9XuDnHqfIQ5hncHsvXI/xRyKOFYALh5lg2tSRcde6qkHdaUKMAzWtEQmTpfslK4WcXpk1T
3ehdYdvV7p9DRTeRrE3bb7FZwlrPXk0JGqOISmpo6UD0NGRt2nd+/7l+/P6HhgV+QG4MHCDB4aa1
CNn5usqR4SZwPazWsRVyGHJfeoUlHYPwqly4hPC9XIHwou+djZ3vtFM0yUeBoXBfFTZxq8scFZv7
Wqk47rABV5BtavyMGJ6VIfhDp80YEi8BWUiWPPZ/IkQuu0kWwpGDl/W1dU48W6+h9ND0oQveMTgx
02TjGgyrYipANzifzP5a9XLu/hlOqzCbcLu1P83UxvIcRjsB/cG/N4G6Gy0m7Fqed1ou6feP4dmS
Y9c7fVbhkOMdQVNfj/9TbxJI2joaT5OKQ8C8P93onpq3W1dDTLKwxlUVI+lvg6pLsvLupQ3N7q4G
IN4tp/ziiNTt/YodjTxc3OinYcOf6pg9L8RD/gXG8cGpHx5wf6SPzJWJYLNHi3oCxCCsOMo+esNh
Rkj4EhzAk4KWO99ihoNPAmyey8RuQciM1cnZi16VrThYhSr7pa0Nt0DIcJw/qvuzMvEP5/tMr44N
HvipHqpHtEOQ0xiigpb4Ksnwv37tS0cbkfSiqzhcMcS7rT/hQQYfwNE6HocGykvtfWsSZDtATLE4
+ORyxtqA/43Kc5sJJbz0z3Q3c7DyPTtecL6iaDn0U3kRM/sAYBw3VIUkVKArc9rpa/mu1wslNr/S
+H0vvOUCklWrjoJy6J31kWAzY8FbQnTARfmlkgjUtfLzLvRQ3pEFelgl6JJFaDBB9xSlocw/0W8B
ac49t7OP4vIn4PEWE6T2Js0Dv8HcXI28ToxECthRb+IsfTdhcCDUWh7AL1PXTeqmCfOBCSyAKyLj
iWdKmyHOflTsp3TZcMBZnwOkLofCqtQiq3xE0D/dEusbCcPrQzoHxBpLdKKLrnN24+Ni/znL6OoS
CKzSiInspObfd+se/cAJx/Z4gQO+QirLfHOXg4P0Gw5MrVvTZSdrIO/lyh9mDMdHTx55NQtU+LSn
3k9BOOlrjfudgx7uagdp1teV/s57n5P6HnuuaDaYw9v69wS19bcQoXBl7jL6bPDirKJy4SgiNe+M
/8yeJ/U0Z4vrikt8UIxg89FBP8DuG8JIxtBBvvlKtrEcmi0M9xdUayU3S8myw+nFimoRI7GIizl0
nJ/TRa3WiabatYYfVdtJd9i9EzuDDk7CATMbdUSvpDHi6WYqEdbSsKJALJKFK+suzY2nUkeAbFt1
M1+Km6UVJtRNcTj45Jwy+fMbU/nc0oOP839srnbQglgBYkb+SjSOIk42AhYcVTuqsQFQQC/0OVC9
UJK/+P7Fzup97OcF8Q512EwkctNXM7fpjLW8Vi0cJFlmSgBmFQ51dnzjB3dHSK17av32zQG6trLa
1Bi8yim/mHwxBt3g5Lr/W58vAUmJ2Yzg+juBqaNfmnjV5ln8Kr8e9wmzQm0z08s2gKc7G844XC2R
aUkC3GybyvBa66SjAMZlzSAFpcGZ8Z57is3wr8g56cBZZfHhKyD7+KOHIkDkPqMCbvbxzZJE5L7P
soaakmlu8i1A3QEex+er4+9WXr8a3MP7TXlJw/BKmUeEq4PWc34yLrW+1vbDxUvMTfqmy+kxW1/c
qKeprrGhnx5FI59CDrCd1GzMDFNLhA4D65NaGnq3aTbdGP4DRNAeC2mX7Ez9KgE9PFIo+pG4quiw
/rkt+fphYrKefpkVuKFKUQ1aSXwpgW8/G9yvR67mu0jeEfwzftWLqYCj7Bb6hGtL9KrthoriPubF
mSSCAVjG2k0N03Pjd3ESt24S2yRV9MgD4/TCSSzbIMjU+wqohCFpDNaxrPXs3MgGhDXO4wZrNdQV
KriHQ/7wIhgDfALVVT8uAtf9IfyQNZf6OXNetkjiqhyNBKHlICI7aqgXSrKl+Uo+/HgpYWxvG3Yg
ziV1jxUaqqlQmChkQ8wczIQeEJdvqMGjTJYvbIO5KQGscuN8kkPNU0ChPOTDBMIUc915D55p3xCa
JuHFvnRct9eDRtgzg+CQtS0mStXL2+JEKaNtZSNc0KmWOnek27hZqKZiN3QCDOrroyr/nGgAwd/S
7kH//LosP31i5tEPIYlJNaCo+/0Nv69X0r96vRHlr2LBmOhlOmuIE/sMeF+5xWePUq5EwNFi2n8H
snUiOyC769FKHkJb5XI62jWXlvBMpvHleEtFdRK8pxQGo6Bh6GuzT9BHFiIFGiW9fK7sPOezdue2
fMT1mEWasBNRyY/uTsdKCE/VOFp61dKU5NTzzs9tCp4rGP4KU6iVQAgGfwdlVmRY3Xz3wAb5EPTt
V/is1ywjSOGFrRxJP0J0EeFQnB3aCD2jw7BzOeZjbyX02pgQn5WBHAp9xLZNP1OTb0KEo7/c01qm
l5ERfsAkBImWaHI6nd1Dc+OUnSQJJ8cHqscn7HE86g1lREPvnMtB8Z36zbHU+wirAIMoqbwoV2kQ
k3kKgCC9MshBIRbUp21ceponjpwIwhNHOtiMbEVgYmd8OLX6LCFW4k3lWDPbQxaZV7XnXsVPDIML
vzLvI6a0wDYB2UwGQBjCBNYFEvCPOdqVRPwQfmeCw/3ZmwqsHK7CbRGPu3rRhFuLcHKfaBjP8yJL
Qb1fiQo9WDmHynIpKblMvFIqReO4Fv5graSnx2fCg+1N5K3sVwkPhrHbxriAt72KNwdaIcC/4Sik
nJ6eFPR2bEjTmzZFO+MXnNIzkYzLO8BFbY8X/Eqyzv8LeTSweCuu59HHZNVyernzxIVsp34/ju9Y
akOioj/UfQtZx5DhjLzGoSwDqbzbCb/TyzHSiO1e5AD4XMBFn29PQS4D598Tn1zDVHYeMGomv69Z
NxsHr9MN7HX0Lf6Om5j/jgsz84f/afG+vFPeXukHYwUr+9WAl6RWJbfFmYFCQ2kztuT/5mkmwFXe
N5uklPys3qBD2pDPhEMsiTm5pWku/WOfoeW4JlNcnkT+YW9yZ2k0RUEdswoUfh1uRkWaA5HeIML7
R9Lwn5j6TgmNGCxHIQIGQRB+wCAbFAxX+NSfSQAmg831lHK8jheZgAR35BmVcMM0ZM44GyTo7Cm/
jBBAGhmw/ih97KEK+mq1GzMjH9Vk6PIEP0uhkRpy3qXWZqBMH8gB5pdlxCQN4n/EBEt15j/s5PYX
Kj34b2oJ17vHgp3ak2Io8ySmEY/3QchT/v0hJMJGo1eTmwT/klO++mJB/THCqDiWQBOku33TWVbe
XsCZ6txc2fHszJ3gXGniHhw6NC8KbF5bV4C1b8Rqt7VXZbbUY6TJ9Gqk9g/Rprb82a0z7ap7ogfc
RcaCNTe6wt9UpkU9yVMrIUGzQHmLB6lG9aY6EMFlbve+OWlBuFC+xGrJ6klvI5ySdU0LpLMsJ1NV
Dwi6j41mWG5URxbS/LvJunMH6uFZew8IU0t0rdnOHRFHPCm2nL+NJwd6DHAXGSRuOnSXns5nICr9
T/LzjxJZ83Sb/ejSf3msn5kgWTsYBkkdoAQQ1uIkbSMweN9xO/wgw4oyTyaBF3TFfz+0JsCRThEw
iJjHhDgamfu45/cTf63UuNkGf+pjFUI4X4iOEF80UXbGXj0bnFlkoAktw7hgftYm8ZmOJv90RXlX
7/cwR1M01guWyY/QDqiWbUNdpnObBtqUZboeAU4C5c7CcdWplUV6cBF5QQWabmGVwefEZOEdu1kI
GVxky1hT3omh69JFZx0pgbTdohrMs0gW8OMvzXrXvEIge7yljxS/u23Nw3dwkCuh5/cBl8x3BUR7
xohLdXb5FwMTH9V8IsUuh7jR7x4UbbMBX6Y2hLLnDMyOU6Y4MICB0HOKxy7FV0Y/UTnmqRwPYQrv
L6965d19gsCPZQnVocXXpHC5BTrB1/Cl3RngRCGELR7bcFWwEkxReIVMxa6U9Dya46WrNnVgUey5
OzGPLazN4jmXyZOkO33gcprDJKJMJoJvxfMnClAoBmb+YhJcG8N0Ma3NqEkTYnfRL8KITBPQltEi
+/jCo44TjVqmllmpJfKzFNx8jws0sYnpWrJd4HGv5mBHul8EWeDKy2x1xue8mGYf//ITyc88Ddj3
F22jkQply1C5hVSPPATfgBoFsNTnTzVBI4/hzMm2Tj//9RQWK8+ekmLVT/fDz3r0zNeWh322usjp
MkwJqbagcbdGw3WVhThUyDjoGJZAbvayxxKtBXpH4adQLhYvpawmlCaVFCRW4O8btBiod2VXcG1h
V2h45P8counSSuZtZ1ffNRljmnIzUl7EqzusPBasdVWyKJTILkF0Gdgs38KuT3VpccUZW2/Ge0R+
yi8sBAM4OEtd3++Z9na71jKc/BAgvalXkZVETyhmbZvfmLdT26HJ+EovOZjK4yShIzwRp6eXDdPr
XnFUGORmJ44gRzz+DlZLY+ASCHXejCKRXCjEiEDa841Rz2FITTOa8vc4JI4xvvylpTYgdUal8Qy/
FvLKJJ41I0/zhwujUZAEe+qcO2b1QxDddSmic/b3EwFSMZHs5bVImvIUZhQDP0cfHssDJNMjEj9L
kEBHFuZhVITbMK3G/neDnuEVd0RbgTEvWQAznpdO2apriLwPeT4cO8dRf1SeuHDmJPHz1PGm4dSg
FNJa5JkBfX5aWovfkjZxfCKqdtC8irt720veCllz0R2hNNMWg1DmKN0c6A/LrtP0Zfl0wUzopb8J
7pcLBAnZAwcBWa+3w2FcHIPfCZ3h6eKTj3UP+pGPUaVtjXbBvji/EHNb8M/Ll1Z0JnFGEaXEZCxR
78XbkHRgSlQK5KHF3KWti+Fj2juqj2e+vr2PPCfSlpGM8vBu6tUQuVyxA1dRVcGj455bQZMH/hp0
xmdQu1JO6xiWmGz5yuIXtYhZng1DZlhsFGJxZCEDkRqAhxRmzEFA6YidiFDkF3GB6TEwBw72pjSk
AQYup0Ybh9PRDf1o4GP1UoJ+H1M/FiLMkh/S9QZQp+rcVbzGtl0YknLWuz48bD0hxLO9jlyAbr9I
YPiCqaFSHqxOIc9xzPxEIX9CeVsR1k1Fse4uunWZuX3RYrWk5a5z8meC/AJD9qnjZ7w/EnZwng6D
QGwKVP6bLfkFP5DqqDUOm2QVsA4u7NoMiyVLrvJojJz8C6xc5lcFva/0F/hvUCZMZnc0CXDMDROq
PSxtcFlzSTSIxmSbzvaLokwG88ONIraNksT6OeY0ZpUnypIfUH+JEl3zGKqPY6b70FSGXkzOCqBM
Uaq7VkY5zLjjDU5N4p5ch2EYU6aJY2c6a8036Nyyw/V8bDJIn3G4kVooVQ64Jb7qTv6SovNH8u8c
aLBSX5V+tdU7W6Cq7i1YQuA9BnUeCPu+OAe9w+IXS96pMVVy+hJ6MjFLx1nHTfD3sNj/OZEbUcsC
tJLcNN0vF+fr8VfcU/IbJeE54j3wfJPzqRKguoxklmpgZ+Z8dKDTUA4ilQgLM0i8YhCgE7WlC9B5
FXu5zXdF3wdJiibzgqSQ6zmJhVSRhg3Zys0ar37vfBBl0O/UU168PofTm6y18Fj0K+ygYyxN+pgF
bMM/0wX3S5+UxEdyUU/dEi6uureZAJOOV02lWOKq3RQ670IIVoEbHknGo5a6Jq+j57FFnEJGO4da
wDAJKvMhyKdDcDddDzNdMYNvUy+BTJpqi6bv4nw9wjVqB7d29ZbDJ+QXCga+nRhDXUCJGea+W6xW
PVn8jqTGio9+IM7LQGoqgiVqhvdTRUUa3hJym5yA7zsT3lqcYmRDrDCtmmn4VadH3TPFI9LJPLXF
kALuGQutpDR82yJCRmuXJTXwPHx9QDWL0ZS/L9mIY57muUZIBzuxw6ZDYMOoKt2oUE0eqZZQpxMC
ScdjOFi/nkBb6bEY8xbRTgC6h4wrEk3ptSsI2IYMJ7i7y/EnIsb85uPaYd8Z58QywXf3IAy4dE8n
52YVcQftp8y1Bf6AaRq0TQujIJEDE931KipwGgLk8ABQCCD0uezB12o11Wy+NAZV2MEoWylLxZ0S
3wRRQvcCO9zoqe+cuERsvKJSI0spYr5cgWrvKLrxpscVvrgMUejgucQZdbM+5zUkNo4DafOUOe7c
gri+bHmcBMg7+HGk60PI/MruGbnB2npVqQNmQ8Cr5GLAtJUcrTC/tyCqRB57zk2UxW5PBbvb1ApC
82CcVPgDzEDasySMu0LdNr4hTSGfMQCNyMkj1daIll6BU/5yCSDLMb8c8AseAOhyD+PR8c64PYQA
zAmDHw0Ujw9Cj95RzAcYJBE+wxlp4tcr9ZrALvWu7zO+PSSiEaYlcGsBx4mC0+evWgDX0gcr8NlD
nGU0vMUXdkLrxl1GNYerV9ftM5kYe+nIeCE+jD5F2xYUki8HMK9wcdBq2Wqw05Hky2G+MT5HgbDL
cYudywLgRXeF29GtOnu1Q14GwuiHfSbTjsboTM5VcwhfgqyHs1WtEYbuMpGzI4j9r2W0zeOqJ7oh
1SgNXf5JZiQjtc0GHlE9WRkB3HlkU8G5sOX6QURqbnVPkO6+zyk9r+ry1XjxcO89wmyADOvzBsj8
mJsrUpMBTU+7soihxlrDR/4S1RwVoBgoMUSa59rxyDqW7KG72ImPePl+SqZwnGeRqgLCjiD7WBtY
vpfh0crPB8O3uplVAoJJgQxLF+EmPc/IgJtnf2dp8pYv/Ej3KOGxuj+daSPxvG4IRMk12V0iBfJd
Gk1L6LzXLKr04szjkKHWI3ByNCDN9YPMhaxRbaNccOdxRspdvV7dvNu7hPQO2FdNwbt4exDOI2Kt
F1D+EcO8L5cNnYj2uJijNXHqzm746NYydO7/EuAXgSx/kQpPjEmBuWd8mUMyj6cALKRzvcPTdrOB
bfdkMtd8Wt1aATfrSKkQWftBnb+84sWUWGTXJGctiZzy21cRKmu76Wl6ICQvK7hAM2P/nJqBRTrD
RgtV+VodJlbLPel2a5So831cXNDqqmgRSgVotHAoVxdMlySx6cxLMbEZBl8rSb781UDcm9Rca7Of
IXgGf7TziGo0e3LwMzDbeP9J3Rh1vhEro9tfIlBtyjV5vjCS1MR2myFrFVsf3XheWanzk1ZH5HtS
vlv2WwuOe+OXjbos2xyfC/PNshTu9E3+y8TJERCylWqbNYSNxqWM3z8Gvm2cR48I8KljGvMWjzxE
yB800EKcuPf18jM3y3RbzdZw0Dsw5S8XcuMknd7LmLlZjyQt3iP+KsUtVAA6cA1Ro1KBXOo8CXDw
hQxWOr7wNfVDEZv+LYxzWTBPGCPgdLZxp5I+lqbSRWFkr5EP4HWK8+Y1LX71xlkOnfo6meoBjg5v
Ip8J0oe/NHslny0ujXjQVggjvOzCTJRpz415wQ8R3aIalnZPhFAiqCBTSEq44Y6AenEmIXYYcSBp
5qFbfSGv0YERvoEi3n4Zj88pZqqlNtVE8x7OR/W7vTbN2FoucU3p9nxIP/zdDWxUJuanyhK/9aqQ
MssB01WDRYIMQduzNi83SRX2rRTENB0PJ14l/l4iQjzquRnpwYbQMI2e78lfKRHxrioxHIkUOPWO
0/faS7BDYR4XZXRYEY7qVDHKCbeYaC+Rscguzve6uv5EKeorsKR2dvJVQ329TLmqmfhoCf1+mvFy
FmVgs9rbROPvB5sF8lnwZgmjDmCXKLc6kYP6HLlAobQaLO8IdhIkQIpUHwC8MqibfMeMw9YWb2Ez
bbq1foTuWEgE7vMBZbl9otdHcTC4F9g7ObJhoNYEBRkePQsVIrNDfqJF7jzLYU47uLrbPLCgqWA9
Nis7f2kA0U4bfXPP4gmsT8CZ3mE6Opn7bquOtr6l/njtWdmmP8hVhFTE1f8xTdsFw0dce4zra34X
BTGb4mCtJtG1eagt6v2d/0bfaNXRpayTYbX64NjivjHUmBG8fERk0CTPJfm7EabxjpnGlMfvz18w
BkicVihRIGyS6lwVDGyRGQJvZlg7r4wJwde2dWta/vjfxhfNMVBorobgzhvSRgbUHMZg76E7Z3aU
pM5Zc2n4W33W70gAFyYq4ikdeX4yQa8dNeLJGYUPbwSnKSXcp9cVX3zicZ29tR9fNdLjw8hNXnR+
dC06eEIjVq6psl9HRc41onr6aUK3kJKCXy8sC/M3i75HWC9lOpVkzIw6CeP2avUyv2fZqP3P2WwI
Sr1CbQ5xHiZzW6yZikm+M9TYS/YUWlj4ZU7BgWp5q/PshW+raCA45v6uwvhGUzZlNMzkfNNY1hDN
EokMdmPDmCCbebPvx+OUnL9cWiYV+0jeh25jW/aNtecI2Ze8U6yrmWQ+mTOFu211Ftc5BIexyGdF
pIblz9d3QxuvXVcwAutE74WKXxae1LGwDqznHH4PC3seKcR3JFi39UZ6P5rfWiYW7whpSREHlPQ9
BD3ZGuRw6ajQZd93Rl061SYihQIxwPG0UmObHDmsbqxKWDhNRvUK7Nc40RymqQ5YVOclUWGRJ3Aw
PLlPRwogp8PET8FjR+w/a9GmeO3h5SputHacVOnKFEHnF0wxb6yJgPaVkM/13XrdxT6GSfualKks
vFP83FExmsgKCfUtQtbeH17wTHPKTQ43/cCHV70Cq8Kxh5Zw6wd1QbOBHJkotS1c4kgmOPoXUOW/
tCr4nkTfgX6WMa4UKegTlb61KXTq2fHidpBqnxUoDuvFdCS+vr3KzoZEZldR0pZgVUSTUxq1vdmo
RJXNJY3YUDp6EARTkKbeWzR5dxnEEaGg/F9r9KOzvrL9D9Pcka3CJJcgnN1sT5NlTz3oGXomdXIp
TG92P0tBZ6Ldf/kEP1T2ca4rBFaSIjCJCh3YpTgYbKj0vBxbl92wD+FtQ7PhqHks0jeRopByo30W
C54tSNKdnmnweaIE1w370S27PXg2FgzTENPScxpuzq3HPLagVV3L8BNkH6yxzm1Q9h4pUpbjGEp7
mrF72Zy49n+eYLX8orvV9Dmf0edfDOUPUlfk3fIxqAv5B5NTLDl40FX/jiz8o0z0k3R8t8uoIbKM
y7P3A2qq3wHF9Hkj83XwiJUIOInyXJlfHbMfw7oVsIr6sWyPox3SHvMl0hQ+EINj/ZoPzFQvdfeG
eMh7ES/UMjK4sK9+hVs08KWZZA82125kn9MFzdcTvgB1VuU5xXtQAbH8rtUJ5pxFSXDUm3TCv2LL
/uPqM8gP+996WtsfBm9ezJGzrAYjgEKtVapYwtPHaTjNE9SFit7bWJpaDy03duALIQR7/zKcwnFT
g6mlmm8T74iq10zHvIYWarVDq98BD7+TTZW+Ln40EeDzMnnGtHhpigBleXZg6P8+LlzETgpxnifR
VAjMNGNqz/JFwZYoyAnZAMlchKW0iUkJTV+L0w3IZPDd9/CrykR1/Qm9MUIto9tv2au5F+YffxyQ
GYc4GIEfbUkgMMM6nDgVQlI9zNQI7nKZHpff1+2YNxrdfTmqEz4+1byfegbx8tT3kS3zdWb1vrYs
aN9K13ZlWX8gGPMgkzFwurdEbmZa0N4g6hop70gATi1V52q7Kzznob6v8YSQ5oGozEgDAEvLR9UM
HZlZAtlNgIw8F8iL4MjG6zxlFRxinynk4dmg1ZP/AgIchuf3qF6jghpz4X5CsBRvEXvRJC8GW+pT
Fwz/h6++3/Vcmw1VX0FWUmJETXRHiPQr+0L2ZOmR59yHxzveIFPbaXdFhZ41tadc8P0zs6wKKab/
jZ7HPbjxYM1eHPuGoYsDy9ayFzmqvBW19y9c70dyfon6cK6r41eHZSahuUrHUh1ylU6w9ZDhtQUu
xoT8gwtNZWARocm3pX8hS/ejFoJt2MdlqaOLtvDsW1obybQgzqBOXE/os2WaIokcAlspPTRX8H8W
aNjL4r6Lsgj4OWvmsh6Wddn2GqfhcBa3a09yrIv8UvhMw/st3IU48t41JR90pDf5fh1VVa8ETiqo
s0LdAXKnLhSTATqu6YBu5MlX+Ia/3TDcjuHTWAOxvvRuz8CsyRi2dDuCzyV4/gwqqYs+VztonLJz
1uZnGEESc5QVE12XlZCPLCbjLrEkI/o2ky0pJA+eeAhbLjawe/7dPSm77DA2Py4mCK/3tZsugM8K
J/l5NAfEqS+Ikg9yEtPcesyhFKtLG7ZYGyrHBP3r9zDvY6fXrWJ+cxj3cbY18GCGxSHEaOwaFMQF
i/Qwf/ZPDf3ZsOo9Qr/WH0gcH3NxQswdCVuN1FRiS07rxjcmFaBk4I/wogYAotzU6Hsg+R3ILyx7
6isASWRqajhqlgdAyB5i2P4kz50DQ82q3X5DSk9N+vhicmtDTz7Op28c/jXIqwgTAEIuXPcLgbTa
V5BlyUbpONFOpAPMZk/Gu80T7i0tCnbd+hugKJGq9WjdBHd8bh4k5aomXZyKhuIVn3Yzl/Z4xy5F
I7Bq+ERo54emS//p92QV/88g84zi9MEkWj5tf3xjZAuX8WdbmMTb9NwefSHzyfDW5E2te9O37zkv
EKdTHN/gL/qO/fMuN17uk3Vs9cNOxeFuHoPaPfLn9wQzwWt7fxOihfETquaq8a4ZIDxCwCzzCJL5
sqgCRjJbUiPHY27DkZUETTvol/eZfUIQGKV7noiAKipxKrnasDJG5pi+/QcJJSncWUcKLVf8Chmg
kmlFV38dLgYxs8XQLp4R6wQCCiS4BvdhRpwUn0fyaXuGHp7Rf7jIIeuVmd58XBTpJ2b2QItL/gmd
FGFEDIJXhgvmDTqpo/aS5CUJcIw5E5fGvQB1WbATUFksLDNaeloeO8lxu8o/patXKOe2AM1O2Kpn
vFOxxR4+Cb2Rxubdq/DEx1Q4Klh6lCc8SmokmPbZXBtCumd94h3ho32V498gaXINi2rT0JAOiti8
MKTK/auCWWFHqhDSXdhrTpWpaFrp2axVizMi9DShYTZk6GF0z6e5iW5j5VmAyd87ywwfI/9ONE73
ws4WVBmT3jTderF38ggfoUAnf38N9xRm2wb/iGDMoGAAgjReMf8xfqFKoAkoXSHfAVHGbaMmwng2
3+PL10B+BWA7dyribXq6TIpFM2BmVlwsvJDVJlGg1INJgUsJi+Im2/AgTXy48jkCXWtkfRv3QBVH
Gf0HeqhCS93yTX36oczXOO0z79D8g5Be8WZWoc/+JYoDQYagmdMkjDANADfHR4YGTYwvApnNRpqJ
I48Qwfsp2RZJghq15x4GnSYm4EBWSTbyVo9U2LQYaGLzyLnbW98910W6PlBYCdMYnHG7TFbagBGi
dQCTJgRw5vBHteMBUHxgkiuS4sYWjWr6j1GGU8Dv3p07oJR4ORjIjJC5bksJ1B+BHQTCVnP7BD2+
NFIrJ31qHChBbLMt9+jr0Q7wh5XwST9lwfaX0bZ2GZnNmyGeamGYwr1ZFcYddOX7RGfwcING9O0j
qHYbxjTtYwoWPGZibQKvLIgIS1rQeiCcLsfgbYVLb24pWRKUbQ0RgBx3gnZYpma3LEiSrY/gJlTb
jOUQPFRQgp27VSnfGkPLfGTqs82gsdiPR1A4hEnXBNbvVC1ztL5eWLo6so4tbz1FhANT3yYktasG
rSyENTUQ9gLQRny1SX76EwH4ytZep83RR0n2YQ6fEnZ0vMrWcrqXTIvGTw6s++8Xj89BOsijuLU4
5ohAFr/W//OnycU4nctKjT5p4eY3f60M1jlpKYfc4uzNwbD+7Zr8KJLt06Y+P+kDS86Ulkadgo5z
rvrOXiqU2DGQ04ezigxnoG39xpmrzZTh1+2Xtp1wL6nR4A7XFtk7mz7IAgdFkPHuj3OBDjGAmkmC
ua/elZpC/EaR/drBQkvHEFu+bwjKU6wu0S7PCJO8jiG6hXd4VIt7Dk6g7uImOXJ3ACZQtpm0Bt1O
rHJqW4Rr/P6Eo4gzcO6+7VpCNGzKp9RssJja9xlW/TSl26vp95OabTEsrk/A6HT9FYkNdfbewV16
TCGadHmN12/Pw95IF1T6bmB7zY33OqfklGrvbipOQSEkpf/LXWzojTOLhQ11rZIFXDnE6f1OJWl3
T+ZIKgUHiiZSgNK4sTgAmOEuyThpewhgWuVCv8UmiSkV8nkIqsr2yCACgjM+zyOA+9RsgatS7LK9
GsH053FCgnJHZjy3YKmPwiOczYwinlPzd9t0M9nrLtPPsCOswBKEs+WpYW/MaI4qwLtyAIFHYPLr
dq58pPrusapMzFnxF6/NEL7EzDoVdC9Wq0jTLz5pBN98YRdCPtEjzGkXxNATmd+/KRZXcjqvnX0P
IqEEzGj+TZb6xOCsQ+0lmxnljdO0pMzteYS5cJ31+pudeDob7htxfj+MgjFQts53WhMiSLS5HTEl
z7B8uBtVAu9ls0pkuzv2Jv5OuzyGUd6SjvbUFoEJbj7RpiMHrnay+x4uQ9YAKMP8Uf0bjVgwOL0X
BEu9NFMA5pr6zCkRbL0+WevuqcGiqcK13ChS6px3mSWoR5V4bn2Rvg1NbWG42WmJYQnabUcd5M0/
E5/5PoMwBV1ZSqLeeXT7o+57muN2LevN+/n73qL9u+DMYgW48/MQViD5q5zIS+7k8dPHZVlF5mdQ
QlSYkOaK7k2kz+TCZ0hbHsxwm8kVBxEm+J2ExBxVxPkZgxMslfpDzbuM1k+ZzqcAVmXcp4CitkgC
Z//LKZFnDjeJvwWtPt4ERdWKq557au1Pd5qKBccIgfJmRq3wTRUEVshNjPkW3v4cf5DE6bQt5iUi
trfCNZVtIASXvVewjT+5GSJOl4Nr4Swtvg3KSXG4QeJ7Eqtdjtls+ZljJT72GXCJKghNxsLnzU7J
u+GnoNJOo9Rug60JeXKWV35ViOk6Jq/RWC9sIEE/wYTVB3rz1Z90rdkQuwUrNYxKYBKoB4dTq/rf
bcQOiGnyrIlVv4lcr9/bq8Bzu9Da4IqTr2lY5yKw+ulMM1oQcLSDuieMr8rH4fSBBADR38rvHhmX
lF8lu5L+iWlpCm9j6+kvjZtjqfJD7fvh2ZnfU3pW1vReYwxoh1QrR9MPfG44F/Su8fgU+5p3jDZB
v7sOLuNFthBre7CnK52l98GB7AByVIW/s0eQZooPORnvPNLqc7RBE5ENya4HTSzRMtPJFxmlcBVK
DMiO3Vltt0phorvvUv3gj8OfF3F7gppmlzPFlorxZw2xh6tXFeCcY0lQ1V6xlw13iwRG5HAp17wg
BpAUQ05w60kXSdSdKfVEKO8ZBYGA/utYYeeIeO6CKOyOoE67x+HSL9bHMyWDYYIjM1cw9PML6xdv
elijf+iqcmKaXQpUleWgbrYAWBoZ27C7alLVa2ItEf2H2bGR9dF5xPvchzCV5K8fdjd4+ftDdghd
Uhs+Og917bnsVrxV45s1p4Hup+VF/rfXRGwCJzWLeyO/rymdGR2KP9Rh6H0gF5vxRq1n1gKiJcAU
/IipMaMSUBj15x4g88nQSwayLv/I14lAWiS3JBJ96H1CdiTvaNpLibg8FFRUBcu/Jg0qkHOaSodS
iccNQcHPMf8ZmjOhSSkNTD5Eb/73jOI1tRD1tp+86bHFnJgA+QpHKTDGY8ZxTE7CamboRwxL7/es
PdJhvlJqRlq4wR9Vrodn7jIhgJvyn8HEOGUf0cYju8xntkFlk3EuzeW+u8Mb3QzrMIqMGfVbH7PA
lc5Rj5p55y8eIOzqc1SK67SbeCm0oWAShmEOfoC9Y0BboJSNwjt48FhJ+NRIO40iSjQJjpwHCs7h
j62UDqEcMIa0Oj6+wAnlqm7zF9cQJ2mSuTtvk8Zx52NFyhS17vPDCqWX9cXpz1puGrXNn7D6hDRY
YJTApRgutMEFbkAxn56iSKIMBWKp6NOi2tzpFIVEWYBpefODaUVI1RcWxbY6WjcrDX4fITYDsnQS
IV/M6/nB+QrMiXaYREVhQBuOTux6kjJeu9Rb7LnDmzlG4byFG+wwROb6dYEt3LrdMz10VpQxAJZh
RCvqV5Vj4DgEG9au/rlArScTd6KHUCNPIdXQWfIsW4KnGmalVbF1Osxrw++F0CF+h3lWK8ydMHQd
PpgBCZ4SXtj6Wpn8DStspb6UrdmtGbdRyMmxjY5l20wteXDynxcdKDayJlKV2BjzZhQXJJZOZB63
xDoIUiWX+kLKASYqwfPbVoLCDrZQSx6Xhu1fSZDv+8S2uO7iLupjkadSu7RfXWemnrmdRdfri0ep
7v+hJALrse+hDcVEsMCJOJozRBJldqFa3F5YY+4cM5VFUw==
`protect end_protected
