`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 257168)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbe8d+E5z3uBYKjPzbXZZ58ehCdnrM
ttlYxY8AcSBhsTSehSyhLNgfK7syuyEtZqtqNG1ELm6lvbuHcUllU0M2P+jNt0AOC2Bh7SlDxSfP
d6AdCWybopdGcw7YEWDkdmvmBH1PXzDph9OJLdsHjJ6gu2Ti6mV+YBYYlwSlvh3UFF+Cg4l08F/I
jwgMzYVrgx26GF5EaibTYpDCEBu6rTUFZbO2oNN+v8463LBO3hO6RIHZ+pOkWTs0LuYpOJMdlLi7
qW+9lxwP7QvrrMyhfAIZ75klq5l0POIn0ff7Qtvbm6wBvoZ5cuJe0RLJAup3GGOhvfGWHtzSWTEe
BYXvbI2NrqR6sCsWban4fq0MDYEN3d5eP9sMhAR2163dfH9p7Z/T4pYD+Twb/LuviT91BhlNcIlk
iH5zp+IGoEYyT6RmI1roMi7M+usyU3J/RwT0HxVaAoRWqy6tptsMwmQiOmbwZXeeawKkneehGta9
o1r8fbZSjo36m24sMRSvzUVFoJO8vl6eK6VTan2KeJMOsL9NJT+AoulaqolNfh/X623XebMU0pgg
eSubkb5k3abh1xJKrJtyZsUaXU1dSn1aKF6N003Uspm9HUDOKQEB8tzj0xOKQAIVewfzVH/sCo6S
idVQhumot7daihAlBxEBSd7/Nlx9Pk2wnQKucScJ3Bzxkr4QTMXT2gNQj5G0mIk/l3B/5/GeiUdV
PY6duxVy/iFDFmz0/krkpdIzu+O8upGu1qihTGlfBvlrgrRzJBKZyXJPrzjW8fD38985YIVvfGMt
pd8Sb84/Hc50oDjHCj+n8DJlZbOWplxuNlJF2XMAMlsTY36kbQz8WqSkt2JSFEK4ukSthc2NOcO/
Xq1TWdl8aEdZ3yhSjIexwmLTTu6Jdai3xt15gB7FXTdw33appn3lzTuMFdx3Dmn7ewy/8l71OGQH
dN07T2/idCbzpuDB8giKdJj3c9gGgTx07zv0+XWaXTDswAKXf7AKE0OArisplqfTrloOJVkFSOJB
KaDSInqgSGdInApFr51bvwPppe0boUTjqzVMVfEgiH290lFz1gxtltsl9NheDMA8j2YxnisnzDUM
8eLGTurP9S8qlompm9Z/WCy/FInzZw+8VPusooM0RhjsszlZfwAZZzlfnzklSWiddJ/od9LCBQ7e
m/9ApEWVPTgXbmzyvpQk7U0Wawg8VRhGjP0zzRoEP3GgFH7KhCsCr/ws5BNEj2MQhtuDpqWKflE/
99G05rXAE3eNHfABOkFdrtj7aTfFnjS42PLnXBQfvkOElUL16UXZHSB3+yuCmr/xUQ3giYp5Hva9
ccKhHmngv8T9aLa0+kayGq/g3mvMyhja0OzRTbLsjSBlWnM2NpWifbU5rDJ+ZhQkwdP7GNjPxfww
Yp2ayDr/4oHvzWwFFKVdp2WI92dBF1PFd0KVCzlHbT32LhWwQrzJ+ForjPlrvhvtE3nBLx7xzAmE
6g+G7refhQ4tWTPviAlpgXJeQ+bfTGC6stgDFwychE5iyIEFO7GjupZ1zZT32ELSNXLlo78/91te
/ejcjyqDaOtCWuwfowb+yB0uJ1tzLtEu1P/vsNqXNHJlSx3mDs/gUn22GYz0AgrIQiK+MO3yUou1
K+gChs0U6Q6ZJFekhjkjWxdBwp/myRTky6w87MWki6WUDs+OuxLU9+PCKHBVW7dkfAA1oQmfaUUC
MyTYb1quNF26NLqPPdMqRHKkyb7AAtNM/w7PCJlvLX2eK+Q3CLf+ep8/mrmlknD9kUZ9Twf8PXDF
ltYDg9G3QGhyWUV9vxmEaA6IVxCpBeE8PVi9+gZagNigEml+end6Y834rcgYTbRG9eNod7GpsPhX
eHUW0XkHPTBuRXTHEgfgCIkamC4DVxlYFEkqC5s+mBPudL0O8KA6FQr+P/ql7ySqlpy7Zjqi/h2E
qzql6EVRaBcmygTkM29LQbtSeUSVKtcT9KZDAxanIRxExOfBF6pkDVQ7uynJs9IQP/wrMsAbMVBc
+EqkP7b/K9gM/yli1NIm9lg0OdHIgXK0VYc865At9nO97O9bJJ6Uj0RLLJIx7UsZJa/gofqUEIeS
r+ROya4O30OzWlS3dowKrVy0WJbss7X5Lfa0oeLZR/efwcWxuGX7O+53YKwIN3D+Ug97LbRA70Bt
h6uS6+OFBwQI9Zb05NZgU5fzrq6Refg094fsxyrkQE3EuqSecQEOUZrpQIUwxzpZrTNpmcSBBdQv
sKaxlT7JcYg728JIbN5oeFbxwZHnGUpJe9Lje0OA7VYOakT9tCmPs3pEQQJryE3ZyXcRau7o7yvt
9zNr6QmqBX1vNYVvs5X5ztia+w2GRYudyVWtOya88HQLMYAasu8ZaN2T940euyEIqv64L0TE3DWz
sHmFRGOShDpOMVNykzcAX4nigyL4u0WouiJYFz7VkAxopvQJyGCQUYIq4hcsmg9BZYcgoCdyB0yC
OVB2V1X0N5AOllOoXeHt+OhYzRGWZH6jG3qci4Uzn6be7vUrMEY6nBLZvE6Oyg6Y4ieLBYM6yBEL
nap3Fip4+0nGOH/VLaJklbANuiyZjnDD8w35nOspVEMSvvwafbbr+7BDNwmhG6h3SjMaIEqXYnff
xdeiFIy7hg73fRXGrk/eM4Mv18EY0jz7kh5ODfmPW+IIOIQyiL4QJn1i8MFEMDmF/1hBvxnVWbLi
a7dKxkyb8+S338rRlCDAAhg+ZZ7nljPM5YK0kG9RVsa/nep6G9M+GY4i0WjfrfL0gkFS/HDVPXZb
yBoWXXH2CrTkTprSn3OEwXX3k55hpGuxREIrrSjNiwm1ijmUdlasjzSqEnAIJLlL3O84CoWQ8J3m
taBFlLx9JGQaTtQeB7ha5q6wyvhaFiVx5prDdjUXoIIyjSBYOdUPiTMgoL8X0u1BmURC0WquAl2Q
KcGR3QVjiCg0orf9oNvgTWBNWxUOITKUKvFiAEdTJJMycsiwZbmge1URm25LORL7P5/1kYcq676d
RFOshd8Y9kSotUxkd3l/ljeD/RhjfkYy6IkNe4OD/IHwT9+lvsOJTnIL4Iuqlz2E/FWmHBFd6T38
rGwKFE1r24gs+FKAaj6XZ9W07rWLUmpi+SG6d4XHfrJ+AVZRdD9HYPzS7TgUjR05wgImrC6XSFgP
hBLDut3s8c/pPXev92nCMAwuwZWNcY1PmpmBbJOoK3e1U/lmd4ujWmVdtIOGqU7MonnFGhcYCSKc
W5K+GdI1ZLciMGFNbVXZCZ+a03qW31WfA5i94V0zIUbO0tH00kv12BXf2bzcYo15mLaL0XP1qXjY
36jsnaq7MBO8ayTmCgCUsHkqNEdLLghJFZalBu10mpbHsYF3PVkHUj3/Kf7+AzjZOsroe0Pp3oxG
VlaGVoQ/pVrkeGbOaclASyJqg6O7w0mCIrouX4qUFekYWELvm0sXw8wMqeliqBBxXWcbp9C44MD4
YFmaW5jfQExtGyWPFnr2oI87ukYo9ksGW8egh4zycSSpSyDL3fkCYDO12pt1pMxABRHqCgGjqw7k
axR6c429DslYTEDuQiYdrDcDaZbetb8H7k1qq8wuEQioaHdyUJi/n/UUwHuEjxDNroRv9+Lm6MsU
n2yzYKsBQomrFJwsvBkc8sXDJxTA9cdYthMr6MZyJmafXY/fiunQOcyf4gQzBAUQJD3PWnm4FqIU
4uc7HPua+HKYj8baQL/Swac9eDSy3F8oPqqZq4m9v/CBv/lzPXvLlKcXcHD2MSznnEYxAj7AdDKK
4Hq8d2oHOdW4YAoGRGuK4Da8dB8ml038vuOtToWKeJ9LrmDrVJhMGVVK2/LfZWr/6NPQSTRFW/sE
g2K51KTiqanu0Art4O3gqTz5nm7YPprMU8bz3/9niuCvv0yIhl72Knezsrn6z/ryca7YNo64lFWz
P654JqNJk1ngwn+xcvjupLMk2YAnf4hVGIvxbI0xEeO+rPZkhN2kcIsU+KYF6I+nIiQKQk+3yh6N
jdZAKx6okmm5+FqwVRst3VC8aDuFnVffNEmjTUgSHk/h2JtVaOZs0wfR0+YqQu79ZbClQnIv2L4b
bkjIv+N/KC8oT+bohsRW6g5igngOWRT8+ut7DnVI60wKSmw0IAwDLDceFk0L1XrA643RGVCF7PRV
5hJDjw86rFErBe6BPe951tIayyAhc8Nw2gj5TPOVQX/ZDmASlgJTPIvWIhx+SJy1S6wUYrdW5jCG
XsWqWdkS48eNeDHK7MW8SnOcqQSKd170eBujrxFE/XHyA1sBxi2yEJwJaxVjsImAKTzyMKjOE4j0
ktj9pkkxGcoAHMKRMjHcZnpTLrpjCLbhuWjh3GDAda96Rs2nbhFLNkQdWXCpRkl42PANcF8c0K0n
Y9+GuV0+57QwgxaGksqWP0yURSsQULk5fDpMq8z/tGGyhOqaOaS0Ftr2uO6Ps5pRze8Zsg4GSMGH
ztvNKDiEd/et0VCZI9Tiks852oGkyDCCV7TotqzJybiynw+Ty1a1T0WwVKGD4cNfhJ9KcUQBgmCt
JB9+qPV2NRfZR+gltVYJr+lEA3/m2LN/SffWFakuxC1Hb7cAil8ivC89+V1jd2WSdS3pQK190COn
q8H2hugCCgzWB2HoUfzMG8Iy6R/oWNQT7b5wvevHOy3d56hQOshSjczIbRW4acQYkB4dwLFmsyu5
CAASafZO48NVqicqCZIE2vSAfHwNIh4HEm5V3SmX1kzfgLnKdcPN71D/UI/8y9AxyziS3GdzhKfB
WjPSZB5HkTx4qvfDV0EwnZdYuTWnHb+KaLrm5VOv0ScGIKvNGgywDo0pXHZWn6Y3xl2Wm6kq8Q9S
5jJ5dTwbjPNDFHClnzhNhbf/Zo0IpxrVqbR1uxcF0qzSvqUY2wkr9e6gbbpf1L25jqA029KKR9G6
0+xWbKZxlQ0NRiUnEt390Qg4r/N+IHX+3nHISEiqj1UZYavoiPI1X3a281IhBBkeWmX63ByH1EnW
sf2LzHM5A7OTaxIrjJQyP4AorT3xLPfuHonUsArTmIc8N+7CgAHkfzQsopGcpX1At73ej1Fo+aVt
CDF9MyEqyuGRHmU25cCy9D0r8Tmz/nyN7IFUVDFeDzPFXpZ3sFkY7T/sb7gF9mIXI9d3BfgmIxLv
f7hz0oaEVEdVaNibm9HxsojTg5vaUDVqIRatJFJ7dGH/iEL2ceZoKhSYmXlINtQeA7dqGBnO18kq
yc2vuyYdpUf19IaMdpQSgMDmRNHqDywtbdIjXGcC71AxuIEKMBdJj2qv3Nafcskf6WLIIimQr6wu
p8KXh7wGntAN8/uynlRukWuzaYWh2zpz/1QF1f00VbEgtlcSOHEZbNzVYkJUAIWexLRxsyVndTxZ
6+Dr4d1KcG81+F/94UawTMkiH/IdlZKg4E4ZMtImUkjTfAP6VZUdbZ6TIoO8COLlhgoaxIPZp6Ae
XS7Op2w2Gr8BkMEizseju9CTbwX6wxgP7mv9/O/rPjnDlgX2VyGAmMEpM+C50dlVU19mRkLp8FCV
V96NIjn2xagApDVq5L8mxrpuWF21yefp2u+9vPJoouS72Fd5xdh4ihdkMBb7KzadeFHLT5jO0XW/
gLiyPpU0kW4nsn2eq2ULeXhcq6L4NdDR9w/EpCtDP5crEPx4v/VaVzFDm/0KctqcKraHfEgTI1YF
qdpHV11l6Bo5kXpSnE3RbYQ40ejaRgytUXNreVzGsGBnd9yQIy2prX+TxM1whBj2uwH9zGA1ABZm
LppV7U8uM1Y4WALIsSkuwU3ZiZ2weH+QLMETfs7C+fcXewlRl72G+CWa1BI3PsiTJ1TUZH1GX9j3
L/QgprnVDAde2jpVXPug2Gegiqc76uLboxzYNy8sQVr6oHFbJSQZ6ck7r1Sg0AyZDsfYXfRUfNEG
znLUlz8AYnrj7Zi7qb3Jp1B18/moOF9iftRid6eQJzy309/UdyVHFS76XH3WKWFdgbpXOL8zAG7R
Vw4siyzmCeN2QavmoWAvQIZI3xyeunsEQzwUAsoew9jqJFxzFFSNdzz1PPMjGc3KxyJB7kjz6Z0/
MOz4I5yfRY77kANPNw87t3c2nNBOTZH1dKxaVYnURiNCTDSTUm917ug0ENwicSeH0ulLFJ6o9eWa
XhcwS0BbbDY8Xxqf6cSseKTYaSsM5rW9gAOrTVtNwzcKo5vitwC7rg11tucH8kPxDqZ3sdMgL5vW
QbRLOyYOItdftlecDjm3EIbtHTRllXrgHIwSu2nY9IqbTEngiJmzlYqD4maGec892AG2punxR94x
Vc4ITQRdmTELlGV3MkgpBhsqS78Hi/MDL641Uzo9xPMQYL48p7pC5jxqY5sSII7TJIctvW+4DBJ4
jXZei5dDxK2x5eauzToH6WN2Zguux2zZOQkS2pOfAEVMZ24l0CwwmyNOms/aUB2qa64EFo28B4ot
GDDAUsa9vlN2IUDrwUjXVBK+UHxDhutnBt1qENrBPDlNjORUnC7Q2WpS3IKWYtlgZ8ADAnjuutmI
34fUgL9BQ55KGtPvRR+YYHNTpD5AqF0XywNHZKsf980mqn3WfKKQStOZP5CwrK3IYHorbd6hDQpG
RSY4LMAfvkCKM/BkTPwfwxRU95mfnMXpheRuCxzyIMfgDorFPz1WebLGQVzUDaPgrtTlGHBENMxY
iNjTOjH8Bt1wGRAq6RSQAbwbUQmN6tRK1yG2s8uRZ2Cp0TlTvcOyFwThU6JnbIACqMO0t0U2r10z
WTY9QBfEGZ0TfufTWTAvfSF9aBUZVMnRPczaAG026+k00Mo3VkMqJTKRj0lBqfBaqVRGmquG95z0
F8Wtcd8aNEK5RD4CIHadxNjUpQSX9QBV/w2vvWROcRzlLbYGx6o3TYsPMd4SGI7UPkahVP5/CnOY
/6MlKV+3Oe8rERAhyNvjQu9Lj2j12dfPG4wExL2gSVYgS+UBOEc1lWcdsBrmgRrPhSeJecYChEof
jiX+Y/y+l5MEEjqiBQ0qxxnAkqgIZEAJjBLyGgAfW8m3CQgcdW9UzAxs//ZvH11dvDLbYjjMoN+/
5vOSzGBKugkB0OmwYTGW2fbw7gpnvZ9fvQkadPSekEl/9idVBBE3DKUWARUkG5vxPmnE4Dv1jj/f
3NCY/7VriTu1TzQgboNKn8N9Nqe+g/9YRIEq73onhpvfLWOchlpwHWuaqVuHC4vokEQBwHFRT6hu
eMX2nmaaKImqHdE21PkPzy43xZfAqoh7WWilfqmU5f1rDfPWwSnmid+rziobye8Jx7bprMh46mQT
KLC2bQ7ROT9mVmTbKxaf2GIs3WmGCXkvXz4chpJMNvb81yXyAKxpiYkUfcouZNwpPWw9r8/CDuSk
luhsjTFZI2XbJcx7TL1ETu2zrXUOAiRdUS3aSnxxKcqnQCXV/Gp8YACQvxaRGlQudamEdIbtzllu
Kdnt+DBleOv93YdNtmawSbKONhvTPNao28OOmPMiNM3i7PM3ur5hUN8WKp2AMMmpQQGtJveyf9pr
UeXL/iV6ZNdx55pGpf5CYEOEsAX4vnSIFL6kWNlYxwHYkHgf/rNBN2hqS7DCARougZiv0U1isLdf
LqU+qxUrtxob64wpGUgXRX7WgVhdaGST37K8KQuG5kk9mPj4G4VndVqC8yXqcu4trNwmGpDZhiaa
pxkuTmeYax5vU/LMYPKI4SNVDYbf1uFzIeZuhvegJHepFzpVPI1UO24B0wZ13MOHVo5D7+yaka2q
9jQhD29Z6L/we/SiHgFmPWEOcaAlOwQeHLIdRnrvnpgym9p15dRj2fuRd+TSizKsdso2wviogWBM
NeBNdrznlry6EkTm+oVJzJHK2eA47nqCBcesZ0ecxmcXOhoiSuTzDCQcFTVg4wIzMaBDeFBr75Gw
WVs7xUG5m+ebygCHHco2cEHild393tLviL4sJchlHbwAM8g5BAMANxTRw8b/vvC8Emaf0WvKePVm
kNpavaFxB0KVhSoeIp9Hr+YtRRmK4kCrcdbjiepm9WLoNQeSFv9AnV7EeuVi9YBDSy8o6Nbp/vHf
jV++Rmvji5uDGNiNdMNfPrgMYN/Gft6Ie3QRIxV9ZdDADV2kIGXVNZa5GAgEK/lWrRpsnV4tvAUf
O8iIQepva/8hJAla7/4HII2/BAv4qiNK9gTeCcWs58tJoqO591xD0JT7MLv0VESd8r5TqtocVhId
hxdLNPuNTCY7yLL+R3sUGQkVm5LkppV6TPj9+gL8un5amt+PyVRcjKn/Ot97jzhtjtQi8qPxeezf
Zf9Uh9vV7OdJHBVKMMr1+8ewRfvAi3lTad6GgP5pX73hCb1+tKdZqoZgdaWdJ8v1A4OCPS7+ws+X
ota39hHiXTN4ewKxPRzY8YCdQB7sT0na4pp3AENemYbtWut04kSSF5Y8VaszQTABYy9Ff+brbt3g
Bx1uY/lD+/yFLsFz4ZTzmHqMmR86bjOoaR3sZOp005Sr79MWALkaUf4Md/XujhlEMKR5lFBY/XtB
Bdkzbugqbi8QYsfzk4cr3W3rAO7n91mB3LJJyGkH5OfWz1ftn7rlexXDp5q6B/sxk+YNkCs9cx/I
68H8xhjshNzADI7GaOlRcFDyfMhcDs9dK6R0cP3jAqVNdtVE+QimhGom07V+OAEO/2pVxxx0wM9Q
LXYYZPxJxIXWMMtupnGfIwiFptIcYkHS/c0b2CWFkuhCjnI4MLfzzARWf0vuWFuIjLHDiYmWy2Lo
tDKXK/TTE6ij6JoWgUEDpr8Qunww8sHDZusPKyO1l+ve1K1svp318bbtV8dhR6NxxpAw2ZGZLAmY
nlgUXh0O4vDwb75yfVJpc0gwUJjhNU5zRSIQcGsG0g8bEQqOg4l/NfTEsg3d0iPxTcwXoVOT7WmW
gj8ux8ZiUHt+xNPiEdzJsIt+muWoSiCAyNm5+1rBMOU+4eZRyXruiiJGOXLG0mYu5dRLDrPUzDr+
4Orebg7Ui/E9rDmoMbv5if/UYSyTADqwwEI2R+zox4AKUux+SZOl6CErsE5ucy9llGBU5+zXxxyY
t7ulL/U1/x5xXbCc1btPnuobZEKrYAPcLclXUkzYbqms4EMsvdZa/uo2uy8g8D2ejImCAvqa4gJL
i/krO6lPrItrEx828DKqzOt2HpZtlkk2eOJtKuZ4kf+wbcCjhj5K+6SIFpWGVXs2gZjkZdqdk4jT
3pUnk7wkFg9Nqgj+4jrtmjtxH+wYRsqJfpPemC3OYcdmX5J+AKOdoeVE2JXSjND11fcUUw2mUhmH
wHCSbuSf0OaJNa0sXZhMPZsLJ50FCiueB7ftzgHw6+Ix/2PNzpxAhgGlKjk9Cdsyf+J0yBgaC2ui
Mb92wTDBDUvGPbpkWJeHlv4HJiD3GZ2N/f3an33ZuX4Hol35Xbc+ftI7ODSHir8gTNPcIPyDO2H8
Jeq+Gq5rOAOPLEhzivbguhhswOQ3QuQYzpMy86RswwFqni6WRWuGifZao2uSG7oke7J5Xz8a+Ro3
yQbSOC/MQBvJiaXMZPgy5LvnCh/sSwqs/0qyuqA2adZtvX8bMOZl2YT/0fPfQeaAiYUXIhPnnY7A
zqaTCsSr9+1c7SxOaQm1Yc/nbWLhs1HCWHGlhvUOuZ551XVLwodfMNM+gqYLy80iJ65Yl2X9+/jO
AEzVhOQWAj4bxN8iV89ACtU6E9UZAPhGEZbneLzyZLJHvBmo5hl1lpdvtChsp3MyihF8qPvT4bYF
LNt0o4ar8BdWzScmjDNP4USoKReMGjeNTwhq/cfkXwAwp40G6ResQvC6uKG7pc4muzXirIixJhw/
bdpbF7ySKsifu+3BjsylFMJrDTh10GVyko4sJ402ROUryppgbBB0FwOtPM7w5OsPxsLR78+P++8y
100Jtb6ctVhaMm7KUUl/aEfC4sNb0q4f4dZErPvbzAdk/tlzYi0hT/tHJDU1TUiG9wAoXjmYsmGX
FOihGA10csNEKlkeFqcAER7i0z6fOsp6Dehj2lIGahDgG7dVVf1wKILU2fASv9c5GpGGV7hAcZ0r
t+YIHKm1pw15iUQy8NFglKzE5ryMrncm8lVHHUhm3fAYD6Use7xEmJMS5ZHbUw+AF+34LAUmqW8E
1ECy3e41eFTYzXkPkZ4BlWqYm0UoWOikDP7L5l6IYBVeg1/HRiTmt6jIWKFBRa9sGODbHVhQ8H3n
SfMRlDrj3t345EBQhZq695kKLlsHw8tedEQRe3a6miaTjJfcs+7VglF+nECmZ0qn4GaZlWiVGMFO
Tfn3RIgMlluGilXKa4XC+lQPSuCvCARFmtQeg2kwkQYeHWkGk6kgvPNzASQszSym4Vs4AIB9XEOF
IX1Cwy88dyNGcGu8hfxdVwZ44n/paFh8T0SPermETbPXG0uDUM9BX4fVHXiqkIP1cnTz8AU7vsEU
3/XtkRX9TKa5MnXII8boTzkGCYCw6Jxfwqe4u5AOZE7m00GMA0u+LIfGqHpZwCMtd/aHfixv2n73
0h8yVjOTKjoI7hIdMVvNS/m5dI25VrQJdilge/4lXekkjgkItqawGatptqJHWrucL2ut6+U88a8F
HUwoOoYZCHwoeX0Hhm4m+Eaoa5PIdHU3fq5gUUZfmUlGtDeunFd2MEhIDjdoFCPe/1TuzGGEMKk8
mPv/gUH2Bq7dhKGDCsmHXSp509jKOOVa6WtTjuLwas49zUloBNKDc6d/QiC/ztddkLqgRvlQThFY
Ef4238v3O/3M/3rnuqGzlTov/D4GmtPvG3F9S11wq2A6RHCHPihh1qMYNiC0nCBwlHxB4OjagZFk
ouCsbmX1OFjw/JhojYQg20oyd3kHcD5htyMtrWY+M0ff9FXLOMq9+5y8WdKgb2Zebq0A96WPu6WA
p8lEJKYZAhbh0OqnMhdMKFl/vASUBfZMDH173H5NDuAhv4a6phUTJFZdP/EY6iaQBqdQ9+3ILh3W
06bBpNjCAtcfMB7CSBREU9uESLRg6+gfeldEm9T9Y1r6vj6UlZo7BmyLv9RaOYNrazTvt7zfwy67
NqBxOcJPF3OpG85gN7u6UH5QOdaL3Yv2GsNXHCGh9w1gGZhEsBSqUAue8LUF6MZGO5hSCb4/dEqV
GG8wQvLcBeZxPqBNGkCqUkZVUr8Z+L8p5MQj5dY/xdt6Pr1nUtVF4Pb8m3uIh7jys2vkbyXo9TCA
zJsfWOyoqETMpHMVa/tf06qoF51x4cyReJtuwlW92f/8HrLd60yiN/C22A8gGwy1RCpebZy5mmIq
PmMLfwslFDjca8JwOG3XS8c3CWS1/dfNoANMFwn68uJHmKWGIR+Lf5B8+NrRL+UuAaZUTJToGAL8
gv8Tkzjog0yKMdb2a0sHCMmSjcv6AOVjjlKeRMhmoOnPJ5HkE+iuIcy23l3spQ+FI1u5hLjK3DNg
TuE659sKE2xtBKDKvUOLUkm1WE72QY33jCQm4y7v6+RRxb88uHcmVwXi3mxID44ehiASIc3tV0xx
hdQglYvJxVTqehXctYsydmvYFEyOojh8gaSS0uAAWD0mD152KQ8rckLubJLDdrBp2yJigyzhSDBn
it8kuw0rGHMuCV3JTBhCEle2YUoVZ6iSHI8Ku48oGwNczHvO/LFz/f5wyllhjlTSm9J6YKXWUIjq
pmhfX6Wol8KMH3Ff9XoAppjx9LnFZ5OQeRZHqwuC4nOCNZ4qMhXaFDCUH0IkQg7Cvsc9aFrrhfx2
SMlxsxXTMxge/7VKbn1CADtilhkNE1H/TMIZWD6sYTES5I9xa6hN7diQ24mOhGkD2EdM3DgsmlFN
wkd8tuE9Vlsxrvw/5qOi3+4n2wUAdpBcyxTBQ2pVtLh3qsJoF9XtqhIRBsTKhSEH0K+TQz0YtB+S
E526OMPCRB7DVJkTT95wuE7M8JtlZvW/PGeTjXs756Fi0x7OvKLlMNaX1b9H8l+4HK6j/pZuVG0Z
/7+5vnut9GTSce022wrhZ+QyUDd+Alld4qQXYxAfkTOg/rpQ9jiuLXdY7tGY3ro9H1fF3lRj40g4
l5oH/MJFS8vIgt4PSi3odFA3HFNg7pVVTuV7CfHnTvYixjlCiFI2zNwODjRxfhysflgmODzcOsyz
VwE+WSiKeY54JP64BHKanvhkyGqrQ4+4w97BbG8C/iRPegvPOrVHptNTH59fGVWh/k/XGo4GFCM8
4BwWttVLkaqEzkdNvtxKk810mFExuzuHZq+ylbBULJMepdQl7REbp9VPn9CZgJxfMvcZYSw9bh2q
kSJYaSaKAUEChC2Er05YYhU0mj9SoR1n+7rpX0VwgpvlJK8C5cwoHN+hr5uwgMFZBmPEXGXXV/8m
RWGrZUP3rKNqNUeja3uwD0KTMvuSgaEFQ3IRyspj/t0dqMt+Z06MBdlT3+OmQVWzhhrRYdgGVBgJ
KpJct8mX8q3qZ4KK7VCJMoekqd/KfE0J00maZIzyYYVB0NZpBDOVl6l+K7rCk8YxnA+sdt+I26LU
OHAdGbtFcu2LtG6Kn1CsW5lXarJje/whjjXCKW6FAcmnRpEuHXqDaGQcp8aoN6YHSat76W9hpaG5
cROI2fLvDb9e4Fp2sdAc756ZxmLdtzzUx+xNhi4zDhogBXj4yJ3END6gAZZB8bhQYg6iADnO83tn
gB8LeMeHam3ltUcCsfEayJsyJQLGE4qdNExm4l1td98hUgaUS4U6LlgCoatHFY/gO/VLQJTC+Npv
4XE5aAouIf3lFOYxcgxJpG6husTRVGbba22Ptb7l6EqPBus0IGmytKVB2BpoluN1IMasZHq2iEBR
TbZcoU+SDh/iiy6kjo0VSXYZqpnSpZT5XXYmjFq87H8Nh1JVuLcPDzzmFqDLa7z5QmCWbvow+hRz
3cvGtpSx8zLnftYBS4zoVQAs+X9zgFQ+mM4g2I83dKomkY/67zYu4cI6nmgtWdpXynV0xn63hNAt
KnsTuqcs19PGjlDs0kDAzVtvHEkPh3pzsAzD2T0hybqHBiAJoe+c2tsjQrubqkEZHnT2IaGCCKkX
hH3yLW1RPClosmKnRrGhKYucRBLTHZPVFOT0Wk3DFjQDWFFga+HEJpUzi2lahjMnp7r0atp/s8BB
IeU/t8pkgXzNpXVmqTa3GejUlwjIkzNevk1LZPXrkFGT8hQm/DjUMO/RsF2M5os6pUgx7b6RgwUi
teJeBY3W2OwOw2APZhuWFtGSHMVKvz/pRaFCUrrJlpAmb0i6onJr1pMDcI9cCmGkVEUFcN61ivxo
DKuqQKpnFAzEBVT01j0yNUDxeIQsoGz9umn9DE0BGbrMwgpclfeDq7IRydWuc5i3yhJg/QOgDNMv
FnNjKINRbw9hIAXIYevTmwQCxAzielWrfFZYGOPKZEsyihSBBeydjWvYVDtFp/vbsr00tJ31/Tza
jjp2pBMAjWpokXWKKdgNYNSE2o1/ejHWh8Vgg9KC0nvrCAyjr+oGVPsSvs9YyzqSJUFag43gIzSs
N1mwyvlJjsoxB0qk07Y77v/hO2RBYQkmiZ2WuPXUVGrc4uLn0QTnpv5Qx+iyq1NJrkEd4QrtupET
53wwLqVjTxo0A2h0a/nOMopI2mhgGhlsZiusLQC46D4lf+YWdTfWpKwUgTG8E1Pz7BoCDB6pzCCC
EZNqOBLeA3FGUfVhDV8xYyoZcCYg1UG29ivsEJQLNcjPgIXXEUdxr7hPG1NcSyumdUA76PY2xxtd
ZZhUck2zvkDLYBWqqkLaZoVk2pUuWgdDwhQH2PsCR9CPpwN8fkJKW7j16/s7EHVC+M43LIEHi7ot
+Ozd6GBuShWVv6kTC4DICpXeMB8ml0q3fSCcMFsk1aiVBrVfL8fKcAsnRbQNjipZrhrVAwQzBQyA
1oMjlJZPyRLvolz3mvrH81Qil0RI0QIBa2PHRPbojCV1Fadpc1D34bhizYjejHxcblo+gQ7AQuFh
44P4b6Nz72Jsn+mjAXei64fVhXBxzzgLaRgNzaG2dGN2ijC8wpgiW/aCPP988dpUMOXIOCFZnqyv
qm9JFqUbUB4Xsed78JYazKK/6fSMp2y32pnaV13vvYKkWLqSzLNlLkcr2yPbEb5avZ4CIiEF42+W
RKMEM2VkNzM+SKKjPRMHbg7/pvexaLD/di7aKaYvb8R7yCp5Pm0QDb0/vTJhNT2wLht+8CzdpPRZ
E55n60p8FnWmZ0RW2sngWyu0xRvyKHms8CaUWkwt6aPP/wndJgtclDhU3Ussl3rWgWpxEByV7+xc
Ohnu0Kt4RssK8qyOhv0aSMmdFDfWmoibHaS1FcVM9/Sgl2VN5mifnxd2+J2vgcKgXe5Ga13xSbOK
AG4Rr/D7TCg/e3+H1LbuZnGrKaVnDG8sQBflzVFqkACtq2wuTsPIWnfkS/BzbXIWWt4EwKAfoWqa
Xhkf66pHijqRX1p4M9XLhVWz37GrRuo0+zsTAr9hS5I6WEARgL7RqYFSYqxUkIZYs+PPgZoNfva4
NIsJM9+Bg8FmKynF86RT1WcuKtCEnHUkyke3QwX6oVHmb81mXbvZKPc32f8fIE6zuHgdqLiU+XTL
wzlCWezCU2ehJqCjq83MjIKTdDFVJOLVnNP4Io5VS+Re7KXgZEbPcmJcXRLERWAMnphIBdRl3OGS
xh4DbsvPD8QLtKL1QNeyRN7dD5sVBaWhDopU7y6JcXEsF8mpY9q9Qc2WyFI7N/DPXWSQ8N/QkugQ
bfqSbiEwHpxU0gNll3IJnYtnAPgz3EbUZMCveXwm0iVw43kUanAGKR89mqZPchvatp49+ZaF5DDj
n+wVhFb3YFUt/UfRGHOByVsof0UgIZDXjtap7Mjpw8TJeXthz5PX5vDIu7VPk5VxEaRgwRm5fr7v
ZY6wAUEuEDHJyies0O0EGY7LvNXKpLlipqDs4b/Q4hVuXA7KlhX61mfxAxHaVPMINcprxydaVzTx
4o9ucUUYWjt+v8Hq39UOdvx8PXTAVGENfQtgOvWClmuPefYQ+ZFEs6PyDbFncSdpvHvi3T4+UksY
XbBzX7yb1LcL/I49+Z2Z6ivWODkTYflnFiDDYGfL7/0vDYF+dk57twQK3utAKN4zgJ7okjohSQ5Q
xwzpj9GK98RLG/jV9eitalCJUZW98/4UzTSubFqoXGtMn4vF3GrHQ8r1ZYCfqn5wMJVC2ZamsHla
L2euwyDNVS4W7u9lHhVpSf36ZdjHkC4In2i/1sIBN+sO2TQ6ShFKX+jn7YFvOWEMEaxdqdCPPqDB
NCY0y3A/3+jkFnS7GUrbxKeSue3YLXuc/GR2qQQY9YZYgcZGPBU0q4rf+3ZskouryDwDFkmxdA/w
SQbSd+pvYFlPWLVqCwPHS9L+DhlwdvHQrI+JxAv0pJlE2QD/NWk0yc7y5AIT4HFf9HOX+3o1QPno
8CvyNQEAyuxUOdODaGj8G83DYWWpX1oQkbPYY9L2vLMm2Y1IQmwOMci8E+rLKrLDqReCrRh+g8Vj
jZdNzOTmyCo5KaUDAFcleGq21s8ZBVhuyzvgUTgIgdf8K8ZHxYF289PG8hztLcw/s9eLzO/wmibN
3RtL9LSDi+zEkp5GU/qrHUQ6WbDgYuTalko4mw++UK75zp8z9qu7Ei+vAyxYd2hxBzMX8cFTuT93
SEThKTgW8sZLjWl1S6Db+3rMcT0ddNPh4zFB8a+dfLxM5y0N81yxumrQE0VPZhX8M8+comyF7BIe
JeUplF++ILPV/HeBjpSvhVsslLgl6JUXGs1cVHC7kg8HNRToHRobWJ4xaMGQclhhSCwmCTIq+mZ6
bdWtUmyEeX6djkZ6wdv4VnQg60ZQcB2cCRWfwxiUiofQU8263f+lbpZw4oGSxJrHgGanHLYNEOC2
rLGFvfEyrJ1Wws3Amv5XSivtrL0nfTHMbiUcBYW17XnRqyoBJZ+4z2X23ftzfyARfsc7vKmn0zw9
wgtdxzM+nwjBt4gNYT8OUUTALk2trIrAuW+HQiEXE544OLBAGZ41K0pyHGmG+sK+ZWroHl48oN28
iQ4uKA9udYCygWHRe0NTYddiNsvuXG06n/PX0G9MuvC5CfLEjY6HnDUfPggQqy04iTLtpzLd8Ngl
ffSEFjtlPzumno1vrW+FObtXP/SOlqrcKds/o+yrEp0yPxaUm0gBBep+ECM5hqzNvQI5tdyGdIZF
E1r25Oi3sMJkDk7BQBLyGvoVqQnVdX1blVHKMGf5b3nJIJocHlXCwum9+4rr5ZIFN9mTash5Zx4w
llxTXHsu/kVXoeQV+Qh5QHEQ6gwWe8ilPuIvSaaIgTn3/AtpdA3eMaCLNtl95iyCmBxBg5PT3WKM
3IwWRNIo9n03n7WoaCb5r4mJiXfNuL3iWVQ43yGpgzGwFCj6SRh6//r9pmecEGDM4LbK94ZiyduW
W16RG6hwAQCxbry+3ryfvLK0pvQXJ3Sz4pa6KuOoWsHmVgPGLn5zpCpXpN3gvvgEFQzXICOg8dVy
VngPT6CbAWKMQuVBcaLc+pEP/dYKGjiydTJzSn7ziP7CoT47A7s5dTlVscGaClrriQzfjHsK1BTv
vv1CN7RHaNJPhyWCatRJCNnINKkb4blrRUwOoa6nG8dS2gDj3yB9bXNtNWw2zDSO09pGqCNaQW6u
hQEnmvYTEaSV6Rh7o5ENFU1rjjsW8YkKplMNlx2rJjDrJ+so0TjAcEymAYzQgQRA1lQuZmQmoBTr
YOYENllKTLJp9hOgr9bQxWmOoFQjpCoFowewqgUvorHee5FUh2rhab19nEwFGDCZQ8lVEdzSEeyA
xnoHsYAR1THja2lCn5R7NXpEUcfbcL8QPTuKUOeXCxBlIKgfXGiBs8TFWyVkNwtQhCu29uwPdv0W
6XFR8s0ZDZuGoP+Z4X2C92FkEcKQbuxIgQ6EE123g4b9YHVmeZXunEKr6VIKj1uGjhWE09ntSl0e
82FMzoOM+alu7BkGlJwow8/hcd57+uWYQ6ZXo1NyCeR6ufj0KI4JiuvkHNh20QBFNC9VVxo44+Us
WpKEfZtDDjh55o8YWOgp7psglLaOEspY9AekDw1kfIXBeE82p2+Z53DsXTUwV2zHLXd46lJM3yhK
VPrsk4bO/rzsYUzBvIWVOa0AjlEgDUnTb5iS14u+geBFjirStzuElZHb9UnvuFA7CKqO8h5ut3dN
pJj+1cUV7cvlC0tRHwJYAWHU1IsqMXKwezJo7p9ogT+LQ12RFqcBuvSqaLZQqKqnUnTABY1jOvDP
WJJcumzgjwZ6j+dcWfLMjSsEE24DH4cgXJGOKqCqYMjyRto1G+xUHbkYURdVLPUUCZHiuG+0Dz0a
P6TsKtjV9adSIVdmC6zCRIa4A8BfAqXJM6rK/L82bMCl+HLN2TJlzPVWVlaCEgVNCQQTUYQEJRIX
i03M3OrGkS4X6j02DUWdQtQhXhuvHKu1QNhtcVQHjyfgsTQhbUMZB4G9U9CMpQbflzD8yTpRaN0f
53zuxMgHd82Hg5ISTuywa3Hucug/Tqs01mEcFDIUywRYpa0H/AVRzFmsFvmzI+I4yBNhgQEOZBUl
SCN38d+T7c1ZKQrKZEEA8TKauLi2pUKNKohSNC0RTg/GtGGteBRNUu8Jhb5kO3cvV8XlJXZMghWD
fTqGcnkF1WofhNQubjSBrEmuj5UTwuwh6MCckVQis6SIsKGffp8nV+UCvx0fSWZEGE+WzWiLDBW3
pdbm5TESDe9smzmvDH77VRQe7L6DSk0rObjMRmoK2lS63zgRKvaPIlgmTcONIjw9x1tioeQFNfs4
eYzBZWM+1OAlPj/6qdJPvYswpkgM9efq7aXBqrGPnbrEg9eRXouJTy1IlnoVdvoyNBC+8hrI8UBj
atiytuLKptRh70pux3+WfCSjDITRCLxcKBQtTRXbvKaK8y1jY2lk/zr4omzf11uZeY4Yxlj1EAhj
cRXZzwy/6AmDTagzrEbZO5dBHUK3ocpOMwsXu8NbSAr7YInzh65juz8TIdwKovrbSKVDc1g+IKvG
DrVk9Z6ox79mHROhXn/bNNvKXOIMROYCXOow/IDd66QMdz4mO/mpH02UuLq2IwTDdktWuagrKrnr
jvV/rZl70SSx5JYa9ec69vVUBN2SY9aMr/dxMqsM7R6P1UyymAqAPVgocNYTO2xK7qJ9JrqjRB6p
9KxLTxHb3QMXETp/hwVVljaItJsyvFclwHtlc+bOVbWOc5Xizypkshx0saufehOYPniZI5iGy/hf
zL9bIjKHWd/9M5r/IbzTc0Z2RqagN9OvaPN8/wWqXqqrfQXZ4CIyATGC+dQbGliDHFCebmsFhK7U
zaw52qTA/paY8VJDeYWcIIQu+wKx4G6lWlv98ni3ESw9fjcjcgeqm5oBwBg+SeoIH428wa/FEwa3
tiM8Axhc4YxEsu5kHbnIEadPFeGmVykOEBhmSyrnEtBvGiBG2EK6i/qaNaiNFXP/Hgupgxg7z3eC
lfHscEllHNilAXlcSFRN1e1lxHJa23P/sOSTIxlPZkLKk51nyFwVEZt/iJIkSAdzR6NEuwBMN0nU
l58xwzVzme/gq8Ig1V4h53zZj9JZfGz9UVE9g22LOLUQV5rmc9tmBnsFTrlPz81QmJERfEvLm2xu
HAblNgXoKCv02Bw5D6VEFF4NA8oxeYZsNkZAIbiTWPAJ2VYSmDuwwS5YCl7g2bBPTA+GG77Y84XS
S53UAt/JvnDWH7UNjyJij1SLm4X6BzP9Nm33N1SBfG+DDOJ1kbKPompsUdJITnXcIwbwrMToK56O
Q+toIa1UPHJi5lxCZ0azKUXwJK28GuMbfXU5uRF1KMQ6v4CyaIyP/GWkeIBFXyQ0HMIBs2DoaT1K
h+rRjwk9UNyUFUnlcuF6tDHTde26SVrk+jDvzdi0GRqt8Qz3WMhChFSGjE8xjBkrSL17ZrmC8AeS
0Ngns2dT0nEa4CDzcMPZ6YXEnZhHJYKqMZH/rJGB3ocihjiT5wNEghF0n6N80EdqVdZItA9Kg7rT
XWNRBZJrrUL+0jbGerc9Mcpzocfeg/IBOGA7Xq94SYi8En/KA+pK4GAXqRF/MZ9KyA2CuCDNHdlX
F4SQYNYPp6d68Bz892albxrFahVXbOBX8iTfh7Uy8N5o1CRARvz7zBs0L1CsYHMn/kRrr5NEvMIu
7DpU1aJeSJJvdvMEDLUYz8EI4q5y+80tnPULuTW4mmVt1+VXThR48Yzw2p5thYA3l5FMqjaagYNR
mhHLQH224/29kxQh1iufurvzOY6Jv9t84sjRcx1KO1zNeJ2gQjMyu2BBACgabyhAr6cu/AGPfedR
1NUM3QpOv86niFxofSr/V5UHBFXNvl7p80eWgE2GLT7Tuh/Qu9HGgMy1eMZTElXCuiezP7SYr03h
lOoUmCE+4pHZdizDkNHkvcw4B2JrU0JvWLmT8t9w4CSEBzf9cv9KwlArswu32Mm0n6MIfcoqOyxH
OIkkDWG97eOsKKlsmivNHSBUWmxYQ8Eo3xzUJUMnNVY8MN6u9jfqAemxoSjraCXTQIl3BwPdrhNR
XTL2dMngKq3wxAxsU4dt+p8L4bQoszbGEDTRW/OFDPuEQVmOVr5K3iivreO3qomY9RAY73p7ENob
P+pjouUGIvxu1SStOveUfrFVIZOeba/lgETgBQdyE6SHFW4m7goLYDPbjPoCGu9ma5Z9NVFTpP9E
quxkd8HXKWa+2YeTee9zpKi5wod6ojqcJCXV6r3tIkWwZ5y3udY5jyjx2YLaAaBu81Dyu6Wv57Jw
4gkl03t5PMxW2TM77b4l4Hs6mwCLi1rTYRbWHj+PxV5P0Rj2UjU/q1x7ad2HQP304oT9z0k0wQlC
IMdiK7YEKryaW9u7UntTGJWmeHb3YV+Z5zhXYaoggGY9+EwsZMIZeFdKJN5TOZtsMfwAwEf8d7Zq
Xc5xjeMz8BRa+sXERXczej/iQMzBKhCcDNDixxp183rDM31sxzCSMh+z8d0vxvD0FZ4LI0dAAswp
gog3WJ5My46OcY+4DuvJJepY/p/JWu+cfBCK9Hugzm3glZDfQTYMX7LGtV7tCrk0sYQWWA/0rRv+
v1F3RFivXBO3wkJLnGz0+XQsfZxGw4beDa+Ft6Eixr72CFqkT7BXJiE5sWwQudx0hShHYYB7s7Ok
V2+nqddvE8caDewY5jJliV8rsz9Ff5pTNoYaErN/Ec0CMlIt8GiJNtUWbrw+Cs0oinIdeuhQSl20
s0KXSHeHQcFf4ds/hoTW9h7Q510JqIo3tn7JcBJD1tyhiV8HnPVFCT+KeZS8JgmA87j8QFrGbCfo
T2KPOQgYiZvhEJUHg1WxIJHYDayYGzfKydMOtBvohlebRjTrVIVw/yKhCr5mEcpQlPo08wZw/gDf
7jzW0f+nsuwIwd9fWqoAqjlkyoRW934VeKb2dOVwMv0RIwRigxcQlzAAVP1VhsG5aEEdMw73O8vs
Jx1QgJp5X/XK2lEOZxfPIu8dUh2KVud20MYUz6TH+kSP0NsJsu87VyBjHLdchPqM1iJuzxibjZxJ
RKgMymrmZIgvmzpKR0eqbZNetCWjvhwKcrdAmOByuUbBpjgTbHvObvzqL2wmyF//T+eaRlM1O/00
PgO+fRX2gUYlJEt0XkERKpVhTMmLHsUQbAtYdOgxZAmIYmkbsxAbOLdEAbUIMNC/6Y6ntA63O2RQ
8RkkI5E8ThczMh7T7hiZn5hIfGBoLNraqm1N8yb/FQxSaFZLfMZJF3mpUYQPkznOdFvHdeFTLKHy
GZjiV8UrUwOsYTURkNGbb3R5yWUXrY046V0XRE3yLpwE3gOhd5S3nqSZIzra+JeXjZ9mmE3MYjc8
TjIFXhYjsGe62Id14Lh0Dv1Yn69mPIUBUHLT21fKfOWwoW5zOGXo7Bb+PFbX2CQbMrUVtG0Gh+z1
WhWneiPyz55Z1lQGjw2xFy6QxwUUlNF1F8C8cGzZfuDMGi7XOYbujBOcZY3JeVXriZwuC8NPZ75i
m/6pHoe6QuGMgH+FZfZjSgVaE0Dw5EhyRLxmSs4V43MZ5D0U80S9AyhAd5qb2LGRXjruwWlRMnhG
SCye62fVgBkh+4MmPa3unL8VmgXL8CzmT9ygORFxMeuI2yOYC9atVaFEIOROwxPcWYKiM+jG9OyY
D7rwftbyEBcYNx0ooePmnj580neBFk1LukQTSFGyfuV3OLJr6ju5W1219qWYqi9oySTJUN9yLWTW
vwu8aTbcfzkIEI+7Jco+fksf5LiFqcEVvwGXyWjWHzJJIhuIflc7qT49TaJNDi/PblATLwXPGG3r
EZw4SImTh+HsopJjwmUWd875KKrmwXexh2VezikRlk31IMyZoNT/ZiPiq6nKxbsIk/hgr2qpYAse
M0YtIzEuoHQssm/EWLyYKlQpoG3JuY4oIput91hk2Dz/sGdrJkSEJxHapqaIUZNZoxBMecDZWmCR
fkqs2Y5WTDaYIcJ8bnqMiSNUbbs7zqJV2IWtQye3tHzva//VDOAMssow16cOqFy345Ii2tg5w5tC
mkav5zyU5argcHg3wu7Q9kQDopx4flhTT2ZmnALLIk7qocdYdX+Aw8eOkllm6vPKTXECGJTkDbUP
pwgPpKUwWJAiqXQwDYz7jrvgC6n3APJaJPqS+cuMau/jBazqQ8WNEnAhwYaDQr0GcJMI9N8+fbZE
EarWBNah2NQdnSR3CNELq4iQ8nDwvRmS/Es2ntq9YOVZ0SJG3Shag84DlVOr53+bNtoupKw04gQe
zPrlorfuAea0l3Br+m5nszfV5sen7jxx1S19iDf7KBL6SA/79ACRahTmTV1kyEAx1sxcCO1qfROZ
dmMCa6TS8XvfF3MPkM55ystqvjGtpKi9TmQHqKjVTujin1eudycXgiJpWMf/LolKXJVpGzAY95B/
d2yspgIl2BSVayIIzjB8P+5/e+MoEu3GNNum5Zx+VKPNQDgVSZoYVULOR/EScq+agLrwZL6rywcz
LFOTKAaFUW0cFl4wmbNiHHUalhp4gfV+Gws/aN16o7pt/Fr2I5wQi/MMS3J1nkxJ2JzZvg6GJT94
y6Xnt1Pa5Eri4NU2GZ+5EvjWBXSjt6EmMxKNCFHPD/+VBYJt28ioPASD70CokHLRLNyl9NmNvWQd
CyXz76SZwTx3q4gx2XT7VSRgAIfSzhIUrblqT0sZfeQkDwJMj9CHNA/L31ejnMf0Njx1cVb/NDYv
eWqKbczfTL5kSJ8vuYJTqaR69gLqvZu5fHqw7rMKGpf9sEcUjEKfMrHXoTLTA1bMaKuHBqzIA+D7
0lP38LupCgRaRm8neuiZ0XOYc26P5WSs5wq87my/hi91DB8FPGrqPozT2bqTwn/3d+Ubrs8DEdzp
IW6izta17A9xuQtC+o7KpOVzosfFMet1euqQrNb25SY22LbX6gEeG6mNPl6RMixLfcTXbpBx3bpi
NXsVLS8OE1ZhNmL1+aKZuN598IHZEtFe7ClGqWyq4x7Jxf3+WXxj8i+785h5X3aKhUo53u/wzzCR
MYRWXIySR4CzccDd4qEXykMiASkFCazVBizvQvPc9j1BezsCyulUtfGGLR/c07c3UlHHiXimfZ2F
D4JdMb1N+lbXwQkujqqrXVkOjWoICgi3wnL9mV9WKEtDfRymb2TbWpCqv/jSYGtaXt4yIwVEJQEo
5pysq1EzrJQJNB5h33bkZ6SvDQPfhnXEBcmbsJB2Olw+oQbpmGziV3rD7tdNieDGcObioohnAaLp
g96Zf3zvWRLgIA9d383snNpsNODQSsKnfJ2Y4uu96m8auRSjgOI6ZUqU1oOdihwvqX21pQqzSzrz
RnFWlv1rjTqPG3VqMLAPhiUARfyeC3SgSm7Twzf1zTlsLGR6n/Q08ZmQ9JqaE0Ces7od4zSQXnE3
ZRX/dotm/gnYIb6GjYxXyDsxqdtN7TE8QJTR+PBayddFiYPWom8FDYJprw0pHeIEF2hYA4SLn3Fz
BGz1zZZz0uSfru8IST/XmmBW8yCL6IQXGOa/cDYvxo+Nmz4mZmUTu/RGK/MAJLEHNIbY9vuP7hLA
BQvdXil4CjLe+X5NbTyftpXTh9xcf1i2VZmLZjtxXPG9nzTlu2/zHQPq8Ab8xyvHc7SmmIlPViPx
TtP1k30x9An5o6m/inFJmAzJKAWyF48jlOBS0xXHHxH7SAU7/4rc0/w7lob+CjJbl8EuaLXJwpHG
3kawfMiyZbwtZtKkWfKAtkO0aawxbmN2wq1AgfhY5KmlHrGYuoIiGZn51oe3jLM9dsq9bPV/HWzY
1E+djHCoWAUywbPHKMnTp5EatoCBuwBFSc6/bQKKpDvSJoJJFL5mHAXW2KS3spWe451ZOvo11253
opd2Lm1yXKEQ8XBiFaJziuLJl3nogZQiwCgrI+BOByfOJn64NlaYvzSWniycq6bzZOH098yzETbP
Vm/ungZnrsnc6tfYSPIeqpb2cCqJC/nPGqZKWKDUgV+tq2VlYmr1jIIHgjZQmP+SCA4XyYmqm1l1
Js+Iby0EhOr8jKH+VhDYJsaAZ5fwWwHtpYwzS42wVe9qFdQXnUi5Kk92qNjLeYCy0EA5UYIzyzmz
op5J5TwbsOzdtcGEg3BHrFxJoq7XSGOov5ai4Kb6sGvwX3nd2YsqiYdtwQldD8VKwMBl+s46eOiU
W3agEEir4Z9IHvQSvluU8FfJJ24mNteXzkXTHciA+IUaDLXDBfuLEdaE+uIJhqloYyoC8e1oJ0Vz
oGnQYPYcNOrPu5QF0d/j18NaUYQMCPrJZBSbFt8aObcY2zN93IM9PTlC+juMTundAwKCiuo6doz1
X0tp9lBa85eraii4g3mV13JCSE/CCmH4y1oZTE+Xb0oAk+4wiosq7abeBIaY7dDqdhWWSaQtEt3m
LlZYcADo6yp+2dM6yLalPOfWh3smGeeGTfWCkUi7S7CYraqfHG3x0JuFi0tnKBEMbXE8IcQ1Jpnv
CvtwXzQ2zJUwzv7lCJHW9curPuouxACxL/s7QeMewDSrgn1BE8rqMomXp4+VEttFBo/VdPoh7ymu
d3l9p/mNsvd547Mnnxx1VghdeLHFDSpRNx1CHZr/sH3fpl96S36F0ORZMKljxWtItDmqQmSqbTSW
0j0M9WVcRHI7Hcwmx+cGl9XjD/LW40vijS4iC+vjf5rWiNPAK/KBdty4Ihl3lMSopAGy/F91jKgK
g+s65+rxVd9cH1iqxIycHMvjp9gyH6Dskojk2Ov99flD4uA12SGw1jksce0r4ZXxTKLzysxyNXWd
/mhKiHgUVbTJvtwUqQfEC5kXs9ak+/2l3DHU5ZHhPngNenGx1S1ysxdVDEDoWgVyLiODQp4B4w0k
U6aDWrZG9jMb7S7zP01fHcdPBfBuKf4XJ+yWkBp8KmAGYXK7fnIY6usO8K/MXejNr3XUApyjsdae
JGRgmo9lITkkYjjNqhgmFiQm1DorSYe1AgUU6pRitS+beGQO3WcQvMzJ+s4LFAgVgUiihcudg6SE
xgbeIItQ5jzMBFKOZBMICRTGlnB5aqfFw3r/+o/JFYGSdAuZQ/eNjBwLE7KwKjS+CfV43UNmX+Oo
6VIrXuvjR5Feg/r3GU49Wj/RckAz9+sESyAB9AQLypuCTu7/hLGAuDHa5/cDov9gzrbN4ESxwUwW
HYCv8VioFmM4OU+gQ/rD5YO+2ZoskAk+M+tn6Qfa+ZVa/t0GRoj6Wtn9p4iEphpoF5g8DOw0NHji
rm1J4Wb0IeGfa0v9yp5UVanlMyYf5ypZyInWHMhYab3lZfxx2y8BP9BENbAYXzrS+a1j6sGEtqbm
ReC/iXdiJaeAyPoXas6IJF1LjDtqMd7HbLWN7CHnrJ7MlHpT2c9RFTrBHpsecilR4BnX6IY2MloU
Wp37EV6jbFF4Hyb+QKLBCOR7F5iWr+X6z41MGEsyf1E1yagYTDh/Uj5rpMckax5O5/cO99BlBoQ9
8OkxDYCNguBKcPW1wroE8yJwcjc6HNVqqaQnGjC1WhDro14uvtFNxUSF0sHUBn4Lb4Z/0MlMXuC4
753+G7FSIcwLTcKv2jCPAih6XcdGlGbkB2/YdmGut5zutzQd2Nl+Aq8vKXVGLAHLpig0wVCPB4RT
T4VJksRr/yBn6IxvjGWLPeM+z9l4/VgsLwatQiVKntZZPOjbdWLerk7VHCnltMBbkQUI7TKodn+a
Xdf/zt3E1Z564PLXYLc3Sx5cJYSvawgYvGnrzx/xkWlsz64BIgBLpTElV3vHEOMeSTMPGzm4TUeG
Ilow0rgdJHw8K50Z2dtAUgIJDHhZBGbox9d0lBu0IOmvn/jpgR/ZP+O+QtUz426ATgED+z+pPtpl
ADwipYQXShCeaV8oTaIAxIClk0wOWUaUo5WJjzoZfIfQkvzsoo8K0hu5Rbht/C3nmO8SmT5Vb55A
BHGm/B0YwZcVGRVcTLWBg44+gPQGlXBd/PKyDSoI5/3FAN/3CL9lQWZLggyy3OQYfWfX1f7bHEz8
kbGK8ZEblTArre5XZ7R6TQJMFug9o0P42Uutta8akkzjIZhb36jO8muSe1CiSSvhzNChoHeDzEdo
jHprCmuhZG4qpOICa7aSgJCXk6nyzZlfoyxxrOHVcSl07N9y/slJBBoFP2FNrL5jocBRdfTEwceW
cfc2qvzQ2TJyB4sV34iq/yn12SOtd4Cv7Fgg8MFk/k5STCQ4Tri1WPUXGH7xCbHX/tjnitk2zCPy
VMu4pq97gJb/uPxgKkIC2VHwv4DKbH0d3IroR2lNkZ/npvDE+9DDL0CgPzj6K01QAAhZwDHNwM7j
Udh9s5cykgKN3bLYI/Is9Z9dcEUbKOlHGoyAgAX4p8ElC5LZkp2sv0eP9aIuABogn2t7CILsNtWk
ywU2ZfVotHBGu2sKtYnt9xWHeO+8dB4SxIlu3v7JS3WIaQ1FbQ+OE6NNTv8O2o4GcH82HITV2f8p
zsC+M7p4P5f7wVRp0s1TZa8/x9J+e6rI8J5Fy1fndZNCRjDrdLpkjG+fH+D6gpZhdeBkLuG5u4hU
65OxOQW6/5mRwcMFJi19yPhsPaKCo2s9NjokOJgUcjeBkV6l7lk+zZaL3Fv7UbdjQUQfW7d5UgkA
0FreUwKDmzjSf7qWTuhzh8lrsgh9NzXyZPREb6BbkQpxPy/0OMtltAsqOnf4ges+NpOLy79JEXFQ
MJTYXqvEP10f2eG3tDzo7QXrIMIxtLFdZn0otyiZA+9OxVQJzHH/OWM6x+9ycNxHGIZoMCov91Dg
sNrRDM+NWrmP6VR17OUSounuC+bjRzep6OuSGz9A0dfHd13Eja79mTjJ+1GDvPi0P4yg2nWlRHTh
2otBW8cO5JZxzMkcFg+1BMk10SqhvYUTQ9GB+dWyj5aljb5yEGjZx/2Zm835Khis+TTIYiPvdZ3P
e7wHVEK+MmA8JeJkfVFYyzPeACcV0nXTNEacIzkIXJTTb8Imdd4XIYpPjAbGqtJhjSZE44ggKEHd
PzQ9Nj+annorlCOLrW+ae1H+ZvgyABn0B9L32+UhEuU7On5DCIO9NSTgAqtEObuCmzQP3ZKol0Rn
H1090gEeuhtSNknM0SgmD4gVLRf/+aqzV0IHEUA+VYrYZYnX1aguFCTvCcE3BEBX1uX0TlbxxW45
nzZHImPSNyAOgUVuSrD/Q5gi+9xaeBD2dlYgJM/0KDtciuH4Yf3Dc3bS6qeSIG7HAwpJscrE87XP
1ANiHPJLJSdqIk8ph/4kgM8k6tsvac53PUC/5pPoyDijFX6bOVEF9uFe8eZxeX6UBXXkYQSa2shu
4gmyCq782bC4zot7w+8cxPKM6AHOntZ0KAQ/Oh/xQAxT5xZ9UZhmQkenzo77iT2VPJJ13ljXWGgi
9OaUlgt45WVPIWpAKIu7hh8qGRQN57QUNsqcgxneWBQpVDoiYVFYR5Is6XaqWu0xui81ZJd4q9l6
TanlbJs4Z/2U7cFcgddp1bs/8LkasVOB9v76NbSCOhcsmDw0MxXLEQZPBkwAOBEDDZA7ibDgOtpT
svoYpc+IJg0PHlmjZ2NA6xbNPZFH+T4zu0mdxLOxdhFz83Dv2HDpamPT39QX2jFI72UBQ/Yl8g3n
H8HwjPxRe164n3RYkzlqsajm9FqXPbIQQ96lKKBPKxRt+nams+6Iug2Db3tmgG3B/rqil/1xAJ+G
wwCDSiOQBtlzRjbc2bDpwGouj10wURc9Oqc7FkqdRn4WS++UmFh/dFivvSDq3r0UnIXuyK3X39BW
HAxzR+K+Zsn/4XUqzF3T/3/JNV2DvaK0OeYYIlqJzwQyN3sTm2fPXOI2e9O3dcFUrNosBGiRq1GT
5TBKEV5YEeoqVlfWpwK4ZSZiPIvVAeEEmDkSFzMB+590qOYPxpR0Gau6A7PycxEqoNj2ZKaakmrS
5XdlmXj5bRBsq62AkO1REpffEeHvfhcahghl7X7q30bxjdPM/Ijn44ABzm3U4xW+DaQSgn2tx3fa
kgpWmm6vLoK4Kj7tgUcIRFJzjzdl16kpNbXF4mBJfk1aVsiKXW8qEa3h15FTr+HSQdfZrlFuoKEr
Dg+Og0k2L4LCCj8uTkEkW1o0/gBLDEjKdcDi0a4wOIxnZgu8DpsPDA54qHGR00I/suIoPRoVwIIJ
5BwKr3hOR4HflTrdpPFqu933McdiMQmke+7wQH8MoHloYdTL7iEuK+o8yyJ1vjHAPzDO1f7mffpJ
L2Tu0LxIrR9tmN+l4ppVVlBjs2xHAK+cJ2oBGByKnS0JYJqlis0FDGC7iYPYFqMlNRNSqQy9jSrX
gNayTIBPidhyPTbCA6P66mhdFMBmt1rzGiwh2x99ncjDzsr0fcqvRarUY2PNP3MfKJMIBsS1DkOO
+WIZuWAwseIWBYxTpMGXmK24X+sQcSiEa/7VbKxJesjK7Cd9ca/fZtSsSYTOJJx9fIC1k3p7Y+QN
VuLaYuzRK1j3eQUHuoqKtJr9uMK+KQab3vcaJ+eqxEBukjOVc7X/OOhNn6uhCUN1HpFrb+bfUUZx
sOwiMm33dJXUKlhrnEweVMfWYFK912g2ZRfVAjKl++gOJ8qXHnVYv8Gb9NKJKHShBi+IJWYzFNWs
BSsAw8j8is3QqrwoGjWjqgk+ZQYbCFOFDzV+S+sf2Tl1WwfppcqjjjmqJAmQ8qC4HlDkH7jYYZZW
dZHi0mlDvExnyJM13WIGS3i+ADA4NMYUqXuAwYb5XcrLDyVAqmHgo+dqZBneYo8e5A+oRGMFc0PL
7ULerIH4yzcyxs6NRkhIkfgB5soTNs5bi3rKQob2MoMFkatTTa7ZqRyAZXkmqG9Y3ncyWWKt1wIh
IjKi0fvdFzF5jopKq83V6LJ/66hWmhj9ZmBKjgY28FEjlQKglkli7Ww/GZtfP79HUAu7+bX/zyN4
x7A/Ya895ZSfWHI9b5zhArT2+Cd7AAgoACFZR/8NQE3WQWQQPLteENSenVMAzYgNgrBZA1A7lhrl
0E+YZMQ73GnG9T6N4mjMfvED0gwxD90gwX9k+rEb3bT4P1lNv1tWIXNDB7+aOySkn9XM39klViJJ
XTTBgiYLXHQrucykxagXA+6EnN/D+UIVeHPYBhYG+r0RJSjUioUkRxTi5KyU/BkC+anTeqTiE2a2
wXAtp4+cGonsbdtn9l2Pb+paB24IOv7QxfulkVP9BmEm5W3UjHNR3gwnwN60hXssd/LYq3FI/A6h
xFh08ar8sNLxMSHCT7abZTcN0sD6CJO4G/oATKKTq8itQ9ZSoQPTBdxYqsKj1PvMK+FjO+cSEzGJ
+l+nKAQ6N0222j0z6tHFT7huBAULzWf+X8Ma/Qnzcjw8bolPe4S+uj28xmgXrkagjH4qGlJURfc2
XXV/pC+BI0J/rxvxd2vgvUx1aIIWfZKDISx5CO2TiNc+sRuwpLxqn5E6S5wZKuEJyGyrXznssMLH
RzI9mS+EwvVtkAs4BegJuxl1K/YYHwTLNUkvqcML7gLpG0L1ehnYJii1BNj7kyBLIs5NBf9kyG7N
MVlKNa/swRwepvHmoqODFsfRsGBZ7nUKaw90agdKGnbfAH+7RSFnnETH6EgtOUTjzcyjjlxGcoJW
ho0gcJX1prVHogRjG0Zy/m2xnUlsVQm5WR4TMt0ZvPXx4p7Ob1kQ+ysMydjTWBriowt2TCoJGQv/
oxTp+w3TJwOjAXHBSbpGu8m+jN3J2bbBqY33YfXwplDnTN+jCu4rUmCIyHYfxwLPRHDZXDwFMlIl
WTr2V0RhlrBN75D8lnll3bvFC8Cf1zgoaqgNm01UAzY09m6SGrOcsLALuJlTt/k7DUG9p3UNhb48
3KPBJeZ+wsChM1mXNeJ1M4WVHio6RNeLHJKssGkuZQYXNfN4WvrBAMygPN+XCGTWR0N0KT7En7Rs
GjFl53gi3jrqyE8yP0rChB24qR+zVvOZJW8/RjKJmQFe+xYjSX7/vAiVTBdw+6ee22/B7k6EGF+v
LWbmQ/IAu27XGu8wvSw8wgJ7B30qazKDLU8YBFOLf9rZAtQV0u3C1AphT22JOU/CnoumVTF9G5Ny
uiSJ4ykxXDYOsUDL4izN/dcenToAydQWN388rdI7UWwRdJaIJWrzNagEddorYG8vB6DYex1MczHu
TfA/LILpBe7aTI49IoZlGELNANsqNN0w1GFtYmHMM9GSPOoVPKTYTr7WyPg9EeSKQalTg6LHZgEw
qZf64sqqo5qA7y5jEqJs1YVUuQal73NvxpVUT0Bcfs+sJwzdxglnzVmcWgcitoWR596+uP07W84/
cjcU0+fCV1hK7Za2MxvSC+ML4ymeDbBziSfkciYD07V4GLerfx3I78J/CPiK1zIl5h8SjeQLGE/c
1jndUpLRnb9ReGTaGOBbCmnGTQYS6NWKowkHjbnUoMtnPbJT7a42eDsavr+7J//DhcSe8cfLmFWQ
h3Ai7PQ50Kc2DADMi8Pg8jxZuBDhVhhAiz31rL3sa7rkN/mnaHOnnXWicwP/ljfrb3dq5RET9YPh
HSUs+Ra7E9j6CCaherxW3yM0jzU7jgPoXc/J1mbEO5wGCtLd0lvy2BNRuF3xLrEuk9PWkhF4S0Fk
R0rQA/w38rwVmt2hKDcXW9ll70oOsgxe5VGXJensi0f0r56ijO4i69ehWc7FPCNABf82xdEOzR8r
8YSUaTMYa5mr1zFRePTy34GuaqtUpuPGHmtrz50burnCLSCTnsDDHbxVeDDM+dnQb4Gf7jyUFxoK
Ysj/aw8JGYSqdo/+IAbVIFBdrOoWqV1MaPHf/im29VF0fWzMHKdJB/ILVJLLbX9yvg1j/OVNrTVa
HSAni5wMuFAJ5krr94NeySleOK+y65VXe1tQssSrstWl7crJiuuoOFgSRgjf5ymv9BU7Rk+1q5qX
0zMOeR13KceJfp4DfzcIvtmzwIPi3s+HnhFIXq8AEY0YXXbsaKC6lmSfX1llyavf7GYhDYBxVYS7
/NbTK2gF/KAgdD/CG0h9BWaDktHz0tg5TLU+eYeW3WTgEeVkzbqpJ53nHmXWbvRWfucqqm3xgsRL
zSeZvufB/5U3wUtNARYNrd8l9EsHNiB7dzUdKiVtWc6vBW//tXjVNu+bu3mCcupk/s4MTFA02gfq
DP97jn5dVNJ9YbtRLfWOG89gzsbE/HTGkG0AueHmHSvPodjm7Y2vOrH26qZI9FtIjGF/a8icazu4
I/vgz1Qert7V8Wl8gqQVhDwbJobOXcOg3YWvpd7egUHFcFXScT6NSg2/AmQCl//dwrCyTtlgD61c
SDiA6wWx9nEN7SEH4Gwj1Aqn5VOpZg0guzdpZ7+xKbRZ4MvNGwq/kR+8eWgg4fc9qmUqfLUGgmxR
r3dyp8wy/SSN3Dx72r/zaGmU3zfLOvOai04bHuCg6ZU6G+8368Cw7W+2G+woY0HCMxQhyL0iKy6O
D8RriJarZmsqXYedJ9Z19W/xkvAcmN9klh9m1l3lGTKWS4YHzaj9lhrgsc2WcAZ9y3XHRednHGEc
NuazL2LJQf26+zAe8PKePnFOVe4mNZfI+O8ZyGo5p+MJJP9hQTg8uBg2p1y847pXFcqN8laGttOG
N9q9jU9JUzEgIeAGY3lHdqMJf3xoNCjMVcjseyqcqQbSpCI3fxjlZGV6NX+jFyvmJ3afxVzLFkOq
2MY/DYOjNo1nZiTVU53JDB+RM5rPf4wVo/OmaYbchQdpNNsI21VFD1KVVzi6cnZM94M1Z+o2bcR8
TGvpU8+ORZVC9Yp1Xbt0mfitM4bLCOe1SDKqGdTJrRJczPaJskD2rODx9OG/hWXdgBmsxmHS9JJf
CIh6IsSf9PIMegQY+D4WA7c5lbKSBLCF5L6IkUdY8eX0YOC2a5lEaDjHntmb0rDNxtbfk9Y8/PNu
SBesQhrl/P8GYjCtDu7jEHlyocMww+TwgEjBP1MmxkDbTh9o2j3fU6tOWASJNuMxebjCCInqEAXh
tbaSPh+4uA9/a6ByIHUumwIAuYpLiPQ1pce/nQGERAlDuoq206k8TOLRniL/IyGHvbSBdjpEPz92
a3u6NNao5jchMfJjnO1PSlunZhMMbOeQFnlAjcGCbGctrbE8NIcV3SYFBWhAk1MKwHgdEkGBKg9J
LQUZ5D2FzQM3lglLtzHDLslrB82pB6k0XktJwIjSOl0Ot7qBcVcKqQqEEKlnCv9wSCEPX0BNbIzE
8Df4Eh96G1QowTqyPfLvHi1yf1xpszcLxK2zawcvUOnq4WJMBBxoy9itFmft7EFvXVr9nyqKXV4u
suAz4go3KpKQapCJfhOF++4svJ+g2QcDoahrSiha1rtS2XtACgu442cmgxNBSFoRBX4YrUJIpGg9
fIKsO2PpfrU3Xq/4L8GEfLcF9NLVZOr51U81YpxJ+qENYs3Qg6TEBpx5JbvybASr2L0P5tPDY/Im
z206AlKAH93Gbrml0Tict/WPbmCgfoes+gKiEPcixC8Xi487+A5YxwWbFuANHGN3SvUutAvj+MHx
1kjAvqRamLuUkSf4IMoSn2Q+yBxrbvc9N/BEnj5+fI1tK1qdwLqMAgDrv8C+pe0B3xrcmEQq9DKS
R6FjHKwSB/+MW93SrUdKObBaeJfYtCv57XPWaHTt1Vrk4vFeZYN4P/v4iW7Gy1tJJFcaXD0fhOo3
gbkBnBCNuyGDZDDcPOipULrr/D9VNv3svDRNkPGTW7r9CiTWT3u1uX6n5x22zdUhD6HT/oqP2ld0
2xP/0FRNAVS3mrhS0ysd3DqwI0TUKee82CccFEu2yEV9gJWUjNXYy2xIExDKIMkOgo7oVHUR3Flm
FOEJOMfPRr+CNHGIk9IqcP4Ku9oNIK654igjXk3eu+G+6+dFhDhWiZKdUbalaXJgh6YcMQPn6F5e
4vD7+RFrSafl84ZyxYY8yyO5dK+qIoLqoeAMyxHJ30nTmTbguEy+kwAQpLKPWcHXfauadiij6KAr
/Sy0hkXLqAnR5wiWSRqw5juIrORLw1Yo8KesBtGehisaJHnGKbnEhiKOYWPzKWTZk9WZEn0GTSrf
RyJqQ/nU+C3CF2lXZ/6ZY20XobuFDTw1xEEHv4rpGLrCU6QexPVAKtK3Gd6/2J5u3dKSXGZp1D/Z
cegcJQDdu3Z96nsnU60wAAGGHPQbIzPyEekeco8Tr4rJ0niR7OIqPNSHPk67QJC0P7uTzjCPQwPC
7TKMcfie9bJ0MdnEP/AUGQKBCeTD1TApbEbUKTktBAHor7wqisxL2MdSxgBFky4BLII3kv1FOz5y
l5BIgFUFsycgGXy5hvus3f0pmguV7tCJhnoIh4USRz75xQBlcxVCFfI5qDLVRIEt2czF2LlKLVHl
zRcF3pG5L3auZPYo3Espd/u1j/023UFgi2rg4fWZpoDRA+3B6yJYk6AqNOHFTslvJJhMjJ0Hc0GE
d1e9qbZoaOviBpJvHBCNCh2RiN0XqwKL+QroJGm0GZTkjGgam0EvcaQrtciupq8x1r5DymO6dmVQ
0gBfALe8hIysri5tvCuGZAzx5bbgm+k/+8wTVjaJqp9mu3pu/TiQblp75kWZo2GY+fjZrElSQUdS
ZcybgUW6wo9XrOjtxfEm698QqHK6s4tOyCps60MMPkIl+B6DQ76G1J1CtrRDoTIBwZlT5NYsJG51
cSTy/2wxDzeuDm5Sj+mGfE7I28kuzR/QCdwnz1+3v0KvIK9ymrZtbNWbZL/MfdEDhPqCBumI2rPk
xkf+3+5yY5eMhr2ffKJPYkS8gzI76kBP5szqLDx9wgXMY04TYIBf10dvgctYJvRBQfDx07XBLqX5
JLmkCUezufvz19MGW20bKQXA7GEhY6br2MASOSw2TI+S8dfocSdBdGqh4PX+oZ+y1vsz/NFBTjuE
tA7fdZXx1IJV5D6FBViZtE8/CvKfnecNC+XM7NwkQpiDF5YXCrLCs5vs2YEV9bD8nG9gdwC/QnI3
+s+/bnqvB0ipAM+Rah85O7kPnSXZMXw/paAkMs0jVrzybQFuR0uCohjqck760yzMlR73tqFT8wuV
9CKCvVWL9NahI914SbgTKkBy4AXPg9S/KRHBfdRc2SuZcTe8cccRBc2elYcjnrexc6kFfQrGRGNC
JvzeFu23vfi1VvbF5HXpoMS8qMTySnl+uLEqpjy/9Od6f6QnYGDFS6iDiu9rt3Yrwm3+mNPRNHq2
lg2qbz1f+GINKOnZMsjJ6VFja7/+Blvkz6HbCFRrWXs6ysgHfqJBgl/HOrMU3+gzFnVHT6EKanxK
c1KdADB686tpXh6bmfIiJWb4x2vKAWdpEcLA+LwTrl6F4QctlqwaY6SDmL2KG9bWfPMZKtoTEz8o
N7ixHuYz/DRXwXwoNN1Nj7SOzdf3OG+YWjMjiNTR+EBYYrLkEnIYlgY3ub6YiB7Fu0HquBlWq+2H
suSendjD+V5/8hvSX+RI5eqVClemgym2yqMlCjJCB4RLI7TqTPjMS1X3T2L2CacUm9yy2yb4iEo8
sRpPb0K+U5fRVcxM+kx1A2FzxKTKHOl9IvaWl+bc8w/ELZWJEIHcnYbTSw9VkAjItQXYH3WTtrl8
X3vXA6uxHQ38oae3Qggx/d92zyRD6SVS6F1xjPQxp/dMr5MwfVUem7UVTZG/J/BEZ4g3dxcu7+VV
v2mm07M+dEY0n0uClA0nioANHc4XZTh4bjIjcksyEF4NsFrNiNAtlZG9OL+7+abQrC/LzW8DBsVW
gcV/Ix/734/aTEBTiQZtr0Y+wxV5LrYbZH00zlrnsYV64jioAtNXyflZ8FU4fNZ1A8d75I6/e0Ee
FIUGamEG/qvxfl2xjnAuFNGKys6SWLr/l2BJ2kLGYrX1+m2033lTs0xvBhZENuhLKHe5zQ1by7XQ
aLB7x1QCBNV5mCNgEqiZIMlM7hhI0VQYZvw2yZ4rEaO/qtLSgVND0BUmvlWW0Hv4q07PuUHTIPF5
ZveA35+LJnDozcSiBRXz3vTa202TKV8ETxEVYP4Ji0nkQVAHQLxtoUvosL5AcgWm9js9QU+G6IiB
2kmO7XflrURpfAcAQzE2UY/VcrekzJnDXmiKQGnKcABPChfa6+r0kH0xibtBrSY2xgYoP87AdTpC
FwGhX7wxUxTBqNqRpgCyvcWDvhLd48uUQxRcaK7Fdeza8ckTqkVu7PTst+3biZQyHZMEFO1jQCro
7otiUoGArQebIBBK2QyK8yRRU3smEWvk6ZrvJEQZJdDm/pyAYTquBT87iTJMLn3iNeyIk5VtWtgh
iQvwCp3TATMICMeQYcqn7wZ2me98bg+V3qmx6CSnF/CW0HW8EfLFDAdcSl4FwdvMG5i1vTZhSRWT
R48SEFL8E2sSpSXa5QjkMx8ytiVTNbIiCk/joCWTmqpXWloPpvs1tcI2FMu4QamD29yAsSbk7gBq
DvIz9gsStO1Su4H0o3vtc5pcPH2PeUF8AnV5G+rb9slk4t6VPAWSO7QAlbUKzxxUGE1fvLqNQrT+
tTtusIenFJLiGsJQiVFysFVEM6V40DAR+f9SrHkS2+0+8LRXZroBr5NspYpjdm1ao70uxOMK8vKp
EmA0hxVxTa3lZhyFT8vddxfZrGiD/MYeIyGRR0jA80oHrH7n3+YAZC4uLWu4IoksawrJx4nAp40u
mH/E+lL8HNj7LKRtj+xEvZYeKi7fSyDeECapWEkwnxDqq0LCxiTQ1hW6uIEOEmJ2eB6g8tRgBoWK
pB+ZebhUQHjUM/SbpBZjCj80qby8OOs81KItkfEiUghz/f20inl0KT4pVafg1feBLwN8QNJLyMEs
Cts+ycE7MhVZS9NIKl5zJ1Zyc/HuOjkbKFDfelkQyZwoiX18sBUzfwBRhiJZrXHiOX+4G1kyFEBB
H9o4lWdIcduBdc8E70u9yt3iqtCcXjZjOUy/W/aWQV62zVPtlpIlsFyp6ciCQegOuHY2R7o6D2o0
ZnWdID7l3T8/6jjZDwhI62xgnaTBcDgwUS9jwaYLHCDB+EIsy/wyBXhkVG6Syp+n0Z+C1S9BVhif
khfN+39qOkuRsGFQZ+pmqrH++U2X1sJ7WEw+/UeXKP2YRQ9ygU2koR8/kHZaxzVcj3cA4iodbdQA
5Cm4Q++yXfBreLGKlas9a6XWyUTP/VziLq/goOAyuuDqAxhw2iJr7RneBr7lzc+Pw2Etlhyi1jGM
/kYHut9GjqHO8n9awBCXI+bSJjBycb5GFMNPNc3U5QGDnuNcgAUOdRfWnYAVHuMjyHwI99P9dFGC
7n/JLWvoe09WoNdkN4Ecvo0VY87QWgRsbaLE/wYfWavSZ7lriAD1PwcWFM85UWe02brykVFyzG2L
RQwaKW0KLTUsnZ4qw5+rBbrjcjZz8KLxpEAZZirm2o4PGfWN1AVmZnMgCRc7QlyG4zpz+RfOMdKM
nTeVpHFnVezi9lvPCdno+wWeAZb41MqSFPHmJ7BWAlrZVnYRgZbKQJsJWmTgErDLVLheCXEYOZnD
RWkHmcALRcRrknJ78MR+Wg9sVNnF3lXbQP4S2+oQpjTOi6H4x7VOtvBAhOf/tmoNG2FBVYHVk16w
UnR2bUvXQA/oVpnUrAzYWnRd7G93CwcMnKhTW+bicsnYjSjseRUgypNY7p5PyFp5cnw1Kk8dkAhL
No6JCU02kWUP8qUXo5BbSWTrHnGa/GqYTvBkcvWcQVGITR36Orr0TUjbGkYyOIQ+F8RPhIaC8LXj
JFh10ZyZcIUDayaBwjrONOA5wPq1c57NBy1WRRdIC54tCKE71Wrmr1LUpRPcYGqw10g3oyERO2m1
ZRZIol6BXAtGm3srm1N5/Iml8OFn0GlRUJVm7Anj0gMu9xSK6MrMPUIAXnlNGizDEaDCJAPlEzDI
jmXgWcJSliunjQLdpdzvlJWH5mb8U0cmjKh6qmiCB9a5tC85wD+nALEQfKc8cDeI5eUMQepmlkAM
Oz0kviOqbWsA5KtxnIvbaTXYbWcP3p6pIRUGz6Dvqf0ifVFJLsvc7LpMO3GWxQXHiT384I1+BEPC
NCv5M9AbelPmhFmlL37P277vFUhLQeWq5YUccwlIiYpG33qXXNZ0iMyZ2eomIB5p1HpMgn9P1GvY
4F+nH8Z1tsCClqCd3KEVB9Llo8AGQm2Knr34NqfMoaOoTeNMc4OGrXN1kDLku3jYVwcTBnwVrjSG
ZMSe0jCzIL2DsHE9uTQIk3KdqEedVKo+Gbwrp+hCnxxnRzoWI2nReVUcng1KuwjluHeCdvkkosJ8
rgomcqsUCkXmSm1XovfrVqW1Tb/Ul9TNd72QE83yuLz53T9Q0/wrN6+/1jDJxFLPG4MuSjXBtIDX
bzBHTTUf9pHSH2+WBt+PEGxPjoWnnVxJ1b51La0nHEuEenxnSi9ri1++kydE2oi+HyRS8/XeX4kY
x5+vpR/jxQo/lEQv6JTs4Z405WH4usxkuoMsnQEQT8zbqT7xlUkvjmzHsmuNHzlVRlH2dkScpCDg
eSHKQTj6zPk5ApAfnder0muJhdUXzBxKsrWaQxCnCk7AohcWTDwLXa8HV89UNfCj+wFHgn5zjbGW
Dnx7VP+9QdVh1o05WjD+VmIz7ns2PMOwm8mq3b1CnTcTJuygIE6vqL+Jp+XWbglFuzDoAuWEuU4Q
y6NhYl2UIdm30rDFPyW66JGaCMeBHNYiLxxDc4Ga1S+aC2gtLdqnweFl0rF+3GAwgGIFlfy/3FYq
2zF222dtWDRk3hAbHRhIT62Pfax08pJmu3DfpAu6pdVyoG5eBD8bqwd+ScaoLdg7h2yA5bw+ZxDH
dpyCkPTZvLzOuxqaHaa8HqRpa6wScznNj+iMU39l0CwnqesXRiQYF725ekoQq/MErnLVOXzrbfAt
F0fX38OHA6illsfjOTGNVQWFc3m69BIt1zp0iRm1bDWojR5I/m7UIkeTYOCVgGO7q2HYivR+bbJ5
Arm+LOMhM13fEk+ii26KgfqR5oV80TEWAyjWN/1iynqgkdG8tkIaL1BGsaJePw8i7oHgae6cd7gR
l926RB8qlyrdw95/eXrmhH6gWbprJnYcZvGA/GMN62yschNNRCkfb+PLXA9Gr7LShiBIqMrRvsm9
x5338fZGlUL6BF5oFcC23wMGVDljh9Uu92Gq9O9vPexOvnv+tMHTa3WNhle5vl2SQeIOPa85Nyhr
yZS2Ow1x0kUHeVvAR0sMotueEuBHYWEQ7+8i5h4vLJvkyzZTtB0pHkaAYqmMyLTO5I7fAaNJoHG2
pfjDlLx1cs3jihDmZ59kzjufgXvqWnzaTfrehBf8u9Yg8nS4bj1mUp0S5v3InJa/+C+ZFkDacOL4
hk9E01VxEZeDJFiRZvMVnSE7Tp+b9ozVRTwD9piBid8OILMgSSmv6wwNlGIPP8LkxITmxYlf14l2
il4q9IjinR1d0aKICj4VV4wz0C0J6GxyVIzaQALYYcBXo+uT31JN5+/09DYnhHX2lPNc/zKx/Fus
/2yzmj+x1m3PebMQSXEo9qEr/nNi0zYZoQDd5Aa/Q7+oSmcAJ5sicZmzipbXs0/hXeXpR9bJOTWg
eIMyfIM6oUNahDbcy3B2nc74863U1D5C7m06vJpKw0MLE6RVTyFWJor2L/3x9fqkKwXOqx6UHV6o
9m7L0P5k3kISsGD6x621AMn3ZRZMTLmYIsQiI4XrhuXabNsX7g6VKHTWqYp7CWvCaoRsTgCjdZe4
HkIyT7IsoWi5VM9TMPAT3BxgB5Vew2vMISb22cPx/AATR3HUQh+rezPQBptlj9TEArN4f7YtBHai
mu0qBtdy1RmtV9j+2Z9UIANglSV/pEJn7mRedDY2z833m2g+I+jsF/O5Qz/M4HJFW0KMxn+KdbLI
Ma3RRIF56QhIuIDb9CSbuwMxmdpy5KqHh8iWr6J6F0aOLS1NVNGj34EcnmDiXuc38+5d/5g9wdmp
H58ks5nqYq+iqpIcFaDkTUIdZvM6A5tAp6BL3Q5i6i7s1oPOQrVh0CR4OAzbJq6vI/3aOg9/fcwN
kiupHoZUqb6XdPggOx+bNMdWlakN1whAsjBcOG7Qi8yqBjRqD6veHerx+hd2sxkCkC65KEV2fKgK
hO4UIlyG028xN9MAubrAf01P9ea7uO0DZOqTzQ4UATYcpriNskzKsvqpm0TjeNKqmZmWGMkoCQDn
OvcQWbxlbhBoetW/7KoseDip/CzYtqkTMItVNZliUxYNQTu9YFQmSEZVq0eUYgZ23Ayk632Tdmqs
Is6zvRgiYztbCBhRoqjKpv5zilwxH3fljGtDBBxo9QYN1nwtIBBnS/fTGT7tbcC0+nIgXbFN4/ac
BcgdfqWuQ3X5gnsin6uhq+3p72idzESY+1/NJDObiSodV+bUGiCm5QZkia9dRfreoHqcIr5QBXjB
GGi4fq8l9VnOC5cO9EEAQlYyCJlC3ETNHeNjch++zRdqkqNCDOYmbR9TJ3FD21wPQjBn7L43JTSt
ODMMCiMKYllMXHmTOmkC+xigvsTkqz//0cx8QphAY/7W9Qu8IIvdoXU5k2Ckc9bvGoAvmpigskYq
47P1xfGTm3lZQzsY8qBW5fEY4gNJo4YUk/EbzZLAs4Sl08AGrCJ6CtT1M5iukemLN5g3XPezsesT
zbwcJ9X16ntlg7Xvy3eOpmgSG5a04aqWQFVR5RGLsr5ccyaMFcIa4KEM39JoMwHPgfvc1F03Rlya
VrSOSJGTBMeXlE/kU2oog9nxuW7cQo9zUKS4+LYeCvvFnffZYNMNcMp7v2t40WNjTtwfYLdGqjND
iulwNVBIw7denmaeHrvGwdrwQvnJB7pVMxWvs3JGzqaZIFqWCB4xgw5PS7umyzpDCDBIuZ2eclVT
4oE9z2wWM3BNLn/J5/MM4KcwULfKlpCua3vJMXi+wG+yKG8+YIwvgSgPKKPNsfZ9CnA3iIhUoGff
NTIGXGTGdhcVkYoF5I1SMeiInL0TndO69Yu1IGNuMCXPudUvSsx7YLs44I6yNcd4uv9UHFYBioRG
tzPeRDh7JHOjenXiC5v224HNIql1p6wUOp7WCOPIxtJlzo+bAOeFwW2iQfF3tTBqhyleUMlFhKUX
JuCkO9lAMfKESBtiScaqys3wvqmCiwPofUaIDtq6zVzayIpVnFTeMJTUzg0Hy6l3zxMFTsCe+Wf/
qsc22V48SUZlXo/RpHATBb7Y2Bz6TAFmXH+PEadhf51i2DY/1xcKRiTyK5qOh0kxxo/d7NUszxPt
G2wQ38vMc35YwZAfFJivfNeAS8HwZQCctVr81OKWHJu/cwww9h+bHqldlK4/FHUfBdi3KwDVb1pz
aMsVxO24DKLhxZF+eVx6kzyz/00Li51gSWFEDb3R2xvm1JfzA3htxKR5il6Ezpuzdb9UnKiQ9Tka
yVC1NGHJVlPgqZbnPr7md847oi+yu0Lx9D0HQcYk93OIhjSCadvExw761hCYLKcucFH2O4ssb1NO
I1U8e1ZN1AvQGOC4qqMdhFtqm5XG8SxSTyK++dETFhhGrFFeMuw5yxj0jBgWKcPToI225pCLOQ4Z
PxqlvTMPspWUr3dHhof+oArMq5mQ5cFQw1vMTgvRP1q3Jp+wgSt6YSU0r1X+MB6gbKKHkG/KBul7
UujiYLPZMC1aOlBRoOK/MOwIAqhOSYyAcfoV9cq5jRL0K5FJpvzefk7Zp/IkWVHmyGsgdgSeHxyJ
S8SdE4YySFxivcMCydwrmA/KRtimqXV9A9jtNlfg3jaUvneNli+YVGww1Iu7tECT9NHfaweN0c7M
ILP8rg/cOekIzrBj+crEhuvfpxHRnHdNrEpXJ8ub18ZanQFOex2U6vVzgVd+Ky6vvyBnihvIZH7i
k6y+3E3JnrSmolsikDaGcC2XUlKepe8LbGN/jvTKujyGEfsx37aAq/KaCaTcoVL1nek0HXKmn0yp
aU5xtAkyoTvjys4PtrMisOq9BXA1sr4IKJ+W5Ak6SwVsAloA7IZpbmCRWNM277BBIQM+2JoW8Ss3
k/36ZURQjyvmH4AcqCUdxeOm/CG64SNRYro9grgDppnOSlhkzeqC2uYhECksCrU04es0BudKdGaU
fVNISt7kYj+3MgUbkT19CbR582bNRAqEzQRZTA6LjUvzZtvPLnFhUKubhwfXB0HsjKGyM/1XBF5L
o5zVIlLFfkC9f3E/s4nm7vq4JERCjSr0gkJ5K7d6LTTXRbGC27mRBvu1UNjiUG17y3xG38W5rrHp
Tl3iSTYIntBSnuujVVfv/7sM0NnLSr+7bw3zg8BvyHNeOR2tyLdErquyGII9d3fA0speblCG2y4d
G9dbT6eyDBCkCjk+HOgRMQbuKYqTEjIuSOMSrAiyByrpVviikVCdnPo1DoQuVvzQi3TslPacicoP
5MK1jxsaT+igaCUtpJYa+5bZ1GK8cUlk0Nt+zeQhHxV9IcQSmeUi2ALQ7LoM3RxPe5z04FfIL/xi
OOPViwVevO6yZhw9o/Y7fgXxKGqdrdrm41TY4ylryAfJHLDseq2Kk5BHlwo5hukVSfUMzZoWbGC6
nOT2oN6dBHmPHftXQb5CIUmQHgu01DYBXFWOPoHIIdnOM54rqMGedQYxBawuBCI/XFrWaEFbK4UP
G7NVBlQWqDbGg5ZdGjqPLWkcmiu0mBBuWK9nHIMI+C0Ns8rmQDJwYVLLLXF2WuWtGbIjaNwu/JBS
dFQFY0pIFZc6Su1KyZkyounuGFQ6QMa6+rKQmdkB0Q3PxGS/bVnrajBxWuJ4Xd4i7E+8gP2CipXz
aClh5b9o/TVP83DBvbCXrvP34sos/DGPltRTDwqjke5y/hvcC1L7bIiwBDW1tI395EP4MCAoG8eP
VMoih1XoG/iPszKh4/tyHGJlMr/vBlIzOXl7BBHHX/wO9Cm4087YW/bOgzV9qbIZZ7yhERnCYXsT
4r0EgyBpcDaVkMnWvyKQQ3IfRZyGdq4QZJTNlNTF2hzYOsWz0n1vpCR6YscqHqyxstX54v5q3i55
FNT9x/+u2L7XxLEPh2mz1PP4K6kRS4meykcgbBHq6D9T/6ELoquM6l0EzmCiqpwDdhU6QuYpSiVV
lccp/RpchLtqRGdlx8W2SXXddtwrUevP9pFYfVrlECZLASBc26VfB4IXYgcr4S5AXrlqsTMywiqQ
xVtNzd/1iHayIBLIYOMmPY+72bp8eLzDSzE4c2eiuLTtSmQ0eD4md6X7DH1EUlls4v9jj+uOjz3E
oF6o6oQ9WMPrG/DSk8l06/8wjHHVvS1MGrimqpx5Yj2GylHZeH1wk6lNQrvPejOSyqgunViuesWt
nzZ6uFOkRzJx29lS6emPn2MUTXH40osCFWvQjU4NdLHyLJ5rxbmEbgnQKbwOBQLpJ/wZ9Y8sspWi
hzN3EsOAsUOR4fW6LCXdFf96XDOXYYDy521TVB7uNGC7BHKoQwt0T2AO53qJDNGLB8DT3Y673mFx
WSV87xJ4jrvfgKgaprFE+hySl9Tp6zoxkZYFYPhFk+PXf2d72w7VbaJylF/ZXs2LXHFRzBIt36e8
mJzBld1ST6knx3TVCtKhtAwJCpWijv09rT5nBt1k8bS/Jwn2xxlxaSGS7+ud8AQVACSlDnhSGMmy
F8BD9lBwPxtyFrF6nAZBLF2xZYCJu5kx8qe+tyegpm7JBtHoX/yNHiQxGC7lqh+QdrmMx5fw5dUB
w+5Av7Kx6dOpxicLWPFDg8C5GGmSwh/I1y+io5KNdJYwdgNYtH38wdCTWmTrHsNZKwU74pyITdDJ
ePDLUjXeVbrNxHcA8/8ugSf8DTwYyb7F3m3RzRKnQequfjf/8MvX61XBZc9TV/FC7MmbHu+jp9fB
KxeEU13G3oa/ERCA/7Fbm/pqcuBDJCm1PmerpWQMUl9roJtp26D1oOJq7MnUBHYlxrtrCVRVlj4k
ARkpeiB6+8CvbUfvRHeO/jg5hGDVFel1L2wa8dQLCOEIiIDNwDWYE/HsVSyLjXzUrqbD4adYha4l
Kd1Wtw79RqsxXDAxoEH8k/05tZcn+JFxLbTfyKWMO+dqzIPtNtRk1vLgMvfXkq+DpO4ovi2bt0fc
yLHf8S0S1LHx7qOnZcmSZ2IFJ7m36IzdBDcnajn4qXUDeHDbu3/cnGvJsTKEWUdtfZpD+0RY909i
XTVZ8kxRGxlh8591qjfLP76Wvm1t166d1vxRKQUqLjTWUVEI1qoiciKOULN+6NWfLnWCctsNDOfb
h6VhhbI0tCaPsXEoq2R/NPmlotFxoht7BwR//fYX4MsNi0tjqclNAdjCQJCu3hAV+Gf0lqIYAaWB
J5sXU5spJFfveOUhyAlEuraq9jBDaxnL/BA9SqBD8/+apOdynre3IijJL02RCCSNn/7S+CT5Ptq+
o89tti/PY1Vw317RnGs9rDPnnEH6WK3f4TkPaCTfhPpes2PDz9vfk30+PhFzxA6n7n+pxiK9rvFL
H4l/auKfUWcNFJ7OqE5zEc9ziXPMVQnn7gseupMQXd/mBa4iBO+f9t5wsU3KHLcM1v+uyov/5PLF
AJdva3/QScajgNM8EoTXTMcjxisRIs1DKlfwSoLTf67G4UN8w2NE5EoIwv3e+/sar9GlcQiVi6MS
rx+BYaTDDOFbOZmFJhbCGy6pjp4iVGAoF/feINxFEkZzLGeVHvHwGV5ivrLaQSRTtL1W2MrhRd7Z
s5/02+aMQzryWXzwD4qIEWW0A8qx0mlU8/8+xQsqC5fP8x1F0wQfmp/r4LFlNoYTIF6kMm6XtJnN
WFFBZ3PvCPs1u3ASEAVTSaQaRJZCv7vSk0DHKoyipg5df+B+e9Ll51IzLY2X/m6ZDgg26y/fS8aX
VgoaI0cWrjaerLNU9RvadO/d8t1P7z0wqlhlxKKcCYmZ6bbSo5G2A7NcW7D4hNess/s8CdN+wYGR
ik3Vu7+arbXH2m+uvxTVWCxPV7CopAlEQ1UDhiEOhXxx90P6Ykatjckks40rOJuKw4NCLX5GMh38
uglhzH6CsCX7JkvgTEVUU1TQzmw5xMubfnCE047YJyb42YTSV59Aj3pMVASNI1y3QvZRrqEGPvUs
BMUAwSZ7R53JDVyKAJd9E50I+/0f/n7WGJFtuv3q6yHvRaR5Ji77grO1Uv3blFeVeiL1/h4Xrlve
L6aX7eNk8g9907rOHrOf0xm5R6fj7xXuBnz7PdmyiQnInUcsirb8fPyK6zAtRKGd313PZNBNFQG9
9dav4gmopd73SY8CSThnquOoN5cXMHj0Haz5msypury1SJ0ft5cmXzN8BKXhK5TGbRM0cBGQtqFs
ZsT8OLtkUnEHlEpikCWzLdL1bIADlZoCpomnJ8r9yFP8VSB72TsEOl3kE9ere+Um851MoKb+xapU
4rNxeR9GaOKZ2kX/E5tGtzFh4Ymoq1OtUeoCk1uG0GRxgKLgrXR5N2oGcfjVuDStyFx7jWTivxWw
jNxOZi6v0T1HeL1SfzwF9Ptrw7GlUd60S59csM/pWgvY7YUzuh3cX7hmnI4FiMnfnBeTMuvIsv5g
aTWK7J4L1e3uo5KEbI6ZvfaXS/LhqkvBwKP0IqJMeOqs+YLaNQpSFrAegJ16lYSzgS7iJFKgSSNd
JrZi6d2p4nE8Lhmh0eD0HSQ6F+r2Ws8VB2JdRNeB6czrup3TKop2S9cAtAUsLZI5SM+p/1t51Tc/
2G/x+fSygyXELpsmBOObYuE313q3yh1F81OD05bSerlvxiRvRpS+Zr3hjdR9Dp5rOBC6DOUab9J/
7n8d6n6rBU6jNHnKgxe17s88syygR00C9B/AtJVg4/1grBX2sp19mj2w4nKGZYwcwbqg7dtP7fe0
RXVUGoOuuFMKl4C3yZoOlAgY4KnGLAAt+M3e40vGd5VS6SesxWV1M2A8mezuMWBip8wtN7fnDlFV
oJ/Namqvhukau9s5giacrUmeMirhz7VQaQ4Gj5Ap/Wn/WtLEi1FDdOYTA6eSB3zLFeFtA/iXJyGV
2HJi1/CScKRdR71/L7wF1Rw+z8BCMsQ8su/UEZ5yF9Fiv+qCJAh82bt34adFLPshNtVlMXKAYRFB
4FRRjWdH96k4kF+jtF8vqD0C0NzZycepCjIAlPQNQezL8GQHVQrQTZKsvc0mxO9DaI88QtPbWjRl
Fy7WER6QlQmlySwN9XXStzBj8vqJSlfW8+w3ZQZT4MldkRiGbfAaR2Gbx+6c2vCMRYC1PwFyXeT5
dPvZ2Itp/vmaC1dPyRQ+b83xrZGOsMi3aPpgX6YDEduY7dw2HRLFpK/Bj2kAjJQwP/NbuvU34bwR
SN8e5cGEY1Nh5J7sX3MHSF34M32JcOvc/BxeLyoRcPDptaVtc0KlAg8XBbXf3bJW0krBZ63EHZNz
peYuQybEuYW6J+og3kHye4RWUkvls2WMkTlFFTUdDT/TZSibEcn8AfXoFVdOvrO7jZ0PeyjFtdij
YV8k2tLr9/aXGj19UVHZAcKUxZkRsz+cLkLcW5USxVqx/0/HfyHu3CDT77d3O+INcXw5kTDaXC+C
7YIvfQwSyX/E6HZ6i3mNK8pc48g0Ew+H7VVklNzyRzE1jH9VCpQ9U8xap3XMY6WxUOHyaYI6Gpd7
BCAtSm0UOt+CtStaqU6E/9kFGQvoWjnvurKNhulbLknc9EGiPJYj0qdcicAbfzKhusTTGDefB1Cl
wpI66yh2hToMqPyxoiZ9xDZpKSGACWrx0dzMg1t+ieXBDFHHe2OGYJaNlJaO278bSq+1AF28LY9a
MuXG9OanYtTUIZqLBbd8OwZkH4HKTn1YKu7J59t71+iba/GwYHTBVF9lZKEX/XyCpdkKSjDws92o
SXaoZuc/EScE7PrbZPFs0YXK72kdf7TkXNbttr02z8ZvLE01UxG2A5150Io17KA2vAx8eiGi0kl8
qaraObwdDVJJQ5zt/bVgjJrO7R+yCd7Ag0OPm+jY+QlAIGLeO41GbtGm7ghuH4LFqOS8I/RssIGc
IS5BpALLK3nuxAQoQWCChaV3ise+MC/ynax17U12KExebqskvULbd4JV2Xg4RTzF39V2bbv9wfu4
BhON1Wf6atEM5V/YSHOJ0M9M5drvwf1Z444y1Dx5SP2/7wMY8iTxYVQYxjgokbVY50dWKRa9o6ef
o2LiWOtY0WUGeOHBYpZ9Lb/nqDP/0xDAyDxLT0eJtLd95T7UB2kqN0cR0Rsq7XINifyLcVD76HOf
RVQCoV9IOoFsOj4HiZ14zbcJ922+5UF/CK4x1yjp20WQZugsdH2GDmbfGnAFZewQxF1BPKkLJAbu
L4Nm3YKs/0aSkXakN4OAkgGK2kazNEswvTdV+eftZ3eHTEgsAuR/JfIFakPVGiZ7EQafJheblbA+
N42InV4DvzzIPqnAJeih0CkJ3/w1YBvBJKqxFGO9cvnUucW3QpD5XWyBPGT61Fqu5n6e/PbkloAb
WDcPiYOR+naggpLdgQBi8180TNDvzBlr2dNpGlYcOwBXgOYOlZ6iKN9gE91EhgHNwAqsOR1BxFOf
4aXmpe+kPfzV1qiqL2SxgzDyx5wG22yFJMZ8N/NG4xEjI0zur+g72Au7/TM6O02Wj14Ng1Ys+XI1
7t8dIXRLmcUG7sWrFZIvQ8lVCIKl32knAH3FwxIESrgsVJeRhQL7wbD8keUWbPbq8IiYFDHoju5Q
RxBxzIFZnv0DwKF6b7Ef1z8eG/ctnoejR8ikwmX7Vi7TbW/xU9zeEf5LNn0HMnL4lgfU4Ofxgqa4
bhPpRceSwTC8XXY7wTcu4ntJW+StUClloPT4CbAzuxJQgt3OvoyNh7KpRRrfKnXHShxNciPV1LLq
2WrPi17HZ7mMQfroqiHytDVFYRal5U3Y6GesmPORh4LzOUzkQ5ok7zK59YoG7D5McvNwJ4oDBjdv
UJBj4kRaeloqWydCMXomAG3kt7GMuIkyUAW32UM9WFwvM5uhAZLC1PhjL74H7oj+8HadqpNSVgEG
ANdcJEEjJDU9Hny4Q6ulDxlAu6SoabtnsvsLnuCzC15VTbJ1CsJBbRWvx19GmApYnnzh6w/0BXLQ
UYM6gwklrgWUC4gsbEgcC2/L1eKM7EY3UgHCVDukC5m6PqHyQVCux3MmeQwSOM3nAYFLUmvmI+Nh
jHfX7+IoIy4Ocu6rY7zfo21o/uZQhFc74cJTeDmpWgFv0j2tdilxNs3tdJTLbvMxVqfQqfaz0kLn
s+BrEyQrfF/HV/EMrCfwcp9xF1T2j0ZlEZaosN87zuBUiY3uz5Agr+KA2E+SOiw5O2Rd/Sq3modu
22xgP7d7oko7Bj8+LjL4iLjTCovo6pPSbRK18D8Z3+vG+VBS/pjy7BdDftGmOQcdNKGXI1athV8S
/X1/Mb6IKIiIxKnROXtkYSGSCA38VzViynAG++8R4rE81sLdKNQIo7YywV9K6t3faY5MzTR8Blxu
Qp8VSYEv5C0fJZgnxGows6lJfASSKhkxcxmy1dxWmDKJeXvc6kjYgDe4wBYLqtGARYUJscvjhaAi
C2plabcgOphH+hJGM3mmNZUbpqJhAyFOPV6Tde95xtDC+DecJPEATikvbLOwG0k5fpzgk9+IsdYd
CJT36qEDXRMtdfXMMEQ3MALbUDcVkPGacRsv1DDYu3o39WC18BtzRyxT/h9AoJT01M7ZSRiorHYa
EF2MROqmSwH+uDizwznOjh98PqfT/IpsGOdD5a1Z8m5vf2q8EZMjW2xqeZCp//osjZlElQTFvCma
enm/HjencP/gTg5GlRZ16FaoCsLVWkB98H5rxdxS5A0cAPeN8GdRkvhbOX/NyH0jKdl/TF5D6egp
FlE9g1MeJuSRLU5hRUZOhdDgIsiUWfPjU6SaVwVuGxsNAwaT52UB+iJKT9rPJXhpUScNQqobbAT1
XHBeU5Q8BF3BLxMMRyJhIxqB4iBgLuNLTvjmmX+MuTmRz0pG9GeE2wxKtLT1WD6eHq5Hz359qVAg
eZl5DpU3SPyDoqM+/PC2eDpp2wCPgn+55Jg8vajFD+CZmxLyh0gDw+nMjTwXfQMJdkKmSj/FvX6U
73OXyyURJa/njSF7lEQKjoG9BM7O7DH+cyujcwDTXXORpvgqQu0Vw9pLrvVgmjlbJ2bs8z6FZeTm
YR2M075NIJ0psvyKjGaps7YKmrFPZH8gCGVYUUvDveC1DAre0kAFOvcEdcsqRHI3FcghLBF1jnT8
n1rfGvsdcEddQHd0OKVhWHsSAKdAb0K8H8sRjWq55cyx4wZguUMrpUBV38Okz63ok/VfK8zxFd0F
0SpVtaLfYq1AnoXaKYnzAaDwTNnOOZBG+MMPpopMYu7M1oRLVRFCIDvsHlFzHr04xwTFiCtjjmef
EG6+6Ujeqx8atwdDQ2GYMhWIvyAR5gWg/JvGJiHxEUmugEvu8wpbStfxvqndHtExQx5/YtCyKGPh
heeCKNIoOlE+2B1nd3Z3OPK59j/uPtFX4zRaxjB5Wo4dn1OUQwk5geGiP628dGG35ueMPGRJdYRn
CjrxsqJu0OjfYMDwlwhLkrWVbttQhcm/lN+VjVuH7JHYsjHRSrafotEh+yDs0DKFJkTGMPc6EhUX
aOSrGXKr0SBHw6UmmVJgNJjyTbHiCrrSg3h7NrGNedHTqdHl536KLZHrx5p1DeLxppLMlQ6GuQQj
Rp7E+I7taoq7hqb7jrHuB5bT/ufCZigAfdn/Fovwym0P9RwfA5HyUzzok6E7hqynl03nPmLgKVdo
KjGBcMY9iwMmVjejR3xHIDdjDy97Z8Cwupt2ieJ6SYXsbWvo8LoGs+zYa3fPCGo18hYhz3Qm17P0
GR+c1+QvlQ7e/OVfc/003VN2G+FnAYiCbRN5k04zL6nsjlJUJkiFSFp5H7sF7ObjymjrmwEe+eYM
m9NolSxgWQOE83GHP0Vmc7qG/jexOSGLQgJBY4uQqoN8/cjzS54i4CHayl4686kZM8NhcR7z727Y
jZCsQixahcNaa8Zv3lojrD0ek5s0tTXo9VrPZwcJngabMAI0VxoY4bv8drJK5u/351ODPnPaImJ5
mH67lOc5/EZ69XuFGBmtqkac/xsFvqVL5EN4w4tuHpkcQf5ENlMo6voUveo9rAh8NRiQyo/G/v9D
DHs4V4vS5qNVGWxL9mZjW3DLx/ROCzt8x7g4caPgiN0pQaPjL1yOm2hDgpVEgGsFK5VfEDvFE+K6
w0Wtevr2kL+aoz07FUKhHGt1gFOjCzis7m08Q1fZ5v2i9Fb6BBeTg6FiBFqOKooDbL8F36rWEcHq
4I42Pu4AXMFUNo+tvW6md9G83P4Qm/41uQysGEmCXyGkricU8CLz8YI+iXqnLRMvKAowipmDyejq
kevOMi0HiyVMf+VNyL24it2q3s199GW+n3bsRt7HPr3CR1QXXDxBMPr+XkLbbNomZnNndjCwLqbW
z5jsKRHVuS9wuOpj0r91k/Vme30swfWIkHcc+yBrOUv15VGFnk6Ed2zP8oy8nFEHBgWAfisagL+z
dHG/FlewMQ4dV50y5msmaemtwwvUMZYuKI8TcjJolO17Zjf5Z3n1y1SuLbua/t+XUNgk1HchDWm/
loUAlPQz+4QUpPC7/Z9jwrq+tNpEfjno5ca5LW8EwG3JJLiQWIUYDUPJQ4lsg9U501Yrokpn5HYr
0pQvNyzTuiAg09oXBwBsSrjstmbwJiO961C+z0J9cPiMjQ1AldiM9U33p1hRNNEVoMDkFANM7Tnf
kEUDohgW0FRdLgp5ysq7QwDMloEIt7+gRKOFXaLHp5a00sBKZaqv5vhrQwghlxF0EG5R8nMd9dQW
YMYmXIyhleePxwSNiUqvtrDHsHAStXRkOfjeZr0KC5p/6GA5gxXMTzBDwXfJa/YvjnznXkBWisWH
Wqm1XadCulbFn/Y239pnVQZppoKekVDIopsKnrIBR9jgdhaAZ4zum8wHJVzC5frJh95i5MgjyJNy
ErAUPN+SM0Ef379bb0wGNwQ0ioBkirjjdc5lEtOj9r8/RWLeG0Mwk52QsCE2DC9s1RrYCRoKhk6P
rlcWid7o9PvquTa3Sv4LNbeGlKrqf32/U4n4pcozW4AELnjCCFJpWRqFap12yYWlteZKguGxrWdR
c5GxgbTLJe3j+nFavb0XpHw8YWi8J4Z6g0NmesHlelOlJFfa9MSaAHgEvpG3SpbMfToX82SSn9YB
H+aPEJJ7jxc7+ZofvOSqlLHeRiykDfkIqrPBhOmPneLDyKavJZq5jWkODvoodIYyBd1Zntz766qn
/EmNkess80xwfeUwmvDAv7SfOZ7oFxsYD3cLyUFCmBWCVeQd/L3Kw7LsP3mf3sNCmECy909y570y
cZz3JHxQ9H6RNTWeYPBKGKJtrSt41IcJFkBs2wXv/gDYkzYOdrnRaFxZb9kzgTvUOp6fy9ZRy+kr
L/RbM/1KU4Uga2nbHyKCWxOaDqLQ7T6DxN0oLn6y+jkLOJgRngShHsP09h8cm+NfzsuRIpQwnTVi
cVikRIgH30w2sd4VS3YhJKvDJlDHn4VaNON9g3ReZF2INXU99R39qPdwGO3NYTOggpmdaY4nTBPe
TKjTeNtae7tT9MrJWbq4lyLIbT5qjopMEYuYrwZZF8LmR1S3GGx4TLust8+Q8fmQiiT0KR0TxAlF
Po9lQKnl4+xHJ2ynQ0RzwKfmAJWYUD7+i+HEBY95V3EkRW2Gn4BPzn2Gpvx5IGlFT+LaVPMdVKi/
AMM9d/f9s54YTNwjQSZ7hIVUiFxX2LQ9kc8sUgfN8icTEG0ILGN/RVT1GbHOrPqvG0BJcjpMPAf0
v7AUrjmsqqt+krqRjcr3SY4qFkgy0ZY6KCKtnbZY+Z3F/Ew+totRDKqJ2qp5pjx7vPh7MnhvjgSp
WsK8GUPqH55RHXIYRaw0BhuNUX3dcU6ee1taO3Xp6etmES+BTGejUt8ZRbrUjUOJaLCoQbOoNx/A
PexhzR9zhqVvRYXQyoLyrcPmFadMU39HRNFaBfB5fAY6BOF61PaIOi/BKjoBtqNx9r3KP+4VHnB0
YVFD6IIv288aitSGVRs8e3wZgi/mBhpTXsKwKI6XH/gG/ioiPsW731BB0AxvlYTIIQnzWOB9YO9L
1WHq1YTwT6EmFimL7wNohmaAhgFfhit8080f7HO4eKAt4FkKjEe9HlsOKPBlKlRLSe0TeoLyNGYC
e8Ged4l4mpTDhg4tFsV+d7eFtghC61SYyAxex0gAxwJEN7JiF+Pe1yqYWjRNsLsCTG3Pysm39F+6
ZRCo+Gfu0+xwB/PEsgGcoi9lM13Ac8t2DjW1PLSnYdqbGnwv2Eq8ciZj5lxidLAuhDkreXbWKK75
7E2qUwD61WTolLrYBYJNtMMwn/CB23w1rWexhfxLxoHZW1aOS+5OHAblWZ0XZ49tAFQi4qzZg3v8
ooP1H0AVWulndYCHorUeHZ+xhIokCQKT13r6ZowRciyo3QKfoFMhQSCHezoWrs8sr5yJMs548ezv
VIp4QGmC40DOciKYTkwh9AggIyuOsXGOzIG2KpHN0nOnPOdJOqfpuiSJ3326zbNsJE+OvIt5fGW+
EWHCymIGGW1FxXRg0qXQFwjyOhcWsyUHWjLqHFn1tFu/uQVNAw0B4tz2NzyI9trn+tnazTCJ/w+c
sLcg1ebKfTSwoFWsbphn0TvfpBM46CrNXqPWVg9jGb7WfZzMkohhqVpDGkb/8L5U/NqYeRrlTaGu
P/EUbXWkCJe098Rv4ZAlR8S1Uvj7u3Sh9C5hBJc+NqqQq/JwMvA/bpPO9pFEzjIRyTr78NHynOdx
bNhEyDR1EXi0Sch/9NL7EaVT8T9iVLqXxDVOJ6OF6ZjYwqJIVreRoEoTbv7xMoVEg1w38qw0MY8C
y3mojTXnMaT2/DyCDhQfCpZPOBbVgHKUCV5Ckhul4GzCQgDa4nY3P5aVNAZM0Pcd1/rVaMFgrKGD
NJ4LlhQijdCzhwTVYClZFVywfpkN80z+PqmsCQrH9EoKhFrw9KYq39Kwpb/l6BbX7+zdTE3y5Qzr
HNr8w4fDePaCO+355P7owr0N31jO18npg4I0kLE2vIEhII6k/sxZ8B4mTL0iPeWJ83oJAn/r+nvD
AAlDHHLq4hxwPW/CwuYJbHq1Hol3EceWlG6TxFbwY330F3UoUvkUy3zqB45yHRcNEN8W/4gdz5BY
dgRPMrU+zLdzRisV1yJyKmRaekm7ATF0vZPUB/hHVMMrChVA9kXC49aBlr1LqgqYCLhSOIOgfTL2
fcFout537hEpTKbsczW77BDyC16W7ENMoW2yr0vb6z2BYI161vb1UpQ/NN0Lvd5h+J7VZ6/MBypL
INzvCRdTN2xlZebpx8QN7JiTt22LJBFsAVk9PjU2hRLiBU0nWP8WdBr815U5okZT726VaLUQre5b
UR32YBD7LMsSUgpdHaN/hOVpbT6UxZYHGlGfY/k1oZgF7oUuGpkWLJJO44v2VcqbU/pbtkclsH02
cbHbkLSK2lpFqgAaIcwN4veJf9lEKIeUkSBnQ7XXtvAsKTm5Ly+Q69DFGKZ2kBWPTtND+TYPagRF
IOLTfUW+D3LnR2Xzu0yc2UTTrVvz67NZS9KRwhKojcvAs6BjuWkPsFLGpptle2pbAM1sEPX3Hop0
QE+pEkw7bFcAMtaU0EGDd22M02jJHolM+UL+kbaS8hK7xk5dmw7g0+FBWNAFCgrvcxhuMfKHYkgJ
XFJNlj7bRyJGiNQnj+mToDdj2ApKR0q7XZB1eJyS8rjUm35zoZG0gRncpkVaav2P1eTaJPfidMeI
ITg6I/3fBmZVYHzbsPJWKsRcmBYOjmyspvl6E9TgooqBdrfHUBjeNxiuhQFFwKHdA4aMubvs36Sk
9OgJ3o+vtWqKl5C3t0W9lYMyv9ZTpd3JEUTYOpg02oH91SBu1F6RTDwXdRhcpqgckq7WClwfDYzo
c+dc58SvnQGF4LeQTd3WDp3M6JdOnbmfhRF1Mv2iNlm5BZKRn3zLqG8cBhPQKuaLnSQqmBVAJWJN
eQ/eEB4OMO49+lfgiOA6yP5CSbjaOc76ZvTZYHQREjAH2xxMPhFyWQOo+ZG2ChHNc7ZF+bgcjqSy
uFMKJQE9S1VncrjHnA+rhncknbmRA91q0nQGugEWjpf80d7wF/NfG54hNHA3OzDMEA5x+3ujt6nq
75wuxu5XDnFyzKTpYsBTdmXD8Qat4Yp6q4bol6STcJMVxocA6Q5Bv1rU9EZaqyeFJrMcJ14fRfad
RzR5w7oESHWrn6pEBof1+gF+OTVm+p3hpBjmQLJ+VuTZeBmUXagDACyZBSbvQCmOicx56ZQIBMC+
ys58+OUdRnG9/Wy1XyiJZnHdRzhpI29e0KNEPJ7MlKN/g32RsOfPiushzKLo3s2TLlfmgw/NFTmX
UCcU1bx+CygFD3GNc5bdDXka9AGVoM7kIUGwkt5JrF5PpNuzCnvdmFiPprKHcPP6bO/OGkorA2O7
I8Yl5QUDefMDzByNUhGMDkfuM/E4UDhK3CYCUGW5FsIMFUn09LfgwxwDQ65tCQL9bP+ETNLl1kE7
BQYv2j6gWd9z6apze/JzYTHpGmGuc7+jeE4vsQzGcXRiy6ttXQCFlrn22MSHpTbItWwVm91csQ3x
YkuyCgrsE2n9cr4s0NYPzPvh7BJgYODOqeNWnek2+cMExR3alY1FceFA1RWd0MB9BVdBq0Ox1JM7
wJqliyynB7YjZGNLojHNErtpmh0g8V0UcEvQDtnlxke3nxVjTGr5EgDAAjYw9sBPcBBiMseI9s8D
AOcDbxEaBF5PmKbi7AyhBro7mSqWlRIztwb/mDWF59137VCVA2nNEQFFu6PYtI5zLb8TmBiXwiLd
vgJ1DdgziKiIEfWNB01+ImBZwlnu9PfBKW88SVwAKEleoOn1zgR4eDuFbn0Ngokw3zDUvO/BFSXp
fbh05uEOtmlYo2RN5on5wqXlb6YlsdJ+TYrqjMJtRz/pZ47dn1oommjT4YH74DLXzZtPI9l7gbLP
IUSnF2ChUNkd1jU+PPKxi/gugYYcd1Pq8bPE3awvjbH2yjGEb/SGoJaaJgojLPlWNGdq/OBUdNYl
uP9vpaNZvzaljXa1Tr8SQ3etZ5ZHvMQHRllVv4nglaNZ8FpEvnca6kw0CPVe3uErCBV/BSJd0Foo
fajqa5VRA9aTG/ILN1BSZN8eA7Xi1vo00CLNnL1LfB7oLg9UEaBtuEfmzkxT1dBcwnDJ3M7PB79g
U9NCh332iulvB2QKE1QaW0iXfkHQRQ37iPvDq0DARjVbpufzzOmt9U/E1xKoT1g/hpZ3jVGqMhgX
+vtNyjZOXx5LV1dkXVtFI4IHW/MAeIxOICKIZarLWxM82a8xuf+SneVQGjcBDCACppj8ku1ubZxr
JkuKa4uvasdzaqJIPh0v/haIeG7CcPE0T9HgLY8qyOtJML54AHQvTKGOzWKHivjktAk135XW84T3
zKsEFWDwkhmsjTZLoeyIwAx0YI02z5YVcQqAf6aEEyHZ2IGmHoQaHgCrc7V1PKkyh3Vuurax83n3
8qH4ctePnIur+PMIRcSwLSGhjLLef3DwuqeGZf+HQVRTbgXBWf58+WGT51l4BTsDWrTRJEG941eF
ZbxDaxFjdXdrlabreUlHYf7bWXjHkJK3liJohSz8ipPseOeF5zM3qKgSOAl4UFlGF6it5a0WtR+f
CwFtxNpEyCVqdmbU/vPSBkpq3n3RJXlbagqgqh72yl4GtY0EQQFcaD1nhnXdxDyTQ3tPg1W6a7Rt
L8oCEGCgW/tVQJrfOme5Rr3r+hZrULo4ONtDDC3eLw1I4XMqc02lh4oJCpvfb/6X+d/DXarlATuh
rfMXzw6jqynIAShndV327CfvAeO7AdRe1FNJ1REt6YWjgpuOLd/yCf9w9YZw2ip7uH/+448ofrda
Agms13jkyak00cFCyd6f/5FbqvFCl8PO2FcG0BdaJAR/ZT6K9is2MLVNjHC9kKNRNiwhJSKbYjfe
xqzEiHiTQrhALbUpL5ICS2jWcQz2VKOuDZHGW0Wb5Wgx8BUNDVqrchsfPlci0JAnrYTGBYpFd1Ad
gufHC92grhGnUohpJuepIp+o65VmcvYqxISntB+q5PFBtyKxySl1/J5amU5R3azJbqiQubEhE3dR
iMe06YMyBlFvntq3AueqeMao0cTWpoKmiXTK+Q0Ja/1bzv46NcHChzXF4UdXCwqD/aLy9bVDxKZH
Ro4YIIBV1H51G43T8UXfGhqBqXW3NsBcR0H1+L/un+Z/8jmYIOZ5iuX1j8OsH6R5BgRBqLCk4F1e
AsePYsiXlMPel7fg8wX/reWbeMGSsvRHR6An9Xl1wv+g0X76zHC4MntoSxnwIkE84DLlxOixwKO5
uMjfBVyCpZW9MGaPepaGPGWXyTkhDESQ7skb19ZynitW4E1VKvEilXZPnLuQHIxN9HjKwE0x5dxY
Nj+2ATJ4I0RzGfzaVGGLk8MRhxdtGy1HzYhFprlFsdPXOAaVJcwCrQEjyHt6I15g/eJSRRB7YAfT
z8tzMSMYIRk4InpwgzaY6+ZtMf2H/6q8u03mrobEsCWE3/bYq72Z4CPwsduJm5DVVQ3XIW+NywIT
HmpGQ7mQDP0SL9b6U9SwCn3Jqc60vwyY/exVQjfeIFZXDtgKW4e8/hvXfHII0IW/xig56Dk0UHUH
QvCgkWUShIrK5kLBuWG54DSPIqZrJV1iD59VluSsq8WmTnZF5u7GwBdhnL9tuvupmUYqFrnFaZTD
ZJHo27La+xYdKBGyhtHJolc1v215DdGOb5iis5+0NfbclbOr4Pn5Ytd3yFYm8AAjQUo/4CfQTUio
8xdRod9AqfHM2IbvsKFMkm0FhqPdEwso6AkTZx0qXN1rLNAzxUZxmBVXTRHLvdh8DYhIjk4yc1G3
ovG+rYC9tY9LK7MdaLXRa2tMSlnyw3o1yUOqSIg6y3sGoh8mdL2vsHb5PH1k1ca4Lv4lE9VmeXXk
rMlKR54qt5qhZc6H5iQZxQz6UMV7C5Uk2yCwoYkWewFGV/GBIqvlGxt4SpRrCdFo6XppGOqfVaoQ
1GcmBxqN+aJ6pNqQFiifqxkA6qDb/krVJbRetdwDYdW/p1/139ysXM6kjkihxtqlYL863ijsuT6x
LbceL5e+tQNOvT3v+Ym98SS6xUiOK0Mg90swsVuN6dDPGaVwy4M5k+s9/Gjw4Qxiw9XaqppNOxUs
rezaRPcLHBR+KVuMNraydq1LZDdtDU9I38duzFgTvn8ZoUF3d1/FlFWDBY5IFQ4CO0rKt5dXbSyU
nFrtouQOMBiDEr+IYJLIUNVy4rhsAdWRFiZaccXeF/1PDPRYzkQ8/dyxmiyRDh5qaK8AD/kz3+b0
iHdwdRtzLNAW2UhqEr+WhUaLRab2BRbrjdEQRTeuzwt6MNpmoYuY32+QyIDvjpRyAaD/KTI6tLAV
USHhRwYWC27fYojNDconOG6LF+WoRaapPH6l6/fxj24MNdv77765Mbfo5XYd7TjtA0IsOINmMF7i
nnL+D+YImGoaPXRpiT1EBfG5pcJHjTt6j7QdWw5vPFGKm2j8me7/h9cAiiWFpkpN6VLzmi3zHrr2
R3zQUJHAdugtc28YaZcnEP3JrHoqe3aPSUndLNJqwZLGvo8EvwOrZvLhyzoDQKn899CAXfjAEjSn
RPpuo2b6NUGMhvNht7kdFZvxnIBMskjPX9fkAuAlTtrlhx5e0EtegEayAvkxWmEV+zZm1kGemcF8
DTaC+VvvWFl0pv0eolLiTvxPeL4MWyrma3h5kuupELwxTlIvNn4RWDcrlbhslA8zCps3MCGM42yJ
VGhADkj9BRjtKijDMCoZwqChwU4TvXdbkEcG63drDleRmJFb7yHr6xmGyh6KZugLV6SPx5Vrffnd
8cgUKhEwnXADGJruNXiIP1AcnHfPJHS3Gh7wVmxhT8a9yNTjh3Gc9EqIArAbm/N8crkdsTpzA5Px
cM+IGQEpsFD4nbW2L30gSSfP/SEtKJywz5FShRVunZ9uZXU0V++vwIDi+NvK+yxMz9qLng46zgdT
gaRA/0IP+J/SE4Fp6h5K3is+M3gkwYUyHdtjxPIYS6U0mCZad07810XyNL3/r/hbmPt+uhnT4rOx
lkJQ/OUydLmymlf6/c/VEo9MNu9KtoT5Q4IVLe89MMbmzuXIZtvYnDMZMaGRr5q5el0TDe9Mbnpq
27axiQ4oXAxfQWfwRgeQYLjkxAE5xmHz2lkITOMXkSUiCQN2DJTvK7KieGVtfFC14dq+zqSY3VD9
2POUIrab9RA1V6y1MAr6N/jC8c9gBk0n35qJ3urYPRQw9nyZqD8O/v6Tg9irE2I42nne/YnstO1Y
CQV2NvHiwNW+WAWwEZx7Er60sV9u2oOkZJxXCvtsw/8CyUvyk/7ym1HCMhBLhqsdiVldSd29ODnK
wuscgyt0Kuaw1pFo7kKgWYuiyNMy7PW2aaVpumSBbB6g6q5t39oAlf971iBagkEs6kAIEI3cbhUC
hseLCIu+8vNfnVHYjzrjGZVh6B91fCnkzAY9wSQZqPPdIwXvHBDnSoE/ubg8/quK5LjSgmBmB0ck
/CFuU8/Udvy6qrXD7U3gbIoJFtiUQJ4Grx+4loA1AAxjixpyQHhKaYxhN2kN1gYMlMK+xsD0H2nL
RUtC8QtDpB89G0HMRLOriwYHNiszj2AQiRkrtHGMTrCCzXTrEdmKRuClbZ5rZIRJgVeaAvr+B8JU
lMpE4GjUnb6TezXCoc4kc93GV5PISCyXf2NqNJ8RsqHcdGJWtxFHOlUNwQnu/P6eUsfLnNuan182
711gMtvTLaOMESpBdEWKkf1SACu1ggJkJ2glBBFWvTGauFYSdW0q3IB6dReCq9pMphXIPBaQwDY6
GA+SwU8DHC+XcwajWWeFZWrDxQTm5at9PT+pUo0XbMYhTRINcGOXKE8lm8b78A5G3S6JgGYu6HzX
L/yuJfXY7hPYN+BuAjwLXIXcs+FeAQtEjsuaCXJptCDw2Ca/3HBl9AStUyPhUAsAOzfPkyavcJwK
BtqdDgUPwOk9mRVlv5aehOS+rC8fKTlsJhtn5U80tHmC/rQKLd4shNav5pM1uh0wOW6hx4x6X0UA
XWQYOUvDkvjbklcnM1Q+1AklDz3FoSuoFbP6V1NMCLWsC5NujXhQPA9W7NDnfML3qOK4aXikvpiE
V4A+sMHq7qY+bHl0qu3YBaQsK8vofuFtycxnAWgyA9Q1FWRqWJJMB2Gi1B56h/YnyisvBG3Rhqk4
cjkncA39DLZwGA34kbdGrKxx4uwgm780rH0pJSSSwK/j+rf2epHo0aI7dcckkg3HPOXv+WROPhlE
DLNQerYBwbzseumjT9YHBhj8YHMtDnYAFJBtRGhf5lShiwnA+korf6vWDTntqqWAZwyN5xGdidmA
ODnJEs/DS57C4l/zJI47WE7SqzBplAU8/tO7ShffTClupjFzGYN+ryqMO6zZCNDxYLU/y0p6qe37
3vncAZLk90C3V6imlk8bmpcnzJRJIo7lZ4EprIluO5MYcH79xGrR6Ka+cbT4z2RE1iQL/dBkmS6K
wGBxCL8/fonQeFzZSYl+vKvOnTh9nQnpfO0qmCqXmX4k1+HbfZlfa1lwCtSHq3HvAxg5/kOmMiRl
RYyyLmyJygdzhtApCk0WnoPRsvLtFnBrw3nzmmAF1J9mEeO4gcNG+MB1PlsUH9FYrPHFMn8cgprr
Rsk9lQrlv2fF5wL5sjRlZr42z2CpCc2PaesGOcpXsMvLhgrLAsRA+jBeebW5RDEoAZGdxBe1TVW8
suX1rEJQ57bzufmIHaIKSpXGu3ZUXwfC4mxIRvIY7dR2ar5oK1n6E3HCM2OG3Bau2ppztpCtA1kr
iH2vtj8EjV6hFZ6jRHUPhPVTt8x9Ckvjh/yJQbjhAtnYGDcVWIkV2B4Iha4UoqeCydzaiZSL4KVU
y9XIn5q8q8XBGpPxrMfydhKKVulenf/baWkwvHughmvaCH91WTXkjG+5GQJnZA46LiVhVSN/677b
G+A5ad/XzovvTU2vUNrNhhvqHRIiJgckEUwHDrAIUbuSzzVvqsxBXpxtP8CjjxkoF6TeUXTeDr7z
5fFyRMjd0nvIH0E9Cwlts5ddHcKrThVmAK6zo1ogUJVZuf0RXoUi+l5hSyAHZVFAXxtXNHNXA8ft
fYMFOXBMocsF/dP3y2NR/I6CwbQEGKqNLmExCrj1zDqwj9VtU99EbdGhxoYEDpD1zB2G0jXrCNlz
ya9JqcIeaaHFFskprl6qdMxM5cZeiUzai2o1SI8Zp8y7voF2GmyaVhP8zd0AdlpBNbgU8g9pgncG
rQwWlPl6Hk5N9uH4V87ABe31v1vPaqXCdzmPqDUV6HAokKlV6r+jikQknilvsClxL8I4dtOjRFFl
xSUTx2o0YJQj1AjnUym7cp5/aA5IZmOz2/G1+Uh1lNgaWjkMGgNej0+CfByDmHXZ/+7ltXFOOt8l
PQvTQB4nEM2y4r2SzZWOyqjypdiNAlLOwdGHUKgtB5qa3Px/Hgls1JxeZmEHtO7AzLwFqaJROzoN
XWCBijwv2+lQhqDka/+4yZCAXqZjtyW0EwWzb3zp1tVeW2cbi2jkctzAN+NxaEVMwQACwR10YkNR
FFdYXTLoHbL9l12RDpkh4zRk9IzCz1rNVE2kxUtH46zJ04U9azAmbe4Ahu9metaE7vM7udoDaZaC
5GvIyHSQ1sqFKJKGxYQu8XiO8Cw4Kt/Ey20W0PRaor3fQc6lXHzS7cy43KVTrLyFeWdqg0r0C/HZ
dM+VRgBMlVqvJIDgtQ5kptljAq7CG5jlVuNA3OfvIr+WOWaw8wSFHaL9EZeh9Cdyluuf1C4Cbqgy
diALnQqVbZWo/PVxbgSubJq/gY3yYL0/TpB5Kbokx0j5dCpKv3PNdUeFHIE0px7e0SxRnEpQFUAh
kfX26zrZBwjE0B0A74T/DCnJFQc/OUd+xQTKg0Yr5aqrIQ08fPFzQWTR5sxq8YAyO1bEX+TXNOPX
ZrG5gBj52cqck21LgC5/nZfwGK+VDLaMIhbNsdtov4zPFUhWmxOcU7iPGvQCmLRqB3wZ2B0f6I7r
8qwWGqBWR6k4DGAC8rNI0GkviBUnX05k2uLCm8KmiyL2kFRmXt0Xh9AlkBj0x9xnVo4CPGXox6Q4
Dec9vLNbWc5bULApDJ+vRqLxHbS9u4HRbJLEZ7FdHrJX6o7tvJXTiP9eC0Xl0Ql0EYy8RQKfFG3d
gYBshub+kBMBeWezRhNEp1xWyNH90l4R82R3tyrhKEhya7mf5Q90irSsjAUi/ZNHUjARuzJ3dhrG
6TS7pddLnPTQKf8ydi19biKJbA28zx2lsHWRXWrkv2wfqeGZ7/OJjD/+Bz2fW9aUf++LJwq0e6ux
WiVhAJoyAO8hp58/mtx0a9aTkC4YtEpPBpTryXPUgUHoCzh8z/x/TXjHQo7pEW0eyiSl22svqMTE
lbtxm0aOgkTvMEIHdjqqGsuwVDO3FbngP/tQzZdS/b5BTykjGJp7kgmQkIT4Cm3OJmhGqb59FiUb
b1P6tCTVe2FS+1sdisGrOJ4Kt4YXPyH/PIVkxZJCQw8/qcRInRsxM+ltVO6tjCE5JcTo+ZPRa7AP
qrLtvzLusaRjDa9BO17gv0fLt29vXWnLIUarmlkLWdTi24g01GSmQ2Sihgml2pxQis0wk3HTFOEe
zYOZbMBI7OxMbZk3tmWpFBQsgA9SC5FaZItLHboeCABJhkfYCzrcP/NxuV/qMUhgm9fEcqR2O3V2
LBVRpSZyQx8IleYWlYFbJoOGXcVPre0+LoAYnFHChWR18uYUB9kQYSEEi5qC7Zg/TPBi5boYbGGI
3yMrDFNeJFaL9GVPCScWeCYoyXrUOupIdKwbrFquGABb0PunhmOQ8kKxuYC5yuFiPh1unk5dVvuM
ib/6C4HcMlpYwzWgWhLsAWA62ZYZtqu5DRj/HFyDDy4ja2d1Do11jPg04d9PqN/IUBxoxcVLJ8Rs
3QO5IV5WoXats8XJmjana+gGRJtMgdRnS7rr/MxNW4ixx+ywuujjgOe7uUEaLPRm1xMsk0J9pZPu
gaBDNpBK2WmidDm6WS368HfqudvFi/T6GkbkQDZ9K4Yv6xHK9DLWv7sxfIQuJSlxRwWnc36AqIbK
4ORs42e0nDklkkcW025kTzDfKmcDM+4frWzzpxX7WMLIexZUIsT3qGC1XgKxAVCuVpCUF4fCjsDh
9Vc/3G/69NEXeV/a7q8Rv4TkX8MP4wYjZ2k+EQAcjFB7M2mXLoySIBCCeiHRx5SEdR01NVmpHmjD
ny4/22ie7WOt7rWerYLYU7klycbA2aMA0hFxeuhZ35jKZ+MvNCAd2o+WPSxFFewXZrjyZl6M1LXQ
Lpm+IkBbKR/tDYuljASM1CFtbxTnBLsT4yUJNqDF27irE9Dg6kUhvTpPuLJHEfqoU17J6V4HePEl
vyGoIAzAgqXdLwcOqzTiMluati+WFLohSyDZcMngdhqqjL38SMVWYsyvY6CrIpLB3PCo2+Nbp3Is
jaW6epfW+1Cae39GfD0b6jILt3YglcCaeSj8TWLWLw4R8U+ix716n34tAATdCFlHDzpRBgJygkee
K4oTepeIDqHG8155DjZRnfsYYbHU0X0SvHsA5nzbt5kSCv3V011u15zkHFSyf3pLGGk/A6auKQf4
SR84G4AUW3IGnvFP4bD+yBbjUvkrmaOLR72nJ5ZPcq7X7Tr9dGf3YqQ4eu+jhwvSaEuc4kt+MebH
xVkn1V+Wu+V65js6caALJQOo6Rh/Lkyd5FamTFg02djK8HP5s1w/fDaBvPURatLMIXVT7Pd7iPpp
ao2xVvur8hfNe0fDe3sua919p+ikdZ2pr7H+BwJ2aBvBwuEArcaWKTOX7mGoNl+NQ/g2J8M5clLi
FYQ84sLxsiLaBmW11Y1CavkLStDti+2exgUT+YE0/M7Hbue0m7TcbmjzX04+lpu1VIIp3ezbRaYU
sxVjuegDpYe7wIGEpzivpsYjmYnO9MPraRg4QIK0FCcxprbd7T13gZvRKLMQ8FSxgEpdh2tHD+1c
stp5836koe7nUksNHrgSikzlMZGpvMBhMglssndWhnyxUp44YSahQXk9N9D4nv5K7AyuEFRcyNDh
n5pS2BjhOxvnf/PczdHdWsI3tFcPjNyUt0ro1R61k/KYFPNXKUARJ/zndmIqxSFVQ4nGPFqtB5KA
E7k6hKja/hd/0q4IlIa1MM7UiII4Ule3dbmD7a96AIwZsLQpRJHkG8oVdSKxLZ29ckj/wHZYMsKm
a5WppSYze8Sactq20J05t3K/5NeygfE11EjXIBGq9XOF+Z/4H9bHjUTxFrWl7aDUMv0dYMQ2Gqmy
xz0VSsKJUV9e09xhqsGdpELL5hnuI911He1ONYjJm3acXqeKtVZBcD2SmJS2Ura0+Cy9MUOk3tzQ
uzT4KyZfpKHsdWJBM1InFr2gZ9R5L25EVH86d+4hPA9Jm2rfLGNKOdCKpCrOAUlKb9wCk2e9G0mb
FxSDBU05G5kQtCKok2rXKPprJkjRzmlnJ1SIYXGsN1fR80aOUc8l0MwiAuBjHrlcr5IHOaZda/T3
YCVqOWh+O/eOHKw3ZtzgIO3dzV0YG1QMPr6yDDn1SJX/nQtqv4EZflBTaxHPLZTQeir/9u1/HvPS
Ef1V6LyicJvPxwEEz7RUDyMHi1xV+TSbn/0hRMgI2ikxDcrWjkUbaL2yjJLG65/mO36fz4XEGy1J
XUx37+U33hNPblgWZGISo7as/OX3qA2kxvPQLFtYMRin26UwEdQIAJ/Lvh8nNv7CxRTYh/OEfDin
VRchsu2XOIsj0Q8Nezfu4xy5heMux2gAfJNZm6iWWkBaAxYGAiRGbMIv2BVmKD+JYQxqUicHZVm1
S2s+Z4vI9ita2Tv8GKAk2D/lFU0S/Suxc+vQ0zbr9b079AlGUhHe9teiPuzCEaATJM4xsASNRCYA
NZ039XIIo3AOT8+MrYnG6kefguLZqEOkaljUdTF6AW0qlSMRee/SRE37dKyR7N4MsvMxLVi494wh
bwZS5myZt6AlVCa76WGjxueI9EuFLFglxIkzdE1xesEtqysBX72Dz4KQwhqs1rd287WmJ9qCaaQa
7NuubG5iKDc335KlSJcmoGqSIp/2y5P0GaP7j2kcK940E1ZZddVNe6K+N+J3TMdRYsMGToZOW1pU
bCt9vKm2VTgULdJtx5JBF4yfSFxhYH8/aHCM8MrrhKLQzPlv8lx3kSqkf+HEDJ7i2TF9i0Dx28aB
wwcxpS2EZK3u5tk0zhRHBke+3hfDNmiXU9fbzTJeFrASbpx60+yCHnD5kG2OLXGieBNpdnuka4TT
94Gd0/nDOjP9kElktB/x5/x3Q4RlmS/hbgyrIFvc8ktTA/6l8nXtye+/NLjZVHH4UqPnfvgrRWjH
nnJ78P7eiYlwmGSAI6sZpOqkwt+tQWn4iaiTTWzY8WPL14rgWIOMKnG2B/ETAAnHCpYeLgZlJCBv
brnPOckwE9Oc8qyNq/UOGRNiIIpUQM8c3ytxRYOblWCPAaR00HLoZXhdq6eg4t3xOm/2MDxrdVLT
GJO0OSQ1OI6tXcHDWSRyTAesEn4bE0SpgCqQnxL3//VgOCTMQY5DV4rphI8s+EnvR0aKoxfQbtTx
JrGQi7bLQE4uSRN3dSfxrYmRvORqwdXR+jUdv6IFqrRGagcDPKVlnc7tLr5/iI4tXYy1n7KJEOnz
HWltMCVCnjM6xFYMj2YgDXvMStHTZVFxorTnByOAl7IOX+HUSScJ/NAaRmZaV8AqC/M43aGEYcwh
/WkFXTRSCafQ0cSESdSAmpEXD9oiTlHcp02Br5Awo0IwzcHkJy+s7YUnc+gP5WUmfIwcdxlmePiq
6bQIKkIC+Yam/5BBYkQMiX++PR6/g+o0DCu94AzJpEYjYTceLIObACgSiDC0aWcLUx1UGpFMkugS
sQOtnDfFgjyGO4wtDRXaXWiJ3VqNw8/qsm3iLWWk0ri04svl/rwA7ZYnFK9SNRdF0D+I3QmQ/vNv
5E2crg5QTDPdHcyIXtDCVcbPPDVIR2tkZFlYcymPcKGgXCeFNb081RZOTjHgoMoW183npghfM2/F
xKGy5TMFmn+18eZzP7Eo10gbPmPpvv2y48cxOUlxoLIFQdAzC6moA5/nMnrHe4fM594mG4KE9RAO
k4A7uJnV5lJ45Qo3+24ezDYRhVG3aouABq+1cArKIU8GEql5Lu2mtYKW0kFNxO7vnAb4uUySZCud
tAAOE2xVaT958L4mx4qOmnk1j8lxYNXNyVKmLwGlGP7uQjLdcoteNUkfL3vfji+0RoRXfpTycTDz
DqFk+nhNBcZq7TTVM1uomKjI55V3lMoIFDYDDXl/FlP+i87OCAkI7JZ+0VU8zUx6LHXPEW3w4+3D
4BOpB7oO5AjgQgL6gWgFwgmDB9v8e1abeGnUsRIKlUY0exZuHsptVtRU7tFnt2kFeZY7qeu/GV4i
oSBWal1fRTZhs4WNUvnxCaSXQXjD/nag7Oa8Z239M/KDL+/ZPsmDBi3eitvs2uXV6eT9CyKrVInB
l5zk8ijLaSa+dV++sojRJxyte0eWkegEhNadzWdlVbqfEf3ifAAncOg91wO8gPFeoUBY/J9lkhZb
Qr5L8sjcCUKL8ZS29Vzk/XTBUPSfCYpdAiaGTWQ+QWWO6y60/wsbO8a9PRcgd/fpptU1MflYaO0B
cOGv2jow3iklANrdIRecCCHaNsPw1NzPp5hu4QNIW8JWl7l9L7RU7Sr0Q7npAcsT4jXz3Tna15rW
VdLb0oLHAG27ClkEDHFLuR/1Gzg2QR1Ooyy02Hm1Gmv391B0zgGse66x0UE3lf1AM8T2/hsG0yxW
1nfkFoah0MHOg4QDv19OfKPJiQ1CUnNYXvwujBYnT6AaO5EO6XV+5sgKlpV44WVaIa4cfP5WwXDm
Nrl7Nhz7MAc59d/J5ndiVRTuFRcBgTZvownxxPu2tH5S4YZFwL4swXECz7a+gTY64EhT+4Z8K3Ir
oOS4ecVgLvjcNhRk9Dnt35b5o8oyczmQt2yEeDqXn+u8xfxQZeTmNgXU+RUgxYRJXH8arYfJDN/S
uFbGbFEfUKXkidRdP7bLLs3o+/gjec0seAfO4aumSO2G7uIekYdrS3sWf+gonUTKSZ7qiKvUjDP9
OrlK0G+kcHpdyxF4KZYCyZN1DIS2YXKsV3SDp/kc+RQQX1CFliqrBSvfwB2L+z8LdB5LtVhq7YWP
IEBebbXsSizJBMrOIbGW/NUPY1bAQSfdD8Bamn5CBUxpNUwAu3X/OSZiyBMXfqWj9NJpLyyFRDT0
dWtQezdRzH7di9rlMGuVZY5E6DpM4j/GEFvMR4zRxE0H0sepIO3pMgoPwcjnq+udOEwUUyP3yuH2
mP3rok82bvlW+nkEP7RYIveEL4bWYxMVuqOWNujkb06NzBwDQBMQGGZem4IEIKcx6D1Iv03UHDvB
qOq6SkpM25mexRrz6+KJN4+7BPV7AY8vyBo2AStvX4nh5W8G/lcffDt7FOAXIdamHx+JsoPCnxEb
Q+/uXE8S2rDZSVdcWCkhu7+YorKpSELX0am8I5Rj4fDa6z5XW5O+ThDVc4zVKBPn+Cl/D95HyqpL
w3QpEot80wtxQtQVYE8XaxynhwYfHNwS4qIRfE6gffNEAUZUOB5TEcylYg7zFK3Cx33Nxb+QMy6N
tu5vDehpgoh6DpJ98nrNUyJUVge9pdatlLLJeEMuZjIxlC47hsBGoKXjUV1VwWMNLasSVhvfHJPe
efSx3ZI6JtBHgmwItnzoNkDqg7VUrTArI5KA5Tn/rBrXAxcUR67uAbUuND6l5qDsKEeryPzn1NK/
0KPBFcT8rkUB8VctTx8WsVbGt4gC+V+/TNFVPOtqEi7RK2ObUtaw3PPGxomDUp0KrvrrHgfq2nV5
4CKjy3500JmqZN0w6jZQih9hdENv6hQk81oW8uUy/A6S7ouCohA15C1TvArQOvBT9kHiWptmesV3
zw+a2QiAT+gpnBtEQBO6sww6t7ILIJiqImt1k+sPbxLT40qqBNFcJWq9ok09nzJj8mQFhC8+0+Qa
V12egbkgwaTx2ZC8dnTOpP4WCpHdPKy9hMmm9NjdcyvSOTEL3HlKcB8VopPIN7tYnQYmk1Sicl/X
d2DYe1WorwsFalJEBS0zCRj3dY2OnB6AfcmAIqWQKXh70OfeyA+lp0CFG59/05v71rgZEXGl7bHr
gH2+ONjMDvxUjspJtsEjZR2TB1Rq+6LWLw877a+viM+cpfoSPQZIuCPzsvJpWS4Z9HwavVO/AxIj
QWaD3+1cymiPydR7GPYVZNmyd+I3+eyc/BpU2XvztAYKN7lhbG1F+L+y8URwhvorRSwXAVcIRUeB
O3hPNHuNLkPCMwPgF3HnS/+fiRhQVSYZ7qCMgQvzVmkGcO55zkVlUJBopcIwKdQVyfcj7aIHbx2M
tdbQHiVMaCk8cymQhIIghWFaFh7Q7ET+Gfi4qhl/eJSXkEs4abFrchtr9Vz1G7a6PNxI+cTwGY53
cYgezGz1HQ5lWSmcbRqhUmv1m89t2+/aRiPwuRTVMEXmfY4pgBjVZibkU1JRF/p+H9WtogQS2pD7
REHh2kFaaE84C51YO3TK7il6+l/hGijvPJSvQUNolU9lZ7uH0cYOy8F815qAZrutBtpFrenNRSRA
OrdSRVIPGzmePqdGM7kNpjO8zPje/8elLxxc8blAzvqXk2tBp3PIfkh2qE8eJ98F2WZQXqliWTDN
p06cJEI1rqq60WKPd00LxBv3t5og5H16qw1uaM/uisuKNtIKNv7YeGHnC65bH96HQOklZ4DZj9cf
ZS+mT1uoXIuMqMNvYjsENBIXfx31jcesO20Q1p4SAEoX8kMTJsU8atkmBvleI+odIkXu3M/cMFGt
Hm2jdUmG0859ScF/DBOMWYYrmSRQZfTpGW08Qo1rxN17SJH9wwciXIaWu6SBDIN/toVE0EDlsJH+
NPQ/UAL7SVOQMijxfLEbZ4JSJldSj7VPPdO+MA2eA+BIT7TXHHoQkt47p9VKmL4OlMN9xfIqXGnP
Y+f4OzCp76JYG0Ox+LboX6o4Is41Sn25KlBbqATP2joOvusJnQ25Pd22YbjR95Qk6lvZ8G1P67sD
eoh5eCv3WAKwcK+KlOhoHqBaw6cotrN6U1EwvNJofkFNF6BFqNuI7MfZ/SIN/gBt5xGNPm4wV0DK
rqilAq8cfwxQMC7rR46NFOu2r+kH+NIpPdcEyXrHk71zmNHfBpJF/OFY+qKVeXAjLCQ+Xt4cpUOB
/57OIn3nzw2HVZ+u2vW43H0sjGL2UsyPEU++Q1xhJCculNsVKfQPPBKXqe/XvtxzxlesWxRoNqe0
Oz2vvWpf23/bLSneJiWcy4ND5XDSy8mE9ksujL7M4d/2AYxM/ovO1hfIiwC5f/m/91kg08Qp3Vrw
nrdN2jB57SbgX6FoF1SS1eKUpmOmb+HJA1IP3INPKiwJX9S/oKIvNCfXcBjGmOLvwkbbNmB3N4bh
ciQUHGcShpXNiCfXP7krp0++hC/Nd/EqvyG2gVRC9aig1Q0ox9P6E8xGFCFcOzGnElZhAipTx47K
tyFfJLcGnLBIPRRwAETG+qoN5LOwyKI2ICUdgpsg2xedDLPHJ57wEyVKJ5FWDjmUTfzfF0LitH7K
ZNyNawJAIxx475irAt7NIQjNZcKGEt/UBFmNG33vC13wFktbUlkRRPqNwxIUpLxSOwHAw7+CyGoa
wdkx5KEonpMRERlJpOFSE451jqiS5shthht9J57P+jS3fndIdDBAem6IddUjkSjLcUbnsRkMz9bz
P04LcCmEbXvVMcS6jZBKi8aCOXWiKSR4vaDcHuzaAH0RHRe/Vnz9baB5aQUhB1jPupTdWdHlfDEC
3HQCftoXaPZYnP9PhRFrn6GsIv9614ZJ7uT/jJ3ovkyYMh1xFS6UusrJG8ADFrcXy2/9X5wBB9OO
zbPTBVlqzqmPdLIi7a93Fg6sXj0ph3F+wDJ29fQ52TfEt7F5M5fTk3yv2l3EoAlFngC+CNi0sNFS
kB8UrlBc/KfUzkccIAq7ddD4sOBUSaIMuc9JMqJe2juGf1Ltyv/RQtg/HZ4050Ietc+U+eC2xfOI
MASTnqOMcE3rSS5lM6ugWdQ2tLpIgmKryLTSGza2+oFBjjy5qJ4QlNFy/O7c/KLVg0OCrKQq+xoX
D6I+nkym9wtMwyHN+1pRAinSt0IDo6k0pBq18LRpqXjCn3w8ieoQrWy4+OVOobShTe/7692lMUkr
DpnzitspuXvhjG1/Z7UAvW1MocOTLE16Yn+hSPdcG0oSmDFNeRUNQABOf042+78gcKGsFCcZV3s5
tYpzJBsmdx7g/NblLJhUTREzw+EqV5RUt7BNsEHNg49JbQh3kekmHDTB1Ru4reHERU3hDcDy4S4p
G2EXvZKJHZjmmcTu1rHTuXII/yZ1p7g8Gu05a1Mg4FWtjkJHAI1MCDViV6WY9xw13mlDybpaCqa7
DskW4IaDZLP1336PaycedI2npiHp0E+6YEQlzOvYD+aNrMQfEpHwgocm21hxa+jY5KdYKmRQmDQa
wsxmGMgPmc0DeeCGAKtLhgvq6n0/kFe3guyuMY6X44vM4GRDTPpV2n/M8SDJ23GfjxUBlXu7/ZTy
M/Mn+ehQ3Pmul35c6L+uskl6iT3AW7iqGGgW5jTrqsJZ9I6XsK3AJtKOZUQMKOyRqwJqNSDhE67r
hMGjWidLteI2mcX6zAN9ZZ70g3ryXxI1cnm/BHz/I5FEhGCc+7U0tL6fTaJnjch7Dl5wTXdsp0it
29kzNhaO12B4YAvIDYEfIt10h75L3GkFvcWa2zS2T/IaC9HICizFC0ee7H3weHNmRzFYpXjwOfVd
NdeO3oH7QV9SUjXJEsFQ+Bv6i3w7wjG1/fsnX5fxHONJlAhOLUIMhPoIaZPTI3OZTvAzZBKOvRvk
Ra0ZA43ySnbWvGTR+WmKAyrjMTInBWbrXFHThimz0U3WsVWJ/w1/5sY66G7LRgTlNwtc2GOZansv
p/2fBZ896cEAX5/X1ZvTNOJLsvORrmk/WqFu8KA3v7vBFZZq9qWFo4lRfz4T3cKN7krXj7f9oPmT
TnAVYeyI9ZUuPISxOYw8UOLxbxEBYMDm8PP7B1Z8oiBmhXoXw8xYZPUTIF0b9VkKka1/lIRQBadx
j/HAzepfshsH7QzKOCq+M9XJn7oPmHRFGwl/RRFfD/bwriOzFw3Va9dBcMJSNUXSolCHt16ur3+x
lrxCB0iIuV1O+BwXV8khPg54/NvZWsLNnupiPzUnBaYp9/xsNQlvA2RDn6O/ZI5+BNCe8fppRODA
GRZJkUGzfjxaFxtQiaS7s2WtomRKm7/dSTm8PS3N+Ax/EEGcxhrGe7+ZOpXDMW+Hcg38tXJbdfWq
+REjZZPT7bZB8Afpbgtq0oXtQ6ObfQJi6khOjIoTx8OuHKhp7nQXsI7D61fPv6pzr3i/WagG/gxQ
TYO8V96Q9MT2FLZZLlWC/nskpk3aslXfjxyO36IwN+LJcjHKOKyhjmZCsWPuHJxunNrs2UU8nZhC
qR50b9qhfAJM6qlxGmBcXAY9SbOIrFPc2r4Ii37kQWqrvhIO8ig7/bscJxvttwGg5/reqjxuPW2o
yRnICa2vJgYqWAlWK34l87ji6h8XLgGnpMA/+Obk72u5HSfU8frPpTySGqNY8NcYO7LkeD7LcaP4
A8kcBK8XFq556wMtdeKwECCswt4jX5K1cL1AaOdiZKCrboMgT+ziEbDkpyNvxDYiTKex5DYZ0qkg
HSwio0RriTSPaTsDH8CBrkgPrVN0Sp910B5K+FLST5XfiC06HN01yZfC/EETuw+seqxSPPX0hKji
tFmNv+CObc702XwsTC7+bOJdlP8TE+4MhpMRRHGrURBJosaBvf4xoPcEqqy+M2OcsLHEzPGiALLe
sfcgrOB5dNUNh8MBuIF4e8v/zl8vPRb2XLSsan17MCHsSWl4A+UyiQ2GwN3rHuN+PCtueHT3hOKG
UnN8hilGqxSpisu85n8x3adoPu3oULu3vIwY5ImG8bYom6yvFreMnQYfzsH275ns32Cph6rl+kRW
NNUa+QJbmem70hK8XIB012+MKnpBQBncb7W31N4zvpXnBf09q1f+K9K14WE1ZjCTrViYwMS3LIGc
RtUKASXzQVaDh+4vXBz/k0VGf5aiyNAjkJmf1XdrGaZATXr9Q0S+tKmwZNpTEnUYPSRwx0ChPmyv
p1qqF5fzMt2Svi+JjewgBaIxFtHcfRZEMZDUzdRlPG6Aq3C24D0iuvCvrN32YQRjYPtXmSCo18r5
OBsfdPYw6CtdQOO/bSg2cKLYQVoX7GU5Wcv3dOA2MaF5sX4SLmPiYLSa9yQCgSt+31HTaMo68c1V
9j39j4Xi+sOeqBWNCuCo4W1oEbreiu9J4fjSkJnm6/VHz6o9eD5ytvIiMHvBmvuCnrgZDVibUj+K
GZU3mE6tx97BmAx+QDB0xRqfAD0yqANPsNFNSaCnm6FEKdrMFuRAkRvc5E/x7zsGmaFWe7rWwBmp
Aaxy+F263EEKGNQ3i3mnAIIiqq+nVERk3b76SUdZUSWM3Pe3iE9HyWIlsxzeGU6HRfRcKN3PiwzL
gIW1U5hIWkU7Y3H/CQU7jkBU7eptfj1651g6RmAIiLSCo/ovJPcIrc/Iu2zYZrfD/y0joP+DoqKK
rypesO3CR9c8MJCAkJ7FmCcU4LZG8g/aHFkUIJAlZb5vCoOk8UB095gsx9Mtq33UuRgNVr2iDXB+
QXcjEIXCol9+69NZ6jj7nanHxXoNKv2fSgkNGFTM4s7j4MkRIzBSEZC6IjMBvHbEF4E8JHF4e60D
mnufKC3kmLKS26ZNfCokkBAaQ40XNadP9DzPikW/BwKPdK9IQM3SAPuiM22zgDpwyT02sWioIMYS
7QtT1dFhDuRAyEb2p9OH4Dg0FckOxjlIjQLb0JkQw5zqC5mIMgsijK679sQXL2p4XnDu0MBYT3BT
byWuWhLmHuD72UVRBNZDaRa0/VIXSUxwEAwMbQxYa6U2AvmsVRaFufXGELcOpllNXbcLYzzKAP6C
gGDG9zmhykgrAaH3a9jwH/lUzJQHrj9dgVtD0gXt2j1iCQvm2COH6o6tbHvfzCrGUmJXwX5YpO76
ZRm32zVJN4H0W9TrVodMALR/T0piuYfX5U/z7zq4YQY07hSnSDGB0leKkfEssMJx9fXFaMkQj98f
D0HjwFkB5ds21Z0mKd2hOgjIefv84Ns5bs6+gk1he3Ua5TAEBUiBnbOieKWt5Uxeapm5SHoPzP0P
SjlRjJD5Yl8YUfj1upkExge2kSsjabjQOkjvTklDUHoDEeffjW3pYAfZbOULGXJDf+NDUzDCYebL
JOMpMlxmMqSfNJ9JRXmX8CiH2wvTIpwxFNdEwlxR21TWCCIqxJWV7ojlDbgsa2NvA6E6NkB3GHkm
rSGzHFupLWfWzYGVd+x/ENba7lgsefkObs7QmRA3xxA0q32fQH05Un7CEw1hurzVEdGafLRPJHyF
dFQuRe27YXBMn3TU3wkfVZjjUWM1OGxsT1TQJ5XiRE0jNzvikWWlj4bMDYTBlM95IUzQo5/r75Cf
UQa0D+yYMR0urLm9aeoe+73xWZ5SH1EDGGqeF1YtPkfWQ0T1h2Lpgvte9jSfhNCI6mpPXsAnUTTn
FkSXzY22cTQorHOvlbJ/yLN1OeRM5tegKas7fbh371nkXvLK3pWzBEmdTNlTcM3nRGpSMXTd5x3h
/n3UX1juhhLuesimgbOnCbXX53/sGYO8KBc2C6VLk+hsrdlx/q9QxlodySgtYx/FiaUGDptF5PfA
4FMh2HX5tvi7LjJ9wh+8D7LNOB1ofjb0V8L3AvcC/DmXAHXa9Br47MJ/1Ooh8aEVYteeyNkvH2mT
KTz/C7Trvqph+xlIkkWKKfHxmAYy4FDlUG2f5t72sfNadr0hR7vBFLUFx5e0X8fnfR0YbfuU2+FZ
RNjh05KwsC+VDSIwnnJq98qQMtfhFGYuFw+D9rJWURO/zo5Cl5uxf47s6JEvwQxmZoesW14XoL9O
eI/rdmUA8Qc+7N1931ouN36EvctogF8EfdB9m5sxCViOy3GJGFySK7oDH5D7AnDUlcwl4As79tXO
g2MVmuzdba8FfSPz1aA396IGs2sgym6+wBm6DK1lgqNMBtb6/f2AgaSiJtkHJVY5otnAsnpVFqVi
6nGDaSUfCZO7nj1zNWXrxpTwm8lOoJhnnUBSeoWWk4gwl0TV4aZfzkH1BFeftWeAUJe/0Qcxpugs
CyF1yIGZ5se/UfQi91QUtOulSDXrtXnan8iV0vy5l1INSiqIwJkj4ZjsPuHE1ttOUWj3B2P8oYh+
obRRqw6D2CzH2ixpzhmrsNZS7VH58F80YQ4Ln4eGVFmbGwiYPwcDXwDMyiFyA93NFp6PhBc33BSJ
G2MYBcGdhBsiTd7ptc2H6Xr6sBA7jpzDSvN4zZjcS8YFnlmjrHuFI7a9+xdWkWbAPWhLRHc+JFY+
6EDnXnVCsL7TJOhREZ9qkVWofD1CWbQCOsF5Zb8CArRkKbniS6mmLMsbi6OIYDclxSorqqEp+4Wp
r+sOFqYYxWcDByFiY0taqgIU7vUieg+X+vx782ty6YaIp0NqfKyt9tTVq2obEAoF1uaDNxIv0Mt4
rO/RWjHtLyQ4EX/UF0vK1+fbZ35M5BHK5ul/uCevPxAkPrIQHObmzm/+bDECc+0S3DjbmRSL0fr1
NgSMWRezRiFVGZFrCTk1HiW0hs+uBC9wt2igyvR6pbt29as3p8x0BwEkUW6VjJFmqzrEK2rhnHEL
VE/rqylM6MUUISM86YrxWLGDezUKZUgcakZfF6WFHUddMfnd0zwexFXZzoficqY4El9XrVMhgNq9
4I9i/zex0RiKxBdPoIwYqp2FHlSKIzY17KQNWOWvJ6nOpH98I6ZeCiKiDYbwUVUrhVEUYpoEuHKT
Fm9flzSrEdzL6Iqsc1G3mNQ/VB9SaiORA3faPBjx074Oca+S3EYFgW9Ker8g7jjCley2CJ8LYXAD
SwxnguCjITCs/FdRq2b9fTCLqpODNNmLgvpIT4BzAfFlYfHfewUZ062ni5eQLUUb0OPaJ1KJggtY
DeV3yh2gsqXnAZyoZ9OgGMfzVw8HQWtzMiIEqZZhforH7zEKrNS9heU5arCj7DJUm6XfaEFR1TDR
gFzlGOpZ59I7oZF3Bopen0AasJPtCk46z+vMu06Uyc8lRMruj/3Y8btYRp6EqfFHIk4JVuEGZffX
o9j0LcPLuvwxw5WkX4LxLwOwntA1OHPAa1dPUYbufJ0l/cfM6JgKL1f31QF2fT7mjeiJEPLcAZex
F7T33caFN7/GPTV1B6vflMwU12yvwkaBUf3WCt4z1HdGtyfSm43DqqZxFF/FoDNVJntnMuwMfj+a
NeWhCGSOMhFUzTlfW/GXyWgvl7mNbJuPQ9ZaH8iLw+BIibaOzwe+9kn1ZfUFesaoS3k1XjROvd6a
WMPtAEQO43kOZ3iORbTiSm/lwaRgDLeGIq2TS7siXPdkQJKqPv2FkkKsAzuVU7c86mgyS+um8Ds0
VXe29Zyng6cSNS2g4RTCH47UaAIUG82AHU0nDgxGH+ZwLmmtVLY6zD7aNZJ+DhaqdCAVFhkOGDES
zpGm6hrmaeq7KHZyXQMF7d5u+MUyOwm3tljRdzCYe2lDolUSH5i3Qf8MvOY4DSHiZNB1NAif0InT
dPrBXL3hjLDiHspv6Ke44F1ltPQ79Sy4FIHTmbVpjmdldZFjmCFLOeBOCDqkLuJgaGJtrgdY4lQE
WYPa/+9nupdcoTdpUtuaBbM9BOtRfZgcP8U+ZQzjotE33Tdo5BIv98uawYiYYQg+RVCMS/o9YQQ5
1HPON5sFsu6eUy9OTK13T8PSEq4D5ijL0OiFQWvl+tqQsUbIpaZNTUrhKBp/1Quu+iTqkn01nFxF
RXsej5BT+M7CpvIyqd9sWdY2mOGw89jMh6kH55r0w8HOXFZ+GOv9hDBfKyt9ergHE2EUyZmdwmBp
/QyO/fkuiayrwZdLQSomBixBtqBGO4MvuIILopCjJ/xAVdFhpjndZq8Uh3uAzWlMuJqjrWIeZ8pa
NyRzomQLM5Exwu8WFbWMosLrctMa//7gCuUE35pHoo0CXzoBpdZY1rZ+FxFCm3G/3zbK5uodiVtv
lFgIkbcvETGW1PFb4ugxqDAxKofSZ9vAbYjbUxbiROsOdXsBxhAeR3MzW/NpgGwEzZrNKXcv7ymY
62QRDR1o4l+ZTYb/f5uMCiJbejziFDp2W+xbhpJFjIdnGckRpQvrqvewi4YvtOFstP6bToreht0a
Rb2SjvpMaoxtNWxxGtT7auFUOBRbJCnRdCgqBKrpZ8VPP5E+cGvLNFhAPql5ukgEK1O0XzTG6HdQ
ZIZ0nMLdSwb6J04ZpwpoH6DaJkS5hKFuU0ql6UDPPprAixiaaT1TOQaEqPIKPAxw59dgS6ZQ3xGi
ECVVuyBUr3s+SDBL3SNHQimnvSrFH9j4ddh4Lh9ebK5esGg//VlNxhMerIN+vl8W3aSqbaacpLUT
fZFMrCg1+l3FeTqB/wf8Oc6rV5CSQaDBmPvJdzkY3jM6QW14/3HIVAm+94x0mtfBI27DTr0kvE6h
aMdmbbE+sVv/wH4HszzSXifwbtut6dbgfT3CSsN0it1xUnJZtKnnvHTOhWey3OmkcdlsRsoqj5lD
2E/jpqG6Li2c6/OoyWjxiZ8wY4cR//VMYMx5w/c+M5xy1aIZDJaWDt5EcO5sGOT49HXMfveedREL
c6FsKBKt2rvStmhgjrTmWCgOjWNgWmgBI4C8fXd9wm6E9stpX469MFjTYjXoLyYUVHhq7ADYA6xJ
3abqXNi3THzbxNvl/TImDgNpjzxTEyUvFYC8DGDCNXVBaSiAhvWG7iQEDrmJpbv91apjbDbc//b7
867fhJMz4pMYe/UgJyfc+ODy8d/z3VhgY4UXtUMSALrPGH9Z7zD0KNZoK5U6OJSqWPD8nfVMaNXN
1DgvRGk4lRHGVqa1fs8wUgtVyas2xRAoj4nKlBhyZLHfg1Me+ERFm3Yunzs7PXsr1CGgKPGpApUn
PLDZE2CO9anearTh/OawDuThz+fkaqf90Lv0MahljKO4msd6RqvFtmQTm3yWgE3UzWWlt41NzgBR
UM2uT3YRuHHCMABezgtoiq8Btsqi9hJNCOScHpna4bljlJrXkgWNpwYiYt0Nc7biQfXF5L3zKLVa
677pRTGxC3n7DmCwaY9rUeGiZxjpV/M9j5G1zjHLhesx4aQUn9O+hIzjwsEhDpA3RbDwhx9Hax4Q
tKIFD0/oDa5xDarsi4teT96wZFZhgUalYMtcILbLSINI9JhKZUHWviW2KNFOw4hQi0jqKWgZH9hQ
kpPwNH02xGLUVTBUVZRRJh7mAlBN1q3NwrwrOFWZTVuHEDgfCZCeMd3Av6++ZjDCKjeIsTqf4O4m
bpgd2dL2OMLtA35aPmqwgPM8wD3u+1pSbUGHpzhTJZX4c89EY11oViBAS2qGE9n02fqcKDpf3g0D
mymq0h4+QfPqc1SrXaA8a35k8+LTPnGL8gG3Kun8Z+f3uouTqVg028m7FOF182nFSudAKYBXVdIx
uqCHFGz/jPCOQdF2/DqonBOzUSS4nrxGQphS2zuOGSS3UHvJFkNKnqHuLSJfa0vS80SUHL1HxRh2
wSJm5tdxIJLRVaXiWe+X7UkCfk2e1m72UTmDTUjkFj2s3Adg6fmZodpqvkUGid4c09JRHoadg6Kq
0zhzV7cSWe6v/gg05Ts0OXy9jV2IfnKnnbLVyhHF1A8pNP5hiu3Aw8Sk779d+9CY3MJe3O2ZZVsx
M4iJWIJhsqqhPq1QlIMwLEKT+v+cTx45WW6PSMiWyJ1AGQMhmpMtn3lhvBaqEzscLdKbuAUwP06h
osafCqUuUFL9ng9rTNXKsnPNpoyHfU0ojAVnl4WCvmbSImUJe3La6On6mNsx3mc9JV3bmCBN+rPe
bBD7BzGo7dftsFoeE9fVslSSL+12iS6o/MZ4Jb67bdWoaNKU9Z5XTiLwfNFZz76WLECCbd2jo3PI
Ql88qH8himtHGXk/S/fy38IldLweNsSdUfkWyueuWY5q+ZB2UROaxvOLNcvZFtzfTf90dy4GvH7f
YSpU4rxmJ4puGAL3aSvOhLgmDO4DePrD+1/MpmUpFT+Z2Hb2XdywpoY6/5O7y5V6j/Kv5ep1iBk6
pa2nE1KhyK1lLjWRCSdlJIfi440s+GvGNPcV7nShi8ath5rnAojfJts5AGFgip/T5bGfZikF6rLp
Lw5765uDBFLHy4kqM3HkbvuUR8X9f73qORPJXKu9lZVWh1xCmXL7TSAqpcbSfSTnESnZqWr6smCo
x0RF2T5HxMlRIiKfFreKQcsjxi482rkAfIGeuUgInAwI13UPWJ6CIna9Lo95TnZ0le56gNRBwF9s
IPgMkcVUo4EdXlFDvytJfPw/A4Umj+FiDkYfLiNehbytbBFFs+hfVNiDRfC3XO82ndP2f/eAnfzg
uswnEPfqbT3YaSSIrKbQXMfhF9kIghxKwh2deQMrAW5A87BAsV9f2sTb9eRxRlf2kwMgBtp+UWrC
TuiAqEH5Dg6pCOLLnhTGxKQ94xoicsm2vM5qtRhnccpjhFa00jpu4xUrg+/EfPhiwXeOMC3TRrES
b3BR09mvWQCjNAjcjPlG53Zw1WjzzLA+1y8Y2HnoBJsogwKJUlX87WVHPxnhY7PMOrjmqQMGDaoM
eu3r86jmHJPWwOKVR2AUMgj4dV+0vV0BNUc5/lfaj5gRpcJ9Tr1yQtpmUyjwfTyAMXZ/Q3QJ2sYa
YqZ8ItvX1ltXHnSmR68ck9CCejSm2glW3LfDPiqEMiDtGZ2Fj5ACOXBAjreF53gg4yV8DHvUtemV
DDi/dpaqhzc9Iv+3rpCqMD/9Ty/ajtGHLCB+N/XkKkL7bENXe9CxYy6QfpdGJyMluLPyUyld++um
etwRb8zjgfSV09amTAcn25R/DA2pa8hK9zpbvRK0RI38JMqYD/2oTA9PgaQKuyPxeDMhMPGu1UnX
CSgRkTyVEcmXEVWeXkMDrmkMN9Xt+AazUz1JUG0W+dF4L347jbTpx5EbLnAbSu9psQv1rRl/6uJq
hq5GZsgJTDK9Tkb0+WnlAv5C4TRL1MWfcpJ3ATsWF0IfW4yD/sZs+x0kaDP3SVAqfrEqwHeo6cX8
52btTlwWbqkeh7uWf9J8JRs2n13+KT2BWUjMYwxp3H1EEJXnfaZHSTsQUx+NKqHTxt8gsycALL4n
VBTXp9rWdd+NeHs/wSb0Mndev+MF+n5FeZekKtVgO8d7XQRGjnQunuzCup/jrgUX6PgrqjfwO60D
QYPGR7OvfIBKVO+ownkCgjzhEmtiD/dgC4Jn7k2+U6MlXGrwOAF9mgpQGlg3Fow01Fs1nKvqLeYl
Li0t5SCrHajrYHWJ7m9EomC5k4HX3tcYsaaita6EsE1d04nL+WF/QZC3tfbKo7M0A4hzIQ3R+EZ2
ulgErOoGD0HLkFoT6LDz9ykMTyjqeq2z3yYm9EJUKaFKYiMgXyu46jagvBKZdwWF1ufrRJ7ZlVFE
gc9QyB+3VTrCcGauD+bKoEMoCVQt+otCRdaoTjtFeNcSfuFckd5gHNz+Sga4yWCRDw9t2zAPq8wV
cWRz2oj4k2Y+DTzbLLwz7qMXi+ZW0zCDzGblhesbJuyQQTytjM8/Qtq81htvqQWO4HCcKdJDDSYb
lvkyJ4NI3xcWesxle3Hz7m+XI6eyEkqKwOSNXkGn0upQt/O5BdtjxV0b0dlx5ATFHykz3a76OpNl
aSnnPFIP+3GykGK85KmOIqD2bq7lQQFWoyeQyzACb6TdEVhW3BgxpokVDFntjPrp6NohtTlXt5eW
MsFmoqvvec8hieToJF82Xerfp5IK67qWcxsgmJ/hrbHLAecZ/GCzNnnzBUTNqTPS1QrarbqttiMB
BAiMDZa4PjdCtvnMROBHIcw5aGpVALDsNf5WtFqttVoV7l2aWR69t2pQlZTeS1f5MnlvNzeoUPys
vjC51lCXOpjkCx6miT+4n52CoNyrm+1xzYBz80LpxmSBACwOEXx6+x8TMFqMnHyY3hJ/yvLS4JA1
A+C8f81HajduPadke0CuZ8xzQ7136+QthlXYewA/Bp6/WW38zdhZC9wfV6+Szn4TCxdPR5HZN2GL
j5T9xXC81GYqZYNeSSgOepx7uxk8Jk7w0mEOj1qmTsDyP1gZAdvbQ7XnzMPX+uJnVs8FCJEdgCwB
ECAF4XyiGcgWPfddYntZ3hFXcSPhI9Mcc0MHTaaErwwqiJStqtMnxilDWG1jz9ewP9N9sVYXQG0T
E9xRrPfo1QLg2o/XtHTHcAz1qziO0jl5bu+JQvDbySu376Tq3rDck3prwplDd8PBb5GTfNLLZoKc
83+CeQBfeOtoRVQPukHf8wTlONxd/dmKeOgL+U+mCraXGh3PQ+WAA4j1OdkzcLV5QFbRLokHNACU
hKQKtV6PrlHDZejmMxfBeMEknLIOG1vzh6ad1bv8BVsTcT2g5q9frR88vQGm+A2g4PVw06h4AU3+
1+4UYV068G2DP03AScFTKk80bcikcDnWMO5cFEjjwArswN9P0TY/jYriyfQ6w20HqBvsG5jupvtb
Y2UjTdtdD3ItO2+daAe/EHGXT+AuPh4Az9bUwDODRgBDtga+u7rknrUhmk2OgTmtvET+IeSaRFvw
N57DZitxeqbRPN/2riwloigVLLAzOMHF/AclvXGOeIdx2UAeRgUSQs42oCwjkxagsBRrdeI9T4Du
diWrgBPdRNyzLnFZZeUfkU8icWpNF3jSMhOy1EdvchWFjsLmNtW2N5+XtMuBM0Tsa8AEX66zpQ6i
LC8x0cuN4wCL/MxAawe4NulyXp9rtQfJX8FaVdZ4xYPWyqg/zRNurwuYlXGH+zk7nH1MG0DtrigU
Aqy+Zm543lvU+UywFDJcNOetbFlNMgJkcbSTz8olqDPQsNC6a5sx+iAKDlVGBSNSAPXSWJ0wXKyS
Snj8DrlCIrvYh5fmyAUywtE4/hu8G63mIo6FvbJ7kJ9Gq0wDVTRn3vtv8GO82txZa95IreXaLLTA
jDUSZCPKzThUpjiZlmnQ749uRes040Hx6mCjWGjCpHhAI+3SgyaSpOH3RZTFdGg+jFBQZm63ocX7
kGCsiCP0IilGX0TtQcmGe1bXYi7fV4MB0Cj1NAOF5enhX4dd3PxdDUEy6l1PPvXQPsPInUwJRhFj
olnWwWkzGRN9M14vtfe1Ao3Fvpk9SkkAEBmjEWDnpnbYCOXLKWYgKHAAdPFYy0Wxvz5dqUFRWD5h
PpTF2lH/B7me9VksF/9sOpKl3pDvv4PvOL7Yg4udD+tqHIHlUnFnfdeFD/1YMEIGpsFLjxIhBba5
p5h+WdqD7H5BZLGt06HWyh1FrEL775ygYC6vgoRVVXP6cbR3VwN62scwrlyvoiX05xYEaBI2xaEf
woy/LF9/4xYAt8N9S3VIk47eXiVFT+/1x83Cifb2OIb7dyIxyT+LPc/Z7b5I2n8/ZfUOXUOCkCtd
Sfhm4q3l+Snh5R5eGVrG97wH5oUCrtcHncI2IcrMHKlkSCTJ0ai6i+eWWb9udeDR53419fWyy4yj
s3zL51RcTwMRIArxlKfOq2Cj4zvLqDYPO4+M6Xk5bwYE1yIdGmrmDeg0p0ytlDaaIT3diTfk49CF
SAbENMUVxXbqQ4K2ZqOzwNJ/0vFPnWmk5vznB3eaXnt6lMNo4Om2ct45X/73+Ts1hH3ZEI0HE5cq
b2CumWjKw7Be+UjIoIQwTG+nAmzAARM5vBBo+x6gxXNHYYagLb4LS3Ozk+i4KiARMJRLtAJxULdy
m5w7QZlvPLaPRHorumXrIkWCeJxTewGSzuoIhZIP8JO+hHjyVn1nuSsxP51dWZ7AE6NJTHEcfPuD
DLwOzL5a0DbavFQY+5AX7L8VLilcFktn5dWxEcl9d6p9/OAeb7HGOEe05LfVEuJDrfKzlbYY81nD
KnChF4YY7h8kIDJ3l8fyURiSs+pT2N+Oh8JXIzqg5ULiacqknS5KGa0qWm7PgfLEfGk89yGYeC9y
MYsfgXQ0TeN5eYK+kxv8rzbDtheoOFl8Oz1xac+Mm4Okbn02uQAEBhloDUJ8/HRuBquXRMJ+09Zh
V6d07fkPVFSIxdcvfvOMavvqUqR6uIJECbuXIFFJ7VRA9mIbZmmhlHCPvJm6KG4sV23QEOZdYes1
dsAGFit4aylkUeX+5wiVORX688Cd6B1z8OTvP+mSc18u39As3nt7Hq/ohig8DgHrzLw3KjGMlZHt
nM3EMLVajuPqVfKnGyOUiv5X1qg9DnKLEvZ5tTLAnzuy3rWlxN2SRoUJLUF7o6ob9f+2SF6RBfuS
bgDcaWIbFA1QCbLg5VHHxh0Jlzzq0M1tXhAykik3nWR45VgvYpKzxXWZgeib34SXAqpolWLn5jGX
RS57d3sOhmo5gSOm34O8hFE9hE7qB3V2FVqZrgI7OvdL1K77gDH44Sk7UBUEHBmfCs9g6VbtQPZX
BdUfhiV6xpfdMMqpcZbU9WIUPQBIygd1yJMxel92m9QawhGzTerlXo2npSke9eBYuh1CE88krzUb
ZHl3L4/uPIUsb7svleHm3l6r3EzDugAFUhkCBSud2wY04BKtv4yytw+eXtEbSak4zYGq6O+z8zzV
7x1qG1SmgFVXXNOxx0w/t7/dhCDOdtYyQ6bI5V5ieGWPj2wVQgUdWwCReuDMcFRcfLZNbe/fhge4
ax6LXDRo/1PgF2jPyXtQocCFFR5WA0ktrTZwbB99yO3BWCmSjoFoRR0kfmf1cIWM/HRhOrywwVeM
T4SIX9Ljzhq8E/4aE0tR5p0WuMOwfvfy3scPJt3p6NoiMrckV/zVa/3N8sUNRNACOTq6f63EZYKC
Fj2UVUz2PGofxLR6Rp6ZXxcnVsdEMUdnxkAtwQZIrn+2U8BXYjPjna6Su5imvUiorDzCnBUkOtJH
PiaCJBhC6W/9CigU3bMIUtZqh8GUPrSrn2N/qgu8MODmYyXhgCDy5x+AEiDetOe9wsUh46hvgccp
lQyilviR1i0779A+i9cK+Ivgv+KZo1UU8J6yWa3nP/hNdBcyplW29QkjY3qz95YUpaVGKXZzYGnz
TcHugGeuK5elmK1+SDMbEjr0VefC6+aQBEXmIztw/frUkBwVp0uZQPQbcVa0XSbiRd08wWzZK9n/
lcAh/Qou9p2zMsSE/55fY+C0GsnUkPGxgR6ORISMTriOTbxGxL6lWyJaeL4gvFcDHwoj+PbWBwM3
kO/63G0h8hSU1csugn4pzrLryfiyXDWdDO3obBczEGSWHI1jj0ITySLxV1mV9k2BH8aNHUoZUP9T
EyKUcOfa7fdq/OBmOVOLazGVxiHpHlnYjHCx0y1kAI6GJh40sIygMGRZqHhLE0amm2YwWMCSZgtw
OpR5wfFTldR4urdM7nBtdgAd+ADHrKObiC29Ylum4ZcYoUhC4ZwP3k2HjHuwUACodS2CZymQ0i9D
qN+QCFwfs7wn/YitxZCPY81XeSBiAbke4GYMguQGDqbL7Z6sx3M1GwE6eZCOFtyxqzsX9t1cBDqi
AcUydA/0h7dkbLxDSpv1lJJhvTOK1ktgRzpmDYevf0Vn2DlWM1AlCf2qTmLPMQLz5rojyAy1xP1b
mLeeEjur7pkRGM/W2G2nDI1EmoYKkSd4jl+rWAgotafvznf1sVk3Q2Es0uqkiKwicq5C/ZlL/PM5
sIThzrBvHN46D7NX0hlkmgP8tvlmXEWtLvvFeIie05I/IjuBo4KinvvZ5IhTzhEBHFSVc7DcHLon
5MFLmThmDKELXBjFq1OzOsFSx/qtSmPSbyVU+0/y+8jF0Xw/eGKUuKdSleVUEVXg5qRlwSFcWs5G
L0kIooILK2WIYGQRnwooG9d7+/hFwwUzElqZC6vbYIaURtBw60R3LsjnyOak1OQEKCBM/mVCSoOC
9/37mGbM73M+VhWGczVmjUVVweXfwj3U30L7zUbXe7bP2eeLyA7abWzypZJ40N+b1u52Oq4ekU0s
+wMXATArzQVvjNiKwduI0DWom8ubpOGzAy8VQYrDhDuQ/C7zBrduerm9immzQ0xrquJN3sItVIur
z9IzotIeHddPoAHE0lIWsgWGhoDa+DyVjk/9wwyv+5VkQsqG20bwGDygEYJ2koC1Cdqd4CzGMCBK
05eS0bT8bNPkrBIxSH8MgwX0PNkU0WJvKfNXHq+TZUGKYNeJrKVcem+bj/m6qamwNQyWjCTdXWUT
9DqlO6Fc+skKb+Kb2w822wvZWtf3D2RSmhj80QNjB9f9J6YlDPjitGsym7PbSOq/7EnQ9wEs2Jt1
KR8Tt0ftqLXudCvToKTasI8nUyM3pQ8vfMPNLkPtcSeDJiECd7nvjHRva7SlesEoqb3spHik8ifX
8A1c+dS8df37PF38AjaLtgKMWHjOD99jJZkLLPNFipxWWpoIHFWZIIIGlEICnuA3khH+I/mNzB9/
rjYgU6V9wHZhJVlbMG185tWZxvHB4irwB8Zi3YQh/XLfF5ped/qy9pO6FZd49dlSblMsEWKF4IVp
pNCnf70pMgug8wGLzoj8nqyMr0yOs8dgTgz/RsUMsCSkMLpPSCjhnk0tkwMT/YDvFwpQovAH8qJl
ZWQtHWoeqhJB9nvbEhfgcJC/hAwExQYK1biHqeup6y+UlJ1DJaj+kNrEBcXRxdMeUzX8/JdHXfvf
xdUk2Bao9kn77M0xqre3LDZ7C3sJRIAi70bjHOQYVe8yKFArDRLOldvz7X9EQtV9z1LJpHUf71zk
kqcBpj50nSdeSmL/LCOXo+pClW2rh5EtzounlPMNL4+EykPNuHUMv5Q+KJEI/riwOiqM/zhE9oIS
u2KYBZ2QgcZml1nqG9XZAqtPXvYE71f9OTbGfE8HE5kLAjpXE7YlrTFrCHFkL2Tb3rDV30eBrAsi
jO2ygLUFpWtGlcRrha/PZ9AcSB8YpIxVLfUhv7Cz0ygdIzfacZVR7F0oVjFp3ZFFQZ/9vrCh7fwB
EVnjbFfr5bmoKpNpIYy9bqPc31+klTgT4lywbD8fvIYtOD5WoiV+cnyjXY7xs/VksxT6ke6zDcVO
ONiKwZgkgN5DIBeozcjcQsTCWkyKPxUd8i4/xFC5ho3mYAwhYWg9NNUY2LhbHQcg5v+jBCLYhMUI
d35UHsKVDzlzQAR6R7Kt5ExBef4sK/m/IQOpHC/FanelFA7ftPI2mq03VFYTdSviNHDfWVPLfpX1
MOhr6kIby1klEnhpes7rfmzbb+Nz4NqICdTdd/wCU7sqjRDo+C6gVCO4PpMHWjnsvhp5SqkJvJOC
LMQ8xJ4uHyWhUVigegR65B8V4Uikn7Xg4lBx99WHAJUxs78r08z7VqH1IrK9Vu13EPxw/+2qfmfH
AOnmu7VEalDXLAEJ3oakeLxx7Prg0CMmEDEc5nsIAqMr5vXwgqD6g4q/7sCUf4keTwKSuaem8ptB
wzxKcHRM3P0HWZFMEJECVmPOXKAuM+hkc97dqYJpb6zV50xvyYBWDSEbRXds27gfRqBNPk6StwJD
omdjCxEeC35y0rgi4ZrjnMpFtArKtpldKiykmC6FQaOj6c4Dz0qDSjOA0SpJ1zHxHr/8LvRSI84S
4Vc2a5rV5MY9zLxM6MykY+KWisiiLRw6jgCH4tT+3r4MLKIOEjWS3lOg8YfZIXwQ0pxak8XAj6Ab
xDoqFKE+wHNHzxV69GQpgqWzlKaqT0vFXAm3n2GwcUf+pkISWqY9GgV/CGHwHsCYHzMY0UKaKoi4
8PR0706pmGN9TPm8XcdYjhTHUPNxJNsDqlKzcEQh0qGGkbrpbP2iIQ6XBRb2ZLoHbttD2AsABq0C
e8qWeK3lvRvXyZ3o/LKIUsynZoVqLFnV3zYAHPuIHFxpaMsEm1VHDll1G2tsoWbt74sOIQEBXyuC
3cTfgPSu4v/7JCPh3VS60x7RUK0ybLVrfxVmeEmzlw/th+ROkoZY5Ntl2613eSEtQf5w32GroRMk
7a7xK+pXJ0n0iRxUm53FPPrX701m+JSJ4TyEMMGBrhBeE1ihKcF9e9klwwvBDKqG77qBh6fYJccp
axiKYLtKBbXBWa3xJnAnNGpQKfFYK7kOK9p0Mm8hgWMy2i/TBtj6UXxcVluDPPnc1xDyS+2AbJvC
OjjdSM8XCAnkBaAZcaJd10B65DG5AyJ5nQhLDZ4N+mO9GG7E5r0KClhJ8opn7L6kWg0vbkQODdrZ
YFxR66WtlE018dbaH2eLrj2dgvzrUeY6uL2HvKGmAl4pJZDP0G3oSqMVYi1venEFxvzAE839F/BT
/lK2d+hHeI9QZcx4R+NpGb79w/CGOAG1GQMVmKpE1HY8sIznuVjfGcEcj1iVKgGlopEGpIdFYfre
4NLPG0WnlhwsdqIb679V7UDsg8KkRPOzwrF6O6J99saoQSAUXCEVlEd7NUI/Zj4W82rBaG4QbKYA
dqhMm+sy2Ogm+kxYN+yzj+j5lgYs5GAV3V9c7ZwaKouEkg22uCrG6Zw3pHoiY6tQBWP5+gepi+66
seG9gK4Jin5yOz/k6LkqplxuPkJ0QIrnuHqtN2H02GTphhvv/FmQIeqb/OslJpoBAEUMu+hfbMYC
iHmUOe5H0DaQAWCh0dRCZ+3c6r2S0RtKmp4+ZvlYQ181ivWepEXVLLQ5aPS4bQlTyi4GHB7egovr
oxcXyaTSP+qWQjj9bo7NZ4eFgcg0MHY98FKBY8QwEqqDuI/maZXcerVz8jtYyz3zXpLqMgm+41an
FZ0d3ZjzbNi3SHQzlwhfvA6AKn57UMyQKOOMt8Vapug4EUsj05gIpxmuK0uyRQBZvIaymeexaBzP
eFqvg2K4jx/NwNmS1gul5QjJ0gGwEzZY12ozpPw7cNSLu3uD4HFTGIzkmuA+N7g2QErpEPYNfgIj
aM12MXg+lpSCN1lha9zkj7DDk+qkQE20L9JGSV4UrfPb0i0h5cV89o0KekfG6v64AS8gjd1nr4w6
hzNeES6G/JkOjUx1kEDX6Pi/sJ41yU63JY47zJZC0E//T5+JI5+1JGPHhidZ3Hp/OYxLgWwMWQY+
pr/DRGFbgt9MeitbgoQsklo8LkV5dha9ci2sjTFON1BRMVoYicGsKK06y4TkOlmqmeRR/Zxr7dnn
sQcNTjjyufNhaZHWT+rtnxMjsQJjcxScMl/pELW5MdYE/HQkRBbq/k/vLiZkd2Vpy9kYbVsekR+H
+CyS3oMKo0Tn72j0Px8PrLU0bjAAMnCcg7m26u4Aa0Y6MULUT/VOiu2UV5CojTTGFobV8w3bP8Au
wnH6kV4Ju+jmO8MCxnExrXBJzA8UYiL/KQYoUs+8OTnkFV6l9q9+qSjSAcQppYxtL1P3iZpuGEW5
MPeBONT03QpSl1iNQ2bVtKPjavycSXtdy3C05mebhGAVbUqHkUysgOJ/3duB7B9Ld02msgJ54G9e
W9vleLLd/BYV7qbdRBKebSNTtYRhTWdeRGoid5wfubBvqPOwQn8NLyRKhEcpW9szUo0RevWLDiJL
mwTo+F2ssI7/EOIwizsOlNsSWLts53fKcizxNL1XBGUdkxpvzFkwKAoDnuUz0LEwb86scPp8l+mR
vEqmpOgOO2X08gwwPDUG33o1RkZUpLR5zt/ZeaF4ibJyXAH88LCP8mbKdfBcREZImOQSS7QS/inD
9EvdKgmCcFoeWrse5qg9t17pbP42CZV6QQJXpNLemwFm0q+t/GuXHMDf1L24rLhJeHH8K692vvU7
JuLaSSlDYIGSTlxVGk+xHvsY2kr5rOlTra5bus9BxFyVWPJChZGgzqPW/rXeNX9CXwBPjEvoQmvh
kjO5eZf23Mhxq7Ia+E5Aws5VeMiw8HRaY2KwHV+fCQwVni1217nW7nmhlPMsZMUB4l8/OA1i5ANo
yJI0mRrpv1T21AyA5749cg2elcuLi3pDCDUovIrZEgOg8quxI0YSbQvdNSN6bul8NJx3DbIddcCL
vY4+0K9AzIqkMhpiBatO5hY80bN81fnHG2UCT+t02+R1P8+UtgHeBCb0ctPIF6Yx+stiw5abJ/AS
K0LL3qPzHbdz0IxP++vhh6KsTCqich8JoamiLi2w1sgcdhQHQOUyuMk+MEoeKymCKF6AlwIuHNHj
YpXw1lsn9ARPeyy+cHySq9NsR6wzypHhTRMYUjpaoxaVKZPAYPUGqfZyAasIzNTsTwjAFNsSK7S0
xgGEgO+MoM98OmsBHNYBPSrHM6kQg8YqglqcMvlzQwUnsDn7LXytv9fsBrSCh6psXhd0Cx7w4EzA
OBPvGlJo5baSBPR0shT5FjmQSlNnYkVlJbY6MfWGpPrV2NHkznmd33Op8TPtKB8ZxVxybTxQ2f0l
h+/b4DlbmE6e4/Gff0AQ/Zv2HgfG3jmTIEpWb4/fvCF/Vvb2fsFOdrYjpHvIkCCxnTei9pmHCM4g
NoVdzqKJW7CkEZpcY5JMS8e5lQAdrOSk66b6h8lza03nPde3PxwMUnPREDG3A4xluvN1Du3H4Rs6
wubL6TG4SD2zMvmM7Zd6cXrYLttS1Ipu39JCzPo7h2IjQyr/cBWviqAOW3EicCzGjzpQUicvHvJo
6oetveljIAoSAuMWVgbPuNPwmqpIDEH132xUwbK0SV5R9psFBKkvpbMkwfvB6J5TUItVk/otOsRL
FZ2APR4ssQqhhHLelkp78TqEfdQ/rzJlSUBMCwlXzVn77E6NhWZ37hK41Fzu6LY2VnxpConLMaj6
5glMC1Hb1hdJzOVuO+zIyIzo9amxhO+xZCqVphVncyYu+BlxEiAgGvCRdV6UuRS85HTfuJaWvBNA
CWYYyY0li74GC65tkwGDLnhue1jl8q7hGADNisROMKa5oBXz/HbMoO+R/gl7FYpDU0+dfRl0OY15
DD0HFx0UHWjBQwV2cR35MGZ2H/zVIsfMPN9+oADZTrErOJ91hpPW23XSINGYIVu85MlRDsz1ppaZ
LLZUN7H/qlMSbA2kEkdGma+MCmCvgjkaEt5xtfBbM6oRpff4u166u5uqjH/fpZx1NyIPv+3+pLML
OakKOhn8jtz3PB+utnDts12GrYDAzX1+dhShWqFpW65pZGoUpCwJTKqoc2yQywGQnfy9hXnNxZH0
+2n6oRjpEvgvW7SS1NKXcLCpc2wa0Xwt9YcbRaEJqCGkDaueZiynhBIg9vraxcWcjdaNKh+LxBPF
LEUo3DOC5k7IrraEprgbULBwitkelJCzzWTA5/bwg+lNeiL0XEx3mr0evZuKvpuh5fSAN6ZAqRh3
YI4WY+ZdRC7/muxQhnq9ZZ0PVAwboxPfhN3AgGwFRzaEayCoQPfGgrYBKtom82LAYTJzSlX2zPVK
SgwMhvpYQb2QupAbpCEG12iWS2cz9mIAsSSwRl6dcj5iux/lCnn2y1bQs0x7MIUfcC9OAJJr83qd
NrzfzwUNA9jvUAGulHlir3nGZ3HeCsAeMt6/IOokT/5LW8hqA9f84P3T5TXd/53seG9xcUENFIEB
FkR+5iw1HtbclMFCCUX/a7Gz9gEW3XPQpRVLX/Fc2qEfAtJqxFAp0zlpNo1gJ6HhjAQGJnCLpHHu
nknSOPwyfHqWeqFkRmBG0T5iWBhD63CqpX0AMBlmciPdUtXqgIVitSsi6v1obdIl8L/l20bbf83Y
64DdIc/sHuCwiwt+JZdazTrsnWbEa8+JO0X/ujDBTT9UM0bdDC3Rev49s+MnbayJii1a2ST+o7vd
GIOcRy1QiM1S1R6a9Z40yy807GZ36Iag4OjSzhWJtSasr/9Elqz31w/RjReiDhGQAGCKvGwAYIoX
9TvIObth8cU3xQaUu54TErkFUE7iVJHvTwwRM6nyvZ9W2Tve/K5q66qgB8i1QCOmJmBYWzunRF5S
qg0PBCxv0e1i/o03IbogBNsMhnmKr5gC3c3obc4hSmE2uPJTcbHqccx55zzmktlxlcEAGNjyDPl6
gtA3HsQc3Efh/IttTwX6aZz90lL9mnbEJAiHcfXCrT+rO41CoESEjoMcMdOZYBYoaOVRLWso378g
LODBA1Nd+BYx2Y87TCJScobDau8/nsSSPrZ+LEcEvQuRSy+0rweF3MlqGBNwEF61f9cK72aEwu7n
m+nr9nWIFCxcyzCJq2Jt5zTlYvky6tmtCJ7m2kh9TWv3Lc8Vyg2lkdXp7UKXuD9P9Xj8otKf93jK
m640TFrFNLE52XUbHGbMXhSOKcTnPqfeu2Ewyo43C3a59IrRVNm6QYSvwYGfJMgv+uPxItYoc5t1
fxpRCFVUoEGY2kd7va+3HL9JVDDVXuINhSkB1tX5V1beQcfoff4XYdODzcKJlod0iq+MbuqNHBDx
MxAbDXSyzdOKbqUEDHytP+A2o6VLMpB6Qadmfor5SQ/A4tNhTqo0eRW0vxZI+vRRzVmwebETTNnh
adubVCuzpRzaEXHkpFz2VUPHME/AA2wS/cwarrLvD++fV855+8NloLgdjh+ZQ+3VPynTmd4mC76J
xMQNd+oEnitG/Vwan0wMDhMz0b2EFgKBVzzrCOTCn2ukW7pKC1ahljd96lytKR8f0WvL0ss8T7HM
SGLjpBVul7kTgK9E5X/YrG8mtkdlyQQcnWKH25hRgnJRqo33TwxvBWEuO3yDIKcs/KK3Dg6zFqCv
f5G2qKBxBtSSE3EVx6/CoyOXb1Pj51zxRikTylQL0hmTLBhV6EqZnoLE9dAYmsU6cl1tGaDP2fyx
B80+be1q3PhibTSVprFhIlRPF6IhFA6MzsvlSKXhGycGhu1RYJaRLCoLWcji2om8RXqeZgVJvJNH
HwWbGWRAIkgFcGFHiqxH9BueHHmUcEPLqhAPJ/B5ZRHfN+Bc9r/liEAWmuUJtAqgg+U+wCw7cy9+
P/bp06CHD98SMt8HqUyEXm5v0JXwZCB+9QYQdylabBx0MY8efEmTNiIkawlyfZ9X/9Hz2kzu3T2Q
kBspB+otTPLNi1dgNPbOLSQK0KY8vxhXBuuZxpbTEzn5y7H02nZdGmScAA6g4JyeXi89p4eY/jnS
IQIa1J2kAsgjoi33+J8TOwZaIsPfWKi0fftT66JfgqoOVRSik3BbBTUEgyZh423IDv3jNA0O74sn
U8S/R6F5eJIlWmt5Zvk9x68nxaKOW9K6n7dq60tMGtUM+6HSEECBcEXxMb30t5P7+Qrd703Xw0Ia
oUkEA01zj8Qb5wPPF4xbju/iBlP6D7RaNnblgPqL68FLub6z0t1rvFXPpe85JbAKvPYUggO0pG9K
uEMJO2wY9Bx2oy5H3ieDjNubWcej2cohxklZXPVT4nVzyzi5cDrcFlyF/8RwiwgNAJDQsLf/9od1
bTuNRJoR4acD8bhCwZevAVA3caXpdcT4AwyJVDngYP1aWLW5FZPW069J6JeVlP3+lW2DA3Wgzezv
pggLKujOfLeQc+LG1XLbT4yuK0Rm4nuW1ivqOeeOUAVThORFfz7TnzDd/2xQmqVvxvrib7KAi8Oo
tSHtBbFRhe9Z+hHF1xGlob20IOCCW7MRr/neoscDaOzqR9E8k4qH8Cy+5c8x9njvOLVoGdrc5ExD
lJTuFXcx5tqTX2wyHQsFyJvsP6Y4w+Qq8kC/+qbohH9auc8nuzE7Rj/xNw1hDEfieYZigWD97ioQ
azfOL7/OrUWaCvqrKFC7VxV8GC5iBN6G2ZiQVDZDPgC8MTpdhbylZxn6uraVPCtKkzx92k4EzZ8X
iIbYJFDbJTDxLzCRUXoEDivdaIMXCpGJQ9yO+/7QSeS67RVJPySTGPpPPZupV8QdBRAvBKqijUG4
3e+IVfT/5BZytn7reUOquxjb6/mJCqwx+8Q1ZZGynYhxkUeLKJJasj9Uaw1KrUwkHPL/YlINBN7N
/Ev579IJwGxvY0VTgS9bWWKXs81MKT2PSbpVGds4AajNZGjEyFa7Xp9YG7mtjHdvRwOGu+cNfYZw
q6WUL8wOK3tXGjlygIpwqvbjsBZV4IFz31zmqrR9IV5ooS4KvVm0J5Dh9OussGQCuzydNJSNOjnc
a3QUUowCB3QV+asbyGFo3m9sE4+h2jDD7L2ddIA6AeU8o/vraJTEctOJOw04rCLBnE1QPKili10c
uuHNVJQy4AYon/3IukpGnQctswmHnVdb/HTwr7pjVOr1bGWyv4qeSQN0GoMaTP0qXnhvGfjo5oL+
IVi9I91vU9Fuhi7ulIB/se2NsRfn6znYxwh8iBLTLPeWp7iUjE2HUT6MfUMbf4nhrIWXW2cY0Ew/
XaORETXG3euckvVG3cdKX0bUZ6I82dz0Vrb1ZC3G+TYgBAFzPa7T4BXKE7pyGIH9ehJq6RTmTQWL
O/ZGBznBVjglZdPJDmcnGS6Qk2iMZtXfdMrt3NTtB1UTe5qWMtw2UtATKGEIblRKvFGX4bqTpfTK
QEKEove9IKuSJiffD+p7PBKOy6tcxsf7ZCLPT7a3HUD6EPXJ4e7Zp3SWNs7fAFHcZEs8aC3lKKeB
DX1H4ErU+p+1Vg1vIyui86jvSg8bXM4kBDZr4jPqBx3/304w3bgOZwi1Oja4tdxPE6O7vxklMiHX
Li4i2pDmg6TOfBdLiVmFYV9HebNB5VLxLoL5Wp+U4H6r5T+MMkVz95BATopsYYTWCkuFLTM5qXXD
dtrVI2FR7MfBz7fzuTJ58oqv1vIW6UxpU4AF244MsXBfGXwWu2VfN+J+G+ZhhiunFzIc37Nijj/y
AhC8wKIEiE8h1LB3kkNQB+LrdolmE5y5qdJLRn9ue5T4XliDhPk8Hw5DxlOQxGi1o5ZTwxI+vBk4
3kG8e7IBYjLx7+beOEvJyDc4eAT4TzcL57x7VpgavSTJTpP4yABHnLoih8QQMFo527vGqNeJjMQ8
cEWYXwB9GQEKLfHtqoU/u2tiJaHw7xouHnBpMFzLq7wwWZMfRmBtjjWcKCJj4L+aLrh5Bt6oc2Bx
5Ck6iNBiGXzMU4/4MVe7SBxvbSOy7EQ8fvPfSm3eDGz8tQ6DoeVde6rtd6ofKfwJtY3LnsEC/1Cq
NookTOWuo7wNeJG4gO8py51O0t2KKqdhQKslQA7GTWtK2on9XBr+p9Vla5VcOuh+FuVMPD4CssDl
zVAjvB9JMWptj4Fd6OznHV2qRTfkvZdqYymSe1cUevCOU8Zs7S49OxExPmy6CgTA1yhMPirt3I2p
agcTqhHcpsh814ZL34ic2MD6sBspBkF6FCqY6v6IoBV+h584V17b+caNlqZ37dsfTPNtm4rtsdJb
7nZ6j013tZNCE00llD5YriF4Lw2CIFFaJQgGQw/tauX4FcIoXdbIjfrsah+9zSsGpefbLUqm0S4W
4kGTcFfy9/ntN51plje6UXUx4rL4FVnO9rShzqlwmKsJUbXt4j3+uCSTi9OwAEG1nWVq62GvK0vf
pec+lChmQBc4gH+AC+Hhxm5LxRuOKtYNhQjbFhv7+Vk1LnKRfSF/QHoEwVDuOIJ74WOcKe2b46HH
zLCgl4dObqOghNtQOpge9ulk7kdH5Di0apXRd3ToCxnoWCa3KoBtZYu9bAzwn3SH/ry3EfOaDSn8
yATNQpqRGbdJIBG2U/f5yJ1Bh9WZ0Pues6oCakZBkN1Yl81ktkcF4LbvT5l+PjcIpeaR120VipKa
IjIBWIAOE1RKjDeNQfbkqWIZ3WNNUSfdnN0G2R5DJvmeUullQeqpL2KA04pXUeFkDC/YOGLlICIA
03zwv/Bj2TAaUV2c+Vk5dl45LJ/z/s4b54kVfhgxYgu9eGqBRXHKJRmwW1hTIYvVTiKhtNazeshf
V0wxiQfXUrfWG1F0OA13aqOlXGrEqK76eapslX4Eq44l+DH1vCR/I9dQpHW5k+q53wnlor/BdFpN
aSukokKEkbTriPp9wL2otbPm09BQpp/xZvs5I5JBJSr9h8mGVW9BqrYGENwEl4Cg3tDEAZ4Z2Byo
ZmAbAzxKUkCPXER2zQqWw6zFaPthTQ7fWCtYwwDvR64wZkYgww2B4Lcz6FFh569HqcW87B9TCEeV
W8ROlrmjvO1H3oooEWnTZmF0O5ner0oIg0YJOdL+FEioiIQGxWhnm1nLl85OVG3IAD5L8Kvp21JX
Km1mmFa4enNSSKvaxFx6iTWbAG50zoI4LmBDseekH8wziO/6UyV37rBFYqpSaQw01tOyDsOHXyzv
1P8r7BEH3K6SdRnm9ioPs3fLddqxvRKhOZosSPqgB/mIlMUuBF6GcuX6UmgH9892caitpdN+jQEy
RqyGsBmF3STrtOf0UHDPWa/qaczBLKxFOoLLklWBz6GU/d5DAzpMfxIbWTPhsi7LqtVflg0M871p
HhbQtMEiFyfktB6oPGpMqZ2weUaAcolTUK+Z+YhTeDbMbcAHmX+3NBVbdogJ/NDGy3z58erSKsst
R1cSG7JLKKWZHz1zSxBBqY9AKWOYtbTNvdLPgZV8zL32RgdIF15UOnh5sEeUe/CfEadC91q821ID
V/hul0HZ5xU/BQUTl282GGoDWkWaeevL2GKJmVZqEvqLXLlEpXpqIRjdnNvfK3WSl1CfrW2+6R3O
Kfcf7rnJ07eH4FnxwEYE9JYJdSDh3TBirESknF2zX72SXDFBxZKJfSgxvxZQ/QBMiYfOux4XqXXQ
UV93R3UKAdR78xQo2X4ezFQjwUGfMTbf7zxoZFLj9zOWUXGn+psHbxnLITpkZIJEbV/0r34+3KkF
UBLEyjLbEIQ8zhEH1MHmQXK0xDI1iPd4318Lh/trosXC41oIQjyQq7enbdi+1fzUSwDnaRfVT9kx
yoRID7wx55r7VDwhHDUauvVq1eqSRrrcSmFWmvtEDTMlC2xFZ9im9GaC/wFlw7GYcyik3DOcQODp
Ct53+mqwVrAMprv+JqEFjTwCgaW8dyKjkhSxitMf38RuHj1ZxUIp8l8Ns3tCYBl+Zbcoj7vgNxxO
zt145osSTNMlJzczFwbgRCO3B0G98XUQgBd7ac40KYBB3xMyNHmKJKKGLBZG8NPeesVp5Ljpdqpz
/MEhL4jzyRDeq3LEOIvuWpPtQn329f8s3QpPiLvTVggx8Pn9boqZNT751lXUgyJVRIc8E3tJp8Wa
hV4DB66TZM/ySfBeMzLTuyHpeFK7uoA9JKZJS/Gm7Y4wmTs+4ymMGJ161mKK9YY4Kqc0jpGlAjKx
ilpzrsxNw3ERk4HRwQNhO4R/jX0AYqwlGLTI4R39nXmb3RP4qgMyxR5MKd+lVDm+0FGFVYQB2l+1
mqnQYkLrfKuBYpS4jFYfCzJ79lJ2cZ60bOiIO1kyrCbdxlThU7xBA7jau+Y+a6WTKPPANyK08hjh
NmeDO5qMkSpGHCOsFcW8u3rHVPcvsyCSpmGqcbyZ0Wr9xqR1khdfpS1M2FcsSZot5gmWbo3r5I4I
6vdLYEBv2/oySf0mzi8uveBXfWGsyansdZ/zxHubIpw9Pi9PhlmhkYjVxztJChXqdK8LwjZ4KWIi
xX65zPY0S/OyUNC1zaelyap/t5sPuWl48LlQ+jDfNU6mf90EXb2l0gfMXctbcjN311SrDYnHZDXn
aDw8+Wq44BmXtMu34wsMYlQiE2xSB9cD3xFtrz5IsuY4tLHRI+LiTCPUAtRtlCv1I+pIvqaBVVz1
lGloZhslmR/jLjqPQoEoClepGQSSQpUSeTDcr2r/j9dC9fL01S8VpQ3Bk3dzhKy252jB1B9l2JnY
Pc2BBNzvThwip5+eLJYPgabXq9ShGrZz6FSW1Jz+poFshL4JTLU2ZSVVsg9i7scYQPsv+v1gn3Eb
NS40D33rfC3QMYDXXiS/D5b7jN5XSHrw72goTomk4wJ4FUjKOCwUlBLrRqF70b2QeuosfGxoz+/V
2AuPkSTDlfGwM2nlHX2UgBr38frq1Dy0sHSqq6p3axSCCza5/TPlvUqoz3xU1z2CX8W2JPLsG80F
exy8xUhAh/dVzTgQrxeqi9B6bKeHBaoAnrEnRtkmq3d9+JiBF6d1NeElUyPnL2qWcnDwcLArGgQ5
pjTVbDS1ewAabsOu+IVPD2eLOIvg/dIPsNF9mHgxE8etO38Z0M+vYNFMw7pXk2ig1atZXumcuhN5
gXr5JOduKzhwWdYt7kXe1u4qxV6fMAqxQW3qQa8Skm2CwoP1oBEHk8IPYtKhndYOMTcqW/ZnO6bE
HHqSuMmyly+z29Vu/n+7BCGMu8K8SQKL875sK7NMf1ofagjARS6AbV1Nu9PkzlPhWR5cO9l5KfrF
ipfT1q0/5or0IzUiCEbTewyGmOKkgSSRZKJMrHUJbZHjgKW/SDApNcut6MTRxGJ4s9XRCPDwCRO+
C0fJl+kmlDG6f3dZgqimLNBzhpoHO34oiGn7TzNOn6UCqReJh9Mb2TRgrZoyXqnCMEJ/fD5/zPA0
AtwHih3/GX8sd06HR+kfjCLN0gCuDK8P6zWCEkibskv4l9v5w2D2LTsJKgyEgzMc7auVvvUPlhvy
M+thlGyqF3ZSNYh+d/3s9rFYLBmUldwFHfmsKtt4z96oztDNuYO1PKkcNzAXtiyfrY+dr7qmSW7T
CUCLmT5h1trQSSdjsmDixn+49HW2mFap6N80Dhe0ioSYbWHdm18vyEmodrE+HHJp/GVJx1biQ6dt
tCTRIAo5KJS5GgD1vVGqT6n2vR2w56ca5UReCBry7LPnwDcRSWICyvKmfYrQYccEhnTFLbWBQY5h
Nsuq/cceNvs38P0umW68TdE1v0I5jNoyjQUspnhxg9VNUFWUqiTkAdhpgOyCIZrU7kTh42p7110x
f9ROmEnQfSlFaWDdro9I9Rq9FHjUhhwD/QqafX55NTWJXxEZY5yZ29zOS3D2vghcJrFL71pxiu+O
6wEyXyoGDdN+SzNDQQ77DYLgtgUyNpdMPgNGIB3K8gzUjjr7DgSblHlcwrMKycVwMONrm1lK2KTL
xRVS5RHupaUXGzNIU16lVvy4Os18PHg9NE1mzF3iojLzNW1yr7f9DVqf67NcB55HxlT6DrLVkz2d
XyBN9HswESR7Sa/Mc3Um4I23N+sOGtsTo6jdaKug/d6tItfL4U72HV0ofYFZsQLCcomzZdKMF231
g2haU4n8NEobojGcUDFFUomozFDC5Y0WZg3f+J+0pRm6RLM5F4yrv9MZ1Evx8MAFbH54CWZB+GXk
7aGnPC/TMhqTfYTrwaIyGsrUl883QHBGAhY5ddawfu+FStOz4dH+iCH9QftWsiSy0LQsQlSmCQci
4W0YtIjSkaaD652svQEuGrUPuFLoxwl5hJCgAOl2ZUjmNyqLfmwcffTZcNk39pDDXkfrZLjKwQtY
Y3qnOD/jqkcc9KSn+W9HzwxMMNp+596STbdbhQb1CLyFht/C1rd03extmYS/7uwZuNBRDJvdLs5L
esch1L3Bzm57caKnaPcIbPvLZ3eDu5lhXE+xCWW7JgLEIqdUMzDl0GgvfMzBgngC3fOjQYsohaWa
tiZBYEg3IWE/ZewyQrijIba+UMhgQUn4RzyXLzFx5GUVLOPodubQ5N5bN8xW94nT5+qpqsKtUZWU
K0v2mYeCRRZvuaNGsw/7rzYwFwROYD5IPUjIPNl0cfQuSBN5g6ueEGQT0yZ8D7pubK2kXjsylhh+
Qvs/rmd5dUUicRXCSDRDE2+CWMC3+6vtfALjp/rYv6Sb3Od2fZfkuR8giVu0ice1F4YTVIXDYIZV
NdF4CR4PMP5QMwzcni/P2KcOCrLXJ7HDVy9GSml7km92EumiTxvz6OKOMwIBH9NvKFjO/XFkK/zv
iDsGsjbCJAxSfgRJKIXYxrfFIpm8K9OcqjqvqSWDc/FPTIhHmqR/cH2OWnqYntbqN1vUMDXzIHCn
Av64kkCffA/u63/ph1+ufxdFiSYsRPXI09T/4WZLegB5gcbB7DIB6iF1EfOYDHqbc6xpo16+ou8W
lcHtHx0ZByKGXJ/C4IQ/5Qi58++B+de12GbluXzzsPMHpcwnFnBbP8BH3WUYZ6snQy+rC4pJBQj7
mnqliekkOPdnPeWymY2H/6YsiES6fRgQ+2xTk6Jy1TWvqDHH9m8E+pw6ttaj+1OTLjk68MqtUu++
nicvGTZfKkDiHlJbby+UNhaUlN4SE7D5W5PBTFb1Plo/LwdflREGxXasynXp2N7Lth+o+QV1xrCN
Yyq9ClmPXHYcSJuZ5ID5wjk+yP1Hs9z6qRbPu2PqDgz2FD2uV2ykt6VV7zqtDbwJiAzFnE0L4KZ5
TUFXHDae67rc33MpsXq8dCFQRJP6eQfgGga8Y5xXu0od4lAPd3CQjjS2533tTyshH5k2QCpnm0gW
XOGUSgX5ps9DGv8fVUApl11joB6qd+ntmmR6eD/XbOzzm6hbnC5DT/BAC2ppuPYoFI8jLRDTk9UL
ALbWcfqf0HWC5pOiRnhGbrXppBxRU7rpgLuUMYQs+6exHVjrazp8BdCjXL7W+mVgQVEwA9c6gRn9
+bKipmZOqVcrSZaLcRxS/ohkl1/KBbo4dvbFWLQcztqdyVsVNgPGiJbgyMHXt/CVlqSdlp6kkZ0s
Pf76/P9C77XO92oiMuBmemruDnC8prd9MunV1JIF1V4afrL2omNqN/aLHAMmtN8qAhE5ybjF1Vr1
FsbhoY3YHn/XcN36r1CR8uGjgt2Q+Ih6k3BV0xm0Kaxjp80TFq5gfDuUf2UeD4uj67h0Ww82TEuj
UafBPWMt6neogQRFayPxMDoBRyk601ZS9K7CTDv12X1A0wWLjXBP2uR84hVcsvLIlb3zMwJnQMhZ
VF9Z2E/+GJyg8IVjLA8wN1cvpIKjpFpqA7tF/YHWJWJxrwb4OJh7CO77YQAKBpS/vxljW6NtgJg2
Cx/NVJox8RNiREEreEJJneuqVoFbE5N5r3bfW+1rpEIPWjlrx5hFlf18E7ekeS+H7TuYVZ89QYDF
e50GvETxor45Vhz3u2JIM+/qlPoYyb5SyGmxfOegE4Py4+bjSl30uNpGfdB75qGosILJP0NJGLLK
8Y/Du6ph3kHOigzwGOQ1VaNKJ+6YhxMwBFIGFuxx0p+Rxp//ly/vyfAvNcviVfCJmQgtyEZrUKpA
IsLzC83XtSGETZDmwA5VfNro4/077P/DZ4a5bzX4W51e1stgmQ824IqskuOlCFx1YjugPlGFTWiQ
ASbVm7Unwcbr00VsF5U89JQGeaeHzgQJj4ND2hmkDpBdtU3xKE38dOIFKFoYEe2qhZU10Z8dhyMN
8MKU4CqL2fP2qfFvQ0Z83U+r8O1DU7n3qropJwVV4ToLhqKMV3BEsw6PYXELveiSqB0Oi3w0H88F
xe1Sp/5s+6LbV0aBFSFqR+35rxWtQ2xEF7lRcOzq/Rm2fht1M5XBYZdpHGawrTUFi8cEF0UM7FN3
De7W4xt3+Vts3rV5+th0UellEzWnrmv2dT34YV5APBWlVhc/sao+03tndDst8NclSnZCJdFL4uYO
4FLvkeciPZVy4LTgSy1Q3y9977QpxgHz2Fzfwtedd/Uv7UZHowLZ5ZWs73sI7D0lf+ZhV9S1OUjQ
9JgsNlMQkeHaqTNl5XlKMlJWmAhE5fgk701w6tI/zx+6OfFXo6UnsYhfYbg1B5p4bcWj62T65hH0
Vi0Q5WsNw7WqDQ+1zJcHA/qWoKCBdBz8o7HiZH6Y5MAOkJ/Vak0xkB8cVzk8AMinPejupO6rffzq
KFpc79u7LQjdxX8Bg++iQrNGseXH0keNg4jPVAbcAAbWNSUlCZBj7yecjB72Hq7rKEZomEQAzf5t
rLcIoLbTSMSQlspSp/4GVC2L1TLM8i/d4B2qBbPJsuw0vxHgMIs0kWV4hSW+AenaPhcPT6Dpm4Xv
3ZbLQKuVsUUte4VDLXrQEcTW/HGg2iZNVQtGwBRN2+We+QkP+841/fkmdx5vvQQLj7pF1IGNJEDU
BIzzq1yy9qTZ72o+8GNx2w2vGKmrXWwGPNRG60/Ofh/VmoEIBBKQ1HibWzeCrGrdKZv2igkPAvb5
+ysy3DfoKr+fCD1O/8My3GOQxFeqUkOq5LX0ECzPmSSd+weSnhROo39q64v/S/ufngYl3isCLTKb
FRbRJsiWmW9t1cLC0kImpOWXC0RsPEevpp+iETHnQY9PLu7v8iaCwUFNCR1sBOX41Wm62rH3tND4
XgzwbzLUtMKu6vBvEseOq408fR6GR5Ten2c8S1VAasQQLjSqXRKT704tYWOhY3fuK0DUwPnzcAH1
MiFdevokKz+3Q38sCb0d+0UUMAVLM/lW0FkEQGx5bUtF4ehcJ9FWYjzxidNFDeogVUp9+SpRnPU5
hJxvU3bYd2RQEIxAPLQ1WQWKxJa7R1VK2pyVMU4Cl0CzElPtMP2ij4QIsMNWywR9tdun1IaOG4w4
JbRNGXn064N1M0eysGVLxTpEaEsNzU40+9lcUPhvMfzENILs9iiYKMIAX3wvdVhqlEF2xMlZphZo
6CfNDWnTXehn75H2LcwOldhx0Ep4tpIZ8+4v/9j6tagZQKOiETLfwn3MPqdGKu+V+e8vRpZzmjys
0d8M21Fkcit//Y15J86ZtlJR0yNr8gDS/jjEPOHJFaq9VLu7YLaczRKTlXLeirr0cjA2JxVjpkTr
gAXfp3FXdPihF1xqS6NDr9ULaVZQ4bu6yJiJmw9sFoL2kJGU225lQBMJeWP8x1qgonvj/Q0OUdw2
s03tOUq2MjkSo9AsChue3VhbUMNpoCf+TCA1a/9WCUwMIje8ScZbWDXI2EoXK45RFAigWtp595c9
GgkgzlPb/Cmwb0B+IfJnO4Lp+aIrb6Fs8c4YuPL7VZDB9dC7kEXEik/WUCPeocIV4+bIP+lyJIDy
QpP81N+IFJX6+/qdYw20csgNwVKsfiSmkbXzxZ8/rFV76ToSapc0LsgqSSp4xz+asxpKBKd7exE0
Ls1K6i34ynW6Pnxr4XER9TZCJ1AbcclcCiM5b2D9wXvyuuGbpm5ndmigznKKrnjbB125ACslWPjL
qW7Zzy6goSUTl6CZDdMXbgQDGMHzZU3leGhc6wI74TZl6xzKo0mHwlmVJs3HvvRNORj6v50DDho3
85mR1aPReuzBJ4hzVfDVi5leNeXpZ/yhz76pFeQ9pGyl3xXT8jYh6Cg13lw18lpW9Ddz3PbAvC0X
E0TwQYDYseoQ+lpE2Y9vF79vQIEA2sXZvIao0TbUY1S3DjRAIwp//6gZs2jYo4gjraI0Ku8RgK0r
lWit7g+vGlx7jxyXmLd/i2jGHJdkXMy0HlsQ9IGEUSO4KdYl5BOtyUbxUfOe4zZUrdPOaMgzAvXG
rrY3YeMVXGm8IjxJx6+ISWaP/i30yN1ByuywYrkeV+Gj/E8wtthTdMezb3/xPwRLuIeiUHnGSxEX
cVgsDETDnKCh7Aw4+im4e8OP21M/lBStvhDRX9g1C9t4a0XvfFgb+kh1PJBW6hyUp1lPE2JMSG76
SKYIMLcCh8AXaCa9US9ajkrULGIFmI7VAgdw2+e7ubUyuWh+QizGeevsxvvQLLAIzPj6JrGwjLKl
mfrtbaN2ycV8p1fuIqIphOSf5mnU//JgM3l1hKngqFAFW4O9a5bjifllxrNYubSSS3Iot6J6PNSE
LGSpKu/fOOxhsBZK+We74/ZTQ9Q+KzUgjwMInkT1g8lRCvtS9BO1ae+ffXdrjqcWbExQHwZZ4X7l
Fb7oOKLnGYtu5Tly1tRRXrGYDujGAv6fUcc8OUJ4YL/lj15dEythvjWKlOujS0C+vmzqHurxE5mk
Fz/ZsRw1b4dO+l3ofBaYjfhpnej9as9w/UHIcWRh3ELMp20pzBzo/SlkEBX/lZqNqoZR3oKqUssp
+2eNAaP4Pb01Qsus3Uvl8bJGlFJk1ra/ZNVzkLDaqf9iO+8U4vfoAoLW2qutALQ6DhXBloVJoVZR
iKHn7b7Hpmf5o+Y3YcG8BH5FzMCVtWOFtU2zAzgaVFZUuNSF5lPfx+a1Uq8qiMo+OZ2IHEemV7e6
rRCLgYd8thEos81dZoW2qP/Qe33OKlS85XxqsUy3YNUs2jY7aYmTg/rQB+BhtvxXhcoIoUoCbLgU
+Waudz1AOw/OiS9zevfk8MZLNXFlZtD12WIOi7yv6OL74Ovo6pc4yR5kKwg6T9GoAb2Hzf/wDoRI
83XsnmTj8euhHnZ/LkeyDCjXtTH/OGiX4NtfhGKtS5W5MleKtE3UuTAvbGrybvgQIm3Zo8eK7rwB
x8TNVg7usvBQ8K6UBhlkMf6RcfXo7zEi+gnrovRJkVZE7LJhmpVZZXV32Qr+3Seh1YwkXwoD52vM
d1AIy6QgdDMvgrm2Hvsjrd8lvJNe236p4tOja8dWPkHeCk1snG16STnY8pyZaRX7V8XT0Xeiy7S/
gxRzQD4zGAGPT/ijsJM6XWKu1z09oBwD6O2/de5+0RFO29NIMftY1iNwZd6bGa3X/F9HvbIwBmKW
MNcLZnJvpO3CMLGbrLDipLm5N/2kE70PZuBziUZ7UxfJXvofB+4MEFCoBHREMOCG2KsZTw6ox68u
YHloyIwDFzQe0lRWKVcpeGI4tY/k6I3BHxndtZi48griyRGkiSyHiKJF3Ytlj9nO4GRud7sAXunX
92bGMudeEBfkadRyR71VlMvTP09n+6/kXY05CCeYdK6iYy6h1nkciQrZzUptRtEhjFfKDQQfgAeA
wPbd5insD7ehi/IvAt3ja1VNE7s5RHPGSe2qxmm9/5mP6fNOmRVI2A3+oOUAiM0hYO7eaNzg8TJd
x0OjexKE1QVNkH2UVq4dNOA5rBE4x2QRYG+1PfAsWqdMaRPUsxhJJueOO1d3/OePgVWuXIC08BK/
zfbsNG6GR9MoqmaPv+BH6KlSgm88vjDUFlBHxTsqSlQlbrlyTFMfI+9ougmiNuJXkrAH9ezmex1g
4bLksFvmtuMx17G4BFgi2v5xy2XuPgnWUuBYRCQvaWS1Hrz0iXdTgY0wat3oe3FZqAmVqhnkWLCC
s4/5et9W+x63H6/EK8fM+aRBjjv0IpqOnSC6zKbreu6eydTbyQ6KpMnc53vccnWSW3wX+VCwC3ww
HL5EeImDPxT7vNHA/hnh3QdUfmkLYfqAAACS56hKBp+uvc1+gCIZtKMk1ASqXsAOMqge1thZbDuF
HNktm4j6jlBdctBlRoGRBn87DWVNuYbtiRxOQxV0yQ3e3WT52a+go8b48bAED3oB8i06S3C4Pv+l
bL4FNVcr/WyjmpDv4xkK9mvNCGE8QTSGww/Bm46gAZ67d2cJoemQ6zYHpbB17lDc6MoxPozopkUb
4e6VRDBsj3/WpShEqzsIfcbQSLJwiil4m/GPaUCy2UV4Cn2Vv9C5w7cc56COrGt0okqwa0xds6Kv
vLDHMat2/A4PqWEeyPapbaemUUA/71xFFQ1s4+EoTxe/g7p8hW9A/eSMlkvxn9BO8gcsKQO6JYiJ
8fQyvzk50C5wGpns6NUYQ9wTN41lcTpjvbB2NIXnG7UjS1iqeBKOKxW1Kqm9Eql2Ctw2Gr5cd1YZ
wCLl2FKURcjBsjYZpdTfKCGoxZ1t1ISU3wQjZEyA2ayMnrM3fU6XYHSxgnWHeu9SykdXgXdSJ29a
FRjJd3WvFyelDm/2rDbxl3fdoCMJ8QHRBrCuXZpEdeL2acY1JpG3jO/wKt7FrZmCgysBn2fLsUtV
lQwsG8xyRAVe8wmzwXpqZAw/jMoXDuf01mVxWmQEkJdV9XaqWrdBMsNoB55A4KpPH36u7sbcS4uD
KCt/Zf08PJsBoWbKKRM9u2xAwU8FjrkBh0vZtfae9gd/Qj2DyAJjML4BNk43ttbMFx+3fF/AaJxn
uMeWvFyP62PhsaafImSS2YVynctX6hMxU7+Ersa0UVhM5fhRMdbSMypb5HGShpunpR6ZYgmkstDd
Dn78hIZ51M4HQWXdfgDTh7BAkXhqIWUGeYcWpmbpRuD6AUG3aE+nr9JEbdJNjLQv/dz1cQ/IPxHu
FAynERLIXLFgTMSXXh79E6svM9TrlNqEboY92LvofyuOzfSorL25f35bvQgn9AtwjzBeDD/Wywm2
yxWdStVa852WdwjCZJRmEOHWZjKKIE4qy6lR+fE/6CYDb5eeZD/qt4xCo5cSXc2bwzp+8clxSRhk
V+ysoCmtBoKQ09hTXZ88nHbNy2ajAHX6xjAI1739qobEaQgLxm4VIBOjuQyTpwJTflSJoi2AYeuQ
BcIhOYvpWnnUGmiMHMo0g7sp6YNYpG5FvjQWbek/+ghPIQCBAwAVxCO4NTnsRYXUKGysdJHU9cjS
+eIXCKNWH+m2/apiOUd/cacDYwydGQIdmIobtuwOMXzyMvTZvAW0+h1OrTS58YoWj3ZhDXmIl7o7
fdXd7RSg0nGcXyJHRP0kHofqBN34jpjdOr4MNieupp7liU2iGugO760JVXaCHvna4ReaTQCoqYZm
RIwGTo3OxHvOw2X9pyaK0pkJcKNTJaWhvhZHEmp9kEZqY6QzomOY2AK2s9o5yidy4idp66VYKVaG
X5ImWHfIoF5f/LIdpbbYTzqfx+DIlVPGliuxh9klmWncyDtqpNRXJjJ5SI5olU+KpAu8+m3BFGWa
5/dgHmH8RD+bXa9jdVQ/MJmFU7DyVyxCQYh5Pr0nstW4T5WJw4bdnnmeXCYJ29IUoXFaP3jAdfc0
rPuMFgFqMX2BaK26BBVET8l52aCQ69nWJr0G4OxyqJYXKltV6x9fkBrHTtNR/lp9PQRDmwR980lv
FgU0/55UyZ+m1M0vPCuOxX6RA5x0k5VTN344YH68TOid+I1lo/bp9zMWoH8eKKPwmhGxa3ZVlCrS
TaML4lDTV+uV95qvVa6kbRb1Tpz4zjdMVYbvllAyf4wHiGqgZdwrzhvOJHofJDnRjJVR9NYBZeoZ
E0804wSJMqT9j0gZflcK6c8XV0N8u0+eAkn6+t5VO3kojr6yBZoJsQvvb1+KzEVz6iBeRaGyoJsL
jBTwoo/7RxjfuGM30Vd8nAmWTtkg1LJb0POhdoGdu7IjCb2P9UqKUMgOPWMXPEBxqKxr3a5wbhdK
clhvQGvXfS4d0bpwFw/Gt1Gmlre7jkHstXl0opJpmV9eVeIM1e7HL+2+nmgIK4N9+5Tq90o9+stq
rb/7MHYQbHQ1vwojRGX6+URBGZ8ZtIlrgV6fnqvmcF5OOq951BNik9OU6RZe1S2OOxHh2kC5J1GY
d8AzGQRwCrkOpyR+KXAnP/VK9gEkkwu+y2Pa+XoCx8742oqidHMCQ7islp1XhmncDha2xW459IQg
zPwgW02BGZGzudlwiAqUh0KJirbDev70y1AtQZF+Eygrvu1vxg9JsURkYDU4w31l0D43PdtVJCiP
zZM1B8revE6c0afIasjDSP0s8ZTLpD+VZxR1cqwCgxjt5AucROfuq6KdSO2v9lEfwLh+5wttA7Mf
iOiwop8K4STsY14RqJWpbMw2wezU/Zq/UCDfNu1zirPYk0ugeZpUlCA4x/NN0TGFJy9AKnvgsEQn
BqcBxYg+VsWmUg6PsaRd9e/GInXIpYVe8owDGiporz5dI5DSebZh67pGuNSbAfbSNPZd9NM784gH
WosbONW1TJEXu45uX5XGT3iyR05pqLOa62IG7QBXZVeRqhkEnBqe8sYzPWuLYNXHpclfubG53zua
UCkTyENBU+DKNaeIMhMFu//B/+z/O/MtAKxcG6h8Mf+kftRUds4cjR6ctjUVSIJT/mafgZvyyhx/
0IPi8wH0Urbl6vTtbSg5QU93I4oc+1lUcLpJyr2XxpF1bW78WYS09kAQJIBvJfMamU4hq6u8QJub
hVQHa4SNL84kiTM6mcNA5XedqlkA53c4JQ2akKr3xezMj0BF9981pEr0nYKNtOt7fX6xZbLQu4rP
lXG28+vKSfAEekiTdNDZbCLd3jFHIryaVj0O9smfiVYR4fRj5Az7xmBJ1rtZQYIXHHQTUhCtMvPv
ceIPinMO90J7s2/vEIvlXRNrBiFvhno3sApOSgaUEfrRSKyWchxM867RzlooTJDuVlBs4Iaq+ZRc
SmOS2DHr1hYvI6q3QCAMnsKsb/wRSH6ykJhWjPxVeyoERvsTvk9/KqrVQrbiB13ZlCpSwd3ByL9e
jubT2IefVZRo2LtZxsFIJ6puBeiKxm8wpWB+QiQWmmGxoqdX2D5Y7Np9Y0WmCCAwNELKxMw1uo8g
JwqDO7Yt/3NTjb8vnK8eBGBoadIg/DnJy/yHwszrwXqrqiW5udBOXx6m4ALF+0EsrqnI4mOw6wuy
y7faBVOjRCH6Xdie9xGmqeTosCXh6s0QyHDQfI8i2gvcf7/8MtrmPGjv3HYCkEHt8b6J7YANiYyh
dxGfrDKyXJ/1fQibMAp3KNQ+tNnrejrHkwo7L7B+yv+9uXGV4yv3BWHgtupkC3cI2hLN+v03bIrQ
7uQGRjo3X3bMYAqt0KrlxiOQkSg6i7IJMcOiRfGN38FHIviDFzDjuzlvhvnE29kDruIUH+XXlrl+
Y6DdYD2R4lBu7IFG9rM/qq0Xy2+VMKHmS4i5jYXKvQQK/XUuJ0Ovj5n4aiQbQ3hqD+yLDONPBjaH
u4OHdBUaTffPr5ApvaaJjdy8zXwDci8WDZkicrwVBM0z3Yg+4Reze32yAKfJlWV1jExzXynbk+7b
uGTj/giwL44IZ6w2IQmbjkft3pxckFedBYI5vp+b6fnGyYjYgGkI96Qf5Pkd7TFpfaXuYwq9imIh
K90/nxQP0H8DSZ7qcxJKNNoJIrh5DftvelTXs4ESVpyawKQiHxUd/1/Rq73qI0q66ZrpIrB02PuT
T/5LslUUx+JdtcEKh9VTfUCi5CIIbY6YVq6hjxk8gofvubAhLExXsk9Xd4HBVboTcPk7zNGEnJ8x
YDLYmjrcELyXRsCXGYGCrItm3Fza2Mq4L1dSpkWn9WChsRzMu3XJoOtPV9dY7Q7N8Oj+32YB9wOK
WOQe5f6qnrou+Led6/EejfazAh3NdEmi9djSL75JMRIBjknRJC7iLwjyMKh88d/Y+aW4jUHTwoRY
7OLfahSJ1GmQURs+18n/TDuOR4zCQRGEL3lsQBQCQcMZW30R4g+yO1fkOGMqqE1ns88SDDMsNowN
qbl+ZFRp3+52e3fbxPTy04h/xSyTGczEABLyX2ybwregArz8VB+HmD81ct09kaN67wNbACBQixKc
CJ/rpFRVsVK81KR/SVbDWFzDyx3JgHTzAGkQb+gjAxFs9Fjdh29qrzStNLz2z2IvIni8ij+96AW5
jnXOM6nbiUk1E5EGQ3bnme6TonjJdvdAfw7QqPcMu3c8lpi43JrsZoQYUlhw4wEQLxe+/JsDSUcO
1oRUY7GDpcaTxrXofK1/wx/bHAsQSLJnA3QITcgmdWWPBngp4Wi5uw4pGQa//jbWicIDHsiP2iXy
Sc45mM7CJlZHl8ZSpk9g4Z0WUFeWobukTfWGu2RcrjQHEzgC/3eoRe+V1Y2cRe7UMKPQrf1wuFpy
QemIgx+rFT+G8ddOLxTVpgvrv+hPIZSLvvl12z74NFyXftVyuyZFiNrF1S525Qk6ISuB/I4xxZlz
nM6TI+fjn/rHub+bJSBcau+yVz+sOqfpyFWxL953ewNf0F6ka/637gowCUxVSvk/INszzDAOWWfE
AwViTyfFGScAsnfmlXEEbBi7yqftiKlxdDw5Zr9+TfnIoBLRsUast97YiW+1e5Xf70muHUOYi/1M
BF3AcXzQpNu6Zek5x394diG7GHaNCh/LQJgzjh31E2cNgQasE0Vxpg1Jh89YvHif4dg0qcUznfx1
L1SEzMnxWLLBVxeKJMBfXgX0T72m/7JierIzSlf86UkP2ftXjquuO4HcxLjSPJMwddH4XXbhs/0f
FcCAC5i5rf6nM5jZf213wxFornrbiYYbgOG1rAIWYxHHNgbqVga8jRt4PW8EOarXsGtnHdaSxxZp
x9BEehQBbpfBcmj5Po/ZayBF88v5Wl6HQm4amMcwZsL+MkfPeYja2DFfx5Jr65sKfgcohoybTbvD
s2ATCEMsI86Z7ZUx7hXoo5RLbKeLBSmN9LyA2e7jd+LJfE1ghxFQeib7kAGh9wFFNuNFL7aFD+e2
82CV52+41JdUKEr8/cfySaIQ+UkK3gb567NprHFT36mtWHKxl5BOlD9Fj+FzHp7kCE0d8BBHv0BY
H6PF6aGOBEO8Jz9QGWCMEsyFbLFv3sUbIe1Xh9kafFrPvPK3KqeDbGmwnhgWwJVZGIz1pQ19/i3E
YzpY3OyvnH/pWVE+CiHBXeyZSgOJ3rkD499SKBywf9xXlK1dEGM1lmVgOYAxLzF7EoWuIFYYLYdh
gJMdShjqDYwN2JoMdb1O+thc1HXQ+Kye+xuWLmDGyLCLseKOBgD0wfaOKiWrIkf+9HwmKqDqvmUL
SVRpYTNiBacepTsPTh6pOez6bd4Tkv5ET9EypUESD3PoKexBUUISwrMY1T7JGyELNWFwGmVzDK04
E2hrRRQ8fCI7Mgq0V84bgMSRTjFlWPGij/5X7dVjhd27TG2DOQvVAUX4q1m1JAhH+/Z0G3XnTYUA
LFrnlIKmjzIZ4TzUtHvWtYBXBEsco0Ii/htpvN2Uvd3dmelPOiIF40w1vjbbQnggd/oaqxB0PAGd
p60XGgRnkmeeg8/4C9iOz4FfM84HC6hoMH9vUJQJ9h5DTz9g4KQ78HhKJghX0poLPBjXzhnTnLXr
o8ITi7s4nA+YFiPc+vLcxguZfPZkiNWPRStc5RT+jw80Ei4btftgHGzn1Qcf07YJX5a3KJLxPByT
rEa+jTCSc/YR/1mu5d8CHmXrPh/gfPV4MTiHyd4/MNEEdqYeYRBP4nvFfuoBxsVzUWM5i6hFTpLJ
aV7g008Ioz6GSYiThTBS1ADMQU5Raw3cPqvKzpmpv9RETCVeZQqsnYeCCQirAzFbmeWrdqOeFrNc
IfXe8/WcunU1+bCSbJ+mGget01wM2brIfk9Ub5UQ+1cVplkPvJ56Mr1y5bNw10VyN1mkQ+fplU18
KLygUcjwHrzRp6PSfG9cMSU3hrflAf8ertS+0N1mxTZ3FOS7uc8YSQvZgezMx0Mx24zXzd/DUCAz
6+bTLDfTcFpEVYvbpe8DJhHIpmwnraiTwyC+/M7gyfEekW8jS1dWCp43YtGBjvolIYyUVYgXitCY
UJ9/Y/RokEuXNFTgMRe18pDoZsOKBKKzuXAKG64+JbA2N1icCQJO4MJBJqUudr62eD8a5crKihmg
DXy/QXW7qUvWzVO6Q63A5suZjdSaFjo+EEvGWQxcrTwrUzWxhshsae4aIjQmEgf0QY5Iz33A5Txj
+kSck4BaDPa9JH8xG7lgSb3ahqemWN5JZt8kZjOQQiWyUxWHPGAlwwlE8NP+0v5dmuVEJPTEyAdO
3v24Yc4PhEyBHE3ckOTad4ay5UFFzbqGsQ6aWQ3I4esYReOUKDpS2JWMPCBowExwyHS/jjmv/sQQ
Vfy3mnLwccpGqEAsAXKuhHZLEOQKVCVWCnGGrRrta7njFm67a1JyDcWaUckSmLTC5wbrncF32XrH
29giay68DWNjlb+d0T7m6QD6SF+4qitFmfb1EyutEN9VYp8ELR2PRL5nN6VzzGMqHdPp3xGDUB1O
Cvyc3LvOlqCTzGKz9gMNOSVEOm7T8zi4ejo2b5LS6+Aga7ii5O2OjUqBTWS0lTF/M4nT7b8y69/L
6T7mt1ljkWf6DaK9H8jCYAifn4dcUZ8DjQzTWUXtEkARBFZtCprQM2BUnJ/qb6DeSxqcVPoLL+DS
WlyeP+g/S2evhMMYuU15zu9kT/XKhB+2C9dq7y/0kMjM77iYUMR/OtoVc10sBJNWu1nsCoC6pHcm
DVotiWXuAgmOuSNgyZug0Gnnl/C0hGQ2vVMh/toeJbMiA6tlavzUQllFYMst6F+rHrzUgltCr/kW
Ua5X8QDHKjg8HL4dd2cUlq3DE4LV0DOZ0q+847tSu/vH2sfxiHyWiHaYqL0X3TNRJgtimFBeo9fL
v2LhFdy6wvSdmUfJusRdgwGx1qJn+Gxe7/j3PGCMzfpMVneFkp8SEerpP8DCCc7xaryYq2+yvydH
i1KJLXDKnJPjbO+lasSmd/LzG9rFEj4MAbMq7BvZy/qB0l7TfrT59wA0bNYIedgXzUx3Kox5igxH
0U5sgZ81XjUCamA8nuDu9IAuWAhcFcC7y84GRA6xAKHM+4BLMyO1+UpG7JJfocgKOQFffySHU72e
NbabgiWbQLBTkHXueZNQpjjk8tmkZjptpQ3btz6mdOb5nli2LRPOMK9f69sfCMfn5/aaAKPSLub2
yRUpp3iMqpm9HKlvMP2qvzhtIYUcrDA28qibOCKFicbHg3Kl12h6FM1nuRJMTpHsQ6FCR/7aPLUY
1TPxAQWU0O3M8ldvdREibJN3sPAawbXCq+C7IBvkTljkp2xdbGLGjUmWeN0r7Lx+5klmgHarvj30
5na26w5U5S4Gi/Q0xvrybzBg9uN9Pvohfyz32vlBGuDl3MoYG52mmF7jgzpD7uHzseCKc6NZ3SBu
bKcMe7yvKm+P5pGkxCN64fmhHIwvYZc4h80HTZl8ZXJyHJX+y7Bw/eawrw+BvI/aM4h5IxhanGLN
0Ej9TiAlY0X7FajKe7FpUiW1PyQjQvv00ZFbnSZl3bROxqW6DF6vt8fgnXOJ4FrAyRAdbd6DUTSZ
bw0CYqJDPUgp5YKpxZqKfNlTp4aq6KxhB9Lt1u1e2KHA/7xsS/12hJk1QxKJVqV5tAKMc23WLknC
aHqwv8KuD4G7u8IjuRYO9p6bQaX5LWnnyBPtGxSGJpX12mTqist+QVSzApFqoipa8YutJ/VclpnZ
mQmr8wLCgG4EGh2kqsQ2invJxE8olouu49sZW9UPhAdwPA59W3OznG36GzavW6yFxL4K35WjZXwd
IuwqmrRaeE02GT0EyaHAKUEelWVllAxHvMv4xwy09Mv6nB859pJomLtqdLVeMcmAai9WuaXVZa+V
bcLdR9+/Tfu2rlgCSBbJGcnenuBDnhhAVkqUEt3tlwCUoOG5yaRdTCCcfouxV3K862izpQqOg6N5
3xnh3u8V258SiAv34tVwQIlSTt2T2wHinu6zvkv+Eb3EGBrLWHQ9G5XY7oq/BeZMcM0egi7BQ/WM
5wTJT83IxvP+Yxcl7sYjCBMHFcc44wHW3vlr75b4PxdfmcKr3iXLb+nm7XokrW7ru+fmKk2WK2E8
DAbl6clhAjDnDHy6Os3/8fV0D/q2w/9yo+7gJsmGDMhgbsaYJBEuScnlO2W0g8DBod7C6shOwJ6I
HMQ6S4EgmJE7XU5Py0vOh/F6Y2OWqWyppEHPdy5oXAgvfRzUTGcvUibD9cbTqGEG6XkO3U5pGNlc
KtqhgKFJ9L8xmtmneO9Wqg9iNuwmNHNKxp7bJKZXTtdCZ6PRFPiY0zb5T/EPjSLl/QunBfhNaBB5
OAR0PY9EB7u9Xq+cwb2rGytsvJXy3lTsG8upUqvwtv94YHPghxp2I3R45Ep49z4Jay1H8R9Fp+cV
twLRRJ2G4UtcbSVstBUgrW5fRGK+x1K6xZoRDfP+B9AhOyr3/lMmPOj/pkc2lzSi8NSprKFXZwzn
dOKLAsFhs+M9hnfliaAXxVHS2Txuupu1B/NaF1n4oi4L8dgP0kUlwu20DrFamT2StTHSvBWSeuIK
ex/TgGZ09gTRymtRgFDEsHhDMukxndWzaneUfHgGK2xgHI8yxaYukGiCcyg2H58Ays86BnQA2qHF
2xp2N32phWyd5x8PX9PWiFi8hnJMsN/VKNC26rqjV3ewpqd0hSJ1/MZA3JkRANogbcp2lynLN80+
t4wuhiOo/O8ZtffkmMJPEpJlJq/RRZCQdbxtgs3q+jUtKaQyOMdu8FOBMc1FsADE3s1bpTCbgX/X
Q78NHA1ielSQZ2zw2/bEBjssFVYGEuXWGfPRWfgvnaatDyhnewsKuowZkfjtvSW1Ddm06ligUmWT
Rn+I0V0yzaMqDD0vUwWF1YnfQlsOE/r79eGoa/R6lpptqBZr7ZnkRexHYqhNxum0HBrAXT88G5lt
h4sZ1ZIkQ90kgP5OUAAxWvHcaXwYmhv1n7b+kE6FMpmPoIDOcQoVvvPnJLW+eOUVq+jjJrAqE3Sb
TLM4tci8rkjKHdNyCejoeHoYu0yXrUcUdAbYh4D/4z0G7j8k+8BKYseRUKlSGLrMI5nGWxjcBbb0
CQKAbIzEkkZPPBVCpIKA9TxgKY4nEWU7kOTuK4jTpf9pReT6Q0+p+WrjghD/7Mg+hpyl7npErRYe
SCpLznSESG9fZz6jyHye/zp+WV6STudbbGUyl9pLHS0d7B8lVnhjiGwfjmzojfxVrIGWPMHnH1/S
LvF5ktpJC0qR/Jav0Y/+MrPce+iheXCDj1m9oixndh/tF/QbxO2pvayxbS2YCEA6nUgEXaC4NS/3
al4yn6LplUNvdjL6gHnm/A0saAl/8WT2kqw1BxouVGqG848dDtG8AbXCbZCf52LaFDwz+o5ZTA3q
xqKmnvt0d4Hm327iTDFYBKOh4UjZNWKpd834m7VEjTsGDg5fdq10M+Lih9K1rW4oYDtIadXKkIL/
sZEou2yiohK9AlipSYaX4hJjHxb3c2CI1XYQKVPmw9uu1ai8rHMENkW1a8jWdzBR9m8qVPHvRDAX
/DwjbLLiL6rfzG7NHtVirTWkT1x7tawBh1Q8yYB5Vu3s4ectwKQHvSkF5JN21V4oCKzzNlIEYp+E
bAA8LwrS7yJeP7qEnKfn3G3Vz+54yPyAX4q/ltoQRMO4rW9kTr2KyfGaFZ9QWsce38fgFP8err/f
TnxUJksSgdW075er/OX6dOEG/jazXkf2BCZSSVWPqzq90ZHGXCrn+1hoaX81q8C2SlUYTgBtvQYT
8CKjJaaiGO72BaZL3suc1uhaLF8qXvVCa0epeN67xJ3Nq6V6nVHGkaRs3bPU8HXfhiTGimHrspBV
RG0KhZ49lgfabSoIpwXDQeCPURG21g6CL+Rf4Cgnm41GkyCbDD4N1jgouBi5mN1Yw4b4BpBIqpY5
BsowIYbwQHRmnTxFJyfCK/V6JlESKGfuZTAZUD53ZO/rkbVe4BTetLEvIAsMCK2U+jEZGWLqJnpa
55ElL49gwqyIVZUlBdc6g9xBNwdS9tj/B1eMtlJgwlUN0MqGh6RWihGmifVgizUIK9PjIquLVxTH
JlODcZi/TsnMRDS7jG904a7epPBGaFl8p51c4EugBzugGrfWrFy4Amrb82lqphKg0jp5ym+MJT1G
vBdfrqHGWREieuCkN7aW3AOrSFB6zFv3dzS9d7SE4Ir1xeozdfHvkdaQpOdmAhiMicVfsABE1Pma
2iHCv5BSl3glz1upf6pWU7hoe3vw1DUaOUrXoLvU2LeskjkDHNgIEpIAazJWzHSNUe8pTNeWKZq+
aZVLUYg/ErbVoe+x2IGYJcFlpnnsie93Ch5NuRmcyQJwD373prheBVjBbL3oNSMtfPv3xvHYkjvU
wdrUJ4aJLwgaPxhmvzLJukGgBn8h+kzOQ40G60Fr78iFNl1N4Jwqm5fWQ88/zZzFhweZA9R+UbOB
J9DiBsc1Zy94mJxhNX83P/Q3SvnpokZqQ7kyJb2zKiBCvT2UMdLqFsENeeSLcPlCFI6Q10JtcZqB
Ze9eofYBEV3goJe4oqMmejJaN2ZS7x07lAKNzh/XZXH+iYT7v0mL8qrVDKVOSz6HiRW8A+yZYaEV
gKvDTWgBa6Ko7nqWRxRTIN9XUburkCPd0Ou4E6S/1RU0vT4/qFnO+bQULTB9prm0dATnyHjzjbS9
2XC1yrLsAVym+Nj0DKb3v8alOgN2DFG8kTYNBHURdwjGPv89o7lzuIfOIRyLcz7KbIYat1VHzAkP
0JGsyZwjf4xc2lkBDljpJUFSJ5r5Mo7BGI2HCx61PZVN6fRHjivoIy/Fabkb6IpsWFBlPzVBktwq
k6iRSoEwK0f8Kz+q77jKqQMbPRi9+GcWbvPOPtA7IxgjlgNA5r5Bl6qn+WEsLOvntrO4PJ4iHMy/
VaTLY2koq7ZZxlijsgbu7Iu1U7oEwDiKfSRHmpi/5VG8kgKmGaXt7J1GZNHaPhtC8V5Jjbma+C9I
+dYtrvh7mNfSGHqf7E6HxpdVK15aBw9ZWw1p3DSBqsVDKkc/+QSkZBTrTyXb1gsuIGJGhsZHn+oE
M5SFfvLqQj05AN6jD8L26RCeAVph6GfaaAG1umHL4QffFBxZeWl2UsOrNvzwle5yiB1tScaM6OEc
h97hsyEX04aWF20Zk9n5xOVRKFc2n0w3jY21hMsbmtND+rtTMXVnduzr1D1IDGTKqsUpSY/6Fuv0
5l2bU0QPgSj4rvbGNAE4pcu4fWZqTqh4wXzRvVkZqHDUdW+g17wJwtcvX/vuNyf5ixTm10DGOU3z
9GXZpSABjm6dO2aV9dMMhGjJ2uu5Kb17sPWBa0auEi+fkDhkZP8Zu60tBVda/tXfAfVp0x6a9HSp
yAOXUpYkVx3u1dZyD6FnQ1yf6IkTUpAkGANFjsSZYkYexQWnL8gSJcSXPYLDKgd6OFL8W9FK4CKo
S42cC62g/FeiGFtF4gLO58zrkMa+RNNNCSuHSR7Y2xa9m4L+DCAT4CmXVOOODG1zIunLi14c4sz4
/WZPsK6pfcXAyRih2oo3RNpdogW8qvjHhwOiKlufnZhfehG27/jwMZEPEx8HaMOXZvP+FY54GZho
4ZXZdomBJggzezAf+T3OVzOXDiNm/FRqZUkBA/K1T5DYA7ollzbR7uByrlJVpIAKkDPi7wuXhjxK
BHCyfc2c4xpLB6YVg8fQhRSeuJyySUKG9BHHpmAeySecKJztVpu66eKyuG/OPjJQhC7qX/oGJl3s
/npTezW6hahRHQg46+6dashMPrS7j2YkoMVLv44OWUqu1N+iwQ9Yl2qqQYV6whnr407fJzew+Ky2
qHpf7J6QztmYRePOC+RZWbRI6YcRcBDZCNXbVzv4bivP0IxTmMNYvxlgxMu6BRy3f5gS7jZw+aVA
iwaociYhVARuvCPbKPBC4Ck8/4+QXxS7FQX23RIxA6lrQKnVxY6Bj35dr32IYEp+AVrPnbpBaLFG
wL383JnNturHvM6p2XEwQd0CNqwXfGrAjpsJgpD4w4s1ZqxscKJKltibbZ8s58WIdCBkyGgRUXlq
Kyccvlrt/6m40zEDyPe7GuUQilF+mvTnw+2zmiifOPHblS6z8DsTDKXXnMD7nuPgd21Cdlm5p0bG
j/uMIvFsuJKEO56n38bqqley2BiRcOzcuIzs2jh5OKwX9hRVwLlcDrlAbbULP7I5ilOGSDvr8hCI
qHazlcaMW2FDkZamt6pF/bvhsSJyWr78fwnL6E4hFKqOrqhlYZIg2YAsvGdvzR4/jBA5qO7FHyCC
UJW8uR63kzMEmP4WN30jWv3/0xE7TSGgA4ifBq/+axwUbwVbAPkw2NdXXoGhb9qqMK9TFP8VNQUx
dP+euSvuYFjY9RebBSt5QiyXJZVW+UPU5jNxV7w79m80UdYFVFHDe0xLjHmWwPVRz0RwCR78lL+k
WPAK10a7mY/K87dcGvrUk3XSooVxsTGVedijin8Bmhpnx20pb19CTYkyHYIVHSnwxFghBkHTX7Q6
RWCC4I2toKSYtIglTM5oyXGuevJLFw+9hRSVOrX77hWb2/5pVa2Z3QVV3j9a5VXni+I98NUKj9S2
AEafwzrOz6r+DxKQIsOuEMqYGS0k3vOp/buBSZFlvcCQ1lxv8PINPSfZ+9wNjlw4JDOOdB5jBvj7
BrALGyyIyci7ucOudlt8/buFsuFJwdcTZx4UPcJIFNQLOwDxywaxxbkQ7uXJ1TEOPLAV9OUWbbB1
a6ur+EZTWAwfEAMuZayf7TbqsSnXNzl3NRt2Urk/NBYT42i0SQXkPfSl3Kp436mDj6LM+MOvUZo6
VsnPKf3Sdxvg4pkJXqnNqAsnbaof0M5pt+3W7kFIwka9OGdlEkQebL0bbDyT9L/eOhl5urG8QTqz
KpMwd3MeRGFdapVg2viYqqNzixUHMbZ2vdqjRvAyOaEyApITJgbm4KEvQzmKTh2iaF6dcQMAtIIa
3/JGhHfv8NGC96n3742eYhKMgbxHoqw9AoB61H3vC/kL9gfDjsvQj5qjkFghPIDXVnsIgY4P320h
ZJnOqngsbJ5A7GExr/0kZOUyrruHIYAeS6HlsQI5WfBoOeRLegoob21822PEDHl01CYC7YiKKcpT
3CYFmJT9LkVIxc69HEozbr6JbxvyXuYQSrssROpcTtmvUDPaxm161B63Lpnr1ClITNM3y53sUeJg
QpOyDIYORBdZU1B1qwuM22o8aFMe4bOrDMqTpGnUg54DEX0gPye/IOGsgH9bnBEy/76odAOaqCyZ
BLK9gcN/LCjlTgCI8gvt4GhbbkbpwY/fim3mgP8w3op4uDWAStufQ9CsZLwoRwShLrg2c+IyJhPw
5sr3jiJ2esWXSO0+upd38tII3vTWhpW0b/wEx725DnqTYxtqQi9qV2Toclt+4klh7PMPaKEM0xZP
mLAFcHJ/6rWqhI1D/tAQBjimwScri0l6q8AzqGFvqfMBp6/51hiYrfJZNF73uRGK3SQPs/TUuT+X
SjsvhVBP7q32tWCx2P+EuQbgA19Y4es+6YpuangafGZY0pFqMbtvxH+sQPUs8vUwBYhhKbs0smfR
TpNwlQyvgSfEtTPADXUuIGzktwrxgQTT46dFt7zFQIjX/psG+/eFu68sQFTffsiGpGuSGhKZSBtS
mAus/iAt+VJRhiMcS8npyPxwLT7DZHmoJpss7s2maqOV9LdgiFKRAIiGIOcdwYneXG/Aos4hnEEa
4HXhDuYOxvaf42yrqsfsFBxdKdTGH+IEy8nZZsnMWjXwMqF4Cna9szTObAZEFFmleu6oIzviIjR3
cxeoQqEFNYgTMysG+KzOZb5eSwGXk88lqBvnD3/nh5tSPUdOKyQyE4wdj8qkRcvioE6kDYpoOeLb
abebfR3ItVsI0ly2j7+GKObTXZS62kXT9m1BlYM1IopZgfTWv6+qleMHbh+SN5cMykEAIHcc5VSe
KNz1mvKJoRPDLYwRm6c5KoXw9TRDDfEF30gtSil8/iUN/N5dEX0UK2B66XwDAPD9iEh6VcqFJ6fq
7LXjGZq3Mz2Tk0PmM+REUMff+bfpgeW248iIMU4CusX3szaljARQWQPdhZZHDaQdL+FPlcYSbsmJ
iXdj9135G5CKlc9iFiXLs0BmIGErsB5c5QZNoZNontLtWNe5AsxlsqOGS1sePulq3EHFTtDLGIcn
4xrJ/t0S3LF4GN4tFYgh6W2dK6O0Ttnx6GN430qNeVJnEow8Mhoy6ZKycHbLMP9Vv/4tXnF8Ol15
fyfkfCTiuZKrtatj8qlOWQBppoUYqgyQLA0vLzynpDxYeG/Pwz8WJ8zxENp4x/bY8ynW3B+Y9Tci
pLzy6RA27dBrExw9irhiM2JkLSimT7VNvPSBiAyreN5n9gGdqw2jyqQzFtTMCPzxV0AJ7R9MLEyM
xA+1PFYdvSE08d4m5hF365i7gDRykBfeYXm/68Myvv845QcH9ThQwuGNzG5fh+ndk+z+4qq026dF
IqMNfXt3Oyfgmp8uFD0lfIensbR97ZC8dDVFCpPIdztlvW9kYbLcTpanYZHFZ/3gIyBUbavNTm50
vhcRbSFGfmCwUm/6ln8aQ3PsHhXE7cF4iiww1O5gUO/FxqHx+5K1UtOZJOTUBRhUOiGRU3F1R3sx
gugs4ktGN/bMlXLMyE5A6BaVMNkvd21I7gBaY85UOlfSJ2jfBQ/wLjJAs69KoDGkbbt8qfFFus40
ZL6s7Plt+o9X31WQOc9AMXI3VbxU78kpTUcD+eZfK3l9rwBlk64WFp9KTsmeL3PAPg0MsybqLi5b
hBdjeokKMlGzK5eRqahZPNTzjpaWp98fkKwHdyQg3ER/Drxmia+0ZttzfxC+4njguNwca81RSXku
Mif4+pgaymMdvex/zUss2XQu3vb6FXI1M/S+yuLznfGV96qfD8gdlQxopN7gUad/usf1pg4QjD2o
kWGGX1xWpUd2DB01dndUJ80GA0tN7sG7pYxEijJNAhYYfdg5SX2XdK9kleaOls7DeQHZDLewmkBz
n8NFNw2Aklzm0ywVTaELnXTfgi7LTtsFmB1/2FrwDXMYoRDGTY3GXUngVuEMnCVBosQ02YQdmOe+
0f1VpNy192uZ9KaenDfKmz/3lIPRdvaUq/jP3HiJCQjzNaiZ8yDlgzz2r3brqk81DvnHyCZuTjP1
aG+UG0urPs8++rMUlSR93atGQQVU/OYN9v/7XU9wv5CHMIUKemdJ3QDqcixaggibNo7+9vfNE84g
7z9ZfL/T3goENTSE1kKMOC/CJiJX1XKHnwQGioB/AF0/1pasKNQsy/pekvtkZk8teqEGYQhz0HLO
SkqZoMKj+8AhLGuFmrTK/dOyYDdSe3c1PwJPmyNIlg7S+VohL7ySdrK9xm5ltxxgl5LKtnDab37j
7AazDzR92gEPh8YTset9kft8eje9lekbaQ2+qyG0CzO3v8xb3Szho6xPL06gcvyRXxYLq2R0oE8R
oEqADyh3sDuWXJvYeyJzGWVyodAxQv8zJYmkKSTePXkDLlJAz0Tgl/55D4LLPtY+zekZZ1C7QTfa
UlMQz4x9CyijUeAucogKvfgmcUC9j1ZBE9PhHXDTWT8GCx46M0LDM3K9P0yOMadKt8aTlonX8tiZ
GgX1gxE+yayFmnomUaUb8290csI/WA4Yz9UfAmR3/BKi8w+sXtg4gWHqEXFAmqOqXuSAuXFwNITC
c7gFQc8bZRMPao5y6NfzqUD+CfwlAXFDTO5AMgjBTSrqrXjj8zrPJYQXY3G98svU/FORw1ELOf56
UYFMv2Dn3A1ifDOClBdBmOSno96DlH2BfG7f4DyqS5GyChuigwB4f5Bcoofh5sSdr8x4TYRACtus
zSl1n4ThXxBSH1F2udbg1NquRO1q7c5FYIv7veWd1gN71U69TNoN8pLNYQbqzE+amSWI/yy3I0dp
X+2q3de6QQxfWSm4V/tl9xQcmGQ8szuC6M1K/Ul7UgLIPRVMC5Hxse3S6Aygg+gROEsMcFASzF8b
RdqAkjE5WnaNZRuPtLX1iAOqxOulQSh17CSjvl3k602XxXWOa/0Jg/ARV0fbo3zW6wpRhYNpvFAc
6qhQ5JVwN8smwk+CP0I7+mFv95ZcC7W/fcjInMjs5VEOtO3RTQaPAGSfkcptRQPlBzF3UzPtthEk
6bXvzHH7YRh2PYGrH5wPHB9576kiXASlIWa563rT6S+16t/ERd2YITHvygjpqBciukSRzYnY0FCz
CQHD1QclwYAantqpCbd0hb7V+C4p+NzM3Fa+mLGi8fAmGSS7gPy+ibaXUwsbdxAfDTS8Kpbrsj7v
aUvIFIIf2IfOh5a3xiY60kSVUcG9SRiLLdl4Qy3aHTURJopVfvNY+9kqmZxEZKoYG8daX3UsL4Fh
ijv3/dMES5s4CtJhsPM/WMnGt07EIkXzPLkWimMmFGymdeHNC+ccijgfIg3eb+iPGTCN5g4JlwLG
OBlXqnZl2++6KasbvRsF7o1w6K83/l17m1SnJLzNb/2YjtLAJMGX21vOE87o42xADuCdSDicifH4
BAXRhEG7Sa87CPDyrikc3orm9ymlwc67I6jyRMx2EXR/Mu/Bdj4Ece588teg35UfGaBSa+6LIAf3
MfTCoLWDWQlRPhl4oFikrgtH0rKJoTz3cW1HaogPkAwJnPtrb6Qz2/18OFP06syV3R2eXhkl/lfe
sFGxx9fyuv4CC/TSw4dSRUg/S3pja1od2oJDv+FSOtuI9OsKVdiNySuzuy01BzV0w3b18uEKgiVd
e/Lo4lf0qSjnNqNwDC7xeD9znjmx/xjlaRFLOmyLf237gnrzNn2qMpzqQbYVG4A2YIx2/MwgAfU/
UG/V8zC2dTE9kr7WIGis+kL57yZn+TT7xl6XOXSyop7iYbsXU848V4RRq4CGxVdlH3pvkwyvvdoB
qTg3p9jzovOPuh02J/7v17QorQkrO7CnLgum0t9jIYxieegCcdc6XQaq9YnC+Ql7R2aRgOrukBH3
SwiRRXP1xPuvI6gksmviz8kxP6carj2WJlvwXh9BkcKHr0isFg6rFhxjX2rvP8PXdCYQnCcB6IAg
e/8uQax/GRYWMvu5qAAiV4TNMg4Rj9jW7z6lU3ifnbdi5skr71fTrQouy6nGp7Z2OyLpjvw07uj9
mPQ9mYE65PTuiLhFQ/NzjDTrzAW53FdIYoNRUylI5xu1vW2TJyUmYBYblYWLJo+c6uz1A1ap62C2
vkMJ+20MaNaTZd8D9gZjOMDs78e8HhiQ6Gy2bfvsQI9OfS+a/6lHmUg8MJ4Nv/3kuiSfxhumOx2p
v98dlwmSBuNLGqs1p7ItOlx1PQjEpAlpMII4XoU6r73e93jAzmECIG/gIbvYZZtXtcLm+VRtbbcE
AEBIehfC/4oYENUI7n0u5JaQ83KbCnZBFLmo30Fo4n5TDe9nRqV20zws1Z2tAEtAXC0aRAbE2+DT
/8QglCRfa/koopyrWvd/vekq6z/1N8WUMIJgjse28f17snuacvrG9Jw3CVIfFweQ7R+nbMPz6Y/E
woPDEgsJkJ/pv2FxqkXnZoeJQp3BEzhUy7+J1lqvZncw9RB6v8fS6bkSE3TVLHkM92y03RA+u/NW
sJdOZZKCO2kJUD3qHXGdYE+yh4HzrACtrrGS6zA4j/6T3yfLCGhcToXDX0fhURWlB262Nhw2fsvO
RfflQPR84hs2wlhIM47XETI5nQ3M+ZF2dkpYlw4jI1OcuarCvjam56sbBzcNqGV9U9mq0N4Yy1CC
qcCFJKUA50TiHafEFPa2f0q1rYjLbQYTijK6mB3yAqf8DxbBKB/bk9I/hiRPNa1M9Y9PkQYoc00W
wsSbnQAPM5dxfzJiqygO2bkefThrV1ZA7XmoyJs842m+3Pt4c2SRt24cywumhReiHIh8XY5JIlXT
HfXZ5BageZNp3OR8qbfiWPgaDKDxR7pWlE2m2NQg0ky5dVHBHSM4w5sP+KBywrJt5VcPhu/ucv/a
m7UFxhaTPK8KvYoY2BcgJ8LOVymGQsZ2gHKSlw71BZZAQXq+6iDE/XqSPWQ/fJKcY5BFpNyFvCa1
yvzU9n2JKFcr+6XeQYCvG3o9efjkBeW8LqVzc8RCv3SEpVKpkhQLj0SAuBz4VPzAFwZLUlOBszWk
MOcHGoUocC1nwZyVgFz8k7uqu5a7foJP+JOtx/I+QVnE4Ya7OPjB7vB5JMapHE42AdK3zY0NtTyc
toOvgDPgLR8fqB7gu1/ZazhPbrqRO9q89PtfMgii7lnGvrucx5t2PPdbp+284pgVYD0odYeCpo28
UamBCwo6grvPObzXH+cVHt/uaJfCen+fufc12m3syemI+ivxObsQnaAtaGnR3tOCzMMOk4pNLk2c
ReoLNPY4gEK6xqtWryJVxRxt6y/saKW7+MsPWsngulJiYWAKGvIqj6ZyyCR7f+iHb5otWC4skkgh
YY6kWmuJHEm0LRr5RttTC1uM4IvO6v+dsAXnCX0TvVVgnY1jhYJcXhWvvlDZGPugRjZFaY8lzN+Y
vRhnfceBcktS7y2uAvzvENobWt7h5na5Hf7UI8RUCKfiIeAk1Ziiyn4RVvMDksg/JUNGmMrjnHWk
fDDmgOFslafpEWs/bRGUYTug6puE9flwhpFjQsXVGnwogQA12Wu7vQKtlCn79lsppz66CVijYM+a
rGQK9VQNZ+Mx5ytavcA9VUdZq5bzpMAo9s2DE3HqoSRhk/Yu7jrjXOqa7v7V7wIMWc39/y4BuPc9
yn9PLtfu5/Eue2Z0qhnK8i+QY36HWV4gxr40V6HVbABMcYUX56QvHCtLPIJHBt0bzBngWRZNYEtA
2GDyp3U3boMf6d3q3eYKU7JYAsGX8lEqocR8Ab2lA7JS4IVkqHCzIOFJOASi8V5+boA2I+0HedO1
beCe3MFYW31t/MHT0L/qOx4tfbwFNHcYEe9rzhwraPDVOzbP2/10uc0Bof2H62g9PMb2t6Yd3zJR
Q7KDJavQk0Jj+qvrt3mT4S59o6jeihf67z+ITvmDfyigNPncaZdjzzK1HuFEOikFFvGadVmZzjlU
5U/h7EWKKzfEBcw9AntixwztQFgwZ2jMJy4kIHNsj4hJElTXZKe+vwdEah1BFIy2Ij0HgKIgIRb+
owFsf0hGKo4J7sk4ci/rCqyS2RouwH8yPPZZ3mkl8XRJk+ZxFO7J7Bu4HZ9CUCf7mshiE2Jjd7aW
gTI1lN2M077sxP45aI9/jwpstMuMoVcymjJieo5qgnt2HDhGlEbNSIGP72Cq7mA5dj56VNXfbFfP
DCKft9aqZJzyGxqXWQ71/C+xYwn/pDi82gYwgtZlcBVJvaMajaw+FJ/0C3WLKJDFh2foLULaTk65
aHF4VAIU/x70lb9t73o6tsjyXmKW+yACxoBdyIIvQr0PmZiG4LBc1lmq6xAG3yUf51TZpYb6pwTb
13JT9OAF1v4ukwKfNu50YUY059ASAMy0r3lJVTp942hhMK5mOeXZDlacRo1UR80EQBSF8DfGUsfI
VPwGhFck+fXLTN57Y3YE2Wf5OcUOzupCiEN+xeKQQ3iif+j7gYt0bVY0zMD4gVnQAC92MUsLywWk
kp8S0Qc+BRoFL7IRgYvaQircgoVBvbwNImBtDcew9pgco61pELrx2fUIXBka2f2t6FOg8Alw33m3
gpqQhTcZeZZx8SmTwj0/9G4bapK3siIf6Zgkznb5IDPfCd4xbwLFrPjb5Ix139nbKb/CiSfWqYdf
FPNLjZtTfp1rOY5t15Z4uv/pSiYAQC8C6DZdpYp53WQhjc6NbsQbwpwKLf8GzQDfmpgjMf6yVJTA
uJBHJOgz6h3tZAEJ41YdNFdAqQLrYBVDOG1GDiLVjK6Do1EJzf74kNM187E8C9r/TGpITVdSisj2
beiyRXF/6+x+BZ7SEZ9trLWeVD6M9JvS1pAOZeo5EMZqH8B5tqPDsV7hftEGEGqC/K3hOrHC7ZdK
cMQTy5LDTixNKTlUtUe3oAvgqAqBFjtS+2i4XZetNxy/f8DCl+shIsOImgDwW0744l1bxQZPp1sQ
ZAUZ14LLSoLF5ORj7/v1f8YDtsnxb5wu3vQGl3DAFLg+suvQH3m7GZmWO3hb847bnmd01H0EBQ47
fSxMmcqlYfbQ4lNGmw2h0OcoqCiQODSqnGdxC+tqeP9IMdDnj+CyKIudaRsWYrUj9o74oTFmt6qH
qx6PUsFnjuJqJwbAFdIwDX+GL/XUW4QGO7AnsClUhSZp7iBMbi94SzyHQG9lJ03wLAFLn3AUvFHx
yRIv+TrE1I664AYQGHW6QzmUf0NT2aGapq0sD3nEfysqCof3FS6jaYLvRx4fV4qgPjWLkBGWAWr+
3zkrDByD2Qb4HwEieZWe6tsEOD/MRh2/ZpMbyELJVJ4kBGypXc79kgBzq057wpZ1I7GprI4OanWk
1YEcJVUQZZWHadDoCDqp7aVcYXSgRACvpCvzkpmXsfUQtLhZdhkAAX7llLz3sjMlqTsPi/RHjtgF
CtXH6byEvoNmc0FvyuQnVifLm4Klv8MWLiU3n8+5NdHdEMyk1uMm5v4wbUsabeq4BGYl2127O4UR
jVWODep/rU/0dzHl1vgu6Wp5VOLljnshFosATf3ga1u9D4q0wINC1rFiuBRcdR/N8dVlmPcbjqcJ
hdQY9PK0g4LSWmOKyUmldxwZP0+LPQnqm3AtdjOgYoEP1EtJpKa+E+x3GOuyCQcz6oWk01eL7mxt
e5OEk0n2qR9boo44z3RsDbypdBD6KsC7xOXNQKrec8IJauhbvrInGDFBHNn9A0UZ3AHUE863Zc8e
BBagSB9QB4EjGwlslAkaIkY/3/XQHTYkWhhwnzZ2v9p+s30ofvt4EmSPxSHQzJ5y73258vwr/qNJ
9gvHvuHY7+MKj1Nc48lTKTubjYMT0lkfj61qFoNQ38eDZWq5Y/0wBjI3jyCYPq3SO6zzEm2+yPII
FcAyQb5RWPcGNp3kBFHl3HFoiCWW4MjFx6kLs+kkoCxslioETKNSag3PAub0tgl/Aukq2jZZ/tBS
zf3U78mIXJVryi4jHNoriDPCB8K68hCUTjzQV30wvydBAKLJWELAgTydajAfUZLuUfiC54tkQNJR
dMcmwGBPLivE7ihhROGvZDc5rxf6Qi6Y/jZFI+bp+DvNOLwl2Bvkpbug1n4wLZrmYHH4qby7i56V
sVowIFnF57Skf8lbIN6W5kRGiuNS4Jmrk736ztddzIfjt+PCOy4gBN7cWECB4sSLpkOqGC6Ox82B
IOUGeqwZKSDrXuQF8R7llrFBWefXO/A7TY2FZYeQZZQLRTIXkK5MD4fgtaLueqD7nIvgB8tRIDX2
1JTQg25jdpBgdUG40Qs0DWG19HEobEysPVwGxgGyv2+plOp/5C+we0/vT5F3Fp29tQCzyy6gIU+s
pHkS0aYNNyi82GX3DY08tcVjwJbkhDYuhzexk5orsRLXGjFEAV3oTCrw24KnhO6YUIdtS10pXAEv
kbee69FkaL/MDEjgVqIWVbP3URwmd7psXRi4EWFOgD88UFzh/Fi9iku5wvsGQuY6Y5DE3jIam5YZ
KIosui9Qv8oZWP5JWIMFImASQGV307pEr1416hDWOTHJ7+FDywyVRUoJarfhbKZccdoDypG20IWM
EYcRIaRgviOor+yd6JcjhA98SwVP/cdHKbW3uw4pVdnkZJ8S9Da6FTw126GHFhT9khQYTvvh6VtQ
JyvIuqA9UtE5jp2BZFx8J+9GlZcIjrEifTwoGpH3QmHrVTx/FI+bI9Xcmti2M4DpU0BYPtXY+QKm
qd6tXhp6T/E8XObZMwWj63dNd5HuzBLwth9IQX/SHamYQ427CXF3QPZPbXHhFaACtUSRbqOZWAYH
rgeo7JGCITc0urxj8vW8JRkLNBuC6EWOndZyTgb2Fv1Vc/cC/4wkCXG+I5RPl0av+asyJtZ7g9ha
sE87ggxxeQGjqD4RJGBED2cHhYYOZKUPId7jqGCS3ezhbRhAEUe5R4TmbALJ0FBsMq4YWlAorLnF
/9kIgUjk2JkPu/Z0p8ioFOfmKsx3whddZMtLVvsbnI0cIgwIMeeAMIN8JD6AtGdHX3Og7hhBpJ9G
iWCUkJ9E3rwUbC2ywiTkSN3Jmn2M5I1sVKblxGvHz6odlvHS2ZJpJOykkQTCW9HsqwEbtCkM8Nq9
cv49hPNgzCQ2tv8I8PA7AjD1s5zB2ruNIrIpOxmXQo8XKWk+VPjyJp7avD3aA9x2t8MlQ5/g5iQR
6YG4sJXW0nRM3fgaimeeIdsm3oG68zrButQKPS74TROM3flCQP3XQZK5MIdJWpV1mYR0HKShrB0D
IJbN5s9Jl1IaG6gvP7CEiBgZYMQ3QnlzfyzZAgtsMFWDIGMzv9B8vubpotRWZKKJTInTrHPAZEBd
q+GY0LOIuWklUPJ45lGVuHcfVYZrLZVzbqq6fu7pCXEYdYFBR4uKXaKi34bwDly8uhJDaL4ayDzk
0iq3+8sinzPrwflFp8G3XWTvJwT3IBoN3BoY4sWhF/G3+lSgUFs/P6MHkKSusXhz6PrmQcdsC2ay
HLcH1Oj8oXcXwKVJhK9OJX4RukGazXFAN0EMfmjM9WXxNwQWJT2k9+h09iTtEVMZQkL5tavQLosB
Z/JEDJ8zCVyvxv7KuMZ5q9NFsXDvLDH+lxvjK2DEnavB5h/lcSTn37uZhYy7E4dV1a6rNe7DmD0C
Ke12p/2A1kvP44O+cqbaGoqP2lZIY1jFTjI56DPhrEJV/X16/o/hHeVvaUM5z44wSpz0Aub450vi
c9/owdWcrD00emwN5O2/kQrQThzQXmptMbCC9GiiOTGP5cXgEL2lCHubWMLE4WUwiZJY63S1fe5h
S+FOQWzLo/IG2Xv1YAWTuNQKJLSGZl9QTgusjfwzhCcrOL0P8jaOASkJju5havl2p9NfUun85mJB
UFIuTXzXhWdFPytw7FZMc65FHlV7xQd7QX29rHnutYEICAkXqG6hzfgqQoI7B1AiwkqJ0uXYCFjF
n2a/QveCPtGXmQ2SuGFlOmvrcIFGT+VNtwf1rVrXB4Ad7fez9UUZcwveZOCIklGSHGkkEOiTdN9k
iqn7MvClGFy6TRnXWVetZxPvhc7clm0j3adLZ4F/QAmCsEn3H0dRYTPFIczGCW/oyRmnsOlT9R3d
rbWGadNMXoaUaHVOyostTopGeQEVpby3xt5UTQZ5IL5t6gIqYvVgqDOFz6tbded9+dP5o+3e75Ah
LANg2p8xPpSgrQXNI48ccjehgTEcwE3wyejV8ZHt9b9azAnni7CHovFJHBj1Cm3np9h2SWT676hd
Sru34j43O4/N2VavvuL6qoFPPojaHYEHdu9+ROEoGnZ/MAUDruoN1Q/iS46NDwt6TQu/Pyi3kZGs
Y7EgaXQSDQcbXPHSzg/DgQyiOQcpiHL6xTahoGJKLnykr4jDczznx7GdMylFh0MAK66uKXC5eizb
mb+a3ff0VQGDC67CMWfBoVwY3Lmw3z9CGqyFBq2JgHGVz5VcWmobRAG08zziajBy/DuOPcAONvX1
HLPZVcia+rNbyg1OJalIzMIYk7NClcWZ8R8SrLbj4xVP/H4LR896rdvY7+mAp/fo+kDnl4s/lNJu
gi+FvZqdh30E+iyE1ion2cSqiDp5FZ2zNdcpm+5SI4KfYqB0YOyydsHGIr4RBbZSepUSSctRZ+Dl
U5q2sSD9cjkTTZi8pfuRzPf2HN1++lPcLs1WN6O4L91nED4sryUzMIhk5SC0fG2JaR96dj2VKLMs
FTlVSU2WXDNVfLT7N4UPKCCdGasr2A7DJWxPk+LoQ+rdQiUIX16B+/Rss90BfDSdYLFZP0g5p+DR
LWaLBdr5rg5wEIEFxt6y/5udQsJk1uvubaLtvyED35zJ3A+2FQx5UEd2+NFMQcr7NfWdw49pd+/c
CpGO+Bng8IWPBHrgCo/uuU4d7mfdqFwT7jynXOMxJYqy68I07Wrbtr3CWoR8TawJr1bd/bZBnJ4C
3ZQoUp4BDMYtX3BdX/gwKTxHcL+3ikJsLH6m6kuuQ/q/YNL2eiOnQqdF7hiTYmqKcMtIxIA/fBVJ
rpGRZ1H92V7IWOmZrdnnvINf5ndkYTldVa7SV1G9/DxHJTQMsY6NHwwG8GpnBJZNrDgT7pb82y0T
v68lzyQXe/hKLQfPR33Zu3e/g6Uh6S9nbNhtvzppOzQkpSgLDq318csIegVTBM3eBdcqjwzM020t
R5Nm6fsIDVxFW7oAmFfHYSVDGr+XWFqy3cp2oZj/3N80tAvps2VP+5WeCFr/kM3/q5hD29Sua7k6
RCLtW2c0y37upWO15gsR2eLR7jl9vGThLvuGHKNLETClrnzGRdf1wCU4g9iJrUvFLiYeU7MSGCEY
VOeYVQG7IaLm59q+jlwm8mbDsvKaAlR8eqGFWIItxpKOTTJEbjcDuHojFEJd61x4YjOuW311BKXw
qr7lh8iMkM0PrDjZhcDyS0r64/S6kaOmhDOgO8beyrucXoOjh/EFXZVVwAlNban9z4PMD/mhoaVA
9Nd1BymDwvqzqUjpeDV3cEmfciUxNqzaQAdLf4u270eFDWKfrd+NKqpnJRbW1UtJ3Z0CDIRZ2ebg
4tBar1DrQNLEHv6poEbMEcqZGUKq1jdtd8bjrphre5ySSSoVh0pG9KSGnv9kOeCXGsh+u5L9Mb84
COKPOUKWzakGmjJQWsEOw3McwHxvtK+moN8GDKTUbkAARpQVa7NG2y56USwJTrZjEPgOoUb8jx/R
ErH6cCb1Q7na3ITH7AktROru7ndirVmtjQmSEIS0brYwImlqQ3pu/9cGY8fMjZb6dhNF47vIp77h
7SmkGxMisE5nqSq6XBnoyALN+WGQIv1LhZdiiaCM1c+M+qaoVU52BasERfrom6RW5PCgPd2JTxvX
eQlZ7xZyxT0uh7tRx0G6MUcyLUstrtyd9RaYatj/1b7GjitureLYmlEjl5bvzkNvJh4nikR9pMcl
3x8/H5GroV3WC9HypTz+mv/OkCdN0wwq+Lhmquh+Um9b1E3lEatuNY+lTxCQrVW0jQN2K2Migp53
7PqCvo2v20haby7RSk/gzfSJEI1HnkEs0/Q8nTJX163zZc89O+CfZOn/4ys8ngkQoyqwQ0u4qYwD
5rvVYajJcVdcPj6weYUsfdeLEOEaj46GWANhvaeT7iX5CIEovBw2WcLhLxkv6Cd3LIIIKVm2Xj7J
7J8qLM2bLrHjIge0J7Ln50w+eDKe+twb4XdIb7SFRzNoLFtjHG7azZMhAIkAI9mKxzRImZOHWzHe
JnfV21auZjEnBc1ow05nU4THFDgvd8wYyj11anq0Mude8cgQMZOCOqAc2M+eIE3m2LLWliEsd+pH
5D2ACt28a527xsrtHtF0xfi3fHlnLjuYZH9mgovCpWYum+1IkQlwZ1KxP3y+ejbReoSw28ZoB3m3
K0I/igKrZwfGbR01q8w/BuIk7kvjirjZiF84Ni404N6ClbcPl+HJbS5ChRUB2HOCvpaj0zn05+h1
LgFGvIG5CbdXGitu0ejirzCBgSsF/S4FnVsgCwOob7/OqQ7htLvqd+KQOHKbB5NJAfs25O5Qdllb
zaV9rw6C9WJZGw/KuhS3+2uOQHmybXN5V25iADdtzVkmP3L6F5dCeTJaqljMadNSZ4gvKdP940Da
ytoVztlogNqEGx4wYd4aP6WWMLRE+spqVvB7bAHvvbuFGSJWerbTq78AwaEE10WE6IpBTEqdr/sT
W1RbkoiiAM6jGzuagkRRvopzC2N5K1xg4SEZKq9LQSvzutD6TSeqxY9lHESIyZsgNzNaEbWkZmDA
is9RgGG04hgN98gdfgfaS26UWUddzLRucHw9W8dgAlzQ76l6eBiabQQX2f6MHTCSZYGwtoiYYuDR
PfW613+P+2Yoh6tumMAqGiPqW54+Vd8Wj1B2IO8cOmDC8Igpjzf/Ykq/BB/kCzITjzTXgXafvV/d
8UKjKyqpmqObg84GIo28rVRNcVuwlhnyUfnDttWvH97RMNv/1oy+Zms/0jt8E9JG3TrqWI7r/I3R
UjsD2yJ2SreUtY0KefROiLTTJZXqlaAMtHUVgpiy7IrSTKz4GaTUfkJpcjDcrIDuiXx58h/MXERe
ZE45iZixwmfg9ECRWz/VMZtFYWw5ZfBhANwVA7FgC/oYcoJlbjGPcXCawKgsEvLU00V1Z5fSbR6n
9sDC2Zv5ovIbi2LqTqA6E2ZQERoUGli9l8ycJWvj0ggeqb7ZKTYbfbuTIOIdPzalgkcE0K1/B1Uz
xGhJ7OcCPQlPLelqkp8kZ38+6doitViPY8pQ20c9VIhhnROckxPoKqfi3rdwUGKauH4pPPj9UsTb
7NEiJvg0E40L5NPexLVycK/F1cAMwk5t+evRGqZA5IpuMjx+rMPp2DDVcI6EqtWBwaFM+YXeo0Gh
vr/1/3JPud4EbeIK2Xrep1dd5dQ5Q+i/1H8M5BzzizX39S92iMYwBVivf6uIV8O486tdRf7bhPMZ
kZtTrRnapp1N953vYzkwwf55cSZGxiAi4yQXCG6Ywfbrd2zsBTXobtsecRgtQVsWMPDn3FkLJE6I
jEWqSNP6l278GnGVKn3GCAEFknVATwbgKewbfq6poIt52rX7a63B5UL6LVfxoBDRNBCY32JQudCH
eMpLb6KJxOMuMcFTpDtT+lc8/8l7CnyhCMOOsR02w75SGW2O5zaFY0XeMKr15y/EkmjoAszzDcie
5AzIWW3lcMO2pyg63e9ZP1L1tcNIybpQBEwlkrBRawIUoN9HOOr+uNIUB1UTKTaF+1YNE9fMu2Ow
QUARQiVjrgOojMoFGcnlIFhtHSaxKXhzAZvfCKFh1mQ1Z8lQx10pRJ0q6O851KHFX6G/yWlzOUB4
zMoPEYOCokq7G2sQHvyw6JQMkyVWDE5MGgSXpl1/tGrYXY15lIXQGDpPQLdckO8jHUF87y1DI8k8
zZVtdAM7BI96ymth6hL9Tde/NOPQUJ9VTZTTMw1Kx/ZALBj1IxgB4rNsxvwoORsSyEniLkkYSote
ImyVhap2nb+gDY+5OkUQ/VT5tx3HTaOH+7HTwd/0T7JJIgrbk2oCE4RWrWDLjTF/av+t8SG5MGUQ
67+oyrmspGFbwLuhnJ1NlbDzqMvTjw2t8WZfzy6vXArNBkRWOPCiOHWuV5v0Lu84hu5QqrkCqp+h
pBMt36DBP8CDEJCWgUbvlwbF+hiGFhk2X1v9XUBxmgVtgnK2ZH/wjculLhqeajBNYUYK3UvYEWYW
FhvOy07gpZRHe+uqZqxmBOkKWim5eg1ohB8naqZRzgxheVdQ/R9pOZHP4eCo9svbw0uMPEbXakRj
tioXM+1Uw0z+uLoOFN+xHdZbLWLV26MIYLdcd2c9VB2eyye1bWSk3qex8xYMf9vPpWNPyAF0ffzb
F30kPeXD+Dd+ZGo4/B5ceF6xG1Y8aCY5lvBpB6ruTV/6njFbYiP6Z+e9hbKz/MtI06wiDYBzx8mj
LwcCYi9IMf0Kw0OZdWxknJ9bvP8cXce27auYaxY2uoFj8LiXjFAVmncfWlGjRY/bpPAjhCdXc3Kw
ZuKBNZ3Qq45vMQrK5R20RNpzC0KsyFVZXFK0W6CIFmiqCKujaKXY30DIKY4MMw427gXrOTkRlVnM
sIN2U3782HfgKBUtf8lFhmvQX7/HnlwJ6qjEXdOO2CdrrUQxJS4uQMEJquIHAP84ugtP22Sg1xPn
Otg0Zeyi091QQLgi/Iw2sqVsjCAh0TVIADDlSrAoddE+veZOFtnvAFPzThooOkTXXURgF3fJbDrD
0OzbR32/0wm2H54QwIlBhxXKR1rfOJoNHtw6/E+WK+A9+vZjwYl8UP6zTx68hoib+eSOlNp86k6V
k2JECqfZeqZ5cbGuvtJH3ePMHgHqb6ZnQbVhatpzujC1yxRmVg7ESCrQjnFNaXpcmjSpE2xau7dY
b8fkEgFtEQxrcLybvBCPUih2tvrocDU3GmCw/340XYr3hI3yFsELbMH+3cg6tSVHNqSBYc/2w70Z
XmJImhb1+HFoGJn3b7mryuf2Etmx2c/XrlhmtfkOiOV6mPnahDaplGyr8RR5idfnwY47m1rfQqFf
EgHTED6chZbI+NXBw+8zz4Cu5mb93kjGpEvEb/Y2Ov5VzZ28O83gaPDDP0ypak1l5KY4qXmg5nZv
z0zHijRkxw2HsB3vH4wDfoqbABVfBpCra6rl2OZbxrKWpSTDpsqRTDY2WFWxkAQWbHxWU1A539xV
LfEnmyIItxfrYiPvQ/eMuyMg6W6fnOfzHwOKXgTSZ9WQox49MZH62wglbgf3pN1GfF991gUAytoi
zCHwUYrkXPPPgdVJL5otawCodMtb/0usow9/D60gf4V/G2rL8NMER3W9MJoIJJiF9KeLM888ntAG
mqm9Ht0trxTK9v9jS0ZZzve504bkzXZB8owxOVfebk200zEmriJIZZd0we6+8i5/hwjbSw0+njkd
aUdTXi6WRTQgU4u2y3FlGvaCQOO/Ib2WiAgwSR229YxousUF2u/DhQRugYjDz77wn2PdQ+wQbK26
HlU6pD5HHm1gwUV8Kgjgm9JL1/jvQGp4zwF9bKE4W3fWDtZ06inbaBtBsKG99p6CB2umqjIbg/MP
qO3wS08byQ/EKK1IV+yu5bFgBW6BWv4WM7Ix6ue+Atw4NcJNsGdcmUXdjN5cxBeD1LtZ9RYk61sB
FM+OmesnnZfZuOjIEFrgG6tZUccr95r3ldt1nYene1KNOm2LEpW96T2LWd5pvPtvk5+Mer203asD
shx1AB3s15RbPjmLqv7vih+/OUEZ+QnjFg1k5YTGfXMDBqNmGTdX7Q7FKGjXvtBYtzfJoBIdatDA
osScgO0mrZXXiZW2Dwnh5c6/D4EZAz0P+ZIdPjR2uIIz9vM19BTbzj8eSdPUC3N70oCDF1fJ98V/
uxPaLX8Sh2Lu6KzjajC6c5lukRB0zNFKcrXj8oIyCxYNPu0EXs3V19xkRGVV0y/8OKM8tbqHj2mg
ftLbXyE8bABXOgVLYk1vtRlzxlJqaXRV1wk5LqBjD8ehca/pREh6hQa2KWWXnXzJD8GGnbFIUhHK
N6KtmbbfRB4YYghVl5stL9B4Ir2t5RT/+6GQaxx6WY5agulg2Mr/blVtIS20wLZWPOE6bXEAxRV2
xXIb6KlvRBoem5mOrobKbKkZVHTvLl8Dz+HxxoqkL2fa8eLkzhlVArB/fmXSDoeI2zrAYh/7yPbH
ZE1TTAtty3aRdSGJ6LWOLZ3dqz7zPfnT8/yR1CR6PWwi2uELtg5lzpNPaCBMST+xT5ywFy8FSuft
ofJ9DKlRBOOkymJnwxpkaWm2WWR/DIug29esAmCRtaTN/N67/s7uaWR9joUsBtI3tTYFMrlvps72
2ecCLDhsf6N2IgfwR5bqIFUsIOeUr6CK5L+tf8T7a2WpHXBXk83M5fLjq5mGudAUNBWlZ6AOugvB
01fQBW30bQ0hxkEBSeHgljfWCnn3x5ZYjJ5xwdntnfgmQkLEqAuaNsd6Dn3Nq9f/MgbpP8AP7Xi+
SSremOTEkTqwlDuIhWU45e+9Jif1HRxVfGymEk3QZQNFpt9JkjpaNTyvaXURxpd9hp3WHXvsdMVA
xov28dHcibGK1dzhum6VE5H1Up7kuXmUXsBUDNRaE/+qIDxczDshjeRStm0vTgoBpn2lWBMnPCXc
x4m85JZSAtG+266Mauow7ZtJHxpMYFq6Gy8XyCjbMyOucHKJStyb4G47Dy0YuVwW4CWIjQYShxQn
sCLA3D9m7WCoZ5IYrtd9aw5Bd+BJ8iq6YDKdN078b1q571VcioyhpaJB0nk6jEpEG8BQy5za5PCg
RIoQ7+TZAYBKjeNnE6JCszKCjZuWPkiYVDT5isLbO65Kavk8SmcAjXFKyLEMOVqQaf2A+atjJRfQ
TIG73Rw1PZAWNUgTz2A0edBoPyTqGqlmH9Qh0kdZyhf3zE6akB8xOT6Emb91Jfl4KLxSWrfz6+c0
1uYwWFHDnmWHy2XsPAnlugM3mp93fL+jMqEpxjXtxPD/nyPDcclrewxukEFFVqaPuvQoxbVwFgsz
vae7UPm/ZLtOO9v603Vnmbb5MKYULTCX15gjW1RJWQ9B2MRZaaLa2lm01ceHhDKspUh7NuFGIsub
s6wv8llfCrRAA27TcHXyaVK5bhjsiopvMaNHebvlfpkoluRCEEKiG5mluM0urAMd1ZjsL457fYF3
DH0kNvncwbjW2l9/HKmA5jQ4xx4eaWmzDnZ3gEf84q0sX979InDFFsGLwkkjhxUiscjJ1oiD+b2D
dQ1JRt7TXBdPXFrnglIHEmXJwqpf4lmNx9ilHNeWgP8O5sh0M7ZrMT7ZxQG4HVJAptL9ynCG8/16
ukUidJSQNtxSWTTgY8+nUv41fR3/K150f80KwUz8Ek+fIotLAryrcQ7TA+R9tirdamEF5Do9I5Tf
gPD0uEBRIHhCOG400WgIMLzBHbjurzFvCnbVxW0ZMwUCZRMeklHEFQgpt4gb6UblrqIh/wAhGEfg
pwvxNvxQ0Vsy0mfREenXqFfAZDHomwV1f6noA0TvKwRFGrFJ2N56fKWZDfzV7L8HqSrGsa3xOJ2k
RCmQAfre27SWRuSm5yHq8YyK03vE80lZFKiz/VDD/mZDiYHWquNPpKZNgNeqXaabZayL6m505peu
eNLVSZhZsbZAcvC1k5SxshjEPqY2/6w/WrXfhwtgNcc8Tn0YoCNWARa4il+6FdXdxIb+ooiBgyrf
1hMaH4bx8doAwTDtAkVI+klPApI9gG8vtoH3gnNEBqSL54aoQbEL3i9uZhIfW2OZA4sj4IZEU8sM
NT6iANdvLJFq6MWzp4x/MJl8HvfmgnwcgzhlGVRhbY/TOJB75yZaYqJuk1De+ZYHpNfrfoNwejX4
L8qbqbSLksELxt4RwIGfEromOiDDWkXmIh1sgM+Vk3bWYfCwQbicQf34cTbC7SbqmIBmq3DjDF3D
IB8VvtFsLzXnm7QPeS9+k9KoMwqwak1gSg30rEJfmdoRFZp3PkEO/+s7JCnJeNNGRvo2QhlC96Br
CZAcoiKTTMvj0i2PP4DGV/QNxHh4a0llyiUlFfWJG9IHytHQTs08ok+KaeIsO9djmQXgIbR6imsh
qcKa7GNEF2X4Mevg98VyEprIQZCR6vV10yGJ1MkDe3L6dsASeaIp55vfwwt2lf/Xaa5ulS+RaA3i
SgrnbFIcvPkep9xomjWtNjNhTtEd0U6B0kEwMgpl/SGaDS1in7WByseGBIlyLU+eGKfxqFCDjFqZ
CVz+g+VmYscxE7MLctfrYr0Tmd534pZxfhF2P5dVSLUd7u1tKz+ucKFHiG1O8exNmdEjAPaCt4lV
Sb9St0GYm2nYf/f9KG/rn7KeTl9+cOW4tdS02yhI1tHIn8Mz+3YXLBFsR6Y2cU4XIDlZB4Nu2s/N
A+bPpoKCwVmZem6iYbQpLxpB+O/K7PTsyN59wK0qTn2SSbNa6PQ5y4a3r3eyqe6iwWb6Mot8UAE1
PEJ39uIOo9X8qOMG4nounE+Z7fxZYQp4v6FdAd9EQ9TkUjlDVXes3uzTQCWYvXuS2l2w69HxLioa
hC4xSpKB8JsdHG+QnDG5AYwHAJC5escMo/X/Na9cz3kYUERouKwkg8Ku/m8iZYk2Pd/aeOj8YUkK
ch1Y2zB9QDw8g7gyH0j45O5w/qV/ubyD0+CUYNfXi0y4n7Z2Xh1mPTlPe6k0PcihMIyZTAMXMypv
bleLFb6gjFwrFd3N3HbJrbzrX+Q+m9aFAjCjyXamcMcJICG5qAGlwuVOkiVG5zDKqn8PmZX9oRUU
jM5YWJWgyVkDMSJsk/7ChnwFxK/p4HHjpanPyHVbf18F+RxREBbKjiKKE3CkGTM4UekG9cxFQTp7
2Ml7Vs0Mle1OymWmlOC8eI4C7fM2ZiH2wHjHwA8xKcGlnJhIUQ8h7WZ12rbs4XQsysTCjJHIvvTv
yHgPsTi0msVnGx/Cb7FfxrkZrB+ORj/DHhxbjd0cWWixs9zWaQjC+ulVtVX2LmncAHi3Ie+GprP/
u8m3k+sFSJ699JHvw2Qi63WwHEDwHob8glxFQt92luCh3uI4seUVPvO5a1dAHpw7aKpBIejyaDwo
4QIB8kntgD5l4sNR06ROifIr39Gs988KoskhVOgCJptXYYVgzAXs5jecJWz9V3w3fVaBjKyDHPab
Bc8jCIgFUbJ763MmeRJlJaASQ6btb1DNtkiF3zbR7zHcnr2pyaOil089yArf3XHrQdwTRwwpSuIi
r0UfATs1fQrZQpNQ99e6mYN2rusx5252j5PZa56HpCuthPliGOH7RB4ZwUM+J3h4G/VcRa42nw11
/GfKygRMU63/IxoCxX4NkEulMNdAJ7hPhJvWQI5UMtoWAI1zDatLg544iTJ7YxTTSC8NHtXk1VNO
gBQOtQCF0sf5SyVywWUpjh4EEfCS/XD4f4X1mMnbOIFsUWkhXhHJkiQb78oAG5CTnRMwF71pJSdD
mq2RDIes5f99XuYPTpv2NQhP+4pVKSsQyd9VAoi6WVd+EH6GlvnclhjCoiDTbqiyuwx39ux7ZFS8
x6YeX9pC1tKV3L7m8CyjMTT3xf3m9cCRUIx29qcRrqrzhBtFLpPwKCehFwxi8wJ1Us9+XvX1RTc0
mgY5FkfXKW4o8dhXkAIIZo6ihLehnM/h9uEMBnddZrrwamAP+J4qKQuY5vyZmFZc5s5tb44Q9p79
+8XD1BrDF0bgo0Sqgalr5Hm/IEFPu3bAnJDjq+bJhzUQ11wFhi6TJvrxgikvNUsOAt046B2xUkhJ
9eUKmmWqf5TaF12seKSYbOFAHxqyE1zBq8BJQAtBas6wjQtCZPVJXfGhdhEhfBnr+/0OBTHi6dtv
j30t7aAJBFvVV9w9mnoujXdrqQ+05ZyF8ZfqVTxyh0ihoyA/03FIOejMwA2aLRDRfRxmnzVmuCvq
CaF6YOe0pRvtwT/hBgG24yzTQzzy32a7hAl2BrBGysm+vf4KMoRmwMT00qx+Rwn426qEmooBniv4
No+ZZovHLnTFCXIC469qsh8xgyu+uHeAn7gp5WKGHvcbpax0uEh8L6j8P+MwYjfArTe/XokssU7l
Hp4it+6ZskumrNVA33pDDBvNk4CZh4kwfrmZHywPiaupgJ5AXfCgvOVlcoWLRhwie/OQhXxqBCga
cjPyGR901HgEaiVhpWtP2SMkdc4Y6d8csAiNaC+d1extEyftgFY6rZZ+BHHJVs8xoylQBlSojOIs
L5r+OiRhKXkvQNEWmyewlL4kCG+T3n51EQIyhfLy6GENl+5gzdSGaJKB0BaOERjf/dpAzNAbSpWK
nOiH+yY631ZFEzDd2zry5Qy6CzeX7K2kMOyFAaJTBVo3+muqv7NoImwUBHHuGfNeux0VTW3d+hVH
5aWOQqrNXd3MKwIxb8dhlmEOVkdm/lo+87sG+IgIUhbcJoGMmF3R/194ZH5hKZYUdduSp779afxN
ovAcx5+I7swp6/rgdc3/DR5PrZQT04hxUAYdX4GgiNoPi2al7oJd6jvMxdAT0WLOia8blwo5MHCl
jvbx4BwQeBWO8A/SOTZG3AoyhHzLfxt3BeUlX52/Ha9J1UDaeSiLXpsNsaRoGJJrrN0rQAJXa2Q1
aMwB9Z3gbmLAaDr1Oq15RvyFFOCp2yT8c4xREo8OGYiBHTwuSdQAYDswXWWtSSchzdC6g9mFH3jL
kDNmJkxF5U4k3V8Lk5wk65wtXY9WwSZpBNU0pTA15Au4C52Et7atBu50GGO1aJj96CdpjdYGqgzH
zLsh3dcULjjY8I1dfc7eBVVyy/4FmRukmMVls4ynjxXug4OtNNzwqGIDQVOd6D1+zsHLVj2Anqir
GSL84eQ3K1hqCOPf2eGu2hzz5mttLXk1oVJ9VbasCvcngj6m+VfmZKujSWJyn/eWytAFFzhk6NXG
lBETJqhAx/ryTA/KrHYdqiA2qwPZ9GWATdT4zwe92HTDWMxRe+oqF20cSMPxQAYL4VvxrcugNeDb
cP4jfu1NRWvjB2JunZ5ZldP/eUeRMiJIJqZU4hCvg78ErIT+bBR6cW0Q4DofdtfeKtbFvWshXgW+
1shT0xIyYHuEwY3McPH4iR29FtAeioJSsWa6XU3Xls89fvfl47c1K0kghH4NUxjtNNKdTf4n1g5q
z/DdtCefim2casR9mKBtbZflypKAtxy88r9vD0mioeLdUlJ+JiEHWVuOKvApXwEYQNGsU66OfR8F
cUhrFHJMjMdDiUs9D7uWcAJA55b0O73WbKbKSXdzykgu3JeDLHEXaiZwg6NadNFLoeKgyCuezbXo
iB7YKPIrWuwyxZ+TkIiKPmbXRvzW22R56H36gQRIYDh/MEPzy7IfzPtsyIVBNcQmZAuKYanqvWQo
QrZ0QJw37XNB8ga/GH1UH1huY16z6KM3EvlN9Wg8Bn3pCa4z2iZRNNGuFW9WkuAyc0RGX+6pxSxy
IapAoauBMNjUZuLSMHlb13biRSSPYfXrUsLwFoh/xp6e6zJpRZOkQiI6ca1pC5aQI23RE0DwNzco
w3zD02zMFcdce5JiX8FDIdel1oMz6LzTYxBSFm7IX6QxBeZKh1T49NQFQZdvYkKZnQ7BzB3wyIEQ
avJ6eYOZhcjYSoAJcuLD+LTFQIzmwBdMZdIUjpxlKGeSOBReoefLFZvMUUl6Zickeh2UWqE9jjoz
f70HX/y+D/bOpm+1+Flo59XOPlQxL9RytHTfINlAJEFZBnF00I47U4GtaLlutealp9TiJwd3LBlO
hevGb9vS/wdGkaoyZxyJx5t/OIEkywP9IODaXg5ZOUWHZccC+cpwEgIZAjY+TuS4Ofw3VEqfW5Ed
w/pJbHu7I+/K1fIh0AGujkrOhT0JTlwmTFxKSt3SKV5pTezRg4v+Qjufhq2cqVEd/0mnnqxU7nxV
vzBs5JoneskgsYu1ZcKtP40lYMCa08V4UaHq6++kExpG5AjCFeR/Wsc7/jvK7jCikMf148ArNnn2
vEkocrqO8/SVBSqMEscaghBU6NAiHrMb8m3yGXvAXbBp2d3MiMLcWBSHddXnnsGWG6/oP5TETJOo
7vmufYaj8HvHAXrs3LeuSu86vavGwYjdax4AjyY3t5dUZDcFCMkvaTkQ+89VWwImpd9TUnCEfa0Z
Do9CCJLAd774TpxHTmbvSOaE4Qm9Mpwivhx9KTXvS50aYods/8wNj0h6xWvJJrl3XHhZ0pEk3JRZ
P32WyGQZ4bpbTkomCPOVC2pepNhvHoDgt5PYFRdfK9Vv4SVnyMFeDqMypQm2tiv4QnABhCoVyaJq
hzHJAJS0InM3Uywd0J/uPaEUG3CHKgcl+L4kYFcIFhB2D4tHbaY65r3aaWo/gUWvQuK6xHCcmwsj
N0g02TgsGfFq59QTetWvcDps3o3Jo4M17KqYspfJAU+SdCQWMvHOZLL/7TdtdEFlWvoYa1HqK0Zi
TWBP5CxoTLYS9A6qUg8tyWnviVcORJV6WJLo6GXkRRjA+zBMFXcWuzt343E9aBRmVkwQVdkaRizz
imG97ZKWIzIj0KSj5dz2XMpjKTyTxS0LHc5153iySHAkhwmk/TKxIp1qGIGuDfCtFnJG7hGqv9lp
zGSvDK0I0odKXU4KbAR1ugIRWJVIzBJv51OHr5apglFjAo+wOGlXQE3YjSkjPjNyE2VD07+tJqWh
sb296CZarI/obEun7H9J2BR+5toqttd3NEfY/1LmPkFS94LIYByZ7kAeMm2PqVgAQ7Vnqi8Qtt0r
n+wExGHYoLkeQ2z/VTpODtzZZphRcI9dYWK5/aUhvgrtz9yd2dI7mjgeFRTp+lG1CGCFES3XA9by
Pfgn8zeKGW9864b03lJgTJjY6OM9kIFrRVQiBkoRS574iEh0GWEGzzpMYosbMibGAcorbMIRhw5v
um/m4jA1FfrrqzT5oy0/nBQ3i+/9W32OkuArZMgSYAr/9b66OQtXLl42y9RNQsPFWgY97EYJoEi0
0+Ys3lzctoYkL/94aHCTXch2jCFgfyZrg4KUQcQ+POycYeboWPDT4qHjWPKDKlq+9NAU15spR5J/
dCX9tndk3w8a3TCv8Yp7Z7eLot/dh0FV/eVKLrd2DaQFRqPDg1trTUNOQdametj29HOMtqHrdZSo
LXfMCvFMYvvN73Ywo8Wjc7QwQQqTyX78WQFMO6y+pzxJmTRbOdmfm5bOL68NnggluuzYk0LJE1y8
CgB8xgyWsFNajz8uusyyQvVvIYB+My0hAIKFfX02lvmyEN4wh+/DbCQznM7Yp86iT9iO43XsBsA1
QtpiVXewLAF1mzHCixvNI2dKHbTa5eccdKUhaXTlfPAa3UtxaeOljw3IxPYTYQhYQYp7RP9VoF1S
qMMi9N+6ZEhh4UXdn6nTI6Go4kcjFr8nUi23jUWko+s3yBfdZRtpLgp6YoTyWKjpBMa0gpRedCQA
+57B6KIwwXAYNakeOqjEZSQy0QenApgpln7Xm2Il65nwMKlR8U1X7YMoGjXRK9QVj9e7gPgmDEMv
L6PE2heGVxCLImOkzLRi8gTOg3ghv5o1ISA6FfKdlu9MRIROYiYKxXCkoqABA+H1gZwQZ7T3Hjjw
ftpyk1SUJlKkMYgi0RrCp3Nld4Xkyh9ab+Pzcv+P6ctsRU+gKIntRKz+ODCQ3cuuhVZRrvG2z6n6
5XQ6WrGNzvaKssxl7CYnjPpesM6mZyH54YhH5MH8metqIzlWQGdjqsf91rhZLnC+zUr4yNLDCmrJ
Qpn1vxLNJoJSUZfBma19mcymtOfdtnxc4fA/lOzkNQPKl3JBb9cR0jUL09P5aOXo3yiUrXU6Y/gz
3qzAcBmv8sENCVBAKRSuHemcHKmEdqQGxzsQyo+mpjOIV5ihLNZnVJwXuZOE3GFS/uEOiR16bLVM
eeZ+gqzY/JNYMPcqHZdkfO/BUfGfXsX6FSXUQaNkWOSTJkQ05IbfafqcYdD6fiSWZn4otJxtlvEk
slxCL2/Uuey1HQPRj6/9JdyeAzhaJk+NmM8dz0/e/+7fI2Bbh9W6NT62ZH+noh/KQyH1YkyTsu6z
upFCe/2Yurp2Ho6oklpsC7uIR43WNQZSyDDIuInE2nQHydmtzjB3vJOR2dzCXn7wgGJtbLlN0eEh
KXrAxRqmCBm3+fX2vEAi+dD/lNN+DKry/MMjVFXdgMk3H8iMV4lbjPL8mwLYka5WjF5oIzigVnaJ
PaGVcLOeKdiIevW7bv09VCc3FCBDOLYff1GKsxwDr/jqSXp2qfwWcUVV4F50VJjAsFxXDhM7ExZc
NXOD6r6IsJ2sQieBlHPA/RBh90dZ2EhPcPw7cKzeA7ykgG1/SjaxMjOB/HbJhiW2aDufy6fK6ukv
pV3CyRuLR1o4VGk9LZmocr5nA7pju18geVzZHajZspQF9n68eWayppbCgxHUftC9liRUKVbaiA8q
eU/CZjyerqzK4SSULSSeJ2Zv9lsd8LIygAH2BI+P1XcEcNk+ijpvGL4VFtXMMfz1QG1e+rNQiIdd
bKlZgh7f6ks781+IRAbKMBV6K3FR8wXU84RJ57J993RS2BlfhV4EC+zHHTMwbfk/4gNSrC1HWwwA
NFqmcZ/abubCAzmFgu+miYVHS/+VzY3u9YgqyZQp6AOz2jzY+ZOoYZT3pTwM/vW9gaJ0VMsGZ4Ba
ZPol6SQ7J0QFAjG1HiYkFi7OCx2F6qPAl6644J8nPJrC/iaO92oqvHjiEkk0MSIDYI3ezhDGoyGC
SOmwUZ3MNMf2doiMopjICteLNdi4D0IlvFJ533IvjCUyq2j6jE2IbssPYChZ80FfAi4fv0sa8MZH
hfoCUEMUylMEBiZ+hQoXm1BEjElPCKAlxRWjuuz2CtClJILUmEgJ3tc8Qs668j0Tsi+bwCZtA/0h
kGq7IQyqbFFpdQrUqW7KY66XlISdYv/5I7lVaiOxD/FhrHOzdLYOWHUfseJgNz9dGEU2E00xm08e
P5blYF1JDx4q1fbBr3UIo/HnIVSZv2DlHVidJdBF5HV1vNNDDoGpVN6NiHiuZWSiRsAjCXSxdzek
FceWr0B5l9wlO3rL/HLReH2tEHjaCq/5/mJ8YE00uO3Hced1ZydRZR9kgFaV177u8H24QBYdzltj
Ig1RU8qk8Mm9MSM4k7ZxzRzoaR1jsncUcWU33yH4SeucwaFuw5bYU0BPfCwcVolnTUnUJDWErvZw
i67wcb07Qvu1uiy5Hx5dyMhBmI4+hnFwGwkSUNklxN42XQ9Qz6NW55SyPN52FNiDX2T+Gs6VktTU
r2X8RHE/kr/wP2s3kJC9WPCveFUmo+6u6qrm3VvZdFYo9sHG+JeOtUylSzblRcWiXQwz62IjXSIc
mKFL6ubR8OAxdLUUpU6HjRYzxXTHI79fz0kVVkyL8ufnlilYWKiuxH0oYr9527+x/j8tYLWtl0mg
aFrwy0+k6J/l1P0abA58ibe1LqCptD5NOnl2VHPghR4ssmrKuqlySNg8ConQYllhU6x7f4PJc9+j
ELjfScbsG92L8VY23pXoLxY/b+m6bXEL2iBVzpoWqW6nlcCUHI9D4iS5FVp3kenOR0GwS08xeiXC
fXydK828cENzbFoUxpPsvBOjjE04dPekGk6igF5aS8wy05LUr8F0gSjzo49mMJw09mBOHWXKa6Nd
YBMkCohasa0i2OoZkMcMTIeUNIIX7JcWkezcVnRbdSA4DQXBJqIsm3XP0B6Pg0RCVK5zYwWOCyVQ
oaU1SvaBD1KKUc7lcicwDsCL+M+AIoCAyx9CXcT5Rx8GROoPsjpx9GwvjZKRFbvWBayhVkfOTmYM
zNN81l3yR1LvPXYD99KXSLucc4vTf48Or8JOrEVKzUosaFHY/x0nAevfu03jn2PbgjBzPr3s7fxS
FGi0+ZpyVBNRkT7Ba86YG3oFDsicXqt3zdRr1PF2JCZ17nM5ZrGQwU3lM+TG8yrhZZxdzcPIzjMX
PTNDsKxUS2+qPQkz3J+3GKGh87d8eIn47MCcmivWw7X2A8tpCC4fhxCVcswS/eU3Dssdim0w6xg1
/nJRNlCjHrWf5Vx3A8bY4nwRd+H1k9SGoq+PKNdi29u0YihRhd2F1ysbxCmGselAflx7uPgjaOkG
D0UGyO4LrQ74vtezSP2srmacEaXq4woCQ2xsAEbYdMJak7JQ7xz1u2qjGbC/ba5pYveAQnoXVpLo
VFf38otkkOeBBpVJRwSDDbd767og5R7KMBMQ1WdH36hV798lhHjhYPEDF2LGlmg0Ok4r+TTroPED
YLt1so9qK1LTPRd5Yism520H6h9OeADJGV/jG69qS39/1W22S0F04osR9esVg2BMy2kvGkZBp0yT
5iojEyWENrYXbF73A6qx0AzE3iy0XVjrAAtRdERrHi5XVTEzNABtzDkOQIAGdJcA/qFkEH8QLall
lfO3gEo7GnC7fJLS6+IpoMHb7WB/okxpGJLmA1+h4JCn2zh0hZBmpN9sTe1QiAmEpaI1y+oGOc/t
BxxQ5GhQezuZ2xKg/w23ituaLGoriC9+r7R9gc+xFIILOPwGalr1O1UcCwJrPhlmAzzkUUzcVnrk
v4GsbHXWiT1xn4X5/Lc9ob2j+dsrYwT2MkBJJAcDWIPsPFmRmDs+DY6feUrBiUHn/vvqgr6GVjEu
Jpx1jFLTTAh4spBHHt/O5CM8y+qph1U/zcNWTfn1PKSPZGVoforbU4mL63Ogyiz1nZJ2cde4ZRjR
TuMD/FpifRpayk644/Pz9LsJejR4tYuw34SX2NEurlKv4F1wDlGpXCrmwaKM74t2I7B1u13C8VnN
P+wmX1FlY6E9MloyT/dXnZx0fhwdH2r2R1uiNploAZgfH4vyTundVwuIuknbyEiVNOemxa5r0YNo
63qFDdhMxbLrLNf8rS/zJx0CaGuVjXMsfQE6d9c7VVk+QoZjwO/2DLG6pmNI7HBhLmEpYuO/4JTN
c1srSBlUi/6J5Evdn6k8SziUIaJk3NZetKZpCyzAvLKGAKXd38Y7We6Xbraq2LmWYbZ6ljeaEtyh
HLNkqfNfQZiTsTd23GtUeEhBIBDvTLB8lqZoqUn5cQ88avI6ARMf3K0Su5FLmsPBK+5qgOcRBYmm
YS55+P5cU1CTafFEklunusAIAiA5E4UqgvJw5VItnRrMCtz2jjV+CV7jpN/Sckbjrc1DrP/oLuus
rlXQqM7n3D9QhJ6ABxsIW4OJtIP5GACMbwtSRrgd1ys5S1Ce/TsfRliYCtrzWFqzJ7scGw9c8saG
d2HKyQIhWeqqqUDohK4SnewsBdHQjClZXXknVH8aeiXRv80hxI3TzbYeHlcmRNNX8EhrMV3LB2Nd
N3BKoRqMoEg1UR2guDuuu65Zq/g4ZK23phWaIrwl1uXY93EgjnWB+INwb7e18y6M4wh6sBWl62I6
v27jG6qaL4tBRW/u31TpW6Ssrx6IgBbCMOLMtGvpurxYKSAJRkFXT30tmZK9GDN/JHZJTK2VznlV
i2ifehu4T8voxL34yrz4wHosKyhKMFlLDzoOU2nBGDnV8afzNio7vwi90s60PYfA8MAf6ZtKPsdj
PMqlVxYtXAU5KRl9V/ZxsTqmeF7UZeaCND0iiBYlmis5ZciBStWnI6EzbBisOxxmLQiQd/+tamBp
ycvX6dtc2Fxd7XTrasohnbiyBRfX7D79hUrrMtwFWFEWyQf0osrPp/SW5NHFgw4UQdg1KxU3p9Hz
waWEjRlGelkY9V6HbLOsUe6sg/ecieWYZF5EoZ4qCNUVANhX871/wjn8Jlv6A9Ng/8FC6hxWnCZ0
UE66KpcbF6FCCCj0A0iMtz4kwB5yg1Ay3iZRjdAjK/akT3JQEhgmYDAktETyI22tRu3bXEt4XssD
jFN0kigROo/StxT+9DHPxYhlrgSMlKR6pyU2gyn55HDe0o8f0THL8srI2Azep7/xzYryT8l7sHM4
Xlz/TNSbkxZGjWXwc/7iDYXzkvu33bUyKPEhGhoWgtEgFZL48Zb7GeBS46EVfPCX8hixxN4mG290
BS+Ww4+APA4+kITQtrTfOLd4tNkeBVPvD8sLo7YLbg6hH8I1yGsXvZnpyGs97KIjjK58NGISbv5a
/5lwr9iIyZLx+3NTunRaPjnA0QjhZxaMu+0w8SWKAP/X/3li2fkTYI/xVZDXiHsVysdosTa91CZ/
HYP2PCDJSZkNDOappkN+ZZSJmMLZqg4Z5l91qxlAPSaSbUtHu6+MGPwZp57mn2rX69olBWt5ye6k
1hrQJr2wTptsyXhggbhVn2nFP12NW95466jgqdBnryjjUQaT5Xi8CIYNme75i/ehYW9DajuFymmA
9I5VyRGjyduaQJfECzcxjKiYUO64jdVG6EJtBXIJL0qBSTBZTwvaM8Pb/qLhTR5OQjBjTzYhqWdB
LoB3Ct1paIS/KKekD+z7Z7ubg05RH7o7Y2pU6nc+gKh7HkgXKkku101aMZx5XBODBGgf/eLMY+CQ
hMF2p3AsqBKyzwUtOvNemS4e4I5649lZUgln+V7EHB1vwIjSzfli9qxXX5mw5Ev1EEgguCHBVmH3
ymBLYqDh0igUacU/4YSnkA7NoWExIPzJDpI7oLa3ETMffa/FuN5QRUoC4Aryy1t8fEfjnFk/7gWc
Qur4kvx0M2iFvJARLl1L4bxZMgMWLXdY1TAbvU8MjE8yPH5JCJILqNqAotWofppbPmHEfcnyVUfP
E9/OTzE0qd8P1aiS7g9ADcB2CGlOdLlSJlMaxQtdUarbqtYuS1PISNhe7/BzpxZZPlNEUBqvP+py
y6NEuW9cjV8wdIIlLVdi3GTT6LYrvyt7p+0Y91CjzLPXwzGfpz78iqWEEcogAm+o9rxSc4W0IbMU
4Z4FV0R9sS7tI+npr4ZhPZLHXxszXNl6EXgKSPS9lpp24eANtC3H+nRVIRoRWTiZcV0nKIdB+qBo
0e3qNDw8Lwjd78vzvwZ4aBP73DLUGdnbH0p+H9JPSdrjEvyWFT9Nr5ejbyjwqJcLVQM09DLG2Zxy
jovdwb/swHIepE30Ho/2wutlXiA02j60g8Pld3JqNIIp2rWPHoSZYn0P0zj7HOP97lidhZ2+LdH5
qRv/mj9ZA8ytjGknGdUD6ymAcWsVYYB7+7lUmpZsa5kZJtMEgrLDgu/tFtV83NugxO1gBKmTbGQO
MWaQvDAvH5c1NxcbwQL3RX6y8gz/OWL4a39jfCoEICxxsCKO6Xfvc7iVqFKytDyPnPHKddD0zo7A
tSORNvHTev8mx1unjdFSltO7lDXBZuYnBWcDF7e3nUzxnbz/SgPnYwhAWpdUaCD0t+logDGSNSEW
Ua4m9jILTa7auhXu2bcMpjwGNqzrHIysHu01kpDka61CASBdQ4hx800rhXVLQB89LN3aqDavwgxi
RxVOkaUTJB9BiOkVQw5dWWMgtDOEr1o3ClkgSL+/9LhjfgtT335JKoCwJ2r1vhmYq0R07k4ERGGI
cfpE9WXmZ6QUJ4G0/W0vYARKEnwaTRhh5PC1sT5X1zrUE1HEr8i0aoRcBsAs8Pq+jX0O6d0kgqx0
BObbgZBu4+CsNR6yGiZmNTe7aboYwkTD6YDlxRSTISKf7++7V0dtuMIdc7oTvrZ1th8nspJAPY0v
kXBDc32vrws/vpn+BG1BCkK0F31HTymJBDhTsGyKMcAWATuNJ3gTfpNySIQxgshdByvINMTXLHmv
UD5BTPFY1MhxDYJaWAJxjjZVXsHS0TMktDHbm6hlDftOz0od0Hey5eNyz+PDusN8sSt7+gTRNaoG
LzL883rIuEo8CqVqvymnQjH7ohrN15vRdjOYQ7ZxRlZfis29m/GXnjKqDgcrr+MpDCBmB+ym/oww
Ygeijh+K00X+/P5PiQk+bu0Vf/sy+rybDwbmxpjNmVzoqm/IKCenJxlvLEjt8b/A9CdZ4UtrtcFE
0am4Oy2zRRMHRmsjLOmIMnQ4pg+2u0n0al0iWnUzAgICSkHbYfXfNNMMxCOdTuihrBkrjOaG5TOn
eCeA/YRWeSLapLdckIUKh/eCClaODjVQZQoRYlOXIqAhBE74KA8ywhI2wo5UPC5J0gTdKmFPKOfR
Zd8uHVuii0Sn5/ROZ5kbYchJWjV2udcE90ocH5CWK/LGgnpJWLwpYIKYqEF7VEfjmKv0vubN/X28
/i7BIb50CRHc/tqn6tB+2ycIIZLBCZY3xhhcYH31/grLjrFm6g/tsdSwEnRt9DRxNxXCbW6s2yDD
6G2vwxYK/A6M7d4iRkQXtDlKpHLhjzp8DAeIVqAIv5hc1JCXHfriDZXtDEzVleDv1MCKNCZ90Atg
4ryamfOqAesR9Xj/ehomj4T1lVtNtomhOq7c3zNd28I6dKntPpiy/uItsEz5Nc7eBnXdPD0Ih5lD
jPDODVxyg5nT5kJnb6sPogbLvnlDMQVdGefKE4uVbZ6lp3Tdb6hPX0RiHUJgfovDHoaPB75vkVT6
ZVhWzts6IWPa7Ek/sDO7qVJvQLOhPtSg0yLhcSAvyML17+o6YzlMzxgCitsutWE+cXYlfoIDrML9
MKVZaCzGS5vEms6hzL8D9PrFH/xvrk+4jRIfOCuZbaJeTK3Ki07u2779PN0zj/3zO5vWNur2vxtb
3/rJY+qduEt7A69pRqQBYATGgaHerucSHa0AYAHSHCFhnwm87AP1WwoAaV4Qgq1htE1qx+5HS3vL
UocfusngD3UmB03aoj9Hb/mMr4nri0M/0IGz70nSq5dOzURQIC1CGRVbI0A+Y0fWULs1GApPqIZg
u8VnTDRxODcZaX4KeutYbbBRNWT8NvkuPQgnRpxqbFe4ZBdpI8vWgpP8umeGCBH86oxYIfLWKHkD
f6cLghK1TogXDoRENfZBJ7qstnZZI9AySnm1yUZj8rC2I3hhc70QJ3CHZekohPCY0RnTqe+frTza
OOu6JMkhE9fv0TuVbTtMnF0pWSMnlIsYKszS4vOk6oiQS/68MOg1DO5hpN15pX6R4WkwO9lMWdZe
76yH3/NffL811TxjkkresvNEkJ9BXz3nsOa69BGVE8o15JK4mgO/Q0AUor8KuOk6agH5Lj7Iaqwy
LeNgTYa19tMsS9IZ/ix9emo9//NmhYnkkjKIDZwemDmuytZ+SP2qEE5B4mb89hJPyFa5mhmIIAlX
huypVrn7jCo/4DxQK7MaVGrl34UGWB/vUE1DOLjtmfeZLWVVlZ2OUkhS37j2l0mbvVrNFyNXXEM0
7PQgvSAEgQpycqY7a1Z8R8RFDRPuq7ECuo8KQ+rAJw/Z5xsxxXMaPcspLwV3h2QTDFree0HKvZOD
BgJ7uwv8LhopuktNG/QXLD/XrjnydVwH/nJPj8ZZ7SL+mYF4hrJrOVxLzUWw13XjMNQNpaSxVl+j
SPL2QhECH3K9yZFy6xODkSSp9fyiXwqE/01AWdP1Dc+hEmcyH/u+I+c5Nnv+kv4IV1tjLsIcEwpE
r85McRk7yIQkPjPqMdX6vRCogYRHKCR1b01o1CrbLezHoHgiudE9PTG2uEIJkfnHS3SrxqoBvY16
HlBb86nPvfUEMtqbd0TR9vjxzYRHwx/O1eRL/tXQRe3Cbyq1jm3t0HWOz6g/l06Bt5CqrfGY7JU8
Cd4DUehBLLZkJt2dfzedceHnQLMvAlvhkbZ8jF7MP2sL54qRLrwyx3rZ8xlylF9g14UurnFw/TkY
KKRpm7KowJesX8MqCDdvKxS2kqu9O+B0ompngYyiYsy/g69ww7s/Y+yDrPO9bLpLuvu0j6d4F4H0
UZcy4WB+mJCjLmnCL9gmRuDdL02GhWilAuyEoo0Y1ayw5uX0RZeCv6L9r0rWWy/oP2XXim6yjgFp
wFE33OhuCE+sWVJAhcDYWkc1rUIOgATDP2MHXeRZlp6Wc5tGm5eNjsRfyRoAdhMkrskNAb0ZVreU
w/YKSW36ddk67F6hgtFTM1yk4JGDueoAE42V+qgMvzI5RIiDmo0TCUMBA07neGHWTyRfOElnwyUr
kvjfWoAq1NRYwFRjAs8M1hyfkPmVw7ipf1S9fzkAQcFRkjsL6zV5nIv5n1KQUHKU6ZOUxWcrhLx2
oHXLnULLCu0tCtb6606/+rGQajl2uNieShOuEeH0cPVxMCEApTQ/pH9EuquppI+IW4BZZAoy8SGr
A5OqopgkG1qT9fjHaZqzwiQKq/mSTy7sA7D6oq9pW0YD3X2HvO63PEh24ADieQgcbKO6Byz/mJKM
WIHrgwK27Qn5ydrYIsyivk5kM12w/CWYWxIFL1qXERViThetnfBsxnBwAvK4h0cyZlkIGfSz++8f
CC+1fO7inr/bFt1Ar2BsEm//rGIRPW3C1vypRXmjal6s7N1VmE6YrDLLPYrfY9qlbubVymtbGCYp
7ltB9+FrKIqQYLRDtF+oXhZLksL6wMN976RFOaYzXvCt4VTzJ5Fw8qIoM9szvvjaFchgWP00HG0y
p2Z1An4Zvh1VR5unLuX73c+2Fucshbmzvx/mlZ0TMf3ju3uZemhDA+fjbt49mXsXU4CCnY2VYj1R
gDiPLmjnmSx3VrajnBWuNj9dTJRpt9Dv9UjeA48rTT+gqjKkQLymKm2Rk9UCTCzTx2SBgXsz5vN+
IRunUOpYfiy1OWeoaFzVdwej9ooIPtekPG40NyDQJHIQwcnQO/5gOlZMOAypRglXOqrNBlR9yqhU
c4HLrXpp5aSNStPLGireCb7G7Dags78fwZPFTbJYFqG34WxLvB7VJQtIhxpWyvMNpmV+E3Fs0Tpm
FsK+2PIMO79GI4UClupI5rFU//FO1M+opXRshRJHlo7vy1jG94zBD8ZX7I8WE/AceWbYpOPfepXc
amLYxTFBzJ9YpLjQPmqxCBRKbOvEG2+LwwcooVyBWyt2ZyMNYFFT457h6BdILuLl45RawLIkPgQ9
kZ0Bmjy+vkK7tkuUhvVzS+xoGRakSI8a+ajkWSVRf5tUALty9+BfZ2W7ZBHeKgKm+AVkp03y5Gfl
OFy9VCj7q2iJVbmhSQBT5AzHLaoR/7uIGe/rU2GvRqiPQuH0CljaqjAKQI8EPsid69+gwVqDl77J
kTZ89Wpyu09mhgBSdmmra4NAZF399W+7Dn3LXqtJmSxc2aWOO35mcDjefySdN011ItW8tHE8bG9a
HxBioWa5Uk6oCIdqBin8XHGBs/YZpBPkki/KoYkrhvhwXCLkbx7dpHWam3h8JFlRV4x6FrZPepJO
VYkMpzVSAKJRZ5kfqVAbMjplnZ0wSZHQyuYn5x7WbEcE4nfjl+sH1nLbYTbvsRYIP5V/cHH8EUP/
dZtV5kDZel2Yc6ZnOu/x9+dCodDGw6hEY7N3JN6MBPXRSZmWbyPMpKmAsN45a62Up8jvBwc8QZLi
UpOuVhPRC/cLF7iwwRj9qOfFMXLabVqqEYBhBmTg+9oIBt9yeTGMwq6TVlFgFTpdd3TP2V0mKLhd
AA8HW4kO+CAYhgKffa6AApevwLvTQ13QD8RxThN/VMTOAV89+lJ/10DSV3Yri1Y6Gk/CvVGI9efI
UG7WIXu6XvmiBfx3cRIDC9DjUtrrayVxBsKHQtW1KcPOBMVBTGI7G48P/oWEbSeSQ9oAq0xMt4ua
VlfVIhYjBvXwUWw7wHF84XD+o9a0bUGmANc4lv6UbcUoSY3v1qsMIkCOt+NQnl+x5LBt02FctNFY
e38iRqBOYwOp75UIusP1jjKOgZUEooR+DQHOKdqkIhI/AAq/NBTthO6pAldwIu9MO2JQZGuXcJPW
cqVw69bPVi5gBZ0LcNYNuNkQmwoGfdUgpuVDNe4UxyiNoTdVWuny1j44wWugdsKT2yE4QnkSJipT
GWsGK6l3Dj+UDWDeZr1DDy2w9P6lXc2iRjRltfaeNQfOd48mrT3pEf//LIPSZ4SjFlc/qzLNQYW3
Hi+FCh9Q46b4lpyyLvI+rPc2AYJJVJM+3xCakIu9yd/qy+ekci5n7yyu2hLlZ1v7noj69MdP+lBk
gVg3luEvyplRN8qpANmOiQweuA9JmHOkdYwlrYywtWUJd/sHDjrHC/gE8yq0aFxGRFFhc2VHgI+b
Hso2bb0zqodc5lMbNax9wXKnGNgBCxB8J80gz8UhWpboBCLy9t7fgcdrcho7mjj/cdvI6fMzRH3q
vgG8Wmx1IIY3qEIQLHHrGa5JJWO15tz2Oq2vZYrD+t1qsbPO17fc2O4Z3wczryKi9wn/qg/vGZGg
QCgZVrXb/AV9Abqf6jU5ZkEbHQB7hpPG/6HAqdA5WmhflmD1n+9EHeo/B81hmNLmAg2c2v85nwxo
D2Am1/QqYgz8neZ5sXlrvEnRm4S/DVlnyjFk8m7/OL/Ws5+VG5q+WQG2B/u6LXPmETQZXh8j+HmS
2LYbbJohvNXeq4+93hIHkfIu5Ma4dViSJxHnf24fB/6SZIkvpMUsDTn67G7Mmy094Ftlr8OZS7eo
x0rQN/v7nULch3QbvpdNsY/tDhOClnz9Wcb5mtiNy9z5mY41MHbTuNx7dM17dTgAg/lKEdyD47L8
KHWO0y07eiOJZCCrN/f8OBoyfYl6T3wwTeEdPI52fOX9Bfvr3tHp4tWVs57jXu+Sbjo9haUvU8l3
todFX4ft4Ifcg+WAXUkfkyX1q3My8jqehXjZ0SCic6ShvGjv3ZoR27AF1DIpEDiTplmDlFHPhh9C
UBK2B86MKeSEK97+Y3Dr31YiLK8D3r4TkGHVP7NSdghAycZD92eJVc2JLw4wquL2lerXaIFaSeBW
QceVmRgAkPGZqbBS3Fh8xQ/q6aMG1P8KEcy4pFT8fEr+6Oz7LUuDRzqPVRCa+mqMuNjY9HhXJwlq
w6zs0Ykl5bQoniAFjkwbkFGFP1Wnu4MPJ9C7hRzckake5pduhg1JVLXKrZxIsYnM2FyNKG6ejTcU
MdNqs8PqAnMAoAJ9KOl40IBYko5QB3NmwtrGiRtXqn9n4o3e4LJ2XX1/wku5t9QanmoZxIdShDaM
qTHTcosg33cuxLZTRnnUSKRuftTCdmFPWDIc3rhqcOVFTQKn9NrFEAXCs98cEyKzWIfKswMr3BHb
7GQNZGGtLbnNBDTxBHLRIa8Ir+j8CGZiU1zGwUlGdU3ZsXXYj4lql5goRxWtlLGqWC+q9mQ008FI
Lpd/R0xsehXJseYB1sclmBhwkVlrR+0KhD6znl/5DhmwVmt9aO5jD4y+9Foo4P1+50LfyQyvIxiK
dOXo/gOpVRQLZM3ZgSVmJtwzIeOVhQRizXxIsyL9R+LTwUa8nbGeaCjTiSwos+8IoL0LyHsiHryl
E2krLd2o/4VhuctXfpZUpQh1uxcyJG3TItraqxVW92lRnRO93BiQaoa2UlltCxzS0rVrUAHJQa0h
xIa+GoDg+M9ihP8DBgZA76h70sn2NB4huFsv458nDUbSRZM5/FDlxETcufONBKs/arFYPyeW8U0H
Gwz3Usfa0+1Lm4sQOZWREEJstgR+6SareU3KI/yXcFqVWlmNJweu8DScu1tYpnePmqEpFTcMYC7s
BTm6t+qMfueJIbsDeZB2YpLZdsTeXKJoc1lIiVfXbAuFY38Dwc7k2KdJJejoJG/MdyC+uDQxMGyr
EXTCUYz2tpm0TFcalRqK7KGb4hiBPMEs2Cm2wwCTVl2KHjpv0CN0AbdQOguYo/NNnece3nfSbXBd
XreBKhtIz+7rh0oKQufzuZGWhXU4bBLjJ2HwtzdmJ+L7cFqXcVNp6XlByK65H/1HYOoaKKwDt5sI
P/AlXAeBxnsgK5IxuVG47E6wGRNaAyJhz91MLv742zynriJvnDKoOfscGLujb9+H2tMvmGK25NL+
azzP3i0lE7g3Ew1BfpeqLPmOO0iJWp8G/0fEIER9yRqTaoqDl1xcUcQEYxp2qydWHK684BYGDjaE
t24XMKuejYXmRXypROvJc8+i7kCu2q0oLbMB5fK3KCPNI/DLkbBnzPwze0oKMdDD4AzbM4UYjyBf
6Recm7LCVW9Kg05qPD/72THxlTbD6Uzlo52ZAw1tl6mk0SwHUhsL387uHXfk3o09UKzwlL9zMkd5
TcRn5bM9ZGZ9a1LDcUpgIOzbP/fqTnqqL0l2s6FQdPCDqre5ex81Q5ng8DBIZlg5TTitd2rHZ3Ty
NaVtSb+bGNzPz877JIbnn4RGOA0tQUTUKoQM2kF9VECPXrO9rUjvIHPKD84sAkuX7Tx8qK9z5g4E
StbaFRpGKAF4FW5pYQpwh7ZR9lrWToamFNJJvp2DYAO7pgtpNhSw/p5Fpw3IciyZM5mU4BKnSEus
cOPlJn/stVJpBgE9hPDMV+1/6iHou5GDWnvMP8//4l2nnQKBoQ5C2+9YWOPH7i8r3oAhIFmUXKjL
pzeAVLLD1xuNGzqbCie+2Z35qME+X5CdMD2b2zY9kHrOXKufAycLrg0qcbBrB8PpIGiOr1bMg7SP
R2qg803aqQ86IZuEk5s8yNNCMU7IdCIHL97gA+pIPIJVwmMcD7EuXh1gPb2kmibaqVr2TuBryC5C
uC5kScdG21nooyr1YGtSMyatZP5VMGNTkUUKFjj5h0g2Fj/TpTf0gJt5QgJzU378YBygphf+9yvE
ameySYM4LpojSyBPlq5Bw6EWhvTVBzKSjSkx9+YK9VojOMtbfbtE5YQff0Mgjwo8BzMg3ckAUv21
xGWGA4rxWf2cWvur6sOkXDmXhRmrSPrU01KsvvpR/n+SfdoHl/m6l7RXvZ2DODgKq4vaZdCM+TF1
GaHyuHUjfs/VhcL6V3yNiu31jDqyN811hpGPPFXOmZEko8hfGnsY3cadf4ofWv+amCBIEk8Ypkq/
WCeliC5c6MSaPd/kc8dnYAmg+cCs0vsNj8gurPti9F5WKOwzHe6Agwnb/zT+A4R6PzA23TsAnSdE
RJfcTEdwqYZi0tbI7NUjebQZkM9dPj5A9Wl7TwuLP1wJ6yr/+EyvAdPUeJ6QCiCx9GkUWaaSEh2a
yyb9zeTe45gOKFS6ZIdphhLxW5eatvQAfbaPzT6GwZa7yKe8kSzqEaN8tZuPeOzfLq0hUU/FmyKq
rSZcUM03AG98fWwoTqjvqrCg8h5ls+wKfJAUmoWZMAeL2Vn3inEoL5qNmxQ+U5t5+S/blkrJunoG
KN1kgFpdYgNBg0QgPwPpuRbYcuLuyJ0Rt1iE8Oj9PAUxFS9q/+54YK/fqr9nh58JzAtxpj/JwaE3
VPDoqIc5e46oycTQFKbgDxSiSSfccXea7JKBau3+RElxLLbAJfVHP4qwOky2YAmHXiWTAn1X/Bt8
Gm+yAL6X5Y4ws4ec7iJR/GLDiifiLiXN73wjG6byEtcR8K6RtZO8ezUJ2kD0wgLwx4tHKerZYbgk
Sc2Dx1nVhMjX1B3/5lv0kmfrybBS25Vs0qkHzlD2oB5oO2T1LdvFiiDWxhY4xNLmLFRVc04KhIwP
2NL+zEAff9EoxF97oxtZwi3svpbFe78QwJRjFyVNGFW/gZFksMggpFk1caE72dInAofBUWizd968
JB+g4aGJSPf4eX2aTwXDBZl8zCZDA40WJ2KABU6NHL7BE6i6aSsbmxLYprWYIR3fOf2KOCZ58Q30
DfQpFq5mn1uh2ymEUEAjgBnCNR0HyOYB6Yy1MDS9oFLhcZNyVU+Y7Uam+93H2ujPpU4zhzgD76Dd
GmWONYEX1Xg8hfmxOqD9BWgPxq+T+MerVFRm3TNMmb6GpYSXz4Eez6DQ4b20mnT4qQ/uqr3SzGmR
DQDnFLo6JRXc3H43BvmQnl9mcHFyP14KtItomjVUt3MYvGoUJwQ+lsAKNEH+xP26loy0/aTKFjBy
RMy9/W4ziyvAOegJ7+4SDCk6pwRM3rLCPLdF5oDV6Ut/ZcTNz77TP2vtztA4izKQ07UH0ybwiQjo
SjtWAyrUu455K3ENIXZwc5Y6oWPt67lJJ7c78QCOUSaTxd0iZ6d0Bzz+y2U67KaVeEdxnU/K1jF5
bGPHpUm35T1ce0Pq8DLQN9eR+rIPNT8sjObGpLYKFe0lFwIYrfReajwmNaTGn9384gYhJzCo22f6
tOmh/5LepwnmbhyFiDGP/Egx1dDm5U3NHbWzcffMF38kSeZgFBaqCEJH3SwXheuaQUGyuQ0LS+hA
S6JjLZt0/0qr8r8dG1O7PncnA0Eg87/HjAyhSKimPrnW7kq/L2/QpEuqVxecZOCBvegIstOb3qOE
jbtJIA+4YUG9fqiLYKyfp7/2tiWmB/CnrtdANOfmcvmS2UxP93AuCcIvROaQZ8ha3838Kd/vuh94
rNcC7TSgWGDTZjO6DLwU7VRwAoHMv7n1dVm6KjLPYkUWvlkxxK/poT5Ax6qQUROqlSo8NZerEzOJ
8CDk9W/wotheuoPt7tvuo/dzSl21TN6gwH+uyRQe4IDGEmaCO/XpQXg3DmUQffThqk/3KJyipMVw
5nzFGGcJNJwmS9PqeA7r++gzDmGqiE/uMVQxtdb2YrzfwNLrux1kp+N1i+esrXh6MTb/AdMBaPcH
NuRN1kq0FeHPRctwSS/NGJ3SUBMGi/uQsutylfPRhauR4zo9vRC6zH0ibh49kbg55pB7Py7RZNy+
b/OsM61FqJ7lmiAyKgiJsDzi3DTCca+chWZw/Yh45vBuae0QYyis73vPIyLrCDzjh6zB3+rxq5cx
uXIvxm8zETC6N9tfRp1jxxMChc3A1d7iDJpLP7h20OxUhLdcA2c9E7V+JK7YkJtD14qpfGvv+AQr
b7upnLn8w9draxVIO6MLJLwY7D4/TNXEVlTok9Sqi6AkxsIoSBZPxOE96z1o+21sQdC1DCMnfT4e
mUQ7klCvqtvfhFDUW3bZaFtzHaODR2qq5pQrERrVtWccuWAcrWsTvLx1mFDR6UaSjUvO3MI2SCA6
OxGhx+jPAF/uSBBjqXkGFpbvhRdfIxuvTv6CcVuEryGaGpleMGYoBCJrAfkh6O8q5emlIqX93klE
TzLh1lIyIUw02bRpIKaPnNJVC8Wd4xjDOg1h7FBTqcmNlIT5rUgPoxp/9goGQLRBK6lWVyqKwhWz
kZFs7FlQvDryhuTg+Z9fzGQidt8DH0bwZyCE6PMTgKQBgdbZ3GB9FB0567scLqUGw7NLbpGHKHj/
cNec+x7bhSJm2nc5RKXlzQ2SgefTnpy5+O93iu90lCOZRPL5nnms/5UCKGCpFiXDo5KAn7qe5J/U
zYwtQ1wC33unLgqqp/A6M7WJdOj+Cx8dkmITgsBeEcWDmyyfTmX7KKwCIISYHsvIQGjZtAKwqw31
5hZuSxeVCqx797xouN7wAu32R6SHuxLHeuFQUnedo0A5BccooXicT8bbXApr9eUU7ydsRRT8CCQ5
uIsMe1sDVCm3/NAGxSbHprpu8kNJhfwNwsVf0N1koFtQ8AGtWK3Uuv+955/cl39FXkDThttFdWdV
xZytChagCEixyz6HnXbai/kwsl5Z5TYl1tAEnXbnNPgMBX787Iorbi4qaCQwYhKJwmBMweP/LFY4
xZb/TWAZLWVigz7NDyGx9UmaQiPqep9Qx/DEF1B/zgaDL1x65LerGPRjw6+AfMZ3tilw1Em4mzlY
QbSSFZ8uFOI4JUwcx+//cfpI4wR75t2W+i8ha/D3gdlF8s1y9aScFLm7HUj15J2YZzQuZ6gvTGuT
ZWebOO37o2dt+8nFynnypKK0sfBgeutUC1lIwn9d9F+z7hPc+EIlouiJjF69oAamcH9by4O0N6DS
fGAGZ+viUbprJNaQYEw6wdq1OEUbR9w7+f5S7jQXHH6w6bjn41bCY5mQpY1D5wQUyJ12xCkNYT7A
1DS3tZTuJMozAS46rdKe0vdNPQyl7n1hLsC9LKLUzkyc24N7IeIBaEDhqYsAbjU5jwpRQLriZoGa
xj3Wxc5QVLuv3aOB1JjzVY8lUnhuYiSJsFJkCLBdD//x6kaQ02VLHPCX/vx/U+rE3DTBiflf7ajV
FCaBbzvvTz7PWLGRlPc+nd2bAVZN0MYOLNOdSLMILDE/Ax6QrKZ6AO468w4+/6nDbFhgvc1cxSdg
l5GYOdDEZOyY6Xy4ZTZ2vjKDEYhLQ7FgFCSggxY2d83Jz2/0Qd5DDH+d/3nh8noP8o81nIpC6OPo
Kj2kxOQpa6sivsgZh1McyMj8pbJHM9tcv5VBhjTFDaktxUlBeQxPaPlxEZKUUvfsZ6X4a8fnOvJE
1SiaLHhZb7ZbElcNiT0+onsa6uMXBEZFuKlyO2RA7oJMV14WafV/W7HRk4VioLA0IZXQ96B/wRXS
cOQ349K1+MLr4q29V1JOUUsrF7I9M+Rkb68LyJGxlgGDqHl3BrV5VlAnPL1gZRcOh7J/XPHYY0Pb
DGF7VLq3ubOgE0iUb8ra+wMYQ0yez6iWxDdKdV0rp7Ahzr71k96h911ymErXDqpp9O3F2RDwY8LY
D6i+KGKlDrqKvwtFTcOuGM6z0SNjXmfNTTO96WbftTp2//wG2/g2W2JgoLF12K+fjRdsPPnENZiT
/z2eetOeilogAEE4rJzC+ofC3VwfeXWSF+GQxozMozRuuqZTJDV/5FW0CJwKO/Ug2RUhvF+uNAJT
zP8emYChiYs/wt5PqVGggwTpNqv48KvFyuwABp71eOyMdp7QuZqp/amdRpJqmE5QxwDZBU+ZwTGk
xLwL8UZC7H5V280nKfmnFWp54d+F5la8o/CACy7WTZkLpWrLLV5e4DlQpajteOuK4kM5rm6V3YDF
leDLTsE+nbbIlmtBpDP7ybP+L1e0YdbmJIGeAX7qm0QsHqUX55Pc/86KsJB8HW37GuRwqQgy/4Yy
c2cDjkjIW1qz8jhkh4H2Ek+t0I9WaX3BXgG6ULsB7uVbYTOC50bE7j0BB2pXcNPxxWkMMbn2waHR
WJ6mxfTZEPyjv6J0L499EFgYavEbH/4g8VVcUj1hldOGlHtDLHzhYtpDSUqoMus96IvJVN0d2jMF
T00t3TL3XwZzVg1eKINpcSMAtYKy0o351v08cgfRNFMZGXnuyuVfifsxDS4VcN6gX3Vdl2Oi3lVX
Cfvfv+W2QJkg0t0QkrjwXUG7hEv9HAXL/KMRTxWntgQyrl2uQ4AHInqxeI1duBWlAx9qZSyHGdX1
gjOx43HjLRWBVr1dTiTwZEeQ6PEJFp4Wk3jTdEgoenUstAHoXZnogg9Zak68FpQWPky6WWoryv8p
hAA+sWAal9dXbVmusX6NvsGx9sBmhUKU0wSiXjAPkHtABmx7zIT8+V9DZmULlgixgsk+L89DGlkd
Oh7885m0hwlC8mgfi6xbasbSgDv1DvcUNPi9SkO4h1+LdMVBRPNFE4+jdDVTDcdA/HD/neN2Bxs1
g1V14D29snl1UzibvkZcYEHHOWToQ8kOjeTWR6+VYcY2ldbCxPh3M1vDAAcdEmk+lq6sD1vWB2g6
flvecwNRL+K1Mb72MqSlb/SnlzWLIVCqaOjutJAtgb5p3eor3FIw2WVm/YcqJoROTDgLfgXdhuf3
R0k5NEFSvjQ0efVsBdQksLccOI6aOa31le20NNlap8uZAkFeUFaUgw4FC0oyfn+pR6XrbVkbScGc
7b+VOzjfNXWhH3Ao9Q1DUz/PgPtdtzd69g4U9P5Im4qlNlOKENpA9drIyBmsYruo7i8whslST5ux
cd9oh4KH3dVI0wKX+Vev3i/90ZIazSRwjnMBVsrWRAUiUeNlcvhWk4Uqq7onUqV5mqsrttrq/Mst
gMDgpw0FiEV/EFXFYjGoxu92lh08Fiprh+87fyKq07EhjsTVbarKGE1ytb1XnrJ49lOnfqkhES8Y
/OJi19J0+Eeso7Bx23K6iHYb08ATc/dy/1lJsL0imgyc5FLEkYnS88uddthxh67g/q3nOz88WSz7
53ubYC0hnXMaovCqS9M0aMHoMJgVmWzXNGza9SQjhVfsKNxJ71xyVTWvgtmEdv3WHJxlfqNaG3IM
wby6qtRVR2F9s83EZDFGgf1zw3DOOvoq94Wyu1kd4UraE0wDDlej6ROCpMInL77EJbH35q1HxJRB
v0T9s4W4ruYC/ayy41huhVnKZ8H2ecOKKLyYQbXTmu7BDD+dSP/uqUBIY2hxqMTC2REWLqAZtTty
2XDJggvn9xjC2qcTaGGoZFQnEgDcVhc4MCTgKsSbanjCm5DHcrPG5EsFWMCTBZwcdBTU9oFw9fOf
2EFMqwnSlnHiR5uTFpQdNtpQDFrFhsWpPl8nZaIFf/FO//EJYU9cA02uL/jX9wrrLLd5dSzRggT1
EAWAabDTMH08hf5qLakGhrwfJxNh/somb6/BsGRnJunSLdRCeK5wYbk+i/4rYFFbyRj3vVZnHrgj
+ykkQUZlNxO9RLX4Z7BO0dJA4eJXuIu0k5h+UpyMpWm7ZrADwXbXwk32qf+1sKXpzTUNH8WoR6I0
rODg+vTil+2aKfKB1NhTkXbBl6qedQ33CujwSPqI1ji2nPlL7QsyDmr60afak4UfvAiVXlEFhByr
ZZOiTrlzovM/wb+G86mX2YEpwB4e5Ip1lHlLnDN6Gj3N2hwW3qewO7pQHv1sX4NX3f2bmX2qffv2
oYn2TQ8n29FjBRfwrEIY80L+uA2YRiMMWEE3dyCc/t/nhN5DCcZzCaJU5sO3yd4kjjGELwUvA7lh
3DDZ4oCd6Qy/ZIn7yHx83K9UAPKvt18jXv4avTt9FSCSQ/PMF1Rb/NwX40dPkSDUCN+VWVSksMDp
s6ZDJOANqmkWlFUclaL5JrUtUfjL5pRsBAwXqsnVZSX+RDrGWN/dUpYBhZmK8YnuZHRl4xmlOLXw
nNCL1CqOgIBA4kF57P12gY8U8zkdEJsm+JWPI1dn17xvBIccQjvgAanmFUII1SW2pkREE3gzG6s5
3yPhzR/CIrR1sDDv4SNBgoyg39Z3SpxmQKgT3n58zG6rpoxr6O0mThSsyPpyUw9AsKdf1FTi9ucQ
6oLLay3rSH5zN+m5wXE+y2anUCoy/WB3ueVb60XGjsgqFbvfp67F3c852yAeWS/0a7sxLxD4b1oT
SeGb3XFzNdmDFpi8kGu9tDzwGUrtBnBlCFXgKpD6qJ5N0h5Nzcu4TI9FanO10oPHD9XfIJ5EDhB3
6Z+i7fy2xR125JAHjpA476wsx54YuNabC/3A4RlKoH1CuDUPI4MNXhYZoNQ7CDXKe4g8XoqL4Xdh
88tt/C1kEpff5DeGJ4Aa2IO1EaDFVeKpN7fbIihptba0fR9QyJ4vHQKecFCpoeFXxA/E8zKW8fj6
vW6bV2OJQAoIcvcLqT67amddXT7dNgDKRNFOYht1MFOopZfScRE7mpvXg69UGIworvq0U4Ofq49k
CF5oChq51Tjhi9UjGPl8Brl3T4GGgevMIsGgBFB9JANpWVjVi4kQHw/GYeBqIFljZohTXva0FMzH
TnQNOV8dVIwdbCW+Hnf/3nJLUQE6U5t6etpmBf2QNH3Y2iIIR2Vcnpb9Sxp62N5p1TDgLcYztKaM
NQIWiLZyEXuC4Z+2fcRi9FeWbeM6d2nOKKQTOTZytW0qTCHReRjlgmQSkEragVSRqD09bvcBNmax
MrCvlamA8/N8E45NDTKfbUsMwO8eYHKqfqObZopU73whGDEXca8PlJgSpf0wyccQKVSP5tWRljoZ
OYhnVz7UQn6Y7gDrRD/GmGLqAiRePhJS2FWT/M63SIUfz4PJZQsXM1+7XLq7RmzYcuoziOoqv6Ix
sFvkJi8L2CDDdrcPKEvp/Zr3H2bAX19W4YwiAgegFhCjQ57qEwc7n/IYvrofQLQGz4ewsg/F4Js0
s6od9+S/TumqtggcgBpJgoZNPSuSfVpwqjWJNMDzfGdp8m9gIPDhFk7eS97gB5lYEvrTCxvrnr4+
MQ2xM6ENsHUuIgluo8PQiiAOFe9bCQ2kCX4WXMpKc1CZs6s3YuY931EFrJABNDcrSH5JvTd1RSpv
CWRNKIhvCziywUTs9HH8tH0cpv5MEwJiKEb0TAsF85QBK3flHXGwbhS3wm+wKi7pvbXBdQnq+n4x
LsDacMkNaRY2OQKQa+u3t051k7V9pC+5hDDwxHFEkNriRq6KOl8IdASoOexvwARiJd1cYCBQq7pj
fRbabqnq0Wi3KgCCjfrt2BuqySdjiHq2YckgYseCajltySyjvETdsmNFKfZTM0ylsT7/qVa6rD//
IesgUjroI8NlyBZ1OiPqjFvOpxK2Ep/6fmpNOuI21p/a5TI1Cgidb8ohmh7pWDk8ZKdjePIGSQXg
y0KWGIrF3G1eYTzzk9fIx6aqkSp0DcIx1qcPVcZ9hdP09489+05KgPUtu5dx3RHMCPWW/DxWHHrH
N+5LZ/KEKsmGMxK3nb+osW7BzVkmCdKyIA6gEWkYsJZCx8RqNXOLLAl/8WMAKfk66rVRwaIUcewY
h7+7aUWjE5bnAB4tctbPLDXRmivJ+AAvYU5mAlLr2nmZ2sPH1MILMIatA5STJxF8x7KVecYPL3LM
66lMrosx/8D15ei0VyqKRbFzwe1V6XlS1W9AIFCrrVVXwhxkrvjDVmhL22i7p7pEs4fNPzqbbuXo
C6ntGC83Ut81qPPkGE5jsnBhsqawLUY+Jqs8EtCQcQoTNlifJ6mIIeDlaawxU3By0mnq4DxtC4dj
WNrtf4zCwDklsW9AA+fYrah8LM5qD3+vqav8pTR/aIXG2n7OdnZbHgf01D8TFMR55V1SYVcS4gKz
RBo6MF0iS3sXPKGOgHukP04T1LsftBbVBUdZ0a0XbMdGGlEzMF2qvgGylDYhd8ICyfMXJAsRi5HK
6movY5oFE86Yp1duZmKIrCwnYHki7hxonc/AJBhKp+6ViMr5bsxzcQnx8MRR2GEroQzqHA1mHYhH
v5vzgMu6NOSlx/dU8lAkdSF6KDyOz4q31ezfJ9h+01qQIUPuYF82+oPTCgVp51bNSPOJFGsVdi0M
S5DRVG8MjFUYRgm0nkO0McfRxe166VWJLJN2V5DV4aDeBBdXtDqFL4J/6ZpfrSyIVQc1nTFpKtdj
UcKXkj3x67INoARbChC8YOA3vybZDQwM40IaM2cZWaWJOW51lt/CASzbq5H0T90W5NLFSzHFMe9l
5ZyqAhOMP+xKaYOr8tK4AHfX+YuSfvYV+rnJB1Tj/VkTLgruFLjWMZNQAAwAxseiqrz5pYUusU+e
uoRHsVxLq8vdZ8qNhBagEUCJx38Mqu6XGI7NNVTwp8R3GWXrAlc6gvHO2WVvWGhfYaK4GWzy5rxr
1cjC+WB5kZQbdKXPO393wifvAg0fDGRTpySuy0ti/cSrXOJ5A/1fizncGJEI085m7i1pJ1qa6gSd
HSBCeC8+Lc7PDJ61gVNlD2YdkTPNNBfkQ8qiAi1nEys1CyOSZhZHVeIXYRzo51ksZAK9qD0dfxYI
hX3u1AyeyljY6XrAqrEyUlON+wkgUCFYRJ8WBmWIiwhEuIhGj1qjDBfz2hUprFdnOUqzIAQoeTBq
qQ8PFgT9fKk3964RUyFo4eluAJ+ATstC9/muaixTQ01K9mhHf5C+yLxeOCZ3dXQaZjHEhb5zilLm
WIKKkFjc0UmXobW3/Fob7g1N9T+q6CF2LeqQEfFDRL9iHpB5xZWQA+n8w9lTJgeYyZH4BUKvlENt
yxspp5wF6i19pFzMQr7NQ6jQY5uqir3JkpXNKgE/W7f1C/BVsk5MWiSwrTtXWDk/vNg/55ghIWzO
4IDgzKfm9OsT5ASOO/jWqx/z8W7eJ2wPSsBqNZCZ2vwDGsozjZkYFIbzHbH8MLTjmKLDgu2/K/fA
3eQf627mP6AInQiFfnYXCvd3LqUA51+iC8+NqfwMTaVD07a0NRgJyj8NytswcRMNTiYR7rAI9FJL
cmpINGtEpw4LelsVqWaUs8q9P0kZ7KWavAgEj/R4jwISNRs8pfg/Zke66esLCZDTzIeSsIbsJ+P8
GD796A9PO4Em9JGzLQXoCFJFbE+XIja4r4z5R1qoHwhWFIghMmkmdsZpuwX52cSYjAgKime1kKnr
Mv/0q0fhDZ6JtpXXOgp64JSNUHh9ajao2kjbjsAtT+KXUrHV4OCoT7CMaU4xbT8Um56MUJ2YernS
GchZyRdqK31k9knZmpSLSGMWl0FQXmMWLEFznCNdquItJ+h02rTlIQpjmR6IC2ih552BkSfaaWth
qUUPTc3iZI2QlW0aPrWVTxlKtfesCdnD5m+2pmMCTPvGQ+6I6hwDa+TpORC8urNoCLjTAWOcqL/0
PNP0JoqQbEqFZFBD3gScH0YpeFeXOu2fqt1j0/Dv3+Obe+iq5vw+awrXeHo55tnSYVJ6RqzS7JDo
OH059OmGV3mNOkcbAT0yn+yYTsGXlf37n2KmDUi9hpWstYiMe/HPQ6wU9zgx7xdfdl/pda6cJW5C
al6na2sOkN2oZILg1qwpzExzXJsljPPgZ22+c/4HCWW63zZA9P3lSsTcK6znHoCyzWm3Yt7jEGQt
SG9i0G9dZWRi88l78BoNqliaTb6JbeBAjqssQDOaZx5dN2GtVlUrLJusI4HqoVoNHVu1eeNt5Byh
GubwrvoLLtSX9qc5t7cLKItXZBrZ4RgSEny83Xcwv6K93lODUDAxUb7Q19I/cm96DiPvswPUsGBQ
n5wHBiwc49F8wbU41LsyP3ZZy+n02Hx/67MaMFp3J+5wmRBmF7n6+aRJiElPad3v0zDNVChx2WSt
c3EHpuvr0SXd5jTZIJXiqopOX2JKym8dQe2gAzCu8ftA3WH7vphaDCg5a23OgRx91jgrj0Fw5CIA
AzSem2ehPTRHrOXLNNumsRfIg4tmEYKB3cK7z7zIK/qjKpBFM+tKtTWjoyfeu40pc7jm1Hd/d6Ar
esWkysgdkcCoYecr2vxrx+in6fysPjQn3jFNje1iQb3j6T0YZEbu7XwYlCwCa+yala6irgiO5Wnf
gNyIb2oYlaX3xg2BqsgIciNvyh0+tw7fINxkcF1pvQjLEefKMT/IwpTOQcqU3OyQo7fW7VdP/PQP
1zyIcmiUhaJsUBaVvjaui2/5sTwnytOzbE3GWMUgryLvndGqrCJg7VmnmTzKRu8S2TpWVPPJYXPg
rMjjnAekQJqGs11vilngoCxeIaTI3/4O+a7ETGmEvyhxJuL0b4Qf6+7vpJEJRswlOIDYGH8/iwC8
cBCvy3vQZRABpKOxPqxuLJSzMITxwx3aWrSi8KCEQEGCYB2fx1XFXcij3PGYTe63pHFcuQblqnOI
15OrrKRclSRS1f+ylEiGTh9HWxAfXOy5RBtEvGEqZh4sE0pZwZ5tmr/r6YeJUtvVe1qM9TQV8w0i
rHXYhDu8EUeWlcG3vFPujr2Pl5IyB+gcfVd78pRZMAc61LzNanDhlJfj+O/Ab8a3NL1EMf7oP91T
IPDY5c4Eh76K2orNqYOG92mKHwK9wwIwoZxykBsv5VHMswXDAQumIJ1pmzKNwMaf0IZYNqKU8QXQ
HjnQDTvP/56ej9claAci5ZjkRY2f/3iB+k5WUHPb/cEmjxVELfk0Rxempq2HZh1/ut+afQTMfxT3
ZHfo/6oJ1CNIV6Rs7MSWgLI3imBWEw3LPhOhxUck2DxXrIiRJqfYVSD66bQ6rUyf09c7xBFWubns
8RVvIKjHWJxZRhy8KCjlHX+YgnlIiuzntvphlfVXP2HToyIIqiqqqaEY1A5xV7GzuOmbTYhxoHkB
x49piqY9dSbWC2KfeYzs9DxfV9U/0M2cDVxpPzSvcIgCeHavbT5swku2/I2PWR04PqZt1MW1alNG
VdybtVNh6G5a3ITivWDG/lzmXHWgKLlAJrBkJ+rUXJKLHp/8K+rVm1yXC/yTH0A+dQP2OoEWAoJ7
OnZyPFsLcVGIvMfGcSYBN3vRNd6Y05H4Y4bh6Y1McLjWkv2AzCudLjOgRzefW1Oe7TcesbcGIrXf
hvHkeiLj6j4Z2+qkhUrYo+RNAOxR5SDTqqpTPvIc9makpwnIjg+jBDUYxKTxBGoD1jlJtO4vhenT
K4frlSc3i8G3pWFMdDjfv1g4BtexpCkP0Jze9k6c1Jk/vgXXxEn3j8RtxDW8wRg8NuwB1RACE0az
GAfYbRmDZgsqQAhUCIPJNU+yG0xPyzW8fxn1CS53Dk+UvfW21bYMlstg1WkMTa/uucDfjD0xv4Cf
FxhDXvncgoHYga/i9pSjesvU6yIFXACDijApOejfEezcL2lk5kFA529s4jPk4eqR36QVLVwYOLLE
pLJUpYzmTHvaDaEVw/PeuLhN2yPU3RK5Ek20d9thPzIRHzKKXGGzPlZg/EG+sH93wk7jvbc7mtr4
x55b3wdBslFMFirX0DFd3wbolwpp+2Yx6XekvbAy7LDF58VEVkdW+LICKOpayFyoAv/aBZ2mfnGR
GgPVYWW3YaTEdioO8kRKq/Rg0qTkf9uAn5zxx32S/pcoMDsBFZpAX6tLtNH0cGeTn/jqfZj4BEvV
5S60Mt4XN2gQQXZq6nBuG5a27L4TcJ+l7BxH9fUGeXHcQH3rhoIXMGSFS600iL9lNGEzRaVYTq/t
myGXH9pUdx1/nGh10I1o7aUX9e/Ypl+df6YM8qXa7QM8QtomMwbpLhXJ1fHpwlq1QmeoaXNDFDVO
esc9fJuJZ84UwcvcNrGydzU2trK6Wtwgj0OJZ64x4Xh04AcAscVZRom7Bg39DWzxpunwcR7BMEsg
jlR5cJpiomyP12RA6t/C2GkhpiMSeOIPK3367LMEOBt9mCCvfwsFIJwqmDOafD/glgT8aknFCYF5
Vb9tVI+jHDCtKWVzhOtcAgtRXKJm7Wc7TdfKuzBB9R0tpjND/jhdeZi+kc8ddpctJOBrmbUw48vl
3l9fHZxXNtKXtHUAupGO7rCgD4cfIVaL+0CeYM1Q5CIaip+YeukMLegz56K7KQT6buGlDtsdVfte
ryaVaw7tvFdlsIF1CX6VQK9mPberxtRudFov9JFQqk77ufhkfpDaXNYqoGoKmRkP9kXOHSPK0ZAc
GOnhWc5ErLmeNGWldSCMgj+7L2SZcBLr+hc3mruEljDbmMNA4zz0FRMH+PHr3+1/lJTi0qaMaaZf
woNfP5/JkMbqOnUz3KEXCZPboeYTGoUL16Gcm+xxBPWFdWh5R6Iih24kx9JAn+u3j4v9abvb8Z7Y
IXueF3kSOOPqCzCloUv2FHc2BdkJcRQezpB76klA2LLsPBLOhkywAdbhlvKPgITDALxKy9NUuuqy
NNrV1Qa6dxwjFpoy8rJKRSokFIh8BRqBSu+0OlWHgcSNyJfaZnWvw7XAat4ZwFhTnFyp4lrpE1ST
EWFZ/89KRxSNr6eopl5VjNhcSeRihnz7/LCSfKktzWcSwVD62UMPbewxSFV/SXFFd0x7WFjkY4ZU
YFIOMmQpBf+ozAi/UfkmK1NE/xHX90S6G5eMYsa8IMUIrze1H+J5lR4LoCP4Dvb6bzA5dT+KXrG+
hFDZJiK8c+o8aDRozJndWN7riWLLGFiBy8WNeFiC8b1EbiTJsz+1/Fdg6EnD7yX+nk2gixUtAUlF
Pp1EGWSX/bdrQwS8+UO0jteCLuVUWrlk4e9xZqkDlIbAB+hM5m8h2M3HTZbHjR2WvQQsM9m6pJTc
thbwQBR+0QrSynrSciwTXPM/Xv0aAfiKb+DA6/azt3ZVn8ikHDHhiQPAAoV0nowvqrYY7vgbPkhG
GOuZ5gtUy9oQRX+VBlENFU7RKu1EuHC3o8QaeIz1CdscsZU5vo8nOU5zphSz4KVs5poS9aCQwM/3
V0pyV+BaJayRJgEUDZ9Ad1f0Hlqmu+mwUqBNxBHYcn2bMzFYqxYxnBYKLwoP6lfbqTp1HvwQVUIV
rocIL12zm6rRaTPfCFX79kUH+AtqIZ53BRDLPMkGCyVkh679H7s/oFyf7EawOrAUNI7NOESRTm5v
2eDIvwCOvFHCU7/1IFLjoInpdyNsusE+c7W7zDDzDkfnnQ+7s+o557jaF6WA4nBzetFGjJ6ZOLIw
dCiVdTA6ZJNejLwn9ojsEJg+arP64tLy69XBaylnoIIpcwyb1LUQyvliQjMPI+OEN51CynjLOTPI
ZNW2I/GeMa61TJ/NBFGc89RXeB4iztdtYzHZL6KFsqPlsZtVKoRR+dRWM5bo/5oQeP8VEaiRZDmR
7ROY5PkvJYNok5rxmuY/JLkYp7gAGE5ewVLbCTWVfDG3+jcURtur2wh3gfXTOH5juq7VGjipQymC
g5cnl3/BRrBNNIy/rOTmQGLM8QLCSo7OR2Eun94qZbeSl571703ElEI3emP1JpTA1fGgxsVLimGx
b9Pf1zk5tFChWnYiBf8kAkES2X8MJ5NrZdsIOyIc9RJfu5s4m7bD65TXGnIV43HdsDTtg/FWTzH4
rHp8PJoxR3LRng5mrZDZF3e77ULAfDSe9JFYcIPhDE96tfOuJbhpKhVPX3gl+CwS0dyhHf7dZgDS
heK9tbjnyHX3urakBgPbOO0lSBQvk69Ca4XhZf+fcpdibnSR5NeZtvLyMEtd+tyXOFuQjqwcfWpC
nLjV9TAUxHorFkbKkkWnGkg6WkiY7EWdGi8uCVutZKvwXxTtEnqoQUFciusTue2Z1ksYmjpiW7lQ
RqPLEe34oDPfITOhYMDi1cT1jGdvICMtWQuFWyXs15Mkedhlaoglt5aDpCyZfgg2gTsVvSC2DP5J
d2/PqIgUToiwmsuykATRsNLuMG4eSkyibVcDVQ/9LPotaLut6iRBgQNSwgvlVr9F3Vdxr/DFR07r
OjNVuGoVuDZvW2GbtTz4+sxuNNEnWALs9SU8IHHf6uI6Uy+E9p2nVGytONI24N4lLOr33HpjfKj6
wV7LBf79uL8FaIlm+8cX9IxM11fOnKqhnHdtLcRjRKN01pWTmEj4x09LCXyLsMC8p1pnUODOFjIn
3elERjyUzr8gBXnB7kDktHYQMr0FzPlCfMbrw/aace9p/eEorju3jqdqNikgCFKeODk3UGbg3lHT
HwiHqQBIn5zN6JDoPp9Q0NVm10QSl/I6c5Yj1PI2YecnfF5aPjNxBZfvdAaTdlBu3v0B+FKAEdnI
ubfBWOnCcLXEVG43ewfUFPvzDtFpvAKn1KaN5ZOBUCfy5KXvaRZt3Jh4kTYDLi6zt9GsrMqg8VSs
kazSXuxU0lTP2LrzsBq/BbiNW3nIqNhqZUDaxczMTw9vdSHWeXYcBRXeoHZugtqt442C6XVEaMC7
2oTVF3imB98BcuKm1gPnLpxd6Tep5dXpAnbgjwMZETHIruvRAoECNvCGwOkylP8ehYbLWY95PqYm
KICqFmxM1Baad0rDcOIlWT7+oWFcosF29P1Gxsugw/RBqj1NVjkgbmMIH6dwOefr8LPbv4wEPMl1
pTlo0gRMUXsECM2NYCeg4FEmpCsUyDxDDOd80nuMhfJSiG9zOW/yG+QtiTUS8FUUEFFPYYbxJ9GR
7kJ/Y+CVifmg7ma9Cjrv8EXJBLMNZ11KFJrVuJQXQGAbQmRlw3EoPQc8wYPnJmjgo3HxQn9yFTDr
oiLlXs1nG9p6v3NVkD6WxzRooLgTKOsqykmWtM0pvhpfV2AcsaikeC8a0sNsiWjDciaBoFG7wmKA
dtOwPYsoLTItgb69+KWKgDgQmHgowLN5/BLaixCTIu1bxPpMQOjZvd+0rPmuivOHyx39EBFhcrIY
vJibDCCo+5vPnulaf2BTHOeiL2rytsVNHtaWWx7P9x9RPWfP+87Du2xjTsJrXxc+uamqyQARei06
j5XT+3KTJO/NN0C7abBOXzns6hucSGVXLtgcYWYIVvHO8Z2vE0rH+dMB0KzGSEtI0q7zaAc5QhGg
qjMkKxLp9/LDK9gCDoGUOtZl0DyZaoOBTB6ZMuAd+GYUa+VCl3F7aXEKyBHYJHoSigMBTTV9qIPG
ERPgutR7Id/ZWgGKUnJjbtxdFZYOLtW8DqGNI5XdMYSDq0JM8KdlJOnW/BSFbjXRXHNggvHheBiQ
80co32DlMrcipRy/RrZFfH7T/h1RfRBH6DVRvbGyMsN63D5cfOe6uRm9NFEeZwlraq+SeW1Xt9IT
oRCQRiTilS+ZQYkd2XSGn/mneuaEBBpJdYJRPzVyKLbJ5khJycqcX7jyypHfFP3EnOGw2eh0FMvg
bMsR6HUjLlxknc0QbA1FXs6riY7E35PDnb4XSs2l/Dzcgm8bgM4Jt+5rwb4H+ib0rb5d51yBphoK
WmAuvCkyMo0VqoQW5LhI7pt8g6mFWtq/MeIe7WARXKfzqbfnomxmjakTsswg+xaMKLUd62sjDHrC
OKYalTNdIUTWJfMuc7JqRI5UG6ejs8JbaA4GWj/y5z7H+vZxS28UCr66ysSbCxwpxdtDx5Wl5IX8
vpUEtCkYP2X8JED/lbdF1JksjkgTEyHvPzBOBUxgUMcJm/ycSfh/fpYUU/T4Gf8z84XN/HYOoB5X
j98rsk3vdRO8L84pqO+TraAVDSd+gJziLU9ndBwhaJuh+Y3x9Q+2/mCbHSuZOk06qeFf3oaw0Yz2
SCQS3OfDzX1O2cYtHp4NcJvP1EqP1jpFlCAk4aoWscKHp245BbiNiBRvvBIPmkdKVl5m2lmh1Lif
GGDrUa0ois/n7KlY5QQvlE29bnSJugE7mPPtpQSSGI4a2NKxYrPKEdkwAb7sblmq6DgbCIpia+m/
ueGx3h+6BBnwZM35gCvrqkj6MjvCmcbRNsvXoBQvsDeI5QBmACM01jPyZdboSs63lR0yApqdH2It
XNiKtev14CGxMVswepas9oGzXOL6ihp5skeriEjg1YMA02oIV4klh+6B9tD6aQzqXEwL3u+ZvFiX
nN9EslWwdjLJZLp3S006PXQr67C8RlXj5AOr1rRJQy4UbvGZ3GWi9t2EE8tKQsPqhXoqdMGi9ElU
dvoc1nIyK/F94LhHNqSZ/+752QZxwydFWFCmfF7TT7ELZVf8TWpEbK5Nci5VthMmqDwXneo0kl2E
v3BYlKb4CBpB9JeJvXou4nMgjMeH92tMaxsUAUXcPDTLU7RYzDQLkfcVmwTilXebgl2rE0ntRNfA
4dPH4DQEZH07r4xGTE9hmPPP2osXktUFnhrUxveH7JYdXrmGWw0wGkni7Jv80PmORSW09L9tiHUQ
ypjD/gwS3mTd5cgl8bstWf5MXR/RDqc2N0wjx5ajGJaPUUjLNySly/78oL5RQlEBe0DiYYwmZIJV
xSTlM3XGcmI2fvWV8Epti08F3fQo0sjYvrWl25pl3Wy8aCIZzlZ7YNmy1XN9UKZJPvCn5VIgSmza
6Qh7+DU1LvMhDjTSqH/FE+Lu1NHgvld3jcDJqMloaZEph/sfLq8bPPiLjivWGkvLZFwYKgCsjWTH
PTPXCqLOp4eqohMd4W2JyV2But8NfLeH17iHQfYw4Ox0FEdHgE/XO8L9/ht/EbnGfRw0RLOgGrua
/It5/zFc3+Fe5kYpDDkUILXBV+qwF4tMzG6FKntyOM5E52uLdmrTKWtnKTbAvySIO5aUVwoxazHx
Fv6cW4ckVR0HCLHSVchoFQO4o1gEqm9eOrlK9xVuYobsFQgVKwC1soGxSdCwv352aiUWdgvBppfD
tfiwPHlKKdM//v167f5XPsarvbsQ1VgdUaNXi8Ozhtowoa5nnqKn4DdRkzLqrvEqZiTEBzHYYfka
JWsYmiMZ/J4iV8yonfpvfncrpHKtYw9vOn2L4KTrNUhvZAOURNBNVkJLCmyAZsQPkWCeOzDQMWd8
Ak3uElLHbeqhvvAXaKIr6OqZHT/sFGQ3KXMTYioenq7/Tv1f7rmc8wlQKCzwp9uwSONyPClwBvj9
ObKxA/gSnX0tZSqMkyuogtT8sZzHlWX6HXgbKQC9NGum/VErjrw6GZ/XrsxM5UT+RXWc96DkpPsv
2LmSblLQX5MEn2L52jDvePG8EYdwYX/cxduhjwOsPcqV8zgcm73ehl2Z+qeIl7PtXpkBuhYmvKjy
d0l9Sr1X5e3NF1r7lEwr+ErzB1gnrmm4WqkqyjsmjV9+gAaYsMCnYUH2tuXC7jPWIcdXzxRgyT0p
DO/51FDQnGBe+kx556LWvp6tMHuyxgDQqCJQ3HjqyCaZMz2oERrG2I88yUh03kEFYl58Pr1epbNH
6oAKfoMvzErl0FOSWL1QV6FJBJ3D1/W9jLksCAM10+YNAoHskeacgqPfSiwFdXolGHWrBRB0FH8m
wWj4TBIaLDgT8WtkuJDNFRHOl3h0FVN+RnibqhgH7ZL0frw9C3IRHCNe2mR5ldW2+Z7j5QEgYxDr
p8SsGdZPZFDMhytk/I8oQLLDQD5waS2+FmucK2ZVK1GBcOpbj/mmSfuvIOm804WF/5dm98cHnNTK
psXsobGDvlbgEC+UHuOjP7rN67IybAmttzptHvyuKsxMAXSHL6/ghrNQX4UmEPw7zTjco1eYmBTR
SWUGiz8+3YAgoVFYXLDqXA85xg3KuRLkIyre3PdKd6uhmUf+7gp6trEcTRF7AO6djw/CJsJcUi80
WuVbkiaKWnexWBpzmkC0fmg4bqWBTOGAEdl09w23Tj/bQiktFinjxvqtHlTjMtx7SK1+zcffyP4A
qvKsIFJkgGploQeZiw3AjDfnOWL6+aNo68Nmnkr8XtvJKfdm/Yd+hYjVfkPQPsLpGeWNRHmylFC6
S/Axk0c7U6Gp0ZCIppPocVn/oN/PV0/I8iM+wTVp68XtIikVJJ6vx2cWVQk848o/KOf4prtQkbcm
FwwgtUdtMXygvMIGeOQw4KfNBStAZl/Kg7htel1GgPWPQKbOWmUDzFGk1xuOt04J4R8NdMnqMPzo
IGt+RDDi5ZcJUeWtE1J083FQOid+m2/HBv005aMl4KCkwlMBGVFM9X5T7euncTQqB4A4PcKxz8uo
psnlCLNNEXy0+KzI1fPY0zm+bLp5vGsBKiDYfLZP/kWBU7X+VHV2ndH8aSAV5MQs+gzCTlkLUcdN
ThmLqK6ay5ZW59xUVVfBMHiU1eJh1leffxE4t7uyMCp7qMzi5vOWjz/47voxuAc/28KmOLUWi+JS
or0zyCVQ45DN8qmqLVurz7S2P54lsk3Ai+TQJkFqcfEKqVTfj53EcN26j2WvFe55lg1yip80g9Pv
Jw/r3HnTe7kvt0AneLOvFcleICJLHiyscTvLvRJEnuqWTLhTUAgFB+zLl7HSdPrumvTGYxL4li2q
sW88T5pMQD+uItw6PgMIfIsQgkbNa4nj3C3hBB33wdyCJ+8BXcCddbzRi2nhVyFK5ieL9THFYUf2
MEc4URxCCo+gv8doTx5wKc8lOgZs96Chd1BV1YHK/D96rd28A67vY99PROQGLyLj27cHhmcd301K
DwVsYHjgV46G3ZYgDKwsZIM6dJZlM0jSIu39/e56ZxqvOQum7btsNXjGJAiFn1HxZZpk1RTO5RrT
fh9fvPeFCaekoHH+hOryibAXxMY8nSMi38XkNSzKUDk1lo127mv3mP369U5M4MtrWmI9CM1mdgwx
0I/zUzdRVpsRM98778NHiIRTi3hHFOTjThSjbWFEzqXn65pCW7l+AwRsU/eXaLdLFpg6ffhdlAd0
QYe7AY/fkveckxzu+YffQyClEM870YPOMfyuEvpM2csIPy9qIy3DK/s9XGGOuSjjHxpyxXD0PKpN
JTPgDk5ClsTMtM8UdLfgqp1TLMzAU7B7vjSoWxWkMnEwrUItggCE3tx4i2ylG1mYp57v81zg7xf+
f25aMuiq6vVqRUCUVw90ZZqZZoWKMZzmPRxGjepPpfBIRxrxCuqbLh8C9unzQLyoCd3ENO54p9FJ
wK2XwAhE8z3uBO6+BVCNkK6u5efK+LheRCEWoOsqqzIcwzyfW+fOtKgmU9LuUnQ1Vhytllmj3eX0
PO/sY+nPmvFAxM5PuBKtOooz0XkQv7AwkG9A42wHd7MwZRt6xTFF57/fXJVvXDJqF5s27SFkolMJ
+kUFlJUScTEZ/Hk6GPe4pAq9RoP8oUvwc/8eVnhYMPxyjrLgeADcWW0jyqNvNB2cg6W33A+V2Ig9
4+MS97AllbBl59f0ODe5yKaaxG5OrGGiS6xUsq9r3LGUBPmBQd3H3EMMz1m1Rx7QCsXBTbCCsuRy
UmvSxbPvkWY7XdkzHBK/y+jBrlsuZyYdhhlg4ct7H+hENUqxal74dKBohAvYPNuXUVY2J7+YsL7O
TRZy09XU/74jihX16557cLKJj1Nu0UtwFPshige14i6vOnwH4TwdONgfIeVlogMVE6rbn3pZiP2t
mOIXoESOCvyfqJizZjSTQRoIypzKk8CX3SIigo4DcVD/0/+HYkcP+eddJbnLn0j+b+9zz8XCjTGl
yDKj3EZ+COkF4pxR0DVBx8ykxTl1aRSFtKE74BSblYV8gPAgF+T2mNSKu0TM6kcRkn3uVV1evtva
RrHOe4VhnXjJxb01YxARHWoUOH/vuSGEOKjfSBmf3YDreFzz2mJakkhqHZweB1E0KA1QxHbFmqSx
lVZtFDyPP8sJZNZ1aPS9+yptp2iGDTsiwHwf0VR66SZ/XU9LrK7MDlOyPYm/m4Ay+qba0mwpesFW
H3wKQNcjxocg/bhJ3gEk6Mcn5+23erFAL4myPYD1PtrOFsMWeSKqSbYC+qV4V0yCnDLOgAqP5pyl
lurLmcKSJwXCUy2nloDVoe4vFuIfDrLpcXSnj2QMny8M0jo47Kj4oqB6a9iotwOxqGRnaQD6Z7op
KaNSOC1T7UUDjDkEH+Jz5EgG2e1Wy2uUzK9U+ysYqJilHfIDtno3p6h3qDK35y6mM9FPjuUjHwEi
CrpEC201Px0E9jEtNDE0ITiCx2cc6ehRH++lu/dvLH0LiJUgITQssv12yFwxj+LqYI55efJGvRI8
M3vhGvdmKL7j83aHPEeS0g6d5iAdg+WiExyoiBsv+YkgNdSd8WAY6eFplL7AelOkDmQojfO4scOw
TgqO9lSCoev8pOWf+wP3+X3Z2+8SGGyK4L77a4INSJB+4Fm1+Z7LsXiOo3Alg7rgaantFHc3n8aj
kuLwpxz966csLNzxZ9DYLyEhFonzNSqdzCScMhs6OyyECMggHqezGLLPro9jvIJ1/yq0rqiqnTT/
DPBNuGIr3g0JzML3OAE7omP0E2RTCrWDBRj+Jr/sKnfNgfrJ0i+pAPuexVkKxaGE3SVdeVJwV9aw
pyHTuBqkV8S8TU1zLmKNwZhte6MAdZ2DEPSFbeVaw40NnXfWtSy3zYPz/xaTSOZx1vHHdynI42cG
A2Kc5/+MaYjpt32HmMGc6/2F9to2an79ni6iRPWyhho2ECIv3BdFZ1zxMrjRp6OEQlzNElQWDNqF
TD75KauTPKy4eY8QpinF7y6hB+FqwQ0tLnCKTIjzVHqoQkbS67LHLm91u/Jq6ipfyKarh/4YdDBN
SzDr3OJDzUrCwSTlUAwyIKdUIBjIrbUqKkfb36HgSzj2U8nFHSX03w4EYCGrZjUYYNDR6kUoo0Ll
MFoXRPzqCFSethMLzgiPBsxZU8rjzFy5/TIL5zJBe2nNXevvxSKsQ6i0wT8eh9SMLAy/iU2U1AP4
4xucNXLH+wATNDNOmLCWYzb1un6mrLgT2Ofv7/NTXkPKzkI+zqfQ4btBf4cB44nnn6XiTasAurgf
jouZduJKQcM7yC/rJvLUVzI8O+/806fKHgSxuPGGoHqoMdCf9UI4QQ7nq8DT6QC5nmyytE2k+siB
J6nF7E6F+VsCwAaPPNllIVk71fkcww7ecomsJUgqeii3qvBE8thqHFss3dKn1J+rF1+31+mox14H
3iYK14QmBx3+AsGzUI8ROeafnc4qQVfJqzpc8K2xVqMATmLIvlXVHhLy9CcZIo6cyFWOY9rqjeS7
RChB5a7ZJQGx1ST7wAgoqs5iUd7zcHwuKqpytVmUjIlvSoTMWHZooe9KWmXwLHYfT0ObMMyGfd8W
LZ8qU0MJq0IxOOPhQ6oO2TtuQRH3XqlAayr+me5b7K8qLXe/viHMUZUYEw5Goi+7DZAxqzZ9yZ0W
levQpCMyF8RE2w5d7gz6BXlFMnsa5CYhfjensXBcn5JlrudWPfASsS03toijpUEQwpCpzBCThyuo
AvNfviJ/B+fSw2LYgOhjtdIRbvWKAcDuIZRDoQm+RvBBpo8MTZqvd0RWeYANVzLuqVTEo8570Xaj
93ei66HDkOWA7zdMcWBn8dWotNWjryX0ujpqk0ZbiCLcCA2HgTOXFbYzjJ5qheMnLaigGFy+G8mz
oreodDMqs78Xr4DGPrks6WqMs+Ft2cmr/d0F8qRGNaMOWvkHY7DV2zOPG0XNosMNqS6tGNsoHGTF
XvSX111j1cf6dD4jr5GARJ1eg022xZaTGi35IfPj9c2DJrUgeDm/ekckWuSbo5OuoPSG1n/k8BBZ
ZlwcZjoHn5TMlZB98J0XQSeqa/mUy1E81uxMDBY4VV+ICrJE5sSSBEnefH9qjaPVW06nFgrpE3RM
pGVUDtcmLOPYwOjuIVyhDHzXicnjaUmXU1R3cYPdTHcWoh6L0gK8S+xAnAkQe54VYqZm/PPzFuTI
ZJmDhseY8EkDIqjhorEkrrECqaZwYbUnwIsBzoWxp02KW8iJJg/AzQ+zidQPCF75aTQiIMNKitEL
9A2VVh9DQpVMTk3drW+qMVWa0Y4fxsRhmhIx/qMuTSRvAPuGPFZyysZ+7STpJUgb3/mJbr6t3cdp
SdHQp9iuSCMdMt+nPbQkwGM/ZntB4y/CPSjUWR0UCYODAGvREP8i79YURB05bHIE9z1HinvtIjX6
uqaSae8KcCgy6Ue+wjk3iKQa2Yyp9tIcDnz1k/oDZsyr/kCN1jnkm4iLgkdIrluKqLXrBxYIIHob
5j/UBCIPYFfm0pePqaXhIFeyxS/0aDjDV/OyTligD/TtB8L3bdgatOEUyJEupacyaTh3gY8s/ln4
ccT4KVFi+tQUpNFUnANytHdFuunQ4VJD/8uR2dq1skiy7xBjB6JlipGFarc2LCr4aP9vKos541eM
aDPrwG5+uNKd5vOjpo3tMix47sbFdJoPUqP9Mn2r+8x3YbT9GWsxTu0rEmZ9tSyNwoKIfi7yx2j8
LMa9XSJFK/LiJHePiBiyckjvv/POgCBAdVWInu89DtioGOBllp1r0B6OS9T6na71f5jhxds2u8uE
lZCqtp0/q5EhqGT4ErqlL1MpN6wrBAUpUnqsCAvSb4uGIHP5cKHQlDEWmab6qYYQGIfXWpCKlUPt
ZKDrIDc69A6dsEr5mjhyaL9YySLISYfzuoYEUsyHfCSAYUsq7w2tVSfUcfvAk9nQ+FfI2k+ZDF3s
6/MgnNkNkaMheXv0hOujw613cIb2e2QDS4vbkfglmpU+EXUizAse8f+8LH9Pm+iUedhhwKyQDC1k
wjB6dNVYvw6xKJ52qWHp6jwJQa+7lIbRCsLdYOxw3xjKYXyBvNPQZJ4ngxJJGhSj6Bj2Puev9lq8
6xAxWKJiekHv3BuoIh94qgYvKvUQ2werYWUumvEMwJBtjM/Ed2n1Mh1ljiW5dDkI36PXlnhu++Bf
XZHUxbA2F8Zc/JQYyzcNkpDf4sfk+fSejQUB3MDnEqSCfyAEIc6pZpNoMYbCuM9ARBiks2Cu5nEv
TesobdBWJ57wNpE7VD/vUNIcYuS0Je+0/8otn/TPopi7SDmYBoi4ar6PlWU427lWMjDZXTeBTnX3
J4vjfcixEGDuSqRgoKzXoUSaOiExr/YMtcwleypu3dt3ymluhO1Wn7oOXnnmLNYhb5DYgCbol3R6
1Jm5YSXrqCI/UIIjX28g6xSAWC0DaPgIJLBblPnjDAvrzJtAp5NaZpz8hckvDbVnoLyE5L+3bN97
MVfqiOHMD8DGD71l7sfX+qi5kSwjJOn1++8S8JMfWhRIG6zt66g5ySEP5RcHIhz1AyH6MCjnZtu1
F73sYvkfy2/khm5Q1fQo3QlFO73mvWdKMa9319r5sreMtL4yR2QjjRHYUBrKa8giR3+UW4KFPFBV
qD/aVm+zp8bIeodT45tUupO7rKuSj3zLn5cuMfKs9bUlw9PRvCf4H6aJutDHp0hGVDWHUfP0xH2L
HrKiojNuPntOc8g01QIYkFH996pg5szqo2p0zigzZpC/9zN3gwXxcNkFmDsf/X1bnOceZg6MebJj
rWNbzLCgx4dd4MLCZJfVP6ZW/nc6XskT5tJwsxVaDSwhSCNygWxkpXcAWtk+c8eVICFMhGxYKmj0
5ac//DI/qZDrMH8/GKeP+T02x5jdG4hLg3hP6wck7VZX55EpkVZ/tkpzIcuZnhAJOaEjal7r1QGw
FGX25zmtBZyOUcYbv/mLrKFVCpNpez/8fW36HUJGHdxY+R995cq+JGqUIb73/iNvmtcnuAq4GrUK
2Ztd1/PyNgGUVsGXCVZZAsY4HXzKDTmcKhDkKGDD3iHA4NYjq/3URp+p09LYi58GRo5J2xYXPMPk
LRNqYq4LRoQBPw7Oq4delgLvUk272CNEI7m43qBng9kYsRyYzSOtITgHUV2GOm3VpDAOAYs2TJPJ
AGZyAu2d3vYfU9dkfM0dmCGfTT7U0+yte4l1uBCb6oe1x4ozfEoWj0Wysy1xDXBBLKJQ9pFTXJDt
U3beMIlNEOOAn5pA7Mrc+netZGfJGbvBU3kJfahgrVyeVcpVTJXCga4ApfweUhOATlj8aAnccq57
S4JlS+Ft+xvkVu8CNJzYcFAVYQOup/1BajR0u43xpZ5GneFsghVOcajqJWPZZD5uNKR+eJpy10xw
byw8Y/+sY3Vo2gOXBOfrqJRhC7u7yJjZ692vgtplkIUXXdRpoQUccqGVgtLnX8O1PDkxel0xVW96
Air2bXiNQmfne+nebyV8GDjsatpitm7WWe3+H7Hh/IanevCq1/1JUlfc+X95e7Bl2g6j0fpYsJh0
5YQt7BdW/GwLH6sZsfKYOIvre6K8m4+H9PX7ILB/Vmv9R4zLT0ChAdqz3ubkoZtaRvdGEQVlqgzd
PuzoyB2OYq27eMps8I+gBDmOcqPseodeMQTz53u3TjHFdo83QFU/icjanejYBMayE9DhxDDZoNok
utqRZLYKJ4TVyOl1PGx6VTBX/xuElCe3vudVSy727vOie94icHQl0JUz8wVGlitJOMWvWUY713z+
SR8w6lsYjZAki0svmpMGI0sMmtHSUNpg2rAXVxb7gCNImZ+JZ2H+JIDobFul8lqm6gcqktOLg1wz
3Kv8AlvIKYTwBzqd4D80VdqT0sjxWYjhqyZWbKQf+P4K8j3WcVBIC7Er3NaHm7Yxdk53E74mj5q4
kuZMOl3PO0og/JdPml771XKMlLWG+k3gzCTa4scu6sUfth9H/fOBOD1wUEEGBbuAKJwQ0fgNbUn3
01A42gRa6l4Uhn7RwLAcfjkPZWgFNEWKesNdPHQ43MlZf9bsr1xjFpQxlEcTbDPe3f5GQx59coC+
3iwExjFjGty8hRpvn3y//V1es1jbk4sOmtqiI7T+XcvmmFnHnSuj9SWfxZFOioL7x84hZo/pxhgH
9XyBamWRpvrfAjaGPeWgKcYvm9KRLTwI3eRxgeoZJKeGYrCvDbbQuPKJe+zB/cAyKgi9Vj4iBFLq
Vit7vL6Nrmi3yra3kGVnOq4HDy15ITfkJ/p8tR7vbNvzlPEEIhxczJsogEg+hkcgFPDCOz46GenI
os+2qW6H4IEF0Wy2l8AUsmqVybHHVqYCo7efLm+4+M9tBEs68edKCbmZgYlBiMv5kBnJCkxcdJXk
GSOQRnY26NhAGwBpQeLSV+IYN3xTbEwt7fx32tDNk+Q/xmwGJ242BolRi9iibBaPm8LfDBj77oed
7IMwaJTvMPJbjUMZeTWls0c2Hz1LEnCxlQsIRTX2W5Zxl6MW4CT2zVjWh8Kl8NC3xKy2mbWgfFYx
/bMW+qcfQixajq0ufWjVCZk00bqVjRW3bxvjYLuvd7Lqi6MD+SrtTucdLEwVEdL1wHs1lV9X1s+g
c/6N97+POiA2jLFxynnFD59kkbvR6tGzmcjJH28L+u2GxDC3JQI9epFQpZ4JbxHXLoS55TtQ6T4H
ftyVf4jhXPovTwAqLmHmYkGoYZfltGQMWxO7FBuYharfLbpKDoY7jt0JfJlrS/iKPc3y2Kh9KpAF
FYCmcWbcs8SvSBM49aT8wSfKYbA8B88wFiYaA4QPIgqzCmYm/CgnyVZHIB8Ur9KslRS1uiV6mvoB
eOt261mWkmd6ROhwdzWVm9RY+DojBDKDzRqsgdlK1qoQEC61AnZXabUGfvmJ6fGZakmGaPuEqM0Y
onpjSd2hr2k47Tw/J+9mAuM50A4h4yFL4xXFc9szzd6CDKfoLUqOby9h80uAm8aIw0b1z3NwQqXY
2jhNjdGAWoXoCum0cWAJELa9oc+iLjvnpLukDtwFgefxcYZ8HIhQ9svMXkTfEI7YDsdV205YCdjN
8MBcZ0MkKAyvMzFRJk2pi2+D1DEV5UPmGWssg2HcYAd2i6Yjhzx1pmGpnHaVK3Ku63C/p7m92zzh
jwxn6I6qIoyNujOjYddPXNj2dIRd/0TZjS7TDSowMGKGvM7ad0QWj341C0SpQD2VN8UpsGcxYc8B
IOVqv63tIvQcI4RN/JTfnPpHiXuX6tetrq7bmQI0ci2aLN9vn/w1sOaxwdSBnWHuu3ipb0RTnLpw
kTO7nAuXmpEnyXyLpfdS0i5AHQUX5d3SvGtuLWmjSaOIulxj+oZOwtw0nGESVYt+E4ypaldktzo8
rgU/QVztN8AFrZrYVwTg9BFGKLzJDY+FkjLe4o6LJIp2YEb7tY4lg89hS2pWrmd3PIoaVudUHd1e
2f2bBXv559Rpi0Yh/fzX/NlyrqtuzxgLcgTmr2hPpsEHFry0Z55yNvWXNMXvfZglBFEmoMD5MpxK
az+84fRHNYsa6OJymuqhxKBnwGjejqCfZpC/upj8XIv6hF5Z64jGa+7g2iQciTx11fTq3XMn/+YK
AyDPfG3A2qr6o78GaBjwPxiSU0tuL5bYdEyIdIrM3oDC0VI5ZQT+JkKWmXSzQfTOtcQs+R1J6HQH
Zzs/Hm09Z17IjY5TiJW3NaLUfMsPq7cthZZPwVPmwvupOaAPpGX+mHjWGf/JQbvTO/Ktypd1PT3I
XcJ2NR80RUA7q32S4jRs9tuKjGLZu80D8uYVO1EkSEHGSreZxAa8knDja9xTzWHrSe+7v6LSp06b
OFN/NAsfIqpltWEfV/tQo1u/eIK6SdgR6uc1BFd4g0mT0BB0V9Qn2z6AB32lgGUXXengsaIWDXdh
DdAk35D1mby3fi/Mw5bDfwQkb5y5AnkEHdVVdsvuUBpzE+GoxS0pDFHytZ+DWjMNrDxBthCCcnU6
zg4k8MoxbvlvDAIWSEKMQWNhmZjKvO/gqaGCNo1DUI2r81tWtoZzu6JzPKH12VJwKe6MjhuMZkxa
Fy9HdOwPYClAZx8r2kIk4q4JCqDIuHFn2v7VTnizzGjmA1BihZB6taYDBFrbq5Cfsc9aF8da1osA
ey2EnVMYvCDXOElYjCRrwDEEk0EV6sHc6q8VGX+mldVpQkc5ljaGXwtjOBC/ql8I/o0o+BYV0wJU
GPdW5/kgk5BIG1oVR/lK64QJOKjrNjLwCsVxFdCSqwQQJRi5CE6iz5qDbe8cu4vFx4xMUGMjBB2L
VUs+cvQhgXScmuES+RQKumsX7qgJrQ5lu/llbXUvKMXbOQeTQeEr1z3/pTfrw+eQ3vsgyIuC34RI
XCMlp+ffwCNC9mgxDC3SDx7ZMP6TgF9csoK/YJx7bRceBuSsIczkhRNYZyRK7GYONbkY3zPDbPkA
maQwlVkjWC+FLON6jPY8Jx6c1kMFvlBV1krxGNYFPq6V8B9B3E++z95R+pPe/wQP6rIUwnmlu67B
4pPo68rfGpUmVhBs+AX+Dd+ObbCP/TUIxIi+6aQneyedFLQTdvhvEDY9+nc+3w6UkaVQ2xaDqvWN
h4LHBIP8yWaCOSxKEQiEIDSyuDEBpq/ZlGtWRYOFLMP3DCVrwaj4YAjhAyD1S5DBdJ4w777p3V4p
WW+OPMRh5H+nd6mV14uRB44zy3y1gs0TpMgfb4FZXPg1n/a/lAX8+RbJFUfVsUMsV968Ll3TR6ZC
hXYcybRvcSKlTcAK9wsEaI51Z84ZA9PaqRyOySvMgcOMttk9/5SACl68Ug6k8cbnlNJZuhTy2kcf
WK1VtFwz9MmL/WYFbfp1QjX4sjG3vdFCFTTbdf3UMGpouLWcdUvwbtbxBBHuXHJ9ZHu9oH3D8O6T
IzgIMJHGptwpAtrl2rAcYEkduwhvckeeILEWZKKuD2jAQNZUVM0KFkuxG4D5wUYEuwE9DjDWowh2
NFu+rdgPYRO9yLKf4magjSZ3b1XaRJNgbOb//UUibLTlfOu9bFHO/wx3WE/86rZ3FO2pOuYs3szu
YaMozcgfltkQVjBqVt16FVG4g2MnFuKmsQ9DeWmw4wdn/GUZnx6lCrIqOdU7Vb5stk4zWykDW0mc
Nd5xDHQDPa1VOuQkg/x+WkVicllivtVFZuOGN+uyS4RKUTpJHKb1zYubud4inMce4Jjfd1xypYaj
js6ALcHxVTypUdXBG2409x/UyiFeYkmekpQ7CA4qNbTfo9N9QU6kRgrM3GofhkZIu/F3iXiyjYGr
xnIfUcMvo/mVDl06aEZIqVvxSgKzgRGVT5GHxmJ0UQlKJPuSbcF5jvKNaTX4dZVPGqjvJTMK8ske
16C9erbMX8w9i6NvIroQ8qo3bNJQTybm6RJVRELn84BCpELKQ71ntK2zRzdYA+paYJQmvgg0dLn/
0tiYv6SQUic3BYHSivLGkX9xmT/he0Rgplxx+oDHNPDU/R5Ffr2kaYgzPSvAEbVAeRxjMItHR4i6
EcJIXykAZ7PuNNxbUxVUp81R/HX6EC5dv47M3Cd/VmCJ6S90pk9h9tfXw9GwZplmYtgbjZUnMuCa
EiFny5cCpznKwt5fWgMKaHaXU++aInqq5bYgvzKa84GA+eZyH32sr9CvcfyHTCvftId1uld04mxp
CEKDJ3mt1V9NczwFZK22zi0VFMDCHx1kpKsmoqml+tLuhEr3cz2gGTW7P6l/SSpQYW1EiZk+3ynN
Zb88K0lDq7sg/kdvxZdeC1/ZkMiyEZFGrPWLIphhhPM/Zg1gZyyJZeS2vO91YNGUPCN/dkMjuM+I
N9365aJUzSEqDHf9Zci9dc36gLR2/ld8qTFg1SiiZuaeKj83q4G4XGxw7GnXsL5eyjYc9YWqLR59
F4wO2tt2zMUXPxfpynpQkUVfgrMRbCYQhlE3i7ocC6UbMBhrnjA5qSErqggFQyEkkO5jI6jFkfrQ
c4Y75ss53fRwAKNVzg6g3Xujwon6mkmftxC15xJkKpt3CyjXQwKFwBji9uYSFJ7PMEKklk/ClauA
A4Sbjfw0O/Hi/iQXs5yZFwcIHPU8d4TJeWIY/R8RpJjLT4ep7n70VGoriX9wtgI2iZ758H8kxipZ
CscZ719bh8AueCn5EDPPy82TRFkwZgJlAn9VlWzDumqbjLdhVaINTGT/WlL0oXUR/frQ/nQ6hTrV
SYu9XzRTYNUpQEMf7cAaF8py4fbJACW4uo/MNS4AH+YQH3zRSnmLkyc82nIlpS3eVMphTLnNp5f3
e2lbuZ1qfyUM7Ff08XUMNDK+fp2bGxeDVK8x/nvHIamlA9GEfZ+gEyYOp3DkwMrBkCykC+NwhynX
J3/AydnaItdwVem6wB9bwqxtmM8CQac+0jPJddGpaFCo/MrC14XiJR9jU/QAMVzGJrzh9aampIot
1ifjHojj2b7tT4yxOK/QX/s+DMfJi74hPGhazA3s/pM2lLf53i0Unkd8UJDR4P6mt8wUxsU56omd
spGam6pVULPs21BqqyBUahmi4SW53MIPshPjybZjT/lVhF1NNEaLrCWuQwLP4GNJrve21l8xwHS2
74YT56JrfxGkQJe4k3osZEIfqqjLt9cQL+scF4nKZGeJ+/9QrzHamI5t0qm+qhp8/yPdkl5Rasdx
gGJMHMrdATljnTI6jVcbjibfl8EBilKcDQnBNXGM5rX2bTEkbbNtsp821XJGNPsiWigXY5xEwTkb
nW78+BGaHhqvDNy6I/+LjDj3S4zrf7ufLPSaecsMDAxL7sAM9YjNRQ/rsS3MbJY+KRpF7HId9FMk
KAuphE/Li+gTwM8xjKzNiOeiJgBGt+u36RUeScUjNfrCxez3Q/jy2wWWltB9pHvVyYnZ/uwSmcPr
5enzxlXlv4YuIpX/PPvFCRqQ6SideRX16dq8Z0EqBtXJvG/mZHSHegwlO9xWw8Xd6Gsk5T1fMw7W
fa5UJtM/JRDMy+mESZh9TRoZL3IW8XXH8ZS2vAwm8hXQhXwtSPRzPPSoMI9N/d8BKITqi0WZF5HJ
JMCi+XctCIylByucSVf7tQN4a+lXeCic0/1xNskrPmL9Bdsb9CFW39xgs4gOYpHxMZcpDTh0zFQ2
GygmLkph1nrsQUfEb4CLTxeo3cC46gxpeyZH/m1SEkS++M8rrCqmNI9K1AYjvcdxhLyEDpenvdL+
fBNJZwC+MhI1phqgWEu/je00YmtDk08G/A1i7dZmYIq/eZln5zhpbkvWE59ZSqcrwfFOWmVHRC0f
9kkADiEGYHOCopTbgFllz3cmdSwxUmbwofYyi8N4TaglwEntIp9KGrykU8bdWCazm6Bb606425rh
AJMpuSpmB1JfPZ//L03+j1GDhIbHUdIPbuH4gts4hpBbcU9ljFT0V+YfDVKHBU8soz4cNVhxCwpJ
v9ojLi1qzw7hBey0j7wOE2MXyItibqO68iV2oSV4MdkN3rt1x8xuNAgKwwhfMwocHfb3RINY4MfC
20D5QhqwnNDUaaj1vYfqknkA5LqV2QqBk/o7+/PE4nB+i/4eWhUQd0ZcvtLor/VzQKUKlINrUkPu
bXP+Lw5XLq8ygam17WD54BD8Hj/XfTvKQKb/ff+v6Lhk5Ro/SyXXygg5J2PFPlgAEa87uAXqcnH4
65HYGOcCmNz2QYvtOpSi0bGtVwH3N/0vNRNSnj71EikHLsdJ3LLkgUIEDQ+eKCeJqiFHqHW1s+0l
iWg3dfhZKneCmpaVcOpXHRtI5rwB7ocsScVOooMwxPu/yv7A/hY1HEwWi4tqg+Nd/yQlgPweh9i+
2eyljIulFr9e39wy9W0sXKrPP4lw5v6Vu15mYHYeT6kVtKcAQKoNpQpfehH/+ELd/PSKOY5wrMZa
yPXrmMpPRXCWbUI0lQGRLmG7gEkeqcj04Z9kqH4dIsfQBevBF3oXOJNwIEem3aYKAj44T4uOAtzZ
HSZH+xyBnjNmPGVpEyziThz95nnWQcE8zrtWNnY/wZYivWom8bDLNM+C0FZJnBEuFA+8AXluoCU2
LCgZerEcI/DAH/7TMhzyDCgvCr4z0HSbqgXslXZf0rSEYgcxZxXZSMvhksCoIu0wnTj7HXYmveSD
Zgqf4uirLR+STJsjGbb2TXC7zhjj3kZ4FL8R+DcMdeXylDu526JMgR/m2PGV2+IpFvtwAwu0+V9R
0ZfR5Ug3AlL6GAlH+OYRDSYcm5kQarnMNXDhpQv/yyp1x91c4cngx2ALIxuuco9QJikpJGQvFBaM
qsz2vfB//GYmes2MzAFAhP57kMX4xrLEJmkAKytae21GW64QvvE27P2eYUidLQM3fhqJAKlA0hR0
NonubvxFyQdEd7mjOrRUV6mPIT78wW1zHOGav75L+f1RtcDxLdFisNuIMvBg72W+jc3DTshC/7Vp
hbsi3wp7R8tggv1wry+TGwGixAG2sPImmY0By3zvuH42AKXq6JrLg8QdwF/qXdFQL3nV6sYYAxtn
4hzx2UXwHJM3tCvj9C2gjIpAyZy3qCP+nkqpH9JaIrtWws0ToCry98/D5gIg2RIpLUb8f9K4ZVaG
1xwRn0/H0ogA9E8Gz4IgVG+lrFxMN79RK2oX9cMWuRJJ81WLO1kVnU2oUQ78ZNbLlSu+KPdtA9op
oEY8C02SJkEd6M4PWtl0qKTuJoruIOW9qHhydOwFPtj7NKu5qYBP6qMLeDXdKebR0XZ28NH/BJek
+h+HdIm5Zli/i5aoOcZKh+oCviwXX1qjs5u4resxUXcHRmYYOzwxD8rjVuSWq4z57xxjvQdQp03y
53Co2QkMdeLL9BgDP5LI32E1HSsdmzp4DvSkrKIQxfxsPpZARyGyZMNYo/hVZinGSbTMz+lgW03i
ekSsn7KsOoRT9k0XzUXJIZvvv3PoG+eFRCQ2A/2NIe3PSEhuQsfFQCUfV7mfgzIGSF5yRxRZAMEh
NjY7eb/YM2/UpsMk57AOk110pJ3a94NMTIUuJ0Xi7igzVxT8lI+4aiAEeagt5JFmaVQca+P6m5ku
/khIN0eyTvQ+WFvka3p7eVEPekQrujhTXC0hM8XuVb6nJIVnH3iDILbjxFdVDTAPUS1cRFL8wmEa
EQn4oM7+KlnxixQjhDAIw0g3+DpqasEgX1DCti/6ZUUSto4yHQLm7aALHjF9jMe6SwSerUf4Mxeg
IDGAMmstAdclXrj4+I8A0Ji7o0BYJPdHI6QFj9/p1HRsrkULliEkONIbMAnEWRt0lq4GBvetKujX
DEiqneEpm7kVLnfs5oehQLyd3fg2lj411nI3YQwckp8Vjyk9pnmokSOlKhR921VnqIEkH3OCDItf
HMgENdKDM3lZFrqlfCN2LbG5vwl5+VwbnOXLvWyc6w3AkOYpeLZ6sy53us+pIRp6OM0PHT6E6CjF
fkbWR2OchGzpCigYUTWqAqfI9rsDazmxlZOr3FjYLbgJExas94bhwp8w9STcoe2hR6HrrRZu4Tn2
pupzqdrjSG63nxorkRUlL8ZEvt6gHRzyye7fAqBgOZzjLonVH6cDZqFxaJ8gup/Q070hme3LdB+b
O98myWwDvNPs491TpIEHS18xR+R7n7A84RCdH4zBQg10saZN1GnkVKbvpsT5+P2uxmt3hbak4GGN
vDhrAnBobWbxmnezw5sWN/BcJ542o7hoTZwE+WUZUaIi437PvxobwhDCIEkVHF3MEBwsXY7OY+WP
kkjeGIilsTJNfJppncWhBdCS0wvsnexXE9SJR2d4EH1VSQ3boLe5vRjm09dqHhkn+kJU6qm7eXil
fqvwlbuR8O7CN2Olfmblj4QNVqSHNpxN9mWMx6QhYgZGdtgM/WRQstcbLVDNEZdJ18Hh3QbkVrIf
S4EfmenEkNnmENbGXddDgauWxu5jx89cSPw0HscFzbnV4BmxFDRImV122oJZ6EmSxm/iIVEqFSlw
NYb6swmDXyVk35KToYvKsqf+yWkXiL6oyQTKqR74HEtHIdlj+GUFiznXOputBOTbm+2mBcCwkpkM
gEcCTCyNIdzMqk7iJRMddjQjpfNJ7FGrlm5NbaUiXCR/hnGYiJvIkccJ1pURds0/WYvD/0dRIJXJ
jb/7/Cy73H9JlE1VDMFeeTEAm/cf/FTwAawlbfG1iTpYVJYFshpycsc6mOcZeA6e1J0wBr853MeZ
JKQvcLyd5GE8VXyn30IxulE9gDY9NFA20pk1l4l7m2hTPaULVq5hfSRcuN1EqGnGG+H3qKI4y41R
btByFJheaVXYqz7QuZOEONIrxHi+GHYj9HuUteyu1vXLUt/yCiFlb+HLPs8YJ6Tri0kLw+z2Y9HO
hai+gNcjLA0Ni/cKurQWtZwQRO6t6nkkO9ru6PFOmbevAXUAO9bjNKMlVzMCQeNhjh47q/uu+qlP
chnOMGOSrnrFvZLQYmWfE4ZPtcxFIyIfq6YuS689rCvTYBY3Toa1wtnxBIyRID9raf6GgKgHL2uo
mPXcN0V/THEP+st7WqhSRpZA6UTh9tWPy9ZkQ112acO6zWUFAUz3ZhRMhWF+VHGhQ86/xq2+EU4C
LyWBhlrK5DR6Y2izF/HCU5N0vc+J8rfMHxR0qNTA/6U6c+c2POg5/b1pOlMLNVdCGpQzPFvMEZW5
oViv+mSNWUfC11vFu8ETqQOr7pFsv+pJF91XUb10DL6u2ozGgmDkw1FhofCcx6ix0OOxAkEXeV4i
MFqdMNs/UbG6p/etnIbY3DpO6S6Y/IMomTvTjw8wajDVxKSLJr4a/gM7SE/4ZOzhLbXbku2LJNv9
26hzl88sJO/Ot0HSZgFaq/aGxQau+JezHcUcd/o9yTSVSBjXv7OFNfI8ObbyAgpE+6/CExIa93xh
4bBTVgG5OmiTkyiNuK9xl2YPjG2wmM+RfxKmjCwAltPnQJMGT5BuWY1hd1pdesyu9jrjMBl0jwho
5HdUKFXsXFljuw9nM7YCr0mPaQPMO66hPt/vuue9fLnAatxcIg6EDGh4StP/IcspALszQWUdFcI9
5dOqWe8LVLJwPOtcMzi/vcGquEshTVLj0/fxgqLlhkFK2y+WKJdIT2LsKDuMGODHuHUkIr4UxkTu
pdz4LXD9qmJoXpzl6nzG5rTXB2iULtlT9+8iNZG72tE/VIl583+tENcS/wXMMMonTcEsbH6g3M50
AdAlrxKHsF7TVuzbv/UyApSOkbmAvIcqU1v4F2FrYFx4xmoe9mTlvIXKWURAgXiw2TxNZTGBrn87
F5aMPYRQvt8n/Qd2qXSFa5GGTAZUzVOc2Wy46XWdbvxMmzrB83+NVPrdx6a72nikfVgYmFs+KCrm
MyVfyc/Yj/x2iRaig/rtgAPs6pebgScHWQPoJiThrUtkfpcGeEpAwcr/X9hieLf1cufZaa2IbSmP
fVz/UKhueWvGQonL64lxpeGGHB292ldq0tKhjJkWLIXBCdCaK7VRThG8hZ+XDSde8WXhSoAEEUEk
ZbomKHhzPFXNI0RbeBb9plmTaNjyd4sW3DPMXwZwvPxy2+mmee0E6qztmAj3M5VU170AOBCGQZyM
WCtcgXCaIucpff01jO5d9OLxTyWtEJAcx3N0OK2EEpj4Q+0fgGvtQE5Kw1f3UK3DG47IBzAa2nXM
XJVN4pSzBZXLBGMwi6gbsMuI7ApNqHxo+DbGH4CI6CXG7ilP6JPEXgOn+MzhU83JyA5g5efEDw7B
nppsQf5GkdzC4gdHXwQoPiDM0TfoNJ91CPSUjljOJzGG3B8BLy/XtRlEC0eHZwxIeBOnwcYpCjdT
wUYcLkAPTQpp0RMGfGGBiks+Kv/UuA7E9M/1hRxN2e4I1qnrz81dBxdgOGV0hZHtYHiUu90JIoTK
rbOJ/pk38m3cTGVjA6HOuySu7sE3m2pMSvJVbpFjISrdMvu3MAOVjyW6/G3G5Pbd8KGzFSDn/mbm
krKYQ7M/020c/ho54TzgBm3QeS7S3SdIzx4BxmbkCLbKlWoRXCRcl/aP1Ny7mVRymK4/+DjwpYCf
zIrxTQgNpBXpRKO+SZDq9D7a7hP18jvwrvHS1ReaexxSCPg2AGDIdxtWdqf8RZEAPFN25m8SQPzG
VLwdAHGO1wlnZ4zF9q+pj3iBKcWwzHhU6S0PE/cTTSnc/3nAzOjQ1h9rRS4+dKWMBHLiHMsiYa6u
Poz23Mt8UWlqucZCnawOGRZByHNob6ZILpknJa2L1VNJn7ITdvrKxvJ64xwWSmSlkNAyLE5jm7P9
QCUW3Vl5ffqH6uI5fSQ+L0nnmc/n37otQJvHA2hbr0zqTm1X7pZ4ve/Osnib44oSkeHXsWXK5GXc
EmBWRXDaS4yCYOxgFMxMqYDi7l8/yRjnGd2qEreqGjPD5moBhJ5XvMOXZIOWxu6NLaBT9CisjDtQ
Yk3ruoFDzcWTBTYvtAGGHpo7/T6G5VyDdk4Vcy1UietzEk3iYBu/TgPyPEGST6fO8+Ov5Cu2eFi0
8twENEmkwjRNdmYvh3Kz3kie7ArqEqB+3D4Nx+Lw9QLT25WB9qGaLOI9J4oBEurPnDwFzXAW9Q5A
4Ma7kfxYNfWkMS+3yWX1Oq6AVfWkDdTHOw1QXsGF7aT8017E3fRQhL5oH7q/NXpChedsJJnF1mOv
cqp5xpSS+oI4vDPWQ+7tDlQspfLEBmq2fKTtDrsl+tbqzixNRvnXvOXSMIN0ooepxRQ/UlsvGZzv
2Q1Qc0/XtKgVu0WoJmQXzvBpjxkGgJu592FmCX4s0ll397zqUICq4hKN8ibtA752eqkYcpnkRY20
61n3FFf3OA4KWxuFTLKkkEzbyR5oJ/Qko+spiYGtbyAmmOqUJugy6A8utIl/Qsw1afPZxdF2e4o+
oVyWFmdVvv3s4EyE1muffsHsSvuqsFtfwM5+CIbMqs1lpCeSl6mGPwVVuxjf8bAoTFBA0bJc0sm5
gFbgPGMljhT45p1JTjDltxWw0Z30lXHzH4jbclwK0WoaC2PW8WbBHuQyFm6hfIOcEamNTJl3x7fY
l4EzPlLDjuNHqAhulG0uNkcwOuXmlhjiGQg41K/7Afv3zG1fNQIYUntq9eRdgm4pKrIjOHQIzpOS
PaiQivuDHUPdbz1/BFQc+mimbvgiO5NAE1Hfly/YRN99bVM726kiOdwo0TAoO7amNk2ziAIGvjlr
RC+T0xnwaMWBJ8GJ75+1uPlLGkhR+bhft+0Y/a4DO4jrf3V0lzmROnlX79qMcyq7hB6MqjqbyrCM
nqG5YDMQ6ta5hLiFWr/yieKqMZgA0PX+TkopJ1KjZdkZxpVnxBTNRdUPUE5/38oaYAY5SKzRTxTP
Nn25JXR8Y2JQxCxG/9A4XYNSOERfAhO/HMh9bb0k3W0oAyWZsZiJ5bMm8p68r43ceV2oQGwnyLS4
qUv+G+5QfpKCS1BMEnpWLCkF29ns9hLL5c2KjXwnmFHTZCWcGGsByyldH+IRTQ5gTigB+p13WZnc
RuZ2NCyYgCkVbKd2fMMTQt9LjqUi8SMyXcyHSMmPZ+Hn3zvlWnO2+RWPldYkUNprQaStOp1D7y1Z
Ic1OkOT7cM9VMZCi2gLAY1ICFydBXo6kuTdwPZD4fySikTg+a5Im4nCjIHir15hEITlDvNmhtBcr
SanjKlhfdZHd0XBmoL+UOnLK9gipNDX79Fmsnfhw5wjrTjKsqgvOfDF0jl0dVDDBUr9XwoUstNrr
JtbHh3tiHb3h0Z4i1398yOxMQfIpNkzuykRAsEOshJuxA2kQfqUrazMviVofAxcoebu3VyRiGyDz
seLjEeIRzgEXbvLRMVh9vJQiM1JuPNIupyxC40eyqapHXFyhfU62Pmq1xBHdVIZn4mVybxn4Ae2E
GKzT5+qrtiWHcYXoOOXS4kc4O6QnS2RYgrjazUcPF1ihv6pAHaNX/c7tYUVNvTkHYeU2Yb28FKIO
BlL9c7oJOFViBcJdfexb6DSCr3RSBv3WGWsUl5r6sbI+JNhTlVCIMpzhm0mCHeLxwvxgBd7xjrq9
smqwspgjQBhA26KHW1ZMzcrxSRrBn3Ak3MVj2xp0BQRV/brOTnyjXQ4b6p596LPETkjQOsEzxb9J
SOUnFqrX5rzs5bV9GpKKvA1LDxITKOdl8CZfWwMw8qgbTFMz+PCJrC9dSeVKe2nMhf0ZWk90AuDz
YJxXpylQc/gxGoHNKuEnNagU89fYQWVvGaVAryLVxhcGIGzHF6jmUlsoQ/EfBLo5ovtAmTqidNGS
Q9UgS6P3HilLRhJCG0+fuNqWrN1dze+hl5POhuStw4cw3BP1T2O+HqmVmaB1Vxr15QvsZZ3T6XWD
VOTki78BWVeTEYGoLt9zCicpNkodG0lsPSBOz0eelvvJ12+z2oGTuCP+mFW25C+uSvl3rDG0azBH
QwE2SZ5ztqtACpDVZ8bGDXt46Zolvi13CT3nqrP0g6+wW1fcOw4VYlA1DpJrbSAla6VCne/Vsf3w
fyWSuoF3U8kSDkkCPSiBd+GXK09Sih9dS0E6TvRMqOgJ+XYajmK3Zx5NgANJfIz9ArIISSePZg5K
2XVuN4+6aJ/rZi7b8WujOhE2LHFd/+HhdBOaKkJDsOTFemf/vuuDB+Pc/H49N7pus/IeChsprMUo
0fY+DoLZWqS713r2EYerDWoLc7xWAm3K70lX/UCbHAjGTlW/K8WJG3tIZsmiNGcC1w4Ar7FZpL7h
cLPgZzYiCGVIOQE79AmtHoFlsYFqSyhfILIh1yZxu/O0EIfq0DyqHR9dOZl7tQEhcS3QFrdc3omH
O854FgfsaZRtwvjez9cqCRnj/sztXhoFHnUNkZEn39jVeikxkkI9HKpKNX/ZEtkbNhB5+tl8EmqW
LWeYW+bmSpYRwqr4aHStS/25nTSx7tIP8N9NE4/PlZa2OP+y1JJsuznuEfKRPdYSlAqtOPD2r5eZ
YWDHU/RQjAQVYE0Ykg9IAX4r28tTxa789ydrtaX/xplBeM2w6eMxSNNB/EQqetCBPsRrCiOpB7lR
Ir7BoXndPdyHqN1UG+Mrd+XV6A5l6DBLUCbatF4alkRmnvohzFAracqJKLFbG/A0kBFTs5wqItXV
s/z3B3hDvZjCGQvAFiD/bCWxG9szzwfJIHK6KJygnDcrbL2ZSmd1DzoOPrOFfrlq3PIUMsVAN3Yy
3ZlHBt4vxM1PZwnwC8iA6UTzUU+yzR3EHIjqS2M0ogkSsrqKbBiCUw7u2l65QEc/fp45qCmFDcej
7JP8nypwGkJEnC7dl0zUBcfQbfP/WmhZcgcVl2sBI6vO8hNvkxvlNFV8NInc8E5tyw7BTun9mkc8
WYcS7AhQ8VYJCRhFU9IECeKXkcajyax39qUTFsoHbT4ErJQv3p4SJdRCaC0YLNr/Rgotrg9DqhW6
zhEQ5Q/MYJ+GH5uWWIXh2doO+blPYrQSwMgV5NhfbatlKQLd2jpYPJLKi8IU2dwXR2cTuP/7xuvp
Va83VFfQYZYFWqTIZd3ItPBW58/5ESASLfgZ4CE5aD/IHlmOPRcd4MJNLVGJ9j2rJ9nqTJQZ9vuZ
aLnENrUExukjYKpRbR3Wb+pQpFT1UmvE+Xt9W2oQTTkCLKtSoTmNy8aZae49aa3vntUAAJltT/uP
BTzXCgFjr2rgFzZ+fv3wTWfDr8+Tv7tlc0u/brxugsPCE+yk9s5mcLGqufdW3vZjD+KBrq54b+Kx
g86wzN4BkkUZRoSO4v7jCi+8AnGgSnLICPdm5Ye1YM9PPow/nEC6EnwBZmFk4l504ZyeUaDW91ir
K2s2s83ZT95YHjSVUcajTiwDKmHbdVfQbROCgPivEHQImFEjh0dyjSs3wiYt5Dpf7IRWx3GFZOzx
GIxrfaLa1+nnshogME5WlCYbJT+fdOVMSE9kLH5mC801q92ssaULvS4u5UtALjksywyFx4waUx6N
uk4plZni5FpnjE3dudCpLQIIlEhAhFhjy0kLHe7settnchWcELOxtQt+wG2zEWRGC+HRO4NCuFoY
Loyoass97eF3ETNgUTm58xx+yYx3LtSR0Yrf1NkrAsJCONhjC+Usei63PHkDNYi7JjEKGqTIe8Fc
oolnTTbbj2QP5AqPhSrexnHfeWKYJobRLPzBNjH//MbjK3OzDwCknzcrMp0JQCcZ9qxa0Tl+h1lh
cGl0SsfpVc3C5+b4KZ0LVheF3e2PwEA+UL7ykV3fWXnLE5D/TxGk8IsILoAil9LbFT3MHxGXTdOK
xzEblBi5w2LXWFQBVAm1XPnozrD/QCI2zSV9YkSM9LiAeBP1b7hyGYx5cX3yOO0y1JlMc2o297la
Lj08saJilP38W/QnYbxO5X/n/qDDet/ThFZp+tHWlTSQe4u8Q955H8/AdKNYglMnmTX0AK9DUdTb
cVXuWA1mdFdGQFG9ay+2Y1aVlB7N74UuvB5epDCnxEUpEq9EDplthUxikgsvXBeUEy6tsleD7S8W
3V5xNpXCrxuCFTGm8EIo4akQ+yzEE4vMvtuptjXa3gZdsw3g9TJsXSxLMvnaV6mDRfPmRjEblMVi
BJMHgAXqMnz+9wml6qZ5MPZoHDWmdzAFBbMm7Pp/rcTWKWizXxG1nhyKtBN/zxTpoYvjFf0t4l6b
bcoW2NYQiiIHopWBqfA9s1OSkiZjPJAXwD2B2aBHnP9bVy1Z/4g589NnF+mrZH+NVLocjVVpS1CJ
T2vaIczInJE/QH0NkoeBOpiLjOGLGtdCvO1W0e7vbmupWb96Hfoz290zR6KWegb5IcWIkjUj1qP5
7WDWqdaQoYO7mcCT/SpJF61ws1TO7pt3RQ5/7ylSV8t0DP+8CMLxR3ZnzXwGaC1C/upFApDlsXJs
0Uttjdy3XU/QW40MS5+VVCm40EJU+Ni4Rx7QA00x6esNh0vt7c4DFquOld8C5fyqdVbsEv8B72K/
emZ9cYfwlMu9HW+UhqXTXnHHk2IRQU6C352KvqfTsdMtXE+6KxA/yqGQEazkmp0HdfxPnBNZELG9
LgE1F1TO3uVGCUQ86EjFmiRy/rqpvnPoAgF/drdR2ucRlsd9kze4Gq9IJryyXuBeUoqFo84Ur+mb
fGp8ZXealaC+asT6IX+UXohqj4zscyiSA99ak5Er8S4UXIEj789+ReMe95ImrDfxQTK/LSYF7OZA
kOb7gAOaT5wzb/uTWN8SHbOjOhhovWhUliglaJcLYZgnjw9v4f+bW9LVgkmPJbLT6Wm3hVvSNAB8
FBY6xJp3qqVyCidQ8FcJfyXobwrGeMjT8S/EVpt/4spO7Jdr+yo4WN3yecEwbRAHy2GidC/sLnRW
S+lnpzaGxeyENoaMCe6fTvFMrE5gxOZgrMXYXaQc4E7ovBrH8fot3yCl4GMlg+7l/AT8nWHeQpDe
315XXC95/wvjIlFRsgDIN4tPiVXGrLkOY9wjIqHzX8KFTPUOBXMnyguclQITYiA+5Ik92S6xBnzP
par0GmMc+vCHGclkeYbTaoVUdEFJWb/lUPqDBJbeVAABjWQcIma5EMcJ/jmGS+q/auFFmCRSUWuB
a+mOW6Awao7Blo0Dm7lbH2dP7myjSwC+pU2v2ENMJmx0nh54cg1sczSc3d0nboce9Idb6zTXJ5b4
zEwpWMBv+TteZpPJyG4yKj6Jso0rpf67Xs9CYXHy/kjxcklIYViYFT4BS7QExvKKOCjki2aO3G48
9rp/Q1MSQb3LeShNKv6KiK67Z5YakQQr8RdMQu5H+h5BNX8RG7PsidiKe1hEjJBZVWdKtZqxU7T2
3/m+jQtp9UeaVdOVcvZICc5Tf2hsaylj5t7+qBGmVHlinmEyff4HmOHXGLnHEoWuFdOPWoOniXMC
fwH+UD1e1/HapN8bzrjpz9K9AyOWmfXrBqo7xElpnOtsOqOrwNgfdmTD3Di8nzyLO3AFV06BqIxk
AvHzi66L1ZqriWGQTPjB/eRW50aj+d0Vp/ChiQsnGWl+aocq++bOwW9UP47DGzv59gMQ0KsTvB5P
uzoVz/ofPc7OcDu5DZQRW+dm0/s8hcApKOUIh8MO14QK40BMys7NZQkO8vt+34dMbdr2NrAmjlJw
zEsl8Kad8I4TY15K9mG3mAXKjP0cLn84YvzgULcGw1EoWY1D7x5MBCz6tI40syWHnmx8Zp7HxIOs
+sQBydZTghDJ7yM+1UtOZ8/xoRvMyI3SH1tVN3X77USOgtUNhTeABaBOXLlmZpLR9SThFWsJY7tk
shu+xsrgK7EKceuwGuNYfe0yrdWuSv7OE6+ZMHLUzgxaWae7FG/9TM6uip9RFRj5Z+uLEdLgCqRL
/b5f/pn9hSPfFPki0UAwjiZWAU2emKlDT50yvU0THZIjXI/i0KO13o1ReP2u/1HmgvK1ppvOp8DJ
kfCztA+dW0SP3i8WJOiD8y9OVbfnTy+aGk7yMydt65lf4rvkh7BeFPIF4Fs+8caThz2Ec1LUptnV
NhkaaM9hYQjebm9XiFrf9TxFLy63Nw/H+QMRgtUor53jSMTNPKScEiPCpvWut6635+Kv0PD/hZF8
A+4zLcKno5g62RL4ERe6tRpXCBGM2uxb1jdA1G3p2efL2n9eOA2ZyimilZdNtXu1XaVA+tczFwFv
y52shiHU8Kqneren9HuyeQD791fGooZYcSnKwetL5xiBNidyPhuPU/V954I9LLyRjyonTgB4KlJX
1yu6Xa1+ICcUNye7CARO/djn3eGog83n1H0RAH8kpwm5kCY1UkdaVLBtyA3Wde9vrtesE/LMDMDl
jFpBHV4PfbxPuGLyRMXL1+LewSu1+tVupeZjU+heh7V4zlbh0PPY4BzoAZ4T6t29Z+374iMnd5YI
sHiPXsRPyEaGGHBgO+Q0OD9KTeEhYlIYWHXUdocktcETJtOktFTe1gEw7PS9Rd+w0bacXiB4ikdS
D3F7l8CYsBpXRKlq7TVALOH/UwNYNjr4WcDUQLjhySsbMeVz/9kHybFcm2DtCaF7pQu7JdKTIqW0
T3X/26xygLNPFmBGL1qsGyEvaGdDfU3cboixYhdY+gWl9v1BltyDBnSKe71TrCzR6K+a2ufGJ5vn
RjIMXdK3vl6ev1wvmgc8GD7KpClOoCKomIGHji6PGWASWWj3wOH338YyHmCLZZRC1771jncaC24c
zILPLA0cWtxNWmFFwgtmEqGtGnD5ANyqqBxxKDaCAmUDMjGmC5BuY1CcYOrjOwjn4PrXaWXTDT5I
FBbETN+9FLnDIdK0yOfedwjLiIBd6yX3FxOFlpStRYR0NEqBFiRapj+X2o4Po0Pssmmd24I3lm0a
4jOOFLdVqc86otfkbFt1bSqW8aotU7VNzfRK0W4CTmezc3ySp7KoOYpgtvME0eKdRdd8ShHYg36b
WBdpKlpQ77xuRfzQsrPukF1hYvLfzNH/LdCX/YMv87zs2LZwon77OwY4DbUfonXFvJ92QGuSj2iB
MWBN9l5Sh9aEagKwknnFk4h+6/KgaZardlnUCCJ+NMtnaADaPUA7UraDkgiHUhvVGiwL+s3FXcHA
HWt5WNohVCrQi2ur+x5FVwU7HR1pOi6jar9oQTrPuBk3Tocxz44Hnxsr7D4KPqUYbJ0VI2uvakQX
nvwHWJWkrmBOsF7nHZGh1ysqQEEj6oZBVzQYUKE4BRfGowWv46htqonqsJFNuXl2tfCoJW3J+7mZ
RW03hkE3Ld0xbvbLeeUG96+oiMNPoiv6QU8dMFlI96agcWs2cgvlkuETNQofb/TAQLqeM/3QOSFl
Bj6n+rwp90ybTNAj1HatBkkAzkL6T6yEmF76E1xmDTSRTf3U/eByroERjvuVjxVhpWIDTqLlBq6Q
XK/R6771LYj3+OGhoyn+BMk0TJInqGKimrzNXsKmXIPuR/qpqnErxt/TmwjVUpRn2gy156s+rB0R
FECb89hzj8LX1QQsy6xXU9gjy4Iy/SHideX7+PyUpz8LjbLcdaupTALQHIyEf+XcEo8Ceqwm2R5H
hkx/E2/6dkhpVTfPJwIYGEyeAuw797yJgF2NTni5slLvHuVAG4zQTnaPIpYan9Z16SQeCEbWL6MK
m2m8QUWTc0u7wSsOekH5D6+0b4lrrhPerTxpiK5q+3AUlYpmPHh0MbQzVe9rir5XtQjmh1SytXrC
i7nZT32WgUtbdaFR5jG9HsoPm4Nm15eecasjbq6Hts638l/uTqXurZBqFSV0r7QRu3Ht94kO6K5J
C7h0sn36S736V8wo6MOP/eUdpX7LM7dZ0DdY3JB/G8p39xGFFSGzpPyMe5CfHkitdRz0YK9gZhA/
rAMDJQOiTjK2DVg9yPgLfKiaIexlExxb9qxu+jH3Ud6C8oK+xxWZ6QNGR6NfGuZtKM59TmDy0CIV
/pGsDdyJXaEwj7udxzeAf3sFN+PgJnFUu4+Kaj/PdwlU3SiyxdwnDbJo525VAndxk+m8bUzCRQ3b
qRlnjqc34v/6vm8cA7bLHfwJTxm+nUMWb46aWP8WOzJxy1BoxdK8SsC77kLU1EP54GCidOF00yCj
Vcb4mXQT1W96gikWFimqub0jnXYsHXVtZGQo6nsVgKnqqws1DoKbl4sIVe0H5TJ7rdpcbFCEieN0
CkFE0BPKXfQhpUwT9Ix0ym6FaMvFpNI08tf6KNkMidYOuRbsJ3XSXVRxdYvkQPAgFnhdMVwhIqAX
4vxKZNJXh7252YBR3m/uwjS0qOZ9rKJAAsGp+x6+2SsqfqOIBmGAZl0e1OQp1RBbbxpOF05wj8Tf
OswPI31mtmatgwPBcDd7p9nX0XieSQJn6IyXcRNJYiAU2bWq45b8Z8kXXZZLpbzwxr31ZWHNbvtK
jJ2o9lHMuqoLAsdCtVG40eEjOXGt9GydnD3cYK3m0TCresJJZuJ711rjfcFvAsF35DmdR6ZdYots
Y14YkDNt7HDeQG8MrikEdldueSs1xQOKY6JnlKRh8Qyta+DJSKkgfN4NROI7xgHN1udvyiCySRq+
jIwOK/c0VxP4z0oN24VdhTmPKT96TfLlwjCCc8ltCdEgfuEKPi0DpaVLonoROuj2yOkrrEkA/TzE
4Zwa80bf1mqRtUk6S1sURmpcRcrtr+PnQklMTsU4ZK08FKyQj5bFM6Yfv3IF14Gbezvmb0dh7uL2
3zQMi2ncr8FRAViNxYLQ3xPaQ410vGIB3Yp+BsOA1JgZ1UMmPnBzUD6Hbf8/SydLVGLxittc8uJw
rZDHY2LYUrHdXRfsB9buqmk5fsZv5HIg/XFk203Hoi/pCxXjy9IHclpVY/X0U40vakdL4M9+INZa
6cITLyNEycbfMypb8ivlNZnZIrgxw5eLz2q/uMLioMyKCVh6Gi09Kl0akDzDbejdOeD5War7pa/h
B6nOJ8GxexWaEJcVzjBtLwUUVSC4Kc1D1NsYvnw0wtX5VDBHw3cO3dSkFJQutKr2+QvKOaM4Bht3
dA5TmC4+r/HQbXa1mAMGk55hM+xmV6AxszYh/nEe/J+yxjK5BjLoL+lnczQo4huMQI3ucKM6eQdk
ACDkNWpR5Lq4j7+nQZRt3rwzyBFW30Mb7qH1XtN67HCLQqAPcBn23Vw2B5eupLrYudZIIv7wBJcF
5iFXlD9sqRlQ/H/oMzpXmkpVegu4k+DazwcKYxQvzXUuS5wN/fiPYK2kdE/8Ph+5bOtswmgw9lwp
mMXZrgS0O8KmMmtfP7rIEExRQDTCtMvFL1rSlG0xAxdN9mUEPfaZKJ6aX080vx+8LPW4nT7Tbi1l
d7EB4bz0CfnV2QvWC8bYWLeN9XG9sXRM0htKT8vxeFKeS2t74fG2nJXqGClli5J150lVKTPfcBD9
tDdP1ta/QWYiu+VBT+jXFIQLvI7fk7NrAF9ylmwWgxpK4u1Pef8poZIevMTZ8vBtODDrdnn+XIVP
UsXR/YgG+fP90j5wLZh74r6qfts12jHyV+kI9YIZJavDMzHW/DhGMPST7mOgsvbZk2SLH/DFoVQT
Hcn0o4Wi2mKFl+uD10Ariarg2DnLIpByVMtJ5mlaV7A4zVl6V/Q0EBvWEhMn4ahw2Cdbvmw9ae8C
tlZ6KUxWnSCYqNOODahyomqkjLsuVQc9ApkBgvEmsxkfGllGeVB085eTodctniPiQJXuHBwVTAzd
vSa9otHucFobVXDaPMJGqZ9YdcHzyVMBd9XulJOpw5S2GCHPf5lZf/zxoPBkeviSCVqyKTc4Ulat
jFvSbsfhXfJHMy1fQvjvdxQROh1mbi5aEAkMD4/FwoxRYFxYyHd6KSQeQMsvSj8ScdN29uzNVVrQ
tFtz1wU4dslf99E82foKAccHkKaooc4wDSlLo7cPBu29nUushQoVC5wlN2ygF7pIXpx+7euhg/bj
XuyMpL1An95g1W2A0U7LwvC6OzWfQ6Aey3u7yHzaWmOUv39O2gbJoG5j+jal+tdCZvxaN7ii3Klx
k5ZD4AXaZC5mUhySW2JtZVamQLuAL4PsnJXQYJ+RFGMgXKgpEP2W6hbWEs8070eiI+WmDyuwdtnK
ROALNon/h3UgcKqs4abBG4EKqMmLuJmD1Wue4TGIVe+dTDEaOEsP4FdNilLfG3lRRZNcFr9iP1pC
Zt/Xflm3B4lYmat5DZt3GjPeh3hU+4UIQzZQfmMLS/+Hg+VGdVBzisLl40ljR1DMaiXxaJkxeh+w
ltf6KFVI8hGoD/9nc1T+22vn6CjvnB7F2CUiALIlM3OSAMLa2Ok68IRr5hetN3S3YA69G/D8TC+I
QjFuZwtoanHodXZA9LEA/lDkegXDa2DxDitKg9gL87H7dadwZ8lAzDD8bMcX1WGLP6QtGOZHlVkM
QWAWmqN9Lvn/WEHrc6aNKzOE8EkguJWQzrpcbh8xSlOtQSNhqtNx2pQITu5zup9ASW4mo9WSoP2N
JIrmK3/iu4d8CerN8M1HBUNcMQ/Xk9vdc+4IFs1vi0YYm0mOF05ZmOgh2fED0MnrJ6ygyiIFrdbi
DK4MBSIBhh0w/shCNCk8nhDNj2I42c9oaVKfWfONPfuQcEA8aGAVmErsOzYt0OP86l11Kt+THlmK
OiDIUQemxWr8+d5eIy2SGU5yjkOpWLctPwD+d28ZhpEfaTIUcZSES/7IMBhB4fpFfdCupMD6cLhw
CwKLhil1X1Sj4HCE2j+xoLuYJ+H6xxnlbaX4IXXZBcp2Nqb1TIjJuJrQqZtGQS3OK8MZd+CruAbV
8FbBq6KruUJvSWGXYR7PGYSLLPUoVAvjWawVji8LJc/jdmz5vRP5Cup4P7GFbOiNZXXZvZxW4TTa
QFvpU3PVvpZLVWwyWoe6LZC/vtvOoPaIB9ghP5m5AX0nTm/0bxU8USTzW8b5Pfsi76u96REA61da
olZuq/M331rMnOYc8uIhp/O6ZwEgS/dprmKN9gh4KLWJeRIBXvRPwf7euUzDn7R88KyTA/ZWA3ec
eYgqSCcfWYFQ1lO24B2C+hb06FrRSWGbZIzmlbjdiae1vOovwIcRO2epNbSFYBmnOaUfCBCsKpIU
geV+wyp2qtS93w8E3RY3DUO10NG172fB3BxFb0jTdqSjby2a+7GJ9wo/GnPTw0H7WoaWzgKixFr+
HSOIeB7qRNH3SJpv3jY+NBe46n+ygUsl34a9x0Pd8+nj9FTKV1uiP+1Xt1gau1/uXAO4lk05bFER
BKtXEJRZtJSb0sNtsvnBU5iBjIxXXizEh5Rq6F3Eg+XxDv+t0EWAKkluaa8J3868iAoMajj6nR0w
FCBH1oqH1h0VyJMbL9neWR0orra7Q3YfgcNw4nNQsdqQcP4fuR/9PjAxBe+/u68sibVA15SlrpA9
qF0hoKgh6qv3UFKAiUKoodIv9Ph5YZkepw8+zYCrlNOIz09uuGd0wuVmOscD3pEwq58WP9l5rw6Q
eQrEre9HGqAbBWU8SL3/jdmv2WOrZfLw/z5Nj8QtzGHWyoTXulEK8Gdkad9abIFnZZvuclZGNWAs
D/Hnw35cSVWvvJdaGW19NS3klKvOrEdjtPoJyVSbFwl4VfDcrIabmmWzOi/vv5e2fQxr+E5MW1ad
H9ZGfpMYAPVMj8qDV1exNUxWcCDmEhM3T4KuW+Eb0/LZSLgN9PH7caIJeY8uPmcZ/gxd3YZhyMys
KMqhyOp7cG2QO3fcKitxBoJSJGBkzy5H4jYHh2OlwMMTSsuRlPXQCInpBuCJaic7xZlafQqHcJTu
5Z5EtlijQWJ8GNnPEO0CG7LvEg1e2THmo4WrJZr7iIWaBc+d2S9sE5b0IDQMcW39b76CCQhybtBJ
7wg/CZh9/PW+AqVKczCbgEATMayib6a4jo3+KoTbum8hFve3p6TEubjh62IGtav/K9Ya/PFnzE/b
KmoiZQfkICcQISUlhM+ZbrdYxSFViigdJzo+Z38pH3LHNJNJpHtAFyWdu+jEz4DKwDcnTfHdNJiO
eLFYBh8/DwYeAFxHYiddwm2EnAsCJOnR+kagJX5jOMAVFmmyFgvRCtfU3GJeZVW7v6Z2VNDuYcTH
BM4LgO4myfv/ljsYyNE12Ge1A8v/BP/bFz1DrSGN1+R0G7mpnJSC3vpR8yhiDkhqlAmBgS1K1J0O
bdQW/eM1pLYhdEZ4DMwYlvb6YCvYFO4QWgktpJmXvHmB/koXg9fXdUthbsRZf8e9UAE4dEvDYS+1
C7GE5L3yS++2gae89nD/WJVd8gPIhEKqvB4CyuwhFcJUK84jYMUqW5yHimz0vPKwl3e3YP5lI81K
IU/C5OYAdeBsbNd7zK1/FnSilqkQgwzx80HZOiffZhnRD5Gq/h7fqlj7C7zCEoeglK/Mxdwb2j//
ctcbtd46Kotj22Yh8TCtAgvbUfXys0ZeCUYSrgKOXrNtv0vhpdMGA72QY2zmyWU9vNKi+7y2e2RU
zkwfY9TeZYkWOCYHy7qCBBUp86Bw83IziUKrGbx9Eevlesi0//2UoUf+O2zb79XBSUBkaWnkK6p1
98ft39HxxsTeyAeXJc6w/rrTYbA8gK/YV/kJMocUi4+V9ihR2i4GtaP6NdgdLMONJn+EC+MIYbWT
duRWPZHOg+CIHg23yYGFZXl+dl5wkfqNZQItOpR5udULfNiJmSl9O1qXfQ05GKl3c9h+7eeqSnJr
GM8x9r6/CXVeSrzDLf12hm9MZwujIHLsILu1aGvhofCrfLZ9C84546cipXz+pjF+UQGIlTda6t5h
sV0b4/auFLxi8gs7OcPLKHTszpIc4dhQMv28PuZYbdWOrDwMqebnO2ifGkpEVTKNTvm4D2uPrKgF
u8Ct3Mn64Tx8K8lKhd0pnbNUfywi6ibH+nJHOAEX/irdGMALRSnppKoYKJtQlKKVbTV17iGT9IGA
9frgD+WTrzemOQyht7n2mPsz5ShfCrNEV/Y2p7AVzMLdu+MweZS5Nt6AYK4LkDfikKTFimzSm4EB
pJuTkiQVBhsZlzHr4BIIAWBGSc38LRZPb7GDlzbBH0AsCP2fvCx0/oZ4P9LP0ezFbhDWtnSSXfpQ
QXn/X+g9Y3xsQ6Fjqg1CrjMCsZjUxVDshkE7Js39STJWJV3Ta5d5kx5/VBT5Xcq5Y0UeVTftkp+m
J5RqHiPSV8tHCaMe+8OyhD+f9HOAqoRFRN4HNcFS5qyx9jCXv1sc+6j9AaVIAMmkPEZgxzEam/Kt
DPMd4VCIhFKrV0akiSiJW5s21tSYXeWKSkz9ItDJn6Cgd5Hcs+nc7tQzA6seohkQwzuidreN8JPC
kmq8KWOJdD2wF3fUF4W6lbDKliWpucZyJLzj5Y2O+ZNCFlwlekUThUic0IRnoOQkcSCByEoHPnBN
Q02r6QPLy8g/LpHWnRAh//Sbt9kQ2KhhOQ1eCxWmG3lhXD69QVv6LvJNonIOTk7WRjbCusRc4dU7
nreu5G3PEjQAqRJJI7rBYYg7FUaV3iAY9ygpLqDZLeE5V9rV23kyokvaP0e+Z11lOxakArqI8yt5
UD6jSHuqmt0/3KYslcO1rtuduRKISO7ErY8nDwyCPAtK4swR1iTQ37aXT4kFq0KkCmC/UMQtt2R6
HwrVNTnTbVRo3eDOBJGMNpJXKKKGCpAwYR1kxEGUr8TkbRdyimj6Lv4zlprqyMZeSiRgD1/ZtHRm
NgQwEoRlNQpJ37yoMWSeeu9SwdmosT46QRaJKHywiGbq7KIpEU4Gg8dMEoHD2NKd5M459FyZIH8E
HvxA0cDbv+AVPeZG1+thCSMPpgZYdJSfx8kcIyrf/mX/tagqqIK3BwyhsxLqhYD1eN3cSaRxywDE
5xB2SoSTzOpU6kV9DdKxzP/bUx4iYKrAXTgYx2ko1dT4gvZklnwlrll08gekDaNdornKOPx3MIl+
T4ZV1hZqJEzIbVAvckG9pqQxuKbRuGhQgnH+OvSuYSXMC4VkOc34ssCQ+Aod0oXwlcbQXuufBENm
Hr+yO0teiQeXKlyerNEmUxW7IaY4DkLO1NRI52RCpl0RlqwxsgquS+ECqZokTM8v6GU9VoYZ/cbc
uA+1SuyoAbRzOGnGlOxn3Xqg94/C9fsP4Gv3Ih1aw6F9oMugfMWBH6Cj1Q8WqTkjOQij92Ff1O53
XFwjyleB0TlE+pZZlg1FbNvHed1B282/mUnDe+l7PMaTLbb0HuiaWIEVzD5/865UJqk8W2DDoklx
9XFDIrFg5sBiyb4DwoSTP/bcYUXA3mng7Ga5pVfQt+0J8hORLbcMwCUJfJD/Eihqah2r8j+mEinY
jej5eMdZnDMUFNnE0V0Wx3o5kJdTIW1eQb58EFglC+qPXMlBdNaN+9lu3cXWiQdEJqn7eQBQmcwC
1Zno7Y9YSRrFO3+T7p+DxV1DIGjGPkVvrsAN1qo9q2ntaO1hhjuyC32me3MeL+LbzEY16Hau0+0r
XcL1FgqYZHRz0bxiNlijb6XpVcSKdoYBHxne8MGa5CTarrYTO6nlekmzPPQZZdN9cD4iGmT+b78f
Abht7r1zSCFRE22z6EiO4bt0y2rOszmYMTMVXXyYYotqyYvzrzv0tTsZMDzxW62azsb053ygNflw
3xjFPQRHXEGizKZsmo3VnKa0pIBmNWuz1dQp46Cky8T3/WweVTQ5qJtz7NOYuYoqWb1ibTNk27A7
J3a4gFyn8oC4DGxWutczS2lNKEvJlHQPqovWFGU6EDolCikqDNLFKvVyRrdemL5xvuZFFG7PbqzF
P+uUrn1uKDn9Z8hvZaNtqQCsZfYJFFskZ0qrslYkdF/gNTvRjb9VSstsy6neQoqG+6CDgjnbu2Q9
dEi8qQTxpmwVW+FErhzaMcvqrUM4GeCGC0c5HaZKYvGVeBUXb6zcniLS+U2fSLacAY8tGaMq3FLu
AZdEgMT1IPTZ1WakmSa0fIahfRme8xqD0m5SMjLQCXG76x5k13FYMjUx8EfKUW6UY29+6I//O/eR
PTfSX3nCTw0qFo572jrehLg6tUloiITY55oJ7WXWO0iFqTrvKy45RkGtX1ktXpKWExzPMKQTu4jC
e5qh38j5rBOS/meHfC0+iQdaMWwAe7gikj3e/qEuv6Meu9OQzEKtRUF0drfz6Iz7IH6WbPfijb73
3XZGf8zfyJoZMtagQCsbzCGD7R5gKRElnQqm1RXXoFPpgzl50HMXaOC98hdawFdUzMsQKm1JvOPF
zcWCFmHsoCQcE26IqMbiD5mEyaFKU7yKb5ZCMXgJ9RwetSqFCXzkYdff3rCrn4Z9Q939q4uM4s5l
rfilOnizWRGQdtKnvHzy706ZJpMh1L51zqTdcrn9uU67UijL+usJulabdYMWoBMGwPH0SnJRsgF4
x+KGzwsdIeVfE8YhnNnyv+lh4DPxdU6N8i+iQIzym+82diIenroRVUp+2i1fyBJunUZTAFmOmQNV
w4ygW2BuStM4Bdm4wOS7KuA+nWe/83uqrN6Mc01eZ7VDF1+IPdD+0Qq7DFtkJZ9XDbrY65dqJbtS
mlz8Vd23vguA1hlDG9vDKIr7hkealSs2gLXQwZiw+wXeJlMztXVGMz63jvQnvWZ9zo+2lYQtw/q4
bKsdOYiiE8PhNLwl/TBrlrc0yaHFVMOz5NgX3J48p/6Bc6UMfvtbW316uRDDNNsDay5ratHhGQxW
4BzCWBROfcWQ//eCtllTTVbWgTLcVMa65qn6fwCV7Bt0PV+yQ2ysoCdIat5LBChZOkoqGTdsI8KL
zNClhe1SoPLs1J1141HsxPc++d53pYJ1j/EG/QNQJSiwTSkFiR/WIzBAzFA20rFbRf20HJZaKXyR
zBUwNo7iknYvRIt/vnRYcsL+kNaq2WcuaiOiKBqdrs2aqWgaCggJCCX7JYxNOtE+xZpaBFYWtPRI
Ea7ThZjAcBBxcLUzbAZgYiXHXIHvRA3V9sXVWA5zyFnufojtZEe5+R53N56rTnVQYBu61yFHloOj
R/HzNJD+wvIJKIPu6iz7M42t7rxZoH0MhojPk4E1EQkpd2mlfO8CzNjBXexAtRyjnq4OAC+Sxmpp
6hnmAOAbpnpE/96GOoVvedPVRK9PjHVsKNK09XiipcmHm8tfGzrg/AX668eJQcsxaICasOy0lSjl
c3Zv1Vx3g0BtfRpqR9DwlCl9tpkGe9W0rJvR/bkfyQWs6XNR9mnYM7aoPavXr0pNOHEzx+ngBZJu
t8r67tAnvyewuvD/q9LVoFoSUFeBaQRJP7wN9oAA1gftFC5j0vAE+KozUgFN4B04H/mjqfKIXbVb
dBtxeqrH6GcvLddPOn60rAjgZw1NSbBHaNzHbOXCE/xN1y54OO9XjF1XY+tznbhALSleDYG6Urmq
rX73Orhq1wcYyDyNpN7uydDJ1p6p44TkhCwMPEdX6vdLoNG6uVprCGLJtqxttZpVByhPx29cXwqc
Wm83Y+pQqIAS4uOCEBjevwji2ZMyDhc5FNH2wf1ztrqVK0fAvtE12OV7JfcUvQOxirFlhImhWC3z
tuZCgsvt2quL0bxnI00qvZKwXzV/nbJptfes+LqrLst7B8WxYd4Nz3lZ9+vA8pxA4p0yXFEj9oGZ
V3TWu5PLMY7rlB83UBj0GzZLYZNpuS55YvNeCEfMpY90raeEpNvPvBjoxAx0GWcN9ijhAB+u/jAu
fNAehcb6eN6TPreRNPZxs8NGzoUyQHrad0uUlSYyLWUCcrmzqE4UnpvYpGwJsalPCwLfJdf2D2O7
gz2xF9mJ8IxUOBY2JvVDo0kukMZCK140OHETt7VCxRFV9Q4z0Q3tZy5lfI63zm5eAhluU5bXUAB6
oM4opfWG/c5Svd1s3+ZMuqgUVAiTtJWbEKsprZRMyk3nNo/2hpCb83+VRAZjyh+Agy6hr5nhnXWv
J/IbpHenHHKy5skGjHcQT8crYF6K40/JHxy1PaqiRyRlmiSbkThXjNKuXKjo1xhRvZzOe4pjikbv
/1U8gf6BB7C9yPvktJQVdXhW8uX6ZXGy5HFxXgKfM26f6vXAXHp3vhpypC89FheV+OKg18ehiTTT
w+Np7vBLxXb2qAIloBlulMdnawKQi6xo+Jbar7qZYW5PKRmP2tTb5p+T1DwwoPb/yLfUDiETARIz
C2NI5Wo8lf9gek1YhRLD1I0O8gxnUdK88Ec8eR9I/HGyr6269pZP2LeTxHH1qcXMYkxB6NUGPMgY
V1E5x1fcx7IA7G6qRcYAqohPj/PkMtQjsVPtS905VuKQiz3uQka8weDDTapup1etQxvSRSaud2qA
L0uSFFVXeTDJ2mW9EW/GDs6OHjpV9gQqjmC7Et/uHtcQsZfY2yXO1qlHM/I6sXIac2r3qECBG66b
DG6+5iiojUo/uGgpy4kV9ZDiWWRhCa/PUjsbscIk2E2W0BaGLVq1/4hf3k6vuCu60m5IJpMsLWF3
dqEQ7b+z0dLVPrsyrnK3INkeETPSFdQw2MVpKi9m+6kghFPemL77YrxbJDVcEsWfPKlMc3P8Ows1
qGp7LA7088w+G2lgyrJQxRiGFY8fhm2lXBUBuIH4LoXkBU0PcEc8eyDtVBTow52UFtFsQpBK43PE
eiLHvaw6BHhDOpupSomPprzLrW8xuuOB5Rwd2x6KDS08AvsfdCER6pQW8gF9kdb/p7BSWfcQRpOt
gYM4OjDPuu2R2Z6WGQ5YLuMfOEcA4BFKKAp35m54uP2cPmTaUM//4namoHqr8lvdhx/boJ0ouz6+
OEp3gUTI4fRvd93uFRnStDuWM8eJQ430o1O6sTG4k5KWyDnolCfJg7Zf1eJuEC7ZYaUw61pXLeRf
w9K8DfTtgERRMofKBrGzQAzw+sh1ehSAjL5t8t3CmPL1jM6ioiHTFA1ISC76h8kJnlw/IwO98uJ2
wvA8Jz4ViBKQO8/iGJ0fNeS9xE7x64gmeiVvwd6lXyhfGK+N8Q2uk90uPK3K2Cg3RIh1ilh30/o4
BVWQxonTrjGA2rjOXQdCcrU1rJQqOPL90JKpKB0Cv4xFnV6iBvBIT9VYq25iqQm+ey2h9tIUYmg9
aJV4XeXQbQ9Y8PvZ5TL+y9AUrPJy1m9swld19VuFFqnWs8D8UkR/ejEQaGsgpV3+QSOdD5fmf63e
AA/Pp5uEMPKrYXGtU7MhxZsaZ1AW66ngCHE/gBw78UUhMcJM8L0ZgsITGUa5ui4eUlDk4SOZD09o
b6iaIRNlXLXEcuvXKdKuYTY44uPyziPOS8O+u6+iNtzGZIgcxQ86DgsspWiCNNsU3DCueBOKjRE2
JN68rUvzLjZNwj8GDUut+VYvh3ysB1IiNP6jebD+Ah0aTYc/5MD/hSi1qmBsj5Bd1zynQiqWJ/xV
n6ye4RAeQTWQXaIrCPvZkWHrGHYB+PIWCCTG9E5SFgiWHMzMAihiAwCxZqgRksJ2Jf2Aa2omoGi2
62R4xVjWAazG14h4NSm/9bMdWnvcRNgKXK2SW4gEz0dB1yLKW5m4pFQg1w67vjUsugBAwHjMMso5
XC8Pcx3lLJp8W6/C9Kpii9+/Crp0sn0BykNQXoDAImg7MZnDfnG50yAsgmUDVxZNruNg791aoIl6
0nefQEVFVxDV0QJaYHCigkHHxGJaBV3B36m0boBIHFs7US8bpfusdS14IbWrw62YFQz4n2RaNy2v
+0e1pomwzd5/LYcGVusBzgpd7tCcXIF71q+erR26CeoO8tU2Ja071TptVAUttmWqNBGy2gOAkj04
0gPA2Rq7SCscN5Hwg1J4DU76UA3eOqiYGEydTOM9PSD+YqS9qkZL69oulIlMtVY/rU3vjAHLmN0d
nE5s0KovTUBnkXOs54B9wunvvvEjDnS7UGUJG1i1nxstKI9vZnF/K20g/4uXKPc19MGXSBZZqwkz
WecbDzB3d3kefvH6Sdzy8wEnydj0jgye6VkKap+gHjjhNlu/IVeCmH29Hpsw9SdTA1jl7hlNWZ91
qGwRmInayKZZb44f4J5TRVf5jagiDrtra6Kf3/ogJlkOe5F/U7PlVK/KHG1jRlDNrg51ifoipvFV
V+lJCX/kZjb/S+uSsgmBWXe+TSb60wqcMw21j9Uzh1s1br2hOKRbzrpv6oZGU30QudKKHOJ2Kgf1
FOmFMPYXnTorzES5PhE+WNyFGlfZI7XcTONVxgmphkGbYp2YrglOh6edIQIUreWSQ+7T4Ahp6WJY
0SLNwPNVgHy7FaBn4C8CnTnf8fezT5xZmJMP9i9MiwgigR4o52CjEEngj8bsyIVCa0pqwCrZdzuS
pgxAmRyrfxvxhPtBGugaHZ9+Cgyd+3O7uiwczjwmSDqxxa3L3NxOo6niwzvKmTmy9TWOCbUmpCrJ
wW87uIfw9Hwqn69M3kHdvVLM8n0kl/JkAf8WvDZHdhNXYfRzAe/5GRUs3wYYYHVxk+iMeW/JVAGz
hPTKMQuxcxedKKrZy642UqPb6G7oqwdQlYhEhoCoxNhubX4nH4hJTjcDUHyrSOFgCTqwuE+TfdCd
fuBLXsVZzu0PqKyncwJhmzBnZ7ZQxkpWyPF5p4Gir7v3HU08ZiXd8WtmVFj3Gp3qjzVilfuvU6v9
ipgeJkhU2g/mqL6DiTj7aU5bT9GyZMQttW03Tq2X0dk8Vi0ZSe+LBL9dIFn+0b+erHHbAIl4eJPI
qOpCTjd01heEXY63+f0nRFd0PME3eF7wdaNIjA3dqet9qh6e2c3SMek/w5o3NFS01ylrc7VSSmKw
y4PvLKiKVn5E6QoBXjzgr7ADBXMY/Thmtf9k/3svlHeR+ONrz4RKG16VqQBc+zibqmCG7OrVsy+l
8Dd67pOK75KHEhnXbzJvGtU1BvWZYfvkiXhWcvNYvrK2KARA10daZjf0ESGIaXQdv8chXyZ5Fv6n
nKl5RQh57Wj7dpTmi7hHIcjgIfD9C+f9XQEU5gn4fdulbxUiPSeFXH9TY+VtnIiexIkvnHdZ9UFC
o7QABmVvexcHEvmVRbXkqY2TpTO1dZ4BvgOwjmZjWeJotYyi/N/YKcc7K//BbjmVW0HM3v+NezaY
V0aRDs9fHj/jKssuYrG5Kdqbm1ZZUe8JqrOHyqmhELH3Mhe/USkuvpOpx8nRHP9qbkzkgKZvSBwz
TJuHhEe8Ui/kJdVyTD64K3VWNWDW0+qC0YQNsBlpnnrEmct2XK/m1K6v5Ouw17zh5KlZ2+7N9+HL
kmZnerayXEwOE9TOa6u4EBr1wfoE+dGf3oEguv61PKA/UKvXPQnXBz9tz+gohBsrba/Se652yV9M
sHznEjdJDZcIQUU5rbzpY4xKCQEiFKb5+0oxFMObXt98HY7GfL4km+EIx28rELghgjPWPknW0eAr
b70y0werLUt07oqKB7C7AUQ3n/J/pZKTgrftVL60B9YR6mODMUdSUiBGl9d2qgJOi6iXlQIvfNjy
fKQpd3kpUidDvRD09+n3vvKIqFwhtK77tYQ6naq7k7BXgczKMUMp6GX5ka7aZzKgaB5m6VlUWYUn
NyR0RFbSpGx+2eiB5tx2uTf3n9hPt2nuPXmdigxjNzTBV0t+2qC0Z+Z4q6v1iT3t5beK4RM4Jejq
K4yRJEKqB09lhLzQP0Uphf3liMe+bjnQjjWnT4vXfdUvdna0dYSUpBpSa+921f0V59LMzQWON6qL
RahVPYWm6d4R68XI1xO8HqoX+wJPeMj7lRDAY+wQw9iQE2A/zF0/PpLM4GlhvFXOYxFPcRmReoll
wRncNqTzldvPoYpMWm3Fz3lVYghBFsarFpXNOPTUeKdSZiz/Br8rb6e2tdolw3om9uWNw6hv2EMk
xJEZRXFEYv9PPkr64TSTHTzskjxnrOYd5iL0Trd3J/Dsj7PFifC1E7gwP2SQ6cALd7GdkQdu6XOv
Iq8/0ZpumDJ2KZqANXILrpG1qlFgBuL1MI1UaRnc4LMMGt6IXvmoauFeDFU5JFnUXZsvK5oeGe02
4RulNGlNS35oXr9DkqL6ZEP9Wg8cw7qkejlwNTHM7n6ns7PEGF+UbVP//21L5QRoSlz2F3UgCXaz
vGBNpFcthu7e3oqqnrNVQeIdNsfam8z4xOT6UujQT7y86JF9GJnbnPBJSKhGaccI34svjbXrBGgE
WrgGU38Hy3D3y/ZsPZwQ7toFSnw7VwW1DiGMC7MCPAiBI7ZZGJOpegB39Xz8m8PtN0dKv8x2zlDT
Zdd5CJOtf77ZDoEwlbswMFAWHPIUT84Kwf0gyk/JoxS1Y/BODJMAGU0Lxrm40qIVDtG7AEdj2m/J
vuH4cGAnmUu5fpXNTSOY0O7JtHs/AZmj3SV4KDZflaqDW2qlE/WpvdwJzjtcud2dzmxjPBJFAcX5
HnO5iDtaN2Ep5GYSIe/YB5LXDZnQvfVGoe+3sj5pc2jQr0TwEjyef+KhoyPLqmHSbIvojfygzaye
5qF1GPlEnaCLa0SlxS79hBtcnxyG1PvTfGsLIMj/nvSVJAskXgML7SuJfZ1LvrvVNr7H4+JojAAv
JK3ezNjwca0RG/BAhc1TQsRD4ypo43FqFBpkt5BwYVQTGbjuFbJOuMwTKckRLLSPbpsSDBV4BKuN
3AfGHJ+hNhWcZerJjg0QxceoW9E3cBTiH6EgGqltjudW7fkjBkrGZ1YBYFH9KqqxcBLz9zEdajmN
DK1vqP4bA/wsbKyus0j8q8e/fOs0aTmVvwGhOoYjXhyjJRN25/KthT4w+dmOTB2OL0iinm7S+V73
Zg10xA7VDAPcv/whZ21qFsYLyDNR3kQ0lJVkOmaY0jtkipAAYgWOd1MTmEBomSMwR1a7IiE61TjF
JmVrDQfVPEf/zpntxq+QypY0Wyp10J3Q0079oH0OLY9SOpBEKZzlOc94W00hUKfjxOjGWYXu/UXz
j4h+KtUs0h1TqI6423+cacMTR0trOjg5u/hVTbWa8nDDuZzuQGS15DSMFe6JWKCk73f6dc+QGUV7
Btu1wtVYU9WAY74mOQjGE4HQby4uY7p5fphr50QG2F4jHZvufQ/PXUJii16dqF6/N+wM6+udemec
4/b6Jc9vokMeLW4dH+vjX8AW5j794ntF415WQztRbkPvXmiYxQMnYBKuWUQU62DT4Hudv1MBka0B
HLl1rc45pkyKVIGsLChRVA3erlPY44BEzGwEEPneu4PmJ5qfgqxYCD+uD2tUlTOHuOcYVKyCG/um
JMLXeY5hekXOaOkIVPTzfapVqM54KhKiQpP8ZyILVzOHXJfbRUJlyYBCL5B5Gqbtp++4ahxbLvAl
6/rzqEObDOqcNfLsUeYL5pZQvWxdjjmAKEzU6LvJilZkOACQ/xBLeQhc58W9CG6ZcW8Asxdmxx5P
91F9uhFlVAh9nx2/KbFvSiPTOLPf5igP3nfXTr1B2xjavQpQCxNME2G1ZTlXD+J61+HfbP1aTq2u
Vx7juL1SGgSBuc4i0udrOSXQR2RBO7/uEVSWklcj3yZuWc2+/yMBest4HJJPC/kjZuoqh31BSoOu
aAGGUm7V7uwDd+qqAPoVqBWb8WQuZLNrGJZpV5yTrG80AH86nnkenrQjC6ALPoXXAbCs4Poh17JO
Crk6gJjwT8ibvUptnkKhdU2X8LbK1GsgEXLo6CGPgv2huYK0c/JIHliSv7VCtRbLNdROEhSktg7+
oAzezdsMddww5jg3UcoYtu6PoH80YyBi4WpwXhM1eVHMqNh80+mjKpP4V02W6ILqaCFCAkR0gVq2
InbeSpj4+iV5tswsD1nXQq0Sj809r2jhYh1j1vtWlUpueE5tgNa+zv28p95zQDLJCCOOpnRh8VUd
ZvF7DggJ7d9R4lBs/t16icVAnvMyiC9Kl+qwjrvyc+vGZJjfN4ZzfCG6aVbjH27rni47qtga4GeX
dytpUsXBjSp1cKPZmhlSaCewpaAjb34lYvbOt0H0yCLwcnymD/26TH3WIAZFRZcN4MqAmn954EQd
PvPES2S+6Lqa9gDkLVPgUQrT09HmAQhK/iJnhuhyaidSUA08SwbKucH5ry+oAjjISPMSh1qZmwfX
+dHKS4vyZoudYY9L1xgyjilyaNMO4nMhDabVjZbsZR9AUbBz5gwIGsO5rbVPMYc3TT4i4cjsHCP2
xYS0rMwjwLdjLHAMfuG8cPfXAZm9Blrce3ZlvsGT6ARWwZzoG+F/3hoYFQPX8buZvK2lDxi3xGjh
JVkBUJRGuk1RfLu9bS8VdwQvPUEJAQmrPAXiPWKMjCybeo3rW+ihNpfM1jjR+EhwC4/CJttraGOy
FlAdaoU/bA5tNRbsCUhKpiN2Yjr3LaEpC+mEMjETiLG3j+oLVhk5+p+zBPantArWDVczwHQszoV2
fG0aDCFvt2KEag7VKS9jQFrtrON2X6cbrN1djToEqcKRrGqELwhdUG+FScuHz2Y2/v8ZmvkHeNF4
Nm7ely8bI8JxloTDM9w9+MkiMRKbmTv81aR83De6eSw/p0yw1bN75337Lo03N7VKLbRFZNi11YQ4
sP7eGb6l5zcRQRiV3zMDMZ87203+sy0ZAOz8EiRAx8W8mrqJEiAbEnnVeOfew0SAH1qDyC3FZ307
/TC72jBoNoxmDMkeqGwKvQT11S7xJtBF9NV8tdYWgq7RKKscdeUl59GDJ9VMEHjKMrLWgiC3w0QX
xLbY/kuGr8FMjSPVI2wnsOUOlJ+2WUJnKOzS19J7Hb2X9ZqLTuOx8iwyr9M0wx+7hYsGZBIu4PLR
A8czzRvgCJZg4hANIzZNtgcV+3zG2tgNRWS2NZ4SVJ5HH7Yb2qhUU+l6JnD54GNL+qm3hXPk1kgN
X5s9dKNaV6gEzfIweqMGPo+MyGkJXLX5j8TDEGx+75rqSy0u5BZPlMmxAh25y1ucBWKLboyjYnI3
0a3iACAt21w1635I3NbCSYPjds5Lhmeq8rpgM421+wgwXfwGoj3XWAYxGwSWhFFQxKeodgHtfWpH
/3dit7RVHxyzysLr4E3StqC/htDibto3H9Aoy1ySYEpaLcWzIM1kxVq9c6PAL+NmS7FbYySsjcuH
9MaJBqYakC+q/lD227Y1YNZCzJenb9pvNuTenFojkHI4yrjlPpunaCc7zHjJPpwAKj1LMxVDbcm3
sMh/5aEn0u3MLdqNriH2AdhHHDeWiIRWxFQRERN/B/fH616C1YzUHlRQwwuoQcmygfOMCsGmvjTk
Qz3jcIeSeNecp6cxXay3E2DR7M/GsSDnQU+VevIlmtTvm+6EJZnElkGOy0FVN5nNRfx3bCI3HzxX
N5lwnLw24X4YC/4hLkYeSjxBZG0//eNP/surZ0AQOWvvldllFbAJ8wF6tfYkhk5y8vnQKUjszTRd
zJJCYhC/S68brr58qYnZ4Fgo8ngyefvqahX2ntMGV1ANG0cowOTprAjKeJtzmzlmGHJJK/ChpNxI
c9JI1YUVK+nPgYe/zI2wpOEwL+y3Vj/dNBXdRfxyD6LoRrhn9iPQ5U5C/JcNj21cF7wKzgrSEv+v
eNuBg+ki6Xe4R2XIcUvKphLq8nVlmbbbAHRwNTvBw9a1phE7+3KHAPqDLim+8VMmEeUBev4RURGj
Z8XscE7Sp5DVgU2OhSPWpYgywm06oyG7T10DseSkpSRZO6BUWMw7iA2z9jYEXj8M07BHKd7pbQBc
H9g9rKoCc+7R+POkaBbzMe0veTyMngmDXyZ53MxLcPWNAeNJbCzN2+tSDMK2WagtIILkAeVBjBuU
zQnCaCS32aYOpIpSUgS7ysH6y+zNLvf3VLTkluwopbtEQo9u2JMo17Y8deuDr+BVjqQdmt9pZLzk
2xba1GaL7Pq5aByiVBGzLqinSmcjcyaVf2/L0Rpvr2Op8xRdyJiNXGIeq4OMIgBaptD3SG9yi1hP
pXISzCz0kfxsC+zWw9Xzr0TxKqrxA1VAdGqmJ//Mk+XfvOre2iLkJ+0mrFjVxCvLJnK90UJSnTWt
doYv6Wubp4KLYofy13gjuyXPVL5yqoFZVivhQm+McY9PSFyLvk3qg/tzSe791eyJqInInU4t8TNx
i3oQk8ZKsR/hd1abKVfZGG+fxoM0ziOEVkamXSz+O+9CI/kTrK8c4IsDXN/ZYE4h9cS5vT7/LA3f
YNZ6aacMPlAyFJX7lzLThMFBCw7nmcrGyG02haJPdLijdQ47QCUBfjlxrFRyPeiQwnemYNRqaGvG
VI74UA4kjYsl3hrN54oN07EdXu8wXj3nejIXtYgYymHUKP04060GKwiXJIGrrVySMyv6ToCsWxdt
EtZPZqcDhNamUapnkHxBPOCagZKSYpg8JPaMD0V4hrLRBUPp8fkuQ0XynTXCATeUsUlJ4A8sOl6e
Shaf2Wjojh+h69oH9biyyr0g7/cKI0SGp4VwgqIpSX41F6/M8BtpVKV4sYbBEN5QK1ghYehlj29e
E8/y8RYj+tdi0BBTVPmuBUlqgyWXY6n5xlQ6hilNF1dtsMog1RcNDbph5rnDPa91tUHp97+q+ZyI
myHiKWYQ/T07GftRkaoxuTmqeBW3dsDxPK1g7ktPq055q9KujnU3Y77Gz8sGH8rugurhdNiVwkgy
uEqzS/JrofVa1u53amBoiNjCkG74XCPwYnqii7qFP4ECorYtp4tFkcM7r9ba3+18Z4yA24gqFoKz
xpMizjeWhL0cojxiNMl5jZDLDq6QRiGG+XizoKyIE5RecQeHAJyqbyzy9WS7SnHXhvp5WD+m7tkG
9lyOIpmm3s/f3sh5ih6/DIfMIJQHNYwVGRbZWtIXqVmcBKk5cecr+LJcs+gzO6+eTBtKxOYSGkwk
gUbT8NoGcs/AeXRI9k6qYQVtHpuVsTL39BQAay8hcJBJs6PsQEMfnDW+485BkoNUNSXK/AT7N+3a
HPM74zJKs+34J2a2nVzxw5vl9O2XRFA+3BtzQRqzIAwpv8wcXoyyEAxt5Ld1cbmm6DrNZW8hUuqT
cojYy9hdBCLaRJSq9bwcGgopEgEXA3z7PJV5CD4NsQ0dMNXSD+SC5/7LKhSSch7C3m0YC+Gq1Dpp
a8sMQc9CHLc0EIuojNAhUAtvxdeIaWkuv5V1f96Wa8wwv57h+jIcRbnuDY8fB7WL2uuinYG03mLA
PWe7TZGxBBubjxVaORINDwEJo99sSK/kpV44LH8jjuwXiZ42xvkanscj0y7SqGVAoBiO4TTOCyYd
rIdnLXuOY1APo0fDYdfozsAtCcy5MvKPZmv2cwq1G67t5dDYjRdl40X2Pjvmq9uGHTxbaLQ8rtDg
gptyXeTrKGuK+ks6RK9oeR3XwkRAyp1iAilLaE2Z2WbjHFrwpuWeHN5hPk33NQrD3r8YDTpLLSWY
SUAbIIO1nPYaiFSeIxmFYe7FKzTJs9ycHZanM9g8sGuTH8NvWs5wRymVeTHiuWyLFOFGCar3lmxD
ZRMUWLXe+dZqu6eAzObthp6wzFtOiF1+xmsfVBGhjp4sA0s4c1k6O3EaPKwEnMQXkMIO71znOn7d
0AnlJ6ORoLv7LlW9RmLnqLgBBY9TQaRErz8HmOhNjFdxRs3sXWNX49D9P38z2dZFyca9F9Xdleo+
lzgPDPlJW5kqtkLPeTw2LnfvetjpAwjbkrV1+WRlslIStAPPDx9cjQBDW0uesY3ZjxShqoWiV/7q
2TEp63RVu0LT8s/XH6pBSBwsizkhT+SjOwsfJu992KLbRj3469vEdYXBwrsTowwlDmc9rJzLD8Is
5HW4mdHx3eV9Qu0lsvB2BMBZb/udE9E+VZP9SvQKgvnKHQNgstzwmkGZkrdym9L6+unoIZIoOoFI
+UYhUB7eDT+wmBjBrEc/kV5ngoAg7hBsTjZSXX7aXeLDJf997f4vT/DVBna0eawsdhAbVEEuid7v
sAnx+Hy5cya7h/BFiQQzifK44x8jIvaRaWkBGN8Zl63XC8NdAg8PUnm+ujQk0EtUlozhSjsq4kZz
cUF8wcFZG/7pkMKYTXUBvbuE5JQHcuk1y3XlpDKwhlIm7eKcKWcXjbpTHWN/gJSyXm0Ek3cAUkzK
d7G+ECbgxtOU9jQzxU/8iOf34PLWonIrZ+62AdLZL/IZX6/6xLpX8nyWqK4oPOOTetJxUFKhf+na
J91r4RybmkVVWtt/Lz3dPDSPk94aEKOkBgQv61vWDhZ/c1FPlGQSuYxXl7Izw7X7YJWbLeMxmkDQ
y29tPvGNAohgBcX3FMjReRsfjNmkjXMOobr0LAO5Pdizjhhm4ute8f3mpZYdwCRO2R4O6G7t+SVt
Q0beip35EGTddJCI1x+Viu0e0B5R5LxTPHKnhO63mpiXzCxLDvmuNsWcDccEcOax7fWRrAV1Byt4
ViDLqLrjC1uCfzd5y5te6E3tJMZggQrDu4YEECT6A+FiMAnvIBLcAjlukuggsrKBdUWzv6sLLPNq
qlYm/XuaBbHd9waG6eJnfOkKYKyM+AQzx28S26vE7L3+vfx4qpYHqAzbvfzXfvYu514wj+UwIsj2
e+mlJgNn+gNNR+5Zv+NWeMTSL3fhlAaH+hSsvMHZDO+VMPKVJ2MfHiNnC181ymMYR4CLeBuOitJV
2C45pATxCsxlSoKPO8AdasLsYhNSsoyQI5CU2Gt9mBMThmVLCBwe5i3nqHJdAgi4tQEwDXwB778R
Njfq9y5FwxN0PDcGwzgcIqeakq0NBcNr2xrazjuuFz3AmbMUIaXlWm0k4DiiMc/Pl8M4Vrvvy+2i
DYzvD4OBthYAM5xckqvyDByIsVzQxKgjrHo4igJEWa8L/CYwSeaSsgnik/9oEiy1Axx5V2H903PU
Gs5joJ+6VNvhhkfYLnUeyIMiep/YEf7NsPcZkcLe8QhHckvZpcV+WvWFV7IK565I/yhTZW3QL9cn
FbYSTTBmEQOUbyGSOCMmmMFh74fC0P00yK0LhojjZKHom0Z+2yEX4EaKryB3mxdAv9k2aFkHSUKM
amfieKGoffH0602ZL5tC5WVo0dw46eAbuNnTglA/VXS5nAX6ByPOYbQ/AMXZiQLxrOBwAnFm/udX
xx+uOkHvv6cJXP4kB/AQlejgPowKJGJBvSlh3wSTQ261BWHaTCSWNYDU8gMhivq6daeBdeeNP1i8
XeAiQE/jd+ain9kT3tgJIpi/TW6ZnAaHZGdB868vgBPhOchSWnwbZKfZQqT7YEcVj+GMOZMKE4Vm
638DUrM4vjuEE51RKKR4x0wt6rBKZc0zecmb/TsqXlBKQFPc7i2eOE+9N6dhTIgFRgtC6Flx7Wdt
0Z5jxqkhq5GdawXni1DukbX5hjLMRe+ztGRnhUReon+x43f8wlegOMAH0SLhyUkJVGRqmGiZXIsq
DVw37/guegbhjugZJD0r4YOcsSAs5M6tFyN3cuagaqRmpLZgENK7oBQzbgCl+7i1t7bp0aLh8ySP
7pZMrOtG13aNp1b4bLFpKIsI1WZ7qLAiB6L47MPIkmgHO/VXWrKRQH/zeTQmac9VuAsPvHPF3qIG
G9bqZ+x5WOOP7L38ealgcq/7jdPBQmaiGmokO5dFiBorKjGyJ0minAsNfnnY9BkKOOxTvVDXf3hE
RKJigYZ/8zXyJaBWG2LcdsSLDXLc0sEGlygIv0iv7qLlHKu3d5Hr/aWnM4SSB+ti5UWlac3apT0x
6gJ57AC/fE9e5ffzIk930iQc3PsU3CCVychmazDM1f55EIVBwopwgS8NV36MKPVMqB/24V13aO9O
p17O+LMRS33bxWFUo/O/yrFbfBsOylOqj73rJLCGnoE9PQFzIbJT6RHA+E+7ctjQgFepIc1bvZe+
klG0W49x4sfgkVvowu1gDROpisYqp0kaqsHZr6Xip/iAdzsBoY96duNFqcAy1AhDEKA7rIZQ1z7n
9ynJMPwzuLT2SsZx4hBrtp5OJMkxx7V0vB1TZa5II+4TR22U85yacCXufk/JvLTRtRcvgS0rrlk1
jQcBlMJOlUT1BD0Gx2S3FBq6OO86oXyX7Bl+2iPWwkDQFpnXPy6yTrXQ+ZstXyFvUrjJJE8qom7P
RB5CZHUny52OAxpu8wbEYZgTYbl67MS1AdVH5n65ZNcgDja8me1LITXcId2VXvftgxA4f/629gHU
De7T77+fsI6Tamy/SdilwTT69n5akl19xN2hsN1ebZlgsEvBpMHL9VN5OYxeiYSAHScyR+oaIoQ4
WRrfW8Pqjx6kiMfOf/bG+Dxfq+8HfI6Syt6w9zPd+JoiSBctLgC7d8hQrfxnnyTia6vI0159HtlU
jKOz1wuNV401lJUce+yNDPsrjBkMsAoqhfrani0I1Ljx+c/TxZMR6v/sLiye4DQ7lSqOlGeZFWSS
Kpbt/ILLMhMRUQQUmJ449M7v69anmbYAMABH9zF3GoSn/XRq6i0JmZ12QUC6OFglZ0GK+CkuWX6z
eFQHJSrJvdfhuItN5VHtbSsmAQnjXA8HS+we6lqxTmn1gw9oqSNLYFmjBIfK5H6CfQYoD/J/oGur
KYg3rY2ZHOv1lSv4+jhU6ZUodV33yUewZYr9TJiM0mGfV/hjb0A8BocVJNFnqvA2mZ9fFFsxVVuG
g07/giYXj3YHf4LiAoCGWnZaE66Y5CMXQLZgpw/izcHmOzCJ1RWu9MbEKvHroGelNfySgrYQ1yvL
mhJtoWJDNS/he7w04HkI7Jf3yk66FCyvynsnehQl++QJHXgUCFeYujsZip9par+aO4WjxIn0uXRi
jX/0lrNKPkumfBA253S22BeVXslOsKVtHIRWXtQTFwuehWC0VmPbHBcSIG9bvm9IF37Fjf9KwGPj
g5Fw5T39HrPOHdu4n5jFNGsG2w2sv0s8WCW85meKWznmg/Xtp+8i4iZGZDKaXjxj8F17nHi6ucQH
X8xBtr1+PgMR5Ot86ZHKzB6BTfmnnJQptjSKyvHj9u/5CdJNqri0zPuCZpxidS01sH7cu32lA3v3
a4medXCOgvSn66sbvorEaxWds4Mcot/GenFcfW2DbLYqP36iK6fVJSRdAgtDHQYylPqOWR+7Fbn8
Jf2E/mQV3SiP8dThvoQiObunKDecUp0NEL5YYBZaaX8gRiBK4GHVU6Nvq1tLbOHHC0uVv9zcXxKI
aB+7fY2dQgujI5J30wRDhsIBUBtP13IQjpihcXhQalPGiax+WGyoCaEqUBan3ZojFloP1snwYe0X
zs9x4CCPIyko9Ius1P3Rvl28LjikAdjqknTzUTDSGdDpe9SlWbAaobGGm1ji9H+rdnaG7/BXrpSh
shr6faovOIz9DVQb3NwD3NJKazhDMfC1QkJnKuBXKWL3wMNv3plD0rO+8sniIVn7qtfYWsT3zDLf
DxcIYsr5xutwRtnHBnY1X8fiLYL11+b16teUImEZ96/hBK7XB2EAstAFl3qVrq+byZuNLmUP184m
bi5UHZlcZSb/8uajMnge55iy8YZ7Cx9rsisgXtwquHWr78f+YXyhE1rz5D+Oq/XhchrgPnLctIP4
tjHeAFo4mrlajqnjnApWNaRUjfJMutBMwKUmtcAjTNi9fXa8W6sRUf1a808v+7mohr9pgsaVMaTY
J6HclEnChzNKLFzx9Mw1/LcgIRPVYhhs3E3dZ8Ky+WbyONmenpaXQ4NagNAQKATJ/D9gRKyjHtea
BchP7veHPbf5Z7Z7eLgoX21OOT7L2rvrF6FZEGFlRP83ctSoc6eiUgswCofNNCAysVkzlf16Hj+c
J5oZl4B0NW4lr5g0fc7XnJV3C1+dzZcEdzfOB2HObuofdS/v3vxBjA8P9CRmx2De9EQOj80otxSq
LkUhLTt5MMvV9wiW1t1+mHW3eRFz7HD8X3AZnkdTAeJGOB8ZhbJT8eH+bwp6BUioyebWMvg2Shhd
x3gUJt5hrGutU1zzeIi9qQ2Z4p7UYu/sDBTsp/xwoBclFI4ooARSwnKr5aKP7MgRloluTLxTvYVr
4qdf9fyCUYqp7VqBo75KvGKoxRLoSY4bgpA2K/pyRilmihopKXBplhucQj1E8ra3IcoeM1D1OHTN
O+ipHHeoh6zK1hFKQDmFct/t2hpNTBXjLJkuCiXcR3INkow2XK/7HePZ1xvbv2ldBoG0pndLGd9K
CUZf1iiVcRsSdglG6VY1SeAwLY6WwkURSy0uIOE0T4NHVNb6SAcvbZtdg7qeb0g3sh+jjamEUnRh
qkAsCWmnPJMNPXpkYfndCKZsmNWwRSsbCWCTYB4Hj0L+3h/P8mKpgE4yy75KGUS9HdKNuGKkkeUY
Q4VgMmtICfVksJ6cHuRHJyrxVKemOKKgfRMyIc9tVn/AkW5bpLDhj2tkTdz+aQwA2h8B46NtWlIm
+KCEaSKcspvwyBMEMhAcIGYrAJpaBPZWy9nmYmix3GNZKn+oAm8vzKlCh4FViFmQYpQyXtaAcGMB
qpx42/hOlx0oJ+7Uwz9wswUike6I2hYTWKJyzh8zqzb76xoEgMQYRpK7if7iKUZON8faqKY2AuDS
G57LJc7KzH7J6a2uLnX9nWbeCOBrjmwVn0fcHQLR99TQ2Yr6GM8hyFbPYHZljrAKh0el7HK79yI0
jYZOfeqxbbOMXMK7X1f0WwsZAslqrw3N/VssFpOGV40m9MhTPqepu6WB6Za9Q24EUmmYzXnYHO3O
RiJOCGlZ0QZDDLQxFuGPQiQ+oR6nB85ZQi0Ehj1cfYqRFY1HNQK370XLTZi9JKv22+lmycTIBEW3
0SG9SdWyEGRKo81z3qyvnz8hF+A/YjpUREfR0AWwffG9XeDvcCz9qWNZJodsh10N3uZ+D+h1zwiC
C/xqOwR/8LLqQ/JP36Ex78g8p8wqsCbIloi3WWwLma8x0ovfVmDPfcvH10bim5sgQCG1siqi+/lx
ALNO4+AOABx/i9boQWn1H7n6BiURQ/QrAkLy4G3+Zja6xSm1t7jeISUAeVn1Kxwsbgbp5A2/LRjz
Gbo5xcuQXD4gR/WQen1Ww26NT2Pu9qj2Zut+AyBJwSELfbBe2NE0jYtnHk03WHe1cB9Y78dbH65Z
RB+9r9lu4nyOnKVbGp8x7TNyn/FY8bUvLsLL3k7iQXkJCZw/0WvvHWgDjqnI/bTYemmrE6DLep/4
zxtpvh4zcuU2iFJbYk8B/hoiaCkAaIhtUJf38nLtglma0E6g796p3VioCdXyKjKFcGToLm1dJhAB
siYQg3Swzw82ooX3/yi4eftRQKG7piRJnsQ5y7b7hwwWgtFriqNyyX94Najeoff1kbdj34Yqzsp2
wNziWxEMU7ClX5nlpQdVshqnspZXC8EsJXVvmYRYT9p/59tAH5x0jS5ke3wujCBpyzLiQgHwlh9d
G/Fgoq2zYU0HL8biCiRx20TaQgn4ZYY+bVWT0Q5fe9IzU5lFnkSKpJ5GkM/eqr4DUDb3Rxd/wvSJ
tICjIUK1wMpNjXrV6zREneHY6+ALimLc0O+pzwmcjAORB7cQzMjUwlquxBbV/W0wW9C1bHepWib+
Y5ej9H/ZuJeIlH652mD6QSEk2j0h6QZu3glaitY7RB0TOnxLjkF4uTFSKAB5YhKPF4n26wvtqBci
PE+PeV3V0hcRWYI/C6Y10A7JBR30vX/R2N1/3PMp6BUZALtbj0yK6pmqDYkIJvaA3Pax3oVWyP2Y
yWwyw3BSQvAHSdr4xJzrR6Rb2Z2hzGXVsIVcCYtgjcz4eaHso2T8KcAiasy130xLvlXvwybq8rci
M0vjMv4bzxI/hMcTZQpcHUe+J7BauL1jOtLCTjv6JV9UNlSaeb9wTxZ6Sh5pERPpCEmlXpIl1q1s
9esUYKyfM7FS839qOY4Y4eXG9HpzPqSGotWuryDORwdkwXWPtidLL3e2ICN3FsSWfyCFQLkiV4Ya
OGslzhiTA2TCmZcM0NUWrNoggqtPZT04nMePOqsdH9SHx5Gs7/g8NbqD8Sp5x8myVStjRAmCRKB8
6KvQkCkHwHqVSkz7l/e/Nv56KJLIyuMBt6u0w4Mz5M9Ze46DlHh5m9I3QwaEj3eyb9yG/x9HE2M/
xGOQ36DD3ljY7FWj876+A/Uor9EdC8WXispae8E3gbQUs9c5Us7eGMy+a9sSxcWZtzmfpSDxEtka
/jUHQfRGqUZX4TVb8cnJrfjdKEaaMnMDdohET4/HCWGs0bQiyQrE99l5RX3CzG+YUosKjFt3is2x
er8GClnWdVjDKp83nPlSzayIS3It8EKkvLaZlHEw1UkqOyxHb0tmU7KSKK3d69zyBsAMMIHrl0jC
QqoYCFxQ1k5hlnZsEd6g5OFMsWoaqxXixDFO4juZp2nICP4Uh3N/q0d70bPXQQ/gVQhlSb2Ge39Y
q/MV4T//UxH7CynXMQVJIicczKFHtgzSot8/9FdzfSOHS+B7oGEjgt+iHGd5wzrWyPRfYrF3SiO5
E1lbbISV0jUFERJvKh5+lqECs4JXBb8OPuwx9s5rJ/zXSWOgIM8MBwztYJ3v4wM0LbcKKvqw8J9F
VxSDlEwhPoEo0rrqgowXaaP7ykLTMM4b7SLhfnBRC+v8j7OsZHVx7FEM7qmx1/b8Ti4Jg+ayCn94
wGgiMrgIvgJCOgsVShAn1sshuvuFU4y7Gp/qnOJkBUoTlhTKzlZPNpyBAbdOWfIirm9N+aVTahXt
59SJ0YDhTQi7fni8SzK4iN6K3FeYuiyuL3/nn6WmRCzrJoQblNLPb3nPmTXgTp0/Y4ixZ3BMCFKP
gLSl+CvTZ4KoEDifzZIgJLf0YIavWvMKAisraAhjG08Pk7OGL7byKrcsILQEYhYWmAiIE0ZDQn0X
mwtRfa5IWB/rSv6Jhg3le0CLtb8Li2O21CTi/dpJmOsxRahJo5k5mn6fa6l3O1fqgmdp3epOc8jQ
qBHzezPwsvZW/glcsU+RFsvW5420crbIOsHH/UQOmDL4MiYrIslSZtHqt6rpV6HCXTAPOQ0J0RG4
UQePM19k8pyQ4OoZKbSd8rmugTfLDVtq/E/Fh85fmHPxxJpdl35SntZKUJ9BM2QH2f4yy1ZGo2+Q
X6vIW6SHh42O86Wfx1SXDKbuujgbIp4OmpxtXemPUsWSer/mg1uuSlCT8MgwTjjDiK3dtM6EQlcw
SPUQRsHSRy9O49L0o/ffQ9uyCAL0elNN64TE6CHElcbW3dmsVWQ7b7U73ZDCiQ+/OJLjmboYxant
mRO1Ygtn9BL059nYAPRVzNLkviMkfqI11FzKLTUMT9SBGsMukl3kGEMIXe8i6YwM4jMKjK4nF3Eb
ObA317N3vFQdAdX7Q9tRdkyeEVhLVRt3r4L0bvCFrbEaJWFB5CbQGrj7J5eo09Z4Hr5ZO/BILzFc
r8dHsZ5rBdZoZ8hHbcQiSXV6shRqg/LlBlKNO5uuQLYBNeJkSbebx3CvHOzk0zsDV1vVU3963Qg2
OsKdCkRlJLW1K90CAbaLgk8WZ35E+UqXDczNUsLdVynYJ94mlVBVQaQFn8ahH+0Bpl3Hu9BGPZDF
khFFhTh4VylRn1RAxYRHMnIqifRbp40ozhZjzq+2qTeCIjB/U+1BQCR75BxpyLj4BOHj77EVbNPY
zqJrpwUC8tFUgC/mS8Arff8K8tReSkLIXBi5iOs3ezn07K2hACkG06Xpsc0WdlyUK8lzMDPutV2X
uXk3cwtr5xzHN+twgbnzUFkkH7pv+2IA3C3X3oHtT5gULW5Nbz6BmbkN83yfHh5Hvz50ByYDesTy
0m51UQVY8BXj6hN1Mymrw2jHDk5SYgUvGspjb8RZIaPXGpvPG1Gb1lT3Ya7bKXUJuTnS8ypu4a7N
vP+lUgXDrTkDLtmpSERaL4w9om1hl1DOaZx03FKMXVDNUfh4emva9G6+HKG/LMLH2YCHPyafcJAQ
iGNT0YBofvfYrD6c9l76pk77/506L4CPUDbZelpWE0Mg4zlqGzIt7fjXYlAecUYtEkNFjTLIODFT
qj8GKI7IDQcrEro2NQuSnuct77Fz7atQvFIrUp8KCbSm4s4E6QBX1WO0ZwBNEZ8rnt+LUZVdM7ln
Xp1vEqiUznmRAgko5GXMRxUPDJ/dQmaWab0h3lavv50nBQZRKBC5S6Hmj71NTK5JKl2BI5FRoXCG
mwBGIrJ/TgRAwulmLMK6StooTuYZMDAwMtxCCF74hvjvI6O2WiOSC9o1obSZeJtgrNjgcjRIlDDT
ovRIquWlOYP2BpCDNBeu17TF4bRsMJNWsZezQPJ5vUEXlW4jWzpiWV4uBfhB5ZwbqFF7Te6044T5
CPSAlJr1jz1hxlSjZ5SdHUy7GQ5f5NJI2UDk3LJYShVaO4/ns85O9KXABx3uRoLDCOg9Gd48IlKC
joocYi2KAdthN7nfJun6q0GtC5wNNMO0XPJgjeO4pvbn2HWVDUscObX4XPmFSe0X0nfG+/zqgWor
yOw0cQj9RYWlZTNWYYWbE0mW3vchur7TI7kJHw5sGqXWgqLfnZ2wPWMoxRCM0Ocjvb0qs3O6wyni
DhPQmZCYBhYScU2hL3MEb4+8ma9CH8Pye5M7eIM1nQZcZQfRoHNYsOHo/PfOi7dPs9Ptydyy3pnr
DG2tY7LjVCihkVpk0P7CkhvidjnfoOOiyYApdwfhKdMaj/uf/4tQ/CklSSRtUbrdIIUFTce10tFT
S78WK+iFUif+p8+PX4c0xHnlRC54G7tR5uBVfUwIT8pvaqzaylHJ7o9v5273Z7EPISUuv7X2ldBe
gUnkt6GPuWabcCAjJWb/T5wzSlY3c0MIpZWa0zQJYzWRQyaZDZoXs22YUyFZmdX50rb1MwFNEBa8
rKX/PRrXBwceJJZmpEuSj6zSNLyZm1EHP0Smv+9L+KBUqsdQjDlSzb5ahNwtBtEfxqhHrinhG3WH
tUF17SmjILAoZlnXDlOAop02xOKn/gXg2xYQVDGvqqiL602k4f77TuId5RH/UFfEevbegKN2nQuj
DeHeiR0ftFO765ztWOCyTxtiYAolK59qBw+CJlBJhE9SYPiH3brvcG1dDOdlk6+TNAvXxZIEpVqU
LHxH+hbxESgIh4sDFH/pDkVhSmYAUyVFp3zzDCeWv4cX0R1o0fN1fflBXya9ydW6zIRyg3PXSRH8
7j1+uFcnlRb8Ka5zxkgIZdasqHwXqitsem3T1+3Au5YiFT3qBNu3uYpPxcMVDNw3O/JYIPHDPiiE
d+AnSO/kSF3AgGr5ujYuOrgDTsZQLoP8JsSDzNdvWSZnePcGvJJnEik2QGrb6XiGgbKJW0sHlFxd
4c+WE/y82J31hv9q26mms8xtyZGTxO71K+bHpzFdYJYk88ATH/sUjwaL6n8HUafTV+p+d+WCFx9B
iYio4Z2mfPbAgceHHaxQSBOLQ3fjLN5ULcYUrt9srxyFI+uCeTwO1ZXWVRq1/eLKhabt9Ej9mCBx
ULNfwcfZ7zdwiXa7jmvJow/uWxZzNckQXaScUSFqgxBoZBFiQ2AWajmX8ZmxaeBLWkhyprveAIx5
zB4B/QSi3SAKsLSjukL834NT48ixWhSv6KnNEGymRZKJDxt1Phb9e2YjuxH3++ipS4033qDqhwkk
jUP6x0Zz75Svc1h26w9F1jPLGlCYXnxMTgdGt8ser2UZZRHw74nYUH+8H1UZJCatNdRVnhKZt2Gv
cJyP8LUWbvmuotuB6kYPu2GsyHjfqf0kYL7I36h3HRgLxCSKGXAvtiGUgzxKTGB5a5eFemSxMAu2
j8AyGSQp+AER+yDYfHoqFr4bribWaCSM7/LNphdsl5hBcZk1yxM0zhVWjGEpy8zZMfPBk64KYaM2
UWXDJcwmF1WGeDW51x0B/Wt3AP4lHiemwvAqcpeJlft5W0xrE9sRf1Sr5tMOgkatfJWNGlgN02zK
2PXJv03n0kpnTgbxuRdKPBkI491x/LTHIyivuzyR7c8E4agDfLnkGO64cLgthwrcg1opI6+GopcH
k7RJ6rH88N4FH8IHgCSHGJZ6OtxrxhwawBQayTWiUgx9y1lKr9rZENaB6S0OoJBiEyw+uwYA0jSg
or9rZ2HBFJomOjgRTlg62LHW8wuf2krkko8/JWPitZ+SepAlfh8j0HBQ7kcU6TkkEnwk1ba5D/id
akrE4rCC7zswF3+Td8yzRrXZiB5IIvU3x5rli2gE3TJkGifsYgqZcDPyUKSOtVNOma32o765ZE1B
Vdxc5KPvjUdsApdYlujwVjBRBlghW4dsMBgEQlNU1bgrWWS5TZVu0SMaOcEvBE/muw+z122qu8sb
6TekErkAZyBM9MaCX2qUeOLBTP2cgVoz7Xh3E8ScTavobB4/9xbhmvuSCrDUrCKxWTcyGvACsIRx
XH9Puxb+fznzQR8NM0LPLw4ZFk90BU69id8UQY7CgY4r1bk6htZnqW8eBZu4Fv8fkj5cZ1VJchSk
P+RGyf2W59/WBdyqlcdt01fiYb/IgSDbBQhsvUE4p/rQc310cIQngxW5335EyTwlf2mYHsiwFjib
BnKHSPrAqOMGfCHDQdOAiRaQqIm/5sJztojxGIFJq+UoazQfevbdVmMmFA86UaOZ2bCEJptvy8gV
WwZmfNpH5co2BgNrA7nRM7Dacz/zPDrmjcpuIQrPCLmrnX/zWSG1mqpTl4aAmW2msdzWqBeZXjYl
OyFQnwYXyyutP7kB62A1Q6lZQT1+cZ4DllrxSQ5iC/lC101lroLUjoHvxiKfSitYDUg+z1gN6A87
0mORMeC7P/yIcqBWVStY96IyEEiwTPn9GsN7boNnVYElP0wQq6ByZ2YzWpPVRr/kqJJhRnGQ5VAR
qZnFK95xhCsTaasELs8/ha7+1rz77kKalJLPqDcrBW3l1t411cYhUouTC8A0bhoHt/suyrKViO+D
oz6LFIvI6xCfCEszGAPbRrC3SS4iuIiKnhi44GDkO2AO85PAI6ysFZedcWyjRaqhHZ29jNPHbIYV
XFzNCCgqwdTbOsYzdbNdQ7OYAh4rMXaAOhuyeSrBo9GNfxUJE5qLwFfnLpTv+nIvOTSx43fiXGOZ
Vcbvc0ZxNoxwhOuebw2pDRRa/F40UevJKXU6CvOIxUuUT20MYYxX3+8XNf/sTCDW6IR1NtiDxXPd
SQ7bOf1/o5AxH/lwHx4UlADDYqOijRkKJLIw3CSfb43LyeFSlLO/hvicsGbz9CRcPSKGDZVbSv/k
QKtuAYcBXv8d1AHXjbsCVkgUo5LstgUqNRXqY4kc1Kc58T+vZpQX48zMcY8BIkamJdcRm3ZsB+IZ
8d6PtejhVAzx3ozZayRAbV9FrvEHy655/C04/ui4pNa0GizODQ/3kIuXR8nxCIasPxbH0uTJuCh3
/dC1InTg5TNFr6kSQAI6VYn0hwB0vkkTueQ3XYieviTbvVnOgGwsJN/e9u2JsCrU0ctYu4RW2/Yb
gBCAzEBbqxVIA1kiTY4rUslUqp6mG/t/EE4LFRueLf+GRy8XQYWSPJ7XHlX3C7p8E4CBuAE9v7Xq
nhRSkVk63OHT15mJNUjBRp3UkFN9HbD1MDwmT3qJ4KK5d4WjVv1I4ISWFhRoThk1N16lYit8IYDR
JrLNrIQv9WoVMqBA7NGXgW66Ab8ll49jucy3OMpf8vqF8pv/1EYI68MbPi8/kzF7MzAm50YhpTmo
z0/A7ADgafpi68oUo+Zud+K20VnO6t6ttBn4E7FHJwTJv5vstcEowhYkvKeTW6qFrpScg6aoAKif
jwErzHLiWWiQ9GXT6ViTSTfWnNwf3CrO6Z/GDR8kr6+AyOY3uc6X1rc9XnHwD3P06Klzlu41gHaA
uOOfidiZ/5d4E5EAuF+uo7enwrqA4alSBFmr9fA/X3ke9fs/bppn0jP9QDFV30Dn9c5JTbxmqHTD
mzRju0iZLJ1UZkdMn5jRZ4WebgS98cJGl8koYR8JAgpqg4PJedz3yxJo/Gis3h5P8VasEVGyFhN2
/YXCp4EXYxDXq21T2Ce5z8ZYPUaejK4kNpE3/XYwkeYB5f4lhBFKef65VDtetTJzy9e0wypPDXHP
7Y6Y3kndFkbeQh+6K+5m72D559i+1eohwnCaWHDe+j/oNOYmX613VPo8eoEvqhGvbRVy6LyMDXS1
PeQvTrkwzNH2hsewr+qHaagbU+vILsnSS6LiKQqYTBpZBC1s6dS64BQiV/fifYETGEZKLdd7YhgZ
l8279BI6wPtVYBjhS4zp5sy4Xe7r3iPVEGe/SW18fnOioh8CVPtss6QD8nowc3qQ23cIIrgpFjRU
Lg9Uwk9qtlRT19K/BWUR0SMLGf2Rvv7pYBqtUuK/K2evlUeUop5CSiAimV7Yi1OJvL2po8jtArEv
50tsV7UJIFU4rsnZabicj1slrE7aA7MXieO+lDe5HdD1/9TXYx0rH9G6juReFag4tbXv6gzbD1Ek
9TQMTnUkT4zK8asfWYRbSd8HS3Extzhb4Qk3GNR8QWkGi/rTaBzfGONCLtGcL/YkJi12HSR+xdpD
hwNRUSNf+FbSOi532uq5uO1gJzVxLS9WTNzPQ1QwOhBE+AN2+ovdGjq8mzkSRL73hIoMhOiCgobK
PYCKBCglA91fgSZxpkJCIcg12Es8NRWaUlP3pPpYdH3GzqERSaVBYfA95EZ5sY6qYeLzHOw3T/QF
8HykW57CeOQKxgDFQ8tt3Hp4vp8qXHDzx7R4Hp8picoEO8dWdWzX0p1tQV6zdeqTJzgmvuEfdWfv
7M7RWTEHs6qZ3c0+buLDXDZEgc8+FlPpms7sbtebEJOe1Bhmudd8xLuvlhNwlsDdgF3VtwemZnVl
KCO8ywgQAQ3g+9Qr5ozXWIKOdcMq5bL7dg7XpeeTgSo4D4LerU0bP2ZGomkkQQY2krUoscwwav6I
OnbEcluQQ1XBY8uEL8Tw5Ge6fAmAYhAYQbo3i0mJGV/wbAkjSA7EGteOxwUS8juMWzUPHJO9wDiH
HvOsSCImEf2fBE6QZpG4x1Lx2pJxk5fRBxordwZfv1gOHHlIXQKaBJrmhQ/zMmXueq228R6U8bG2
xkD5+IIsq2zttdD5UggBNHwv+vBmpzc7yQPlsTNdOhv8zv8Mm/dBGpAamBOHFogQUGe1t7GeMETB
lgDPJ1Qpwfsno8CS0VtUGF9SZtxMnRFjImfgeTXvyXnMJ4noF4ii2Rr+Ypzbci2brl8bwAoEwzzw
xwFjs/G8VpbT0XeX27vKVcQ4A9C4/p5bOORkJbWRlu61YkwiIx0ZtsiA97qD5DxS9X9StYG9wSrq
hIfXweF27V7PzhfRfM2NfsoRrLaw3Utk1S2Mw2QNWA1RP4iR8FndQtlf1V2vPl8CHbMKSKf03yM9
fKgcTWCtQZ9ZLFLyEbdSiTbqQpPRF64HCa1uerHc3U0FY6PhL2uEANeoAfg3TeU0TqCGb1lO7gZM
o5KFS9+KcJFK1hBX1nTGQ+eejP4Q6ADf6YSYPTlmtCMq0nnNzuqiCMPuzEYGk4KicRe4aJWybjVv
ecezHUrXoSMs1WnE0FPHztSCAiCBDmXtsFoZPE55OtTHNdc754VyaRnFihsPY1sPD9g792SbabV5
4IO4CZXrIGVBia4R9Z9BI8lKu7bFSwNHgOB5IIObeO0YnQuHObymbizHxxxM9BlIB54V/d/sHmR0
fdDv4DASz7tPSOZDnt7RojgRtti9h4oMBBtQQvJ/XU9WsieeG+QuaP+JJ/ZOgfNPPmIkm1wQoPKh
7Mi0QLyxGd2dB7Ruk4ZjiVB04LvX2ASL77qldnuZN+EqOhYWpFkcmBFbSIIh7jopoQvjBvvwyCl3
yD9UT2cDqBFbZXSUztEFXvDJbNeZyt7Mkavr9Gv0EC6EKyld0+zj+a6IIqSKj0op4MyROwpwpI7U
Pifk9HTTgaVH7+i4i7S0lNBSzoTbzOXGi0Ylq00NfQOQpkKDxnVKMYbyQIVQf0gIX8NnBxipXghD
RpltmeXFqwoT469vMakkZJxgi7MZhZy5oAXx/vq2lbDUwmBoECYTPZFO5yCcUsRZapzjaBbdq66I
CE2lSeJ9uC+OBCXn6gruhv2mAjiwhpKpR+TmCd1sqE0gLFiYvzZodP0WGmxFjlIAyNfX/EfCz1Oz
YvdWudIsIJsI2r4Nqchn4uUio+LCRJ5F32K1o+zl1vUezR7tsA38ifNq754iOYIcB0XvUt74OUIt
vDgJ5YZPxMb0soIlWJwe6ZdwNjfKxlkU/KNOmExGl5MPsWRSBWS2mwrTtdinMQWeLvQcuOEdlBb/
Kqyf2X0SSJ/wnciZTvScnzBi7qR2VTNqLmxFdW63fJtKTThv34bf75HlVBbkts47IB0B/iEVIHYR
gb0fA99i0A7gmblc/Zl3ghD50g+hLThVE9GhyRAEqJdGHIKUYoFTj+ZsWtUCzKBr8IKG6w0zbEql
zfonLH9Qglez7BL4cMUPmXBiJ9uy8fDgQ9HrYN67dkAGORoARaWIZksRM1S/AjLhx3oUzDWhBkbH
ZgI7zvNzQ8zOtI2nMx0HGgqHZk/23N10+vL61iJsi37+mF/s1QOYGwIdi1oTRVKXWkKQVxB2Oixu
d/f/BuoKAbLl1TTrhNoBxz249pcVCRosVCcpFNW7S+lEMJhzHRxFZeovE9eUD9TmfElnrOgbVneb
kFC87hUVQ0M3pBVghGTLpb24XLm9HGZRazwuhY3aPwsNCKUK4jQKI4hXG4ShV34CLWJNZlpmSQRe
WwZ1C/XHDMg5/6n1FIyIckXnvP163VOrfm74udhCpBwEVnJ8pRwr7QEpSv6dXPcO7IRVUxoBBOda
jsDTDLcPRQHmCgNATINTOvG87b2ZmTZULbaGB5m4OY6KkKUB36CYehpA16OCQ5HJW1v76isDHqj6
k9HNlN8Xtf/K6+VhryfyBwjfgBckeQt0FtNGqnjJGL3CMJwBGDbEKyJd/Cruy+JlkfTo1s9fz0HP
m63ttE1pbEuzXXOB/VyUkMTdkRQCIrKjxNgfcagqXS07xCJt3nnV4Bj/mUSxHnJdRdXKLSJoLevJ
NZzzjdTrm+Cx1WNjgKt6Q0gn/eXGqH4w4kPr7MnKwGIshs/g+YZAplhU3sCyrdYKVnA9oT0a/8jI
6dvo1jNSYZY2oZGOGbccZ4GpClmIKMcYVKE0pDXutrkRsU0DtZun9TJfOpKw3lt7tdyreejWviCi
J3oiCiyIWpdAbKMgRygrahTANcJP8EGahp20WCTE3h2OMJMEYtEvvwf8BmbOhzWzYNYHZiRGm/z8
7xYkI/n54z1rpHA6of26PAaMn8ej8YFsNRK/SzESIrRSBokC8zhY2U12o6ADqIz67KYKNXbOONDL
xcqWgOHN4f/lMM1sj+myaCAOWNnLPRpm2La8xq9VbKsYTPd2fSVKKreiQLZySy56Ov6EsXsbFzTY
VDHsigQIVujU2detpq1/A73plGG2SSaVmrIoeaI5eePL0NklezIpnv+4ibgJY5hhTaGagGnhH9eR
RjYSgClkkm9X2xzGUYXBYg13c1hJSbyuN804zZ1NiZ1eYijIvHi/bhs22zTr0sgEZg1QcZmngkLd
ZtsopK2JqdXmARdMPrqpAjUPXBLfIEyXXnLQqEP8X53UP2dTPFCGo6EFt/wn/QuF1uFekl2gTSkq
U6i5Pt5lvVK1jipXw44tWoaK1HQlwxjaT/RdmfHDlBkOmJLgObTj+qDni/Cz1SoqfC64QsVETaII
AS1i+pvKaGqB0o7Hb2B2ZXMJBd9bvKgiv8NdtrmZG7axZEazUGPjMJkKEoAKfehpp2Bu8T9thKkC
6U+CaHTpzq17onIvv2NpCQ+cMm4ddN+1l0FBadUijeNkQCS2NUkHx2kAwrNw46q22Lu7EOiTMA6I
mb5o8vtlF6RYdWOOyqI2iZ/AT+E65qW5El2ea0p517SKBuqSbEwWKB8YnkC1hDV2yo/Po8QzqxY7
rkLQt6pVkC2aXySGk9XPk6jZokirJIum9KRJwUTqrG7xvJyNwhbQ7CO19HlOXdscCAhdqEZNNdL5
wN3COXqaxZE7IZ7FeJNVDCNvHHHbUhq82O7KZg4DxeaBU6n9ltUasVNDwts/KkF7w4cz+eelS/61
0QEkL3I4HYNlj00zyMkzOtMraad0xjMF8zlqe3SIDIsh1JGCbUm953Em3HUOyubjRip3VOYp1Xmq
JvADQZuIhkGPgyXvuMf7/g66EndMTkbl09zKGy7n08JTt6gih+kDKCdK1HwcATiVkPdr6QM1+tON
9VC+5qxe8xIeo9IEToB99odpOTwxkxKh6es4lbOhv28kokfWxo6HotcorNx/8psIbYny36uAVg+b
ZRCs/HERT6kFeaFBzy5boeumGfRSDr45G/RNNl2xjwAL0Y97YQLSwl4/n5sLuFf5vqE69lqqsozg
zYbSp+g5y8EqsDXevQPUxWuEy5xyzoo9+/Hyh5YrNxMH7B9y5Nk3+QCRUq7EefahoxqWdYPo/fjs
7+4pLMgNHx1LIWquaEFfXptwTxcx+ESG9YxZDLCIppMNcQzjC2N3kGZFG/2VHCS1wDGmW5/wB7Ia
xj2QrMElLcYeeunTI/7WZEG0OFjkKXyi4xej0N9QdkPa7uzrc2BTwKcVBmXQ8En7C+vNR2wna0kp
8wF0sd8F+AGlUo/oh4diaXBIk9tok68E1AEEUaDbk8rGilSQXrw/NGHvRc5S+DXxn/JgSvFfeaYU
rkLJo2oJp2NQvfOOJZC7O07ldFcWth83c4nm0DWgYygJ86tWCkJHwHn5UWy+XEawWzSH7V0s4Jyu
2VBZc4k71CVBK+hJ4VB3FhC+o8zPcmV7xGsCrv1Op4m/5z21pCh0FoS4YzynscvFQo73jADXDqmY
a7kJ588SSAR7Avq+F4Ef/Qz7u/4v5zJ5I+tjtYIayjC0fiBKS5yLD+iZWgTY5fdJng9YV4qOw+xG
1t9WaCNFRsR3vRT9O332pUD2NWRmT9Xvz7haKQQWWjHgDxCQwQVTyvOJI8YwHL13pV2DKZJbc3Nq
xSbU/JVbmAaK9Y+O8aouV+N20UOug/gAVNQJk+bdz06vXTJigcew7mKIRRt/AkEETLXXr4/jyniZ
ACzB+r27cZAOjTSDaiAm8A4UYQBX6XcbNSv7GoeuyV3+skWwLQxV5Sx5nNj3UwO3oRDX+MvKSEUD
rh6CB373F59j0KBmQAM0qWRcHgEyy6si1lgjcAGvWbMu5luuJAD0sTgwogW3OUdjnl4qGe78blYD
ybii2roYU1tIT0qbaZd+iQL1C7IoVgL4KyGuY3EsJTUfFSgMJ8Ta25GJp+FegtmUmcs8NF6RoQLh
+6uzu1m/QniGWnFI10cYs+tHgtLaPIxLuiPQVdLcCK0acdFAuIsacxDFD0hhIV3zmy9obLp13neB
5P++4Cxay0v+0wSzCuZP1JRZw/w+uD+Oa22NtbNlht9CDiFizuvEQSQifF3gjBb0kRvgCaaz8Po2
lPAQ/nd/eMiwWpvYoHsX/TbBruleaa5U8WWqT6CKF3cJLWMlz0VcW7Qc1LJaO8z+9uYQUzZCZvEU
7jZiAdMX80R826ad2pTeRbGRZ8tRn2VDS7ibP92IF2o7gry7waUFno29+J6r021UAUyDRr7OtA/l
sbHJvyMg7KD0p6a7PVRbmPwFX0INnjkWjOLyRLXbwN+RVTpos4lXBvBFeFLL87XSYVSefY8tBsKN
1u+BydI+g5gud3fSgrYIvsBiH3l5Tze9c5GAfDzX57qQKTMF/tU5iSUZy7Rd3mIsGjq90vSOZ4lr
LDX75gs8tTP5afvRM0tIIbNk/59efTYnI8jV6wraMh3B+PTkqag53Vu1nu61YNYSiJfHca2mHXZK
fiHFeI0jOFcTnU5D2Yof2XXfRd8i/1qFMoLMfyZDX3q9wkQvxVOkNv3oC0g6LLj8bBvKw4pXCEU1
dDD3KrU2ikTuz+uaP+wNGnlOrNUeQzyRjZTC2+7oIZImrtBumPY++xijWTGUm3x1iRNUMb4XfdlR
8Di1POVZDY/FApOFuS9TKoG0mTynYdYRsKKqBqYkyVeBghFBAJao42AfwYPR2g/4Er/hQyiMOJ9a
3BDmfPuvJE+Y50EqLXKMYgSk//s92XsGTrpaPQM6GoPAC4R9AYv1ii/NqbovPkveRjBE7m6T0kdQ
xDCP5BgZfUe7Ez9H2cfyWcC7lNA1AhW2gvBHb3NHhggzTvU5sUXa7odjpknE9rYgnIOTx8oPvIly
KmV2tZvbjeGwL9RvHHsERy8jxcgzuMlt1s43dchhfrVzXh04PsLvPm4OmhKVdZImxfJeXM1c2CsL
DqMwVyTAa3JtUXu/N+1RCmyivKIE6iHr8pwExbjauFNzrdN5mbSxBG5qbCLmXwhz3vQQWbz+buHV
bf/URBuDceremRtzXjpFyXgvOeCFAr9Fjabf4bEqnDCamdEWpJ/lMig7lQqo5uo/3NhUFeft0/OY
GLCJrarLb+C7eFCZe9zYdEnqSaTURk/exGwXvnSmuYrFpRCZzik/ZFxWDqx/YCaFJ5cmoaylcdGF
efedX5DJwTnZjslRS7DoWPfalw/mjHAZ50mBXzcuxDtO0+w3fEVyr/1+f0Mszt/wOiyPk8DIqQUN
3twKfrKOoPS9Af0spQaDxLhpjwvkhSVZuLVUWN+BvoV6kPXko+d78t3q6IKAL7FHHX+gdjGtCjPv
WsYlsS/BLAkWSznQ6oSCJpxNo1q9Em9C88Vphvlf1JzlebdnE+TCsXNRazMMaobXjTRZ7nVJIEvM
C27G/bE6yJZOL61kGwkb1xEjGMydWhgV8MRLuk6y8SikTbNDEOn8zQlmGnOMKSbT/I3u8d3wE6Is
Yxp7i1hRFdzy4GojhnLZczok/U3XKsi+BFiueA5uZATbaiadOe9/wa/UC1hQZSKVNUuMnCEQA3Ca
bx5pMdzRCabIMGeMGY4IhhNFL89hvqwZT+cyUoQYnt560q4cmdBgEGj/0LCLzbsxuThxhcJ1FzWz
uOvgX8ifn5QRYmvu/oCRXZm7G9cbropFaMnuA0L5i9Mei7HY8evLULhhBqDVn+ueBISds5ehzt8Q
Es8+d9yoBPAf69CQ0v+2ez/DgoCYrUMcwNqMW22ECnSbE9MRQucZt9tqJF/9z+xYxr4Ib70lnsiO
NvwwBfhFONvS16hGOwU8Q6hunI6WxnjzzMYM43KEGx+IcTOS18q4gJHjHbIJcY/Q1qz8A/YirDGz
rW37+n1+zjWm8mJCSX15+rH4stahuLWZkm5zxcRJQ2jVzTPBOThgbMTOOz3I+np1ey0cb+2xIsP9
Fzt29DcybJtv4s34nXfae6UKb3s0tdYVTXl6o4LNLe2bdyrV2mPxLV1SeNRUl59jCPnRxxGO747y
8Mlv+piByxfhj+w61beBxjxDe6iamUo0XzV+3bdy7z7hh/kl/rvIpbgQR1nITb5/PxvmBo0h5ryj
4SksX5SiYqEq2MSl3A1tSaA19YAmSPB1SKp/wsZ+GXArLBgYwACuPy1IG1ZZXrPkcAYJasdMG0yS
ySDd1n+mF7p9wRcJ6SX5DkzkZH2es7YciFiq/TdNsdVUz3SMsRFttEu873QyD2+pKcp8KvF6Dt66
py+CDLUwaaKjA+HuXjhbp3iNW/7HnhUjlx7UFNLAGfDeaw2xdm2fSPXWoB8HoclT5XQPpphXE5fw
+elg1PUd9li2DqvBIKtF3OTCY3HQ4Xw2/XnphlsfEDeHSNUccArl6pXcjqHS3erbRhEw90M040vn
4Oys5NtfO/GINcVP2V+r658tHigxCScWNvY1QkBjT8/AIvas1SrlmhhLTbtzESfgsMbSYqzg7zd8
hnQIXWKkZrPBWoSbtqsanYkzh2J8R5ZHZAWwwsTX7J5lfnG5wZnDYlQ1Nb+x7gN28eWck3rtT0cb
GcrYEU/R2E2JBuwGJsemOiC5kHW8ecUcl0nyWPY9zY/vZhK3tqG5nSsw9qEIgZoI0506VqSouByk
ELwURNFwyrGgRDVb4Tx3wmp5qkUllgilV1mRyT5tXLlRBbgrdH5ng+xl0bvb5EatvA7RRCYk1B36
N7V0UfNv/xjBCJSUm8B9+ywQdIrZ2LnRNntUgaERM5eRJ/nG27faEtflBk04Q6L9yXYxmp2/rG98
SaHcI9p7lTgFtXdmsSUGd3RW9abuEYrgOsuW+HyiKV2x/gq3zkX/EVmDYwNpuzmFQB8n6GJOJQFl
GxBR3DWoJlZ+ObyzhFHq0agYpUNq8NX0o/EXOhEdE4+na47gEZNX/2awl+ya1xhVMP73POEV7lpG
kjUI36GP7N1rgQJ2MqpzduD+3NPxFQY9dYgirDBh9KPe9bfEBMU3WdG2vyUH6vfcTXEulwMfExSo
upVWgCyOT6JwlgMHYr/gC+Od/F5dXGWKqxEpssezbKACkbfiDJwFK1AOJ4Tpz1Mq3TZhw7YpTHnt
qXxMAkUkp4/BYNTXtgtetgUyfzmshNjdAWe1pI27hmcSNTQO8+/vglAQup3XjAFnFKcgzQGprffZ
L71Uv1EN/dAjYc6Mds2+qT/1X4oLQWFXaV477Oyt1LRzAqtGV1b/8LfcVy5tO8+SYlUHqXohmSG4
G32WESSA5c6lQCLu7858zCTVRUaieqzYYnkGezEgCzPUHbm/purqG8Wxir0SG8rgpc9ZGQwaCcRA
m0J8Qh0tZZllNx9okIzD3nFDgzxUBDZz/ECda7N73+ka3z90ow2QH7gDhkP8RAflqZkPPAKQ+jrZ
tDuF5nFI2bdEu/yiwKV3gdDIB8tOapVZVkot0sG5NHqdbXKZt6szDgS5WZPcZDeujhR5fihU+Bsn
hAI5BEI4s+4VrB7iRwpAe0tjqyagAyLWFac1dqjeLLfaW7JmTGIKa2P5O/tl3XaIm9k49NmzSy6I
xWXgBQh6mYdjJy7C3pT0N8lMWNr43UvSv8/lqFB89vjl6+BbBmRxM2cdwnzJoH6E8FOtR37Xkxai
Tqz3HXaPkhZexU+YoZ41uTgzmGYqgmNSvBhgSTjlJyqjDzcQLCqvOLwyZNVV/Al4hKrAatTgygFA
fS6GUbPmhy5nUcxgy7RhQ/7DUYDmS7pEgTr2J8xXSZNnJNdkPCvNQqSNV6IaH503koYMCp+LqAOG
8SV1laJzGigw17NyZEP1YjmkQrHwk0q5MWBp5BIcwbuArjfWAeA+iDIialMHUy1YhmlzEMpAzA+O
CXgerG0t/kl0KL1mHl9mwm95HjYTgwl2MH4Cs6GBzhJnxJypEiQv+9FUzyGozOY5Twi4fWenC+ky
MuVk5aTtsDvl1xndoMHNA2feBKBhwuwbomZHp6qXVEuVjNZ9Eh9cFYTE7P4KUxyfEry0T6wBP3NH
weirXswQJ41VyZZ/FbSMUKowd8xmjvyEM5Xxe6HKfuTBxPUbiXDMcFGbo2546QJCWRVlHGghhzS6
l2FCVXg0TcQYzh6uqUI9gahZBmNz3ysXgd1BdCTWSafdCDaxPb4EBwhb6m5QkUHQLPzUSr1AjqaE
UXaEey0M83Z+QudbrFIou7l3ARCPQvvB9ZpKSIH5dBwrjjEXd+I0GmJdfH51gcGkkhob3zY8ur54
sUJrvLhcmQTOsccvraBI3OvVG16szAv6l/UO2aCKT9xw53x50DHoiV0ayKIn2doVAOkJSZ4e9PI8
40gfKpeT5a3yq21QkXZLaDDpEydEY2aW9jm0jG3+CoyEjI3yF3SQg+JPvL2fs4T4CGOC54ge7bqo
OlKm4ECuKTr0D/Lc5gv9LZZChLh3E6rw0hElHMxdoPllG+FJI1ZczMtYoUMzCd784awheShZ+fvb
g8AK+szVdSgrtzGcuITc/LoB41pfZbwSt/r5UmkRRF6OLdtXotd/ePetszuXcrCBMsWjOoUfhOxA
JUrt0DKLsBCVisRqJOBTF1o/nbnTd8pjeRIljhuts8grKyFdbw9DykSDyms77nLQp8KCKnGoiyww
gcwX8MMV0ZPD5gL8ohTWmEEN51tP1KBojVDkcNfqLlBdHSWgp3c5TVEnFk1Ld0DwoPWEzYFZ1Vh1
pbLoBG68T3ooXifdIRWbLvTXPNL6bpGuXsVfRH7krHTuVkBP6v4t8a4TT6S8WQJlvZ83rb9Yqd8a
eLZKGZ0pwXyIMFgesh5Su3MCnSTmSryPEnZ02T64OqlgDxnF7+8Mm0qY6RRbh+Mimy46No5T3f+x
FqY0GU31iVUTaacCmoNJ378d7hwcS8h1MsjabGo92rwUIHldPm4bga9TVwKPxEAUX0PIQxmBkvTI
szGDWIq+Mloqb17gWA+0Wc1iM58hNgmGKQa5C0pfi3Qx06KHzPGULo/F3jeyfTon8zJuXYAaGzuD
mPtkX5QpnipQK9VDXs+hVkZ94QORKUBhJJ4hCMc8RW/IEji2ON0C4MkF2VeOcwhb0TiVKb9dhvwN
rJ6NDsnBs5Mx+YBme8OpSSaPZi60TA6DJp9aJGKOGYoC3AZ7bnj9OagUjDUq+EPvgIvmI3DGkKyN
ia67nhR1fh5EI1kbrXugB8qooMm31ZqZiz0sTr4Bj2R674A+OZmfHCDZttVqUOpUQXUujO9/w9mu
QoQuRUIWmFognbF5jdFpOEJktAPzinpJg1DtWvS5pFELW5iZ7E1CIPG0k4BAt4mpHK/1OMTZxC/D
EVql8hyeeCrjpWqcz+2Ig53vEimgPSorMsu3scECH5UDdRSR215AcrJSvGuEr1QkJYK7vKtsUnoB
MrhNIqO/y//OsA49bUklNvfJpc3Op5XWj8nULP3bWDxwcA7Mz7f+rIAXjol/VKNtj6q0Jq+Yhd0D
Udw3XNTQadiPqHGve9XUEemzHgfkQgFn/RKykNA2E4QA8Id6YHESJZtaF8WU7Ehzx/EMUiL9btZN
IgC9y52ZEfCDlsVOz7z5YCDrlYDZIrnupsynf77SGB4ZKGUgu+3YlV/M9pPX8B6xxyy4gk5jx2Nc
HPyQk5fqbbNgQvzqZ4Nih1/J8XwVytV+ilQeWLTULicCOdGE0Uvtd3Z6xOnKaOyM6OhcxeeGc1xe
hhU5CtRUI/mXWfxMx6kCs01yJN6bBgINFQCNGYAt7jShfuWCvR+v878voTLFzgc7xT3QK98xP4mW
HCCbmVvndZ6BHF7DUnlBHnYi6tv6UZeYSyi3uTZXiYsNRyFv54WgIqC6X36d+frv5wwDAXhEYyDK
e+wxhxpXGBCRDhnpO0sE1yLqHusBWORj2rm5Ec6L4xHevb8KfugATXkYqUUMEf/rFqdL7077sNzQ
3mRek6V3pSRZqwwuMoG4B4710JiW75Wbqv75t7ot9YLVTbCUJ50gmJdgh1+5fKbKKUFgpJzJAJkk
nk/lZ5FQOLLR6H6BbqrzHwa/AHhX7yw8cN3OW2/ldjOLIeLSNuf2t2fOS3zxkDmWPSInzKrx85gD
pceLnjEbeOLdVWI1z5s3dnhI8cTh0J2n5+0p0iwh8c9fei6KWu1Xx+RBMfpNqAFT74lzMXTBixGs
V6mtP03YXN/IzAL8In4Zc3SK2+67VMZgZQVnzfteL9MUkDxUVA8eA39XXKEedlaBdjrBPx9xD3gz
jTezm+VobK74e0N9HuwLx7ODY36+tzw2mv2JY1xq6F2twW7lN3wj1EbiBtfn4RhAc0uODj+VKD6p
Dm7BEXIqxRoaF0t/SWiIB6oOWEtWxgDFEj9ZJafE1ZfKvj9ofjDh1nCc45hpWv2cI4jJzt0qSl8I
QPqb8HznH9E6DQNzJBQgj+lk2NwdPbKMfXcSRbJ2qpXFaPXPBnGsyAkihH3C/oIWlq9n9+07H1hp
exMAitQxJBDcZRXfsbKteQwccm8ew+IgojHJXqNld2NTP3caY3WS2QvUIvAmk90iildPxRGPxCIz
8yqxQcj+d29+oyw15YgNJ7OtwHwlRNpiJQUfUyZo1m2Izmi1yhTU7dees0345zbuyHHcalolOsN7
X9+QC1swep6XCOUGTgVYRN//59CaxGvEnwdW2W7Zd/6BU5hzq/tOsX4cITrM4bSjS5RRdUU7Xxbu
GbqoRE52Efx0ChTKBwQ/BppaMAIg4XLU1tkYW9N6cT4DLn7JD9iS9LOlE7xg9CyCe7iOpnUZ8nxw
LRrgXTP9ipI6SO3uXlyFiegvb/jATNp3F99vLlSt3R2McdfmGdfF9sxbMSSa8Wa6rcL/HX5RCqt6
FyhPbZC/Ga0OZN5jsG+fas5uEJobe71LsLrUnQgeOQGw9eTewU3HJfSG825VkjTGzw1k19Hs5IQw
Tmibfsy0h+ctqfXBjt3OizFGzRdaBxJ0zWjPZccendecydTEO+T/fcIu5SpsBJCxTDCSKNY+XiEj
jN0i5UDG7fa8jpR60mLlxVYav4geL9eaAbmVTJ4lF0mkkw6TuAC9+b+2Oq1Q5I1LuNG8tz45phX3
hi1BragaL/5ANPP2fVcJ3NzmgFYa6LRyc6mcDrZ7PHgKgCtOfKoYi+4k9ZAfwJ/oN9SnEbnuRq6q
8H0C160g6Tr0js5uacxyjBWU7hb9BPb30sy47dlCVu/I5xcHq4e3iO/+jp+g1rL51dVV2F17VJ0L
hF/YhCAuNGaUfHJJi9CBNIgolKiUYOs84CfNYTxVLe8xsyErVCpCMUzi1MRL+YCe72AlxogjtQh9
jTl/yvKbtPLZC+761TNUEZJ2vxqgq2BugAA2XjQHGIM/Rja+O+PYPPvraXUUKaSNYFeNW8/geMuV
6cclmg+zJPSklVZIdNpJbYomkbiXkzDRFL14KTbrKf0wmU37MkrLKjtOMVaXrOBvbP/l5633gUKH
aYz1Zp92yl03qeSow3NEMAV1EDQUYxfdjU/AxgAY8yKfXAINXKQyYX8as8WHIZIzLWIREnfPvdjE
GT6V9swXoaZ4iaTdST1qkgz6kUHIql2Y6AuAUOAxLpgOlvZ18ASQ2ZQ0eEuAlfiMM3YgEJzxG8dQ
T7l8RHGu+GstKVnls9rViGokJJ42PeUZQliLB2vTJHMULWGQrH5ZN8HBEYiHw7DGMzWah1Fvt1X6
x3K+BHeyhltecSgaLsOLg+IG0W6CwAE4evSX167qhEuR6JLrbJx+8h7I9l+jhFDhn+yrBU0aTQu6
x6Uo1UlHSSiUGkJVwyLGQLMW3ZoS5QuRU7dJuDy+SQo/vd6+Wadf+c8TQJCAy/XrKu6JDf6ASixh
ZzgSyZdddlyG/LAHXWd9U4fu5Qz2QAfy46YQp0FoLIadtBwQvkcrGa0dZm+ZK/sMI14uo6Xlye5C
771nytLP/KrIcNm8r+sRYi2SaOCjLIZ+S8XO8gwVwYRxBJTCD0Y4mY0SFp66r39g/Hyc3/gS0DiA
VX/S7+NhAElTibZICAmPh6SvBbRA7zz8q6wiwy8InMehx5nzkukcpSSbKUeOmjDH0Gk9eaFt6n3S
+8YOHrXMI6t1FRJlpp89e0NamPd07MZTNjdOPHGEguH623IfVFhFSZYFYC+OGGmTmumoyuHYmCwS
C4dDiKwf3yESwoTYW/Dp+idYHRStYvoKLvtBB9E3VshN/Cj7fPpXcIpZ6M9OV9U8U9g400WLFO7Q
v66vtde9Vou/+hu8H5eJWT+/VkuWqKG+4uTwNL6MDELkV0iNwqR6GcbbaVCQtjxVQVbJTji5p0KI
H/qLSnK7SxUuxk/hfzRqVssksoAdozXqyMaDW21lCYCLyBUmL5payodcUbX0vir0/x45muiSQr9J
TmjjezErfJ/vYJ7FWN+r3hWUGHKqcocWA6h755ajaX3PALM/JZErDbNTetLJ8oeZnZvZm07yu2Ub
pDwAXVB7BZy3eIx995AeqOFtAMXld5DqBeuxZEuH6cXYGBJ7+qGCzOIiLQ+25dWyc9zzHQ9Fu6sU
I7N1qbfKIyc8oPc8x7rqCghsQRefkUdlIDWHh0YXVxMiF7/jkXtzer3WNqg9jr9/5C1vbYXMKVug
rS+Mz9SnoMSvoLl4IgCNTsGDdGZTiLRn/Rvw7DUX4IJGbfF1fjOW4tNVG1PWz6NTFlxiHXOthouI
o8qMjTrBhNZgPf6EeYhWQ76vT4lpuJ2HSTTAvwFgXvU8WvCx77gnflOnYOyviyHocDQpWYgWuMwG
BOed4HiVGklzAHttjmFs4JPJDEzK54B/umrnDSOEiHoEC2sY4ARmuml58ugW1fMqCUBz9Tmc4VTs
sUGHBgcHa7U1sx+VpzdXfKtKqbuo3HtPCqtAAZyMhHCrps3t21pVdBngo3G5X20mJnj1z/v4KDFv
r33Uy1uWF5Lu4c2sU+FhHeUCXOO2/Datb8JOzh677j/Isyz6ENviBYAOmdjWM5J7o+ZSM0lOV5Hg
1orSD80POUShHGqhzqeHge5+CcDwho0qFZHgiEJW4T4ypvu0OZTJJBp57LXNvACOrJYVybd9Gwe0
EchtsDakmyA7i/tM95x5T/Bg/uuzdLFtPwddP0Axn692D5OrKSN116m+zz/WL/mvFk+XANFwdDHC
doNgHoP780n1uXhbTd7Z0CI65gpdnq3BUNTGoMsF958/owvr1+x8t+WYCXX6GYxL6Oc6kBYEJ7wL
xhAtrqT9MkS+bVCAZJnR37VjNNohMZBQcQg7YGHzMFcBkKiFXF4vzP7t38yz+bn6OhawxOb9Vz4+
Y+FENNnHcLVIK35DluUoqlGj63e1igfHGKZXPxUjom9p7BmhgJJOipdG95S7MZq9DZfdWt743/fk
k4LoGwpAjIKie7oPEjQUw4jJEIbhB5gnIYFxVRWBQw4bHlcLwohh1R17M2t+WE7M+hyLze19BZGX
8Mg4S3aesQDUk3Hr0gTG9ZJTd9VahRX7qamAVJa6YmRe5UqQkwkuMuiwzMNjMolXaLCRjvZTw1C3
mB7CZ73tR7Vh+Jm5Csd4nHl23X4P+IXbgq8p1zlglCPnl12FkwkR8G+5VCyRfQ8VjSd2dPPN9+/U
0LMsFYSVaR5Ydg4i1+VXm6zZ7cyun+UwC7HLNoyhlMun0rEx63DN49x5FriKkxqsP9oWP9EguS3N
hBIi2fqBWd2knWIeqiWfrM44n5+trxR6D3Sn7ny8FQ2+Y7sjb1TXMRSqGceSlpTL0JiBRBKoBeBT
U0fCVmTm6ZrnkrCGFTMMVPr+zIlwOhRC0o9446ds0dG9RED9/NiQGYxjsr/1C3PqilTfETkIa+tk
SiSPHtnxbSV7/7ihJKYI3tDfvK/IoXThboMDAvlbJyZ/Srzqm1tf9qlCxkHDOuhM5O5lr5Ek0P/N
Min1UvI/W/tTEgAJVi4R00XcCigpMu1SP3RVte8bPe89XHkIRefYLNmjKOLnsj73W8kz5Njx6cKY
2+65IxkWJXzDROb3CCxZmohWxIEiDUIaEGx9qcO/+nyDXf4rQx/0jST+3rmfkESt8vURZw4DMBfl
5nMD8HX6qhWsRhZexlxpYUfG9cUweTZIc+Z+TmY1ZtRpsMDjnRdlImS6JetkBpVNlZg8QXDZVLhS
9fFjiVqGQbnw+5a7v+9B27CL6oEZBjVfnYnvMiJxI4QThbypSyi9REzgWycYVQavH8GA6cPsqDlE
pXmaZ6fXOgXWa5D2IfeaTGuYAxGZ16nr6tWDZzu/HBnIAVC5ffzZO6tr5szLcztDTbfNRGr62hgJ
2SutWmCjaofSSNQ9U0JGxvE6tw7nRMWKEkMziiS1m3Vxy35OAwh1xauW7DKFCAVMOc3mfNaQLEHd
ZFy4YW40jKP2S8GScZafV4CGURBtHHVgn1j8YRh4BavHzBD732ONcHn7iWbZs0QaAtl3VJG28W8t
Ul4+pj041bfihutWH2xH38C/ryPDYmzQEUEBOmvy9zJ+DmDO8ehyioSK97kUsKB4dSEeib/pYGnw
g0NnJixxyp+BRXtXGqJ9Vqwf9ZcfNeIVyOOzx7cSvSpq3Xikca8rpgy8t6Flao13aS5XoWuJYGoP
7hgm7hNN2wJvWqh59EkkaA3xnM25K9/7dzV01qiW5mmfocqHtSPutZ8D2B2ccWllEWIH7+e3SHN1
Gce58umn2T3pfmmDIycpmdlzAUjlxRLuCWa/lMb4xJ5xSfdt/PmQcmD6jec6xMO9gljI75MQGZf6
6rbXQq5nmcJr1xLxcUqZwjxnelo8Ub/Fty+v+nOxZi8Nm0GReBYGn4WNPTslAZycmq+u1bIp13q1
+TrL2tfjWPz0TuPjPn44V/FxjpjZNt6N824HC7imvEoTV9HjRxna2EsTKH33iWoBXmER40O7RWBF
f/gb+o7Z35u4ArL+N2HobQjmyZTz9hwL5g7biE4XHSxCEVs1Wy8YEXM0du9pJNc3wuWimQjcarGQ
dwmTmsW02mRhUJDCf+R8LdsuxfOzzw1QQpVRuiquNPv0mAjMLQhQjwkTN7V+vj0BRkgoBhGK0L/x
wTqQZ+AKgUAkjFMuyMUQnqAQBoFmlDHp8Mnbft3XT1JmY+wJWpwATKZzWn+H++v3JAfGfz0P3VbH
36wtepVapcCC2opzhyRqejczFxDtKkqkGBp6IAZO+ZXe2RB3T/FLMTc8DXSzDpLJ7UJB8dzISFlr
9jwLHyFmnCgMmk+P8C0ibZbxUJzGqipX41+aOI9suhnfhva79fgT9fbYE1He1/mzn6Ytz8VI4xBM
09EdJVJsafVe3lo9hN86GqwnF72s6sFggDRRgJTGmuXqfdNCX8degDPo7NRTQ1+zxQ3tTrYGPEQa
3TYjEKud8llNLdkOns1nkZnpvtcL2GB9yfCfHM3MY7ysyVFMTOtOqADKTfh+onqrgwTFMIaaLMbR
rR3HVJvDZWFQyN5sg07fwN6pogDCs+w+vHmjXxnN/SG5r8u6Rhp0zyJqmueNPcvUuChs+GNTIEFi
I/tuIojIS67CSrY2awLRyFaCPz39dkFyFsL1ksJPohhgVYTi8mUZmTHP741qsYIEGeFSJ71d9+f3
2u+edoMbqWa0aTGNNWPtcsGKHLHV7WNXay5xSA4DJqJyzRTU2UUX2vpW0ig1qouYxAPOr/n9Pr+i
1pKBnmxyMx5k4t8cjUGJ917dpKNGVTHokxIGblyXvwwAxqf8CVtv9LRNLw8iJqWAzyevOOZ7Xm4C
RO/2yHosASazXuqZrawEsHz3Yo88Z5dgJeCGqw2cn2hEkGAWIs67q/CdIkAeUPEs/ILAwxS592MV
nFoHA2Y0mtTqLfUwTSu/sR0OKDH3Xh3WEuSuhSKrNo3eUCHoVZX5qnVH1Fbzfc5V4ShBGrgstGvt
ab+saQgMTQKlm7fp/C9ic61H1x0I8C8YU7sqYm5mJybPNQT7zDcWz7emiT1UDrz8mx2zq72C7D1f
2OAxNVkmhT5SuQR7k+0iN/nxyAsFnRK9LsfJumUFRcBWJMyK6wZMcGV+wyiZnheWLmAm/R1K9c8c
FVBnTFmICWJIkjndjCKi5JdjBOIV6ASQz0t52r1gp5jZXyjG3rKMG6pTlPbLPEtoZDORJ2ISaJHJ
U9FyNXXsox8QD03vvM5HbPGKF6GVBzFkvc5USs/wmeT2E8zFeDwAaMQzOcE5o3BHLPUPS9bJWVc8
oU8KM1rlFTaEyeSxXgItsuIBjRVF+7HDTIShu+JNhpaBiqH+0hBwqYG4L62kOuIkKdcviadbGBuN
HYy5ihFEMHLh4SjVCdqtqkRPog1onfMa2V8ip35eKpmP1Fq7T81aCvo0JYZ9MDo6x56oEDR8DiBM
0uGn16/zorw98sErP8Fn0Io03T42HQay5rvTeWkKLdc9GMP0R8pasFnZAHdGFUBTV84DPddU9x5j
NPMDIZZLoPKulHSFevGKp6Kx4NYDo3Q2RmoXPrII2K8XomsXgMTHnz1wR4l/hBGGH7vnK4rPvdAA
g5E7rWGE1DX4xQAz62b2SsLeF0PCUrl9sgQAvRk4Xv+O0Fep+i325dset5LnalLFprpEguJo5qKN
sDMdfHdngmnQhPXaQDlAAmoosM11efgXk0+8GwKGozF+6u866llPwATb6FAz59RtUIOnqVYFmZFN
vr13ffn/ePPbpDoDOM3TJ2fon4dZ30hxUoDb2ltYlmRCeBHAaNfffJNDsKgmITuxzzKiWRXs3MnN
k1gfQr2G8aVW2vIXnglFV76C6gonb6UKW6mCrCPbevBASV4Rp2Iys9Sb8liCCzimOmVcmWoiGMay
sHlk29lIcllaqfv6TaEUtz4mLsxAoQipiyr4/b4ok0G4POxeTO7LkhWo+C6MADrzB6/S5LZ5by56
aFrXiMA6myytSegDKWCur0Uj5VjCkCU1zdlDyP7SWw5UJoBrQvgpBNwkfE+clPa2fwLIbCJAyymO
Py0dKtSm8Fg9AhftXHkot8nSDifbz7eukLKPR0kLRrInaovTQoqRSiXKsjy/W6L082+ZnUKyMzf6
TQt6PUMiEaTCRSLU6sAxU3CDOXWscflB7K41VPljUvhMmVagEhjmMe9q2tRZz8B2n3CBvg65hQul
3DeavOLeWSTWG3vnEBXvZDsRlNjyhgrAJ6XgkvdU8EX5NgSJrjZs7MBph+kLKdkW9kCLNpahtShw
ujUtAQGPA81eRNZFkhZ/3QaVI9XF+Qmk3DWNdrYk+KAOYPJG82bNGMc3S2g0B3XRQWDuf3HBQqdy
xHranDXgMdQx6PR/cULoOJYrPZ8fppNkg7C/BwTMj23/jYqnH0ZCEpae92MVfzHjBP+ma0yQXLnm
ncX8HTfzz1x7lnlFWOQttS7hy+QAGBXEozbV8jz3+yh4nbWGWRDfwGb1RiGvqGMIzvlS19qrh6ax
HwRRGs2QGkXKx6OWe5Af4YzZ3uvh+tRjFZbyZri6GstlTM27lW08lqTCls1n6Ig4cSulzAtlV0VW
5s5ZWLWI9CC10Xta+UM6niR4Qu9S8t4vauIgjKOQZExk6eGtmZEwPQrphwd4p8ea0QD8IDmCyI29
BqIVPGE+3EnS41WKvtQYKbdIrcnUeUKJ5EmKG+WHHuj10GAuNhgvJsSOFGo5Wt8sJdaxFIzZ7Wag
ARUxSjZLuOAJX59etk0YnUxwM/Gat8PS9SmtSAfh41/7c2tQRFozCADmPyLmivL+q1L9HQ+Ts+/h
IX8wt66yzb8uXxmjo+XpFhzkKpTg2e2J5I5wWQrxeaDicL2jzFGszQ6ruGOv7YPWW3Hm3gMJnguG
0mlfT/7IlHSnXQVaohZWjce+/T8QUE4pjXTPks3jekEgXQYtuIRzRNq1wQbPVL0KWoSh0Y/QuNhS
Sc2+flARcpz1Nrrf3jZcNxklivYiYL4YM5ijPPFowbMzhxEec4jRW61yyNRROS6OE3rjl+7jbatD
iXyMvBFNwOXOvDRI717e2ouQ9XrnFYQa3qXKzMdTH4YsYRxrhap0noLIAQ5xJoVA5D0PkwKA9sVQ
fnybodGJwLf+FEa7R6jOTFEGJkA1nQWqm7uggI6TBffGLmWtBuCh+NzL/uTAtgxu9Ogzn6w0WdiO
AsBbjNzIp+xw6pHJAxV0Da5xbhc76g3TN9+/sOt1rERHnx0tQ/roaJVadYkKkmMKO6iyjjOUYNc7
ac7HAEMlTMiMdKdE6jEqQohZOn48p+gOMqSq+7cAw6WFiyTLqYXhh19VAqRv2rgCkIPvuFLSI9iK
dwokrkbL9piXD4FScwbmN1w+fbA46qmLiL304/OFlKNToC3hoVhZgD45sjMFQTRnp9AUYG2JF89T
TdfPN4YfEWhwSUBajHc6YMf16tBaGwSMS+YUhzyGIWB0Qd86cdwtYukw0Dt6eXtL3CLVq0HteuG7
MD8w710roQpiquGsVPtpjPtRZZHQusMgsCv6zjlVkHDTXqgqufIEvaY397X9cwUHbypJclweMirp
F3Jf0D4m53rmmHJ2OdIEfuMjRxOfUnu2a1j2+MHuS6lACQxK5tpsLieftuoX0t7uWwIp5zw0+SwI
7XJ/q9esXPMDF62IV7RW2KWD/lhwpXVTQne147lZbf1rqF9xAQgJiUY9z280+JkqDBXKWRC8k54G
TkXhABRSiUNOjub3pyegyyrp1Fr7XNKCNyqTe2lpQhhJn9Brq7zIdph8kkUQ8OATxRzsY6w727ML
MBB3JUgy75B6T4lM+SEQIPUGne9ZYez2/Wugt7M9uEqYmZfdKYM/QzfpebanZlWt2E6UxFgbJloM
kLPrYA/8HRRMlStQ1lDtGlnHwf83agfI0JRHnxSX2XRkojom5Tn4qvVVlTC98vuCQ/mjPDASwC7T
7KQJujvY13VbAJ4aKgHfWUgxaiCdEsAIWLqa91qu6hlOQeTTEyIuedwPVeZDRs9tl8yREBn1bB2k
oq6TVcYg32gojrJpAd8ylJ0VdOQkno0adWrcSt+3s61ReGDnv5d4RLmaVMOm41h7P3+OeNHgXryx
kPSXohLEzYVmAqnsRyR67rEL6tK0KFLsumRPO9TzSM7Q2eilGFsQmbLkKdCCMm3nd79BktO6TThw
shRN9fsWSd8HyT+Fe0ItcCmhoB4Yf2RAp7JCRutT56uaazBAj+jVwcREg9Txd5haeqzi/4T8rQj3
NtfF88/x7GKNvwsfk4JfyaJctzWdtcokhUVs5Zz7vchY6SCuGnjEvF0LEJjUvNZUSMg6U1D1ah5b
P15Gwznbbupo62E481ZvY9oKhI89qe1ohpBZjPd3iA4+HOzVwbUfpeSBsTRlbH4bANHJ7yj53uQ2
1Gq8Fsv5iLFiuL8Zy2WlSoItQQ4S0RS2IxeqtPT6sQOPy7c/bHRlA5Z1JGBB+5f5Rf31cLxwR1Lp
93UyskviiR9heYII4UDLzTk77Ciys8y25Vi6GJ6icITyBl/h/J5j4PXTf/2g6cYjQ2QW4TdEemPM
tBlq/SynFAKM9CXPH9XpHJW/+8hLmusNmLG2/W/n5hKppRx2x1qFbVGKuQxStvNd9fQAXQiE+ahA
L1R73bfILbYYTQU2/2sZuemrfrHxB3rHP/z39jIRxN9BG3O/ohBgzij4Mm0HH3tf/FKVj9rRtrJw
2Zjfsx4L+48s3dWVSymUoEYMP0XthEjwuV8RQ329wbHbUjVVYN3Qe7sm7tcbeyhEP9x6k61TY5Ob
uZkhPWzOXYQaPbAKTgSMo45QejHBGAOorTHE3+C+t9GiSqCZT5tlMkxSF5SlFW8Jh0qOOEojqPat
9E4g/C2o5zYzXDtAIY1Mrj/m9Eh74ozbUc/op2ejVaGtWGZJkj4m0WMja5VYUjb3H04rZz8sgjT9
CaZ/I3Rjs1EUMpXMlG9aqIRRXxcK99uIHE1zWPOk5H+v9htYnpCltTwOzy2iTjBjXF84hz9IPyC/
qYlcnt38b7ko4VpZQREbytwX0+dIPv4e8HeWSBhDdeVABChTPVlqGtid09kN4mRXnnSL3vdesko5
19VO5ipSCT525jUE46Yacc2A4AoqX4+aD7hNQoJsLo7k88qsn9ZNgQQyndIRi7wikpqwUtiPQ9Dg
6f40rCeaNjH8J8NS4UQpg4nX4UPVYQIPGVdj0FFZZqqNNBuxuyKubLfq8Xnu3yRtYXlDQC01fRjp
buaXERGrCQvQMyXMkWTVnDMiXF/SDEjZSU4SApi/4kGTndY4Ayc6kdhNa9oJ+SH3K/CpPQtk33Ig
p9lm1LuJZa6w40TLBiOVTIzJ/weoQfQzsFG5SWm0j/H4p0a4R7/w6qcy0l3etRuRqgw4OH8XktKb
eknD/ggFM+O0X1+tlJfi7MjvYshVY7Nwof00rMGs+jVXCk7IYE1N+Wbrh6dtRnTrwfLhHuo7d3w8
LzgQ+9/RtmitN4QFJ8/XSswJtJLICz9JSCrQlTbesWak3W0AbpCMYGrv9zaeW8ULFmabDt6otbzD
gFuTUFWljnMxJZPkYkbffZvbamgK0o19wX+xG2dr2ryd7jaLBfx7z2ttFEvxMYyK6UPyZA4uv8bP
eT3GInDJcqtkAqKENnsSNdsxLGMpLcY3KAtfRbPM0g8YVVeWrcfT6rwEWam8Bwu4DRWggoumDUOC
9CNh+m7K8+O4gBVeraIRJSc+CAmbuGFhzytj68OSTPyX6quT/3SlLRlyRcYEbPIH03F5Djw2KNoY
ShHQQeUugCa0p9oWIGYU+pHXTFE5dmBdJ4heygsKKI1AcLuiPgp1G8POzSXMaWI6vZcpAmHCuCs1
KsHXKH7zH11bKKnw9WYdb24JcWTl91nAA8pVdLtswQpzLFYVZR6pmb+i4UamJjlbijljnJoQ5Cim
suckQmbqnywl+QhXFqVQHGgkGgC9Q0D//OtOT33GYEkWNQZ5nHPFCupEbvlXmWpjhkRQYX/AOv+c
W/aGp89shorEpR3u7mA00pSz5vXIIcALVhlUe9CriOveMepFeGyRepZb7fBsPf4hFQ5J7TI16cAG
lgM1SBmu7gbxf0MA/Nq2g4mbZE+leBIwHx35yssA3/RJB/86wm3hP7GgSJRp3rnrB2NCDFLz2BiP
dNQ35+gMBt5vJvu/jUpPnOf8/yqKdROdeyGRF+vu8NOQLzz5DccRj2xeVXTY+W7PZ8aNFCbs/750
kiQFkmQNeOpg2Y/Wn6qxHUc0iEX9eWGA2R432W8j5hBWYhOkZrNo6msNqR2KPVZ8w8iMArQQycBW
RIN+STDLOPTT4YKHo5+sePMlc9dySrsHp46TiOytyDL9zigSCJfa7oVwYo+DAW13Ny/+g73aqoBO
cJ/xfcuSwiBXch9uLv3/NoMr4p1f9IWAyD4YVmhUDxwWIIxs1Ivqeu5wHH2Dnqoi7bxItH69OBPs
l81NbxsoJ6TwYGM65sm9WGayLyOksXfYTGfWjaGmrCzp9IDG4s6LNPI3o1AuDOwMwHDENeoIxwNt
tpmXIDs/rRmjXApHpwfkXH6U6rVafuRkzwQaLJOwq/yLOqxRThuVY+GcZpr1GVIFxaFMXGGSB/Jp
agEYks+cRFX41RmVI/hzszVHAtV2sfS+h/Eq2ukqAwxO5C9FTDlSZpph+e9gG5EMv3AyD+jSLfsa
trnoZ1cTNHEsrvSK9aQ961ymHgqVPS21vcrqXbL6oaCwGXC+zFADa4E6E9vno/Qk9U1DMtTB873T
eFVTWxB5jnzqfFL5+Xc3O+f97oLV3twT0ApC9JBJFBVLM3W6tX9ECVDCZA9ZmhdAkykA1h1H+N4H
6qTDKzYOPvxFoD9T1tjtLZERlGNDj2mRjJXB+y5WE9mQfmdUlPW+uNyIUYcpqwXm6+HJCke8Y6+T
njrzE1njSn3nfA8d8aFvXTBHxPnIkawdbrpMQ8eEOXUpiMzZTsnbrIo+L8RB4+oEFe3eU8BoPHWq
Th/DuLtEfqHK9AFnkYsUGUc1oX+y8Q+0aUd3CUfYgX6gGdh/AzsIjjb09EZQucgsn15+b5+qYf0j
n9LASjpXmpyD8fQokcP0tHzX+ja130/H4CYl+AB9AlYhrzgFO9Mkf8gjvPnSP0UrdKgILb6+Xidl
7j75xwgBbUvCS0s92U4abu5WfIY/a35SzZT7znI5Tf9LWIhpYBYu8MSJWire+3blM/l+ARlUem1z
e9PTGFPIKs2RG8DIREcmGPf0sHFX8Dm9SqIGajwuHWFppCogvchjjoqPYTZwc9LE4fRHnIsmN6D3
ZeBkrKohBb9EaCITGt/nxCqdK/IujW6m2uikweG2vP4CMRXnRD+kevA5aS8aNaXf3XQloKu6TsAb
U3q1pnZfFk5cFUFUP1KT/19GPh6+DTjvw7tg+md20JUUq7IY2R0Nz9Rr5cWzy2/wjX9JrnxkE7Tv
XwBJKvnBPx5jvYlRRq/5SiZ4j/gnow/pUFb0pn6CIkw/Hn4XfeLcYN0asRrOUhG9GWuK7+TBGDgd
se0c+n6M/6EBfOYaPUF1g1NjT5EW91PUMl6brggUuMa5rG5/XK7ogaWh1RuYXGBgDxYBJYsbyOum
Ifr7nKuhhpslPVukWIuZqWeJg9jHj5cs5oBqjKpPM0UoWmTIjk6v9LUGv50zT8B+mfGcS2d1tPxE
u1nae1z7gHPFTCFNlAq3hLa+RFxfNk0DEB9sjnUu1Y0WjfOTkrS5B5CropBCeFJvl7ggU/PQGFBI
MKvqyPsEOIGYXyHyBG1mb7vPeV4aKpce0SSSfvMOqJXBUB8CoGRB/asohk5CAxCSt7ry5xXGuhW4
on6RWB6pOWGUZ9EPNW1Gudl2H6ebsOqT7BYvmxxuARZsIcy9jwma203Nv4narKR701DSNgV0Gd9t
8sqLVJYRgv5+ogZHy45rjuiQKUb5byn4O+ioVGYeN9U79WWbuBxs1DvaWOWqWrXm9s7t+mI4XsxN
vwNuqGpH0QJYvj6VUPt7Ht5q4h4AM/GSVdDDHusrERt06F4zmlKKHKMveYSX5KjB4/Mq8O/Qv7uB
QIzerCj5A2wQIyZEPtGxA0iZK8eOfraRxV/5qT94U0Cd2e0jIXhg9i2KD9fxO2H+cGZhq5KPIIu3
321DtkF1CF+JM+axBBatHZEAbF9Kcwq7qmCtTxUNKoU8T7FYDdsnDq1/v1Yx8ll1V/neZ2iSWNJl
cK2F6V8UHVWoxf05QeAq998VQT06f/DUD8c/46ZU6Pn6eReTdOs5jEj1IxXBUtl88nxAsc/j3lIM
B24k5qn6PAExca5fV8aqWP4ApnmfwKvlTRG6w0+uPCxWVaCMnUbnZIXrVSVoZud5ctTO5Y7S6gcR
MITSFrFsXYhP9soWoI+eXzKDe3lAN8Fr67iHAm9jK0cH5lrj+0ci3lqE7uvrIlYeRTwNEir9a3NO
XnkqSkwI5EQMLuarusrLBn0DkI1gISQjkjX0ss/iK6AoLfjNtVhDjZ4tntqibAqowrQYsUyTg1V5
Ha3kZyuZiyctNfLxg37VRMlQsdT1N6VtmpDj7EP8w0sVMKsqRBFuRnOQeE3ru1Uh0k02RaRldv/a
+LB+rFppiF2zI8L8TrRjvNf53P7uWYZAm+nYqRLJkxsUeEnn/ngG/Xzb9TgZBS/jiaFPGg5pyzl8
qXYEC1WIbuYIgILnPTcmzsCpfANJPQNBtt4ZQPVOleZO2H1/e6cwFVpk+Ld6tq/nviAdOSORrxB1
Dg5TE3k9SnkgKBJw8SyP3rbV1/TDRFvQGJ71RbsGuOPuRF0najfvCRKpr4pWwFPC82D3qYHZUl0I
ZJAGaWbXFgUgxneJSYiWL/WkSYoVDInL6u47WhJjsL+NFgz9NTCWiM+9RjfUs3amGwaBK2tN7v6g
OKAzp8Vz0kZQNSMwVmyBp18ZS90VFOMKvd1Wd6fRRI6v7RLjc7jlVIKLoWc+WRDDEhDs06VZzvA4
dHMkVyq4NiNJrmcbT1o+s18ynssvOa5Cj9GvMBdzUWDr2pAyG5/qBUEKsvAthSD7Qykug+N1ybE2
A3EQPNidsoFKSdZY7C4AV05rxQ01p9m7f4PwlCO6Pvg4EjrOMecC+ptJk1jJ6DmC37RNIlHnSU1b
njBkSqXMvDMlk/CCoyzvL2LvwLcGVgkgwFhalUKEGsOjG6Vpjph23Ni2kRwAACbOR4Gp9BYkMnAZ
W0tf326gtGKq89iHK+ixXxhkggPTg4ZIDiX9Extkkk/gbY9Jp7o6s/DGgWytNrezftTwboJRijBu
SfRhlzS43Dcfx75go2A61Arg0tO8yMB5AOKr+65HgrHZkjcpZbbVO91CULR7WItksO2rFOoliunU
672JOgoOUaqmJmlO4vtugg3mYWoFKpnQOVi49MzPEgHYYlb8AGZckaoNo6zMxM3O4A/tWbgccgOw
hrVQ88pLuWBDrCajAp+BR2D75ILXWqWqmdKBil0QYh8cRpGmJK/7OtAQobmWm/lSr5uNwExRrrsi
Y1Pi6NWmUDA4rDm6S1aj3MAxCcIlWNvdLG47hBHrCWf5nctajcQNwOa/FBaleMuksbTZ5n/PSQjU
rt4URtoVuWNbjlf6iyQmspz0yc2smGzxdrAXkycIy8+wahxe1rgRShGB6He/35DJPpnalAWQcsEQ
MHn3CkzsVIJOGJ2RMB7x1P1nWlDNH1KokGasL0zO8oRgheJVyfRBYReeDn77Oo6gWnYmSUEvwBTs
gead452I5qYbqmNWiiRys6aF0DTPemRuoMKosf4kpDmdslQMn4w9vkMT+goxaHe9PTWUdeTB8Jm9
eU5s1oHda0UG+Bn1oTJJ8jHAN1dQY0Om65/o70Dbivz4tXytMeFpsuciw99tjVPB05K9npM5b5y7
EcOyXSXWwr5SwmVduBFECVj/7CUsw5hdmMT6PTD52MIafNjeazwnCM8OFwsWiwlJXFKBtROHAUpb
VOV7HuMfKjNPDINnHi3cTL6PAz0EUvwhUfH/AHPo3T3WavG5UC05qPbyBy+UDMRt/0v6Ytx8yD4a
yOwtPdx0vDMQ+faCsyhi1X+lo31oWcD0gl775rya99IX1o/bomkRJ1srFqUGaYqbrn9/BS+oSX95
njxdHCsarCeq3z+cqyn63A+46RlkQr3O5iVeqVwdstPEVgvSPxQs3NItk/BXBgI+MFz14IbomKo1
j4/7Ls5/cmSYwssERGEjbaCLpTtOU2Y/dsa1lfZdpuT/E/nJxRzWNJbt0OvbD3wELIcPqs0Xwbcl
1bpa0kCSiEBPyEVNgRa8Il/draV7933Q658FTQgfnCctxPgBvLDF0Wzie5rdXU/LiJVI1WKPh1de
XF/p/99Wgx9I/Lt89TvlaRl5bfkoUQl0dxKYXegklJ8FeGmJM3dY3/Tu7CzsUXQB0UUF8S8lvYmE
e2Sm7YR2YraVFhS9XE9J+v1ZseyNEIiYtiT+hzc+4F3KGDTboEHET80gqrYt7cNbqp1DGoqplkIk
wEtKrLeAV/Mf6fjxDPy+cVQmpSt/aMQ5tycFqi+DKcfYQh6EdWdOFB49f5G9HSjV1N/ocLJW6oEI
kvdZ6E7JtzpebNdiXr6fkcRP9bSqpR61rH+KGtg3YQhs9349pvEAkoWPMAK5M5hHmb/GFS2nonw3
+nkbwQ/T2mgE18k/x1WRPEhEEjQx4PUnrCgBALhxtO0pJ70Zl5QvnOE9M8DA6T2FXSNaZbTd9DcX
RtAte7S1TNq8XxEXNbGzd6Go5wk5viLWY2QPoxesVFKqo97qK/JkxYbi5Ac+ifvj4Gz/9j60DvAV
rJRG4HNIi754ROFgJTzyHxURRrT7guWy4UkWqDxtEyKEsVYdjfbN8gr/6P9MOpz4D3yc5TMQmY+R
jAq9VzQW7+zFFWpafHDC8lc/+2eNnzMeAXmrHHXmjqpajxvg2JUn5e1/P16yYdqqouxrcRzkgNaj
Fsy7OBtf+roNP0KfaN/752rBiuW8dbFYd3ffQkvNXPaKwaHoKjhVin9oM0L1aC/qg9OL0pBXHA62
zVToX11WCKDd5atM+n+2MroECoPPvJwdTijcEKnPU7kQSXUfo5R/qY+5GYeHHdBW9fMdRX/YEWKu
G+UkTEg9BlEGCdjXE4RBjVcfMyeZIBBMMpCmSCpbYrmJNlOduqSn/gRzE4UniATvkAHe0LEXahrr
39nMLZkq0ad99+sQ76ljLjvvEIr139MCmbYjUS9nvRB1ya09QgKZ1w1fnqXWw4aS0sK3Egi3ZYqm
6EVqrwtphV9PcV2PyhJ3te3HNzn/mPynAslWJzOkqAz0ZoFQ+6QoVs8PiXDwNQBul/T4LQecu9xG
TMFG9jSJrLbTJHGV688qFe7FhnFkKqdXjMU4r4FGEwRG8+8wyxeTGZz+65WjT9pdy7wh8NM0uL0k
4YGujoAsZ6TSJppEni2NrIvV3++gc+BQ/T/O1u8C7hn73YHMPjaSCqMiDEKsLuzj5kmV1OIpts67
kS3AwSTnBqfwRprv3kJ8VPmRiRab01v75ya0UrWQrPe3M/UWmH7TZwoXWzn1Jizq73RrNZMUEKic
g5dHZQcn/qpQH4IhkI8ew38NGukTfUN7yLYS2LOZ8YB+mJMjLyQCjyS4AJ3+PvgG6TjzggNyGTnh
FK/5mT+C8U5y2ust6k/AVf/ZcXYwKPnmS4Da2rpuSSxLw0sJvwtIeLgCYoiN07sByr0pQr4LXImD
7e4I/aXvrFRb/pYXcDg4g0ynyownc37BJX/RMfvwiX8GGJB/t1xt4ljQ/vFjDxYR3zWAarGMINh+
hQYuGW1ICW23JJybO+mMxxCYI5cUSt7wsp8NP4bum/09UNWlBtrm4eztjxIewoR16nh7jRuQaxTD
SHd9dsAylmQUw4p1RRx47bEpmYbXUlTsaBsprNLB+fZ+UUsPsmGumHoj7G8AUuhFU+kQZQnQvzQQ
oneWmaSoADUTQv52zupXYXUsH9Cqlyk0W5KVGASTd4F8aRlVQyTMx8+4JS4JFcA+d9zdOthbe2pd
C1qBdvInvMLMsCc2uBFE8M52pjo5g3LcSMJG6RQGBnHQ/JjXI4RTXr+yeBzVU6LIsFL5U4GQ5c/W
4XrLwIrA1lad1Cq+/JnBiBMILGmvVEC226U/lbF8kafJXKKNyU1Ec/DmdRIWpHZwhTWx4JDDyKn9
K4helMrxML6/WqJWn7mHww303lSuBM9AA1Va8EkoHQFb+qvX+2h9sxcdVjRHmku7iYJBkFihUlli
PDmnHR/IEGEgs8rSQ5pHBo55nrBywbW7/xmN5WEm4ctLmsLyP22s47Nz00RLLkMj/usUvXNjEHJE
4h+wKOPbQn8uWl7VYGl0vRLTu6reTO+ySRmfl4yMXZBuFVEByTL+LD4ahQVhL9/j0/8xozS8nEGS
hwyi+HbHdianmJt5TCkkTwV6PhLcWJEoeU6hB7+ZXZ6jQkQB7YeJMfMBP8ZvZh6zIPiSo0gzWP/G
HDeJ5dF1w+fsnDrxIRt29U4XUz0R+6by+YloPdYKT3wbUsodD1wI0bVQkYWOtkerZJC9I0uapIMz
w0CMFTgs9zSg6kS8K+J/zVTAqf4bB9r3r0NuYngbSPM7sykVcK6FhAf+wH4aC4t17qavMh7ylNYd
Kip92jYX6B8fC1KCF2N6OATlEqliLcjlMBSqYgvlLT9CngfK19I7CrzkkCqTwmoBO7nxAGhvizLu
WXc8nm9ANygatVIhT4f4c0f7K0f2EKyxhgojcvYwAwPcwpT7lwOpx8j2yAjpsb7bdytd99ysKxsc
QUds1aD2DCrOwV22eFWJcjewLcI/Ut67WetXh2Zvx/Pg6uVcLtdCuCKTVQMXLz8JIhVkw1MWwOwL
pk1lRmfzAaA3Zj0Qr0DmfUSEbgcOrxA2fIt7aSLDscmjpJGWKoOGgBCE58kMDdq+CUSOr53LjmJ2
s3nkuBkc5Tt4IV6BFDovcy0Dnd0udNW/1txgnpGsGFAQRLEGByt4mg1/bA5zQ1sr8FIsEd70DdZn
iQFVijeNaaSkBn87VjwcDjlioljsqSNCT8acRng6dMlKNGxFMC6mRgIzwEM+Wk5SGHEP2qBnFEsc
Haul1CEb+k55abKVH/7MtcrV6A9XvUR/68RjShQqY3BxjZsrWtZN2RQqIJDkU0My5W0Krl1eeNIE
r+zHjHYZDRJolTQhscM3M3IADYqtbAktVyM7frYVKPcmladXeCaFwYrz71azRdHZ355LYOaPXSmY
xPVeZKP9uJHqD3UlvYxivGzLxL6W/AdJ4IR+jhK7U3EUjFlwJfPIIHQ1X0eoKpGyvrOdk8S5WGqh
+jN/7c7/BVRkjMPyRr3e1bOTEw0gQjdyvRI3yhyuvtHlDs4kecIkThEEQI8tQ532nqBjfRK2nrwu
UiukMC1MjJ2ZaKSSIIfSzhaIESOhubFIx+KtRrG71s62ZNze/zPWJOhLZgbhUiAdgd4aT79yCiVL
ShhWTx4giu86tbemIiII5P46joKx1WoABO9tWVHkZS2wZsZlwtH4uobogfLAARBpjXTcyrbmWUAK
Ag3t+JFtfRo+laDcuEZv5gQYYxc1eFxaSuHvjRIG/2STwq3WezQQoD4ojzOyqiOfSdTqqApSB6gq
giGpySQtNSQ3Lu9uSwqd0D5KaJsO2DYySJBJaQef7rG0esSmi1seD0ADY0yQJXFPsEVMOxwfRDYt
OqVYA7CK+Fm97jAuMJz5B9LTt0VFigwfxrzpaAUEeNO273P6IYJ/vEXCc39miV0WPqbmFFRKWAWZ
U09xxNwUhX6jcDp4aUtDe7CI5gqGP1FibgiwaIHPkDBzzHqkFA8VCrF2ivX9p475AxljHG1kGdtw
PtcV0IOpE2luxfRcHpUxX3TPp8cj5ZnLuqgvuG7wADS1uhT9lmiCoSSzqzxP4xdx+P3DWfj502g7
Vj6qm2jXmsAefZrRCwZuOyVRyCHKiYUwMsqXtgG2T1NLri159pPlhdJn0K5GyIfO06/zMGuT/3kM
ysOPsHmTiLtx8y/+m7v1sicF8i1UYwwHNDpW/EWTPQkpV1xeKY3y57sXKRBJy1AEtW3PKtJz9XpO
Mb4q6h6x3P9sKMolSrDh6HgLPSmnR7nGqz3Vujxq2A86yRVt6l45+Wm0rDtzD+20P6AKsJQNW/pi
76JjFziTrPYcnfaGVakaR4GrBEeNxBVgyMU9oXrMtCUjLOd3Odk2DtErPG22kGz9/U0nswjY4lP6
nD4ibEv7Yfb8vdnITh2yQnIwY4Xs/Y9QnlXb40CHQpLxgAJCHC5PFQoR0Y9kBjR2iT7ODH1R3xE1
BzxnumMX+Ly0wa+aPhm6oWoIjyleQqoVlTfm/UlMN2ZWtuqTX+poCIJk4Fvj47b15KOfnUt53R34
w3Juu6fD1hyEkr0vALAFq+Vq01SPOb4WwfBXe39g3sJucNn7a81A/dAGOcjy2X6Zez9Rn/UsEd2D
eGpPorRbez0Z3A2B9kcuEo7JSBOZqNi4FVHU3cFYJ/env1Z5f9rqSHzgafeNXps5fuESXlQ2S6PZ
v6/hB1/ZJqu8+2adJ+NtiaLLrT+VZMFBPjLXLXRqLzNSC64FBVPAIp63xYMnQ+cBvh4d85SN5PVk
lQRP5qO9Uqp25xLwlDBbaiOCPtC+0HMueEA3jrrYJmIuJbfx0hd+Znoxdv41SLUUUrDRjF5Q2VCV
Nn+ny8eicSisQHtG+OzEd5Wte5nE2wgj/7TYFNEMPEwT65bzSB9rO+XQJ/o+bgi/D7Mm7YxmxLMY
NAQz/dOYsc9pfAchvH8qFeig5vgHKtGDvcvdW0N0mbCBnNaSPshruA9MKh9AOmP3Erp5aX22mn7u
7ecABj+niY2RK5oTV/GtapwNXDuSMiPyChVUbEvusQ8RG7mS8IpXSpS69plMz8TV13cAJX56qt+l
is0MO69g+LLFYyp8OvaOt8P4h+ItkruGXdNzNTvucXysyI9ep5EO0ZdkloSYUUFrS0jqfbVffQfk
itDXcVmpGHD3p74E24yP+9jC5rjahS+eER5PSG7893q+VAAiMP0iB0PejVCf5DKaKb6RLyY6qCBA
IvsGUkiu2TJj/sa9DpAhdnc50OR/QIF8IXTGKsxxuda0pKWBL2aWrrFhYc01DJjGMk4RNCisCE6O
6UuW6HedA9MZMl47DhE0S+U4Kh0A1dCfLn72FEu3tAYcDXW8v9CjTDFuw1Gu5u/YCchBwVfeCfKQ
x9dlj5TPzMx30XiuKqh3zSOh9Y8veA6razdc6JYBVqPf7asPczzanqvRg8oOJ1v1PJScrAFLXHKy
ly/DaIPfJ+cUu/FycMKq10XcpZPG/JpE3kZMrLg79Ec0o64s0BE6voj/7hLRMeZFqSAfK6Un49sI
JLDMatzei4xIGPQ9OvRhUVJdfSSvhh/FSfvadJ/OPmbZy7XI4/Z8ZlU6uwlV2ZhN63ItX0iSIWDe
uu8d1n9tFoVVV319UQGBVAnAmRbnySNDZGxHs4DEpmDRwHg6LAvqSsKyMhct7CVTCLSS0OC0nNub
SgtRlmsW/V4w66T2tyNpMJSSvbECEVBgz/r3hfieqvKaufr3T2uPbBVvMEbtDnRmmTNeaPa8o65N
DKfv8duuE6+CqKTQ5kYUfVQ3HpM8G1MLSDI2qW7BmluG1g1qjIL/DGj1VqDX9KDj+iLv3+5MA3Cp
9Hh1+8xXilbOQpMAA4tjeTD5N86s87z2IODXpmaPLoZgdXGEToWG2gIwUGvoTRShN6/umXtp9pOW
y+y3d9ZJ3T5GA8t0OLnCSoxlmoHQF8vWX4iotPb7GQ2xQGThMpB7WoOSOvQOfqVr0xJogM72x3Iw
52XmQefl9bWC4zmcJxRJgRwZiMhauKBAaJgEtIR7GKVK9oiUStHuh+yaV6WzZwBu7sAIVKtC4ClA
N7Hrp0Zbm5EDlLm9SFup8mTtuxpoDxYWIvgK09npNwySr5L+p/6oBe+edIom4Ea60rDWqINt2n/o
lopKBYmuv1vbhEXivdgex1FBS89/Bub66FY2wEw1IEw4aEOWDztDHutem1k7PE9M7iqQqr6cqXe8
iEQojmeM5qrFCwu8H6AXKfo/6AoWpnZbuve+Ca1Coy6+2SMmSQmj3SW2adr/qw0uKZ/wtlul+lfP
G61eWhe0fekuL01OKz9pfYPf+A5gUG/M24xHGoPjhYyI5GE0iEA1JyWRsEG5PoHo42Zbweh91Vx9
yADlMZaUdb2TDGHPrvX+pwP7gIKd9EFqkzd024QFMKko4FIi+/Q5NJM7Dk99YeGxojS6nnlvBFpf
i6npXhR4oXWioxfBqvS8hyzD8fclJ8mK/AizDY8JIeCpZGQiAGle2B3VQ/RRPwwGe5tiXpRuchQT
YxjeHXzACgp9lAQ5v2g8HgHuN+zi0oFByfM6MNjTbGl9xcL0dgBAAmgY6j1DecpLqhrt2EbsYlpC
fGDq+itBfnQtgtih8edKgHmOhbVET1xgQcw1LJWeV5IPB0IcLgsR0Z1VenRemfZnNunoYtwVMdyM
txeIqjbLTQEeIYL6SxmKS1TNG7EMxguevcxLWUgLHod2KqzU6ExeK3/oFh3h8CbMKSYG5ueCY4JL
rvK0phR2/egMcMZUHzoSIfr7cxlxOT8ir0FXl3+PeEz2cK049JerXppaJePUru6OcmUC49vNOcT1
XkeqvTVxkLQRPrf00zKAeolErZfnC/DL7zcIy4U1nSou57Ol7UP8Mxdh4T53a9XtYbKNIsb3HyWg
/YvWmBMCdyyHsa1ISwVmjbChMh4R1Aza6vfX8cHQuA0qOzDkgBShBPslBybpPg6iL5zL6SXZMcVr
BmqyYpeH+lmcfK3ZyVuhLaZrkhXPwwqNQK96xup/fvUMPrRdXubFdNwrHUpUgJG2IP0CCM8Se1Lw
QgeiY+xWZrkzBc6U3x33LGm3+6hjTousdkQpYrYIZSlSAzLgrLBQ8XtWmZ0fAcjjpBnF7MxoojZx
jctMYcxu/cUDbmI/xmznaonbCao7pcE/dQ4zE0R4d1a9QUPclvvXorNsSvgfni7aaGR0cfSfJxi2
3UMdiJ9lU6qsG3QDyqZDcMv7pxmHQQvLBr9mB28uHewLsRRS++7cbcrQkrZjc7U2/dLYpjbtq2s0
2Nveek2GQTG9RJHNoEpnhdbux5rxCQFXdz2f02ulPS6nVUS0vsAm+QnXgTuiaNxmsKYKOGP9yAVv
x049ciPN/SoWZZElitUB82M3NozHfWZe38eQfV30Yqvm/Euo86RAjtBU3qwLT5yAcRudOu1GLc4z
xC9mAsuR0/T3wSZTGE3PaDZqbGr2nL7vYbS1kG5q+vk4IBbwQfzW598cdlnjMgtTTQPYZYWKMo7D
ayDsotAGc0shEQeE15QrwV69z7ek42BwL+2gKuGifuPUpJXmUC4MPZ9FXitzAmP6RKksIjyMTnzU
4yFteRsZRG1xDTX1oD40ugDRUaqEWOG1l2y0wtrDFgc9dRV5B/gy0IrLU+BJOrfvIX+wiAHhV3KR
nQxv/tE3pzIJ09kh6T4sqa3S81IfoFFs7311b48dvTyTUDo4yf4n3EvDVEFa3z+jOOKmmOUgRPcm
dFig6QoSj6SZOeFKhQKXqnUHe3tZrVETaZzhcb2HZCr1M3sBPs+froydFRIc0IwwyI7+2IYdJMS1
P+wrsCDFwpU+aWaetuXYZG2AaFt5/p/AKO0hL8JbzhTyj5ZAki/wPLY0rRSYsDrTWQ2X49v9o1k3
Ih7t1selslsFZfI+q91rcdaQ8P98EDucVTr5689Vhi25klEnamanUY7f1Yo9SS5/MLx52KEWrf+/
wtLeMn26evlTiXkWPZ3QCHlODz96laObFyIfn9XTlUzaGJK1+14b6j1aPYYgGtRk6G+rgcCjRcaj
EVJB+SxbBBxNKBp853ndi0v4bxuX3GojvIlX3oOWO81cKJKVaqsC3yWKJk//Qgh27CRoYzl+rzL1
TRuIwZOc8XkR++qXRsaj4RtfP48xIiy9vl2j4wPaazUSRRJlDD5bZHkB8fRuRDNbaimtByLGFUJm
S7j3xXTMUss7qJ/tTz5M0O035/iBYkQFc0+/GXpAG7epBqWQFw4xqGON+qjNSPdLzCuyUhngA150
LHTFbcNvRoTUSQAkwnZweeg/jvhG1EkUkt079EXSud2fG13MSJGE/XR7iOu7tw3H5nvvSPWVIFo2
VppH4zVzRV2zJ2NJVAvQWl1RxOaXBgKK8jMNMc6gjmAkJUDEQ3ComCS4eaGj8zwjJDgjfz6bnHDj
ayUaE34UyejBIWn4/CqPdroGa2aFbC7/RRLRsNXMY8gF1x7YM8eCHby4meV+AG6M3vzaI1PMsrsL
jquxziQk5BpnJeIllreHqXE7VOLyiuIzMbcnWytejJyeHwmFQIemyTdBkhWIcwVFl4wvmERtu3Im
jzU46zmAzFo4qhrpOGXqQyRIRiv3+4utif0a9DCpsKcr0payA47emzdVsTwGu7co03vvtYFGfVPc
7xTtmZ55Ms+u6sxNWypdrwCnbEltuIkLL+3UPbRvrkNlfTtyGvi1bj7qjKZ5gAKWPIG+OXyn8dVa
En2zHouhXVa9ZZvHXQds3hR9qD0FJHt/reZBSnuTgZhba7gH6w71H0lY/v5rG9Q6nNmIC+SEJp6c
RWRqPGcLGfrOS2E3mjsDbD2se5PXdxOwsEGdCYJN4vn+wBuBo2Iy/3Wm2fPBwRDXDNHswNDl1bS9
YG6Hy6CO32eZ8TDJbNFIoIM1WHxXPYxpHTYziUjZP5N3AAJV6KlntkxL6vvZ9TSmbrHWDswhnMty
afGW4Y282BI0Wr4+F45J3IMDgYQkQO00YkCZKuHAQujkcf21dYYzpT33Yfz028bpyCExjZ6QFDOV
EnEnS/sVe22730n/qivLekTkX2YnXcKZE4BtshLXxP0tpp9wGlQfOMrUgeKuzE1tCTPZADpwkVsj
U93UacfWW4NSj+H+tbt0NFd0biKntVWw5PJaDruCH+29aE9gu23rFoDz1WyRBukyvh+BP6W2W0cq
FniYUO8gow0B56W96Eh38zHhFSv7MqMUWx8YQGuNCNfZ3yxo7xpyeXcmKlPVsvaUfohCCbPys9gf
ormGxI1L8dj6Mm5uA9lYiVI/PXU6JJly308rt6mO3wkr0QVz83NNuDx041UCtvmUPRuLasxxFvBB
FuKidSFnjrpYzIdV12lfeax4u0r1Tj2AWZJ2HTK6iGZnjLYeszRYuiDvXToXaoS+X1xGE/NDTzAN
J07tIovynmHbtOurKG+5sOY5rnA2f4vzhivruujnFyT4DitMUWmvLY8rbdnx9Qj0UMhBrnFNMZS+
FAUyJVLrXnQWBRkMNlxo6C298avGWIpnrLgwjK6Qk6fgJi2xsjPkWI+9xjbdmtD5O0QNi2mf78lX
5ppnsb0liMNoClymb6r9L11J7i/TT6jaxl6ExFM0//oj7j6lZ4K9tZh5lJB8ha09TbsVR4+O0Qvv
G+QMVRQ38jhpjZGOmJKEGyz0ynH+VZSqBiATvC96brmTE6bR87hOJuS5gPcdlz+TibqXg7pbAQtf
8fJa/ipa0ZtNVqHuvcgjQr9pnZj4q/c2/CPAKIloiNgPOtcbnwAvYt0hCa3FsaN+kX+yqbt0obUU
A2inNawkJHnPNpuVmSKezyQRUPRFudoHfxlav0kDLeGYiHe5Q/k/dCIByfXILOUBcZeHHTnIYOOp
MhX8Egwc6dK8HbaN1YrUyU2PUMLcG2PitCFcOZugXl/nQlkutsh/VC0TdYZXdDSDsr2lAnMgcJsL
fc1e9+7Hy+FElWwPai5ZrAznFwZYsB7zhzBFjBwn5mUPnNdyYy8nraLTEUAl6BRCNi3oEdcgpgNF
N2UTKtHA2KUjAIl39mVv/HpKxoMi+PV/5CpJKttfptP0DwFB+cKFOvdM8EVr69Dsc1CeZaGdLyL/
y3z0ndp/PlMd73D4Pgk+Dg5n81Sx/3NJI/ZM5XVCKWliO6eJyFqfx53C41ZGUEEgKjQ76fw3v5bR
ycLGc4c2l71Amk6RBaKNMYiZiHTJ8df9Nm7MnvXlQPd4+qYqjGwFgUtw3jagJclSpaJL2sfOTzKZ
7mFxZdhvdSlfR0iccPt3mWvNwHugXrNA+MHPIehlzg90nBngNkrBQj4ZXIKk95AKjaUncBlYmYMQ
ai/l26Fi5Q5No3zXdkaQMu0KrvL8lvopIXgOZ3OHyAOrobeYn6SpsFto0ikrs4+pwNIREvRrdcrj
UFQOWAhkDo2gX4Uo8s/ykWau1r0k/FPEMsNklKUFNCrmYOQ1QsAeMnYGPYGCEoaGijmIa5MRVHFS
3Hr5Pvf9pG+fYIB68afMWrzDPxodhffRc/m8g9KnsywhztamW0jJGHWViuLmP4fQMHSLGCWr+6x+
9W3n+y0owfajZCQcnDMsmikBC3BkL35RtMzZd2sAWWfCJPX655hFhEdA92yfOwAntPCbHZ/av+6m
fI73t9ugyA+mgkw1zpMF5azw15jt6BhPHEeChsm1T1gEskKc77TKY0/dMs6iFUCA2kf4OmaMmzcw
LKaxccvEKYBLbdJGZNU0h7SkqL3t6Wsh41w/vIhklaOsK17MidSNoFwZFpgFFodELsGH6CzRiYdI
rQbuMl8MKcU6U4xQXk0eIFodN9L500E5apWMbcBYGVHdpSrp3B5zlVSBhY6s2AYkAGruDsL7Z6D8
3oZWDFvmDY1oC9GgZdTUzoEgY5hGMfFzryQHxo4VLIS42BdEpJX2WNYfqD4Qo+2Fh3nrfVF1KjFI
n6BU/DHcHKxiywQjgNjH5ggUu1T0omBSbwaDZ3vtM6evHtWZAqauILeaJIMIYFEqwhS/WafCOpM+
qwcYtgHJa32kIUXq+ZVrfBW976mkOcpUh0JaicuGXdZ5RoDm9pdBfy4TpXPemwEow+AFsLWxrQOz
cEbX5MtGa7djQK+Y1oqh1eADphEJHWCUSfWcoRBszwJsI6P3VmurDtKM09z+kh+5aEOtKtm8w98I
xm891ecrjXGaBqnu91iIyCQRvLndJvrbokKmV/yDRKVaDBhWuWqjafTbC0qDjgSpiZVMtKIt9q5W
H4AVCBL5s6lin+GwRscpTsyDQj171aC760p+1Soek8fGOJfme2ZMn0jXfrfxu+YuXubmXsZ6T1QX
kmxPXlqJz0Db990saz/UyXJFf0juJ4gsr7OZ2ogIbnThB8zyLUAedAoDFNspSrTs1YRSec7qxdl4
pzJKiyNJpl0bCc3d09oxlYbHUUAPaEcVHmI3wB0uB9AahcRQwLg/KwgPsQPxobyb2DNPZXPqiCOR
m+gPeKBlOmLcAcFVOmn1RW4yNzNP/GyQLPB5s8kS+F2skumebUOIY+hecB3ea4swV1elg3ZhvL7V
P8rth63GfDv7CDN2kcUCZcleneMeeEcAQRlwC9qtozLj/Udnk+OgddayZfkMSfbwqkdKzCLK2m/b
r0VjjweuaCOVnvx7BzHciUMSpFL3dglaBH69HmVNR6NWQYmhoen5GRHpbChR4/lO1M97qqcIR8ce
3DQKX4EBvoDsenVQmjgsVMleBA0qsdZAoBpwHu6/5TNSs5FgT91gDOuDYSE2YY9nYvgHx25NDlY3
g5SNWdzr2Km8LmWSy4r67b/bg00C8Vq3XkScqmHz7M9ttzF4pi7qM/8Pb2uFgf3MxySQ0mOhFant
d08djQWHe9QLwuoPFR5oY4ls8ITuoRcyOySJmbfq1NFp1IQ+pbNG7gBHCCzPKHh9iV9z++LbE37U
FzfzZqdkbwb7awwFSNG1bHRwmWZy14SUG+O/vQd3YnwLSeu8fITjkGaHFC74qSaCz/DNZEM5DW9U
WWHubpvfuLD3gnCSm7VqaFTodG4KJ6gOHlTsdPULukWKZaDhAUglCoT0wIlex7gb8UP+GWOzrYXV
oELeQUpuRqKpsxkvrDDLAydEjldwar6DspjAjV8tZ2g/6n5cterYNreQ80iW26WYQi3X6AzV0wZu
Oat4lp0YEf3kgLH8ubX5hQQsLt4iUFWgY8mzfWbgrDp6N1gofdIcLYodKiKyDWVm59Hf+6VnOWRR
QLR+iMSKBBthsVvHQjA6zPEfxtZJTkCtrFThnW+vy+Z2cFsXHRL0miTI1Nh2nSN8XlpTJmBr5OlT
JD9DfKO7Vuw7Fp6RI0xGCPw5dZwfbRafcLCKIHp22010SmiKPp2lFTLfqHPZjMFE6SkPg9FSY4Fi
AutFGTQH0/dyAYvWuwwWU22eITlvXKHtOyJeZzuQGmCEMTtEuzqv3hQumQNs7o1lXwA5gGkY+brQ
hswL/4eoJG++tir2zYlir7HnlE61nuV9+vR0lvyROGHW5loylBVglMRJ2hY7iJuS5BfW8QanZfSl
GdC7a535laZQ1Bw7TZ4ZvuKfl2wMSw1Z8r9h7g4Rhi3Fwc5jnZXB4UErae3L+30WRlq8sVTZ6tcZ
BGg4mm7OdPiQ9hk0caSi1eYwwHgXCjAoS7mH47HfW5ZSTC1GOL9SLi4hl/IMqPToxUaB1a5ywKRc
0M4VI7ZYlbgfIjoXNmdHnR2uKz+DOxnduq2X6UihSDdDeP1jmF4WUAs/E5HzJdlgLoYJ4cnzOjc1
9Cb5V/Mzn7Nu2B9QuVgnk7+RZpwZz0ElAp7CqXwEMlcohOHbUAZNs+zEwCAobyWHNf044WSuCkoT
v5HbhQdKDYdOMqjM7GStVHH1PPy+Acbo2nW1hwTo/xAHzdU8VjUxkKN9FxIs4Pv7a5tPioO2RXp9
QaIazt9Wh9VAMr7Nk5KN607BOMR8N9FB5ksr+CqMI4NSC9MVK1Q7QtgZNPg8WtjRUfhS1rU3xFct
42KUXNmQnRX65UcE2Q/rzJb2lJzxLvPzu7aNF+pI+8PY/jEDrG79wD0wvuVJVizr8MJSmVj35HMA
9KuuQgWleu59FIm1Oyh1xEX1r6Bz/M3vTwP3nN0PMupSyyQCsMPJ00wX9x99lwmA60ngyvoCiZoF
BPJWIhK7vLvDStAlPbFsCkVu6hNG4HW2+xcGA5X0pvtCFKR/tVDxiE/UOHLWpN70l3CtjdPfvXfX
+lAJpMNGXBUfWAn/xkhnxsA9i3ceDR2p0odOXCEkVvSSh122iRj8fagkxyZB+L0qXBmtHADByrOc
+Nue+OIHFeOqNPzKe7iDJdzdXZRplQpENGApCc3o3z+/d5ZlRBYVsCDFPjRy/EuTJ8eg5FLamDIg
Jx3lPL+FMwW7wbPt2aDVUSPBQPdNWpP5GtgSyWa8aisfyEwPUS1fdtkwPx3vgrwuWvniTJYGhFLx
PeJf+F84yLa/SPCeodDh9L2K2kWNaTo7keYkou/MDOgr16/3Uw33A73qm+7kamIQ51QeB9fUp6Pv
qAdra7AZOTkVVsqS3H101E18QKf5xegLXAUxN4kS1Vg/XktMPbQFnaArXAn/u98lQQ2rwY8VhXrZ
e+rEQGz39TZ8l2vq/EXZsBkaoJ4XilInFXDEz3L+Z3JKZb8O5ZP8eAZYnAt+kjL/IN/Un35oy+vx
brFwDcmtIZbLnnNcvuUxPz4dionqBYQLU+Uzy2XWsf+WVTmY7NFkbphussnBrik9+P5qT9cw7ENA
DLVFOKju0pX1ZBspPYv53mkF6A+rVOHXaAqTv/wJNI715i6Umy0eKgzE8CnEvXsgG6kblpEp1CrS
LaLmkZa2EMiKfEkIgC1gjelJ25HVQ3k+90+UupQL+RUn86FALlzx3q70vKaGMRVHi8kBacHklib7
B/umhY2JU7mT/E6AGP7P3ayXggjcbMFq2QQMO1hq1fTNGOcNdNNIVQjiwhkglmRv6bJz7pr0tQeS
3XhlDQ152KFKptH3EpuDR1dAuh9Qf1i4d+gpTynzTPiqs0CML24aX84h8xMIEbsKxLOsdEqQOOno
SA88G4job1mSIandeWasc5CAZcLqtYzOYUgrRwDS08h7nl512Ntubj0Kl8edzA36XMweGiFUn0AJ
/KDu2OBblVZWA+03otdHrso2/lHmPGbhgdW7EyWeVPLBIjKBylDob3i0HqRizcpp7Yg0kRv+Chls
QVkDtork2hrumEdVqOHVIxJyy6tH3/U4bDPYkTMaHDMtfr0b9ui1YJFtGM9n21XJjMBwhqTYDYun
TkxIRb/ANmdyZwhovwTu4n7kBmO7rNzVx57Bg+yIzHOv+13GhkZ7rhv959x9tih7xS7luNHihWEm
8y3rWif20jZXsrs+xLqrd6JPQlzh1jveHEhlH0W/BHJ3jph82N9jFXFtF+wPJvQ6/+7T3/UfoSEI
iZQ/E8THhtA1vSZEN7iuow9tnflyl0DEkziSJnHWso0i+h5eXuyAODZPSpbXDrNKB6Yguj/q7L86
Qk4slAKsoP5ZuvD+RgFRGFi+3nWNhJXq/jbCMToDGw9tHiQ59C+PWs/UOcrGJ+HXveoyaz5IzWkI
zZk6Sklvf1NZansbdcNPuQLGqjcUEwpgy7wlrFJpIPBpM/jNybWZkzayO9plrT8Vymn2HRVp0DCz
WSLnDV4TOuQ0ZdwIQrmv7dBCGIHtATlU6FXrEl+y84A7zeTf97d1+/NPoJzW9AnHRgjOA85YNqIZ
QvxjimWLGUi3YJEsPegMYkdTk7DfPpsiXALJHiZfRXEm8u1Hj+Pq0bfqka6EnNKkpUxo79sNnIdy
THlLK3bsjJnjziuaBFe9N7LrcHcBKnkKGhOOhd2wtjAGdwS8Y27fXRCzeYckaxsUb49DznDu1OPo
R0tcKvEqFH/COkdC+3Fh+FvoI/oexRev25xhDX5UZ3ytd2smBJayhUXz97BCcJdnL9hupxXpvITs
Du6kCr6R34p/ig1GVxNtLCw20fBnIZ3j08yxvnKLEIz9xw7eUBaTG7IldH1XTNH/La4kyOBVht7o
kxjh7q+D+LfZVuXGKdS1xDJ5C9kqgPY2CpV6rejX7TWN1Th1dkB+41DCStLjN7hU3C0UUzVVuWWK
EEBi0VRiPjIG510B/wG0DTmlm+R56Me5jSYi1b22L2iMrXh2sFhPZZbEWUkPj5YjGL206yh02xtH
DzpgchgTEqUKbdsuzRXY1uhL3ka/zkGyLfxCSJZDMIVxnqzBVaZ/jYrHynQsooHrZXzcLi4J983P
HyJ44S8jbvh/jiYBX4WSSe+h8zSRstcdv/0EPOYZpv2iVTNT7QHA4rbboCgQzlokwP9ujk2dNVp+
RgP+zhvwLuDc5KO2j//1992yghg+tVoUM0RupPVfB1N2g7J7zq6vtU+Iwg8yPz72Mr6Ow3N25voX
J3CGL+T1hc8E33GrfJ+YjTomg3jUcpSt5XudvPvYGUx7WYYwhRil/covdHHpNNqBg0bg7mFfZAkB
TF0H5Ee8/5FacXrLY8baRhJ8DtkmwdfPWakBg24w1myqjpYm3y4THD/b5MbIUZAlA+D9NS5spJA5
b2gyqeh59G4zXSJw2kbyRps+FpvkCrTHGDb7zEzRFEBNxUAz8G7BSHURVmwvI1wgye+oFd4Z1wnB
eL1jjlz43LM89I89zcmxBTIV9t/FRg/nCCFm2EWtaivOp+lH9HcKHHLwISepBfgMdWqrzeitMrMl
TMLkdFceAujba8gc9m2OMmmbk8Tbf5CokLH+iZdyKh1WCj3CisFQHTsNp7adelkt+6W+G2XuDc0L
oEAgbieWeDes4Fbu0Jucv+rQA+Aot1oODcgUeCGU3nFdSXM1ydOuKdg01Q94GNq74v1jE320q+OW
kklwE/xV3OPhSU+0HVK2jZolqSBekXioikrgnTnRVJcjPz24VXpeSI4oxYjnPm2VD+ILnw7Cskd1
QkXkWbqPyVkaAcxd1Jzmtu0s6zaNvAUmQrNgHX71XsiJl0swAR0vBP9wDJ8C5+wBA/EINxOtAmWh
jIjvla3zuRZR+QEe7u8RLgUfDWL1yn9eqt9CEz6YZXnnspF8yHWLTOtq+cGYYlfmyh3qmp1dJtCQ
ZEkqrQezGpbSBCGsWqiXBN/ziQEsGwQJnyITqWBgClG/xMXTBthupAqzm0YL9BYurxatYl6Be+HJ
91NsfDL7tjJ4/izgBlR6m3FkZ0iWNJiokOSrBo5VP1HnaWGQ6wX7mf0UKp1Po+n2Mn0eABKxBeCy
rluu0JopokTfLLtZVLDA1XgGI5K0BpU2OY4M8HXWweyVtqEc9EQ+UcDqeHJdy96JdfsGwnja/z5B
C5XIwKINMLPU75G07cTkejtdG0vKAPffWtixfCtJwdKUh5ebr+M1JvHaypsoIxn9eQLUdWaIJwn6
axbMLofzzslvUskaSUoqBbQoholQb74rLDuk2tzxolUT4/9HEQqAU4EZtBIvk4qg0UOq6q9TbMZ6
j09KIHl5QV0Bm/XhbwxPcZ83KqeNI20tuNt8H04aStLvWynpJQGzFUCns8z74aTfhMfT1w6xojyS
MCotcWGmC06CIi9v5YOp7CU6ft1uJ/z8gghvTlBbDkPj1VsNkQP0FF/8vtnHN2T9a5CTVPx5sweV
a7vZ/MW94hvMED8hgUtaNTSbcmF5zMwp39ku8yUwqfXIxBSXAIXM0SY2dH5yrpbF9USzxH0tIZa4
mVBeFf8MFTnSru46ZOL92fsCIKqxehnD+B5lbMBzC5fMqw59Ug+9reQBvudZJ//4rgCQvQgBip8o
Oiy0i1URp6VW2MCo09nAPE0ltR15tLQWZqSRIDQC2Q8K69cDwSjXwWdiyAPdGes6+pzggaGmeXrf
4O5Ccel8C+lziP2gBjtaFfy9YbsXKlAFTZ06DYBVofoz3HtheUy25pcB6PGDW6fZmaG+ZWnSl6u+
dI8tueW9MW1qbocFDIEZrfjWGxq67p+u+UDwILsIq8tILxWb5VPhuLlQVhphY4BJ4uifOqwiFt+3
zi59/8wxsg8XYmWrdfo1BofIRU7OyReSh7jmICTtomHgA7PAGGk6Ald65B6S7eUjZLXNL6K7ASit
gIowweTXqQN2eUbh4keQZBI6/5CP8i4eoxVElCTrXYOdpY7pAGkvhOrd63GWgWZrzwRZBn/Wt9Vg
5nVcEHCF9GYcOGoLjYvgqwEdH0tiNeEIABkisbYjacRlDhhd8PPqP26eC3krj9As6geiArf+QZyY
YidYdiMLzJ34tuQS4Sys4//r27ZfYIZLLe6tX4dHtifnmp/7M2WaKwYptYd8CK8NVFllaVQREIk/
rdwRr66rZrEfHTcbUyuGmyk+FMHgbw6To9WHaVOeYsXW1DiGBVNGPLeAM2JV+UMXJSMKIYFRaiJ9
Ptw7HRUaB2s5uwWR9qjaWIbBmTvPmI+UDDnyg66yIHpmiWLHSsLa4jwc5rlHwrXpfADSQD0FUvYA
iQh3KalcZzgdMPYeJQKnEnaHxXHo1StcTHZDcbVa3gj3+8pkOwaUYiPiR7L0YuwN4GrTaakDkXxV
wMcLk1hYLY96ibgnuIAuTcMeJ+iMTZh/CmSYwlUIY+pJylaZlBeu6Mpd8IU+qlDdXDNux4d8SMCK
cUtdai8vdYT2XK+JOf2DsmJFTc+UuBILnhri3czgKJafOtoRO/WFWZ5gvbib5l2g+QG/CH4cFDzY
OQZykWUd/vjhGfIq8zTAZjRQeUvEsyU3+E4DfP7ebYHJYFtPyhO+lHZxT/eI8XttQX5STHXKXmPf
XqFuf+anV3qIlCgL8jCLkfaT+Y64/I+GgTMIFh8xZVRitsNSrOXthUik/D5ZJta/5O/gCpOgxAEL
HPKZ9A8FSySmxnTBT8Ows22JpN/W01VOWf2Ux76C2vg03/lLlXG/5yz4eiHYCUnPfuTsm/oRkv5D
3KIudx2eYVereT/Fi+qn4gvfZLe7d8gEDQX85H4pEZR/qqxlYLL7sXh2TsD8MLgDtkU48Hem4ppR
enixy/5h1xXJNatKHwof0E7W9YLEHQ1YZbKAetXqTLXeL9HGlbm8abzasoITd+jvBrdkF/3pyXS0
O1TpUnFIXyC2g6ay6waK8IQEeAP5q4Pg7IxrQNYSeQo7cGTSthHZnhd7ZYRGMV9tAutj2wmYUCBX
Di/Ez4mggySmMcmzWI/TTGnhu8BpH6tBC2SrWTOh9QsyP7kVhgZrAOrf77lR9BZrAwWb4A4PqGyI
pRAVhGYE6r62BKzD4qjrO0hFtU1V3664OkemVWqhETFn38KIdU1dMRSPirewDPs+cOKfwFzGomk6
uJ2Y56zTyqqalHsRyyqbGNCIan+VscEG3FO8Xjt1fhpMW/35bOsbytIUknI56KM+8oqqKS06YfLh
QXZT3OvZIBKqXKq2MejjnVgldkbv95zJvoF+jzjnN3qrY8XRRBi6ayXrnxIiUPFxDcOqvo+TQCkP
VYo0P17HN0zT80qNfvpYeIn09PQOGPOAzFGBJR0QO9SaVJToghLEOJ/LHA9HPHrM7qz5+bMkqyM4
QSOXxWvO1C5Z0j9atuCuxa5dcNcwN1FlH1KiGIyssvd0It76GGRdjXduMI8HjYaftxKx8b+7TGWI
y0fH2+/xSeuhadI3+UwlI313SMOaSwbbza/zum76V+Bqr5xjt5N04qZjR8g+FxtlLiCsxLJdFXFV
cPr6anvlMEFnpHC916BDvJk7VNAFdmrwXtGK45BTjOSvozToxEU/C9q9pIjMcaYj6+2rk8XDQJ9L
AKBdk9xwUMCsgbeSLiQFVbFA75mj7vu0f9+PcJIg1Yk0lxOvpPGtwnzjA2cFroiyNz5EsNgZNc+t
vNW+b3JBxHq84zDqoHIB63EsAPz6snQ10qunUOlWPeGDwb6k+X/g1bvOgsCrtLKGtVTlV8q6GhjA
uQlgW6XhmaJUJxu7DmkDBaPaorxqAYVyVVz4FfE694c1otkO0pO4JBnX3zXwnoUOnooETuFpDH7E
ZrVocM6DS8IhcUtMtMXZbK6f7PFMnShivNP0cgW733+pC4PaB2NbrOyqPEWY90Skt52Pf4xNEcZb
+slrfu8loJKDyLJIuFk48VOyEpYf5wx6D5R9ELlTGGyAfe4r5kjZ9d0qTYNCjSwIQuET6PQLZkAP
NI1jF8Rs038tnHVL/99Df9gHdQl4d+Hfn7F5o8F6e6EvN2BLwA8dHUl15CkR9l5FEkKi7VDqxI4r
fPuIde4qIRnkDiFnP1VhyA1fqmU0+RKEMzikxmAPmv6LnrdB4B6lF1PQ8JK7baNP5kx9XheI5ckH
XTa5mnA7o82q2U3q5bJu6qgmeAuqD+k3IfSDeoQJxpeTMtFntHwtftAQEaHT9yOH92PBKRzcQj4t
Ta4pqICBrJrhTkErtKj3ynFFkwXN6LquW1SEAwvusxwYB5D+uxn7ZcaHjPU8saaqvym43l1UMzRy
/3B54FwOtF8HXUSxIpR1JmyxGH5eZb/e8o661vxf61TAsKQ55XYM0iU+QEJSK6pO1JIhhov9AQbz
uu3/XLI3AA3Lj02zJWOrvaFGyEwbXB66RfI88SXN5OaMM0JPvTmE2raeY7GIN4FePCKcBEC/caL2
fWsxPcu0vrwgL8x90F3Eo475qw8HfGym0N2dzggy3DroPTxSF62c+XhUmFABf3V+ecDkE5BGryMd
Dy5D0pS/UrLvY1Ht45vy12P9lgutif8XZgbZKqCuvIVaKGiEuCjXIqve/ByTACoN4tMNIoxGqxXD
O7IB46nmFI2vTyldTfa1XwIe7BcoRjhrS9mAxJcMvqMpUsMeyhotjXfDfltDNBH6E8d8lbtEbP3Y
By2dLYhYGe2kct88tiGayXcz6mTy+El11a2c+Jai32Wqev2f5cjzneieqg5yBLLKA2h2PeUM0hJs
wn71EzhIfCmS8wy+Btc0FTL060Jx/ZCGr6p8cVsYsL/BfdzaS8qn5pRsm/JFtnLj+iOdSnbPdtq0
EqA4/6q5IhOIRbV31rFWqGxbtAIUTk9blGJ52BG+kL5I3esXdkrYQAZMkEPb+8rX3Hv9q8xrlDBE
PcgrRqhqp1JE5HGz6qCCVagpLhNO9tHg3XIyyWXOJ4u3Upa56nyOSgOSP/TxN2ithhR3WqZieagq
BOdJq53KVPsfZaGhTU+NIZBRPfOkw50S+iI6cYM28PX3ld5LrUZFrdKozJPH/+/adc+pBFhhgxn/
fFAewabPEFezcnbHJrM6BDy8Wi/QFqMboBjstMxLjhWg7SWneY/6h/dehiaCWQ8jskKKSrz7gcwe
KPKUAuE8FdbBIeggYWw8nZP/8ssQ9EgTiEH5X38/+noHm14a/XgQ/UH1Oy0XK8W2yu+xFzeDGLoM
IeSvIPj4x84iTMA5kQ4KfngcJAV6radU+6mibqRcZ9BdCSvyztNskdOrn2DXNy9wehUp6kAoeEeT
xrqdI6n56YLVmtwD4Eag1z+lmMujI6ACR1/zVIdFL+K1NkI4c0Q6DZwXymXZ3UShubV9r8L/xFoC
/EibEGyKBt6jgZJ0I29JivbEfT799WCQzWUfvsFg87mYOTXrw+YhLb9rb0lqgiyCb3Y4Xy1AIyJ0
+idOVU9oc8EHoB8RoN/C+xuDoQln85R+fF6noTNVzKqTZuzzS20wkBiuAxD94peyf65N9ZfwQ72d
rFTFS11i0/1yabtP4eHINssp3IZbUfKurWZNVx1x0soeIpIUddTTLNSevM39g6qjAunkV1fnZGmW
MOMdrndR9I7eGxdU17aQvHDGYrkHEpmKsxQnxGYiilYe2woyj5IOyGrmnvZVAFz3zzG/6IdXujIR
R5oLNox2blOn5vMQfyehmNUU16Uo+00EvFG78lFLAydBexPdZTlF9xG/rkOLoQ9ABZ0gIXkydveb
qT/Gxss/p14eocOylLiCQrpDKhU92WAmuaahq4s+Wd3oKA1VzonRTjB1Gr9WOxJxWrgDnciV7eyV
Yd+3RHG0FlQDKFeCSUKmAIlFov1H25sQnLvBzWHS2Sj650F3eJ3YsDL8LCYHKtnP8ICa/ruS6XNC
Pr/xxKODn3oY1Ts/jfO0M/L+Ji6m0bNXSdsTPR3dHNpRV0osBCqF8I13B0Q+Uwh6Wzyed+aHYqI/
wczrVEASaivBND4ElVhDMP3gVh8l4l07G3bWjA4C4YnOex+h3CUqQGkbYbtwexG+6+6o0kX+P/9Z
kjGTV5lPnZEf7DI3mo1kb8U0pzV4CH0DqT+t/k4NUpwqiaLmyqIKEtlncCPkktNJUhOrVCY4V30y
qzL5TXHyACiFWKhXahW0LYIW5PRwtHTg5scbEgZuZ+vwkqlDCO4IHRbX57cd2TovAEYNoaL25wTa
j/5lpIFvKLArGSd6p6iGBH86k2QwPRINGLXWyg6yOwj6ehZ+VVkbxhpSjSP3HOtxhz1p48MO1mwC
mSnTOHEx8BpWb3h94/cMDpiz9/4+UME6TD5S/YtWARjrSn4hlG7PrvN0axC2LunAglnDcLa/Sga2
tlYk0prl8cqzIMjtpFPHXi6Ot7jxe1p8vWJrkkVS3BLRClKEVV67i8EPscRmZM36TlLNWO4YDiDd
R3K7gRhgrfKawqhXiRhP8QnMGWrtBW/Gt1L7WAH0ur5CKuZoVyTVZ6dKTAtVJcVerkXfvWHFcj5a
76m45xCE6O5DqLyfpd0cSlaZ1or4Tvei1DT/ni0PdwGjl0FTEL1ltn83YFs94ob9FTH7WEk+BKUo
BgSuyxmAwMrX8Hho7zm8JK11480nCvNIwoEWl4vVAcDBOGPggj+7GqQ74jlad0J/dh29HW3LvwUA
svQ9pzgUIZUA+P3NLDQw5QV/gCRTPIPa6PC5DzS0BIUoRWal9vjBEAL6qJCg9CHNKsvC75kC7A1C
IoDt1W+sZ/lhv7a/zeCYkXF4Lu4cAL7cu+MQK6b+X8QrgjnbywbRI/nHXyVPfYTHbRhTp32ty3da
0ZucDda7J87oSwa97d1X99HMgZm8TeIIWHlZHYbFc7AuJcpMqD/ze35A2Q/pXnr+KGWrbulfnSgj
enBJXo6y2+b5IpLu8QBPvAdVVFu3cMnVFK7kie3WhXly6VgZW430+pepF3MJeufz8GcLuSgh9BQp
UUPb+GA4GYtPWqrBpVUQPmeaKyVzJruYnZlsGozixP6Nr9BNptFWmmNV15uMn1tFHE5YLYv+rIxh
Gr0vhY/rl9INkNeAqJCgnzuLLUP2FeC9Qoog/r8k1UdrtP8ThS2quCHk2QXBrX8w54oV7EKrjJTV
5KOuJAb2c1S68HHaIdE81IQbM7wq/ie6GYDjHGkw0xf4NnK41sKpAplKS5AKoMJQ+0H/kZaHrohQ
eiEcdqtUiq+cKg5v93GOB9P6nXfYMCaNUofb37XltnEzz7hEovaZoXOguZrM/IFE0bXHgFGhXCIO
4McYlPdBwz0s0T1YWh+/pagNWqOFry4648cMccw5Ojl8SO6/AbnCDvSGADVXQD0VfJ63+9sDBPoY
ybSW/lbM+11ZSPdEULz9QaE6ao3MGj+bsvYa2HEk8w0952h76mhmKIoSv6aigIJFixBR0xtA9o9M
457Ncl6PSo7ffxn59Mudk0PQy3Fore8ZEVIcRDx97DfdUZDQ5bugYe8ojVN+nnZ2twUOq5VnkzSo
szf3MZI9IxMlKs3TUYzDQdEz0fQoqKLxKtmfuy9kuhIVmeEqVKZ41avIkbcZENlYuhUyedwIwvZp
iIZ7ImDTVTQUyLcrkNZks8gOyA/7dYeZi5xjF+sV0PjExEKayGu2xsuDOvgwverh6IPJZ93xtAGo
YtwmJwDnN1bxunEFvHGpOlAzxcUJG0bNLTIe5Zbf50Anyaf5Eggc7hkGQ+YS0VsbSkPJsiFIJptn
dWBur/IeYAC+qN3fUjgSqo5e7zq4enNEzdeJ7TGJ/Iv8AXnz6tiNJ6RyEsTfHg0DEzgyIWEK1yb/
WmDlaxaE10aSI1+0rFHCX2WpuGZfiu+ECoCIQe3SyFFIiqzJV97m0vVvUMlcJGJo6+0jDJvPJuqr
hpaXD25E9mTQis5aCm6aXVWWkJCuw6KS6YOPFcuDJTYn6ASFKu7zoDMokqdhS+1A+3xolhYiYSRK
7I1+o13nsqf+j7cNjYNBBS3A/y+LgJUorn4G8NcLX4okZNzGSo15ZASZbIsK+6/diDA29eiilOqI
rdokah9vQoJArOvBhL2bL/TQSxR3nmEd9aaVEJ7m5yfzu/aTMK3LwVbMdOHgJjOwejXSc2PC6CmC
rCPe7mqnyoZS/2QYg9LRB7IAxDXQwg8PFy/o1xAnqS7ohHCj+uE4wlYWswC1b3XpvRKSVsRLRkey
tXSFb2RUshXRlV3u+16BoxMNmJdfepqhvFwDFHlCh0rlnMuTHvNokqk3kZFcBMWk1MCIiH7E5WpZ
aiSl90g3/tqQT52Ap9NXsPvjztYu3KDZkfwI0ufgzkWAg1JgaSSCz1zG+G9bSQ3hSnaMYrkKVUDo
LD/0HhUfOM5Chxfz4zJxh+PJ9Pc/R1nK9WQXb/Wl2fg5UQrpZmmaJl38fldPTlSJPvsaRri1BbKf
Srl6VyP/u38DOOLG6mi8goUOZr6yJmnnqKdQJjKgB0AMuGMt1dSjr7b1pYn6aGaAOaylK7Avxj0O
0nvD4GZVZPGsDG9VrONe4nHIbCvw/cfsAfoX1LxoqLoVsZaIj0Ndpy5vKzmwyjilpErdO06Sr54M
fxQk9UwrmHM1dG+wS2gRFSK0ykD1J6BXTOusEOxkckzy78qV8lel9LZ45ORKa/EqFjLVUYBp/hJX
dMTy2jwQTtL9j4TwHq/7v594IehGMRDyTtFq1B73CrZjeex6qsGkx4R7h/2XZI1mQZeILnPD11VQ
64jhIFqlq6W8UExiQNzFN1f5QUZ7O4DYNfZIkd4VnlF/XZBOaymLOdJxIxdsMsWq2fD8YwaKnanZ
McdY4QwAuvU9ZHaaJvyry7Lydhw+j2AyHvnaZ+TqsVfYgn5vSdU6ObDYQDArliLKmyvJa0AJBhtL
I5NoqCLDuBmkGWUy3dkWwQpQs/K4EeiOKfNGnLn/DUpIXfPYdPu7HIiP0vXXid786rkgRUnKBdr5
AP134zb6m962ag8QkWu/oKSyB3ihbzSr5IsKlNOZ4MdH0qAM9BpzUrIXQfP9GVl1L2fQ7EqnHqQn
/y0yHi3f8a7BEd/YdciQfAXz97VZ4F35ULZpDmxjLIPJTr3sA5U4RlNVHY6uLWuWkvBSvQmQIdIT
ZCP7cSRGn6kfEeF5XT/odsgr/JcFNOYNegpTGaryrbVeFfWco8PRJlWGQitqGwOcNIqHQMftXtok
MZdwMlybZa16Y+NPUQzYybqSOZXBGurj5VVsvf5xrWINT/D7dGvBm1YjQmI6Mmj0oQkwz3zLRvZY
Jgmu8MBcq54GuJUIUQ2M00r1aXQNOw2pxmDU2rL+G/uwJrnPBZlqoarSlGx0de25YkZiSNLTXmkh
04unP889cZTkxg/MHfbzRCE7x71X5OWVZwFxE6YfIgN9ECaf6DXIF7KEFBaaZZIklpEd2ace2u9I
sNic5jhTeDpCtUU7RGbl3r2PfYKC+IEkS2h/VYfJfPaMTCpp+PhcmGQhVFD5gSOoTArcpYXstR0w
uVdLKK9gWLVRnmxdDuDtHDSqq4aPL4pxtgsFWK2+6ZIrBzDnR9bPh8NVLMAjaR6fj0DOJdIENgHt
t0SFhMBYFfTE6mFpywO0WLIp3115JgAX7o2Ps8ZdaolqKtrodfIjys5rCukYpDwcX46aQ/ah8tbI
e4uOpYP2L3fhEj4iMa10ktin6OeIEXcq2ftcof5pynIuoMmxBYzMTQjC0AJ9cBX3az2e7RkmfCMx
xFqLyczGjcU/VIeASq9TqBZJW//KfsCaIJmErWCGfPt2/zWvU0GG5XiIlqlGZnMUijTRPM14lMpI
x50tXaaWXDNKwRSYtswV2VUKmNZSMhUXK8rINWoRb21IxdmJhjPcz6dlEPYqXxGcbqYRTVtexQkJ
d27T4jxQhXnLwnqHZgJvAM9gv5p3A9/Gf1KNb+ltnn6tS//nTzZG1AeAw0zohwhyo9noS8vRHkPh
uw39wz84NnBqhqojpzkfTNIsAilHV/uvwtfPot/X7x6MzaV50yILRFGXMDuPHjt+QsNEeo4TBF6N
kEauYqCPOaOYb/ZyouHRVPgMZkgepWaPt1aSAYv4boWD8oDpv3VtXL55n3mqZe9aaRZml08p7pIQ
WstdjilfBAFNezAiZ2U1y9dvywEpguWk44yLr3cc4g7dURa4oFkT/cEoUDxrOE+IPNPAjH5+Y3Og
Vefx2TZpt/iW2yBzps8QVc8kfEzzVRvbmozeokzCl2l6SL1PZanYOgYbg20Zp+36bDPBYVfVdBbI
hHNPziYf2HJ9axcgtCysMqAGP9JoL5xBN7VzWFV9AtKaS5l+uqOFgxT8ciBBsBWJlqqipUQiQYgH
/7x3QZq5suoQhmaDU4vJyy1rPQKv5PtqSA7yIYbpznqcUoaeOgD4yBfqLHukyPcS7jZK5OzdVAAL
bzyZu17OHn0fUM2pwl3zWJZsqgW+2lGBXn6y1DfxCW6WzCKEcjjJ083w5XuN9H0rajIOCLAWL+Zs
r3WMkuV31Q660i9ir+jsH+aWYGiuywUjK+ohUccb2jELfcOPM4znGaai+Tq7ZcWQHRtbrEwIi/Fw
2DrRBAlYTpoizhXxMPjigSVuw0eAzucsuPdvojqQj+/G/FsJtccQk2KlEgLqDgHXgaNvlQp+2nKY
eeytJYCEGafrKIBEDIUyMqatWhtyG8/j3AeYHMZES6cCI6kUCpiJvo8I1bmZecsgfN80cskyY9k+
58F9Kl2urrO+K7hzdtiDpr6O1TGZL1X2oblOiLOc3mCgm8aK6Yjz5Q0Q5eV1amBp/JROh6NYxmBk
kMUj2VvJ5G5EkpiKBxiWC1pUgGT4mMADeVgRCB/b5IBQgnfJGABWlEINXuRyZN2P9JfqCaNteC6C
8QzyFVLA9vnzEognCB/HHIx5dsDnpBSTGVb85uVprRU28wJr0ZeezeEfgPeD0vrYekTk0lSP90uT
U2HbhsLspKRHWS73HGcPoS4Z5H5336woRGsQYutJ7Crfcxo5xgjIK1t/KwwQfHI3wCM6ZAEI0yoR
17QkVzj/vatNfCTCzrVu7mshuqUfVMAVQ46RLl15iDWOtbaPs+POhvLJhqF5wik49+kXiefG51ll
UYyRlPWOUFLaPUyUBghniEarbRjPSrEUALmG7auQdrUG22bVMHfNCo0cIGHsTm9giUKv2lDIxuG6
7fKElRAhjUMLbeowZX+k6tlQ4RkCzqEDxZLNVMvaCHCO2ycAHU54ZGXhUWkjPhbneClmKIaOiTdy
mhDWGPisA+cQOs7y+Sj5meM2ukg6iN3yFXcV11fEiDG2hPYNhzKNsc26NGkTrJzIYw2sr7+w02CB
NXG44nMuBRM4p0Amj8AIBCBfRZpaAQw5BGDZMmfOb2dAgClxuCBQHaTjq4l7EFxv7sZ2Pg/7InOr
yUTNSbmeyyF486/6I4m3uAgkm6PAdbK94RobitCSyoOjmhQumb9W5OqolgSdPehR3o7wAyb1qCJn
n+bT8F+G4kYrHxgA1bECWwcUUprBR/59QKS67GmtVUMv9x1SqFg12AryB6jPKqnbb1usA2xLnNhv
nPZ9/43ekHpcRTJ6l+AcClPRN/cA6Z0x4VkslsqIh/dDVFE4ehmyShXEmQYR2OrxLYGhfxacb6Kx
Fdm42ytTLz1K39hFs6oXv3pHphSLXnzRjzXnN1o7Y87Ps2O6127Ir9LPhdXZYg99JiXIZdn0HFdF
LSJVvSg1gA9QFANFiOgP2YLRMCCpU1xr3vmSfS80VkYXKSow/paGZkHKmNuoZZARb03mem/Z/UxB
wCHJ1WBFHqVVgt37YiM+b/wyUA7ZrlBOoFrn5BK5vtBRO6UKId3PbLGuCR2PqIZHdeKyYTyfjOVl
T1fXdcjV8YY9xlRcI0egLR6JUC72Sxf7m98D0PxnoHyWZtCbWnfFrFd97pLQnPQL9gZxhH9ARKfv
c4Cuq2RUHGfp5WcHI7S7uEtM6DalT8ILSvHcSymAX96KW4BWntn5IM4NZ41L+4NwIixLoXAFwWfF
W88N46as8BP/CfYIZQM29lHRne1obTElz3QIUIJ+u7WwH6aEwnRV9erwdXUDS4Gt7UBUmMd9o9PE
NRW37Sy/Z2pfTzzjB2o9qHSruZ9I4oGUo0YRFT1USf0dMolDq5j8zYTwR69UqYi84aiY0n3Lx4Vx
9B++yaHrtCFfWLYPY+ZoRDxlXe4B+xPl6pwjHHhLOecn2RfIMNyX0iHomQ7jcSbQKq80R4JUOCYj
zfTpRanhOkeQRRH3B40+icW3vEcxMqxFdI7NLw2eREjyfKdlMqzby2iiOP+no9r033h8oUbh/cvb
tvkB7Z6gBVrSzitQRvfSS40eFBqbR5sBW5Jdxwx/ZtuSR8PozNqe1a9+lZTzUNyyCMHvLIFykT8w
sx0vWR/g805hvae7+jwADYvfIhkhtduObEvUIkltYIVrhyZyEFryNZUD0XRUjcbRXP5uP1AbvZH2
UhSIXYV6EZatvVT7hbKPW9rl/IkjjwMq5x9h1ZtRuIHwsGh1CKCYpc3upkIaYHiRXHlbXvNVK7/+
J+2RzHbnGyrNNgS8/pTQAoz7GsbxYZ0TeK5WuQWXoxdceocweq8/2m6x0aRLW4hJeWu72LeRsuN/
2teMRK0PaOtSVKOBBvfBOmyuvh5WEHEFvF+S2ib1YDSx1Zt3tnteM2Iekb6FRocL7YVK3pZpGepf
PPq8tDU6ADTRRrR78tfproF77dJWohxuE2+5ey3odKwZ+CYK5CnjO9fayBK278n92Nm3qX8h6+/Y
lQm5KdZ9ly6WqXqNgj66HGzItjmjPuoBPMS+1o17xY4yTIipcx5Y4Ahax1G6QG43LYYgbj/Vdd13
7ra7YwRnVAXlpjqZn5oCkWxAbwhk+aW8b9lxeszX1B2TsxkXDPXw4m4Kz9YrkC53puWOOD+5PzYU
evigSklbOO4XMWUwjSwqi7owRm8HHvVq03iqzyknezF6wgxzfsKMlYA+zgkZD9uGKkqS+vhSGiFQ
LYoYgTo856OH5qIPD4MlI/FnVA7oGPLig1eE+avivYghQcvPL4Z+mtXOdSW+0lop2aTEN52IuzOD
aIymjpHJ4n7FD6GHTkdiG2V8ACtzKQNTmSCjMxnnh9Mj3z7abTLTrSi5GuPt+eXW108sQbAr2FoN
+frksWzM6lOFSROxCAxU+eAIOXUBLQ62ouIBPdCUySH8uDAyzLPy6fHZsDuj+l3/RKCVljegQX8r
eYXrqhI+PkQBS8sOzJSeUvfEHDRruu/ND+fQGnxdorDe6YVQpnByPiI4AJyq8YcIF8/sIgikGmWJ
UCYQiDhYAfhTlpNSbfYf+jpR+/0CMqqe3654gYGjoe3ZA+Y3uygN1mgBsMh4H1sYEEjZfLpEeRr+
Ybx/1YvVa3wvg30VqpxY1PTrmSAr+ww41fproYr3L55nb1ciobgAs1sbPKQUT8aVvhVMshZbeB+c
bLMBqZfNdMHUqChi1pSPTd7xG7wO3Qp9gNSqYGb6fI93JCvBMONiEFZQRpqQ1r07ZKYxEN5KErgL
zKpYopRAhGBwvG7ZXCVifwAYpIicQEMgkkE9YiEGTBNgxMKZcjBIeILA6pZuTP1i0VJBTT13ooUu
xBKBpNQ9GlqYWXwutgtuEEvDDVMJMN56hwrbgelgevoXWRrpu/Q4oREHjQIV0o1Lf10OI033ZLsh
d9CCKTq1dlgSYSfnkI04/shkUPHfQJwBZYhZDC/HR/xTJJIV3BOKtt0d0SROUFtvQHbjw1LWKUyC
TB4LBnn+SU8PwdI1ULFlTFQM9yR5lE8KWhaTbxPNcyJlTaQvfub0ufqdJfw2+/dC9mNo9xSp6dVV
RCzz7WVkuYe1ozQ7eZYISu2VMk/qepOwuxoFTx0VKccQb2H6DRZCPT6/vVer6OqOyvgmT9WYq2Gz
e9Paz0ZMD1Vet7hOfv820v/IY+ae1ebsmFWAsKADHTXS/b/eJ1HbB6yn2C49eN/ko812sjt73wdN
yO3okcFvb3gOHE0PPng9/QFzwKGpFT8DVHe62Snu+OxO8G+73hK9ls++8e4ewskJUkHYnxQtpJsn
hOOxPXdIIs0j+HqGNmWvx8z6LOM0fykTMX+eRRxZpHEC/F+StKNrUFEMKTrnwAdhsOjCCMTzvNnl
2yT4ykGYT+vqjD/CNdWDSGbQbOHpUt6bsgXqCuahzhVTNzjqKOdI7j3wBYYjKZIKVMI+YKG+0IS6
T55Yp73O+41gu/1tTgLBpiQZAVoNwQppdVnPg1QzCJVQspFgeJr1g1c8z3tcWahiKtLhTqQJo+m/
qkEZofiSktT9sXztpx5O38O+Apb9xYf4xEQrciFnHm0uzL0D6mTUg0DzjbAeYW87ZCymwZubH+Vr
tocggjaXOVq/j/B97ZYDZvMcySmtY8PdM/S+usa83AAwRyetaSdzjtius6EXAmpUZQgRCXG04YEI
twAojn6qYOfvpKKsAaB5ibQ4FzjFybErtRqj3mTCsepjpICOWig0pssSTSaBqs6744YY7IDsqv/t
9boNllMiFg++NvTylyS1gKjL0CBEVhzCN5+AIlZMIV3yEWYqgIhzfSvOP15UHNL/VTn74+0e+Lwo
kFlOhoXmnjwypdgyNs5AgK+FRB1vQWZgkxKmoWXEOe2T6RZP4GRtMKLUFo6+gffJi98QDBLyWa2g
10h1kF/tIh9ZswPlMp+sFIsvKq2VUdu9vWlKp66Bn7qgiNQD4hZdpDs24g3zm2dVfB+4SF9gCAgG
+RiExrT954/pNNBZUgmKxez2taPwQs/W9mXIiPE2WN54i/iuXdmSUjOzrLIuJjvb3BUne1m1P5X7
rWomjoThLwat5fVDouqc4tHKb2FHrsseSpNS/yf1qDvY9cqmABZFNhMRw7cr+JLzrpi96zj+ZrxK
FQp/mcC015UV3k3hDdSxGXoKWuz7ytQBFS3D70AifUdTQ1LO9MTDHRwjtGXGhR+xChUH7HcUPAsS
oM/VX4E7T7RosxkJcRStU05VQOR8ZSNdPryZjmZLQNmKKZ/lq/iSs9RWfhYEjVPjutE1whSAef3H
Z2Wc1x02vW6VT/dkYV85ceyJ2NxAIBO69D3LtAgNzYBtGQk8A0KSn3OGERxhV9mfLKPgNGMkaDqI
E1pnB5K2OAnHyHexF6kgiriejUYAOegNvgZ24cLlEMNq/qB02KE1Q8Sd7gE800TjleTurIhGsbLh
vmHoraoDm0jl0XMBntkFQIepq7bPjA/rkZExc+pY38LMP2Kwmx1kDM68HBdp5fYQPphhKKJKogto
9wTNPrhW12S6scNHAspTcpJn/vKJ4OO/3eWgEjM+/h6lauW0RFBh8NNymb0bDQ4Ici9nWjx4D88n
Rxh0pK3BAISHi8bEDY5Dx3aM2ANucBUnZB5Zlk4elNqje1kiFx7qRM38vCKvliiIPKzRDxKcXE5f
V00rgFbwDgyV6m1wyjkkOGiF3AYyHHJINrebYb+XMyvzwm7R3WfOavxRrQArIGjYGMjUP1T6dSWK
Nb6aVnWtlXDq3oT79EVE1ehwbep2gYRcsFEWJGL0t4qOs/+yR2YdYPtsnEpubbnraqffLN7YMvmu
hYZtoPMNJAeZ/sMuzmp7j4Rh+Xtm/1to8xxucn8iFr9RHfhgMHDoDsTILnMobWAhbDAP7gykeznu
J7bStYazWEyjOpgm1cmHyLe7hzE3guvsfwxc1XahKjp804jbAYeXfblbeUN0W0hrX6PRUCJ0ThGN
uqpthMOJVBBygbWr4Op7KujNM+7g6mVy0nyGG3Iw2bTAk10PS9ilyJ6IV6lITLJI5qjbKnrLw6dI
MWgoBY9omTdpKRCKBYc3XKlf8IGuPVJPW7CACHSf3xoWoBDHUgNYVnHZ3U+TS7o9ESX56ECMNP9M
v7/H3QLcWBlmSdmYKxqJt1OIAXfH9B2lhuu/s6zd/zEn/uUm/qrMNSTJMd66oF3blA9RN4qCRFmj
x8pIRR9jcQ2pqm57iyAO7jd3iBy6nvEPTmA+TOrhTALDsxvBkoXm9mFufinhaGQ7ekuCkBDNS6Mv
GZxn3GV4TNOMJmLWJOiFcMzhpWuIB31FMBGn9JjMhwVjyEFLaIwx4lphXYfJT7p7Ph5q57TLE9Vk
k6owTZcD7JFYquObSJyzZUqsdnevT4IoWkYCWxuKl5AXoeqbS5Amp4ykV3FgLCkAb2CrEvDt8D9p
cQQhVM4PeNDRjV1XdXp2ST6O61hKTFCBs6/tZrktCvUNXo9wTBGJ/WQeC/pMzqz19ox/yU1HsOgP
eP/9ac42FKwllmptT0lo+oYGLnxYQMNjNlNFv3BWW5RPpFUJ649vdFmYiD6x7oYK8oWh9gSAfXFQ
tC7izXX8Omm5UikvqXLrDpeXwc3uxr7Sd6ru+dvL4TkUJ1fz/w0SQNpOozhX9vL7ahlz1m5qH3Xd
NAtdkwgjl2VUY1MuQovDhc9pMCSAvK6I3gCV4FnHbsV4Wfct4nHkNOiF1r5kyLoX53ydmhnmPeiW
ZWxtBHiJwJYWiR21BYX6HwMIZ0TlJbs5woN0i3uew+ImN7rtAbVGSno23EcS/H9tgAuqNINqcCbU
LFJssFsQhv9ofRYw8tV+38+J/SJgDVWRBSSKYbf60OUwEiL2Qf6qe8vYbvGNMf4BQSlO4r1Qxmou
2x5XGJ0mVkjh5iwsIwBrmcphtl+3aDIdgdYGuPyi2JLFDt60C68GSkr6pDQmvOpQlCqVR//4q4nK
lkGD8PXIMx+naFOW0qGrZmPDNJHegthNQRL7Yu8cGkkB3hh26JdfJ6VlpplWexOQhMtdZaTc0rsP
Ocu/Fi3Gg5hgpJ77BRPB0UPCyHvE69cM6+/riVt3D6ihuRoDFI2Hts+cZAogJLvAefBigjTDcpQU
bcvC8CLZfL/zrovOEt4ScKDVspWuciXRxbhDuLOFkYlqbJ+mbyhln1QBVkXHlOjzSxbECA3w1S5f
TihAYKEDCp9+NrsNcScG2MDmSySbL5MZjMrlnplwNLuRPZ4y7g+NnxRD27EjG4xyTz8qzryExnDx
NcyPZ8wITWjRbEBUVi0rxH+KrLi9YfXQbP6xmWmhPCtIDx3m07KCvlg2iKsrDRkqnbJEzHIDRYXU
gEPgSYxWH37t+3+j65XRwBUu1sal5HWITZopp1cjKBIjucrWGmsDf/JJWZF5FbdKsXwT96WkN1uw
p/LpoeQKxEg8xwQecEMnSNn7fMLxfk8ebX1Pn+PR9xgAsBZVIOy4Wbs7cxr6kpefzeqMsMQrwlZ8
C6OlQRa2XcUa5NuGQWkF512yrnYf+isRqK0c4S1nU0TbV+6I5WDROnjKkOwLBlN/Ga2cAwVpWquG
vV6ZyptUU4J6lESCzEOEawfW+mFcfPZdcdJf6dnxKq/oYJVtQI2lS2qIY69snFhGOVWT/Usitnxq
V1xFPJEOtahaQqZcTDrgZkkigTfli9FEhHfgwcjxIndn6UAsCsNoSw31d9N1cLcENCei0UTXS9bm
Zbo04aCGBiiTG+Khqeuk7j0puDKot2RgTs1ChmQMscOfA1Iwl/T4Rzq85Lfn8dE6dQYfRkxruHab
nsGLr98O3MYhqcSvBOWpdyTjJNoic72dVyPceXLqqa/7Jego3QSuvx29RGQDIN/UXxlv0EMIpaQb
kKohyYIVh/noIBHZDejoIo5EbZYVxKv/+uEihfMG3MyzXku3mcXtMaO5xZb+D6Rg1hfJ861qlOi9
xzluNxXyINVedmWGt7z6J8JLFJAdW9V007+tADrHz3jzTRbG5AXFxmxy2OK9qjLNfEpOBultXdi1
4L25UFjgYbkh+6Opr9mTL9z8nsC91O0zpkAlIXawavSvomLrOtKeHaO1MqRlcYUTsSVPbD24N/eD
npDT1hIc1uC3NWwfEq0n7JKpJYY2A8NieqsZivddeZzd8TtRazpAqMAGyMU8Ot+764DojyivTfby
hq821P4J9TnmU8r9EB/bNVZndkcdDDzrE1NIXMNOJHG4tZyKb6rSw/Qj4bXeGeROcl0+KMsFoaq3
hg/EFCcE1tjiZvNYrUEw8Uamfei0m6F0ZFg1nza8RatIIeSUlT/A+sMnWlnDES7AaXcSXzd7PBwq
7fgByLQZK02E7JG5LFzclyDQM+sgKmpwyuQxNDgEIqdKBCSgUFbGs6bSkZ8YpiyKN9fcgRS+uBKX
Z7pPwb5fm80ORw56K3FVx7wWW6/9/zJtq34E7RNn68/MlY1BcMiUY5ihltcyk5D98eKso1X9VvK5
wbrFQs+f+K12nQKIgfwshyuIc/WeSd1nz1EjBn6BHV+5pFnO1cPZNVSN78qklk+dArqplaXzP61C
zuHu/FS5IeR5rdvSyNSkx5epuPi8zvl9pVteOj4cGmw0gtR6cyfAdZvNq7jfwpxFuNiHQbVT7kc+
oUGgKosdu8ZAcSyuPcFaC0tdoCNCyYaqbAzLlCnNIMJ1d+2IxEE7PSLCO0ToXZYxYsb0ist0n3qZ
fYtC2VDyaEbjU0JUVo6uyELhv3N/+djezdL9H1GvHqpUUaN/SjyScmhNKO0caGpeEt8aqqvj1jMY
Odjk5KQHX3DB72r/Nw90FjQfX7GLTvctArffvqeT4o+AXtefTeN5mPzaKo1fIuyd0xE28d18wFO8
//MtR3TM7wvLlrgmVELGXd/hrRQiSwuMuoKLQ1qPCq/rukE7KHY0VqfQZ7gPP9S/O+s4zNxRB2zB
wne4E+jBuJ18JiXPb6mCD+bcuhNRqhwgU1iU2QitTFqVWQF5AfYOawTptEbcBjpMu65XB3CNPUae
8kMe2Y/ECuiN7Ii9g3uvCz+WCRXwXBlwqGgcLgOlf4lqEgwGN0SEJx/mziwDuJ5vCLMdbYcoVNjU
qPwlIqln35ldfMl/7+ZoLZm026MgiKstakwcSJx1d94gdQ+SaX4sklF+sHFiGe2p6NRMnsXDcdXY
9WOLszYl4K9aStA+h5hx+30vqvob84Q9+6xZ5+N1aiHvc88DbFxAwN3EvQxWlXhbQm/OpL4vEYKa
JP11/AmTDWPErPo3PayW1fEFDDK9xjm71MhulWInrv3NNEeH9ivMp7CkMMSupjxYWSw9t1+c6KTY
mWdFHGyx+rXMoelhAUTIjhlUUEru850MYmg3cFQbCtJs+ZKMw2GGjDx9EpsZ1cyTvcrUvi6gpbfk
6Xhj3HGJXh+Kp/HyYSpmkngEUCvpYjxOIHFtax0jDMffrxvuxIBwI1f0YFpWHFBl6tSFGvcVvY+M
3hAzMlHz3YzTMm3FM7M+oCv7GsBNEFOPuYPgfHkA3NBmlINNm8fVEtbmtjORCfjQxC9p1eUIFmvY
jBZ+NPCYjQi/FqMY++crOIgYj3jDZ1nd3gdvrudbjABWaYp72ljo7IA23coTL0ruazFgXWxr6EYC
07dgcyYQgbUetLhf61/9h/gqh4jxjdWBm1RFHowTTpFmp3am/75H+i4r5m2nqq1F0vFY4Sf6UIxR
u79EOdy5rSjl0vM35nvjGOjIlAp7KXjEQ1xEbNZ+WsrhbMHTMzh0qQco8eO707EmGIz69CaxslLL
cKwQuKLSF1ZFk+TOEkHHyt+vYKpVDJxM16EY3ulKjje+BxY0syqWZP+bP8TMl89DDJTlCoDVzyg4
3TXh8ky7kif8Ioj43/s0it5Q/iex7Y8WFuh/LTQBUtLCBIUlWRpdHc7sqXhMNmz6fqt0Px14O1HQ
6ugdw80XljB5qj5Z2jhlqa7WGduWqu9TywychsLchi+4Udlrjn0nYDymRWbnxWu5Ii3HZg+TTPwW
GTFABYw8XrwINDISsWdHfsvw+50oglMLriMNAgwKma8NVgulX+NBq+5aJaIOSKT3I/nhtvwMnMPj
UIpiVi6ciPHqu7+/U+0lcv1ugwbQnC8QF/wKnWwqj6wjEprRdjHbMjdr+6k6Ve3A6NefuJLuKXO5
KKsoSrvoCQhp6DC668iXeZviEgTyYdxhqZuUrhWaIKl0EuZaMpKt6nl5dXN+Zd6pm4UCH8YJKmq8
ghm2sAFUk4r6F4rtFMAm0mgNYAqiKqOX+R8ZOe0pdkDR9AFtFiGe6vA9MUXqdOscVxrnUjx7GLZe
l87PAlyoR30T5I5LtfBKPpNcJ9MKb1JI9c3UOwnISDpu9LejYV6m/jetBU131jgF0JEwLFnzvPNL
E0nQXWW+vq04Fa4Zt0zeywcLLeFA2eDBzs4dzrYc1CplqX/3AyHj3hcwDfRl7i7GHbM0kEdr426R
zjcxz51+KflDlv0T8awX9bAUYEejf+n2wDaX3tQaY1fuHqeWCs33ctvi1VQFYLIkrnPJPJuY2WAg
Dbcn+2WiRmVunlbbkhkfTUFQjmmyTw9zMhO4x8FDFDa47qttJr/RrZBeDfdBCTp7OQVT9HAnnQTQ
HuIJb6fTQOe+Mw7mFOfrx5ll8aTbpcw1vxpNPl3yk2idtTwkOdppLBVqhx9gdVvJSh16Z5iQ5Eaw
rR8eYhh/2tujUEifnXVxGM0OZI8imIDT04MF+jD090ddPzM0GBQxA172hifyLXoIU06+jFXgjY+H
JWjPBRwnAGS3iHnzt/vGBIqf+KUPZxig5/ah3NkN6lFCI4ESdbt9JtpAqqli8DFR2RgyJU2AOcuM
2LM0RjnCaaoT1OfuWyF8QlYtQ+lap0ZU1ekXSXLA3FghgrrJzxd2cQ+fajUMxil1Bc5gBmio/hBY
zkXaedCkxfp3O4u81kkpx2qtj6aecb+4dqFXSwxc4ydsnpDLSNI/31ZPr2hCI42cxpr0xceSRv/a
hIlZKPThPGuT+uGfC/sKYAXCTo5Nti+5hRNvWWCVzE7wlQvAqHdldsPfsV6XvkwhCUwkP7nfd4tU
bxAgIBOHkcenqX7nLPtlDavuJpHEAk2bBBAGL5Swo/6c/4pVlmsrjAAaavdF3w9ZtJ78feTTinTe
BIxWMBiyl5dL/7LQJgXDm0NAdzkDGCbVYgKLH+5qWqDogLJDR3blC47uTpEthG1DD4C/kutrDaiJ
GBqYb6isUabAPX/V9aHgflYZDjpktxD6NwM+HHP0NoERSnwSPyHMs7E3qtuV+JL+A3iwXNP2RBkM
4bbBWSikMEzEqLGAwm8i1sQ10BkO/RjSMbZewlq/+2jLOsrYNjLdbJdjS09dYDyqkff/PiA52d20
YB5Y710qqRvh9EHOFixkMNQgqBm/5ySoSA/9mXgN1wVJy72MjS+wcoTaVC4r50ziZ7DCqJyYY8si
hQCfUBY6UqTrDINGd/KZP80jxufVbDaQRGEJ3vZF525zulmhmVTpW+MkEQz/xiCsfLpiM3USg18F
pT+uqBDA25Jslk3XwNAT2OtGFNjqZna6wnGswarrBYookqZB6Dz3m2PEvArZ0d7tBTBdfN5PA2qC
UYmKmXhfdh2pKzYYVEwat6ykq29t+xv9pK7a13OtZ7LRTgbsftzSqed3DM6honwr44Z/ETe2wST6
fBib8kCjV8pLqbthRGPoX5P2ZsDAePeYUzZQlg6w03xmazc5v+84hPLWpA/6dJMm/Itrjv23v4pZ
SfnTc+FctsGoYc43oKSF8Ze2rocl+mqsjXmnWaF3HYIS55vlKrOsGnv/92erkEIsHUJXo1O5MOFm
trnvsLl0NGdIYGkZIFLz74B77dBhf4Ri8sjDxN+getcUy6Uu38mVQiU28QCkgXcLa2pIBVuHuraM
aQiu9iGBJnSZ3nq6ssYo6/9o/yd5t4qzQ4O/yl6zOLjNvKYy8MDR+aOZpmZKpHbajZHb0Q+d/Gxk
3vJaFW/IZvuiBpfeRkb6sYBLjFagCXVREzxIOJNW30biDvpQpEbYrXE5XkpeaJ/3xLCF9ACgpLA9
jjfEiiw+PBKCWzexExu9pDk5q9NrJPUfG2NDC5zvzcpzq6Bagoa5A/CXbeYUSxNIIitcr4f9uR1V
Jaav7p4dA6MpA34jDpOJzGp9GMeShCFHUo2NSw+2OqD3WpRMXfS9P1RemxmpTnAQLW8Ebmrpl9tw
9fcgSrA5b5dxh3M8irRxu7fddnW8BOOkrR+sr+sB90JQWCiYsLnURa6BLR+HU2Mo8uE+3frSr6ix
u6FlyuqzHUEQ5Wyq4YWpXsDdMDVLsNEl+wZltgRsDK/XxZvdYVUjGMD7Ge0322eg4J33lTlNlmLs
bp/SYFYdUtGm2ixmpOmcQMvTiNi2AzFglVv6KZXNzl2RsIxl0KxUIcred2gW8YLlvafnibvtZ1T4
9leYZrvnm6ElcrkfQidPbB6X/hE4NXarCTShEJ3o4YMM94GhKFYuOQA1+cJfMqqPB2qcNIny7GLo
Q3E1XDOptipq80Ynq7dbA3bFhjn8fsgPlRgdtlXcLH5ljdtoxef+6pls4RfYyJVLJo0mBS3hhLNo
BfzOTtYh6G7yNRi+B012b1Cz2GEvOAskAVlDWNDmdJRP1+25rWuSbpqJJn9reOdWdtEqdT3VfCkg
qhyHQxKYUlXJr7nEJCfS9YU2dUJXvOGUf6bsCDS372s5tYr62F/inPbeD/JJCyT2+7CpY0ydPfkf
uAetfn2XwPuRQo4NeHX1R0LypU36QfzITo302tklvPBL723Vehx0PctlNR8L412NaxSDKah6At8F
h0dMozbJCZD9YJZ+R7nU61GltVRJyvfDkLlYOOYOko3sWSE6k0BIrljaHsPLr3p/cANNF7N9e80z
XHZ1YQDECAllvHhwnjIHr9ZF81AvUHz+5jonRZGjPs/Bnh5kD3cBJA5rjXRw7rTSBRG8Zri62JtO
IyniKLUEkcNA5UAR0AF2K1j9oG3WwOFfPewZgCmmz50jpfSHgNH8gYXPl3V7UQxtCdHvr0B6z5F/
mfmwd2gQBidor14vr9Y7d3cuaTM9A/9ZOnWiQlw6GScEjsVC5fI5rLhT26ouxeUea4yXIh0571PC
NobQy5spfLjEIs2n+gxGIpLuO2Lju8RVRV1a7uyLlNFmqf35ecLsTkJurGukbMJU3PRR/zaTZuAy
TEV6MbntZ4RVYaXQBL3dFz4PHmCfJeqlOV8y62rUUXB8dNyt4Kue4ObY4P3+TKisY98Q3P4voKcR
HCSnlRYrTorhbcu9bFe42FuQ0BVjo6zhIkDfl+6K/tH7IR0HQX3+xX5u23dFtE10b9XCvOAsnZm7
UVuUPcPVeIb7tWwlWCpnJL8v/SXcsjSMqBc4eGFVESZ1scjxHcWMDZLdyIk8K+D7EURzhDRq9yuc
fC6lX4vVqvHm7qWNQoKlYXuqEAc8vmvvQ4Mywrhio/dXu7EUcqqUaMbRAab1Bzj2YAXk/2Olobcs
yx9EO2tuojAezXm1yLbhZTPaNh8t0m6um9ehaEa6IdUqrepHOBM+gI0WuuQjB0LUSFk/dpZQUaS7
W/V6BvSPSuc/59pZUxJdK1LGsVS+qeNsvxAahal8CVYd4VkrWe71qHb1Q6zbbGYCQ+QIkwzZeIUS
QgChG9QAYMTyTix7UrMZPX4tUSjA7VcQZa+bJfJScQ41YjeDVagfO5SgMIjp+fiamC60WA+i+dEw
l/pG/Xhprxu4KNe+5F3YVpvPzwrWvkZ9bz7ITRi7E0RGxFyUyDJCflRAf0i2fkxjllKkAyZnnrXt
R2H3jr0rXXEft6hrpZOwlSYcR6q51UETcYIRNSgJzcLdU2ewh0+UhbSjAqtzJ7hqVg8jHFQy74Fj
L9E2mXEb0bd6kyArMWnSfN/2Sdlcwyt7udpa8ttoYw/GuWhhm5fpvgffJpru9VrpVgPVCMeF23fg
wibVJ+6kC97EgkBFq3WNrTuuCD4+gzHGxC4oCVySnOvB61QRfcDbtAZAKiKPGU4cDl/mx/8HnA7/
f9rbrzxE8zZtzUcCQhiRkJOLX3QMf+tD9yaZDSVgEDEM3A2oYsnrQUJZ7tAY6HVzHv/i1nm43hNR
ktVBSxaVsxlLybAA0hEm8SrF1tuZa3l1JvmhPUOhZHgEI1Q8SR57XmE14nDyS1/aKVhB4Uz+Ki8Z
vo+MH3Qg93uzUAEiQfNV8/KI6cIHE0CsjpJxVwgcQR9RU9Nz7Tuxg0i/Xmu2OYg9y4rDDQ//U1fD
J25QomPJIktBx+hd4hN5mpetQFe6onJx6AifokwpIqb8+zu0Hf262u9uu5sAysIYaPyix93DOiim
YqXLEgrfdPT0GOPNragUDUTE8bi6LsSgIWwqQcEbXURAJJmvacjHdsf6ZiLlXc6uXtOASbkoaofE
JyTazda5M9E5Ee0ilmQHuGDCfnFyaWUGXWzdOPulsraPwTjoImoShRmAH43rWBzwu0g9woUtoKxk
qafdgNufyoQqaQE5rqRWlneLkK2i8RIviWzzHiSnfDHICHfCB06JiEQCkqpH+WyQR2zPDNf5WuKg
ysgHp6L3aEqvjLQA60UoY3KljvzGyNXiGHj7HFT0Pl1dpDR9EP4TMZjQCNfyH4G1vMbpqjio7+3Y
/tGuyDv5hZP0zTI+BLQhTL8jkp5uCQkOpY5AMJ7HD2CZHf9mCUqzA5yF7ekjsMZhe9qg5zsckA7P
XTJmpC/sVAX28/+4A6RhsuXY0wMh5Ijj2yXQ9fHiwSPG92CL+UoUPdv87dUR3kBDv37yYaLyd5J4
yqq0vPLL8MXxv07kL7MRFxp/34yKQWlOHsIjfoDFnRxq8um3YhGHtqYyTroMWLV2Irj/8ecy2EN4
bQYYzfe8G8cgW94bgTwo17eHDK6GWd/2tqz3i/tVcA7Ez0/6xLP1RzytNoB/6XDo8WWr4emx4sjK
tvD8YmUfD0kMU6RrESmyjWy5sh+pP9yObEroVeRoQfBwIyLIq++omZaXpf6bHmsBtlA7QGDoNvMr
pVQHW1Oa+wUTL7ZAvd2mQHUt1nZ9GZwrcy6dXg3upacGOqK5kYS6ABEP/JOlkz70mARuhclUeNK6
JcEVWdbRNRYHvz/m1sHAs38o3CB6wFTc9YNFxgihzhkEqQ9qKlgx/kPCxBzG4+jcYW55zb+soIkU
ncDOOQzTiGbCYiFgXB992yR+nVBSaBDI3282lO3Y13Havl+5jzVIBfqxVtpGrjUn2dfRYK0VIeiO
RrFGAWyVXLtId3gpFmc3l4RW/XBUQbuOhem4sYvFyBj6Ap6zB2SltnKRUddGFCjLv4yfl6aMAIbp
Z1Px8WHQFGv9gBd83bjqKcYWKiyEBtKiTA23oo0ZJOyE9k/dWDw8s7DbRE/cxtVxT/PxBQFhE7ly
9gWcRHmJKZYeSiHofehnduKyz+344ZG0kHiNi3w9vIrcPsPJFTIr4l3yRRWPxVNyKF2s3+N1hDK/
1B2AWMLL/RzCI7nQ4ZE2Dz9xOSwatNnfndsRnVjq3UuxECmL7M77yySC4Y85vN/4yCwXDHYxJLLJ
OQQqOxXfO4FZpx/iJbftErTE0A3lIhtGByO85q2jkmqd8q+ny/9bSsZdl+1HwgTV9jYKMV18uP0Y
cLjpt5OTexIoZ8pHLqYs9yoJ5kGgwOgGxJYPH6P1m7t1Xs7GCtbpbqtQ7Vp92CHcJmeYcB8BOOef
sTdP8m68UDyNlCVMYMUYTNLnfhlrz6FOSw8ismReySUAUB8jWv55FinUmBl4JFVACeXdk/qHR8gm
Xx/InZOQ5vi2DPaPBd/sKIuRMaiXM2SzFDwxeVuJldyT9OMiKnAMY0zqcokUSRPLIz/Ovx/Ylice
TQi+xVudZtB0prfsSQDZrSDfIK6AWybmt9wcRuiL/one+px5QzDG3iu5yATFc/ZBaygQEeOp0HYV
M2lEdRGPdW3wiHj1VyJY1EYFVlCgR8u7uCX8JZcU0bdlfCUwgZ1neTXFqpARVkEjYXLPenvOlrdb
tmqgQ1rBKkeR0Y2mUyUSAxvTkNQSyaIjTlr6H6rjUMjxK4SiocPF66e9IyB1Vdq39lcZihbTQn8d
tLA8dwY7+X7YtNSHbwYlRnPh+g1gKd+Zl2MF3RB9az5EGahdXybiQomPkuAvdJWR/T3ynCJOP3Ui
prrjoZT9Z/EnCnoXN+fCBu5JHkarqDkexh4DadljhJxJrWXsclDmPO3jDCho/EBcSnTgt56eBZi9
3kHmlLa15D4CTVmErGj2gdL0ZAmNyXHZzG7ThPOXYTURPji14KHklA8rGp/5joCYvhsHQBSkM66u
BFe/wzEGw16QHxkwVD7WDn+pQwEyr6WlbGQ/ca42CkihC2T9c4lIAfGKeeSvYo4mSMKo5kvS1ghZ
MkFH+3l1Agw6BMZQ0EfGcJTeD4covp2RKY11QdaNBKWJPes1bL3IAakPvmrRGoEntLVtK4y1t5mm
Q/iVMzrZgXfFiZnpz1WiZcB5Gp6XE3uaMULzZBhtbC9iucUV6fUOyrEus6rty5YZ+K3tPDUZQy71
S4Sac4beMFiwcH3+2OTDJHfqZ5a8JbVrqlu37exngJRC1iNVdnskoj1y2Ap5boEKODtT3sUyhxAV
1TPXerZMyaS0W/xZ0QAQH9nsyvUwd4AZ7XEw4Ry9qugeWDGVyhTuK+dG8gSDH69RlP4qZWoausUV
LXy/wyv1ayCutVhjqDAD051BdXU/YWk+D2Qgkfmedbp3rs+yJOAXvq/gjX/x+qSZRsC8pbRr0ozR
fBn/O0ejWdvtmwKKv+m20mFpyp3CUX5VXJiFzQMMNQVaoBskETsCM2/fM8qQpqJxFWROJ6oENy81
zA1tydTK/7/Sm3eAkaJeR+rsUr2BscdQmnzU+vLA5mDc4N1WnvYqspIxDTh3kr16l3QgSZo4PR9k
cfRIiNdoEB9oNvn8tLfSegrAgf/x9frTA/Md3zo+wZfmblkqZpzDNEskneA/pzj9+7210OCtqx4d
y3dLZ17H1IJYeg/pAaS+8JYEhHHU84DLGbsfTh8w6wIfrIxuWnLpfhVaxY7TztylNl87k4ZpWDzL
kqFe/lgDWVVWjw/uibeHrfBepEINwVOiHH9wutFaNk1lLhwZVCTliG4ui5R7SsiJAFQoxKTf2p8R
juhjn65azFjDCvc7pvxkVlQbYHqsMKn20bp1DIsgPgt5jiRnHc3rsxzCmWRmsg18UsmopqTJ3G72
9iYl+3LZMdiaUzNTEY5BS1k6bZFt/kPMK4dRmiV6xWs+l++LF8UYXe1HUcrQL1iisut21qU3qU5/
iTz7K+Nyym4Z8loJdoCKPQM/XIsHM3tNDH3NfTBOAnl7CvmedxhyZDWan/KLjwmWY8I8Pfu60sxt
4pmB0rl6dzxiqycsRjA9Grx+VwPVoY/kd7p3y+/ubIKxnTe5QTmmuI1NYCacjQNLxVca1shcoAgE
Va4ljDXvInIzP2S909/A1+PZJCHHchvSz0R6K5raOrSOfNNDurcRD9c6/8agAbUKD5WpURKZMUnx
7FJZFSUjFYVP6Iqf7nDBre5OiMemlPbXECYQ7AMSOUTR+GFzwJfbkVY0/JFLub8s/jHrbxdHzuDB
nwJHFz/ExR8wybQ/Dm4R7UePVDN878SKMfoapWr+tL6H4VLZ/xB7ixOzv2cCEBETrBJRH6oSbc22
8aMMqaAim47NbDP530rSoMibb3NkDik0EoHoVtVIQ/8vlp+WqVIm1x7tO6Pktfh9FlIwVe85h0tj
0O21Mh6mJxxVcwc6kbAXfJZ6mRKLRJL20cFhhpjcqwsRvk2oL0Xirb0rYAG8EFFkukKcF8KJvXtC
MDOE738SMlXYUsmFiFAxyCoG2ZIIQbwKVhQ7kfbUEkY/45Eyyzd05r7oIDRqVvkJYECya5BwBWdb
fzDV95ojTLxTIjYZMfIAqjSkUg+wQN4MQz1WoAPSjZFCRndpR843v5C/XubIRohlZM6kKJpAwcyE
4VAWf5PBj6mQLXqFojuc6ov6Q2xQUUaM7Iz7JqMidV1XSQ3xruDI0b+ltZtSOKpBntD6PJA1henL
Gznk1jUzwStvHdZiupXgp+i85CusH9oRw03p0mx95xOk581I1l99Lr7JnvWbCleRCZYBM9nZODhc
86/lmpgtFcXBKU74fwCpuaPZqadN1j68ZzdeojXZSjKgXvp+AuOpJ/2nXP7dTShTpLAIVLL+6dRs
Euk5Ijk6SzV4kWYQmCsrP5lyZaPIrc8EkyrhFSrr3tihyHw2Uv7O8PjawLFdM/rueLng6VvA7Fq+
OLlPY/iXQUP/P4ypvTyJCoWB52Qv7Mkwx14lFedKwSfmYnKZE3/qMvaBBwpB59h79alYUb2deKXF
BECxauk5JQbshsyWi5GklOG3arzehegZzmLQ5RKU8rRS52vTeSr4Xqs42NVqoAG/FTdRxH70ovqt
ELJY7fKY6BMjRydiR8ccwL2sQUxHl8aYgbe4KsF+gssUHBThue/4cEw7eRTYSKapNF65EI9U0+Ld
545qkW9251UPrfMhmW1d9khogwiT2hLh8cyXDHZOggNjJqJ1Gmq/nKfpqMQrpJ14Ds3TN88TxnXg
VEBzx7i3+xUpeZr5+xevJhuIdfXconU6DEz/XhHnn6Dyd+a6my6DftT3JdZXPrCkqobYa/E+dOWa
uY0sy0s4COowMjbV3bzPejzMHbJBWqqkp22jHeUgRF7UTWNWWNoAohIzS7FtxEgFhdHLbgL/EuzA
kvJYdMfHIjQBGij5110taq+nI7db0N6cpt+3jdDRlmG2F9JaYdezynw/CRgbQl/vi6HgKlTVDzXW
MNxtzDSxyQuU+ZhBeBUFynrTWGat/iawaWxkJPcjrZnESbpvq+yVhWxfnUAYf+cCf0L5TE6Mzv4z
VknyiOwHdHktwQP27qUUG3i+9g0K8UsAhZpNhKJCklOJe/9ER3xLRxwHWUz+J1LzWuOhZbAi0tsW
4lQOJkZY5Bs0yZPtlWbPzJ+LEOKOQtWZeILh5PjhV/0n5ii15NmTGsi4vcUF2FMgzWIZA4Gm4FtN
azVkh0Pls/b+vbpg+x6OJPGG3s/5YpPgGM+Z+Kldwxt6qDpNKp9nf/4pPNw6DcLHHMPHMHvw1ZYe
GhzGXS8iNA+N/0YcyfE7yzLCxy5B2bVic1kXHKJQmkXiBcj+wJrUgvSg2Knpm5xtfCaVFvh6QnaA
A8g8fYXs1gkvSQDuS0frRw44G5WNSIe9PTSo+6bTMpEtw+jk1bVo/5YPRsNK17M2C3MuC1VoY7zI
X44LWRiBI5cevb0H6pMH2f/5AKu9WXijARHo89B2+JQzq4sDlP9L5/qXyl4FXI3cue78RNWd5u58
Axxyy9nmDwcq1U1ss1SVsW4QSmPA+2WoofOj88WWEhCh1w/vLGcRmnWm0leK5P9PDCZoar9efRAd
A1eHn368kNCkyzsIKDZgjmZTzGNe9nKcjadHPtc72ffo4pxv3Ztyh0XCG6CfdJmnFTBi2mcZZxV5
SZfQjcTL2W8UENJzfbfIowECUStK8OekzcSrLeCXWAjav69yo3EZhy/CCxOQ7Qqi6o7il5J2Q4SE
ysj8yNc+rWBeER93lkaIVcx9d9qm48FxkdkeKDWAi0avtjW5d6tSffbzAJQ7EuKHOnXaZ7RIGOnk
NH3+j/dJthkUnrmz3tVkw2gPSFTTT00zkBEV5HJ3+wzTijnuXAexTqUKVnJzaaUeNveeTERYbmcI
u3lV/UII6xwlkV0V0pvHdpg0vmee71jeaArc/3GtJuLm4e4wHsSFLLaFjDS2Gk6Dd0s5r0Ske1+K
DbdnLKJC1KuTXT9XEEDN5/FKSLDfsJZk5GG9OS21GWkBwFSpjWBoIHGJLynRU7B8J1CvZS8pPBBN
Bm42+9NvZ58AhYtbrfcpXC/nueusc106x1bsmgFQRsJNqvkD+m0k4KSEnCjUw/nC8wFRCoo3+wkN
vWIP80Q+WAD0BTOQzEohRLE3rmZUOzQiPNsbcTjo5UTc2NmVHH4QJFVgV9s7zDQfjSZo5I/JLs06
MNUXYqaoXXq4dWIdHAgDsJNSigBlrvB9hi+juJ3d+TCRR09LKskaw8xU/qYLwwDyy3BPYs7nJUdR
SZc5YI150avJDnnv4ByIIy5Oeerxn+n4AahcenfTs9YxgCUmP+r7hItEQWGn/vzmxaemuoqpXUbZ
Y3IB6ebH0eG9XyXnFnf9A9X9jZGXbmuQeWgQ7D1WSdCTHwXBqyldY7ogcwNYxaZiHlyoSqbzOp8u
37VFfiCsMbHZ6eryDadSsJbUf6019xECai8/TRAI1PowW74ZUUpEtVvJkD+s/0dy0PWg272hfT1s
dLzut88EdFEKbiAwfYcSZKt9w5YX/PJLvsk6f1TbWmykomNurgv9Xs61wiHWwMHsMowGUduiP2ns
ycXD0FV6eYD5npZ39WZu76XaunmGfS4PfKjKpK/lNaqcz1hPrE+u42EWVHIY2wOvWx4Q85srj/9H
CJZRuhR7ybOiOMK58auqaYU1csSjhO7oBC5Dcpqs0h6UX95kTFXY+atVkkIURYNr0c3MTby8rBOL
dJR4uNp8C6PwtLVomiSkbL8JF7rHgc8M7ervS1S6H0NSNvLBmYCd089bnV0akK5j8ehDn5EA1r4R
ymWg9VE6vK3drIePxCwrIgX0bxG3+GmMJG8LQEiOPButY3KMrQDyEiDPxpdoyCvOWnoHL5zMgyc+
KxuRVSnH78t70qpFdLE7aXcyq6Uo+sFg7VtsD7DfHPjDGPVKXnKP1x8qvKrRe9ZSafCfJZjhWJNm
isOYdp7tfHCgx+soXd0jZGxNH8sEarwNf+D23OuwICU+5JLgCYlSquySMZAGkU9qpijihN9uOQT3
4OD8Af1Jlk6lELyC6WbDzsKlu5hCDNfOnd4YZ3bUStqg0f1jyBeeIqibJzMCpX5WbVoHIghm6vEo
LZKX1c5+Q0TJnTRa9CVq+VST+UnRCXYPSExb0xYQPGx+OxBavb8QCAcwyFCBuXUd/G+iCzy1V417
IjTTHb9mxhdNkVbu/APpsmLXhg89KJUOv38bd1EfyXUzFu4yzW3U6c46Vyedo34wRGuSXtUjacIa
z/XHIjD42s43Jjbj/TV5D7KRIsC6UMx2lF5hGFWKRZlGVPRlk5VDKQIw+4hnaDOR61I/lCCYGNDH
B5MbVvdxbHwNPsPxF2DBe/ejrJHGj62/AcMji5Z7vmnZXhaMNvybuDIIXBx/zyqozFjWSuvXBdKL
5YORxCsvfW+Y8CAFDXIsQSs37O2RgwF8iDMNv4c9HX4Wlll+WjLoDLlk184vCi8V18pUV9eoB7Bw
q+NjtNrqYxwZ6C6rPgZX/Ntck0USUpa0FNgnqa6TJBiEx/tgtRazr5iLUYUJvchOoERNxvKQGFFp
GpilvCWH59VW9O+4ikx3fv5HAC5n06sMkp7LeyGAKx5UWiG1KLxrtW8ZqiXY623e8x/3muT25eeP
y7MCsnqwUjg4FZG6vdVdploz3P9S5vCX9XpOqWj/eSSiEl87PGVqjly+SspsBxjeapafJwmLSaA4
yCL+OODc1bnkBPhl3qUwokRXZkIOkmYXOaa+Oio0XagIZVNYkvF/iEUpiQTn3YhTV9eZvfF+hH5A
T9NdqxgkJJKCpIDaehEU6hnx3vbNcxjkpg5x9fSmRSs1QdZY0xVpvA71ZxZvLFxmP+N3J5jj5Kb9
DZBJRolPfj9fZx0FEE+eglgYENRYxt4hm9DgSLRyejk6mJJX3lA2+rS20aPWqbARNLO/duMWUmd7
2ucGo3KYYeLxhLtc4nwSMnJW3WAozxTqk55VctSBViDQeoxxkeeFSC0/mVXj8PigWZLIHc7pFnYI
EyufZBLql4N8C6Y2gvcBYYr7AnEKetlcOrTTz7weYlQMRb4OddOuB0wnTLE4t4pm3noQz+RtwOVi
kcZd2Fq9XAwxNRdrB4K/rXK58p6RdRAnFRJXf9IIj4ENyEPHT+zPJfKy2r1FYqqdnKIHpdYAjBOj
D22zv9eftoX9ZW5/oWvrONy+j8iv/c0lv2hP3ZUk+oHGq9efmX/fiCgNcM5ekms9XPk8w1g19I0a
8nII7iSIokK7IZNPguO5b/UG81I2OMKS8hzRm/VBtVnNdpq/yffPyyj2qL6h2UKnFOexdf71lkuL
FjEv0urfG+qMpbqcqPijHsF3xS1bQPlaaS59NNIOtI0wWMR52PhfqqSmbZwLowO7RuS6jjUoAkeZ
aLVvYom9lKTcTGKzmTIyQiBASIPyTODgPgl4SuZ8Jb5nWtBLckkuAc+zZ1vai2Dd6U/LZpfj2mJj
B1Kyes+8vl+F62yaQ6yYNL2s6Dt//7WxXgDiHmvdVKSipI1UFxPte/JH6WPfk/W8f5n6HVBK0hMG
OVFdhWOb4cmICkfK38lRViw3vJVymOw3xYj+pWUNjB3AF+6vCMtPy56WSzxE07928M+nozYz1X0m
Jf0RB7sYtUb1592Cnc56J9ympV92qImp1dY4lqKoH67ea38SOMRojPW67vXuGE8oaYBnELd07slW
RQ7L6WVr4SGu94tXd4mdce0s6W1q3LM9GAsS7M0biGc3XgX6rFA4PsgYLu6mPsC1EAQvxzDzgtAD
3FTNBNctqx+CriGkzMGdJnmfs6+C8U9L9iJuOSDXurmAHLekRcxWBk4mPEuXCumdk1jt04H5P1yG
AVgRBsMZPCGFPxqI93MZSC06D608Pqplsk0l1xIQRqc1es02zjdqYjUKzRFDlepmGb+bFrR24wZD
8F14jeNj1+vwJ0kxFdu64EDWyXLobrFkdQpc8uKmnIbS+t+FwfU9wmZfdFD4mifNpAIOtt9Pe4m5
Ty/pD5s7YIywZeZDoA9ipOyjyBK7WiFFhH+1QVPAyCSVcT/8vW85QsluSLofiomwmNAGxMI91KPO
/tk5Ugv9rG6tRIs55qiNmwnbvP6gzlS8+PZXmjjRQaVsKWO3ctpRATd4Hat3n9ilVC16Q6b2LAIL
556RF0YR4fB4NDHJTyfrn1NnSpU4rDEU60g62KmVfA8QZtqN7THFgtF6aKpPxUM9kysVAR3dfZNn
Se1udkMZR6DKdYoHcibJfkxWvf8IfvY3tqHIlaNbbupR4+WCNnnIWQLVJTiFVLRgVlcfeQFRRqmk
1CWO/C6ioy09L1oQMGEts5cbJYLZyqTq6RRIkQwXeCnNnwcqiqvKK51+yw/MB6/ooGq1bLpcFoz6
h8qmKbU/CWM/nMk8CcTlWcd04M1dnJdw4AD1U59WdweBoizKGZxAgahH7/voTkf6lR5EX6HheoYx
Fx6fC9sfFTBAmlV2hg5gXji/T7ZUXjijYLC5P70y7UiAOK+VOxnq0llHcjc/oQ+lzQ6KFGZWyYyN
HgJBeK+w9eN+OyCVkDXxd7KeNEnpzOMAYDnhhKqhCTmZSSYwIFkvD9YU+PRc3Pm1QQdy5jB39XP/
HElwQ09pPHtNcXIcTFtPSMkQYmhWB8Bb2GZY9xvvS7R2y7p1MzzcPy0YvKD8HWetUCfGa/2jPzhF
3S9+iKC9s6VFpLdmuRAAoACxsLR8IAo2fXKJLAx5EWsQ1eVDQ+tEU8ghr0dxW88OFpkHLAs4xl5b
/uETF6tZfZbppwwskbuq62WZeu3tLT2pp5ziX6KlD1rm2bVQZG39ntHi0X6Dz2uYnWPpFkIDLUXk
8Al1ZPUDJcBWQYQzMlyGGbf3i8mSGWhvdV/7QUiNATDdyyzY5g7DFzyeCfLfRx5yIgqFYs7l2Y9q
VW3YJd6XwMTLteax3s3DL1WQhwo2OvYXnCGX1hAh0F5NvvBUePAgV/bA61nD1EWUpBD82+QKRmw6
gSQXYTmzSfWvqwuaqnLW1caLFNF84Q/rR3RJLuD+HiPJ0ueOmzaj7ddXag3v/yitaPvp9VI3Suul
e/bhty9x3SZtQSAuZT/D8kstSAA8ZjLtaH29Ui1hypGNXN8/1QA2EfB/JN4540FHKcvrcgRlaT1h
34by0EHq4YT3PVqYgFwWaBpA8ctwrc8iwOm6Xeff2NgJIWFfSAWu83vR13IPPQx63RmrCwChjh9x
SrOEChOq+y3hUAy3A1j3SC8OFzdkql5+dUPguklc4USq1vhErYQNhfKJHHsGpFv1saDT00mfDHfv
uMJmnccE7WnEagoQf6QnQehw8H0ugUo2Old8EYMnZic8dqGcyT23+zcH9HgW1Hq+OMWQ/8Ga5f2V
G76TkyD7rv/p829cmXzW9UuCcdmmDQOtvVwQUhuegtJT9ZcABb9D92takrCLdiWeJjUmrTvZODF6
1F+Sf7VDIzgz9uOzHV02NPCyN0AUzMW4OE+VMFB+q9u1MS3Kax08ufmdFwFC6LD3y7gRkYwzn9IH
5E8Go8QMQuW9cwBToMweF2RbmiWiC0XJr8p3UZQnVu4ulWO7LYLdZuk5vPIWRrRAqxALWNI4cNHj
jRb3TucDNvY0vMiuwG4AfrqmxeYfw5y6DQrkC4wp7EZKJpGHyPuQmAQPsp/xBCpmKO+qsuWaK1D6
3ZyoQb9jmkq9nILK7ORAurMF+F9zx7+Kgimf2DT+XhsfhuRtYMXGCIRnfzsCcyu9/D6cwlMtQ27S
g/XHaWaVwFb6BcjIP30lML351cwkRgRk8184/tMOvP6WoHN8+CCM34UlmyR+PoPPWFabnXSbbDJf
akg7OICHtivSFbn2voPJ9HKLHO0hOj7Bs5mIvuNkBDvCPtPlRk6X16anwQWv3ljHaTzmfpiz1drM
SPsUTjlhmXYpvbhrcbP6q7z26rGmVyk6JiX3CprRWpNJlDhY8FTbotdnCoX8AKDlwcrRzuiTaal1
c1LDh0XhpNmdE814BDd3rF8OvufmvTd7oKJV6ogQE4UxAnlMJ/I2xmuRkCLF9ZAgC5iWPX+ALNkH
gGEM2Iyd1fqQ6iGKsUGR5PHto3lXgPXxPtBGFomH52fIUWY0B9qzd+IniOEAhK6igedkLWZKMCsl
jB4JcBCulXa0lkAgPKcIW7Lhl3CrAS3JLftitMltCT6UvBZOnFPaMHBI3rl1KtQlHmGR/T/DRTEG
EBWZ5dLz/+nw2OJ+6qCACJb3yCltlhbKlQIM6EVwCztGxGfjFZT7nq5bSI6ZxRe8edborPVs8zd4
/YsG65D7VshlNEb9JEgLedTkofZ8lo4UiJtXeLmorMvfamouwvRwYucWBLPF/ugHpiHU9W2OVi50
7B+cQthq3LWIFq0iBNByyBue/Ei/d2sA3V+oDX3B88sxVUAY1dWy+JRd5APV75RCO4cfViCv+Ut4
FT2ISoSTV/F8Pr8XD8BtQiXEFK5EmiBhgWPsPhaQVUnwrlXRtntGAI9kGusXvFgRwLdVCLXkg/7M
+KQXyG8DpRU7hPeU04ZiF6KRip6aEaCMwmlVD3IMXEoSl/63BKDCqp/BV7eIqtN0FrBQPgxuABtx
SVbUB+pLhLd2/1jtVvBAInn5O1um3SoA8OJ68Al36M0nQoqMl82LeZBPdxFGaipprIoTGyfT8eEt
wuNqP/M7FXBvZK4LnNMHLAF6BbsAUuG7+4Cd0s+QCX25av+m1DiAWyV2mcnIXWB6bkPMfslSychr
BDGXyuHTAtV+VPmn7tZResfzn0BUYO3TCkszxTxU+Gq5b0ngDRh/dArV3ywUaPndxgrtMbDbI+M4
AFDByNSo4Tp9EW6dl0bf+bHU2Ls7/0VBnIXw2gmHDJ4qKSPwNtLsl4P7QYpk0zM8dpnQ6QV8J7A2
cW3Bw2rSxmVRXdj44k626hXaUFl8KrFZ6V9NDXXP77bDmQKLUzs3lEism4GfW2drihVzWEyCng+Z
e5x5r7MSKEtFwCsCTWq+gXg70cJwlTpkFs84zmnmiXGZ4GBnROFkNjZ8A1d5NCkDFuQz//hVcZgm
zs1qsVIpFu3P2TUINPNUk+oAz54b5wC93SY1+noG+NixyIEO+HrBnyCnqkDJwNZfJ9oAA5/mnggB
sVwObPVytmdax1J8WkWfiJdCd5/EIz7tYViqkoBpcMd+o1peAEEc3yqDxAEu6USY5gQDOUA7hQVD
3LC+pDu5ajnvjHBh3meIvftDyCdxeouyr57+dWWYWIu+dp+H3fou+Y0OGGJ7p6V9c5BP6LYEuP7e
o3kI3j99O+zfJbwSjamyybyVca7Iq3aakMp0QaWQO/rtdCnsLvR2Ab4Mn+P9oFfB9yqtS7mCyqoL
CjolpPUTcLX8t/fkqhUACk8Y323tF0J4YVe8M/OB4Xr212vveQmL632c0GVVy5DLvTlpliSRp/zR
sAZr9AwL59YFAEHfrUnu49l29n163eOe6d3hodVq9eKQUHJcMyn+XnXaJ0lgK3I/ELgXRVEjJ0z6
5nOjVx40PZJKbKIFrNpGI2A4P5IY+7+9IwlNh4tH+2q8TYQay17XCENTCjILarCcBLI0GOUibl+T
XPUyjWyXXUSMx1dLataBvlCCRdBTkpsa0FtdEtNnYVYulB6gUH4vbmPrrj0Go81Vvr11Wp/bP3C/
W0mdhZNkDh0MTgtpImwR0RxK5ugQ6VsizXH3TcXjT6wcFSS+NPkJfFoEKmGMgKg+lW6TTq03yNDy
brsm8aRGWHD26iVsDAh3NjZD2qv3Vn3s5pVMB1gqOlhH5A0Vr1au/wtZUrkl4F94RvJncUPOevcD
iXPSdGDGoeujIPZrMw99CCe4ZEYO1IJc0C6tQDAZCyrktG4VGvYdjNEvPTHJrHg3GR94d+P99Eq5
DzoNoO1Lr/B4Jf0k3LSMjVXlFeWWQx/u2UjLadSPYHKPSBwQ4Ttn1r0MXpG/fUVzAPLasOLyXvGR
ob+QYA2qpxDgB9/j0+fHEjoXJrv6/MGHZUEZ19lqEwGVspOnc9qj9hRi5lvG10QQq01DucPsZWDN
FE6gHf/j6qNW0Ea289WUzpfLurJ0GD2emdlOZVgeFj3Kz/lajMxee9EHNAnkltU1aXBwepeFhi8E
G5OgMOU1MPDPXZow0PED1jv+/ZjmJod3+stCqCB3hNnYwwk6fwzEVF0K9wzYEj/if3wb4O6yt3YY
ZfJpVAuAyh6bobw3yOCTh0NRoR+VW9YGnRwsqFLncRgYHSn7SZbhRb66X9oQlYPIsyMoZTBJhQ2n
AkJMmxxxS2e9jMdg/dFVnUqL8EruRdf4+ttlH/PNW3kmjju+YFtW78f7ClYHzYBN4P7jFZU7wS2y
C7pqFX6FXtvJ/qUCRHUCBX+vVa3/RBYgXneaL1Bp+/aXBVI/pdaPYZKOSlAR7FO2ThytCEIhDfX/
3RiaV95I7mnWo1vrx6+Ioc1zp8ow1M/xXapGKct7rZxlTC66yeHO/+AteZPQkwaRt0TJmhiaJChH
gOwlpsLbtN4PxkeibEMcuoqsGDkVqA4wFmP1qW96BnXPBAvChSaYia6aVYavI36oBYyyB8NVwASS
D1tHlVjX861XsAgvlXsnFkNhecI0wec7OqBG/fJjq9CPB1ZNVQ0Q7ELo2064RchZayN5kxaUsJmE
nW0dbWIMioAGbLOKTuMbqlJsuvc38Ca85EQCBDWDT39NEmsyh7n/QqbLtWRHieAfTgV6hinFRAIO
1tVAAgwQFiJSuObfN5pHQ9YrM177rcrwn2q/tyiDKfdC5/h68aKe0GGnAmeG+ZjdAcdAmd3V0Q1e
Yv/Meg6iTieQZ9zb6mYKI0RqmGZiTgv0mtW8DGThH9qMCX+rCwrlnleIUAmw5AjUxAJiu5RvEjGV
i3bm36NwzES86cqFp5bv969sA6M8Yw5HaVHJQqakmhCHxeknyH/o48y76EDs2PcaC6Q3nvxh3WB6
kGH2FJfT7KLQP+DpzHUFfa2v1BiDhIvLj5COBJW7P6j7QED+EFIGX7fcj56guzTt4hJ8HLwVNMpp
9havQ057doRrLNF9lHiWbET7/4yR4rvCY9gFO/R+rfcJB0XLii+LA9F7HRaxmj9PAUztw3kHN25M
mqp6UZeRoB7vwqMw1rR8N8JkGy3jeyTmaH/1ugjP5JIk5i/asBLO5fY8yDCpxPGM9dHhkq2oG281
ItezVeWk2vCslIRTC2fz0xrJYS9LJqs8U1O/fbOYqCggt3HhbdXAIk2NeIzu9UQvbWNVExIgf7c5
lNLsABYlItbk1bsHo4W5XEPAKnlBpATGV6O7bKcs2z7OVCWvR2uQjFYzWxQheLyPhP7bpv8rni4C
R7gk5YgwFAepvUCiONOgGpQCOBAG4jU4QB3CcyLnWvfrTOh5Przg6tIdITxiQ9/xjgwdIZj/Go8J
rjl0CKAcZ7fTLf8ZZeVe0kCl9zPp+exMoEhM3bpBqzxeg0RsJBCcZmSg05Acy/Vmv9vz3YWSrDOW
/sXsjMR9bfmlbLwn6MgtWTUjXdsQ35y8OPEnC6qDUn+3Yb3+6uViKoP9b7l++qSyzVCjinr+rg2b
IkZIt0L/JsPIj8Y8I1rKEGUKmeP+m8SdW9rP/AlK1pxyvRayFdyvPu6iUHFOFaUitAEcBbllxVot
gwq3MwvnmA3hMKos+/WAMTH4H4bWSEl7hNAmExNdCBUX0XfEdEoE04jb/JH5wW3/EMpfTOfEPBOM
gLyKaPiJDDVvHKrjD4SszpplnIbCaOsXg4ye8Imd1kajypdDqWCJlT3ijqzz8ob1A65sbgqdleIt
477tYNP1kCHeXIoym6JyHPWczYcJ1DooYicn+4EafzIO/H4ttx3INTvA8bmEGkHh/bDnYaINHwXE
5TS0xUZa8wGUfgK3u/R4fEm/csYeGtvlpGb8SQbtbnpJsGW6puCx/x5Fu+IzroIEevXr+ThRxcvJ
TEhs/PL1YCLJqEwbkQ54rsQ0PepsIGfx8pfUWKZ9fYUq54J2uQcU/B18tpG+VbgcfiUSjisabQLz
2XNlPtBXxr/v65E+3KkxZKOpd9cfUL0am9J73txolAnfgWVTl0C62+eyGPNQnOTMEJN6gjEjIgja
KyuWRhfn5H0kAyR1uKDFxDIKF1glJ98UUq00uq2REGjAXGlAD7jTUyn7xNojsVoiTseB/PADWJ9S
gDrbmvWZTtnmm29469w8IOCT07QJGpfNZsNNfdIVl09gE5+/i8MsorPi+9RA16y+2kbZ4nn4XanC
iN6tSZhSf5SArTP8cUcaJHJhUZbFBjbyLaX6YK20ClUk0F1IjFvBYHI/tZ8nBvI4GkWfJnzFELV6
knWfKjHCkDWyHOogasKkddyPFnYCqlmvGB1B1YzQG8db8FE/+xJ1VDfRtUuUNuZOxr2nq4YsSfaT
1Zgu9J/UXkxHkQcGwmHmmFT7NogYKO2F3xknCG4682hXzu+Ve/NXkarPheIcyzsqppx1jFFIhk1Y
/7+IlbYLskwOl1F/aLFyL1xHwTOQUJM81Cw4ikVv8hHnxlBIrZirIM0/H1Pae0aFRejUXpJ68hYs
Lu9ZD2eLDJprry5ay9maxixvFHmnsh0O3Hl42E7af2ri5zET0S9yImd4qHTpAZ3FDs09lINrbHfg
L1mSvH5Znd6GpkwZcgcwegsKd4vdvL4jO9XMBAEJIuqbsgKHzyn0ECeW0YGtyUcuogjK2505gktg
RxdcTMB19hVTKDkiHi0pJPGITWh9bbK/7jKbRCCPGsxH6U3QG+qTIZSJ1GaF/xZ+88SCIr3UXlrf
rbURZw//f5BuFCLlPfzsBAFCB2vCOM79fliv/heRWJSRwSior1z0FyrUcdlcQGOi5T5dFyjrNo9z
Ahr7H/vvL6VXKzEsLNpmAFSrub2uIgowgX9+yYwZarn989X/eGQHr7H3FpygMhvFQQuW1IViiUdx
pGsbM3XTCzLZDYwuHiJGdARZGa2VhAUB9EsQKZQAsEKZWaGsX7sslsBv1URU57CB+jmEtWyDQxMw
XzTa/zMbkVyfgp6dM71VjMAZstiyy/pVKSQfKsdN/MySNu5W0Q31yg2wR+BNyl2QJuuOJOBfOOyy
zYpmmf9krZgsEemA0sq5RW+IcfOruMqo0im28xg58ilquysjDrUkOA34h/OOaBf7A5rRjj4i62jV
tVP8ADceu/MpclY92DkPQkB0QNUC8rw9DS/EumSv83ElYRoq0b2gOtBmSc+0gtGDLOugK9LhQdCv
ao91iThpc5JFgadNA+2t6sJztaDcXCGTPY7WllGaSLsm0YzKFhlMjTL+TLDqSLq9RxaybU0Qref8
3Ka5Gw+q3OGGCuKjL8eCoUClTfVvQtRGsuKpAVcuyMYGwDsQZsp46D7p+tIBynMJCO7RDaWmLLqx
9ahc9zlT9Xj9fjYw7Y+Pk2uLyaDehKzf0z2uo1Bb2RLSAf34A6HrQO67aEISc0bwNHChKvg2u++g
dQYOoyKPdJgHagOpaeWP9Ybx1sUy+R/UFr1Z6JQ2S44nksl6Y76wz6jsRJHG/al2lPjK/Sy4KtZq
abhAIG9oQZ1uvmqMewMs0f++rL5jZtMYO6vG91TInYqNrlvJ7mYUKoVGmxoj53cvtgwMPxo/SkbM
KAoORztiT/QVgLNdpFJj4bcPRuMtwfnNY8L/8cHuTrMvGWKX2phXmlyKVAv50ZCNdTxhLuGA3zWu
h1V/XGlQsbA5TWH5HfK0/XdvWlREOGpvEBQVTTTfeG3hi4GHxVuVfe5cHpNvtd7t1MpcetXImz/s
Vf3g/hsG/R8UcpP0YHmIaH16rM8t7mhHrUGPwyrOu/HToJdxvafQt/C8UsRA2UFVbWvDOaNQzJ/f
MfUS/XPobO8lpEbikt4l+P+7kJVLW7Uub4WwzRWIYmgj+iXyehAkjV9HMlj2+q4zpF2mIv6Vu37E
rfA7LmeEyLE0U8HRX29YAcnkOrXUQedyVAYNC830EDxCx8KPPZ2Z/E4Up18p81PRGU3O7LSpOoqL
gsgusbR7ZT5A41dNENXjShEAqWCTXuAlufYzmEQdRvdbXgSRs7utjJRPt+VKoXJSBXPSEcCr7cgl
igtdjcD5g0DLZn30VHjiVxvrDH4VreJEfmNqYQN8TAX9R/F1yzbju/9JjQPIw4381gsirlX5nj+V
fAUI1xYySz/UavBgwzC3N1ryUGAOJ7Y90HseNavNozaAG4OVsY5aoq9s4vt2GaBQAcVx44ftZGld
pYUFXr9R2Q05Y3hUi3gViceB0YpJBZa4NWLFHa+JElok32gI2O5bvlHivKSGX1xsOXn+CccKzOCf
dMH49bJl99mrjGK77eZEbejvlnxX0Jd9ZGdfscWFlPUWYzqL+NIAorOC4T8ZnaQYWaUriYjTqis1
OVoR8woLJhYhLRMzBIl9wK+hH/gR6WMo/w9tBGDgjWiSh1/K0y6hJJqdHOR/OBiAGlszvYZ7mfsZ
NbQFLrYvK8BofRRlYYA02FS04EK2Cf7CEm+vUZZUK1LBSIKdy+u5k4oqhgCR0pVwUW4louB4Htpq
beWtPvlz428x1C7SqQhejDWPRa/LREdFTL47/lwRiIfaYgRiurzKSEkHpzg/aSdHAGyP6Vln5kwZ
9VebSJXa36f3rYo0hsBXHSIbeKCNivxqnItCDaqMHoXn53B2rzbpue2HBzcMiZLhQ2oDPeSlynxl
7kWue6WMi4WuyVlNaaWGTJVlomxyaOdi6+SJBU4wvCNXyUlI5h23HgmLhEflRh669Rclxiq6b0le
zIgylEY1NnJYBN9h7kXOjT/pD5xiiAk+f0fpfGIJHcxYsMqD+phrKu0wKCD507dosb9rwNrUgDmI
rooYYHrifBdx3Lj1a4O9RdlPnA7JEZGPlp961BPcFE3X/C0tJc/1xr+LNZ7pH/ioYI9tBOVskBPs
vqgIIaXPsBcGGgvrlYLnuz75w/dKVJB+w0LkNcGh2bOdgd0D1eY5a+uM01gWWcZkxj+PTVX9qWFI
vEM6BsFlcnVsEO+s+/6JCNBX7y4YsrbRpHOvLVO2K+I1ZIVIHq4JVQOn6Wq0Eu5Wn6jDKLp6vKn0
yRrMyeAw7f/w6hB0Hd4OBsUD3/VhOXqoY1vUEBFPYHnhFLuuM5yq+WFbX95YRm7D7t/xNfmmKLpS
9MHpMXF8IKdm61Pj8QMf1IhRHyeFpx2FemQqCT0yXlv8vKuDyrKP1lgFsY7tZcRgzkK/uzmHbRvU
sbfYikk6Kzt+p1Uh88kYGk6Yn7qNd8Jg7zFfkZqaAVUbqjO7TNW+2RrcEymkD0BV5wGqsSS5O2qJ
gGqijkdqPSGfWQ/ZMfpV1H29wbYfo8m2bWDYcj7wgkWIuRonr8i1DMm1n+GG1zSbPP51cdRKZQcN
sN2dL7FaOHXnUE5n9elP6KzQY9m/LcuJHvnoJ41NfLeV610cNrNisXHA1h8roiofXmibNnBIh3bk
Qv/4Ro9967wd46xNQDT4VHj9+8OzMRGuzTIeeGtvU8Pb/LQvEcL2+k8nclI9ByEqsA79ZGbDsO0T
BGSwBzwox6BeOXooeLn7gw8YeAJC/oIN9nOGtqHQbAFDA/TTD9+2dhe2JgQ7lp7ufx+nuw0tDnDf
Xq1MorhFVh0JKncyT4zBdqYrAwWBIvNcER/+PPSjSYfbx2+3jnYmW0pTjo+m+l7tEMrX/qqXG4R/
rJDu+zyIVdp6Ovn3t+7q5aslr+Ur4q/dPrF68HCpxRrMVtYVld7Yb6LYQQTJzrzdmAKrv99k0J25
3Kt39wIViOdy/AblvOLps6KAvzqYl7uStoKF0mNPnb2DNJhAYT2cqPW87+UodePxKjiQnqoSm30z
xJLJP4HvO9XldBbu+MxkS0ayf9PkLAikkN3qkobhnuwrhYK5y0F25TWNLkQtcH3cjV4vVbAu83Nv
pfgLSVbG0iJ36DZDrn07qS5rYBqMtAvesQvNdwuiBN1KzjKMY9vrLrYrgD2sIYFgIDmdKnpyVC3I
ICw9XukP0DwEGi7r21P7SpdxCQxUGuknNuknd79buA1dLOo+I92xUIPLlG+sSc4yGHmmwOMP0S3W
DWUZbqHNoaVP9LsMpI4YSxdy5jGPB9UttZKrU2AXOoq8sKJ0KRLjEuu1ShtXHR3uf0VLtT59mmv3
QFnKTyprzpcyovRJO7aAFP8fc4qo2YOpLICyEdLUgJ3+Gw34gk5sJGlY/FwYwmEiN1ad/UJZid15
sZTdknK3Qo3L2ZKjofZdKTJWLLSG9HnoO60W72D/vCrTgNgfIshSTUfDTe/8Ac+V7PMCc8hnZuSU
NKajmLPO02H81VlKC3jfJliRA6hKkZ5jZGrrW1uqkAtzJkTmyO6o4RKZVexK6auLCY3i+17qcR/t
NwQ5yXHq7LQQEvQrVQFVYGeU0rTetknWBdmQsEMFbCZbkez8S10EQ9x1SydN9X+CiEJubBi1Y7+g
MJL0XiC3jDWloskE59UChLXJ0u5hlaeGUVcZk0OJpo5IXbviGVmNEvUwQUbEosP1ykUF4S4HomXG
WhYdH5nlaf7NEAwMfJFKVhey9AD3WNj+Xf/97Ruob6pIKfDDT4DkU6IyHojeKY3ocxbJZqNbEFh5
yz9PfpKXdHwj17ZpqDKbj+nQ5aQZU//4fXMHMgEDiAm3UQyEiNyZY1r9cFBoL06fwyZTfplfwYRA
EXL3qJZEMEzDdgTjR4+6jTcOPejggB/YF76lUxV4FKZmBRaTUjyU2pPcz2iSxZjPQmW4rIyX/dG6
8SFnpE3JW0tNMcL4eapKn1xOhL2fhH1SrWEqXpU8w7IPod5hxcRF9pshM3AePU+vlxbzTuL78/tU
vZ2CAbYJboIkeW0r3q3Phma2TCr7EsZ0JA08vKNMCFIQXEJHLaUaYS4wYUMAki0eJHMFdlt5GH5x
1EUo5q6t1z8YV+gbrIjEt+YXY38rrZ+st3zS+bPO5IBZP5oL37ZnkqsO5gRpW9c1mJAf92WGYVzF
luUPn/sL+irG8yHhqeJo3HYZYw8PBgR6UEsm/8FqfjW1ivGq5sv0LQoMWIWb8KDnW5vEtjoIhPBO
8TVUd61zNSVgUuOyjLCOtC3Pv5N0iciHjS0+F7GAza+NjXAKUvBwyf1TIznsk/ltW2/a8API6sOG
5XR06KAXB2F2JFy346lBfvVtjgK6YvZLpS2k0qJpCWYCm91dCbcMW1UG0xyG1iYiT5XnILeMciXA
3jgv5LzruYbQ2LrkJpZwFyZhydT8jSW93qNIgig0Vv8VNVIEWKiZYcntZhQ9H3YVu+PoQt/lykC2
LX5QriKe5SWNPbZ3GPSzKJdkuq16Qjr4W8Af6jL3e7L1Hpkz2yMlarV1D6IfHvrhlibn9yV0eEFl
hNMEOi56E3GByGh0ccOkUw6wfqdyvLk/QLom9Mj3CtgAQpwL2DFmAqIuIbEO7qJJh1UptPxraehp
khgsiEFXYoTZ1NEGJnVdeswP+4fGvyQ1hWJMjijUrQ/IeKsHOIhQCJ56vP4Idh22htpN9b7WSKmK
Z8GwYiEPW9Pcz4tK2PK2qa28PPiaFvevBBR48lU8UsUD5GmeYaqdbEZO1V7tp7BYKGa0aUajM+pD
koomnazzLxwK2shgzYYV+bG8Ybh3aZi2HeGqm9eg5sHttaqcVByBIutwN7l+47erInb+3b5ZWObP
yBvNy/qadGuy6D6SGznmo0J0qbFHojgo37acVJb/hnoDBBEhvy/2o/rsbbYdcLghkVH/WT4JdXI0
XW0QPykgQqyzowzWIASDk7zZ740XWNJxB2u24DvOKaKLSAvYjpOK4OgXNbgxbTX4ro93nQyFWhKz
ByNX8lvbuJ53jEeE1xh4J7COOMH2w9JD/LAsCD6Q5U81eUjoVGjvIZOMz13eCbiMn80SMfkeOkZA
O4DAv2oDlWzsu4iOF7b1nFe5HqL5U9MNRiXDngCOtcQAJ3kEeL8pM70nZWYRjiUWgjoUGIIoTTLS
xk9Ufharc+DBRfD/8W+XezSYUemx02bXSfgug6hs1MJfXPZ+sKjEG1JC0XIT/UjEdlq1fuArD1ig
AEqsDGCndQzyFOjewzGiiCIDa757yOerhpLqv5CO1oSd+vIHX4WIEgFM4++UYdkHn2szP7vdTbi5
Stu9BuyLcicklAcyKRI95PQt8CJs1GYgOAinglEEmf4U1ptsfp7HB7PKZcpbXIrM8EM1yrFuESI9
6vL0weaEs/BHvG8WT+tiL1sYGkNIBAWDVNJ3x3OU3BRoG9agVu3aY+Dwn0jPYS8ufq/Kqul3SfmV
d+3vNv5js4wCyV+XqHpn+Bt69T4+WWsfpe9l+616xXORPB5tDtkezIdLLyHFbzJAlwVj1gEBhmMF
VnoR/Faf8sPo2Bw6iglXLNCat0WjWguGZ2ksjSUk4QmCpotPhX24gN138mOcqxmmlVex7Bex/XuR
W9ezSgEeYQmrw6j5E+GW2alyxGr/jlHZuTfOwdIREao6oMzCmtS94ofl78jFOH+tRXQnHTjUiSeD
lcovD+/1lxQcBguaGZ6+3Hv+jasFfkAjTUtwIG64HvfYidH46s9F/E8Bw30aryDZO4w4+tvHqnOa
pqPsK6eGwGCIsRLfKF/Zzq4jcGksI+JbaHU0EZhigUZGsr62BJd0YVzUGTq2U6B0clmjwCW5oPzv
dHUxLMMrmUpg9OPmfX4jZawzy/u3Yd9rBZmo1LusU3w6h9h0gxidRqYC0T7caJA8KS7Ns8/kurKK
Ifu5G7xLDMrOsLyKOP521jlMKavDF5bzG0/TgzmsonfBAseGh71NzAwOCG+HTI3O3/4dy/k5GAMP
GH30EMMyYcETvp1tGlJefSyr5420smB5c2hA8hKrfX+oyJvr051V34muwdO00LaVP/PXwWDM0pp9
9rwWjmWeSB6NNdUKdMhkb/TTO04qzXn7UhhSBU8jVx9oLZ7fmWigrGG9syxIztLt4cZ7KrV3YSL1
JwQgJ8IK/Hm0v87u70XsQMqqCmLIcAGqERhq5dRbhCJFgj3CB3ap+wUXKjuTAz/yh+5ElYgmR2Nx
3K82tFFrLw+61G1yby7iE0rAX46wKTuOODfTohzGNYr9TricGeZqFXnwioGT3ekJjBQMfNF9MPCl
Im2TllksFdZucLDfB9nbgW6WovjBf89d6rPTHws+1aoLSlZ7mhv6WeBU+yGNHr7FZdiixFDKfncx
WSHNUiiHAZ/VblG1hCXk9U1iS7uI3oOHrGMxfPaSxt0yjH1dkSze3Za4CVy9Tk14LJ14m0yjtfGr
s4WWqwUiKRZWTfTI4UFXLSzV78SvxteTvs6P3eoD7XqNjh8K7Of1a+041EwP3Z+AC1QrrH69jzVY
dST6TWQQNDd9q0Fua/qqJ4qpOgx87vadm8VHxzE6P3MrCalR6mvh//tTFl8fsM2p6IzsHU2ij4mG
hoNeYubfktS2xbLzC8KMjU2ebkv+NXoTGmcJcZJABEF8S73SStkWYU3YKsaaqRzkDy2T8I+4U+j0
EuTyzY4A0ag/Xi7o3/Vhjs42Vo4VrrtoTSOVlIQuwVbUi14f9strPppfJGdKxp6qdu+L9d4rLlVO
TLPdpg+JXSaKx8L1Mzryy2pzZauuNJDZ8LDmT5wrGiAoH7I6yDmSZIpPFJ72XvhgvmIV3Rb9pAXV
V497DQtmm+MKuRzMWn2xZbdMblkhOsMdPQSTXnfe4ZqRZn0WmBDxgsy3sEqmqWd1/Xp1lbbRM+l8
tEQxthVsKHh2aV9wcymoKlpgyox7VhkJdCH5DluBZ8sVzKZYZTNxdeMVqUb8cQY682ByP4PfCXdF
7NgtFXJsTQXSZT6plbyVsVuSkZPfLksWuDY5IkZrz5Xqflg3vU7252347xPTVxpK8eNg8rshoEce
STMWIwht1TVX0Z/5Gb6PogR6fr4fh7vGyMYN64LtspQf9QXyPzPvCkG12oXjIiC3uDTF/YjbHo3D
rhZsKsjVJM1opPODi8sFdOzxtCyqDRw95TquT5KxweeCddkW7zsIVjpz9Yeg+Zej54OZLFAbILHN
Tq40fMkwccZe1KW6tbGX/a2hrGFT2X+HDKdi8xS8oak9dwrf1ZM51bzYs3iBtTuaPStd2381hGmU
wuNLyOJpqQd2aDuhDMfFYS5ZW2jMns449k8vui1oq5kI/UWmBdD6HrZRc9tiYnaR1+4T8gw6B33K
+/0D2HSer8AYHBAlz9yHnRrP57S1NYk15ruUfc5iMDL/NJscF7aaKfTaJRO5r0qZBuu34SoC4IYe
87uxHzRpaaAsgkzuoMsvTkCpeLjSiz3DQQbMWPu/6lfuv0WP1yutB96CPBLsivUFTxBS+2WKaTzi
HewRQXKKy9yXnt2UPewnMM/ZH5LidsGAQmgymeZ3Q7LLR6y9waXclegYRSszbTHpvUJd9qcuKZ/f
qZxP7y3e6wgBlALTEkSg3tEvx6hTbFKA3taZNhOxMKtGzNJKpIWE2p2evQW4LYWRJyPoK+JyUDl4
kL0LrUekhC3bztWEK2qXXALKmryzYSUjlFE+jJYn+/bMB5auVaNhyZppdPooofV60rZ0pRNmf847
uGLXwk3bZi3o9WMf90UvRwMAHUQzNvOddJvL6sCZ7+Sa5sbT5MIWN4JnyPfkpJv1rfe/NYp5bgKU
drlVuuZHFutrOk7/erq+6XkxshAloNYN746+3COy5pJoU4z9YghPv2GU0FFGl+8sAKulPsPMAHdf
zl5x2gPT4sdzsiKR8Gp09vfXLCm95lXtiyxctwiolg+ukWbXQi0YEPsOfirak9re+dtdaLSzEkBk
t5ElteSqv5/vF9ZvLesFTvzb+YhN0t6AL1T7X7eJRljDLQKWwjA1ElOf4mouc8mtGJPmMfdLHUzP
0KE3mKHtwW+H679XFxg32D7v/LH61KDkidKCrc5yZUnnn1OlcM9P8wkWEXIvTySZ06NF4rO2f6Gn
xVwLaoamicazz9PHGzBcqhy8vJcAB3LQPgBLPQrv4rm0B/OzP7NgXJrP2g3zZ2E1s6x2VNTLqL+E
6rXvEh4PsQpOMywG2VmoVdmucLXb+KzCn6NMDHsIHV+Z+kNV3G20ta4TRfJHsWUaIqi0np2n3v/E
Ul3ZgoeG7ApWumhDJshEHeO5dxWuDsa77MYYNfJB/WaDohF6E5LWwzZ36TBy1mfozHb4BMb9q10Q
0c9i8BLaEQ9hxnWQ+9OP9fX3xgluoAar6W9wioJ7uCGjmOeUXT6znAQ1MR0SHyUlaHJpbStdRYNU
7wLjs9vwC2Zv6Y02jAeb8ldW9G/84yB60jSf/iBUbu+ifnoI86k7XZkwDOHy3yGDELMtVNiRbxhN
GYRw3Q9qSU/yFKOQpeVwXeOIcQt9EyW+uaBqYYkm9YoXt9gN680bktar3FDMOvHIrKbHyHwwhCWK
nA7huYOgg9m4Uu/+eKYzb8pmFM+xda+iA8vP1hMDWWfJ2voBsLw7Nvoa9opILEyDUcHConS4GZWN
0OqmhuiQ/GoyaLWhenp7UlCRcOn344HiIBPkhl+0Ys0mD5FxmKKWuidB0qaJPQsLXwoecdWWc8AJ
RzkzGvsAhvbsog+1HlJaDt27FyCCrE4Fg9zz0EwfO/cqppGRxUlm+pDaWLEMmiIKCZULZCtaEx5F
VkAtxRE1reyzYlxtSsD4Vv+RzPTcAByvYmKgZduCp3I9WosAmKI3cPqq9Y4f4oCiX4e5hMr/JH9v
i2uWhFIaZtUr9CxaLgdrUXRIXl7/xnou+NxQN7pqIqjDDX8jvI97UnAgFKAUc46Yczs4BLGY3pXk
tmI/q9j7/bmPKJfQ/qNCfG3HvtUmzr9025iXTPTSrI73d9Syk8tC+O2ZC9WhwMmjCKaIMhAHoFTA
YgY5WpbAcnRhfqv8yaQOjcmRHMteONHM7TczQlxg0pYq/f/V0E+gAKY8OmOxvi6F3TDom0FR+EkI
ePGrBp+jqmnd6yZmYU+3bA7lh/ZUPNJGyuyAIE2z864JSmHt2vr9AjtrArY140ydS5riA3JiDjao
nhoEcObwVjfLHG5uVFv/B3RcEwDcP9c0OgDjfphE77B7taCVLqv7gMCQQ45OcL8UVySTfP2ZL6PX
M+iG5+7GKzm1UDxFlEuG1b8yswqjCGzQKizYwwHi/JuK0aaWY8JIq0JPLcu4SrMl8Q2+9UADeqDj
hUSroWIK7SWlSVubJY70XpiiZHFlqNoRqOq5zzmN9DaHEfEzGQS9+3G5vEDCLzVUOp616IQV1hUN
EDfNgvcpHG5u2PdAhh+nojGBK0NjNRT6QhwsppLYRPiw+TnOv4RPyC1d7XDQ+9YESE4KrFYBd9V5
vWUCbjWx4jWip1VNWS4L2+NQCMFDE2G1inIe8JXMvWICU38XRxACc5s9Fx7bQTW+mFUB7U0Sbl0H
sLVHxu3xSf8mEp44pTYYko5OZyrmVIt6ZiGYZ8cGSHze+7UzFX0Ji75OtkiE5fViX/WtB2xsELb8
Dof+JkSLqt5AZIDvKWdq2pDICh4uPxFZDOveWnEkLwMJMAlR7tjJ8nRDjqvUG8H/CPc3dh3j0ZO4
+KTk2MPzrIBszR0R3cQp6PYdvO4M8N9cXaB0GvOyF+GGsKCWDPc7ATqK8LKqIXlOFy/BIrO0dzt2
iUE1cgVXs45xxmBs6STP7wgN+e2YxLdeqdD+kFZ5jr+HbbGzAfKvktGny4EdIrEfvPC9Ca6QhqJR
O+y/JCDtsZmmsGlTfeXuDIWbgu0HcpJHR+wItVmUxovqSE65sQXSYwjOTVtYjWTditn2M+Bdqcxp
zxSrUT6Io6LA3YP73wryXQSSopazEvCMfjSsf8J3gi0jr2MzrF9aIJvLZKxHZUxuGdhmoMTAR0oq
Q4hTwMQO7GbJZodzzT6Uh+S/am7/P4MiePAFiT74FHhHRMtftZ+TH6DRtbnMkKvsgD2AKsxUTD0/
PqNEM2gLjzgWYE5XJMLlirBw5DiSP/dxOJs0y31SYbeTQREGCGP8ZjAayT8Ix5VkOlcAOkqMNM5M
jJtD81jY6M+2359BjM/2W26+9X1FDiAv3ZqfMgX4glHMk3Q4GJYrWQGrdv9GRZxpFNb/V5mJNR3e
y/bBWREF0Bw1+ITvpv9duwpAA3QJD5lj7gy8ZdOaRxC0ytmw5eraFD8TEF1TLzP1GzDYJ47CoFYV
LSxNrwf/dJzIZIUTKo0E2T+aQuelfcEPlqhzNpLVu/KgBpcaJkou5y6T5g2gZeJ/SOrQTJXSAKt5
QwNRVs5PqeTZDJ5Jw6BTUquvU1PK3IwCrlrfXYZiS0cU1mYGG8COj8ANSOkFnvfA0pDuWIBY77LP
vEuzQkmZMS9WRvip7hER0eyFYgBxIBN5D9aOgvU08IlOlkzoqDym/SgbYWs3+Dg1IIFCZVUzxyxv
RHCoLNf98vgixOTjf/ox3+nGGAtWFBflLuQy4CHohrVRFk2NJZuKzB1i5HABj0gvmGj4ejH8GOHN
ExsZv5WNwL70kdjUoHmpT9UCHHbpt3NAMwlbUDMwWwCvXtoPIXFpz2wz/I1Mxz4vdH4Vmh4YHKvW
w6hU6TjoGjxDA6kG9mnkAIVKX3YjsUOdiI/7vkNnW43j88fT7YDljmUWP1ibmgUxRauNWCVYk/U8
MpfmUCL6+POtFAotJSr/47VKvyn8SLKsvE3VCSWlusIBab3kdeHqHQUoEQXqenWGs2M4fcGpmcti
lrli+LQA8/u1mO0xYYFfAw4VvMsOnLxnqRm7nA6FB9xbI12UNBLpyF/YxrO+Gg3XB+lIKla6O/YK
b6LSH4uJKsIakncMgO+JD8l5NrCN1YkDcAt2bF4ybAK5lQeyeeRCD7aUT3tgCGmOexoPdmxZDvtk
gy9vFBexZeRbSq9SFhDmYmvgImG7vffmcTmpTLvrMsPlkW6IDsFa+w6wwes8djWqmFC+hy9r1Oj/
r1lRgZyeQXE/agaUIhIF5xE77MZa/0z0jY3Yn+7QeJuGH8mBKpjcJnVQ9/td5I5CW/JefSoCVT+H
aoMhtvqse0hoizAf5PkA25GI8a1sx8aPV/x/h5vPdx7lxQqUnt8zYTytXPaVEqWaeoWq+agL2tJa
NOsYjkUL1B6OsejrlaCB8sBow4o0NoNM9QYjHnYub9cd7dVpB+9kfIEfKX8qzopbm6drjn2LMYRm
wJ05DjqNVb/HAPBCexphEbfwWF34SU9MyL3LZuio9qOTOccVEf8wt00VFcVKY6hxsLjZ0s5mBYO2
SfemfL9qx0/6Q0tB5cWcuiyRZmO6zWW1bZGnkBwRXvoxoiyyxwHWk5PjnJcfm5H3z8oVBPVI1Mh4
tbxhwXCK7tjg8r6ZCxrEwJbLLEStk7B1k262Jvd/MdAvZ5NxQCX6Mkzdt5XXPcjjmbQtNmAPoD30
Op24mzOt7cccJZ22Ma2D+kzMEljFnvWHNDG91NKyIVf3l5JZo22iO9+NdUon7+TI+IDBs9JUZQny
fgBalWr8rIzXZnu/cSIn4V4cvFQ0YF9T+FERQSz6LqmTju16sEEWo+6/0U94gfDZmH5ZSCg+Fk58
aJMGTT6JM9yR3pTba18dJERLBnU3Tc2phTNxFygpzJx8ry9dlsw3MATBFLsLJsx/42/teOVT4iwO
Lkc6TXclu3ESw1OXe3YUePMvRjwnocn3BzIhwsVrUykQ19LPz3hWJ1ACtMGkgx43sHjSuogr29JQ
JS5ruiXjjbVCUcWS63ZGWLijpZoGpV1Ml2vNQy8fLLrIhgPKTCOb1TbBc31avmub2ttlChgf2hnI
ElS5ckvFjefAl+DLOVvmrcfpexcFMNyLqcl80ugrHEb3jM9XYLv3Pck0XB9Nn18FnesJ6csVDmX0
3UX8Gcj2qVTpaR3fZ+OT6sLTxto6G+MZ+XlYfXeFV8J3sdXC927Qz8hVd/C/m8NWe8fl1CyiUv0q
OGy+56aJlNrtbfciPblYhrH3VP03BypiZUaUYQoUcinlJugiipHQFFRagIzHybqOEcfXooGI6/F6
GtO3l3QjmQ/eUkNreBG2UbwRqIkLBtPMCE39sWLQk/hvy0coa1KjyR4jfJ9gqVZgnB5KS2MnAvJG
l1E+ARfktHb7NnuKfiLZz4bU1jCbk/1ttT5GdLvHwSgn7KwaMICaMNjE4V1a/HWUnyIYcV0y2Bqh
bNuRtWIORmRvg8zy65TP9LMu//kjmCgnRs5e09qXr0azZ93F7KqCWuOtj1KgjOdRtix+GUAQ3tdn
mXnLMT6kKzLNLXpSRhbJ+LAcwv9HXUkf6W2i9o9t13uDtdtxYAsPHJu/3mdJDptToKKXLsi2m1kt
C5qyrF1S8+Y+/RtqjhY1n0a7BehkkaD8zxgdJECW0ZANDw+lVuPApkMAO3ZOQXmpS3w17YyDkS5N
/XlhiVK9yCmYojacKKhcd+vSu33iGlMjHaojuS0Jus7X0doM7u5idH65dNfu0+p18rA6d+R6le4s
0+isc9rFJ50YT8WDME2zTp89QPB1/dZau4Rqy9M+DvOCHakK3ITtFEcqGhmMkQ+8pIlT4obGgXSl
/hw1DJ08PpeLLJJ9c1rJxJCC6OM5jcuzKX0lN/iSjIxbeyp0kBrHjOjo0hohwNAk/mXcXkEU5hSb
02NMf4TjdiOnbE4NlKFMEMDYw9zz9BW8I06CMmL47tdl1pK3qfl44hnpFg067BYuzEUuHd5t0NWZ
NHPpnjQMdL4B2wrHj+3wG9EEtYjUaC2cmbkK9qRnw0Xk1xl8dUxWz/eUXOLMV7Pv9f1hgjzNuXlc
MUiib5w6lPHZU8G3VV6fOWiKm4plSlWVJd3obqv/5NrVZrTx2fccjez7K46bp2gS57Zfwsu/eQWL
byRv6bzaYdn+WPdzXDtf1N6DCf63B0a/Ep/vDhryOY0BYVg6pmBFu4b9SODUzYiMRm+JyWtPxWLT
XF+ZgtI6R7iXbGXwyXGpo2xTNVVTRf2UV0Pr1+v9nUN1TMTxx5hSZOubLwEdQ9di8uycHF7R/sD/
ZYpUHVEwagDPqglrn5NTRsUAvpw9FJK+/PWoXEiVvLteBaPbQIWEtbSkzOrWGrxs45OxuhmpSf+Y
6L3zbm8bLmFRKuJEJHQfhQbmkr2osywBulJgCYHIEAecZLm3whziNfPwUPfhS6DRHH7RIvQvzHCj
49FUsfaiQTvopQdjxkgn1IaIJkpFc8lNvxpgRNDya4Nn6oRjdmDBzpaDdNfdMQBXSuHfNMKOEI5S
PxUVqMzXGuFbQ5u7Wfaz6M7jaezQHm008TLOAQRcTAGb/IAqV1H81HyjQ5TTnpIrrOwyNN55+lxp
U7HKhGeJlnLWInCbaExEBRyzrDz2WevyoevL292iEMV4DP2Iz/E2Mip3e1PMMINglmk1aeW4shNm
J3ax8PsUNJOcNu5AXwVSJDKzTXk4NGfSS66QCz/bBcGs4+D5gE+0Sqhs8yeXsyJTT8UXvFHGtWCE
xRzkkhaQxWbLs/wRcvhJNcDXfCB52LVUefqfwTu8MJS7v40oSFR6Fu8l2DlG49xmUVmdohIEfl+8
lfjCEdEc0eed4Th4ijND+VwSSOd7CeCCcYNeTShMfpvN3/68ElM6UynbsWATBu4jr9sKx3h0APwM
eRUtWAL+d/bhhDq/68/y5jqD6kBeBASmX9kMJZ0plVbVXH56cIUa17M83NMX3I4MxsxfSu++2usv
HCsq9JIIgvzMMvEnX+HKkZX/GkfIvseyPa4GRE2lVBBVaJ/JgPf2GMP/PI6dJjFJhgNI025CLbos
vyl6X1dpFiHOrImbVmbzb2sU5zG5L8kgj/9s8CEuQnAdwfG5KsKimLMooZ96hckpxdXp2dtHthLw
ATYhq+4ehK6w6gD9SscK/pSRxJMY5iPDiD3P1YkOLfDkPqZoFoRL305bhtYxY79SqDArFNKqBTqS
l3vVG9XlBc58NB/8ujdJdKxis6nXqpyUcKk7GMyFHq/jNqx4X9CNJPUbZdm8vgtNBniO8oADzWE5
qfQNH+ySHhpXXvjhq+75SBtn8a1AdcvynqQPlaQGPyOskk5hs4hiCwCCW62C+BhkkvPMJxpZluze
zUfOitidhmH7EMJVllKE3BLqvXYcTw4x1lrEBeokidxSTbqwqPwusCBbaryErdX41Uw34ltHRq6l
QzTr/UThv9AuQN6VCgRb7AEJVuqdj6n6pOZV/KgTLVqds4kMzryOOa77ZHtgoWeEJIc4947atC7h
DVa36Hlrw7jY4pA5Rlzh/vtXxUB3dhrhmR5AhqNUYCwiaqHhEEp4cHAtZ9n5/d/mcAIK0rtpy4f9
lcV2jsAF/dklv48HsLGDH/qi8MBL6a9KDDqxPh9+y96r8k4oqjHlon7fjAZNf6qwLNinDLStTmbu
QS6/yDdeeC99beislQNxqPsc9HfHfoAzAOKKdiZLIPQw6FNvlHVQA39Wvk1dTYRHUp0oVmsXut6A
4cCw5chx8JE4CEcLYUIsCUwFbtBhrVS3LqSwVGn4OvB1lF+5v+Mq2PFjHVdiXF05S3FVG6OEJFMA
9xFH9ACSdD3A3eDN81tyqzUbXK8yxXKYWb1VrzyXxQrcZSkpgqd71CAT7GQEFea5Fd/7yH9ywVgs
e4TijOUH1ZezOmV36i5+cemQpnuySYYqp01XQXu+IFEf6bOx9Plhm//eXJYfx1TH3J5mhmE8HEEM
wZgOBnWW2TV53LMND4TGQ+vbNXi40yGukfopxtg7VG+dUohXSIMTznkEz5yRXqbtk0/MrjFt4XEF
w0hGWLUmKAaRY/M4uNLXCSC9ldTmkUAJoN2IOoGRr1Co9WTx1chWFS8qpU7UkwXnb/hqUF8PNGwn
EfpOst1OavEFjse/2lFHR2wGmXpySQfonxuoRImA2vVAtMntVAQ38HnX5j+Vta8/rd4XcA+2un9y
SNJV3T8PWCXZa0L37S4Rf6/9i0bSZt4Cs70XLVEzXuUFSGcbJfJKD+yDR9fMiFNOYAbCVqVv9lD8
nPcQzm9haD4ObJeZQfFDb2IHuLBTH/y7IXEEEWASatUWlEIOGyy24UWnLOBrcN+XPMGC7M76tSym
IIgRBjGwVYzK3X1fkCnx2RynQm0ZapELiX5cTCHHpDRjNQI4cTjmjOljWLkfTO1WmFKqioHuPPCh
ChT2UmcaNJCKjh5h65fActRNnVjuKptWizcY9QdpZoP5Qi2RmYYLCBxf1c8m+9Ug/wp/k3tfPvD/
ukvThYU+vmYq8GVA7F+cGPWMgnRk4SVio5hTvCMWB4EEISAcist7loX2bWMVn/hf9ns/pdbN/NPz
VHh2DBiJxE1Anm02mxckzZtX5NN1WjX0vTloqiYCxkX+iiB7yMHIcZ5/Cfbv/8LsrX6E+QdEDelM
ZMVxaJm9TsezztY8jg75eYLeN1nMZmH26VNKBRSa0xJGJAbdsimQTvUAiG7AYSvodmYKuCwfMSsG
50dDqfxWR/T2dm+ZMLLNQ9TWpaqqU69qLme9TkZ/qK4A1Ugnn68FhTvvqo+DG1uko+ZIYYA51SZI
iExEwSfheNirFclEz6Qkc38oTYjP0wKpIhb1MpUvo8wia9yvoJ81PmP+CJWpRW991+5oO/9qAyhW
mhmwNQ3KR+aDh9gOZoL8/lOTmdRxOL7eG1XvQI4Wef6BniomSU2baWdkqgMCzqjh2mKhmYgbZv7Y
JvSwFRuS5sOy7LtSBvMfLaqcs+U2gPusXIWQwvTAKWx2cp3tXM3m8nIcWDbJY6iC/H2Xt8kT80v6
Rh8tMYGujZdCUTOF9bTSln+WBbfGcpeMiJZHKwp4i6duJm7WRAPHeAJMHUMmz42IzsVCF4UqGVzP
/7CAeOWiRw04FBKxaZMA5+nhOv635cI2ZSyykt/UcK+FtSy2ynIUlkNfwQJH+wipP9T70SpyOvbR
s6UAPpwCLybDV/JsXxDJjDEKUbXPvqAoxuSMTk2s57vljkcSgqNccZ+eeIGogd9TIPgSBskJZHNP
ij2z/FZWsI/qQnApeBHOwIMVfCQXiYYAJylde3bfn28Cc7YxVsWngUQkwxAHjC3LMdi8WqIRThEk
931vsKey+duMKbMwLtUmwXXePcWxUqw66kKLDupvuXwHesU/IibZPCwwgERU/DPixjwoO2JpT2nV
bwxyQqcWCYPFLNFIZkCbP9Z1N1hGJlOukZOkHnx+dxiBcFcLejfGCLowXMnJ/A2dop2oxW9dtBlw
OnJKYCmubPDeo7+aV0/hXZNP5Ab1kuVbNsKWRGkh0T8but1fErDxSCNOTUk2DbiTY4+Wik5sWikS
yvem/UB7TqXekcK37Fap+CdXj+gWNR2iwHt9XewIJEGaaqmYS222Q/Wr/dOYOXFeggUB5TOs1eID
49ec2xwx/rd9EN/fdEGAiOhy+YTEvZtS5fSm6frFgzKeP5HfvRLyySeXSujwJrabwY2G8rci91tZ
iaKGgtkxoKbm4PEu1BmPo2LV53qw5I6ZdApZN8KGC7FMxM2OC4P2OeSAFPNXutbvg1kX3qg8n4V/
56vIg+StpkyLWrDvjO4B6JcAqY6l0vVP8FTpClTK3yHSSuZrBxx6e9+OXwgcgKCuKN77lJwf/fDq
cKXj/s1ULESh3cF3zXTAbLexblR5J2Q2G8To2lUHYel5LDbxWqHZ7bqNDkrOSTgieqWYdujSg5QJ
LtB/TM6a5JBKSwoSKmbI7lmyeb+wgY6CCkOjhuE1JrmlV0tCAV1nMIjWyN4rXo+mPjebfg6uwPQu
xd6OxD6daogQsC7bT/wJcfEzM5bwCYZVCFHHlq/NLi3f8vJDSi1PhZC+6dIQ8O1mQh3CP2WqMq62
MZ/h4llhY6yq8ranbSthxV/Xm5gH4bS0GDcPwTfk4tp+j3cA/ME6BSr3DMQuQCvO8BLs429cq76D
E2oy5N+FPdnUJ7AT55kBD8cuENGlkfug54TBeyKssX7rsUgQ5deZPhLaFkVV7mPfIsQMsjLoq2jm
qL5Xq7YMy/K87xw83Ym/45DOI6RCJscZc53O6xHN2o0C1fgBtW/MLS77krCbeNuY+zylC66xmSFG
3NQJ84+ucwf8CVDo9QN+I1x8fFtYsnAamyTQwiO2AW5+zifl5TtYRuuc6B/YnrNIZB3Tbv977Rk6
HjpbxMAAB5q5l+bp7qWXAw1x+vHOPBicnNAP3U/7Vt8fUImyNkgwIbFgUbyh/EHHbvfO444Mpxue
Bw/bn6FiE+zHyeRHO7kn3sIyAql9ypAr/HdHCUjpaACi+z+s2jsgcE/jYWuWv2JQkdzB+zB+qOOk
ZE8fX0SEPUAiBpb4g+uHe7AnQdrEu2wbCS+zsuMjH0LJ17VSiDgM2AoKOODon70KABOfgZSacNOQ
v1ijZ3Bn5uVgBnUirH2XEu8d8y7zrxYKOvqnFcH0bLiM1TJLGYbH89AAPDoPx2sEpa7Yt2BKBBUu
zQpGVjX6VhxWkIlA50SzwJlJf6drnh1ixT5tPY3iu5FklJAeiZ31poLoav5HYyPvUZo2kkknUOt5
QksKk9ZfaDZ2UJTtU/DsCGAuh/nm5V3wwPshcCX8xDbRJUI0sSk+aTRoAHrrMXuVrpx/4tUzXB/I
5l3bDL5RnkC18/1oX0QPqRZY66TZg5uJWK8eIhXIXZUc1zy7UHaT0Sd7PVXxLAgeYIuWXUb89Q4S
HtI9h+42IDdE8X5kWRotdg28BlcLk6gj505Ccgr8pTgpK7RkxvQPuQOuyTtFYBrFBKdwcxC6n/P4
/dsi4C5vWkqlnPX1N69HtGxgdoBvbhevN8nQb955P5eOBLc6HLH6OToXtnyr4We18HqhPdnznnZA
EcYxNCtHZG0/yhviir5WzSTj4T8n3RGRAG2ce7IDTD90M97MI4oi4dqSzlr6r3WUAuBMvVyDUsLf
ka2USamD52P8+C1P8ZXJ0PzzW5NKudydnO5aU63LfXcLTgtXykzjMMlZO3qjKDfp2OBMmr2KV/J3
uuvObBKBf+Q5dP+5/YJaVwSp9S7tcEOuIv8tCoZVXeuRI1Qjo/zeRhzCVrqsKpDIXrOWg8z3a7RR
hQomS24qGs70bLCB1ZSimFE3vA+nqfYyD/mvjdGSwmTMd01+w6XSFB7j0hFRl0ic4YyEGJilsrr7
l3jjzs2r4wDtCgZVXG9zWdUqeETgbDrKbKJkJzn8xPbhoNWOxVybDeI4RD0sNrMl4xAMj0zSfElt
z6HUoWBDgf2JxS7pimICrbogeIEtgp8yVFdfP9A/Pfqe+Mqu/bhdjSz/jjdZK/81Iec10aTpg/Gp
GRC023/1HrKLg+oplCMusL16oXZbi0Wg7yPSfH+BXVOQMPfhQAcP/sZQ6CQ4CznADQhIZWr6haoh
VHcdcoXqV5ej3a8FhziUJQKRm6VZIIKpLtPTC7iswyqO+Ug69EBRFJQozvXIMIemaVa2ZvHP0uKp
E9eGZtNEnqUn5Nx6eR4mIezjAM06hhjEW6wu24GmuFk8f2Bn90vADt1esEJULzo8WaedC+9QkOWA
3WbXtu4ViDHGimvZVuTXLoTaMFVtavAgZlgfUlArktm/54CO2ovVzj1eGByB1tYQJ1Eys0It8XTe
e4CoTYhfQX5hMn/4I1fCL02V7lCTOLhrsdxZnD/1MmjP9ZlwTfb5voV3qbboO25Rb5x4spTFtssU
JbH5yAWA0vjtxt548yCbt9m65aXl1kbdORPSWWwFitlK8y44UU/9FBMZcfL5d1lkt4P5tA7FxjFg
OY42ukr6EvkBPwBC0LhWtTxZRCKuy4b2NKIlYqqgx5VKAPWxDFStTcknEPdisB3Ka2qWbtp7Cmkf
Knj1jxyK2aCmfUB34ubUGb660R+PAwMsUrIFXHA//76txKzgSoiLYn6d/v5xqZylTOYsqtg8aitE
abfXMLdAmnfFEb8/nz6ORxV0OdgycHqL6+ke4ecyKHg9OkJmm9Ol/Pr5fn4ju/TuclHKD5OOF/9v
eAnf1hvmPiazThRKuf5fab91cqaPscLMKFfJdFbT5ojT98NqqPYHYk4sv3Vkdsi4EyOcof5pP8IC
4+MpXgDNF86NZ8muUztAqxPzPNmBE4ecz+Uxzv5/1FaqgMXYXhMmPBm2HjtWbvStab3eNQlxbYuZ
f4w5ikaY2iT41Or7uUHmJ7f8efdwWKJaKiyhi3USo2kL2vWVT7xT/UvUv2Dt6wJ/IsXH7hnHo61k
P5J67CK+ZoLyLWSLobjA1gBPJG4Ox+DrBy1XV3YQaZrY4RCP0AX/N+V4lkbvUs+kcDKfWt4m+zhb
ct1lp+N/OWaW8tmD07xFj9FT99wsjH2+DL6Rt6yCtRQqNourY7xBfC/T9P8ya6qRcnIuelyqiMk7
9zD2udA1xyFcg516cl2Qysy0tQnE5EFfvho11DJoIuNGiPX+gmwZD+XCdH6GbuvJvRGed0OXD4Re
NUx0QfjnissIXwEVSAfm4jK8/YHEAynnI0V0Xm1IntUUC46jsA5fHI3StPYiJEA5jQICDI6DL56J
fwM6oQO/b0of6jOEuJBGI0gtnppG2mjjAkWLo7vcSWiHCAJGlDACYLD1gaGmaT+uGvntMNPHvChJ
ToJj5AwXZiPgZOxCgJRLxhLjQ7PUJdXJTwcfV5PXiIhtXz8tgQylqMepPOzymFe6n7XsxurbHvyX
ZottHrxFk99US5Lx1jYYH/0Hiz/zTR9OYd8lzzCicWHlog32y8mF9bnn1ZldGb1ssGFyzkam9oya
ezBHvCGAZfV15ilBckP6ZLbQXS5uuCyyUinGyZO3zJyotTCvm/ZWmyhSiprh0DLt16CUNqoAeIBu
S4fWY8AT5E8VM3h4iSJ0cmQaZM6JPDK68R+FvhNyhF/tZy59CMWDb9m5yEfPBMlYm+o3ZLmW/tfM
Ye6yLiEIdHguuWopjAPmU3q05KszVQd+wEgfYLK3UhBJG1WwO2aEHu8vAT+G1Qmlp4Wty7mQOisX
LYqTdR+25OteWEytK06+LmPVhT4+jahBKsRXN6eDZ0O7fmpV5/p6yvqM5A59NB9S/ZLHYEdyypIR
BHsqo58HB4PnHByp+IysxMbvLCBA92VrvQp1RABBurHBAcxky27s/AqI71MT1/ZYGdnHDN7U/YU/
3aFji7cN0M29PDM81jgA5tANoqKGP6PIRAYI1sD0rGVguRme/jjDg8mkwFWIE7mYMDGUt6KiHqUl
UqVhFh5ckOxZRETBe22hVAIlBvPS68jjemxuwoGbt8nvtNd9Ssbbm3A2XwCRmC6V7u34zNouBbeV
tF0nPTRMNsKRaAkfhJNyuiq8EWwxQ/jE6I+kUaSzNkHne6ekV2PWDKL1aHAMTL2uUi+9UrSNB7/C
s+cQu/wW0UBlfZ3AFX9D/mpLl2t+9u4hVyXKmr34w9NkGDkBe9ZACUntaj9aMlT40A2lLYAY4zox
1SZXEFy8h1+wseRnhHDqu5PmYAd0e2oByoC8pAVj4LrPQ36itiMOxTglhyAtNHI1sDiVNR6x0xv7
frGwlksteSxl5F5jmlLzFvidMeb6hKMX1pPqvfxAPGrLMVCOBpD8d1fnEW3g+mOazwhgP+Fp40hZ
T5Hv7G2MGNMQugKvra2eLp+QrlEC/Mj+0Xi0fc3YDjLAhWefG8z+EDTLa+kpGJ3k5DZw4jVEgDwO
ZCUfts7+V0gGfaDvDcmmTn3+QA/kVrknIK6CfciQe7lc0Hs/FhFC7RQ2GdIevWK7VTWgBh4918kR
aCqhQe533jnB7U39Upvba0e8GdZdhMSSwWAcSAYZq4YKTNMDZzqaVyZkSKjo2MGmGYija1BlhKJt
2wICMYAOkj/cdEqd5A2ajcLeOG18Zw1ZeyIASfEMr8FGz9ObzwTCHonoCfOEZLMAfdO3U4PjXuz1
0Gvcyvn743/yelsqQvOcYqy41ogtGS9GtxL3ydGtx8L5FaDwysaP6SDxfivIFG/+KEcS1m0LpsYd
W9/sXIADzYyJuI4/euLBzulTqSi8CMC98aSl/4GiSOfc6Fl0Wbza+/blLS1N3buq4uz0aBp6idHP
RNFVio0LQixa/AMkRaUoYG8ZFgq2jrn9W/S2Gn0aj5PTvvuCOEJyI7PXVF2oVfoRO1/zBPUwvA+E
3IDa7zwro16zIdszu4R9r3L4bD6y51tbVGsk5MkfCiawDOawhGOrYttlZpFXjzZ2sZ1p13+JPteB
kML3vy6GS1jsItHDLGX796Z8ZkWAlhbGPcgjc8Es9fBI/DL9Ingd+vBIAHm5ON7UjH/+UdAF049z
bqYr4F97FwGkpDFOReT4VRyAVoZAifeVwKC6m7x2A7DGMoOfkcxJj832pTSojgeFJcISafKqsY4n
a8qKJ7Kg0ry+aqF3j245P3D+USDhXYtkuSp5QGECtQGcHrUzPEdBrjpsxAlntRdxt/5McX4CNWMv
Ndee94140CAdfLN7ixPPTzfas/eyq1sZ1jQhf9oKXPDudvmVzNURdWc4mliLkKHNAuUNPOzzUnSX
v0KXHOVuoJydaE+3IapvWAqPeA0N9iEwjIyxnTx1UhHntDfrXBzmg9QhxxU/rLAspX5m+frg5+o3
6/s12bRKydoOb0Be265LFDbVyNYwSIxSCyJu0PzmgshFbedLhcySXmtF5TgXGR3TPiIh+kivhWHk
u8Ix6T7sviIM8zC6if/gwtxP9KZW7zI4WcuFFAtVaR/2ZlIJ058Tj+Z+MDjVWd8mkQcUjLJfwqia
eKyUluQS9/5jzE/E2QyTvWxqHyBs7502rs/JVkSgcKC8Z+Pj7GpPnIhJC1n16esnxsyE+VGier8r
IwHs+ugUPHjvNyiuXMdgyFCbY0u5lbIUh2CfmYImTFMfjyhaJ0GwCpJwc7nbirRh9UEfD6SQKprL
DSFoAfYUMsCaqEwwZOex79LhLlqcUczCk8KKYb60b3yf9HP0iiV99T051btl2mSJhf8jnh2KBawi
IXIb2JTEDB/7FmEQbMpiVqN0cLM2XVlhtLFyFX2mC03EoGXZwzf2eJmtI34c1hesi1NVpk/wU2Qx
YKONNqo+QxqMikzE9Udg4rjDMeY8HogtLU/zRD5VQ2JLLoXN1IhisyvQCvhlONwG9XJinKm1ndsW
G6QtF1baek5gdyUA4tIXHamyUw0Tw3NgkBDT0xeHfLLABlHE9I9xGylDJ6dck7WKoc6r7C19II5j
IE5D8w0/96UvULd5ZPvtjxUjpqoXPdSK0Q+RCN1O7QpTaRA5WlrVAgpq6cUhRSFDdbLqyBpsJdPc
Q7oG9MQ6rjAfZAuaNyPm1Nqmds4irECgE74EfQsacSvEZdpogQ1y87hWhBwQQKmnwJPL1B3BviXy
IlLRhekBoROfDkcw0k0sZGJgdCvup9NlzaYVDWUKwxJqvKtyJdHRuhI4YODkVvi/Kn9A7X3g2XTL
q7cEZeEbf2gIMSHr0gurf/9J5Yq0Ee9N7Nkt355wyfo8R3KzXzKS1X73FQpfpi3gEYPtHsmByq7V
7zr4+ewfxhDSgR7zGgUL1brN1MwD/6RKQw6rW0eweZ61T+D3EoQVrBrKT6Vdq1FFVeGfVV9hbfTO
Mynw8+wLPTKLZrIiPghc87T+xwT+bWyvAIeuMGuBfNwqqMwotmUgbuFHA5P611frrBU/k0gy1H9T
SaqpFBv09R2q1bp5VrE04iDy634JHXkCgrRVYRqlhFlcvUx+mrjbqp5dBgNsOKkSBd1mpmlJGqfV
9tf6ifBYXW9zTw70XJ8umTMbSgtqs8081+NSyOwy0QX/nvqIoMNukdAbm4/f2vttTO9aimiCRSAr
TmWctMcKVjzjh7GVsNpwVjRXg41o7hzUZiFx4IQcQX2DgTvSlfaLFMKKXjXm6gZLUp5cnoK78YHU
5VXjfZrng9E2UAAfzupsVr5l+VWJ1Mjw+5++SqqvOOUZnVXy0YV8EcsoypE88qs0cCtb51W+3xTc
cNn7s2+47CWS6JChsXYc+amuldEK/58SukceDgMS/Zz4MQ0d8GcoGLqA+6EB7VVM3BdWhcs7rzQ0
JBhH96Fot+ttwaxss6gDp8OwXyUTNGMnbj5tp0QxpOMjW4NQXfcvFtEV4Kqxfj2GFgitVEZz+iTj
R+o9JgiIF6thjAykEpWfgRKDHcaxy//Dmkztqk6jUFEANgstz9Hct0nDJLjBSulz89NHkTeJPCuY
PFlewoVqprKFMA9jKs+6ji23gKVCP/MtLWYXtlbDOumtTfV5kLz4rzl4Wf6bIDAVuLlYh218d7JK
ON/+8Brx3j9BE0T4a5SxZ4XMw6hFhIXXoqI7Sl0Mrx+APDv2FpG09FebWHYWt9Bi/44B2hgN8D2v
i95pjNcf7PQ+Y8VV3sQRoUoc5LOuZUsW6Sv8s7Gk0F6jF3mxy/jCS6jMg2OPe4JhhUEF4twx4NGI
cw+8KD6fGmrSyR6lK/ygQjAbn6Lpj3uEh3DTqhmfmcEMII9O6Uyhwxn666SFeTc3hQdDcJ/V+BvV
bV38LuuvSL1bOO6YcHI94bp7zCBqlTD/ogPt6DAw+Vqwdlf24iNAYKfGNdHZang+kmEjFT3Gbavx
zMMvmA5MkfRAACDuaMDSDOYqsMK3w+pKRUj9ZGp/oyl6ItT8T7Qm3Pst7ihnAqkeVA66w3YXnPFk
wJT1MegtCPRvCVp0FRB7moyF80RchqMj5UWQ9XCFReNkLXXiLBtSRtAYqkYxbm86Xy+txTnw4tOE
izE1O/cJGagCi/6jF4fI/WFPgN2tL1WWY9JnLbuC3QCTacPED/A4DOHa9yXf8f8U06n+xYoHC7Ne
GY7ZLSh2EzkUw3GR8aD1ol+zPALIdkwjr8jfWOLn9ALhH9rAPJfxNcKGJWsKmZ7qkqNv3khxPWPQ
zz+MVbyrH9c6ppMGf4lnrxRgX0z7CeJFVa0qcCcPDdZCbXGJe2krhXoeTUvWJyXupndTx7pn4MT9
onOz6KG76gkaPzd4cgBhEyM0s82FpCRbmxEOe3uMICjHnrjkVaZrtSgeU2X0tmVmmEKn4DNi69o9
kQaRUvtlU5BZ3Iy1aCTJKh9eN7+i3ouuVPlGe3q61PRuLGrcjrHCqpbjGesy/FE9jJDHoh3qghJP
rz/hwmCXXqjR1d7cON3wesL2hb/vSADRT/TO7xM9I8fGivBbNKCm85HMH3hlxpMIVEgtffZaIRPJ
V6OswphztepG/3A8ArUh2U+CqyuNAUg7xNY75vgSK/MD1KUtymMSPJUNIkaB2y2ZXra9ZvQcar2U
vsX4fdDGhrQhBlfhcYWgkgJhP9vHB6d+9JrLaT5Mz+zkP9Ub8ScmHwU1wu24qSUg+izofFz8UghF
4d9eIo8AxnJzFmROb3AH0auegLIvg3kTjrJKMtOa151+7W6uQh7v5OkKqdoM528NC21R4V+Jm/aJ
cD0axyOMrXS95xY/hib7l8eWZN1m/hrjxe8xZ4q12Aa78fdKAQ+uMxFwhJ8Zl0+7IKv159A4I5ae
I28VS62SdJ1YvWEiTXfYfnpog6zxYlHhjTOiQ+JmcQk+B0GDVcZi7KG0LJ0JCFFy4POsf7HpBzbG
7wC203TDe5AoWYm9KsVfFU0U/W/PDwGkTtkQ4kRsApx6j4kY9fvTpDiEwRnG1IsVVQ3DF2I4KRce
l/WRxuKNXpSswlv5Mo6641UI5WlXyqoJ7NPTUry0UBr8HA32119s3b1vtqxGgp6fyQn4tmJNAbQy
tjG1EDbCn8twlenvNOyupUrxmwGTEMgeqxYjSxYIOgG4Im1xNR0smTFHbnBdrdOTlLFDXQlcMCWK
4xcHbXRMAIy7rIIr6/Aysk6p3UkudhOf7f5qevFxWipn9WACgrH2HFStxvGtV+iioffNltDyrrTG
bPclh6cbtcdyiU97COnTPqU+cvFoG+YTXOEowvp3ftIIPnGUDuE6NPLAytglKiObb1FsiiZ4gWzG
OTJbrQriizfulodLdSkd5/4ngkM2kbSg4642LdFW3dO2F3bbbseOJyLgBWrPxzMlUIX91aLCtUtf
jZrqMmTSJEDeS4B89vyLmwn24h8OA+Ut9X9vKDAbOSbSOXbqdEtzMa0kcMpw7KYf0DaEpPjfvE0d
Ui9fu1YbubgW9/eQ6bOgRzRUmTH3cURwpNIgX0bDgIfuZ81HU3WFrH2WhdyBJC51rSh/BXlucugP
LM68koj5CAjNY5WlI+RWRMDd3vq0HZNrzFT+jv+/QCaGnEjR4+kVoxjCZG1ZQ95Lowk4atix9UVY
TkrGB8eavxaSJKaWeenCPgTIwjFOkM9lm/kWIQx2ZIbEoMSYG9JOBgHtPdn9AyYAHCRfnNh2F6eO
8HCrKI+XCC/ZXBVxfzP7xwQtpH3wdDMB1QNZLGsCNhItDcrHTSLRXHEcRxNRRTI4ZqbH9bTmEkvy
0sLRWgDXPtTDJxROEEm6UQ9iOygl5KyRWX1T6VqwX8Wq4K3vE8ug5Qo8AxGjXBHBJoVjxEtQyWDx
MJGPp/HgW48Ptk3AXnfzm75HR4BlzSg/f+t1lWxoi/XHCH86zhJOUKUiqSE6uGNRodYpUcz/cMBK
oh2OpsWv5j1K0k9ZypUj55frggNTWGMwtbeiubF4wz6gjM0QDynjYrd47/R7oShQyoZ8v8fSmnmn
SkpByly3z3Q4g6VxNn84gA20gnL88LAR7jIJ4DgtXK/T/kN+GpiGCaitPPuNTitEGT6lT6k9wKhi
FHcsm75RRYJzoiqVGZ5vzfJct5OloywCHxwVS1lxG7ndYvkYNM3lpIVYuU00ATQb4WDh8JAQCZmt
Lgudxj/2JGj0xE977kvbssu0K3LpgwE86EeGcSPvWMBHOBN9SyNiONtyZlwfa+wxUAj9dWT+E2P6
rwXPhCcuzGdzLAj6GZ5j9x3ReNKNWOT7ZW0sECA5DJkimr9Cx6mOupZhM8nUjo02UztFSdF3o2sb
NJls2pou4PjDNTcf+CY1gL3ysQQFjqTzh7rACqwunQ2KGEoRH2fdxLSId3m/POz9GLvI7RBqCxMU
MCU0ixJ3G27tETw0q54iveDyEVrJVRQ0YV8RbaDnoacVmJKPTnV/8aWYhdLOz8Z8ovOantulRrH0
utUsTk5mLAkluAbePX/dX/nBZ9lXNQWIbnDIECA4snlVO+nyYmw1nligYolr6KW9PeIcC9i4VvYG
3KPQJ+zcDaDa8p563MMpIJRaLM14JabWKleDxDx6YImAfgQM3ieVaJegOH63k2lXvEGJNo2qpKc/
gKsIlf0sp9IPhdZi2msVRvyUtralbb0wfreX6lABDMl69RSe9sCK94UoGBFvfG2bP6sRN9yLKwhB
8HlbphN7u6PtRml5R4ligP5hjZqu79aE+r6iPh2RlX8aszLxZcyha1NwUTzzQeQO2lWtkiwouwoF
XvuVvq/4o5nbigbQV3aZlZxgIykelFcwE4D5HwTcvgJi6uvSiAW8a+IL2lGnRxVht5PltcW+EWgK
nncLlRUNbxXjk59JZ1jHYeQKO9QiYo71iH5VGJ0e7URgiCskq2q4KC9byTnxqvSSxgTCWNqLuo1K
gK1bXRAr+natpvTW7FDluBaw46I9WSP1WzOZoG2BVI5K/Obc46hCsTCIR0zU6Q/6Ua+cCMs1V+GV
Fh+R9S9HEasLXzFx6T/gZ8rGFB6R0tpzK0CW+hZCm32DTLxps661Z+wi7V+l6DKcG2FEfWS0iwSo
GX7y42S+QrZoeb7uTvvNsCbTm2rwJVxeqHidGEyB1SL115IqrpWgxhcqtRi0JmP+Bv42pZcUo4jd
k6xQNl6EJ8Tuyp/nxBwRFHZF/xdfyk5d9wxVGhS7sbl4VDexPqLjig5hdfGtqC4t3SFqEoBjGkND
s2SqiVVWMmUrd+AHKSxAFKwacEvHB5cNl+WOiWs02fE25caAm/wLqeNUsSo4oiyJONYYdGGHwu8T
zC/fDrqAbV1lyRF7btYOeHY7mEwesMfpsYn3abTQea8C/d4v+3ZnWMBywfKESw21Cpa4nrVSrSjj
sDtk2j8vqsLIArHkpJZoFyDRDS4nxsRmcxiPvlDozXZamQZCmL/+20kqSeT4pOn/qfseOy3lMjP8
B5VpuLGNnlx5h/zpVGtSQCJjbKc3ZK/I06hQ8AayKWDU06CNo/yVfkz+Tj48CWFVIBWltulSV6jM
wTf/Wrr2QtdTFHXQ0Yyd7mK908PQVDwH9de/pvMX4S10RK0uF8qQO2+G8POzWVlEgE6d4S1ET3Dq
FBcXhvck/0aOJFieY3HevQQ8i4v8z51lDb0lQgjgINXMssKe+TSDkm7BfLSZ5pIbs3rdPQ3U5Ztj
wODAMAG+25Z9ooCfvpvWuhV6Hx4CKtLDhYPawSlBDaeabcnyZkZuXZcc8vs4LrbhfO41AqgGlpit
pV3/kucqft2VuS1Ip7cKPLWBRDMWZzhlIpz+n9kbZ0ZGKsPa+NqTf0QlvjHKCfD80Kb2fhnWgx+r
CzGBlChLMs/A+bK021YHRZCJddVZ0jh+zfRee4fUFaE6mmd6NNtwjs7aDMIR9Pmo+ZKPETWBOJOf
zPMO/YNW4zfPdQdNq00hdau1HuOHGUq8CvQY6wWoO4Wcbkqgzfv7XSuaHjwvlCX6ux8Kn25R/Yf0
kv6BRnHqDdqCEwo0ll3m43rEOmbapDjlylgE0tY213iblRiOQaaioWSG32qlkPaIEZTO/Y+x8qNt
nCVISCoIK59WfGZ9gKb7Fp/NGiVJ7Oiw/Vm2jZWGce8+KuahaXZTe0S76xg5zNdObhtNgBXGzDiU
TFE/dpqoBrXGTaUC/X9gN2B30spBsFrWg/3mAQCNjBmfEl2JRmgnnk5SVQilFs7H5lLAkKj2Qess
ttErWYv1H2o/usj1tRhyjWioH7Vk7BJMl+SfHOlWIyY+z+e4yGgd1tj6vVf6lt4j7tZKDYSfFerT
UhXc7+iSflMrQuD6nkG5ZW5kZc2edoxMxVzlDTJSjG3V5VJI64FxUhU2PyhX3ozGYmpGF1547jj3
Cw4QNckJ5IdYz6p9zFdIurjZPGNWYsTC+ja1XsQSeKRkppu3ZpD+3XBPwoJf6wj40izkfQ4R7H5V
MSXS5hTbULh8W3Kb3XGYev7Se0Y18MZPBQ233mubQzG0XWMcue7+Oh3jQyGfzGYwqt/WWkk991Tx
0rQKc5jDfzjjBev1D8b8tgCedRxvpE35wVJs3Ma71ljOvXT3bfBs1dDe8FmF9C7Y/yo0YP0wz2CI
wl18tdyAgnvUiaJQ7P1DKKrZWfy6VWmCneXt3ZE7ZJgaxNZgOjK93mtp0D6LNzwDBDqqoO3Q+Vsj
axYyxwejQAGAg0/UhE2UokDwR6TO4hn1i+ZOBgnDoYXndYMUx1CxqyTjivnp8IEbiaorTiRjb0PQ
U/TsuLk3L0uT8i1A7wIPuQewXJ2VpHP2GiLq9SQhoMJAfvHmHldQYSipKkJ02yE8ioyC3udJlnZP
tkhJOv3CUZtRPR4V9HeewbgzvwvydRoJYw8JNjThK6uVjZYPAx1yCyiUU2O5f1iuwwng6UVTuni1
ztNciInoYEtnPA47Fpey9vKc2yLtX9GjYqCW0zqCv+2yee1qnwTMlRcHHxCqtHA8eKW+keL6qjGH
plE7o5DHypUJi7up19L4QQf5fiUwQe/irXUyjqmtqCRY2PM+XS0nMdjif1qPjXnNPBd1K3JyxwDQ
eZuWA5C/GFGUkqqX6gBg/D3HaIGvbF7XrZkwtTrHy7HqwgOkpHluRcgnXbcN/uOPoCAfQZUhB58Y
fl4SqaiUL7TS0fhMIaXXT9vz16bryH3J8RT8JjlW3Iob5Yvb7EwYkjZqd+gjPKhqENixlVQGLOFE
scYoML4qH7M0yotZo3g6BMxf6eOeJ5mxAd8NfC7CEGGwz5/FmxpTxxFjW/O6kPsfbjM61VcHyWK7
KIC+1m6XWbOq1QGKZ7Z57ZM9zpkMmq9LaZrJgDBfZUiWt/Z1Qq0Jwklh44n5ooBaTsKQKVxwltVd
6MnG5CCQM1ghZt1Q7LM9ANpGMgbVvdRXcmLGAskjGb56wp7vcD8slwRZ30g8eq8saYipD3V+tzOv
gul9P/oZJdjn8t53Yay0KJ3bH9LIaxL0g8jmH8yW5OipKi6vA807M+gmXBQiK5kW447WmAE0ZJg+
qWqP5LGlFadWh7LZa+yO/++IuZVEoTSlC8IIfcxoKXDcX91FhKVNU7KOonjraCeHibuO9BfoYvEe
GJhaHWLXUrd7vjy5dcF18bq7/cytvWg/+e8HhOb1QaiMYp698R5kPVELpyIEG0Uw0e+SaLQ8L193
S+ccm341rlvob6w8oD0NhnF1kK38YOL5r58zMTPr4X4DPulIh4yDZUbE0qgS4alymcw+chHayzsY
6meV8oTLSoRc3Il8EUwyXJ7h3siYdIeBexA+2biwZ50S5JRPM3XkZBLTzvnP2gySAUfQCFdE8P7C
f77Bju611Vy/zUx1N381eUESmqxN9kWT61tm7jd9aOaA9k9OuXIEjAYsSuLB9MEComMCX6AxDFrr
w+jTxnhuc1kBh3etQfI7LZk+aF4oigYamwrCXnHtxZj+r7wu5v73iwHSr+YFncNvebRHgrHPW/7+
tT1UMo0s0hOjwPNdBJgUUi6Pov3TvVwW2/JSm3tHTZgRG6y99inB5UXJUrwCfesMiM/DtyV+mk9T
R31Y73vLX8okjQyq+HOYqcstqyqd0KSo6rbjYsLl21NgekC/qqXgcbL3bEpctyM4jfmsU8MeHlvg
FESmblGMsetsrgpip5y8P2W3HxyvD96ILbOp5ohpNN4dvIvXmWPdwqOBQaoP7fM2G4zxBpisAjlW
jjHo180T39mLjlAyU4gUvyUokb9D0wuHXgXqkpK57YLVn50/Eg9nrEFWLRxKzdooeMMmko3arDUF
d2oOxP105H717Go6/vY9z3Sr9U0MYmLbowhYX6RsNNvmeTKbYzr+R+QS1D7X8nzDpZybf+JNxBOE
8ea/kOx4Dm2Dulj+zr2wIbm43iFg++Vftz3MdG8DqS6R4IfSynuGiid5bugu/lh0UjxUO7Pwbutm
m3TyQIH2Sg8t8OruFkccM6WuCtbKMYzqYt6dEEy2qEjiXjH/02xIF7RlQ3DGlfKbxamBEbODanZv
+pnRVD8YrDlDxz2q0+vUh+rto7E+cUboA/3iX93QVWdFoQ9+hoUQxgJMlRhPQFbJshdFuTg2iS/E
vSeDp56xJlqToXus/K0ogpwCsOLUe5w2uGHsZCdmKiUM8EUPykkU3rTLXlUYUI2BA75rognt0SWB
oRA+hj4M2D13bJ0ZURr2hTdR7cziK0M+N91oGSNIGAfaFdI6qZCrzjRgA75iagCdVMaHU7c7JNkB
cBVbzuDvmcHV2eh/tfdGtmTxHzMnTj359nAD38xUv2eCoS05jx4T/ZejDvx2vVRcTqVSn3pF3Tq4
+xVVA9qfXx33TISgQc7cxPQ+6slAHXr80ulq+WS5brKt0W++jaavUv8LtmjTdSbkGoLpWEBMidCI
aK7rSp2d/7SPWUHOHmW52Mn4Br3mT1p65NnBsiztij5g39bP7ZVJni82EFnIaSo+1QIKDwOjkZBF
HQP/oWeOrCX6qEvFq0Wplx19Znt33F6jD4lGyurMv/i2BhLMfE1FH9FzGPQncOfeCFFlEi7HMWu/
Jz6yPFwp0vyMXhJv/JsN5Lfv+H/+rbe7Awb+0dIJp+3PNR8Pze/Glzc9nC1l1QwQpteAvZNMcVpB
7ZxNo4Olt1ectXp6EZiNxxECssmNdYF4NTr5vqnJxtDieaZMzoxOTX5fMYif1A1axxOoDomAj7R7
xXOX/f/zb1HrnQdBdcMMVP1Bowemc2TUwde/qLyt4vr2akfP35oYgaHEXmUxHWvlk8WkQF2Zfs3c
972/FZHW9U7fIt8gdvWtWatAtOwBNO69UjgOmu7KR4xWQuehikwBKrHwatQYunfnQzi6F1iceBgi
B2tVwMjZIJAw0dCIaiwksZm3Aup6SJo1JBqmzvsoQO6uc8AEEYaPm6LbW2vPtoV/YTu6n9UUheJ5
skGBKiXXsRYBuz/510zx5mQ6m63fDM5l9mj5o5e3pFpPhQL/zMdlq+HmnnDfiIZk/yfA6AjRRqKy
X8MdnJLSV913IECJsSDm5DlvVzFA8a/m7QBGYHclBKZBk8MbbbdImdsgta22Q4d2z0K47WFiB7R+
nOR7Sen1xbvQg/FtqSN+RxnnSJBrmM41449umd3WPDxzhSzAT7NlJdLoeZRB99LN7Kl4ZR5i6d2g
QKZmsJuf9hWjon3Maavejre5BYNTFtkeUQ5FrtwOFHUzNWmUnanr6N6LmPF2PXLCaGemIzasHT2r
9Z5ZIApv8W3tei/c9UfDMftLwG9yx5hTu4CJUO6PW/86CicHkFQb3d3zSfXWlKY0CiENF77iTYYv
xIyrBmmZcLZhvJM4aWX0/sMKOdk2Ga5/bZsFGOvnyungXHdzUz/9J+FnDknC0fT9nwcicO49FJIM
1I/edeBRibnLE/acfp5xkMVKiCHJ1Ni1jFBERThPku7FYbg/xGhQw4ariICCcktcmfuoKaMbNnDs
R3PdpPcWk33C1yAOAZGKkwhOlsVUHxFUaA4HKW88+CRXsvBXhbDFnlMKCzDVRMyzByNRdAz5Y9ei
McsE6Jt+qm0rHFiTGeftFgjERblp+1oWPNExxuvYdE/RDHZmc8/xd+ZHZ3GL0XDtwK5oB7zmmbmf
q/3OKaG6NqgC2N50ltIhBhCNKmKsyRR1HHDvJv33y3kGMqyD5YlawuhxAU8Vq3W2u3MfLfwNB8Ri
T3sKtXxx1b7e9o8dJKVyO9zFw2UuQ5JVgpLuLIAsv7E4eewPXpQGuXF6M5HuCG+xriN40TV4ludd
Zn4LMnQOJJqyz6hQWpYLO/LhukBPWSOq/YN9MQjQ6SoZmQaqBFNNd2CDt61+259bdoUHQHplYZcF
+9mlKYwXlj9Sv+2n0MeFU1igFY9mqHCQM8rDPUVB5Gg7KuDIvlXjU7bbJbjxl+zl2VyhJmfAt/16
LFON3IlbJKlm1bYwnnMVg4M/J3M/q9HSXkB0njK+vs7GmSPUcuizDrkyXGRifswrM5/lChptEdss
QZwhCSej8nJomHr9JHRV56a0KYAkjHc0gLmcXL3c154jwB0guCi1JdVGRaGtg/GY9xjeJeHLDgCz
IPAErc5OMp+4ho78Dubxo0gJO6I/pfJSO7ZonMEow5okMtrEW0dJfJIq4eVsJZcmvX8JwRu31YCh
815qY8fc/C/lh4rN3tZvyZrYMM2TSQVWqjpQB/62y64SPhUz8kthPuqYMq5LTKuJuky14Wmu8Kde
qsVRbdMuT6vTtr2qTfn79a0FhFAzPl75n4GwsjVLdvZ7876WTKK+55TjBkJ/6Rm0sdt+JrYz52V7
JGa8a+kIHvAOI5aqCjSpSlaJYMeolj+XjXLafAhJ0rwSAfie6qzgej/sI/b163aMYyd/aFieE8Pn
4dEOGwl9y5T0qf/bDLKzJ1/buVE6WWDFxBnwo6zmSbPo2bS11X1YaUOoyRXP+NEYMRMAEHO0l8B3
TdzssgcEl0zYmMEkbGYDKBQw9hJonkZ1WReM+c7jtYMdCtsUx8V23qJ4t9XuZuqG7yvxY55JLA1z
nQtD7XAZ+0/A1k7a7cv+vux1RHvlzmhM3u6i/bNA3hJ8bYgNzVAgQWXrWs2CzvZKG7E83KwPGAMm
hLSFUEIV2refDjdZblQKH0ChiS4T1HtaUF91IDlfjJBaLXnz6vZenrycTFmJ6ROo8sOFysqYQb8w
lgKGdI1iz/N0ECFUeBbHGMmNasmeyPOm7mHKO8EivzD45HLr5iECmiOD3vXOQn4LIpKniCYGEL+j
+jB2ntKE9raJmG5wMezW5Ma2W9RKLicVbV4UB6XdPH3urHUQTHjcuDrOJk3fbhaDwwFLk70uQa/S
ePHjhp/aCBqPRuxvLkuDJuSulSaufu6yQKEyu2+npKSuzr3L+68PS98wAtqjTkny8hjsFspYNEy9
XGD59eRS1RLWYWcAn2TzXwPU3kPFYQYCwrawtzZc6HIT5w94rN8i9i3KKGGBRhjXyy5lAhIOwHEb
e11Sa9jxIskoYMPGNqd1mAPSLede/MPbkRmKkMk98CJKxnUHLmQZKN103+8sVK7kgYYviFwq+xM9
C/L2mUMj8GUgtir75yW93L5ik9agTbipIW2BPWyVXPuyOqzeQNMapzRazKkT+7mG8Z1qHVnMmmOv
3m3Xixlx3TSnxEupxxkrQAAAIn7ZVDyLQfmsUVEAGQpXqm2wUoGrkjdZTZoMNawB4Brj4rEWbZId
ae6VlGeOqUomJD23R+DaZH5kPvoRKUcANbevGv4FrBAKKY6g/hkJsIg9G5mWKC0fuN7XdpgtjMPg
mCT22SHyZDig8GWinbQdiVNrsSp4iq5MurfJqmA26MLdKusHXBZkgU5g+Jl6+NvEPEZymJu2mGBX
KYFJpVaCQPsNoNcgpsXkA4MT8lYReTSWNb+5xBYOHUpy/W2Hu1r6gss99x5iswjavnTCwHi0cZVu
e0sedEPk1dZsI2BXFgwRHjVpIjAE3fzLt/9uMDW/YttDCPOiRl2zVFEv6x7itWOmuyo+QrLtQ12G
bs7I3G0LQq4XLrUzo9zqRaZyuFvak0l1UZhWNNqcLhIhPNp2i1SZmyw5z7SmZ5MbybeErmBVHcB3
swfNAUdlOX2j60EaC5GGTUBvj3oZoRzob+Dupy+dNzyU+MnSCz3BInTMjsP2oMPVc5yifBwzNSzD
/fslIylQS7GM/cFgz3HeLioqK+uGjfcS6fZbURgHVNughDbsEPEPFVg26gYyzAV1yIb4WTmyIsca
d9MKWcVZzyGfHotRal+btuctF3ksA6mqObaJ6UnUyS/topqStZGWHhiuzblYqYXn4Ohn/NGE1BkL
lVO4nHz3e2tnkSNEa47V4mn1iCOqBLSGrk4ciGu6XbtJEeNFGuT0HJzGwayQFyVt0cQdWc+WsChp
7EkdjvPWG0B00dOdaPzJaJ5VnyIolf2BUP74Z7LavtDBOqMTx6JoH9bCBk4xOE38iAn8QvwvIBNM
Ymgf71kUXkZa0WPFu1dVN9mk7tyPNfOyafuNfZKa5vV+ny+i6e1B+bAk9ObRXLByP82bmwYVw7iS
2p9igIpdWZbOMajviuaC3R3TXlYtmyKmRwkrp+nXPFMLmTrfWmvlpVRCPV8vaJmqnkHKAhM1CVsQ
PjQ7EDDKACd4+TX8j2VYDkwoD+ERrPMfqaiihE36TnPe48Kf/0qUL3NBLtLWewAUKtLqZGDTyLqd
b5wpEq14+SloTjNmJIoF2so/IpMfmfsZTWRh0xGCX7ApaYBQMIX3sQ8sMLodHNY5yQXfVOehHFPf
EanaC7EQaJ3o14tScbQw8hF4LH8f2JMrFpiaIsbBfX1sRP6RKuuRiF+FE+QEB8A7cPPx7HMMSKzb
SIi3/SvtGRAQJrnwExQHkudTOVMM915zt+lnHQtCibGgWY5pj27qEf2Ii8hbqQJ7EoA1ZDoeMeqf
2AZwsA9dTmuaiH7C6FCXmg/DJ/JPmFxPOwVcFM9f7YxY7OnsxFqTyh3lX16obrhdWZZgVZQDlaJV
W6zkm9FnS0LclE0Rt7DNMwK586q6NfRYZrRSzOaOIgvlDlq46+BvZ47c4MJjGnnqOciGhKckxB1c
dXqY4msVTM+7XPRTnho9Ujhvc71BJ8tk/MInxAULHET7stSsk7xHs0cwlzObYnIHbeD5QVKECYDf
lOUGROrRCoslTRTQf4GsWWTFtBzN1alYPCiOrvjdP+dHaH/cia7nWowRyyHE3s6MPR/mQt/5DzLV
68G5bUQr8K3EzulW2BVCiBk83QnbdNZkhb8gDmHakgRG1YI7hLVwBov05+6bITSosT2YARa7tfUi
dv/UL7X0NelnWqRUsw1u8Lp0drHcmiivVdjIpTbWXpUCDDT8XF6rWJHWTqe3Op+R52mXGDBEKxQe
O3tDyJf8gGsUatsN8+J4XwAcEvm8CUFlzNpyHTgFHaluSSeZDMvbgp4r5bQpiwTeWPaDa9j1YUAE
bbAOnMuAj5waJa5lVM30oSiHawLGgu7qOyTP+byBk0sCJ9Afdftp6H8PIi6Pno7Ve/kmzQMOrtjc
JwVdM1teCYvELAqhHRc/EXyIPYiMiscKOIwB6kkymEwwuU8OTtX7mkdjUi/AuYsMmNSm+25wLqYO
ug4GSBFUfbV5ggqXoXCas9EC5ccJmzM7dn4K2GN5p1V6FcmLEiaBC52iDKMOVLobM3UXGocViRx6
rCc1Dnr1g/uYekfiB+3OGvWuwl/gmVBjIFTMNpvYXYWg5eeXXdWvIwKCH8s1iHfz72mECoRB4CDa
xPXYPYBEX2/wxCnspCWC6Usm2pV8lnFfL+2hVIDGZ0GtcDujCYx/ls3TCZb9KGFj6e1NH+2I+K2G
xMTU7EExKC/xR+d+b1ZGTLtGa/n4sY2tTKSG7W5HhIcVz1O30qtE/dXgPmwcS2C7igDueuUiUjZX
JZEFPNhmDrO7Wph+2sMNjKyVu1ovqnU2LjLh8sTN6mW8+BzcrX1uWbHY4GoqoC7yy6zyq1QWLjgZ
PkeDbxIp4XK3/Nydb7bQdSkdLvh0CO4hlJ9e+lAfDqyNTW0VeV2L5vM=
`protect end_protected
