`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jNvGKMNtWEUNKagzcg2Z6WIUWv9gWJV7my4RvssH/ux/cX8RktigUyw+RYrzrXJGrNW7g1x/nBwF
74yzP41Y4A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cve4pj2EfLuhqfhnGnOz5iUJuIGWUldTY5TKWZtU1S3TPZ4r9ymlKXit4YnjR9S0JtAX1GoFuudL
h/jZOj05rTC9CmxzpO6a4qp621eKZhXdyOHyWMf8jPXE24P9V+aRttTL8nXifMfo/UFfsvRfUHHL
a0V7II16UbNY0z/aQ74=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FK+UvGaeunWTo0SP2EhgyPGTZaNb+A6fyrB0Pb4mabhgLBujusE/NHHToooQsIrVtG+iA4L6uoFa
xZk2qbFfIXLgeHkE73Jf9tkvOVSfNHKkwE4Tk/zJ3hux51whzpeHeM/jgYHXV/AGxAjK7wYmqNEp
cavJsaWgLnwe3yjG331MbcwzkmgERAfcBrC1i6iTT7oe42Z8bgt2QuADWtJa6+y6yzc95b43/J72
7JqV+DovmhlKbNR1biVaDlEMoR8wVeDr0xj6PecXn0O/DCkFw3POXJoaMT+xrRj1LksGsCY+qMlG
IfvdA3kKCxIRZxGcAPvET4wf6cGXK4CAVBa7IA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
z2wDansBNwtedB12HDIWNrI0jJ9Of4AnAAv+qKssr7e7NujivlJDkMFVu15DOLNgNtFvyO0niOHn
/kdDAjIwQtt+ugBkFsRzbHtzg25iwcWgxIDasTP9xLaasNHS5B2OfeSNk+sAZRujgTnv16OLLpuj
xCVg+ocyScQyJTN2fY0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dHaEE44368Lqz+gkjyTg7OMF1sLix1urvVlzCGNFKkIp5zxC5Hb5ei+82XYKqaRz661xkzrxnXIz
CLpQVXEZh1wM12r8fA1f5G/ZuHgSsoz7RWoNbHd4G2GQJUG7WVKCnogPJmbAQZpXthW3KW14NIsi
E34leEwjyTjx/frRrPczvVKGoZSH0tKOZiCD2ER5SRLpYvlTJUkcUEXx3CipAjm/wVGV6SSyQJeO
CTF45Rt8GOFQIMhL/GO7xMB3lpMvQg6M9+8i4GbdQOAk3MmCg7nCiIL/ptz2eDE+txQ7xQlXt4Cv
Iz7BX+6KUqHhfTCrqRi9bRB7HwJgifi1MzfmqA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
dBSVDAWiIsOQDtztSiCUKV2dJjLLY1u9cgJNvfNDnv0mQgMBDekawHMwokXMXnMEWx24JgeBeilB
9g51nehcuGcufqsah5rsE1KWunv7ggvSA8TUt/gj3LA/b0EWJ4nWQLOLqOQI+uxvS4A0ZKngETkK
33MXM2lg0rENmoKIgAkJAPOdMvhRlPeYcwMF/MrjW0hgZhles4NxqG8w2y8U6wkAbEWs3AnGhZWV
ZrQQokZXz5gagS4TAavFHsYwY2ZeiSnzfVeGFObWMgrMzRbcBXiHPfcWOAEHoTRTEj6P1iOgJt6L
5JC+0dp5WrgjnUjb567Z9nwMi7qLQPrXaGxUUE6i7LCRwKcGIe8G+oRC+YSaJtLU6+Lh5g32KDde
bkw/JpLxaxIRgtWTDivpGYXfdcPgF2XoqNaICD0kEXc7difRN3S1t03f8msW1b+vOX9DqJj4ScNq
SdFKnKKFdw6GRwhN8/JNMA0Atg5ANj/ke9iBdn7AdAJWXPvpqX5Rl8ys6+hRuv5ru+DygnMPozx1
v179i8ggwmLHnkHFNvPGpVbYLweqdwVxr31+BpDjXRccxy3BH9hogti4KMpASx0+Pg5QuW2mL0D0
0uIM+/x5Q7N8VLpofNbjDGtpdycFVwKRjD8UTI9r1pQtURIwYNiVTJ75Bqhg39zu4p7CEwqtOGPZ
9B8YbjVIgFpzkoBpYPMHP/mA34N2eoLVJbKg6reZ6miylwEUcpN+vT4PlE9mWti5Z2SxmTIRL9Zd
+TuoaxLKnDtCdvlfVHnlyzzU++NOOGkj80ifmVgVvzTyrMMmasn/ZI2zXm4FhM7GlaUHDxiOuAWx
aPem7DiZ96Vaca87FfFdgNugv+WL81bFrpmRB8aUHH7+88LNSIjv7jy+Tna/fAxrdN2ycv+9Ud9k
xdFY8rgGJw6bL66ctYEcx6cliZrx14K6sK68ktfV9troDkruzcinfFluLCZpDP3c7YMcTzgEHBYw
mWBMYppzM5nCpqII0XWufTACKjQSq8pOg6G8yZjoHFk4RUh2myWr1rgg+1sC011ex93DoMAWktiU
MjkXpK3aTixnqbhtNMSAcuOVx0efIFErt+HUpKNGlDZEjTeiRhX2KticOaMQ29uIaXG0QGHr+Rvm
WUjopP+WNqfpk3L+32y6MXaOOmddtLalXBmkNH7v0rEYZdcOhxIg3TpkUqq7/6ciz90t50zqD6DW
zCKQgFlecNsEDQ3SmaP14an7Ip6GmWZW6CJpsvDcxvsfvwpCWjGwDRHjkZwTYwj/XUMn49UVkAIf
TaeEphGAN/aTr5G/ZeViSMbyVzg+7LmKZx8zRoCKfNeVRpahmGCodPte+DEh74Pgykqxx2Coq7JQ
efAl3pdrmMQNVGasE7ijFGvyl9fy4vg0p36r9hIcTuhVEEGzySLOg3ZMIjSrtjTnSXKGL5Sqa/Nf
FFPMfCxqwlM6vn8/s3VCgEAO/KKwmHyjU6FoIL4oOWvTEFm7oi/sY+aRKY+khxpt4Z2V6oiNxVYL
P1QRqB+ZUItNW73TOvPkbm/Q8ECrWHAM0/KsYeBBxTf9W+USUmoR9GXGXAl/Mpjg2yW9sAoTzZEh
DWHSvwp/UhoGCR7C+BOWm4B1UqC3ZNAObYIjlYYe7TAYKaZ0HUBCtwQlpm545vGNiBynz91vIlY6
47KIkI/DjDgXb3qlAtLsbKgetTUnkIrB/HGKfAZb1kwDFYlE65ZSqLZqnUhwGsEn/MFj7ij0KC7T
CgbDAwSEkzxN/UENPnBIc4qR/KCxUJalcbrgWrGlXcWlFfNxjmGEif8Ehj2ITajymg9SmnBd6nxf
opxJQ1BJeIHJEL3K6LVxOH3/yQYZOMlA62HB3dw8wo7RFWd5PTRXSTSmq7TEJiH8g2wevOvp9Z5j
ptpo5M+cZoBlRA0xYgCbUFveG1ry/L8SDTYwBDGt8gdwIlopumxEusSY3jXS1uIQiIIAwjANsCul
CLPvJ9rzr7VV+DtNdE26kiKTib/5lMqcZUHOgerDaBVw280cPDeXGmYDeYxXLYUrjhhsZlb66Npz
ywS1S+b95rAIst58ZZ+DIJLjAC9UYzx+/3YCtq5xT00hWjuzm5BEvzI+MpnTHisw7pkgb08kiIi7
iQeYuRzg0uw+qYvdx1/k9+4/knYZN5db/A5RwJgjPWhAztEXkGfRu9Rv2CRTgNY3S3OnK08mjTUQ
iPHoJiC86JcvrHpkswP3n43aTeAmBV7EMqHrVO46ayw5aoDWKiXV81+uX3MOSB72wn/XwM3AzEej
6V1SBFQnsOP2Hf3Hvh8Op/+It3cMhpEXP6Asm4cm6GzbG9Et4ZgscTKOANGRMFuMG0x6KfGjiIuv
Sn7728ZpAp4kaZ332N7Qbss3M9VEO0xTYO8/3hywTqsnPTjOs1/d0g5N39Au6lvYs1nnHhegLB//
/SHh4NpkdYwvxYzRZcW9V6qvJcXdRrUX4sKx8/1bIATR7CcCNF/xVEs9ftMTGc5kxja3i9PCHuNu
GLjhs/odTD0CMDt4zOaS5BIRgs8XDFLitKBOfiqg+7IfFg9rULvYqxvz7D6boIO+XtZ//hx0IkZG
+Iq8zIRUE8UzEp9JKadidU+3NRNuIWtsq6Aa+2qzua2PpChJESy5ynl2TttIFi5hdWmR7fnWfJNH
W2NgySKMeikjrTonXf+IPq6o0Bx0lbwbzvRKBC2Hsoz0i5z3xbtiaUAfVsn8teBXw/M7GmawMe7h
3yMMPyUVXNh/ywP/0D6Hm9BFupEKPpwxULeb9P8UpkXJnGAqcr/uqFIbYS7RN/nw6PtrHvajt49A
k+0yeSMRNn8xga85EtMrbY5L3VirbEst2KVSYEnagR03+uLhkSvZKzyf4+3I+m5k2oomewsW0UxX
DPMp6ELYLTuIbVFOQ9hFOD0BQQKze4e/Pes1v/RRn/mAWYtNfjk++zMEwrCtu9WHJaIPZQhjx4pe
whamcF4jh1eIAKXQusMtV2nH25LFrFdWjpdQcbMEmSXfcY7cqmYsKQippYmmGl70HNOhUKci/sKd
2ELxsCKGEABbDx0hMfyrHlB92cLyJ8ZxECeAh3eEfEA6nTECc64t48/rvl5H1FERDwk9IX582bdj
lxvveOUwm6V1GMXaw0y3UWlDLPQ/QCT+Xsq3jw9WhOQFSFLRh4cq9+3dWEjdH9wZbRgexDU9/u+U
wAcyQnHcfJDfch/WLIfeqQOeM+p3IGY2AfAWm5NotAybSr2eUQ6XxDNkCUEHk3K+7VrHgDW8ckEM
G8Tq37rAFsByHzbN2ejBI5iQlcyWL6M1yvQankGD7AW29LyRWWYr1pVNCjWWtJzHPkEkcJLPGcZ+
ReQ1LyS3fwretzAehroAlSMeGwJDY601aeaYqWQ5332xXGodeYdcIYvvROkoqc8k884NBRQzcWDd
aCJ6788Lejn/XAXZgqDYMm7hggMZIN7qL2KtRjCwQxldv5WIcuUwJozBev1BDBDbfyaVR2tmSz7o
mCfIfYmtKhlScmIebOa6IXr2JjEIS1hJXAWlEp6TSbs+DislQD+3XqG9YMqYjNuk5Xq0ZwsIjvBQ
V2Xw/+bm0vcfHawBccuACan0+LHme0e6E0MSfUAsckoNdEW89p9ZlBGaPZZGREa+4FV4v1wyg/q5
L9IQ5FZixwt1sVbTV5byrZagYI8gjhWu7jO4pu4rJnRx8KQ2g84SnHtppPj7pI7EpCLieNMbw3Kq
rIbULLCPHeofcNARoDH6o3ZNxAjaMfslzH/u9WLtxJNTdq9/uujcvZ4AV/llwumov0blhnd487mP
2RPKVUeB/L7IJqZ9a3FPB/rlfRrOiXjsew94/eLPLlbywqMtKyBt/YFZ6vhuckVbrvtr/kSevNQa
lQT0HGXvz6+gHJR8q5qC7j0K2hyP0RmlL19uJsENeXDhspolknqMvUEZj43So/B1uA8qwkKOOsuT
hcDvt0zbMioV540Symwxjr2rqBPLxR535hMuPCFOrelGWUpTBifI+h6ev0TuMbdVAkdOMXThiz9n
SeXujYI+z4Y/YV44EgKdOcLbpys3VcWhVmeGdke7ogLMKql1HAj8t+sfHdmU/xhpjk6gK49hz3f9
v5OdjWz1da+tyNPXjdSiWFwUaBV3IWxuCsYkoUx2xB4ImLAwURLindNBu6dQ4SOUTAnfKKnmw4A8
PyQRXl+Asbj2YxUt8XjhvVJ6T6QUNJPokuW1WKXc4AaJH2HR6emAL8xmQaCjbB0GogxEeA2rZPMD
YBN1LnsrzW+PK/LwRDkYS40QGQWjHF3gYUHF5OafKD7eO9N08YCX+WbkAbv6TCmY25p+fKJ/V/qK
VjvKY2g5pSeZkluUWDX6y2VyoxXmePOJFeCDK/T0NavnprgWGpSjQFUC9LdkWh/BI2qAb6SrHeGb
vi38cpD3ImXpj3PmOA5JFObHNKq4yzy6ge1ZtH+2KjGnLQaApjmxLsrnSjWMrg27saUw3GQEXQuD
Mv7R8MMx0wI4mR0k3r4/QiIp9ebActiHvRYOIWl+4hs6i4TK6FhAU0PFJnVM1dnm8RcOvRNbcREd
f55RHg42DOWWChoPJW0mWtEJsTvUTbjDc57uQERQEMM6EUCVSl2b8Ngml3GsRW+7LH5h5mpM3+ha
EOmFIZupg5gAbpFFQ7bt80j4umZr4MN2uiU7/1o+7LcWo7StFlEU0X6z3wAa8q7sM3ZXQ0gTWwUP
PJ5Yoj61CIGnKwOvPKP9w1EN61c8RG0lHA8WCEiUvWc0PazPTIG4oD0riKVfONX5BYazVfx0kzAi
uemc1fC4sZLQlXypJ+ubZMca3r5CiN370v+sdwg8Acx6c/LpVXHsI4PQpIQLOyD3f7OqAjvlTQMd
ZVVC8nl58VzLwDuqDhFGfH8spmTAe1SGswqjg2Cgue3+NQWhHllzytZX9/o7hw6B8prC6rk8baob
7ozNGi1vPknCqVKxYZ3ARrPIhLf5p7E9Y4Lptb1RvIxyLM/SpA690TgMFH0bok+fCN/b8GeBH9eB
1jv8y6l+KuC59Uxs6I2NVNiw1c0J7l1zLOgtFbo2xTFpzWOYnedTbfS5kapKtE8ICm2wE6mTvDBb
DIriAG+FJnmyG2Xxuaw/zOhkArj1
`protect end_protected
