`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9584)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosb+EqZ1v3SQM5cugroTK0Ogv/nKwWu
IP3dGkUeW4FH+9YU+CCo0CN+uO6kZ4slP0LVtqG+59ekLqaba1VneiaBEjGRt1Gz97p/C1ncB81D
lvqjp/OeO71QSqf2Zhay4ZYl2tiy+Ew1f0ZkW47vQINNdKO/M0B4+2Kd2b2OwA5iNh4jb38Q8o3K
fFSQL5clNodY1kdOeu5Xj6KBtyhTrCkKd8EBaxyft3gKcQzAMEwlBsVzPJE9l2mlj4L2hrNPkABv
Ey4sFxsQjZkD60tKlLvbPKVAXxUC/ibnMo82RwaOmGntqxcgNzstz3DH5w3wJZC7d51S/N/EV+hA
Xo50eitxzlUoU6NgzTzFdMOd0hQyDs4xoDhfpDzKkPk/pZSGACtZDHWsUA5j0cJvzcNhSq5PURNS
oWlrEAGpsNEhb08y6QbwiNynOnWHVaeGfQ4oA18C9D8nM0KOum0AeD1wl4dIXpy5biqf1NbACamC
7BbNdkGdHLVVr1euBdu0AFCauwjDRmEmFd8DNfP3w0k+/I14hl+vXnvbfLEut928JCFmpOyzX1HD
0DJHqCTni4867HcbmIrobdDD9zg6EncF9uqDnLxtBseSwOHARwohapsDbgBXsJw27r+6C7vuOCkh
CDNl6aG+lNb4Xh4SFYi5mY9v0FzbNTWOE24I470qgSQ/vA6WvHyiL6M/4IqKP54VZ57lSbTSc+QP
6QhdMn2KHFp/EbigDabmmcsc2mnSDCF4qe8HS8lMna4VW/p5vvd9OSLJdUKetkBxysypKgKI8tbj
cqn00WVBuVreOaGPga/Erb6GNmpmLMfylBRVIM/9aO2cben6hKfDiuGzl4d76tGXc6O/JHLYlzTU
M/hGz3zrzHt4M8BaJ1a8HOSFP4Cnaz0QqVP9V5wNAqol7GhNKQEV8rUUqgHLSrlPfa42b2R52a6Q
1+hU/YUd7f65R1HyLivViwcEYYbgEnjJYPQeGco1wmaTk5lbXhgXUhYniNu66AlV7QTmTf97wWlb
xYXvcOqWRyDpE3hPAoMuDPm2oLr7TMmZOdBSrvHUNhmes9dcwd4HW1uQWofsRCzX0waBngNo/bOE
h2S9P45ofwHkZM+2Y/2wchH2/XEVgQY7z+7Bu3IH7rS7/JNNjMpx13702mc2moGYhQ62kISWCJR6
6WP2zGUQBhxExSAGFddc/QFM5eFKOcXXXyNaF5b3dfN3Ks7T3nb1jOdmxzyIHKX1bQCaj0DzHGc1
wY2fcdQO9GGbWcEjZ0/ceSQ5lTi+JRAE76fY5JcJWq+6VUb6tPhDtlEE/lPOVKaNwdjtNgxegiWj
UTAKY1sy2Gtw6caKfWhV3RHUe5Ei3Cz7AE3xJa60j9EBxiWpZJRXnfGE8h2D9mv3nYE0MiucLQSj
0zb15WyD+3I+9bw8xiET/IyuqQ9DsYqI3c/CcdDVUwjStPbOekw2bnVJTz6iaqLgSxMLMElyvZgp
B9tRFMH+xek1on8c2rSmw8EWVXKeNhZLWZazTfguWla1DjRPkjGIHFyG79Odplhkg+aeoHQgEzX5
oYKPHM6eItFc13ukqdgnUdo/grPtEQKQwTIifpe/Hmz0NJeisnwj9j/qeZ4G2FhgCQvHHEAvG7d0
XaEINyabHUUD0n+Ko5dvpJZQxEc5GiCTLrn/NcrEVRO6VU4+E/WZh/IJoU5a/YRn8EETOiYftmDP
q7WJm6peGzn6UqVGc22wzX8ERs7XQHLTPUSamX8VTX+vGNFOL2dTPQrJ3Xbyg686yVAoGvECuTj0
DlGyLrTwYlk40tFfmZ1D6oo055BBBHgXstHJ//ZnHlun8bp0/tNW45FNONuwRYC4VfoxuqQ/Dzfd
hc51nxtiIsJsyvSTXgRLFnfj28xYiTyGX84W9BWh5Ps42kym+2v7qpbK+xKOyNMdgr7ziYlXbsW6
2d7xFCVe1Sfe+dZkTdEE3sRc/uBbrWwDsPJNdvbjT4LK4fsG+tptA8KP2UBmHxa0uS+XxnFZNDuA
yRgKCUbMjAp74mXjC0OQkmOL0WoDXicw9dgEMGzdYmpUSxMWdUubMc1jRv7GvBmZfALoALO+pjGv
PiFZ76B5wsbhEzngLgKGAlK1ar7Jdw5tWCdCClROxydqPoa3MvMq58fE4YFjjwZ5LjAT3VG/npdF
pYL3yWYs2d2kaN6khyEX+oP/YpFLyuFLZ3ctsMdyoe3DVwDxO/0Ek61P8UIvfQCyMTUZEfnKUCoR
rP2/0c8d5R6JU6vCBqUXJbyGiSw/RyhEcc47D+FsvhSCi0YDLGqJtlxJ9xTzT9VsUtRoXmEyGjny
YkUFTRNV16V7QqCJ258lN3ubIJUE311aR9kHaMzMR6DdPK40q0eSFpMYJhwJOgyxOp8RrGxOrNhV
AmiFwARwn8T93wEZBX/BiJ1YnzN6G9c2oKDgWjb512o4S4ZSw2+KaJXiCnsYMwu4wgqIgAFyy4yL
xY8s7NfHOAeefElDl98Gs5qJfHtDMY14Lgp2iY2kBXHgYRFpBss8aZivWgSU0cEJCt9uu2pK923c
Lpax+Ml/ZmlybhnsMRpQCWPlDZP9dw8/h34W++SdBPLheSc/URpbhknYToBHoRitb21gyxMRjyka
qz2va2WOPsHtfSSByI+bmXiNF+0upGvTIG1QWJdLYVDjlRC5wq/DqxBf460tlRmLZgvmMTCDPG9K
yHQD7jvAk272SopJ3zvtTudkIas60Nw19aTkyFHHIbY0stPj2v+d1e8xMb286FbvZ3ci6vIxAECO
xXylu8f8DqGXx8VP8tuP5cWVPeSgp57SSp0li5orPHkDU1uPkh8Ojb2vYVnJBG5hm4plPto4g41j
+u0f2+vLeL4y07C4THqC5onWzm9xawyHqPoEsC+2orr4r8VlFLLplWbQIOxPnFyjZO87eP83E6xC
hSMZgfM7ZZx5bgjqxsugmyNNscodyt9vNKZq+eYaNwxw1S+ub5v8+LLJLKmUZq+zLo5jn5uQL1XM
7AFAR09pMz2bXbXpaANxUU/yAY+w2A8SvmE/Rd6N0CCEZmAGZfUF4zTws4u41LsmhKsz7n+XILYV
P1l6VEUqat/vRgoKkGzVMKPrr5Nb+s/ebAWZpHLvL5h8LhKkMXO1Kvt+YU+qW3lt5z9eQBpShLFB
BkMssXSUd26WPo05aBlP3bXrmP4mgXUtJr60MHy8H8/5HP+EErxNVVk8rE3db3RVJ6GKMGk3jrPw
MdroEAR/fjpOzaqAJ3FQt/6s/BupB+wWy7SxXwkOhyCb5u1zY3BZ9M1Cg7rZI0v6yXaigFznFg4F
NqwyHvKrcj+7j/Yhwd824VOv3FOHgNWHRuDGqTZv9tvyU17lZppgSUqO3pzf2aRSYqlXwzOJrMb/
kCaF6QEHDBiJ0DdOXWqmtNr++HyUch5tEfvLujgkJcCYqzHbORt8zauuOJmdMDg+lcYlcfkYbngL
ToRQADSSnzCoiTbImBu5jHnnJQwxkaWpS3RiAXQWLM7/tGo4Hlw6yLakFev0MLisT1Wf5Z2jIuXW
Ldk+oL/CWQgSowySEtwWg+V1jz/Szy3Am1LQjltmUtCyXHwzFHjtX6B6NFlhZeEJTXs/cGS6znwu
vajyeZa/NXrjDOPopN6WHJyIOe5rsRkh2rR30djquWZTeMWh5KF3HroTAJ24Z2SGUdmpafpmbcfS
K4xExpbYfkm3rcH9lQchl10c4+C9+wuT+dV95w2ASIWU56FPOEzwrvmsXfImCHQ0cFyNLXfQVoKw
DJ3w8jHzx9sYvvY6OHsx4SlolPqIdff3SwOI/IuI22hJyylxOTk9ipfKtsfS4rAvuAQmG/rqjPW+
ARnoOxoBUrhJaKDJPPE9vB/rJpLSL0oN0lyP2hwatxV+2QuhKaVwUL9x890wojuUWfLDOaJ9z0tc
5EPJdkWTAF6ujidJjZxf5pns+VwvH+ilRNacnRLmApwBbwVuwINdpf2uOBseQ1lU5CNfr/E0jf/b
1b3bH4jl38JANj7sGBGAL0JmQvpTEYTgYJTnpNmS/1Fy7LxvR8jsacL/r+WBpxIGWI1V9X8OiF2P
g6PmiIRVWsfD6DkzIxwWobcpqUJGTvZ4EAvT1fNFMDYeZ4apKkJc8blbEBVXnu7Mc0xpTzucLc8c
32Yc8SOxNc8RuDMbPycsIWFctkHZzBNC30sFiNtqY3yu0OtuHnlOnXlmwH33DaN4pChCLYdDNzXK
aMSjvlq96Kj36URDSwO9vT4X3vKWx3Lw0BR/p0ofIZnpdGXHDrys5pNUXxuM9HN2bwD7oQcAoWpW
IwfAcb2L7CBVhLnk/15+PRJ4h2+UmgCHyBw16GvetUfEpct6vjkBdwQ43jKLOabgBGwkv/PJDNGj
XE3EhWiNXCd6gy4xQuIdpV2i94isPb3yWdj2Vm4eaDOQa13ZxKJPdS4W7SZbyNxYrFR3FeIRTZt5
ZyzJIHLV39Jh8RuJBp+pqsqaPD5667Oe3tx3O2brWR+xNpMmc7hG/Y2MZwFwgxzRtJY/+uNMVVC5
pk+0RRYLFrlYGgKR2Ru97+Wn5UPeKF4U+twBqTmKQz4++/y1wWk9W5bt2/mKFH5SElcnH9pn+Ivq
eIKj5i39vekW3+ZxyMSbEG5H2v0ZWqUaoJ7P1Xe+S9lIrbmh/DSOutpVO6lpSEMdiMxdnQO1+1jb
fWzG1xPr/Ca5l1L/x462BsBxHYM9UEDg63r4O+sopWud809c3EztmW7APau0DOjJis5JnnYp+XbU
dn6T6XgpVlMaTIop0uNBMHe1fZBUYbo9wdWtz8iRWI+zlYVlJsZG+FRO7Yslu7wc6X1CTm9DUNP5
E2Eq6X7/iys9bwFXraIHKpQgURCVOUMoTIox9N9F45/7ToSoJwnF+TOW0iiNV9OfHlHMo8OFMYUZ
H0Iq3ioMH0ua0JXTiJGQC804lZV++1BDhGIXogSoVE4iquY+34qp7lela9MYJmNm+e1eoBhSrEF6
PT6mhrmosd56KruiVrLCy/NOlWOpklOz6I+33uwGSa5iMORb3qfar9DH5Ts+6sCCec1Q/ozh2CJi
/8v0LiRysLhT9GhQgsp+fYmRjxaE19RDDhzU/ufWR/dQGA39L30RT53Pz4nYNVYxk8VLgxyO4bI7
1D9SFmN6k45c5Qz/I4jkHOgG4gWCKReMJUIaDk3a8ZIjBNanFhlnyqYoy/xr03MubEIRuPu3V/6O
AemreFG1bVLkCQT8mBkge00CwCr8yDPEuggyuvfBYiFsRw+Wk1LjyIbY/j1g54ar/W4WpmSp3Oe/
nZSwpzrg2mGKFk0WxPElDMGyy58dasN52k+5BDTH15TrVZ3y5hDuObdNnE/rzH9+RL53Q2xoteS6
Ao6m563H2F3FfooK8SQrWOOH5Uf2KuthmmyXWNeeWUtearodalzzl6v7slvNzwIxVdAzs8wG+/Nj
9fqOhkt7OiQQxyOA89O4T1UMDKztNHDow5o5HMsocJ/XWLfzqWrn/53py1wfk6vyW7OuGtNPbcOP
42GDMBYwx+zJPntHQNgiXYVtvWHNipRgBdwOhiDPtETZIhwbrLnzTvpFoS8FMRtSNdmAxzkCOYiB
u+/+i6NtUZ/ZrudKmNP1BYpp3mk9c4ZjnMSowGcGqujI3HCIoAujaG3Kwg8485Lq/UGD3hVbvHgL
aFPyAN3I6HI/X51vcjPnSWnbbXCNWtVXO7NQvLIlDLmN3gn3l78uChguGfWaBngbrBO5GAq84cSi
ZZ1raXEpZdQ4mE72akF9ALgG/3wH86ofRgWR0ZQR5JP5NKmJ3TcdNsCeNJxBGY9l19u1zpmO94eR
O6XZwuVC77ftoK51RDORV4LDMeJatfVxNr40hTIeCG2I+Cr8fx3usN4g1rCp7oHBSUzMq7IByHg2
RRjJ0KcOfhhFLLU0Lxn1c43x0uFHSy5iE3Vic4Rtp3j9M3jloBG7U2O7R4VUKcRLoCoDuoTUgdfD
/jvdI+C6zhBjB67j6aKxFKX60iPtXIdqo6zA/bCYvxSjY7nLJMPGe78Ka6OuXQKC5USTkv40WH6z
Tsf9tqlsC40E1/Rgnt5dSxpBnsM684RU+Czbj2Ph6pIRnFHxix/INu1PUGAif1pda7FbdkvkMP8B
Yv2layYu5/IqGoQltICHdj4r9MZjVyxMM05zscIrjAwZu0tsg7N3s559EoeTBhbgk7aBd+BgJDUb
t9oHVxEWHBgYDIvXL8IqieV+8EE6kp1oJIMvLkfG5UWxxlChKQDq0kP0tsCiRrWfgtWzNMmGmUyt
MGYKJi+8Kge7CJ6/VE8gbQfKYXkZ9/R/rAkJg/RMjWgIab6vZ/xA+v4q2wEgBLZYh7yzukfakOjv
Wb0b4cJfZ3ghWIEm3pvP8a6tpdWvV5N7YHaDw5MoaSFtyH0MiHQ/hyMQw9Wkx70KGTE6LvQ2TvqN
zSed1zml7qpczoUn2s6vIZ8Ih0cV2+ZxKfwu4MGypsd2ea4JsoMVh0KJV1QmMO3w2lJ/n3PLRu/c
VuoNtz/nIBTKIuZonpy7c4p+9hQYCbNzilOKo9dPDoxZmfn/hnw1XicGxr4m1ZmsRx1dFn30uasV
XBi1pLfQ66LYwCILMzk0vaiCp0qBbhUd8tCfV9f8ukXRUPRb38CYHzxbcBLzRt4YBYTjjhRm3tOH
lQLGCCzXQuh/0cvbzi5of5PXzpQGSFCMNBF/p43+bqHbVQVub3FyRldOZ6GlJVWaOF0ogjQyfGJ3
EychoI8EYba2+C7KmS3ODGm9k+q6FOyFXefRLe/KMpMRxH7pEdjKMFqRiZNxRMDrHG2LJNg66SCD
lY9bODL2EBLdddM8pJqf2Zg8Z1ZX9b/Qsa2bBhPMjAXpe+DjuxziC5JS2aJAkNajQ6ityPQCyZhU
uN94MmF6eaGEIGB1fVQyOFKEwBgWQjaXlOD+e7g1NhSALFalV05FBIrqqbsVj+yadQ/DHYB3xmTi
sMYCUzhU0utfi0XCE0QxeYJyIRhrPMPgD49YGzSzV0hgLqJyeHLOZGkSUGZZDq4NU9UCaqHy4OjK
Np0o+drzIEMI0I0bWY4Xa0r3bs6IWJWolQ/RloLDYdLlVh5kKDEWVsK02JFMSVDW+56jNy1zJ7yp
d8Q2FmSpA5DuustSvUKzUIqd0Lthihkgg0cazPXjnCp+3kEkFVce+9/GJXMQJfKLGT9UMl66SZql
mVy/b2m7BZCQoY3XE3v8uPyqE4WTqDE+4bmcseraxrLSD7mFJPKuBDlVrwxj09P4Olt1yjVpnWdd
ohP538S2JDa9wKWEAdsj7Boo0IyWn0Mjaz+PP5pLb+g93f450BOh5M6J5bXvSgI5iUNHtfkUSTEE
bmkE+aXexC4OkAXrkQLTU3Vl/oMpdHKje6In31VFp4e2heZi4KkfqvSHd6OZ0GSJ1idovLu9ApPl
6SGyb9WXtJDObtR793wPghuKpEhDObfdY0xXI1runDKObAyMK/zj/SMTuJ2Y9yJufd7j5pjFkHWq
ysLQ07Kb7C0dHiFixrBQIX0N///rq2+lG3qUVrDmVpY/tj/YT3zlvi6mHe/txnLMxt2rPBr67Z3d
XoOgrFLfdkLVbU5xZPtXMfxhc2OX76IQG93+ik/rq4K7CBSFiRcvhihFq2bgJEGqj6sZj9y5crh/
GQYRDeYsu69UzjTHKxaO8UCBbUl2Hdxxaz2mDKSeeeEwmKJ5dpcQed/PrEgV34ILZ1Ed0gd2NeX2
dOZc5Gx1LPyu74TJ/DnGakyegcs5VsSyaLDWG6RbQqMaf4r2MUd4Sq9JUuhHbhS+37xZLVSF1m9c
8EEn1SREEhOWseg1V1KZFZ057ffD2VnSYsmN2lrtK668ZokEOYpr9vzZa1YnZctYxQalHq0dvXGh
Fy6nEH+pIyb63ogDcmJdte2Zcdlqc8hityH7hUjYTz/3r8U1B3r8g7s6VB1IOzgepnpZX1N9CMe+
enZD6NjLw5IEnXVAKeTYvHCKMncNsTsuGth59BZQeklPV+5lBbIfenCrviN0yue+RcxrIKrbMs0a
kGIp2ODSDaZ1fpdxH792Hg1lV2O1vKWMTXVDGDtso7ZhlhDx7qdvAl3E5lTf5OR+hFrBFWSMkGye
IV5l9JRlLYoljWOss4LMTinz7COGASFhWCBJxDMWrjOzNvVd/UPPjpPvXztuBEn+F5H7Y+TWJ9fc
Uwd4ciBvZP8qnWNRjZoWbCIEjYR88B+DlmYWnBiP7ZujZFlapILfz6fwuW79a96wM0BmgBNhX4sV
Ge+kGGnFCP3zGdKPBa4rz1EBsSm0+VOILu3II4vtDHwUPG2Ip01aLlRUNDS7DQm7AEQr4ovhqVxR
hDH+OUPo+8USczX/q2ZybzUz6lTSSy+iv90vqv2t0Lxyj+S2MLHkY70+1MFLwcNga4yUfupryLuG
+98VKNplnmp249pD5xmnMn6MH8EQG+Pxjk7TCwd8fwIWT/QtRdA8i06TyaGhTo5BLWFUe6emvVzC
7UpihL1dSd+XIXPUBWEGPP7O4fU6beYvMkUJQidQu7rBktSycZKJFP7sJqtJFoOrPJyJ2VTSm/xF
9iBB1TJn6N+QRJn3kZIpRskFhwoaGkteaJAMdjRsbAOBHtGr9qevaHb8PO18zXHaM7aINtsSrfRq
1S3X8QA+jF+nIL7fcNowOUbT/MXqy4R1vZRX1VEd0uHAlAxmZkqX4HMCpCEMTCWP5ntnuW9XlYL2
Er1zq/e67Tzw2ErWBoVkKdbV/VEGnaY06UrGErxBeBR1TN30OCwT4//bzAzbB+E9CI6/0ujCa5Wm
axLR/6tpVVSRy/0emrhWDbUXXFijhsZEqAW03VH9poTe43G9hUhNzyur0pvWUdkhDOBQzLuwGzlp
NySxQMMQJwn/BQcTNiSlADG9K3yexhxaf06MzYtqczC1W6e8H8QaMJOSlnEGqvHrY7aWbz5bSQb8
25ageL0s1undOb8566KtBJdwWy4IJhA85w9xqIdFNGkzn8/yN/NnUYKwtGQC+IKNotfE7dzseaTx
I1m7riITgZ5NMCJRvdKwIvABbtHIfAG4rLHCcRb7mv/Q7AuvTZ36gRzKbre2SaWlJRv7htIBOloa
blZVesrU3Llbw8UIa1l53H6Nv2Bj3E9Fv2qtwjG273L4AwCdXk/rLSa8x/X7NfljyLyEup5dtJdl
jSB3PLpXHo/AJECMs4VPVu5DJEHIltPAYvMhxP72LLVK+9ULdhVQIaOMoA5eYdsFBj/WYXsRQeE0
Kw3SpzoYA4F1pJ43dpSEuTaAWu23Lt0AZgz3WdSd6WBmGjo2KOFWXEfnCdz3TmH9nAFbjgVQZbyD
FwvQxfHm76y/D1sR2ZcWPoUOQ67b8eB/rWIVpVKD78Pbl1kwRZtoyJ7eK8MNBVKate9Inzo7kDPf
dCFTPfx88Qk=
`protect end_protected
