`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51616)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aPkk/LZprZljgyNzZTGF6gcxBz
LkEl/7f+3dcASD/i/KiDJHjoLg/SYtHgqFn8AoZY55gFdMJJA8JI90uFDulIUqGvbwJZIByx+L/S
+bV4MXjniE+bWCtR2EfhrkDBTkO7weLZkMnASeMwFX/46+VACoaw7QJ8FiJ2l9sd5rvxYGk7fWAL
JNQJir4zqZlhNlKXQDctEgXQW9tx2Pu9L3U+KSLj8dxraSVN4CizjQT+IhrhLs8bZ223nkoBdJC9
Jc8f60ukG24sT+BDrQ7K75B1IJ5oC3VEf2xy9ACnnAZwj+Jf9l1B/AUheJbjZlHGrfnjmvBF491a
CGNHjpBcNHhosvT6r7rs6ndLJz2KDlR/ULp+6xA2A3XYM9m3FzCNqiFh3kURxovd3II5ebv5c4Ua
5XfKy8+ZMtKk2H2hJo3QcocHnS0dbN1hso6EAhZO/0OBxA66LOuONoR6ZZnI2PqJmvar26nYq2sN
Vs8bXH7IF7H7E/EhLXAvFDIlqEBodPMhlDvqYR3fnxqQhkynK+WMtFtuIkpwkrkTwUNzrg8OaC7w
rzl4P2CSPCwfg0kOpcDKYwTiwrAaT71bHpslPIkUciPZT3YeazAJE4XAgnRGY0vSMPfEOeqPATPG
Z0zRSj4u2qSXA21CvrmOXbuRWkBpHWmnSQSNmJMXKaORWE0SXZ9+a5l1cD/mmTTQP8yDNEls1vqn
92irx/X/5UQADwS39EH+MuIYE4LEXNP47aldg8NeJtkU3sNKWXwM1uP8km8+cWGlizlXoKbr75Gu
W4TtlJRr4fUFW3lmBwE5keAT/JO0Zt9XUsmD14Soj5RsIUshSKm2e6erFLAmc8JdPgDtyxztsQE4
hkRQNCuCKmKGKN7oz/Vjpvs9mLC16IEtHlw65JSyktUS3+8GRi/Gvi56v67xqIpYihmqCe+bFgQX
nbDFHuTQSC4A/cVl37s5bE77yGvyoI7ywdpJ6koqpjYarbbGC2s0e/jUzfPRF0bMqjHjGs7k++2r
lQp9iybwYo4l9Jt4sPm8RWU11/GVRm763pFCPZ/t2PC7UWt/Sa2DYVMsRwoxGT4TX2drFDkjIp5o
0qOXq3jLYUTeNiN7PRFosocYunfB7RAQawboLkaMqiMZMs6ID1d7VwBXk/Di0r7DoUxD7ysMc0h6
xOuxgzKm2NvC5xdxSB2Bj1BtdmcV1VjSfndC7VedKMB/GwGGf7gV/2IUXuN4soqpO/Jbgf8NU1BX
ERCGsISsrZl3dAYu4JnRq5B2J5EZ9puY7+twmHxKSeHibtp3oS9VdF/o4p2c101Fnsln9far6Ot2
oD5HR1wb9ySy7f0CHbCUrSGLfIbgK6yAE9GiByrF/9CuCg1sswvLIZvOI2mnuVg79UpbbvqgY71C
oeL9gLeGXUddTvOF2uFVUnP3tJrg+yX4An1MOKottASrXVm2jXnBw77or+IP5Ll9w5hVitYYJ0w+
Cvz60Sht2tKnbnvg/eY6tr/ncYgsIaEls/Emnfd5WUrIyYTsp8m18JvTRAj5n0J9WeaB9lgxaS+H
rkliuXOr/qkeHpodzFZTZew4eIWwsvicx46zHmMua28uelI2KKTKyQfK2CFy4XGL+ZBZXsi0gui1
Tv/nw+c7z81cg7RFEvjbcknfL69iVrym2HQAR8qdj5I+63LaXgELBgNnLdXuOINsnLOT2KacNUOv
60WNROOluuw7CGL78oqzgz5lXkJ5PGUc+lOI7cYOSe4NIPM8MXJNHBQwDNjF5t1dMnb884OpPgrG
IvhcqxOJvTXc0kWgCzyrDh+yjlYK9R4e3px5tzjXO4fEb08G6THas2qolXOSLx3CmmfglQctS/UZ
A2Z3TQG7kqqvQ5RS9oT2oo/1W3zv1fTmh1kLVsgSEH0o47oXraXz18Wn/bO65PpTvwa1G2EWRQ3J
GvU980qF5WNJXNp3Gi/7CeKy4xHqcJGW8Ki71XUP8Xdun1aUVamN60svV8PvzCm0/Wj+VeG3zsmt
dapB/XW+NVgXFo6E8ytg32/9W+q2GH+Dzf2CHis4U6dSBTTILCN3VXWDEyWsq+uP4oX4OdgNqgdc
Q/UsUIArP+8o3Tny5k7brG0p1+UdLU50gL0LbPUrCajAvwJqZW6BYtuOFIXw0c/1ei+rR8naE1nA
w+bcyz+tgWKuRDAFEQdip93SWEoT/zR33yNBtEColtaTmBVCFFq6ytj+122sS/2n6eL2A78W8wl7
cEOL5cMH8voQSAR0Is4CgrAIHPb3gQJuuF1meJxxze0wziUz034zko+LcRzy5g0iZcw5ibda1gfi
AuSJAV6OP+nI//U6lu83I2BQ+5vdt8M2ZtXhCfK0PUEKmNl91yw74f2WNe4u5kC8xjH614MgvQqY
LWRnkbi7t5FX/1NjOsvo8NZJ2oYtZnPxXizzfBGfO1xNDwSWoLC+oOzMDfHgjbHBsqCU6zaQBmD0
7a85f/ayOyTeqpiv2Edb/LGjjtqEk36yoZhJAiV3VmTrjgZeO3exdNTk/bK0DaZLnyieIqo0AUKk
kWhrf2Pk/KpoQrR5gnFN4h1GqPIisTZS9ywVleqwUPFEDpvOs6YnaUSIw8MSVYnVaSvD6OIccylZ
/8kBzmQJMSoO6Iavb55P4KaWUPrTAJgiBGhtfGfh2pMLAmYTb35fprZHhhi2EIu0TLPPVCMQ+BR+
lbMp+2fCRFRpctUCNJHODfdRJKkG61q4bkWad8BEQ+laBKJQYKqjybnwVZLda3wYXO8Nh1Hm/ABC
HusOCYUp4eEdjgQNt0Q/gszs5pDTzen+5kvn8OtofdqipkB0rrMw5tWWu2Wjtu0BvDBb4oZ4bZgN
hCaoI9tMbiV+Ju3Fw1i+4eklhHmvRXwFrCJMGu625Z0/k98l/N/QoTWeg1Rqcv+UdIsPhLAS4xyO
HswZCWcOHx2a7z/2rGdcSPN2/nLW3U6hE0NNvLq7HdXIkkZAp/5wSfXiopD4uCsDi+b8a5KHa/D7
Eg8WNao0gdn1rzWEp7TCx+NsQ2RwEt9VGwXmVGy8L6Q1lEWVd/xOuC2/8G0udI3UolUuq0uVUZR5
KNKNpOO5evJWfCXkXsznwPWyhKQym2VN7tMLFKpmg4Q6xuEklF6qygQAJ84QaJX0hvA658IrR9lx
7zznc15oR0GX+zYvqOIKNMtXFpTE6zS8MbxYeX/J+13DyivQjhGH5bDquhL/OGbeCCfP13+WJqwC
LPWGzXaKMZqZdc0s/OfiQjQEwQS+720Su1dPHuBSKqyCR2Zy8QA8depCO7nfpUF/w+dN8f3C7O5x
Zo1+Bgz1Sjwdx8K8ST/4UIMeUkJ4HbOesySM2FO34UOJpnzA4rWx5CSg4nk1e5aDboxbG4ZboXto
P+GV33csG6AVA0lOqXQxbOKu6JZO1JgsrD3TiAuHO7HawThCjxxMlUj/jISdFAdJ8/m9jkypxk9t
vRWTN0BHepzI63laV3+KXMUb45YDV5p5IhpEdDNjIKZgGwssXCzRLyfupacc9OD0eJC3huJwDJN1
8+DVOg84qgeSb5Fp9ps6Pz7YwJGx0Ypm5hCmxKjhqJyhNtxmOaezZHJLuJxf6/h89eamX3ACne8Z
WuFZi1sxAJo1yyLr9CXqlBHB6fUXR2fJiaDRdHBRh23ykJSF/xwgdVGJ1w3OH/zf5lf77105h+vm
2n4mJlZz5Thvuf41AO3qICNi8K3/5hpGIZEkAsfTlJJDN1EKYK4Q+JoJerwOy6mRvaGa7Q1ZIpSC
3HiKcBoCQMYxguJ7bqEwYFvfvjVZmq/SBydj43UuwxGuICf3ZRhuSp+G8WAN5ISrVzBKPcGnv55A
qRjrUHFLw36qRzNLpHiGrXrZNmHbrECoo7ghrM1IKSm4zD87JAd19da1W8Bez5al76zN5IyofdV5
2d3fbXCB6vo3IQCXxF+jo039aAlo5ZxuXmCMKYbLUke5607j+o6UxzKHLjGTYeYCZtXCmNq6Sfll
nbH91fbETCyUAVGNkMrQza3X+TVytFyyqdbMXl4QEMNtz8gzrOBD20V9RM1ADZ6pMzZ8E3O0PJeh
LsD6qdXh74tT+i4bi/phzrgIuHGdXMO0A+sBqBW+5sMMcOQTXSm2ahhyxNZzqWX+xzrHEQs3eiOb
ZDML8o7sW8qTsGLNOjZoSSxBWdvoXIPfKiCUOl7MULH/efZJbtAK83BQoVu6gAISDngaVADEubQt
p35PLL417JtsNv0lmazZmc18m8kJpcdtYMHo5ReAtGySbRTDgpbiF9jM//jMxUXBCfxWTfJPQefP
ETVK51FTFnASGRS7OGF+RPS0PkirQE8PtyPzRSLyNsfVIRlnX+MRyJi54K0FZai8tvP5M69uOx6A
0QBt04Hw9zkQkAE9UpjZas/NQpsp6OQ/NEdoHU/8pi55jCLPp3H7gGiYyzj+gASy4dqAvEZyDcqY
4omfpGC7NQCkc2L6fXC0dylVzz8hhfC4bBOF8Sho9wQIDyqHXseZt+vQk09uStO+OVDzYyMUSjvu
hVLxWyfyhxIqyZIXTE64v2zqGHyuW3kk8o1ZGGnlcWrU5XwCqpX5CN9PsF73ofrN+EAPcFirpjux
S7+zDfaurpZieo6IVUCwBKIgyyn9j8xfwgaviMzWkvvk/g4kOJHWs+T1ihuk6Dld1itBNJ/HZTIC
D0Mu91olpEPCCQFu6rvjCMAV+3CaHSNICv+d9FohVjICyS5N5AE2ywav7XZwzDy1CRPMsRw/iik5
IxJxJgQMSA6ioo+Ssgg4jp5Arf4JLHXxVDMKN7X9hivCuegUBeCqd9srcYxb+dKVS58HBmek9XQ+
phHVqJH3SsvhgcVhLdP6WOKTQWlLvng6vH9iouP/RHmQaReofDu0qb/AR/koB1xNeLX4ul4TBAEg
zx1k+JJhn+2WmpimP9kLqxaN6IHs5Rbblv0EXHaCRKjMVakOqToT9usc/toTW1eWcYNrJYCR+2aR
s62wlfTu81UM8pyUTwGvip+t2jJiWmZ8VqxpKoE+FyB7SW9rvMId5dd49DbkkfhCh0DU/nN52UTj
A4vorDd8/6WPAA9p+9RXtH3BoL5QaOzbSquIkK2z6KDQneFJHQcAUEjP4Usb1fxnaxccb5aGZ7Ke
yqEB5FOCwp53lHx4SPvnQC5QF/CUcTYkTgJhj+dQ/zuYicVGoNUkrQ0NwaYeL4lfaSpEe5+K+dKv
qqRt/12mkUw55IIcX4FpRBhrmw3x48K+m4JDONEABOwyYKgSYTlMWHo+PpbI48DRvwIs+oS9UOf0
4IjlAdAvg9ZeVsu1k1NnAgrGxniYTK8vckv4vR4xy+ZL8je2upNOffMPlxkneLldpdUxiN6hOR5h
CHoM4yShIPmMUX+jnanjeDOvMNuNIawTpBQXpzv1LsLATA/M9VkeQMK1wyIsIWcbeMOvrSuQd97f
zLQZpnMyMDiCxLE2r6bqTtu5sZpAujCXd9ImYw4FrcNVmdVKfSMCIaEmv/jGonJk3UIOk4jwkCZO
1hNnzlU/zBxbdlyNoOVk6SuOQdDNq0acH+r9EQr9HGt8rNxih/rl8yySmznvJOe0pA15g1YN9xOg
0AevanXuJYeSFpGVJBRQYVUG7vaC7oDk+dFkYgHYCKEHom1i2VcUE/ukrnYQ+YpQrkNzbhXKi7mJ
IfFXErpqLvjutxH2Ab2CHl9EIvZ7U7RAUI0k3GBVJWi7T7UgJgQtoJPBg//+BmUW2XXS4XlKzgJB
jYW+saiwPoyg6x6Qo5rq8h3D6l6Mqn9e/c3pEKTpjDv1yvDbcYzyd6YRjmsQNaZr6RyHZ6EClW3O
pJrwVAfslBY6Px15JMlg9O7dR0qB9B/B2PoUXM8HC3N2PiTjoZAIaPSkj7Y32VFa+Nys7zKkSk82
ohhU5iJIycQDJ4kMj+Z0cxpy9zBjpc0JZjZOU0+ECfItnU53sfeOuQTTjesCb11tTfCFrO1p8k8U
RfiKoljYBGsnEZGo8U42luC3+1RpYQj9rMV+re6Yu5oKNj8bCP1zqqYgjJfapW/9N+/6q2q7kKyz
hmo+kSIplMjkXCimIGBIdnrdhzYExIphUE5dkmqElXI9MzHcWDNKLkuP38UE+/exKnk4a3IBF+Fb
m08nzQbVZxjA0riY06R9in/mch5G/JTwboonQ3TleZFDKXNmq21eUSG4Ou9ySb+o4GjIfxX5gnkh
uupKr+v1arG/6cbhwtoXWa7MqigkXeso6mGcHF1vfm7KpBdIxjJxrzo+onyZqdpC7rtaRJVFXNkJ
F5a1BDLp3vRqTp0rQ+ydZuMmGHfZlPiQzXz39hkWjsFIPmL31jovUCPbNmt1WFSa7DPwW+zj4/FP
ft4cTgU+HgLxzCS9EpU1t9Qo+ABwQ5HHo2YE+peCSCvXbUB4JtRaBk35myts2MIMqyQudkySri0A
XQb6pvU4I04N4xTngmZEZC9TzvnEq+bO3pVS58rmTV637X/aPlajOymTEEVn+bfxvT1zHVCPNrFE
OZf0kGEVUShlZGDoQ0JjPwymThlHo7YPtjX8c2AaEhxgdzuH1SO/TysHYfid84dk4+aKn5Oo6c9c
7Wiuj9Ug+V6kYBls60uwIW/NZXU6VA8DL/jQftAYG1lhIRs87/cs89bocbJsm+nHQLLxEr6KdNUu
b3icbn41xxR1gPJ93yiMizuMs/mYCyJOZOqcdTKU3n9sAU0SAtb4G7XiNxnDmbCv5OeTsryexkVc
Ezpkx9PsbNU61m2E1qmhPI607wvjtpblDzij0K3Zll6nWE97ilf9aJrabjYdVyT7osjPfH9V/bfA
BM0EOV5Dp2Xqs/a8WSyhk3nfTJSzhH5ILrUmjS/0jFhup6NWMlStjJfVxsLpPt5xTURqr1VNzE2G
2eImh8bTasfcB7t1GCdxlvi7x5zbj3vVVVf1TeUDLfD0JoAtrWuGH0adE0C+nWWOcYIqI+E9asDl
BXafg8XFPk7y8SjTRt3fLQ4w5ly22eZy8gK3PNDBW0iJEO8arO0OFh46rC5+1QwpKJIngOJsuqGp
pcj0Wr8oVyRrEFyhWvuWl5NijMXnLbDBcWTw7EwsDVK4eoGhHd2b11Pn+OH01msdLFeiSA8SBlbU
nmOdqet3FRkYXRoDTp9oSDBdgaoDRT5SuN+pJwaHSIkylqTkJgapAvuKqczm+uW0jt4TFeKAq1KA
bUtHcwdhcaQXJbVEfkCx5fYz/Aq4xxUzEPTbAPJ1lZWYDEAvscy0uLwH4jxFgiY2cAR/GT12Yv++
rGHWKGJmDlLyieuzYqrTwgCctbGLqtS7Kcxjzm4UhPLcT14I8hedUl/W0iv0BACxMpBVBeOjul/u
rkFX1I2/LH6eBYNsAGDsO/wyJeXWXcE5eUHWm8iu6dmwDlMlcQxWD07AnFeKAAJbVZTNs8OWFX/6
ZHMTN0dhRD6DZDN9aXZNAdZ0OwEpOUDjaYn1g/j3u1eIiGnEOqHit7BKtf2zTFkiQ7/W3jKM8DNL
VoGH+uSJcSnRfzc9AW1jSt6gLYogXUcx6UWekQwDao8/Y/7OjBSWl+HZ7DAFqmwaF4sLt0OaZCyw
1gu+TqqO2bGdVhK/Sw109e/AMMZlWUHszyRFJbg+Lf7nVd5Nvi69town8XEEjreu0zcKa9S03u8V
6jtZiM0mU9TOWtpu/cTtaxKAuQJMKQHim4pB5PR5Q24mBRwrpYGl5Mup5mwJPrItFXC8Ai/LKW6+
5g4eGweewmY+1FxX6gxIG6hHLzx9y7/HoORk0NqI2c/WF7mKR22bBmVNcEXMTRz5MeJMHdpVkV7y
9si7R6QQIf5VbMlhc85MgVRXluHrwvUeIgqlUXSxeA8i069F7d75z5PqK7ME47dwgl7ngZEWcjcQ
bJgKZlTMY8QeqCCa9SN3EUVocECX0x0zfdIjXNzRRYZkEYaUKNpAUcpCb0t4qg2lNay+d0be58nD
aol56Fw85Q321Gk6WwI0qaFF8SVaUrweZ6VMdfcJvfL5VSisAOnaLHRLAPdgNjtV1WXQuGptfZxo
oL9hXoDhOZZ7L3Df9EfNK16vWtJvTQdFql7AGQedXtuZajqWiHRJHKuMqYeFdOCNVJbDKvsbUw2W
AbtvIY4tUd+zR2a+yupeP0q9ZXUDtie4Um3ZeJf44yijXtr2dAqdtUdpNejBw9VbDMqoZ5Rv+wyE
b5E5eapoBZzUTk0VYYKQ+h4byhV4aI07mjbPiDAQD/BB4ssEpNmN33vQgcVKzGbh/8JqMA6xfUav
unBJdCw7iHhh3fUhcQEt5Ut5qFnkgHo8+qJMdu/eRi3R5rFE8e47GHgy3e+bi5rVWP68q/x33R+d
TRB2BV1koeLefsr8gd85YXq+HD9/b5IiLIETiMeUy3jymkrBEiHkp1+F5XvWcDcfDjXMUB1mkJnu
Zljl0DJnCNEg6WDTquBvXcdg+xVlt5fnsNqaz0+FuLveana/mWDtUKoah2nUIgLJgZSCdhFb+Kbt
uCG/gFUA1a0RJHG+s5jPfZIXYKMf1L9HsxR1y/CLRkfriJ5ModY2zmuWjR3aSKxcbTjf6PqoEiDb
aReIa+wnWyUSSOuwDxBICQu6UcFdrp3GTqk9qIpbhkN0SO2llCb+FgTpS83zwMI0cg3u/9ZZXTyA
2WoLBN+mDDdDrHWG5HH9/td4JI9PQ95Du4MiDc1Q76oo6Wyd18vQN1FwJP7E0OHP1WwTXC3miARw
TH0MTtcIQl22lGvzrHLnMXqy63A17iCWrlLIXxlGgnuTu4qwlwkaQhSXh7QjYAq1jG8X0nNI+LcN
m5x72ERlT1pGfQfMQ5NKhZycm84ZVQ2e1HVwK1GAK4DdiKGXHuHg0dlmGGROpaKfzKsKslk6ypE2
0weEKpxj9UnEQq43Dkd4cvHzpV0Q8WFyU43JW8ynSxVZokl6I9JDSeJ5Og71Y12lc5HbAZ3v1+Qs
QThE5WLvfjHplsSXehkYJLvo8NrmiixAP3l2ZQL5SZwCj1j99bx8IqM+Zshn6JbejE6s5Pmh22mD
VvUu3qpjQerNNQn0U9Lm6qx+cjp+yEYpj+GYvQSFEfXUL5Gqb29gYyWq2y/ksrfC+ZUU4DxESH+3
uvMHDlHeSqsuYOfUp3ijqsRSoCOv2RVRORPpsOcCKIw5IMoL2dgPGJfv+nHbAKKkqHJyVmyr6J4v
xkmGlZhk6YHarSAVqgpHQLDewvfFtEk6vb71+MEFi5xPwj1QHi5t8BsKdWXmrrPaAMxB6oTywT2q
dSemKbUO4IHythw5mPh7mKM8liX6yqGyPtCV+ep5NP6Jb3FvGN2jMmlYZ3h4M/tsK7tyNntiLXWO
IhQzMO7eEf7htcGPkvgpI0M5uTYGMaGZB5Mm23x8XN7hBx2aVZr4+przazl4UoBcHxG6be+GT0bv
dw8WBNmNs+0bnUsSm6WWl/nBJDzGQdUaDh6prNQBABEyMqPiHceVnCEBuqscIbGHF52whOFf1UNS
Nkqss+ZGkQppqmNMTBjajqvP6YRbtrbmPArammiv1USjejHdX6XeKX3w/3QPD3v//tNwX3aW818p
nC4uIRJhKsMpoiTTqX04iaH+lPAjXAx6q00pbp2tZiaoTQ+kIwwcKi0L+mT5O0k8/4ufsbkTi1iZ
L174P6tSjvvc9+ezqvcHhgGVSDdtzQd6BB7pva63bbPvPeHStWh53MAdQYBhOJdNKcXyn413nzmm
3D4JbAd1LIVPFRQod2JgCvfDCfumbKdkdPuV5RyuH6kkyYi76HAwauyzp+YMkXT3SJrlMWVNTKqn
4rd4lAbDmM8+rH/EahtufF0RKr4Q6ufJ1LRV+Id3awcQy0DReG193ECY8PKnWIr8lWtF+jfvZZZC
jwTKh6iSdNaRHKU1HmMj8Cjg2Vy0yMsXqBaWqGsPhLQZzaIU9rbcNbXPINAZKk1m71UQNM0RP/M1
qvDC9bF20OXkibrsKdr6dYHmmWRx4X62fEV4bv/cU3sRZJXKwXUtJTmFnZTzuTWomWMQPkGIfios
KbVEMLsGkA8M5mcsILZwrg4a850H8z3K4IOSRAcKAs92jAdhyqIVglSfBN1kznt2JcWp0XfVLEu8
DqdUF7vjy2glgctKaVXK2HSlGc75ktF4clTU2aYVPL0V6Ui4/vHxmqyHLIpBJWzfwhm0arvMbH2I
Ncwy4ZTCta1hqAmj1KcF5didD55HLQ6hgcwEkOKl7Mf0EXXLOcrOmmVFxbkkJI1yCr0BiT6zgpie
Aft2z+nNNGQcnPlTBZ8vunReaOTABY1U682tUVD28GYSZkFJ9Zh+hJ4pgrs5bB72kqwV5adlvH3s
9l28xLU8GY3xVIYFnN7Sql7VfdC3fM//k+2GiI+Wk7eRNh2zMEAKJ5wKlEbXdoFr0A4D8s15r7CN
qdkNS7Ynam8G9MZo4Lwq9qvUyw0pns5Ji6+uKJHGGEThuy9MQ/ztXwYVu6m3rCGpU+VynvpHI1WY
lG76WtjX86tSiAxxbIHAEhMpPmMMqXcnhJXcN4oVUSf3BaqS0xfkyN0f80Sve4a05qTJAgictW1x
826mZe96qNHMRNKH2vxPynXj9suTguYfOzuFCK+aQNPa79cNDuK+54cq9N0fNpfkl5y2pvcAe11I
RUj6wsZhNcy94SekGqoWJYIXjVy8yldO7cHZxV8hOxDxei+ZnLOFYh+tuKM0fwieAFsxEsBN9IaD
98Sz9do5vnbWTL5v4+4dvx8b7ZgjJ/EwziSEczpgZTTph69k+KunHbW7nuuDmWhcKZoW0VXLUZb+
7c9LmRuNnyzJF2AQe0uuSFIQtOTC+9yf5/KOHlqh4KL5vUvbEv05GHTDUD17IY+P15wTvwq5JxEj
WUpW5NCT18H7VQAloI1V0+FXa3EYzI6BlLMJ/wvS271913EkBsAqADoFsutssvXPYGlxDJpQBJhp
NxWrdv+lVHbtmslo6X8Skr9Ns2lN8xFb4u0k0SKf/6GAOrIKXoAoOlNrjbX97HFzEz1+hn2vssLz
miAtZwB4+xvnaEQFDpbc2jpsalV/uydjwWejaIviEP82BVcKo8lehRNQO9XwIG/peJyitoqK5AGs
9gqnguGbX3r6g5JNk8uaIBZa74bQ6ZGIOXB/B7PqIiP4Y8f4PbrLvccO1RHTHpybgCekWKffqIXM
oiR4gk8hnLXbGt5IDSTOi0l1X2g+Np7Xf288zTa2ilUOPltiTWMzzj03yeyRMiwtbs2A3CvUKm0Q
V8ndfQ+O/DJrMK2mokgFuqEHutfAZJtAAVgDDUgKWvHV5w9iEa44a1nzSem1Vw/6cXvJiFSwvZ5K
TMMUNUzk30OgjVaf6gKvRWQQuqhtA7jCvgEO7tFlkfWrbLDTYze4zVZwnGVnXAAfVfEKlZSbgiST
csrUhlyAL9+arXWAq5JYCQKeMBK+DU4dLo1s1R2siKx1TQkvcRsFGZ+AMvI213k3Oywo2kUZYR/D
t7B7I6I4dWFRspmZr7prtge2Y6uu8+b238FXJ5duDS1b32FTFWK6iqLpaBwPbymwHg1RjdUJrHqK
XtaswUO84iWSgFXvhYnYOHyasgcICWfBBXk0KuJNhWr5KfiDxNlZzLkrg7PqTl7f5ltko8+DDCae
jNK/did52pxI8qbetb9zAO6wEsE6o+lrQT1xkdNqxxYY7w8152LXA9T+5q9fMx0uQQazUXQ58Mjb
xPZ+VXuaX6eCHU5BPMZ0ddVv1OVBRCtyoXFEPOZGYU3E6C2JPLWnwqZy9tUpQsbuD7v2LTkOXWZb
SFHoPOiyzS6nXSH+nMK4jbdj905TEDXD7wuhVc8rzXGiHETtJy/l3CE2twUNeURbyGC3PzymZko/
uyvBhLFETRfk3LVXSX2jwYuyXGwMrz5NdL1/dln5EuzdgU1AxJGEVjt18hP/Qq1SXSxsjoWzRAka
lEFLljtx84FF6WPVVETmiWASNgq20HKsFPFjAUIJzEjghxhW/O0d5T5cCRtSba9Xda+txviF2VNB
BAf6cBqMGaLkJAU0Os61RnFDC2UvCdycDSyYq/HcJK1CRLx/ogzGuuYpExZ9I/70+qO9PXS8OzM5
ufOfmBTTKH/euL1ElbisSIOsKuQblK7fqlIpbRW5Di8Zpbe2XVjsrOl9Kgkrr7CeDK64caU+TGLC
7KRXUWdwS+cN+eyUcY2DJZtUtQaWNxAQEmZ3ZiJ4yHNj51a5s0gtlrUAdaO0bQ89BUvwvuUwsFCE
80CNhnI0TogvZS01FkAfa2BIpvpvw7wt1PYj7dCVYEOYfZRmfm+OCuWbq3uhKTi0HFB1eTEya3Lh
qXUZMZncCNNHRyCAglpPSJqsF8yn8heY/A/UoBrtd9cQ1u5X9ocviR5obEKo+6nw9H5NpGX2xY8Q
7WefK1OhxBL9/3hrzlgEiKxs2bbnSSX6gZWgh0zK6vCLmYEfGzXdGAlNGv/Ood1RWB+oKsW3ab10
7MrKy7pzNqXQDlv0tbVDsPy42FdqYjabj5MEAg1YCAcrYC2lZivcfY1K4BVSoLOVWkG+qm5Yr6b5
5beKmbUlfY9acNNYShR2fnvJqpkfOaR2/ks0FesIdh03/b03N3Q+WtTaut7G3p1hySlhLAiE0B/E
/t4zrlg98rPweEBfDExRUP72+vGkFryASIHH4iHUhmtaLulxuA3b6KF9tdkTRiyKLJ7woI+xGEWk
gKkj1qKwUk2zlHxZKcsLq4iTqlDBkQs11FZ5GprZYf3cSeyY1GIZphEpyVgDaBJ1dMCcLzHwTAgF
10F5wH4fvhQt05bIt2dnH4rtbs3zPreg3OBF9KwTNZDCYg+9d33f+d63EDh+iofYI2j0FcXhnRTc
VwuiQzwpjdS35quuK1/XJ5+i2UbMA8e88GWs1p7cFqiIhvISCzHPsTHyeSWFSTzIX33Avz1BllNG
BmII8IKaM6bYTCYeHVKdvGPiq2uMpIfBOp1vqPKynXOdzlogpuLPtcfZkyoSw80lzEC+jJ8+ClZb
X4iFwK1d6bvCeHZLyihiL0wwIexMy9XJp8gI69a7i4/J10+sHTNZE+HSaah7ZF8zBdcN6xJHxoN/
0bc5eTi0pjBETC6lVNzf6fEVnLKlPUNQpo07G4WgfkJK6OEAvimGu2h96Wc0Qu/9DmvDMTRwacKP
pClIPvj7JeQeixVaJKJRiDfdEk55MGLgT8B09IGbpwMNiXALv1tba2SHccJ3nn13+LIbIs4SOCHP
VwlTghaFd4fiK2mC77Guj8CKyij1Yb9gqCAVYWGea3XAKgzzjmCPY2JpRONtxowQfngUFeowRGpI
abLqWzh9vJXJEQhsCxMuSQpXQTL7QzJImcdoIWu8bLdD+z4jv+Yid8BhP0WQHtW4Di4YMcLq4feF
i2wEfZ1RkPXRYSxPIjxcxtT0v6BgrvTDtyEIOU+AAIG3G80ZUHD2JaIB1sn68Z6Tluf3GFLJf0c5
yuWeD/4KgcbXonwxS0XQWlmURF+0t3BSm6qq7XM8bPPidnm2XGyy4j0rNPGBU+19ctSN+x6eDCeh
8lOQsOt+L6tPv3ubCdaQpq/i8sMWrjaDzlvUL6zlr4wS6UsGa3QcBl1u+TMHMm0CJouKbzd0AMqk
R7BymD35q8kYVA2wKyugsHXdqR0sS9gAobxuJkk1T4hkHychKU2mnO513q3BGcsLWpp8CP3LdqP8
VVm/wADiO7b0jxV8JNnM2OAtB2w/HgQyfngOR/vznETFuXaWMQjGVK91bC5aSLGMvzI55OUz4lAr
kCxM/Bn2aNfrOBYi+5CUriuqlZEwfQQkAQ7fYYLy3R7ybZ826MNXnEGFo47v3mVMOU6U4FwYXrHU
Q1trSQVk/eTq93uelSiGGAZfgPRR1HKtauBYRK1JUnBUgDONWQwuNaRR18ZtR/035SRQOxCQgqcI
Cg9/SjsGQlvzOFKwCK83EFRUaWgkxzjtMBfKLrXGNSQOa2pTCl2EwG3MmYAcXFfUK+ANXXN3/G7Q
+jfM9Z+3WkUe+I7H8CUmjfGqppRjH4R/8D5tM7NFmYQlC2NTnPXP/y146nskPwnbcPjXVOyVadA1
j6zLLJ1v0GH5DJogA1oj1uXd7Nn0z0Tn3IwTp2C+6NgkmKt+y+Iz1ds6NM6mMLFRwgTdB4OZTf9n
OsJu73RqS5WQWII597EEaMFjdn4sNTx00W9lbUmRN3vnusS9OSRx/i9k3Xjmui5PtQ1uk0j/8Yzi
b3SjZfzzuvjPKlXtXFmn5PTf+lg3HUXFTN3qS12Pj4UcCSkMSd3yhFn0qK568FHKXTS+s95S5hkK
0tCNWjAJq+ZWBSf5VSkmGnl1uOvODclOHebdaawjXWvUnu1R0r1ZxRM4hZUtiKDTDRkV9swFXB7y
Pt8G2RMy3I0lIoWgsqPDp5mWDdDfR6QKWm9J+lzDDEMDwvq8TUD//mORSpmE9uaUhA8FvCOQzw5L
95gIvvnv+2N9RCH3FKvzT503nPpX8o6HzlJwc73/VCUUifnjVudvxR6+Ojon1vLLEZ8Hb1lTd59F
N1Hk2byOiWn/5bEkjJg1BTiOKk/5AwE520juLl5so7IlTw2/rL7xwvZtHNsn4+IbUZ+0E+yQ/WGi
YiL967aBYFDfU8tyzDYTc3U5zicYKwYzXddFTdP1iPer3kDpjsC/9aGAspjW9+TZzoQyPi7txsjy
RxUmYTlCKwFc+Sh83O6QxYbiV4kfrq6tqLL1ADo3YkkZCmZLkGyf3gnezkdptNlWFvxR7dfRMpM+
vCo/OG7gqnAxzswEu6U5HEzpqmd6TESy8+IYEr+eMC/23NHXcCo2oYYRt4jKS7PYOvK7l+gWkYe8
Mqoe2QUlBFd5KrViD0NmV6DKGpOp96unISjRMQj+XhDIajSXXjXtrglKq2JWCz4hcBJ5LNuPzpaE
dM/8dDQyv/5c5VJDWPabGhYkeC3gr+P1qOvP0UR/FaJiQzCp/R4DUe5TlCGrJfnK+dZfpjBo37tn
4fTVU30Jt0zFk5vOCguLUSrodPAMz1Z5dFBPGIWB8cp2vmxF8X2oFbn66a9bPGUcTRu4yLkz4TIT
1MMJkTwQc+qUjaZ1nyaGKBh7DaV5oP2OlMgi8GH6AO8CvRvxf9a9/mcGaUFtkE1Iavk0+PoYMWOD
C7zCynlv3WMLqGy8YKAO0UCTV34vkoLRf6jNs/F5cWhCSg+t5LyP21qnBmoIRG+z9QuoMEjDBmHV
LyBAicCWoDKGuEqo1nkbJoK98ztcirHBZX4Dl2C7B3jrQl6J3KLVdcekdWOPhI4xICFBOiAa+dcX
Mqpvx4T11kkHRF5y83dj/5lB0y1TSKGtkiWYqIPzgXTjLfb0mWYzAS4cHHpKDFqhEcZDxe4p7QpU
S6LO0g+raK+RVRnbvDMpgaGJIGYPaGa3rWSz8sro1QPYytvsRGPtMCF4BuHZlO4bqgCDS0jt6Yho
VU7eXxwO2NhlCdi+Kz9e4+kSut/p57EmayvIadT0+ZIq0kx4paOh+mnkoS6VSnhzk/JevyIbXcQc
e6yvulviMA5kQ/yoc7gZSNOteskduGuEDXNgrwn2m4GjdaJiolGxITWNoq0W4PMz71060OwsJCyr
d4uLP9O5+pI5CBGZgsS+MH7MtAo+LyvECWhT/V+Iy+v1mf+xyixHKFHJ9q0z0yM3R0pzmbNBOcY/
0CNkqoW2PZJGBzYScK/hzwOAeg2UXqbO3eydfO6u2L5+/O3lxj0vMBrljp8LPsiqj401NShy5wJR
V9KQLMf7EqMr41uqibat1YdF9duik78aP1ZftLsvoTMDmNwMgDL6x4CHj39Iu+n/yPkCEmRZb2M2
gaj+T5m3QvXP9b2msSGz+oOG/EA/j5XVDNMXB0xHlmvwO3GQKuDrEcgOPF6KLnnoquAT+MJaAAnZ
eClkelzDSLlZr2DaOnuhMW0DGuUag3g68uLmBPrKgwPljPVjYFKhYhalGj0L66bXzoLRFiwarHgp
iDI1B7/9Xum4cEAPgsk2uuOh10CPqPpYsaIcZSiULIJdUhg/E3XmI3suxjlQNGj673QUHC7zYsqz
8ZrN2pkAWudW9AnH2pJcghXEbltGhkDj75ofDVIIzKpv01IZxDkIwahLIvfbHuWe9+kf4TBILB0E
jLvOHzDM0JBj1s1T+9+u6og//aLotnPb3zAS0mdK2pl+PyX/VPfjT4wJgJ0GcswJ0bzieuMuuluC
AYhc/Y7jyjge6HjdeJGSQ8oYIlR1oJ7ru1/8tnu+AJCY5MlnxQvLig83913oZbqrieUZWqtY7R4g
lucX/Bq+ukKg+FHwWtRxUwr6NGsAWKlsJxrnm70Ow6TqTDBi6Yn8RSq4jxM2peoZzQ7ILCMc3KN1
2bJADMLuZuMqZOwLoISCdMdpLvsnzL6YXB4kszo4GbdwvP/qjqe25RHlWBfv4L2Z3Ji0EiHw1Qku
TJe1yXhZ8DL3BuBQhl+mbU0C9Ho05Gbp+9p51tGZGNjfs+hJYOIEmZrRziErUHeRcrPoKLYzccdE
MaAT6M/57uke3p5IRVZyin2q411jd2m3S3R/99fjpKYZRiu/bqvhyNfKNc1STrdIGfGTxX2B97QK
4lVRCtEjV9tG+/o1lsXjTFhpQjS/RcyIYh5LQfDU7+7UQEJWfjLOwWIr9MQc5efT3XuIkXBQhTUn
jYPSlRiWTNGuOGaKRuD2WTZGmJMey9MMX9ak5Ogja7BKs/DztC7scGZiHG829KNkgZ+9aFftQUg9
sQ4pL2WrSaG2e+RWAwb5RjfBNOejpiGj4m/5u7+2OSTjQFsxiNibAEE7HAGTLRGkYUl0Au5pEjMD
dWEH56vCt1/FYDQ2JVOl1czp9B+6w1Lx7wx9rLTaoNxJzLMBFMR07ofoBcrvtN8u82PYxouDM1LX
CIbp35mI5h+laul7F3y0GA4rwC6Kigi0rHrvjIT/UzFX7XPMSRvwtkLIyd/4PJhF1pfsy3BaLMyE
lryUsTawEbKbokpM/ZTAZ9zia1Wzdjnjxa1MnlTuqzaNRJ6zcJxMBIFQPEpJPewpnKqW3p9sKz6B
t+goQI3UwANej8e6S6ORsaFaYiY3XyM6EiXw98zo4Axz/iJKu+TNowHx5sBx33d7nr3XssvuOw5Q
uoOsCVtMKljH6EmOVc3UHxApWKuaC2t1jIfAPRZvCR65GSFPY/gMWw+Py7Qb8SN+lI5bUFRwZTjP
hpi1hkeRRqyo+IVkYm26NkOGctlI3AWIN2sgXDTOxJoo6nXTJUVgXPqxY1ArFrzhdJn3Gz7LnRbN
C6lTiWXOrxBdP52SsBrOnbiRgY7rLo5hXIt+htAejreeuXaLlozx6mJl3TSkLL22EvO42Iw1lwGD
9JH6q88ToKoEqwoSMCDrxwxcrwo3BE4046esp4HpSLLvPkyYlJDZu42P0TYOUUSW2a+yNbpsR3yh
Xv3OIwGI7WKz17yJ/RKNn2L6lcIiICu5KjjCOXmRNPS33uwbRhEcrSA/WvTVoFHOp+lLap3g8bae
NKKdssJOQpXTqE3mwNsnUX6UnzcY6FQ8MB2cccr5fqwEs0lF4hooLCjNVvT/bVuUs8Bh4IiAEzSb
o4oYJ4KaeFH8FxljoAU7FwrOXq9B/OlDOjWkLavSij8t13/UheDZN9XEQqchILHJ8F2f8lfTCJYi
Vc+j+Fhdk8nV1mQSin3oi2e76l4hgQ/iqh6XBiYoeGEvjZhOcvJqwR8FaQAruH4/FS5H4qHyHcAb
PfbC2EgLMc78b53LXOFT5uDbvrCT7Y3RCbTw8rxQXhwE10ab7x8sMl7UCsFoMSOwRxtlfLvLvpyS
6bBd1eaNE5K+7Mx6mpKkTcSqLCcuxrONXrmXE6Gq1RZLSHjwRS0Gbbvfu4NMMgFCzOfFRgxf1ghf
F5DxoYJw/qtyM7eAxWAIn4aWm2Pyt+EnfLQNbGnwg4h7UIQnaZhcsh+CcuqdO9ED8hlevY/A+9ml
JuR6s7tjZojyPEx6Wkd3qN/SsIIyMvqlQ5xT1uoJeel4wUhEtp8UhoQqSpS+eT9dKXoBhwugwis2
SmAgWlCoxhCRWmE3sEWaVW3WSJzeDdXV7kZRXv5k9bt6ASLLo4P5Ruepd6+rXr6TRVSxWRqJRUq0
ym5lw8yCBkgLxlhfQhhTSMFxZRzyyeC77zRb9kyNY3fmXwEzyOtZXujLSZDTvEsa0VKHuc9eSgeq
mhMIa8FKOAq8QKoIcrxazyr+qTAwFETsRgysmBlZOlBQNVZR+NQNk5Z5bY9/Ad8v0c/urzr1c/KV
3OIjBJgzdLbML9DEVJvAzMYd3UZkip5ebHIxLoytiSHqJX6vqjPc+A81RHjQwLoIX0A19a1/A+Bt
8a1lJW1+wBFZKAQSS7ovF5QtKnGFKeZH/AAgq4CSABUPzkIla2FRtdzNUeHwNOyjoMvMOZ8dmHLW
ZWEQw15GGR/q/wSD/Enw9l2uktTd17Fr/eKbjAKYKmoxr876+zBmL/VjwPVyfcgSnaDsWsIiL6RB
aWKOs5lMdC5JE1lWKQqwe8XrKPgCEdBXoaeLvyM/mUJhGKH/kzx0buEj/t2EHlenw302jc7nWh/N
R8rka9v8PnicR97DQjLec8LHwyG+c9aXzOyYp10Yofs4M3S2nZKgECJON9R1aaKPe4RcuCzBwJH8
6Uuz7QMdETbcH/S+EzUQRS9yK/vfrNpDqtGuaxTobnkeUeoWsIivZnXq04xqWGH1FgTYL3Vu4FNf
A5Z713Q3fpllXUIB32vpeBrI+gV26W7Y2tdfOESPhAhMK5AUYJjJ+MRo1gfrAb8ZkFaqMmXxeiy7
0ag6/fpW2jqiP6jOJ1DPbQAHkjh1SeaL3BmRrFPg405EqollfvbgxxrMmr69ZGxYAfUYmo54kr42
aH3eyDcEa5uT2UQ3MiMeC/jixlI07sgm8bNcLw2hi1ZzsThE5uEP20hzOOKVdQ+VhUDZNy2hc6JM
VzHfuJje2swwewTZIlbnK6P0OSTyrLeu+oneqOw6izF2n2bCmDnZhrKwOiTKa99amkrodqKTGYRx
gQ0Wiy92pU9EbeH4sckmPbdwjNNGf7PSxzwAcmYGdadinLwNez3oea+P925mfy8eFFlHYpRln1jA
53YL7Vt92XLX4TCcTiSOheR9O3afSpsRUdScsMTyA/DGsMODJ6L1FeT9dY1cnpXQDgz9Fa6/AfpS
BBy3UG9JW94X1c2XgTrbqA4bz+7xyNxtm6a/VaXhVkwyBvnrH0fVVJMC/57RN5rWyxwcK3jPr4Pe
hb28YZEjJe5sKkYDy0LovDv8lnWgCxUELB9LIuoEX7/fKrhuZpq/kDXR87VmxmuVMfIJY4nM6db8
sVOmD4+qubHL11Dpsj/DiZJe56eSd1dvYKjVw2FmgCKAulFpV17RhDELQ27c5AuD7i2RMtZqpatU
BewzWm6htSbskV0W9U+QJsa0PzIHwKPMLlWCSXSerIUUqmbhV/R1PcfedvnEnYf/8SBwxWnWb9Hf
9dda0qQyWtsPaPBxiGiEj0qAXdr5PuTtskSX/XBVvqzcvSh+Yl9tpBuBUq+UsPLA0z9sQIIdeeCM
cRCx04SftYWTS6RojKSNiUOeEnUy5FxbHyklTZn9nTg4X8AOkw8EMWCsDnqUYq7r58u9ccRRqFCS
g57AeIBNvKoKswCn7ZnXclhnllWr9VtM/b4gNeEmhClcEuf10m0RLzxya5+ZsjRz5K65rbdxKP6i
7T0GBKp/YV+qBIoXpd3U2F06cgvOjglf9Kaju0dgg4lvJotZrUPhvU/Yfr6ZhAPkD8Tdwbz7tt9E
Lgc6XOxm2lJxAJq1LRDRPv/wOhfdnEGDOUeWbC5K8XORFzZYEVLHrjrJ5AbxNLyn3VAwl3goZam6
/XwuaZY0zJANR2Cl3H9arOPzOHTefGH8mrwsL+hvXSwhW17CRfYr5phi07jP0meRVeDH0RXQFJ2v
IY7ulXG6GMJQq2ojQr+KlpehcryjhxTsVktRDWQ9Xe98L7TunxZkOfwXUfVvGm13fokY8U5RPhAn
e+8HxVm7bXXQDMlN2YFhIfOZvHpsIh9jJKuQW3YvW6QrSKvKbPkV2CTGIk3i41K/uDE70LAKJiyB
rMD6ZKlCDBRKLnld0MDS1MmyGwuzlOvRV/wj1AhfFBp5LivGgymYKMfdRB3avl/135EuH0GHNJJb
pyLkkwP82Gbauo8q0Wp1m+9AB0Kyix7HPxSkliDj9WX0NDI2yXq6qzsZGqiDYmzMAB/sOu7EWFzG
6oLB6NyvMdDet2pCbonCY7A9mmD6lqVD+dnbMEQG2MvHavieDBFKt6MsBOF+4iYJOU7+8jBRdAiL
XRu+f70pShZYIM8+eQnDaIGP2oB+ZCerLTDSG1a0713kO2rOKh0VE6oMAO3iTizOPMF6QYOACHQd
7G8R3QsdW2rnJuKuw5ZGXYaHl66EeQfkHYTB2K5TQSU4ygGslPIrdt55nU1j/r7V+eEg7DjnvSB2
+tVZGy6gkJMOhYzAxB1OLOvwHmWYBCoyxX4HYSvPil9yLJqlJw2rnmcleVyhIDhC0BYXyqo744vu
iKpIdVB92k1+7Ni18GClUtrYkoAEeaFeMt8+UxgFIiom17+bxvLjn48eOmQINh2Xy9L5Vsni9Lju
2I5qN25HHfpw27GUMen7lb+tptjPPbrT3ZglQlztbjt/aqMcaUn+2m1bGhABedAJqRjU0mltn4ah
/XWfnj77eMD6SzaYouARAHD47g7TDb+rgFyzBCwpNcEDJ5cCDp/InMIupqwdlIkS2f2bg2W3GlOm
CpQgAx5a4E3m+f55YNFmkp5b2WHXLg5Gp1O2TkGwFMD9yRRf8PqTPUpcddJ5PxUTuM2WK7uTr83U
bZ4pNo6ks9a+8F8u+VzaEZBYo8orr82L44AJUR4O2MtDVX23tpaokh3vJ8Cgc+u7X5vKmUc6AAl4
GjgjgNctu4MubJOD53vDh5XRd0l+NdCBvzxuhDVlPDepS2A85zVyrGUfYg8SKP609D0xewornCHy
KZ6TOx2w2iHrO7bfSVQI7JwkQrl9OjyrAaoFNYeK/2qiQp812a3to/GBwWTCpj6S8TN1iD4eZEn4
lBs+ixefaHra/nPchv71SkkXoyl5L52eyo583nu32vb8KaItcmpB/YI8Li5jBPfpxa2oJWC0PvMk
eDcRr8a7j0vzGIBGfY1Q60Rb+OfqorAvvzrYi7HG1UnswtNEG8qu5cNNECXoSHhfnLVRyFfu/lqF
PR//0i3J2kISfdgQ+F2PAAdzPRg0bRLiz+ojdHAtDLTiFNrCFUWGCxhd0fWjL+aXHDyB+HScWSwG
45LXgnKJnx5TioeVZfewVD24dmSj9JcxEaLctU6ttK4CXGYGrHbm2+og0dgzBfNpycUNQxGmwOuS
YEBlSlIOpp+fZQVxAOIDSnx7/XG+Y/3848tGUV4Z3K/hB+En92yW26bkYwOqYx5U2cFLwXciG9IU
YaDrzubXUxQ8uTGd10tDOkBiJ0hLRe5s5L6GpbsjdLzUbhqUJ9DDQ6WqjDEUdl22AG4a+F0WeQ7R
RKU1iwWtoAAxfWxqy7DWJsp2+wujqneTM2gDkjooFHFOTJ38JDOlgUWTvR0dJKI4DtnYBHz/KbEK
IjyaprdNy6YNaXgW7LVl5zia+PFpowD/RXziWPJXYQUPxyJ7ZJG9q5fHACRaZno0zMCW1IYiFVeY
W/AmNhVsuMs53CSy6PjcucF7W3/P/IkKXJTpQZiMWys6nGqCzcIs/XRrEVKDjsQN31U8w1+eEMdt
yGiPM8JA9GGbj4OEx1gVCUT3hDbXTeuND5uEpso+YwienmQI6Nrn5IgnpWxjcm3GwsFBb+KhYITI
8vU37AWNgwiOSxQciyj202RgAfKAsZ/tdsuh7SG1CS/5giiibDtizk+lKNq/uBLTgzSGVsmoPTTo
VhhCcOSlCCNau65jtW0cH+4btHiEI9TXqZE0WjP+1JfOT3Ekre96nBvax7X1DLfTg1YK2ceNrUQU
pMHa5n57g3rdA4kfSDOtjzjQ3WRQjvaxxdw60XIMXwLsMgWBiu6CW+AJWK5fj6+X3gmFf8T4uh7i
503ARyHE1XFd/ngXsIKWLB0368W7GeMu4e65wxyon0v7ivkLV5qoTZUKkMF2Wlyn3HkWYhGlMKgq
V6IwFkWwt6mQ4fcphnm1KXXUKwG29O1k1VoAaFgJXnht02SJi/pAU50dSM8WO4fRCaYXkOFTeDuH
tmvWrFVSVRs4cLQDqh/Jw1QSmTHalQRhFQyAtQ39Thj+5/OWF8mVomPgqDt8iWwiVFGDAhxluFaz
nLLodv4ZKc7RSsRNGhhtcq5j7+LLGajMsLL59EZm8wQWtqWUGrDzD6On7VgDNoj5qiIHPFr1Hgjl
CdgBzw2Av5GpkaHD5Kn11dmHOgNvQc9FKvaaN9WjT+JPT5b0sSESnz1PufewuQB5mdByyvoQ59w9
pn0SwSSiHMxbBIJQi/hj/W1Js1Ee8LJh9FmvFM8/gBb2/TJFZTOokSr8oRsVnffRwzcQWxmSt7E4
GGwwlIgCSZxyx62slogItSouqbXXt0vxiZrN8GT5mMgcyDjarMHWS/oWXZ9cZRDHNeNQ6fFj4+qz
7Og16OsZ+RbezYYkcbjj7A44dCgKnRwXc2S9MeAT2I+9t9HPBptZwuVzyzD5jFVd4hbp8LIP2u5Z
9zv4S7kC9ReLZzMi1guMlH/KlO6yGU0CwXfsuOJycvUzEtk8j0mjFRwRy2KX/CCtOLblHdR4zrp2
CGQyULljn2vMxoNcBVal2QQktitVv/oMxff69fovAaMR8JYsgi79MIXiyn+iGvTvymCR+2mDYfic
9KL+ZOmdb8JalS3BO3kD2uianp/J9Q/Y/BcJ//lsu7ftYV+y3H1Pqv0Mx4Qya2+G1g623N3Wg0ij
vh0dsVWkvwWOihRWPuOj3Igrz/5V+Hy05Upi/0o7rOlveYTFk1RKXDrLgus70PpGjgK5lsG96t4N
isfAtInU/i+xMWin/uHbB+GiX5MyRdSiOIquQF7+/Ho9VYjNbLKxo8zDATEKel7EBG5ZdJqvQDj+
FPRzqTJjTTn2/MmEm7FitNuMq8LA4D1aajH5pdtsoXQa+FLiFFmGPEcA1V4Nh6SOK5ZazPlUU6qM
0jQxETDaUDApD2bKkLAMG5ykuGFibbVj2vUaS1nVlsJ8HpRBy/Mja+1jNQlrqKThzPnHo8dJhFSy
NJ+1bhjYIU4HUHBNMrehPzpgEmARGKrwws4xK9vRm5pllbW0w2AyDhuDjb1mjmQ1KuX8HWDdUMYI
xBIk8dsM2Eo6BW3t4j5dmnydcoZmsthOdFuUEOZXZXAnYcrF0kKRMoCXGJceN0XpH4TdVTgZYTW6
vSp/PgYvSUK5IXgn8vP+pf9jzOJG44du9QsS100M/sB5XDg5JIz7WVsSB7ZJv97VF8jC0vduhu3S
EeAtcSbHrUKIXlsB+zaxRrpscK1jT6M9Q9+NYqbD6PZXE4UgNHJxGBj3jtyQfAJetP5Xyz14RFe6
HD71628pJP+xBuL7y3pFrc/dAIZXQwuU7Hhpajtjf8yTuEUt0gJLwaBqVCVL6hTjDnXNlWccI1Gz
BnRERuvF8L5PSl6IvxChaSvQwudHZhCLaaPRg+u/Y0gr/BOEb+CLIsMI3VOkJfQ9PeoPg/1P8VEr
1l+xgeazp/mgGvlI+N7R9yHK5cHynL7JGGLP8ESaenqwFsOCR3GNd1vIHemxGQVPUMV63WZMj1Vl
wyiNm/JoxD1fbSOe/qf6WUMfDxy5AVmyNnZ3rZb8s2/UvdL2Eb6undrt6p5b/9QjB3C4bWsnlrat
JzdIieX0KntFyQRlNx/Euawh/ZI/hfr8J+FwAmAJaVqYfiE8jL4Kok2pKuILbl4MhbIkmDbNc1lX
r8qz2i0gDAXosBByIzyngniFwVWN+nydOutGorWEQzq7vcKnliaHPlpHMCYOabWbrTBWfT/4Ht+H
h46qei2dSlyFJntrhVGRNtp9S3MP4fuV0SmAxxXg2O3ka04rt9IDvLlNOi4mjH+rEVw/87nZr2Qo
V3w3X5dXfWl12QganlYVFBooL8LY08KBdQsDxIUSAuSkEGIxZ27YUhGMarcZd+6iTrjkUiGkbUhg
se0GvWBzKrL7BZ4hhaNnnJsouoOP9PDULlmRBLL0HPPinoJMJH3O1/yjCq8LBaEQVKTTMlYJ2I2B
sPGuXO0V4dyKKt/ZCNE7FsPL96Sa0JbDjK4PE3teIy0dxeu9lcTiU/jpt4Ym8d+VShlwEw/2OCyS
YtTLuWqMetFNiQHB32WsFT8FyaY/9j7mjcTgcSmVsKNjuDQewiY43vMbnQtq1fFVOAz3nIZMipEr
tH789NQttwKZJ+/SvygM4OwH7NldFD48k30jPySOXFMe73tKryp+pWWBnBO7l0BjXRNC2GYjjwsS
FH5DJxPWzTvu/XkOseNNN5FKpAzpHgC6MHE+vC381pqoBNaEmHXt9fVCrfIFLefGqP8otgSjmFn7
J8txuxgznrSU9J2dDUaUSu8rERALNrIe6fSAfS0/jfzKZiSp5Wu/IkYd0YGaMjTa8J6TkvSkLhbP
ywgFfHWC7AhRh69nDgZ/FpdweYGExNu/n/o+Lpw6CIuW1DazIyt1SRAEnvgyLtDsXO4mmXqgZN0s
BkysWyANMPr7O4+fBoKB4kygsrDGmEe77bg2YQ0cUYZEGge9cJMg6dI1QcCK4orIY8qoLPI+ynp0
IB1MAn738KQayBUdT81SKIvmP2tEPsvCMi6Vxbxs/piA8YazWd9y3pJrDJl0eKMeRslEUQHbwQWR
8f1ZmB76ePolLKDIOeVlwMu6m0FL0C+DLj5rp54oclKc+6x5lNVyZj4Rha3/qWS5a5n1OtGGk0oh
P+5albwNG5/wWd61ye76jwCbnq3bMivRUo0W2TlAkNDZLIaojhu6IusXIqqEtoslKrl7rqx27MuZ
dR2hfmKWjs4zlMmomHqMLSAEzL5k80FRDMuFMe+c1b6i0T4BCIi8zNZ2FsUnBMHSVgrXyRw8ZMVr
qvQaI7f3sjqsXboo216728kJGljnfbTJbX6ZoMoeCKQ0J3Tj7ifOdgoJMcpFO8vaLocS2pff6HHf
9O/2ZHaSAnVrxoRsfar1BPOBUz0r0u2f/rK78S7XWfHkB7aV9tL48qHPRw1L0bYlwBctILUH1usH
py6qr/vpzwZg9SIQ16zkEnb22yMMJxFq/01LHh/5kp2DgKCbEiCa29mDJLVTRPNADUJFJh5O/3TE
2YfQdZp9tVyeIFG5hLytWcFS2oUjyQQnclBC8CFCCaK2Qj4oZ2j7/JPHZ1FcSK8tgoitAonwtdqp
6M/uCjYeUIbHMCX53A5MYXEtN+gC1/HpoOqQD2nPh9Amitc7Faq7uqjmbUlwZ4pabXV8zE7iQsXy
v/6blNHrUuL9s4Cv6wd7q9BnlJAsFaWGaNf9or4wMAB/P6zC/g8uTZON37FiUqImFpL7NWDZEntA
Dq87v8BpTgznjSdf46J4628byNcmA9LjUwOxJFfoDbotRblzDbdTN3SKd6tvKiME91euy7qEvDTr
IWlsmIGAiQ1I5Pgaa1Loxq7+x4FUY2wwLkMhxhZs5imv05TjALltF3GPB/vurrZI42tYxqf2BFkr
zJTqlkPdm6MOz9myx2kPCxT6xoFENRREGCrPlmSK9TSOOc9kjSycnXFen+8c5Cz2KPABpxWCrZMN
wiwVPeACIlT2qbS2/DhNVn50HAMG0y4YyqaqdQfxBnYG9pTpP3nNI3V1/ifklgtv8lqGd+aYmlnb
F5YC0Yt1xwGDsv9YJ8VgHDq5xyQX1GJkEZ014OLgiGJE252XO+5NYIeWjeaaaQOhzpPUyck8Kic0
Dx85y++AbvgxRRmhbpsmY/NAK9hyGKQz7AEEp4UtyPv5TIxhnkOpicmlUL5h969lfnfq7t2ZQfGV
xMTnKHuQhHMnb6r8ybFjfICMVHceSuI+apUuw+I8wiGml7bixh5eMJEADxCNkjn1NUhwvS8dUCTj
QcgT0awjBPimBDWs1OA8Bw1yhnYBZ47tdhAFBalolRfsM9qVYTjNrHeov38xNPPzIbtpLFAnetCn
N/CMl5gh8yL1mVg4d3Xxhp/JmWLaUUTcM3KivJB3YLZvQyQoxQZ8vXvpE2Je85tnyDjNLwQ2xVca
YPZTwulvClp3LrRq+xhwM/7zlhaBGM1IviBfaxRjcVBS1i4RKFozTlHHDsdN4LbyoUPjSv6gN7T+
VZlPur1Z5zCQUCI49Eq8JVjhJSy3ol0jTuGl1XUNVpYef0bkG9aeQrj3N/3fj5Za2LsFZoFXKuXB
qxokyCl7NUKYdGC86LJtGordEGJxA3FJ6wvDi90Z6+1+m6Q2H1nJDBTbu6zcECjlWCq38xuu/4da
ABO+WwCXLEmpVWan1u7K2Fn6X1D+MWiwW9Z0YxIGztMSHKBpx9KTCkucEEi/XC4Tp9UHObSUm8HP
ijjtRurY0KWOC1p3Tw6PHlF4zR+OAmjaoFKXyoC5D3ZX+tyQgmepLvsmgFqNETl9p/Sravg/OZEL
D1Cs7mIJaurvJaKfKuz+KEU5REl8P/p+bb1UgxiCLJo+sl3lbpaYwyr50lwQ/gZEMsEYmSZHU17m
O98XbquP8bv06GqeppmXsJlQWRlYkkkwB6Tn6h6RzSYWx3v8eFNWWMJzI/bQQf/I6uCzeROYySXf
vmQ6zTz2tcTP+z1Oc3Z6LaWoKNrzDEtMY3Z98YSl7QOlkJ+VAWuYXp7e6wECEFBzKl4CwHT+r7pA
SX2e8wjiZSsq0baDZp2/XSmqfDhhdP8aJ3yrE3ihsPoDD4FDBjplMrf7iR/1eS7Q5UoYJsMEHgER
DoreItdWyHBobwfRvCLkUlsrxmj+Al4c23PqKumFolOkRP+dku1uBHsg8EsuBPAfgoByBGjCSH7J
hEI++X8AE60SNK0Q7k4jEgzlnp9hXG5tUMEsDDHIe6/2EIaJQioSWuzH31ISPBXb7D0UbyzIETqx
7GONCh76vWw90CV/HK1QUy63rfpB9Tkoa8GLLMcCHHbK+GL1P7gqNtFZFc2rpoiuec89A5414qnZ
zmLmon35BKD6w7iU6MOdGyBbjaVKvo0csFcRcZcD+qFHoE9/03ccRHZndYrwkGf+pQUcJrlSXvBO
WPRXCi1X9BvRwdIIPlnYEjFY1aJMVxl+PrHrlIJgZNy5AFoX7ljj/b9iCbSMXgy3kL1DE617Hbp7
7X/ZPXlNIot8vS/MgCMRvgnSoJPtbFPwi21MObtx0dbbyupmlAWKuS9+OfG5g8mZhrdnyBlQFpDS
DgmrAkemWXLs8IuVd0PSnB18tvLq1VlAPIjUVoOBASbwDN8/40tOOi7MofGEqUR+1608vHuz45il
ijohaoyMVZX6qynVg/n06/YSWmQHO8MofDtOJ4+K+2i5Zm9LG5XRTsHjC+64P/n7kOQGB+iNR6hz
AJdYulxgThaubaD8EoJInlyW2tzDlAfGVzQQO78VYNXVnayWoeBWMF6wcV8bwr4RDXmtCp1++Ntm
I+3dtoFVjn13RCrNHp7akZs7cSOYqrBP5aHsDk8ESykVyfWBGvkkA1Z+0PJwywJsFpPI1USgTocy
orYoleYSY85IUFOLoU+pbLIa7ZT0MXT+2x3hifAZ4ypVG3+Hl/yJY29glEQOrsw9W43wZhkf0MbP
TZ4MW24OHjL0h6aiUVkQHMAu1+PNIQAx0kH8rYSe1CVSAwgz8choGHpvizVVsurLcSJKzgAYRkGf
uOTzj1LT2qV8DWg2R0dBy5mguAigiQBiqFegMcqr23KU/lHuhePAZcksEDAKOgZemcZSm1Ly7CO9
rT1rsUyghngRsh+hWmNwvdSZBypV3jUzvlf+zg9NBEhibwLmI3JVHve+uC85C5MxURMXsVB1JcPv
eqFl49o3ygkXzNn3mqE/gWwchpt4L6XBgESjdrUvoK3qGD7C1b12eh0rDBJXenrD9mY4icweM35N
X7BNu3YvctreAEtdrwdwDVMP0WHJasiW3fx9TY4hZWu9IpJA6j0Vgym6XYlsuJ94YqsD7Fa0VQpU
Gj1dABUenmH8WPbTyqdXU672/8Mcn70RVI8MakMXYEGCbZz3ZAtvWeTmGG/7Tperq9e+2abvnWs6
LPchg0CxTe3cBfvAKNF6K7eQP3Misy7PReSf/RjGFPK5uew0I9Bz2zr9my1EWQ43kSYneMwFCNNg
/LSEQMx5aRwJDMeh1yKmCjGSxeU9/1/MPRZgLeORsAuhyXNxtYBwYR76kRchVORhk9gAgKwU+fAt
Fji1h7xOLu+jIBpFWMmgcYyl2VuE9Qd2/2JXTmg3m6o33jVnUhzcOgTVoB4UQvEhPzhYFTXNuXIe
T6XxNt21aKBB+8KZR1Plcw/kd6TWkbW+/zbD1ou0dOTB3unw7Gtukk8/U3kLzxqmWhrMBrnsM0LQ
hI0gBov7LZ8BBcQ2aSDvGvq2tCrAOdAksuyCPEY7BkkVFZUwjUrJ4Eh2K3DXJJ02HUCyJBo5EK8E
WCbw6FQ6numB5SfeQCU2KbtN5mrL8UVFP8N7/1VutWp3/wbSk/am3gwoXecS03q30fVak3tETAdA
mYL4aFRcrutL+rwh7BpmpVcUj8EBF/Id/W8CayZMHyrMCfuJNZ4NcSg+lnDvPAR+mWNay4emsGl7
L7GfUR4LQzzeuIY7y1g6ZVu1SnS960F0dfI+WEDxl9RhKBf/z2p3J1hJcgjv+8ipOStgzObUSc9I
V6CSre5zqJhbzhEAaj1FsWqqy1OAwjtVjwwm8P+V+CwFUvq6IEXDU40q1ai4qPujCLE+A/ksb1tV
sWriFLIBKtFhvMcZ/PrHOniQ8WuV6ofWqrA+gT2dTwbxZTCjluXgkIDDu6H9rG7h3hoFE3qmvFix
RJgWn6SmI636bjSQtz4KEDoVw6rHivKYUAzakFts58DJfKJG0vLTXz1KPilhduob0X/rCxU7qlxm
0VhOYWZmHQ84mUZqcPSIHEtCi/AjnLAirMllhtPbhc4U9Jj9cKxGpZmR5kyW4n8X1hOEHcZ9yBvO
YQ7cNQH7Ou6G9JLjmq6FS01lAQ1gGgy3tRW6VhHCm12+vZ7ETIJRZko4HPubqybcel08XyxayWsQ
HDEyzMvFbehx1nrXPo7dWtNSoUylfKTujnmNGD6nJ+cm3S67yeJhh+Z0bh4ZO6w9jVVTS6BQx441
Us5NNCUMWKursEk+3tz2emRrdlM0RbO5hUPUuiUkQSXgJ6GPbdH98PPpbPBIgikPct3nsO1tanXC
nJMXJTIgRIzryWZETi+u5P6g70fNxdGO/nK0+Iq/TzqljuxvySTJkf19hb6Hh0eNhvbk+3R7WqNq
cONkZm9ZzfMZyDEXMZY60XskVVhVh0+I051As9n5bB8BBa+LasAtJyGwZ9q3yy53g0A7N4N6kDOU
S/MonqN74E2Wbtie0wocCI58dn+IMMorNjqtBVrbENcORLIcBT23eKA7e2lLkrE3ZQoOtTIbeH5s
T9NOdyKKc5NgvfgxRqu57xzuuQmVGdboULc907GI/TH+TXErYcha034njo/z2u2osFR2Nk0AjIBP
leANXwhjh/zvNjV+teVQl359flo6i8+Yb/uspgRSyls8oNHLF5k8OOyoNzWaiq0iVlSP6XsyryhZ
ZY/Dxjd0tTeRSl/E4Jwboa+cPzWQsqO9Gjiugf/WnW5wxku4JnZauORubewRCCzZC6E7nq3FEmOg
BL8/IQqskoUa6cp2y1l36UuM8YZZMRWZXgAew2utTOt7xMPzIZG6bgdYxxSnWZvUrlOXnmBMDF1I
TmCKlZYByoJox4muFzPh8eGFZ1aYCqUs1W0MXFoNvjMIokwZCkD8F/Jhf0gyvkzJ54bm9SHzyD0e
KYVlI9bAqL9z8hTOdAExzmU6Y1W0M/KrXxFXr0Bf1KtuzdtKPU767X7+V8EPmb8YuQNbV67lKzxY
GEbyJxX/C91Rbe8YiRNT0bdQtWGLffvK2f4zrXzxgURVtvHZBLqWwuz48NMBuyiTFdp0Ddzww8t0
9H6vfaUJm9t2+zG2Lf4KSVbSRvDNqTf6qU/gDWgqUsdTDhNklfFvh6UdPHdilBzfKES1HQiA/VM3
VMua1uRaYhmqE9MLQDqDwhwoMg4X/X77Io3Ue0kglOUUJw2TJuXTQurFQAhKj5sj4Rbda8x1MrNk
UkrzSWbXMoy4Gk+sC4lyfOaI7/n5ApGx9k9koQCNfPc7V3PDZXWg42hM+GHy7XT9CmSnD6wUyOzk
EzeSOraofPulVKRs8x6gjYwSbleMMlNZIR9HFa/9ijYwej3syOVlC/40Bbu2l4D8l/9dgox5buYo
cxqGPjqzBtXD0uo3ZYMjY4DDblYSMXtK1SQ2Aol2GF2XCJdkTkqoYFDkhlrcAH8RoHPoZT1A97Rz
l4FQHyVCe2znsDIazBoVNZ4hst1dIFTabRBTwyLuQSj7DXRmsjwbLjijvWJJ6rO78n2eP4Zprveg
YX/arIGpY7+EvMTMIhCd94xF300Wq3UbhQ5YApt3Q8rl+Tx65y1ZvHwFKfDzLjPbUL4OHL2dJrFf
49ivJ7dFT+/QgfNVTE7l5TXsBeiHeZinZ/91EYgGNKa9lmecVryyr4Xu9ND+1+OWQT/3xNSl2nPi
YXW2D7t0Xfeg8izvf/Zr7jX8aG6IlyCGOTKTwnvSm097x4jMvSpoXBeR+q5VlgNmpNHi3kLvCDym
5xQdhOGN3k5wWb+uSgm5zgP1J98RuRevaQmDrfW77QC7DUTBpmi0HJM0RwyGUFM/rBu6IKzJAw9K
rkPZo1+AwH2OkJ4gRValShlR2qmdQ+cxEWo+0eSNfzLR7DQzgiNpHZsPVXJROtlTZKCi+2kckfVM
WDrg6WUIkf8IMv31V8c8xXpTOF/Z1a3/gfn2nk3zxZRISd3woRxHh23/UaKjXfIPH1olPINn4wxW
wjg7ihq+iQptPacLmW/itEUeTS5DKkKpEng+e+HHO9L3CYcYIsqF5HNHiub20rGYCl+mN0AQLJFD
M0B4JIMsJY1/yknviMmDRGnKmWAxo8gohPBlYnR3ClcCrVgK5Nnd7USRBGjzI9CmO72zS8tCVfAu
pZO/MOjtlQKqWrsoo0p1nfx9+vMweJeLDDE9kdE27WFIiCRf4fSX1KW1w2QsbhUWEhbF56gC0kDg
5LLZ3hjqJyid9faCaNR/gl4R64l8I6WqWusQKWQFe3IZdWT2ksWcBLkSxi/sH9NhVLp6dGXqB7eB
IoTEsP20eGQeHzUVHP/6AkJq+mfHRi58oXGqSm73nTgV+OnRs6rHi+j8nKunG7R60QSwinFr7lTt
isfe1LWMdhURPA6Y3PmI1CNNBOzUEphRnn55eue+KW8TuoupLULE8W+Oc9OsEAjkKKQ/XK/Onf5A
a6Ug9ck3xFxhK6nMjj/YS7KFRm3I8RyZzeVJW0gl0sUJknD6vtnLrH7wG6w64dUSKxI6kssxVU2s
hQqF5df4WKBoBlpKKddVC8AYxWe4Cr+3Iw6QHBtaiiLydE0yk7oDAdhFJRGLbdlrOoBhEumN37iV
rqFAWq9f+Cw+mkO/pENqhh2vh567xhQMaKomdF+gO0gXQSlfMjfw3UN1BS/Wn8cueIgphhh8sefs
eJ/MjRZrqPyVfLy3qEIK1gaAGHWK9L8YE5fCH8n4MU8wqP/ekusE/6kqdT7Th7DrGHzgJHe93Bpy
lC4tmZbNghG5g13OzzrbadvBGqf6c90MDhejReriIQtYgZlY/Z2RhgIUSIIAdb5f76Efe+ORU46A
55UwPbT+WksW67/bpnR3zDaqzsR2+8SXUU+2NbKg4Ag40H2UUGlnlmnnkqqfbsv76XAW6xKD236J
cIzFXrA8KYQoQL3Ul6+1Iyz//+mn6tQCvaLyzhIqkInh4duTOLzcMiaQl4p02uAXhqK6jvaC0MoB
BdKCspS5QkdYXLYnT/ZatCcqkvIO+mGJ2IBrYMZQZuPqm7/jpe+4KdJ/XboiKB7dhWGFSJQ4xB1I
7GCutmbYwNXm4AmBoeRaSdww42bi9sfZr+rux4NC+4GDuCd6OfJDpdb6yE8u9JNX0b81ApmIuPdh
F26S15FF3nwPzUuBn8Dgbejs/Z0SsaFHSnkn76tHxD0uQ70iKYTRTLTryMfc07BbpWtQHux3vPm6
a6/BTAzzdPgmBSHu5AM6JUKSOqqMG8rZs8fMymB79e1jAAcdNVVgrYb6JsGlDaytPJnZb7cT0NmM
y2JXk8dNO71TBqRALdEOU2VuXFqF07HZFjoXfVdmm8672XINEnAVixcy7YSqjzB/dyXN6L4XCukZ
/gXkH7TddOI65NHF3zhkCd84DKRLRdaFvzy9i0Bgav4rRXJ8bnlhCJJ9QLnX9KnmDBBsKEUEDWIP
CzYVjcPGKxSiWHbGIbTWo/eYRGiuxzMKSE5SSwkY/7rNBVIR4nj89QYoWKs8j+3m04WJYKxplraR
X7Ewl/wddnRe2G9EfDRh9pGCGUUJ0/77SVdPJqvCoKAhaach5+A/f+9UmUbW6kpJA1Fut1rukD8h
AOqCy7qyeCYhLi5QQSsRpK3ue9ASbKq8qGnjDIRys1FSwwcQjyxqaxU4HhR8whBTFogQm8PAFp2s
SfVrOoutRTmm+eeBPPFw3DU9I5X6aA3CB96wc88GI/7sBzoOYfpNRM/wQWVKNqiU6i7L8sbomOHt
Q3CeYgZI0S2QiAuatHGRoqvvS+6CGCFxFvgWTEtLZ9x0IPJDMf9VKm/GcEYPQalftyBjL/7ExpJB
6ctaBbQW6/rj8iOqJ7DfefeSEArR3I6vqH8jYAEXS29JYQeNEMEn/3qtKMVp8vId+ZpcoTWuDn5d
fYUEY1B0zoVjNsUFtxkzC9DDk0W470PNksPOCE43TYlh7uQAchaPl7WG5UzUMNAIHc35ZMED/cSo
Dn1egoCPyU8NEb27H9jX+wU61rjwut0TyAdiy8GgNQBcln5pkyUwuy8fVaOCJU9j2nxL0f5oUswg
jym3GUoQRb3+ZuU+mzoSSfU1EODTgkuXAjWDk4nUdBoQL0tA3Qa5w60IG9V2383UeCHovEA3tA7B
kUehgMtsdfOC+CYS9MNu9b2CW+C7L4jW+OCYPxUr3POyngeDn42LMFB29CVR0ZC8TrWQvbiJ/9vJ
OXskyyGVdhAWS9fslpBCwy4BtPn3ksrEYvxBckmhUD+KDbvpSs99HuJFGWa2rpcT4bZX/CdzysNW
ulqS6upWuKOHJB4BsF20+KYRby0tbObdMrzrCAsTZ9Ys6bZi2kXgf50Juu332FUwvivZBjcUnqcN
GD6XXRZ94qzDDNKoA0ZDX5jXsIcVY/zh2ObVxz5SXZ4SLeTmf+NEnUDoFDYE50QqeJed+gSV6UsV
AdPiIyFWY7d8DoLK1S/5w3eEt8hHj4cCItFDdgv2HGOV/FL5lAbRA9qzLZ3jHCV53Pm75UxzR1Qm
h4so99xGYMYeBW+YLKMtIIa+6/fJcJpg7+3fgeJkU3E2rxqMpM4xgCBj1eSkmppaAXhZWMSD4jrg
BP+iYRrnMALCC5eHLfOpPXOTSYPE5MWqtf6TJ4wCPB+eg/N2xxL9PgcALmcgsXLXf1djPpXipfwR
SENouP6b6yGMoefXQl3p2uQ0VI4IZFW7CTDSKFPJwthItWk4HRCXfIuVhfoNpcV4OtBv0ICsRj3M
KjeJUh6imntlJBr65Cet07663XPTlhaWZloTWikLp04ofzXNZ7EbjRWZZ+l273+HtkCQQGfTsx71
wM+SH1ugPdDlbTzB6hDEfNwDanCcNcOE0NYf9RBCyu4lk4QC5G1IZYxGK24/m9DnyLedmUct6CIF
Dkv0QFrs9LiHCyU6pdqt8OKhDMLNY8A9bT99wCRbQ5P680X6B1gIsqpnqhKlQjXSOWM8k1xibm4G
5itc8hFVYTifGDitcBDQ/3GfFKzYzvNTxqliECOAOTlBYQXcZWMxOTvTogsnmW/pp5ba2zQVYm6Q
BzPMfaX2CdZNj3zqx1wrHV7hKbDtyZIxtahSQimZajXJ88hKnWUszbzEB5+MDN1yPUVMOPE+efKI
tvz728JA2HqNrx74Qc73cnA33TovjV3VR7GvHqa0nycvl1uhJLibzsxgXvnexeP7FQBKlVHv1L5w
pceuoUWPyEoeDi71AYlgNBuim6mO7lcRD0wMfYKLO9zD3c2oFXF+EqdMF/7L1peLG6YMlZoiKd2Z
FP8aBpTQjNeAarTPwL7X6c7hFYPA5dqi9Di7qs6V7OkQ1dWksvxcKbWhVC8dhBJeTxyf3RP2B+TK
cFgP4uX79l/cHo9mirQpkZVdJnPPL+66sfOoV/pMmxDjVkmocQf9Tlpxv10P/OfT0plKrYCFRBgC
8TkCQTIA/nOSm7MubBSJHc7Zn6W6bM/F3jWLXDqo02XcGIc28CHvbGJ4pGp/vDBJGKwICH1rTM/s
CA6rAk+oBgX9W4w8xNZiwvikGfbtG3R2UJYlv9k9LEc32cKxBK5wCj/cWo3aGw32SnDLv+cvlzK3
y1jiiPl2wZDfhh24MFwJUJAJxqk4KOAnMDsC1iFSmOV0MFsPUH3kBYJlpVpwCmR3fWnAYT6WXeyl
dlN+yf9WRbNs3PsG6RfRlhCXqylXgRNPP8IJgN6WbrfGLJ/ubZT/E/l1+O/LvyjQoWu0uyIkoPss
RXl3QcSWCRflZpddLp7XPJMXnt+RKFPPTFSvEEfg4JV0wn8sXNVWNfCzRydWqlGOe54FZJOiW8wb
eGoVPbeis4GXSDwTTdj/qDrJy4Y6Tliy6CAxfdJcfUPaJI89bFMzYh3bF5oHJGvr6Xgjk+Rz9tuE
GbEisXiCKeFx3m47Qh5f3wfljyA4kX7DRuWZlrb952Y6kpSsqjbQt/niAknjmwMfo3+DWdjcLU+v
PPactHp8fFkhVxXjtCbcgGzzhFr3GhKiqjh6Nm+89CPscN5OeEqj9oyWfvpjdsYBl8AMWCXxyBLa
s+Bm+4CWqGE1BPblK5e8Wn6GbquAZ2vPF73GN7pWy5fDBg8il2bPyrmPP20VadGFPOkQ9i8fNcVt
B38gazQu5Mc98+3RXAOmbEp7yygj444lR+8l5TjVqZZEO5Mb2WSgZcdYNA0fY6BlN57cyzOEYiUx
fCX0EUyika9Rwb69oshMQZWK6T8h9lt9f9Tfs4dqOMFM/2e0AzIIqFonqUf58J5OBV0U5y+iMKlc
CrXpCnVEXKlnA6Jeb74401pK2AZx2t/mrMIZwlhVOTISXUdyB8Y9YfLna6faRrRGpU+jHJgHA6I0
iz3I3ubMXeRxcVCVs3D4Abct0LMmyX8MZGHWQ1BW+56TUZShGxlYtUrAx6mONXPbgkMo2BhoO4V7
9QjUaCwW15GUTBs4s8CcoATzGXYkxodsrNSvJOvZjJCQp3hYgR92Q5ge+TlmaC0ch5g0UyT55/MV
SaqpVjtqUZc0wm97AknHXelybSilwqXQpLWQI+h5uCUreowLzcpFlgBOsBDCw0ZQ6NRbect9M6vB
2bg6a9Mog+UqPleVhyzUp1BJ4LNX0qS4Wae12HO4GITemnv93JHLSQeH1KVbPOqlOqQDBpGcq4+X
X0vPTOUtvKGrJKuB02Jn3PjgmEXGm5j1YPnBBoEO4INToU+zI1G2EnRDggFFBvIShEHyaUKsTktz
2wwcOlpiQ9h9EKvn08bfpidSShQLUNlXcImd9OR7GYy9BvTy4uupdGdbzPQSU/be0fKeVEl1kriy
7tXAFmrXKUgMNoCG3kTj1qtDrKZYQytZ/Qdu1bXdovNlO/b6SueMuPF/M+5N5MQIntgvQ6fsvvO2
nFDWUONS8q9lrnZp6jHLhVdxiQ4H6EMySHVEnR4Jwf31XLdiLnPWSF9ledjiIf8fOkQgWEA/jjnK
oZFBbBzO6RvtRO7Dv8msmvgZEN6QNohgwklRrd9E0SaaTGwcDA0mjhzS1WJnkXUEDauB+gAN9pno
7eP92EWz+vFskMnf2X5nhhxViPazQaIFqow9Bbwmtw7BDPwofVI9NdptKRK+r+iEY7IybRAlpDXW
F2j1YeFCgtpQzD2XRfx7Ef+U2rVFNaRRaVgXpLIjTg4kKyoLyu2g1wOzsSQdYMXw5Z3xvnYfKVS0
5eqtho+5eXMXvTGXDRHnZQvEgdTpYXBSpuVcJcvzs4jsMBvgJMbK/DAVYFibLxzfz2WYZ0RA2GFi
gtSeOvIlCyOdgnu7hEsa5J1nnXfsAL50ah+kIJGGAN+5Dlq6ddMha+VYgqnoXhLhbEmlc8oPafLk
wNToHrU+6cBqlQZfkDSX6/v0+sIAmPSDIfDvOQ/IIYCI71Zp7vofXN4qKjCAW4h/hhKy7X7UW6aZ
WRNeoqJTJzkKre9t19UJ8kXXA50npZ/43XGpOQ92qDm8dBZhq9c6lZKeZV6oIdNrx3ceJ+RWjQYc
bP7er+inGBFk6+2qBNhzcZW8H2hIK3X2RgTh/2UPUIGs3ef+26x9ebW81Aq7tn55sEq8iU/+iCJ/
116HdIAn9SgEUT0BixrmIcCD+bFDaYkDDDrOiBqVL0QdzExeGwu2PZcBaRVF1Xb2yYbqV7aKck/W
cyI7mSZO+yydOfMfkOAe9zRXpznXmjRXtnW70sKUCf+hbYkl35ntZgkFINDVNYU8E81reNtzyFPo
HZhLU/ofsQqGKHgO9ih1OoCRGdfldZQgE5KkJ6jQiw2JgD4QAAL8uHrLoxjbggiCVliyP+QjxEJu
ftk6cOu7FjMH2twUmAk+A/6YxlTrQfkC+0E8pkIXY1piDpny34VGbSnjZKPZBTWqJ7B3dKDNguFZ
v9buoUQICcZiv+ApapO6Qf/euDmNtb0ZqvYvIQ6kRQUPtLwFQOYdMH+Lh3ercujhoGFmPXab2sV7
HzrDd4eiMRYxz7LTWRahXTuOWS98fVOnUgpGExiXJbmJstVC9qjfgZLx8C1kSlNbEmUWUtxb/sss
VLHctJz6HFuWdxJxe191eLzTRsOdfALJcf5+nbu6vO+Kl0kkDVj+1DI70d3gzyg7eUZMosL4F2+h
an1xLvBn/7FvEjJvnhgXEa0EK6Gh57Rtq5ZQsiW/uF48wIk4DZQeSmp9FwvRsnNby+DZKUCtI0US
X7XEUTDI450/iiqRR2l1xkaEAls+5mtDSSXxg2prtMcQXoyLnfhWN2bDUKzsOontTWsC6asp099P
rhd4OeboIaQ0XKkfxHUsCXebWivZah4sry3C3f0r+e2hUJR219Jg3CRsa4xsjUvNO3wt8LhuOGB6
NKKcg8yCUuN9ViUjKtcbn0ijwZ4x4lJ87lRAfCx4WgzMvghm5ZeHHvNMt4ZPzva+VJLOYamGkmAz
15J2k1WfNHem2xP9qX6eir5ZCKNx9waGrNGRMYHqLlPPI6ewsgtRzwIAal/WcbAfSFgO+M90xl2H
ANGno6CqwKDQ8D2DgOc8g3l8IJ5PQcoBzYzC6YsNdNxU0YNU1yy7KqtN9GpuCFYUUFzMHB/qJZcv
1mDSeNO1uaOIT6NwHYTtAKx5lCJq8iCZzIyDyTpkuiRpz3Y1aPhEgnZaNzvgtxzD+0DSlUo0isrf
Q1kwPY/WLH1FubdXqL64tRn+SBs4AyLyftmp37qrCnHFsYk0g3ljgxZrL2xUfx7BO8T30hVhWQ8b
wWKZzl9GglQ8VNGjvkCQk9Q2/RBgiWkfNGp7dn+5M+iJ5Wz821dpU3A8SraW8w2UKLHnnVAf++eQ
FLOXxD+sXJS3nENx/8hVyuvVTNl8DRQ8rMdyx3soPeghOfyWWZzSjHRQYoEUeC6zC5t4ZkJ9GVFc
xT33lRlabSHkkKJcaPvm+dCqOhSq7i1LB2kuc4Qha/kD7peimZI/RTM8iFoPs8S90JkJ84P+H3O8
oLNWIIX6WpR8hisxgYgprem0CETjx0SFtipVKzF+uE7CTvYmosCt0+3k1EbHWEQV4xuyd2pRARi4
MYD+InvUxTTAotuks5IFXly/x1HYFwNqWIfF0A55iPhG260Xo0MfvZk8OoT2o8heO0O6CCiF7d0L
4MaPaRwWMHG+AKOkKvDU+rah6noNJkGF7AjQNZ+CmepsG+3FOLsldfVRk6KKxrOeXu9Ad+syipVH
lWKAz1i90YIFo5c+XL31XP1XTIAU4toyaW+dSPbuI3gzKG1kmOSyT/hQYOVt/8T+ZPmj19/VzDR/
B5HsFS92ltuhQoOVT0+zZOo2FxJbWkHZzeaT+I33Rfhdb6CV6kWnBhY5duDoLgOOxzkDAgQB6Fv9
q4Z8d6RhOTnGUwwrhTBX9uhgT/thXkNPG4bxzikm1g8qUS0im6CQw85i7POxt4Llk1MFzx5x4rFn
pFGi7PCBhB3V/GJxxW2ZQVkdiQ1cx9aX0SufjpaOdkHohkMHG0KG4TOajc8ZuONwQ6LY/oeJImlm
99xTaHp6xMHtoG9p8omc4V3ggQAIAzdqJEPZseBmHydt1k2A+27k62XNTRG05K9LL0k8cfBNN6Zz
ZkaxfjU8ugQzh9QPyDZv0+6pGLaJBoCDl3lM7njyac6tQXDoLXphSp4G05R6b50pe9AnpAY5DH7q
lBp00xEM6fbVsTIu8Qnj0zHwTFxOVLjaN1hcI+I9xppsJCT8mi9kZkCqaNdi+5l8aYWNMKdBaooI
jVGNgFVuXcGYEzAUKzEmxq+rCdBl32h3e5orHkHxebzXLbb1LbiwhkIdz14bwWyje5l2GUkodJ4W
Pae8fJ5Q8b5xO2MX+IQ2ZH8Jz7P4V5gD9OrpyQFVGAfZUibtZZtX7D361Lm/RGzsdZxqNuLujgEL
2AilefzwO9YjM/3qQwjyiLLI7+zkRR/YKydIpLfQibt80uH8B4HqjgmjZaWlNLlYs6p1g4FsC5SY
sC6/hmOsJufUS/513iCOaj9U8Xn4pPztn/Hw3QlDkhvy9dr1M3LgyyqPAeXZ+kjMh3rGl3TCmYSN
0q/X4dY+5bWa7F15SPHRr/s0E6OyRVTcf+5OsV3G52ApsA+LszOVDKKHoDcHAGECgBjsjcrikB5s
M3nhzG/FdFyMeqFooM6jlHIjUcovBhJjfAGvVBCI+rNyWBbrAhrQR6hhbaTJfaVLQvRHmoOAzlOP
HADXxKb/s1HeWttPsJk74tR6U/lCqvdEhQg3E7lys3ZOhuKPji5r+K1G7KNj2EYX5B0LTBslilY0
BXuqeJFdBx+SjBgYmXurGV7rw958deoYjXqZJfbr/gy/kp5cL93gUbNFGSKvKAjQtWAedd7U8JYv
fMGY0RrU8uxzpOPn7gfxWXd3LQadklVlmQwTX4KndpKh7UOL6RvLJUOGvgoFvE1Jj9C8b+OplCyk
SQQ96DGYBHcWeCzmlrO42PsTl62PH85UwtrXQFV7pPS35dWcSk5lJ76Z4oWTKJW6P+HZdhVOFrpe
gQZCIOv93zyJfOumfkxXd9Vqt+2vx3XsmjTEtEf1zGzW7S6zsQUx7brxA4cZBzf9mdEB0DjKzITC
XeNF/N4MeSQw1KthgkX9wPq/UCLMegetm7KgsSAVnibi8kFLVKATAZlm9ImwRuPjniJbqHT4lbAK
Xj7pk6mTdk5eJnLODXjUwec9lQmCDzKsjMBSb/Jdbkszhn+Ybh0Nr3HQTLvP7eNiyfXl/ZzJg9WM
7hTyKolAV/vQp38bC/5z3kCH7zgJTZs7R1iq8tuzBS//VrSqlPTxaDDaroMhHZuXt6Lp8B1H5/tr
0P37NAgaRbLboYJDYjrXdQrZN89d6qVHetk/zvnwZzpOkyv3w0T8M3l69bQnz0svFFmVslOqqfuv
e9IXppFCG2jYzQoHFgUzrMaM0s0qyL4XLQnMK0qhVk+zCZGJQ0GaRucaPaJHAqfpieRQoTNT45ZQ
9eph0ct8eFj746zDKZU8K9YFIZJDRlpRjqQHbQlmQ2P4QhpLZEc37Y1VqaZue7IkvVeSxMD85XNH
PTrab4kbgr3FHn5psN1Ws/PQ2NgDxYQ2sZahuW/hebyTgjtnXsCHMv/bejf1GvUsIAmWEMbxJLpq
WiZOIFvIOEWMoFxKuLbxZuJ0adEE3wkMvOUJG9CrUv3DGWgP7cdsh9gltIr4ZSljnydi/0/uc1yC
8RelcFyftTJQv+gOQ3mAk8OXnZppolZIG8cyeZQ+WqPb1W9FNUVHPXZOWmVYpUiOqq5+KRQdVtvH
8j/dS068908ONZtA/kEmaMnl9nhYJ1Zmrk1i7Dmx32QFB7vbwljcLpR+wEjU2OecJf9EZajJw0Y8
1L0zXW4wzAYk5mKayfMF7Z3tCLWRGPf3ARxw3nX6MrcELvkWSsl+FqQQgK5llqOXeR/G/hJDyZh6
0k9d1RvLYIwa1EwFquprwpzyN2r/GEazVQ8dkrc1yQBj1mecB/99+y1sNp0gugkhPdemfNCKskHy
xifyKPd+Qrj0pD9OdU+RAJtQAcsGApIGV9vvn3vVAnBdTHs6T5MgIuX5IHR/CEV1gUWzkXaa23es
JcjMq3ixLqWUKLtaKRzua+FDzcJUHR79OgPakWd5bhenyKVwP9yKeiYFSGiJcXWZXxMTZVGmX4e3
Ulb92GD8mtkNGaB+hoOFfk4w1CfyAEmTpEblm02vEFhosot5+/OMMFW6O0pumEHScq7k95EhxSe8
f8hfOfptXPNMZje2gGppsT8PehGCdcr1nAufRp+9rpuYbcENITYBhFnt9+Z46aEVIqKsikcpGiIm
p3ZtV8fJDCRw8fDHhJhSAxbyYuUcjntm2xzi2dIEw6RJzOZjh1TpIEW6i9WVCjVrNidqSttrvpy9
6ac8sPkGAOTUA3bgI38aPG/YKLA+go6dYAM5PHDDs+XFTcTsECd+Xs+yiiAaZwYFWdbgISLJuqQn
CKf1nRkjz+XFAg6alhiQwiuMdQOazHx3FydlLCXVHeEwYCBNbJZG1Msk8YtO8hIIvmiCItgREgCm
4ybPF2RQUJdG3SHXZXyqGDemV8amAZSrWdjlM9qfncof9FwhXQyeNUdLu1WjSG5FNdyXBnkPHp7N
27qNMvPcI/bE2CfsdgsuohaB/uXcoBaUncs7FUDAkZoMSi+E0xRUH5wpt6TE2NZHx4WcK4sByWrF
gafy7yKMYosNVkdMd2KKJDTF6n6NMgjVg2u9whSoKNifK5gSQmguPL9aG2dsdzPtFPMIkl8bjiZI
GEycGQAhNH1VLVUTHFQklgldhGdi+1485hLBd+BHMyucdaNND844h2Nj54cIQ9yqtDXzcsgMFTdt
Pgbs4kZKT0AbnrvjXgyzaWzaqxnG3zJrXyfRPJEzYmEoYSom1YMxHVzPBx3nPQkDcqIJ0ekRj0+p
VwUJ/Y9H6t/EEeUw4pvz9tFmgEj+ZFs9ObVJJku6xGMpAJKKTNF9yFQU2nMrhw3VhmF0ylT1iXgM
nTr8u2HKsxBX6SryUr8HzqHplVcTB6hVxZRJNQ/r+Q3P8mG4sXQf7gmq2c6SjOP3783T635CHhRR
cncPXuQhN29Ijd1iS4Hexkwzi8h7s8gWzaNa7poftEb5MjsKRLlBPAIYRuV7BZfI8xwrAAphZt5F
Rff3F4Tlq02vAr5+HW58h4b9flt0SqzHUoMkbkQqXLm0RMFVURqHnI/5ScUsVzz0dri0SK4PderR
6LJ/spPyaHYS4oRaJMlExoZn9glylRQURr1qNE1R0jl7uADzRX+6diVBbX1U0qbUDHwN4tIXZe+I
4u+fbePinCKpM9im7FLDj2WOAvQ4iUmte+tdDCQnTC33ao/aKYNXZC8ZE0Tf8T6o+aAmn+focr/w
22wyGdNa7mrg8BnCLo4G0DZ+o55cD6yE4DUeEpOfqk/MZn7a2txie6vnsyJi73NF1b09aGdxPgTn
3fOdYdVpoNpCGCC3a0oNQ8nXRlukhSZ/kDqv1/YJ1NCJLNFaMbDh5vTL0CjX+1gt86/0nu9Y7+1q
ej/3P4nbrcMkooFBeHHZX2Sv7GKmM/uRNlwwvtH9CTEW7EZyXk6V/HLTQyo4Oixo2odWJwrY92D0
qq6kbqkHxMOTiMd9UYWGxpULOlpyIwSAnH0wKSUy7U9X68Hs5j//nZX8V1USSB2iNkE3/qpJuRFd
l/xhFf5NRlK79+SkgI2elVZnJObht+gH91JArsQig3/qqjO/NFX7PtEWwENUsTCoo6zIfniZQCS/
JHReh/vQWyWyfngPoVKmAyv8pn7iJdIP6ZOt4/dmFaECDYkTFiXjicV2gKjn6I+BjTiFyza7Ncvo
2BRvUBKjax443NESqP4ct6uFxUSdmQZA0mcl1UNepcUi6yJVuxtCV2SSxzZnuDKUs7qyJRr4MXXM
EGWX04GcbpR4tbbWf1V6vnEcyH/UNcj908EKVPz4+YqPd54J1rKlNCLNe0I6QonTYTJ8Rx3eIBSL
njQojOcm1v3fOgVfkHsJbTd8pGcM1cUgbvr7P+mPG3KwmOq58uldOUCIybWxa4BCXWzAWQpT0/vC
BungdcaZgoKYsGGRLw9RbhW6iCOckMv1sACXsDmMEvzXaopjbov5p/ps+/LgJh6QXUfzOhintr0J
sigmdKJtCi8SnijeFUtBHF92tj1yHMThXTqyGdhS1cx+sfwEe5CMDWz3jirnwdpLimjZVtdvExOq
xyhM7olJkw4VC4uvpoWuo+o1mKf1Hrm6kJ8XDZEid4BDSzU6E8t0OOHE2Y8RBSdZQyrmZenYjgoI
TuRuNBuLefgZg+QmFitLn6/XHZwLR19q0Xao26MdCd5gvP6J//qGonPRjlGlPDRc452TY3/EaXcd
geSJe6d7/izVnEth3uJws9UBzSE7uSmhH7Ft+JGGGnxlE+UARD6kixrIAJtuzd2AIq2erVdqrBxt
IT4bCbaVFELh+TTh1JuXuD+k5iZl4WBvOWuUTyLoj58frjG/89FXHJOsQEFg6I+wHKC2cVEAbeiy
NstnB8EDQD+7O58/YslZzDsimhNhRZPipsTKLqtv+Dd63rN67SZT+fYRaMMPFTPRAZ+kOs1OTx7e
Y9XaHSX3vUmceAMlrz4/y0lmcBx1rSoS25Pb8BYVmisHsjswsXxRM2MtiigtucqC+vawP63tWwE/
j13ZED1Ks7Oaoedo5LlttFLynD8O4Xp5mG+76PXjxHhmUZqJ5Dq8k+rxe39QwJ6DXeJeRTYrDx5P
b0KIq3/RZNQerdcUNOXN/aq2YoJvfPitdgDX4n58vUQaJgoSEizFUWFjW99noKByU0WDorraU8fu
wMwE1vMsy2R/DGmHtXd8H9gxQDefMk0APzsSflphsqG0WDY9x9F2hV8VOk1WMUH7JNcGKxr8cKNq
rf+zqG9PGFT4JtOwBcoH0OiMFrRVFsoow+RIoDI+ld5d7/NISdeJOwmg2Xe+ARdX1epsBHm+GYdI
wobw3yLIanPvojD81zcYzZWQS+MKtu55cpJqhBSoTdYc6710PAhqEGMr9DodA6v8VpjWUe/RECgW
Vk5m2ODsOt8+ayuV9mqfNjj2RBvedYwZym6Ypsnl004EczoRemvIK+uoq7XxI8l1gaeIYE72Z2n8
tlnbQxV7JGS2oTdaOQ3MauW2VgW1FPFklz9dRTEuitaK73JJss7g1zFbve1bv8ow+MP8tCnfbMT9
gxFNxfbX1st9c39NAz2RiGygey4ic91mli25y8Xw1D7qSdX6I11ORjMOzLufksgqKgY1Zg+WDMLL
Lg/xQ209T7rnjpvKNvyd3RTZychq6/yXx3nyJcjMKB+w6XHxfLngYv7Be/jlW9WDKrGaJOhDk5Y1
KjU+cf+zQrztvynRO8p202HrJHnUQV/pZFh6VnW5ZPRQS6DIwbuQacayeqK/XLDMCg58my0w+eDT
VGY/Vgu8taNSFUaVyBdz/Hg4r6jRTU48yLmGcOX6ny6fLGSAuPIhqL8/QnA3fd3bUKasemsciEPo
rPuHd8hnVreU6Acv/1nZ4l1bowQPc3TnLz46yynasAhIXIS3vL5Ucih93Q1VcjmJqUU9nE84iOI9
HhK7oRz8Qns9CNhxOgidVjDjD4ytv2jbhGVFStVl+MYsaAx7y/t1iHrhOhRHhhzlMInalVrZzN1z
QJ2cy0p7q3HwvjQ/Gim5kICOXwuFwlmeBM53Blv2ivujblH8dJtkcKvwOwQ/wZqSoqL279B3NLFr
u8COaTED34Y0Yv1VsjFe6yw5csqOEPWUiIU8bcjE7OVjyzz/Dx0gVPfDqrbb3jFbqYybxO/wnlW6
d9hwW/ZfTv/zfqgiTH7duWAghEizlJlfOmUk0vwJNNNMzf43FwOBAgICvmqbfJ/OnkaFWTTxv7Q0
skwyLeu5JOfNQ/oIwqSnyCYN6ucdIOW3tAbmIYrYl5y+wXlQe8or13DOJ4xKkL/BMck22OprSznF
Agl38gRZbYjnwKXWQE5B4IOOtCiDcy9+uDwdIM86C77QOEBzCAkVZ6RTipICj/QTYeOct0ftts6R
7SjVVSvX5R/HxUqxWN9dGumGsoOQRtYWKQjC2mTqN/cVZhENbOVIE/6RaHu2s7kW3nQpJUH/woIR
3dQ4phoyE/SNDmgaaveeAs9yvR6ft5EmTpKVltsO/kKMPPuVyyid4gR7XtHLT0PbaDn5HGPzlIJa
K7JYhbVcTY3jjcTTbk46RWOoYwO/YC4nyk1Vpb7OmNsxb98AsDz6sSgsK7TTH9im53/wLDY+cc+F
5B2z5A9cn/pNKtXO92GhOCG8+Q82S1KJk2wttC35p/r7s+NsGEZGiEfPJX1SOPxEXCtrZuwHOlag
N4xYB97CSk+DpUHBrb3N3PyA27g4BRk6zlBb56rZt768gvmraHv4BTgfIwS6YwOx0hr10faYdurs
Wl45k+RjpsEPfJ1A0iCwHTtoiJlwVt7+wehGo1T0uUFRenPMMKWji1fP2faWMWdB33U7VIe/dNWs
zQwyczClfLhLz+lTefALEY6qyYedDkwooEqdQ+GfKjHpsW7lMciTs8owc6QtJzvEHI8IIXRbB23M
1wN7AV8Lq36yyLPVSbHACPD16kVijujXaHibE192BLyTZx5iPjXsKx1LOBl4LD56WThiX5XMAWMt
duDPaXanterc+gtUFaQYsZThATIIlJxYOZyyW6nOFQXDMSbtSolakGn6ICnEKGLIrsXNsYtSfByI
O6yJL5kM0s3HbL6JtC0J/oJSFm2pTEjvHkRJh1C7e/lnpny6dmaHcpyRL/aOzpv33oEMMnsPpSFB
Lt3HYuan+yHYyRL5XRQ5iwan7Ae1iCYuwUqPjZrCA78u3o+QhOS1YUafQ2HsnWjTFf8H+AUgRl65
jjNHzYBl6xlr9U1GJqhMn1OPso6X02Dt5n/FbsfOhgK/VJNOZnkS3JtzSoIdFleIksa6wirb1O/x
aAv0PmnQBYZRXOlIN92d8ykuRcwkajYn9hm5L2cc2ms1lcRy/YZpYxSbtbXrSBy5sQ9Xkm7JUHol
n6XYzPN7wWMweAcFS82JWulrmad3mBGllYZGRyZejB7WTYHfjkx6Ie+n0G93HCizw6Yll7DBusNX
qgW12UzfXat4IZ/sb0sESM17tZxT1JPzJxDO3x96my6DHem5zakDriJCs1/5uof9i9hXReZrMKUz
mJAkxmcAZ3o2YtIIQwSi9iVrz2BEZr1BC4NcxT7Omp2INDNX0qCqfOBpSCq+H1JRUDogsdQEMsyU
9yJaD8EF4ExmbkY+YS1kR6sptE82/TozWJ7VEFFL/qKDNMMULy1LlOC6DqofXibJ9ET3QI+xQrxY
8NkS+D5MXUHAxq8SGqGedSuRv2dyRDFM86i8hUclWwZd0nfJH6EQUEJcRFL6YHY7Y3oCnmAuuCfW
2KxFfqaf7yVzsQ31HjN6IY6ijUFoam7ErhSzsojEGUdGYxXUfhlSXXZWRhq5NcMGXbw7UqHXt/ax
vMKfMRj9rH8KVpaRVC567Q2N+8sQHHiG4puWPEUvLHX8TlwT25iBIHHMLILaCoyKBECUZ+qwQ2II
kpTwFgOomxVkLlylOAKeX8JB7XmBlP8l/yuD0eQVFZk3Fc8Ul2K3nw3U69Uj6irZ9At1BYMUMw8U
5YvPSRDRwHMpBo7wgfyMKp6C5ODcoHSom5W43oeJk8VzWNP9P5nHQiGbnVrkXk1YPdHa4jEk6fMV
pnWSG6mVLMIQc7DbsyT8JSy6V9fCMwYfP+7YQaEKXnimSKc9pR+8nk36GvqnCqCKEJ4GaH/CqZDw
4UuF/D5hro2Hb3eSk1cnTbD4zCYXB+TZzLM6uEOrSvyfc3kflK8mgqmwlMC9h+nRnuBNBU91oEr/
Z8Yfq6fq14z7m4kM/gfG5PStB0zK52LCF+NU/jytVqbBB3sNNRxTUgIfFyF7kYtIYNsjEt2D24H6
XjwQAKSFAqqr8xBe97NF3GLZGAiYhy0el/EcNje0+EGmrxnZm8l2wF+9p8zASB30YRhRXC4sL/qw
+2LgCy5OjrdT4j7gGv8e5R6ebMh1zG2wWepSqItKMbjoLB6vqucDDUM8zhtIPbRkKrZ5XWojHj9J
z7U3vYOLldhmKkQs6aPo0LYlJ1l9XDwLuwZYa2vgoPL/F1hnKDbmHn9rI5nFMB5DnEfEtL5g/s8Q
ppTd95xziwXuzDYB+e1/JuMrnIMIf8W44f5vLyFextQzw8BBVFl05ivV2p+oqEYuq7YvvFYSjbjI
fBfThXVpyRBX4adlJg/lHfF8jLWEMy8LpSfIKMcWlf0Q12oKOVcrDFECSfRAS1qX4kVkkJuSPPeB
sduaUup0cjUbO7mGeV/S3JJjrG01r1DeZGvRFnIpyy1E5QjnXLS1eWA8zUVus0I+AI2t0st00JeC
ct0vDGKHh4qMSF36PwUAExWJYUENKvaqr+Dz/GU5Wz4VZaDmNb/J0tjGgFxeGFsj2DAu6x1YLy/D
lOs6RFST+BY93ETOUEhmkSEez86eMYUxcQ9KKegJBo5/Y4oSalK8ognS+2ad5I4gpGttS7dW4Zm2
lMUNpgsntAx3UTvdM44f9QzXggRxqZ75V8+ALPmpXOBZjMdEQl/4KP+WKNYYWM432OxWOqU/0Imw
vWvauLvF2zaqkfef/cGIG/zQBVm/kc9RJEKz3kBGY/4MfNX8rhrBQrlZWUD6xs4Xio7tcDSpIOiw
JqbV1nTCSMs84059/k0DauBGAh0px0Jt31BhO25mI5uqV53vJkh2nrM22wHhkuTyI1nchECS03hp
pb963DkwgtXs7ihpf6tfX7Yw4gvckmXz+gHV5h/NT0r5JYUprrVrw6fFSDoXjhV0oweaInkT/cTC
r88zC7Bp1bNBenHdoipwV+JrHFFJlNSsOB0Nu88nWWAY1Al9prpDH65Vl9GG7+l04CZR8MFydE3m
RbUtq+bY7tBD/58NE9yhWuzNrNnQH9ipJXg6cnYXdhBvU2+T87pwLbIAOyrYPb/lIRcVmsylPht4
P3QsXv7wuacVmpwNiTHcbxfrvMCGll5sBzdLXKHM+3AV45IgoLM08fJaqCu37lIqB9G/zqSU/qPU
z8JqA3C1ehKTkES4ebkq5PDYmwis5yc14GNK9JBZSgI0Kt8YN/51kJkRDXZWKWYfcU5hZD+MYxLZ
o4wWAVUGAfcBoB0y8OniDR1VX4Yia2tFVmJyQvqYzQLffm6l4mZx7U5pgugGoNoe/zQA/CsofvFR
vjr3/dgXr3hxG2W2yUHZabPhs0X35/hvgXzRb4iMUNK9sQaupHZnoMteANyiuGA72DaFJWQWNfwP
jdIXj7k0RJqk337C/Xr4dyjODOMPWEzZCi4oBN4HaHYZkN4Lyry09TP/O+giqiq5duKJd2IAaMpJ
3XXXVrVfbhjeO2KYa1q++cB3nvLFqwk3HHLHijOFk86R9vu8agM5TTysEE5YDG83chcuIVHOSRUo
55bXBHHCGW3aNn++B7OU5iTEZ4jpBAD3OWOib9Leghq3hbPHgHy+0aECAmVD/JajYVY/t59k+dxw
vKu3SFaIrxaZyP/gyUsLcKFiGMEmQh05s5u/W/21NdAkLfbALehEq/8faCpjuDGJpUGW+wfT4xOx
xLeyDLEWyGAoq5dmUPEXaRmo2McmT0C7RQXE1uhhawFUKEG98h+pRSyWZoym/NaXRTMqpXZnTZ1Q
dHzYgNAgCT+JhmwogIbQxbM/0UKIUNvb6FuXTThRYzYFvo6x1vfM25PXoXpfNssDtOPuqVhBRFsc
BdJD//HzkD/fMSmWRZHtRy5pEEaZ0NYAUdfO5IQ9yeJHVqQOYKvomjn1S7+qwAeFEVqm/dSywIPV
OvKRVPhzO0QUBUQZtBhRTHuU6WqUybEqIMp7QZ0KdYKLFaCnN+pYfXTBveyxGbhmqlPQgKRUYHoi
bN7OX4hfPqJm8gcbh1A4cVNpVGlRS9WOXTmdt9yKIdl2f8buQQfQL8Y0xLTjVgRMwZX63pea8sgB
YDdYbqpxvQX2nFzP7ZyZEF1yJwMEN+mFOfwuc3uoqz222NAP6w8R1Ib153nYMTUxGjUVTh1iaGxN
VIR73OrVqj5wk4fnqpxbVp1P7RYJtfSAKbH10rvMHsL81QM2qFIBJtjH4whF4HBsuwdO47ulDWeX
0pyl/mpxTT30JvlkXAxdtOudc+y3VT8+4dJpgecBvTMSWkfS/87CoTfbqfi2yPnc+oHAaRdwSGyq
0faiACAlmoxi4nqN4GsiXKGhCmUlSZ4DUFN5/sN8xyjkv7Ib3jiF4hW0Aw5kzHMNzAC4PYhRFMIT
30O8LXyYesiy4hEpjKwUtzkY+eWZT/utJ5WIz7WRkc1efnI6vFyQLe4wv+PpVdihr5b4MDAVOHUH
UJJ1d+rYG6Th0+o34K4VoLdG9T4hLSQ0j+E8338F7nWOjGuhAO3ZJlB+ACML+U8WV2z3ZqdvP2Io
JyNTrjg9xZJ4mcpL0dUaGabYI+sFMbo92ijFOkh9EHtO00AKsBtuqNl2zDTgNDl4u/EEHsXijJH5
SLYEXCfOO/mV1PdqEeUc4M4LkAzXKEs9CVjgdchRzdQhMFRTGFgUxUSKHh96BC+V93D8DIEUIVJy
N2K4HlKYEO+xjEGPvH0a9gklHNYQV/6067eVzoEDQfJffzoanJvN2WGHFDNMX+TQTKXL0hXDkwgc
vDHJZkQZ927hzZP0cve4lOaq8fkaGZO8vUgsMDe/WoFnpeJ+kiCWfei2tX+nbGXS1WqiaR6d2L7a
B9tBzDWEjy6vFE21W70BzwrG7BAu0B+OasQPPGxsam+cBfinpofeyjlrXtgyT10pQ9+6bG22kreY
i9eZNpXjbdh58xqBvtZLxk1KgIqvDUsKeLsImSZlFlVoCSuJQDSIdfNOdAjA1ixnTIInKAXrrcXk
wn44Sicdq0w/qdwVuiinYgAPSe41yYAX/V7IBSQoPOcddmAKRnOMl4WJS0hDNUkoK6+zcwYonkM8
TAqbi6halojcbWcTdLXQ5ywGT/XKyETq6AK6xZ0VVtjCXawMsqIo9P3qvMrbCF1oAOQDoFKFrP+h
84d+RYSMI3k8frgdNiU9JYDvEOgE8LTttmnRFRuuL0d/n2gqGaGkcIzglckmGgDDa4X5CddBerbV
ABSy+HMjxFXVA3YxYMzdrBvGmKG2ggiNVtQQ1NREZx0i0xANcmckF9QRZtoUHxiFXscerhTw4jdr
lCzAtvH/0Rv5pJwOxwWi/whKDDgy8MDMIJaEZzr0JFVbAutmoAYW6sXT11ocPc3IgRc+sUtAEXs/
m5fFTluqlSUUro5gIL7Xo0MJ831Jyshe5XysJ/7jMp0n6IRrFd5NWFLGxbn/EQ4OumEDfiiJi081
322BAauMk7XpWk4gWHW9m1l+fl2sQrHdn1SgtB7azNueo6CC+MMyw4o4RXno6Jrl13VHPtoJJ49G
ru4fsLnhikqHqas24go5UTvQ9bWtO/1RwVfjJcLFjU7cgGLJDIx0Pcs2omjJxgzgXiudp8/GCz+U
KGrD2S5zbkR/tpBtlcby7dh9/73PREeVN1rXp8nh5M2cQy7jcBAAu887lXrcj6G+5DEsjIId01li
bI6vqMjIJEvsVC8fzpvKR5vrohMF4ZJoKkNn/iCLVcFgfo8weJ+I3iHd3J5TlHt+Vwwz4aJCtTuU
ZdEtyuqV6apJ6FVyZegy2wzbIE6niiK5V1wu6jKTLYF2uNXVxJVEaUC9HfLThnujtf58w91lJCms
gVDKqVKUIPym/B/7ejl+n5UtI+0ZBtnkT+aD1GOoVQnMdOvmMxMSo1yBuF8idTwA6g2jLjwdNqaO
0Q6PxS6kDKYjtbpmgVD4X8jkgw+Li6dqXpfMNNLZMfNCiysP3Zb4/8FssPX0OD3zZIhcbwbAcHK0
nq5INqDMweSQE34fPDFJEUkwKzntiHBRruEGUgoRUSvVDzdejrug/XTD/hiq4FWJ5MjfB9claEOR
2xOlznmbuWrEcpmJrprOC2uuWbcdL8LJ8kfY2WzQkBX4cwGZDbAflAj9uSg/kEvjXFvFVLlu3w51
ZVvwI6SghS2/CjCUkpn0MLXcFn9xjqHwndCGMmzBchg0vSYJz9+R/K/kWddIre83Rz4Gf3KiEd32
1aGJYmomBNxS+lTRVbi6HHsf5Z+nn3I054mHCd+2+oycNvg4HQA8xOaXbi/bPaCpYmZJwlm9J/6v
WKDsBHomlDD64b8j3HaiDGRI6iLGj94CWa7jc2hHkI4B4visztkvWwrNGJmIjq3C+904R9Mg7o87
EScjKByvgtGHjO/qoHeKDJnpVZblOoQPcjyIYOlCN5fYRZYhNbj9Lc2AWvl4YoHtDhrr30ZSFf2Y
EFHRPqwPJkRfGll6nXcMsVOdFibJ+OoWpBljDIrIGopI3x3EkxndQy/vDYl1dKH0c8/poZ4tqBas
ajOfrnR70KDGC8wdTzhiKUnHkGAfoWImr/hX+GP79sqXDkMKR+D5qvTOTMKysFxDigwhgPaOpZuU
/819IBY13hntxPasmpJXEagmtG+eoW9ocUsFTaaIWWJo7Lyyh2rIDGpwlaq6quT1asIVvgD0bRTb
RpnoopoTzKZ047oi7E4TtEUTDF609T5m5gDpWnj7LSA9xwH8aoEaNhNrvivn481QGX+JERCPNcvu
NDypx+OJ6H+8SuYWFzfFF0wMMWTKw5ZZK3rS99y7j+tsx63yrqHD9JzmV8bQ0qYKBZevf9rwImHB
Ojy5WgWy/lUHZlllJ6gWWAQJuUSB8LkqA5F5CUlQ4d6IONPl1MDXW7MgZXU/gBa5fy1X7uYSMnRR
x0GGeAyrr2sOs7rj+QIYy3KvY8o49uPLL4Hw5kE4IsK1DWwbOS4vMZCOnpDDve4yfO8f+hz2/aM6
J8Ohfra0UlUIDUJZS0atAQ3vgsS+VvmB2Tm9PlqCAFGcJlISsazbW54CJN2h+vgIcyHkl0MzjFoq
JvV5sRiaiXwr6QtfYamV4Xf0O+Gsoft5T2bt6c27BN8VrBbU+iUEa+YxgZTF6VWR03/lMFhjmxf7
93WvzmReAYwUDtp0H2rd9zMDbAOL9yF5mWngmNNZI2ET84sSNLPDeTf76qjXNtMnaUDq6cG90QIc
VHzD25W5Mgo3MEXLQjXjsBJR4/R0JEWHYdaSyuVw64FjbCSPjYn+oG+ZeWefRxOVQbK/UmitW24Q
TzvRWbJOo96g4eJhMHEvPvB1FUTephwixM6YDLLIVluJhdZ3ZezrDr/GR3QIQsA3MRNoZ6/FvQpJ
PePt+tZDUqd/+Z+6SdOfw3MhE8nMAPVoW+2wE1KLmQbzHrT5o0cpIcp01xGoyY8B1X82ZglAYYtq
Q2mV2pn48m9DBp/5j0ISfPf3NdnCM08Kq3R4LJExCe1m5Gt6Uo8OREwvVJkXdMaxpnry0YfPm38M
TWZ7DzxxKm6eKzvdJheNQV420AErm9IRhyI9CW5o9oQZMHjWJiVqGYc5xBCzgthpElG8Sv1gxPGP
7uNBncr4xrGxVZdGoEyJygItOXYkUmodJ1ODBASm01qVeSB8qFlCVV++ix6uFdP/GB4OzvQl2D10
4aVHC2wzzohXL45/W7b+BfMIgGQ7n7MvV8jQCBtGGeGfw4mEjhnCRtF/7mH6f1Ol3PYJ4Ui5kvzZ
8wCaxuZjxvbv1oe4horlMFrZ+bulIuxhGBnirCvGFrB4YkxDsPyqzzVAaMIBjb80xEVzao2kJo2D
gYnQpSqk24ABiBoO+CWBe+SvPDC7KEsvdCwfYA8Ha6lO4Ebv9BpbmRhxkQYYWBRRS7upcvwT0ciT
Gw125a/etnGaRlxxnA8OmmcGoZrxVVi43qkzyw/fe/IfUC8GtSCtFmhgHEkY9zy0h5+6HytLWK9f
njXAKcIx7SfYzkNa5aIliFzZSxDsNoupvKNgaCaH0D910BqP7ZVwOEHenzfS2Mh9VC6utpFVTt3q
2Aohu/96kxVDbX7qY7UF2eL0sOe717IIDzYL1POlNCR4CLCU+rsFOP/7Zdr71m8B2GEWHd/wmb2t
03HOlog5b6+iAoMS6M/MELcHWp5l6Jzx38k8ARm3trOFaT7SGRdaodGW4foI/Kv7ujENmtOxJyRq
6ubV7Q3fHLvZA7KqAfKXVAE2tfXRb4QVZbMYbzS/V4W3l51HDPpPNov93GQEAXM5RpQYlg4j2sz+
7LlaaT5YYaLcVvWHViQ34WOfUHYljOVE+lKL49IPnO3kPXji+aJbVLopI2TfH4q80mM4UTVkdW44
+YrhHQoomoOIczCUEUgQsNc1cqE2G0j8dKH8vAQpMGrooaoBBEilGNcdZQmWO3FShJFSgAdrdnAg
h6pPaAhSvWlI0myYnt1mARG8mfpoWxIeiZB9Sce+ukrnEtuQ0imdGdoLb7jJ13g1641WBcDuzQdb
QySBObslcYwuZAYAw8IgNdgb+9qsZ7DDfgo1ivvti03MRuGTDAoe9b8MzLRfBK1vA/6z9yE5IbKr
7iCgnPYDpp9MVDLT6D42Jd4kbRjE6JeIlT4WVaAVC3sB5vyLxGKoF9CjAn06qaRHZyDIhEQCFQpU
WujAIG2PJHLhiU1cHANvVPyMvy3wSGnnorNPAITUJbdqsUsOpqHSzV6LKkrfUKiyairm+fPCaurI
NigbDLsW5a8qpcfYtCUuH4/DOgJhq1F/ogf9TZsS66bzQMzVGR8bUkIXe5vp2ZYhQ+/Dki1a2qNG
rvaHEPUfMURDSfydIcL+/WT/ctmt8SSV6XC+pjGdbdEyZCJNkJASg6u0nuKXEU0OmOMVrm1KXU3Y
tse3MLazu3SlgUMegqVAbUuibR/wmtTaEQadmuaOaZJkLy4VX6R1Yjv4xb8b6DjMDQ3Pd1UQXj8K
ZOseVBWJ9iUIpdqaGmgmw4fi/m3eVBjL+xMfq1vTDI7h93VHwsE40qA8jeQs9ZbAz68ghQXwr3n7
8bQBfKCdWqXlGcc3XbBV1rxBx/DQ1VK3eebSO9vW60jeaIlmtC76A7EugqQ6MzWY186AJPLklYzS
dVZBrNaMIxnjxrLUOUs6E7voMPnMBZzosBaB46ZtQLhK0MISIp4Ty07d9ynRrn3F6aELXoMit0g3
vTBOTP5clPFQz4YvKPr0vm1xf0ZmopnxwDuHj/K/mH/9H/MpamtUmlzeEx71uDjXedQM0/9tg2Xj
cPWyJCwgsQlK5hOCPveamDCDiIpr/U39L8uVJf/6ohW4ti/QbycEMnJaHifdCDZ6ZI5tAFht6GXt
bagojTCa8rJtPh/YAc0g64P9LdLQG3pskRhIIND36h6CPosPvE56TgVr0V/OJSh+3JfoRyTzZlOG
mPeW8SHE2rXY8QdElx4CrqxeMVqvf64K+VqtEfdY6sY061JuS+xvV7/JGyDpnlL8DX3pe7/I7yVu
hG7U3nFAfHxzGrt2Py8Rdl6BWUBYAmncqSYpgodBRf2XLCVMIkhY4YD7DYCOhOmO6NjzycMJmV/F
Sof++OhdJQxEUfJz71s5UBJqEdEcXkvF690lB2Jr/dDYsz51p5chD5lnUDcLKNa1TS7ezrruZ/X0
1w5rb8JdHFkWn6HFL1rwktpI7E5LcddlYOZdFbF5Zg84sb5IyuwiXulJqYvMeN1Tk5aRN9Q8XJXy
6SpkoPaIIvEI9bMdPpsaDcydjK3Gi8yPq+RHSrtMiy4h6r0LcmzcPzkgtRQUTaOYGFv1gylgJNrq
cd1dHDQzgeHh4kOJd8xKqdjZyuAA10UF3/29KnyPiBzBRjp6z63CoAkNP92G51ZHhrLUTBFKR83O
fFjUACBjY6FKpGM6eN+LXUlF2rjNtq7dX6bTBIhjVFTOdctg8XZn/kTmYPnmdK5gH3Z93QFN9SyH
ItO80xVK0OjfDlgULz/Fbjx/g05u3/etjw1vKMS1gHeAHk1hoBXlu5oMlI7IcKm6zF/UqKDOVhXn
/BkLrmuLaJYzJCZ5raYY0haxvDLC2El9d/ENQgdDMy8nZ+VZRmZc2oGI1alKcptFnDbryg8LfBNP
9SOAj+KfDOo4zf1fMqwySmhNVAR39akeh6QnW65sXUZ3ULtlZUzlKlXZeaTrjARTSNxgLSPS2nyv
hXXNU5SgfQu6gFXI4t9CQAfRDwQvx9omCwmXvnn27KcRapCT1e6DOvGasRoXXxPS7RNrtVFqjM67
FjJQLcvQs2VtJJbIp/WxqFJRqWoTuckfIYALkSvm+QxDDnD6gX77deY/cPs35FXuGdmlaJ50lb3l
LOJBxaWG1N/hQdmrd9HU+nf+LZh9M5Xgm2tYiBnhPWOwvVAX9ewlLJ23Sm13LyFyKaDSHTp8E8VH
NraOfrTLDTCm+WpDHNyVWJ3wN+jDpxc8JUfN52BoyDvMCXuifCa3M/cADqTU9erqBkgVb3GuzjBH
95UfSGwJUX1W0C5p4HNn4qTmBgl6H0R0I7YxciZ3MGfBePOvISR5348nca/CZSKLeESUrQXW94q6
0kDEfcN4Hqb+tp3piOonR6J3XRGWCeup1pq7QaiyVJ9cjNQxuw+3geTM/Xksy4rdULYnnHc+7Qqo
7Pptudpb0hz2C7ehIzBIl2oyq+aDjzlTuUaLtH4Cyym4N+A8hZ4FHuFX0nM8dxUJp7Uzt3UPRCcV
UplTRKOaWQ76k6CXGVDBJqTOFoeOKCFVInx7MIgRDVYIa/bIYxlfWdz69lYThEuZh8lptIYZTOeX
6dz1nTXWUQ03eZ8wFNHU5awJRFUSr5NDmFULZKFpRhivYg9fwZRA5w1ZxS8ee3hPB7WoPphheEga
74O7uqZwTJGuFRA3hR0ih26o6bOVi7cm/p5uPbf3qEAEXPrRIFNDYTxORBIrOMQSamw/dGeplaVz
hzhfC/7xgIj29Rit5sqbHAGNWSZNnub7aGuAON9G95dNQVxZ7Q4F+0IscCV/eghqynRA19/JbWvv
RaZNOUCRcL/AALXq9+dz7Q3iq317l0KYbx9KD5EE9hW+zmW4crGh3yf61vyUV+SjRS8v4meJiUrZ
1aq+IuCh/Pl7vkn8vhng9wDxsqsD2tjBYEFeRHgd4mEQZiZPrNIa6H8WklZM8F8w5w6tPn3yOGEG
17tayZQckdji2Uy1ox5kIREVhNLXTuVTDj62Hl9xMlVqsu+fWrOyD4hNUjnrw0XtmsKbccjPpJwT
uMgNYkFxa5gkpZ1FbowN6PiLoEvhkLZbZ0QR2wbQAHsUI69nmffC42K8aMUR6a8A8KXqZt4ceQSz
99LhiINR5EMeyIHUOzPfCzUIHpO3K31B/cg5Wc8hiT1Xx1m103gWgPsA5EXiKc4u+DopeCVM4T1K
z4RMDzgpryeGKCwzfOoTuPv7k4f1XhOvzNhbh2q88uft7qV6y4b22ne57GMWHuX2bBvnaid1Dll5
9OSk+Z7iOjQW3h+GwZr2G6K0nKULTZeUeC8h599qIJFbnoj3IHGirDKubR9Hr61OmNQjY2ugBVvD
mmCUMJlZ66oQXuZaIZe43fsjPyyd4c085sRcS1OYHlYmO1R47uc7h8rXaxrwP8JtG2okXUmlAiGx
lkywze8QgLIfDuKGXvo9yAwrxzoYM3cHnwIR7kpx7wAeAuzb+k9MAoJscQ094JD9N/naxEz8k2Ar
aDUeQ22/6034a7/3E8jRmvo8uq0SHXWvFHWtS3vSvSIJDmo4gOlTeGBNPwoOTjf8WrNIEHJQNLVL
IbErwrqsPjmhRcYSTRF0V22bqNDTRVKQ+xOHDeTjI6VFwNJJzr+bjT2k0T44q80bVwX0IVi9qhew
WxwBY7/mBwS3roWR1vapvzIbX8LWVJeygM4As3PdtNiXzyf8gBhg9QKRPVwWNvK+5o967BPx6Gz8
Hg+pmqdgo7Hd24nI4DhCeIoG7lQZwpWaFcUnLmT+e7BtCWBrvSjgohCAIhDTSOqVI4MsS7yij+Y8
QqED8B+0OpGcgkhMNkwAkIiIPfMO4yW/wDA6oQKFsMDYXmwtGoNe9BWOC2FbWabpKu2ckecy9mMC
g1tvuA+GrVwuk3U1nC4+VSH6XGo6cxBvB1esxgasbDYLgoZd4Q8rMwSDF8EJZ7BDsd6IVY/2Eh6b
AwlwiQIWhuHeXgfj+VIY2liX+2y61Jy3PFbsQR5BCHJmVypS21RxY1iB21ARjCNwKHg7bqLKEciI
8wyCpVT5Iqcrri0ygmLxwelANdH6Lm26PI0vsWVKdgbwZcV+OAbaZ3xigDpRFxqQfmwUhhqVh21/
Iz3YHsoct/IUEkEs+zVO/WVnBzPIbyERgooU3TOHS99d64N/rIFHixgjdYdWya4TX2Cv7bBpEnPM
k/wXb4a3awoY9FPDVRW+3nEJnwwUkc2zbkgNagQmjB6uk/+3Dl4VHShqHjFzKVYKKgKMzjeUHtIm
HzsX4iqlKFH7JsJEa4LGfMSrpabDdntF6fjjnSuMrfn/1wkWP3W36JhBZjuZD2QIbukdtJCSiY05
VQwKchXLVwVzewnYdAUOaOFaEhtsEkrKDoYxYvuF28b7Z0utbei24BXs7XMjMfXdNQzTfYcJ6Hmi
22iRU2pS/tqXXfUdR5GIcHSoBo3powE1dfkyLzlxtKWqb7AXmyrvj3iJPvmIeV2Fg/scuR9d8CyT
2q7Mi7Y0HJx6pnqkm7OOnBYFxu9OslDgzFsT1rFkTiZJZNTlDME1XZIV297OMy9P/fe9OFVoYggu
63ZR5JtH+kdkkSUjWAG96MyQWM/plxRk2Ct2RBiWKnYrFB+D4cokcUyOZx5PDVTFh0LisKEFhAs2
9vSLhjN4DkKIDLOFpIY2DFsLG1bT5pCartXINP/selFUGiypDrFuwFOd2xVSg8F8Cnl7MIHPOF2z
iavjBOXvVfwa5ob4IRvMCUKBQnsffTHxzpQfU89ob7wGxR4N3e5IO4YtQN9cIo0OKrhBtFtIFfn4
jFhSsafrvCF84a28NSiMS7IoVyA7kWN1d9jFw7iGl8dXgOmTx7yGjzlF/tS2WThr2idiiiwojJiV
GJYgd/N9nYDJJhkPcJDBfcy2ygHdad92tIgR8+qFjb8PuRjOKJCvhRxCv14EDQ0Oe19fjt0MGdpg
G53XZ7G6nYz4sIzon6f+bCsUDfGWk40WnqsKYZr1yMoiRaGUN+KfBeBI20PrGJ/VgEtRNzgw0lGH
h26lQmZfDcFXL8pzsDQpYBi3KgoSYebaYDeDhFxZx6uqs3Pjl1+JMfBOCPll5gvyPd1Z1nDt4V7H
uOZu7Ev7NQMo2oXSGilBtryVCPubmqjwbpXy0DtnHDulkeEnBO4YaI7AHAssAbCQg5r5L48bZ+dE
zovpBlbuFhLzWiITOLVq0L/h2tDWRl+nbeM8rMHfI31H6qOO4EXbjK+iZXRHTP5eyHxrt+2Dd5+W
3etIPyyh8k0BE4981LvK0KqrIrgxNlZihpH093K1WEnGz58EnXLZTHcf79rbJNUvewPtmpX1tEs6
UATQfrhdvRP9xGBDLWZFdgnBkO3AHkqa9i7aeS/FDU/74So7E/dBVUHV+KjBvxSqiDLpQ3hAVkLH
wpJeDu2ss8g9e3qGstAlDMOyVIagz+9oy6oIPnYPUXx1xzh5kLas0bxvHT6baUATJAZZkL6j9yzc
6wFeR7SCE76y1m8YstVNovVLbEIWVTjnHlCKaM8SkpsQIKv6ese/GRQAA/kY1PzNVRASGYcNMEzh
LCcToI3UUkQWPQGPzGSqYKM6T/nEFHeOiT7/JuX8IO1FhBK1cF6h1Faj19qpdHQNYoNoMhIUCJdk
eV/lpolXxSMlenTd8LdwaLry2Pzm02owd9ZkEp1LNWmVuN5i4c4C/GaV6wUm+JvWp/hvOIXb+GEh
dvrxwb0k6YTuXXZMVTDLfPFln5kLMdVArJ59Kw2oc16R8Gt6aqfYoW631jwUvPdXmz8hw8Uy+7k/
DwPAYBvyrRmV+qokoSpF8c4NOpuxfybnvBpWhhg+5DAXsr+6pGLhDIz6JsEdasIRn93WyF/wXQJE
GW2anXphjZxNEQJLaLOXIR/ewuej+eQwNGfiJ3/FQ48GApAft3dD0w9VAG82IZ1Iwko21nO9SqD3
uaWR1u5kXb7lc/aXnRCkn0udJnK1Eg3L8FURvk3vrBqtCUrxrFYvfyngmQBpN9CbQ1QLVPuuAtwZ
OZw8uhs9WGnNLIa4bLM+KGAeUb+QJfhANga4cRKPfiBtusOIbMq9TRth3OLR0vva+Z9/DkI7Tv1c
lO36YFaNstxCX6CoQNN4MaiAEGr/kKnJ770ZyW5puwhkt+RntDqodcDuPBCIP0thkkcF8C/Azcbm
9Tw9H8tOFAx+iYvwuqCVklrJCUsNeod209wy8TTiB8smwivMw4tk/jnHCHDtSByT+tF4om3F1Cw9
rn7iqNXSqT2PfydkYs5TyQujGuWvxwe0F8WHzTodMoZ34P6KkzukEEr7nkZYKMlladu2SKcuNrEi
n2HQEL5Jz1D9yCQ/yjV2zPdQFsDjiTXNsZjxjauSIMMUyuTgsvjJMhltPZ93ijcOHh1/GKJNKwPc
o5tZ1rfyOuEwfutmeOZGqi/PzWepzb3wu/RIB+meSrMEN6dpJkI/ESfKPqKCOijpBdzFk0O8p9dc
V6i+1IypyCmWKIbhtFvbZO67p6w/7XsymUgvmSJ2j5+5aS7p4pZ6eyNrQAIr0CJYLqhdmZBslYUs
Y9WFKT8UbZAQHuZu6XniGR8BNgQO/NahSRpa4a31LeySBXJInj+PIZx0ia2m5Gs9F8wzrR3vuXg9
7jZGWxGp3VLnW3ivw9CODVHRnm1WnhMosOcc5OXP8mC5mavxtQ7QDHd1Yr2E2I7tt5QqrJfZYVv8
n1S0Vimce1TUFRBds0+wX1Kjr3/wtBVndUuau7n+nY+r2HIphcXHJJ7FvACtjdiwMsHxETDziu7b
8Hk90Gq3JftAd0rJ8wHbwTCij/rVdHDiPPXTyGLDVNxgeGzXbn5fRc7ZehHwBuS4KPRwP40yrPhZ
6MOrK/+8XAis7NYdnNQlJ64Kyy8mNiFTnYEWSNiJOGkjx9cy8ScWZWbOkPwF/80yjoLGewA7HG6Z
L+oHU+uCrq+AYoxwUL89kdCTGn+2ClZM8uSJ9QHGDA72xmy01fEpbOWe2SfWKozdM/+fMz1xuAkV
tChXpg6uTmO5tFzT2ClbMNK/Yvio4xtvUkKDVsXovwfOKwbTacxb1iOOdNjQ4ToC5wiWmJSsxvC+
rV69RbTBhRx6p0yfRftskh0zZy27SfXGB42Kz+C4m1w0u+cf6z0bzPNoJOptOFcC5Lfh69jk37mL
wyk8TMEDgL6kZGsRNs3iL+egamc6dpGG91NbwyTl6ziu08n1iAF/9/CxSqQKUqovXcZ5SYr2ymA0
Myg7+rG89aJBIZZ1v3XbFVEPOhAehVdqAl9xOQ0Hg1gEGRiX2vZ2lluyonbygvIVr/w9CoFzKN7u
ClZH2uKgspVoCsNDzpFm6/vxXwBzsbW36D6RKlD90cX7kSijTcLPnZwADO2UDJj7pvmkoxp/w98L
HmcFf/HuS6c6TVT+0JO3KW8gSxsCqgfK1lxKc/1A3buInWQxed9zFJH6H4oYHSce6DAE8EFH3thd
P3v/FpDgSyQasUmsxD/oKltpkP5G0zG/+CFQ+wxgjz/LTu7eFzHVQVHl5qqzu+hB+AWgarUpbXIr
9FIpgIpSPoMkdHmytAu9UkVtvkfClwn/ASp8ph154Jld6A0dr+KDg5/Q/STdL6cDeIQAN++Zw3AT
gtU0F539CzEixBSVt49rsQLpccqBJJnQt+uS1MdmQwrdmBGpKGScrp9Ku1wx4T3Q9LxBFkZWkpNG
l3faR6yKaQgQ1yJYagzoxHy3dW5d2oe0+4+eBAMy/WGRyhqaQkdL0Q+o+GtgB2iTMOoykhRRO4Dl
At5onU2mGmIuaF5vWHhmnKrYVKq/jwRQH/uH6vWxV+ucrrorBoYP2vKk9q+Zkgw3Gk9upm1kCoqe
gZ18QfX4I8nZgGSNCP60/nQJ3rARY3SCwTlrvAIka2rSH9secivLc5ipfPWtRq0WsEzhypSxSqJ7
LzA0A0XLYidXuf94osZs2ZXYQNWHFF+lCI7BHirceVtHnTf9HfxqAQnjWXBkuhJWEZ1XoZbNe81C
Q291/KTsItJZh17qd5Bmi+vMpHVwxEiq8XpWGgHhjyRqtqNDfH1xUPE/akrP2nKm66sg2R+ur+jF
dwSD2eTN5phfboEjT8u1wAVlFB/JpQGlCdGhnHuxNI5wGXruhSDnNzkoIo3VdtCO3zqjmrdSRnrP
xFmjmb0JGXyKMz0YsGxlHT4eGFqnQz9nkh+MJoSoD8lRKVZHFlX5sfNfOmCyOqm99iq6O/CKVnOW
iUprSmCWSbNNoKHXI4FhIPFtJNs0z6K8S4fvEWfE3exfpSxBKyiMxm0cAcKiIIoBUQxBI0N4O9hc
xvoxuebrc0MVdiA4wiQk8c4kt9rDcFwEo65Uan/ztb9M/94vyMGH/3gbhHF86gLaG4mXBKF5FZ8s
V3B7mfDNVYTOiDwpFWelN2F1WUm6H9GK7kEmjsgggHOUyhjB05TCruoszfrG7eGk5uLRTgXZHi/f
npPtyqyLfiN694QmHNo6NXCbMxouK6e8MXJevMoiSd5nms2eMLQmBNTMZGCyeH/Rradtl8vktfDZ
hVXl8mWjicpbGj7cIHmLcPTXla65gRzAmv1DQhZXfX7JxVW+aGbvDqYv+QsjXmrubffdteIIj47x
gzdC7n40IhnPJRprRO/7F5anI3k08OmBuGtnbJjmmTj+Kzunyg3kZAA+MI7JP5nlvN97ecrdjh/C
nn7mflZLK/UQ8twO13klkSWtOq1GVxA1gjH3K5DDKkT45RQ6VLQis/OMMOmLnz+hTH4CP0jzFxi5
kQqNH2HtvB8YfxwVf5JtvTZ0Twl60Dtr3PiFLaVLrdBnokq+bZNWqV0/fOJdT/jLgMdbq1J+0UWh
zTlY4vb6cziLRm5WYT4fJPxHNHzrs/c2ntav9ua8lQXUhgnagMuYrenUnzAGl8b3Z2RyZ/rVTTJb
Yf0d72j3z+GL1ZScDwaYmyJ7/OCOKjz/X+eocojyFUh9/yOqK1DVwGMaBr/zNNLhNoTM4hgfahgG
HWTPOWhDXNtba82RCvOBvVvWWYDz5Tu/jMLeIMUGQRj6EESpEXpKT1bqpdeI7mXcnlLgMLF95P6c
5pJpjYKL/ByGXdc7rsHhRF3D+gpY3EyTi5mXGqV67c/V5kbCofxBgElwfWyPIk1ksX7UQ0AVqYSd
APyemu7bzW2qvyVN8eRa5U1dFBcYq/KLrnNaY4nROgfKQwF5ZuHFl68R6wtiztGmVfd4JDO+jKnh
tyGJ7KkhEMptxKx1xDwO+m5H/cpNB0vxz1GrAwM/XY1Pf6lszF0ScysQm2Qc06trDGo0rAiM8sNc
plidAD2Qh9kjMoeBSUclWcLxlJsPBfdkTSOch3Rj4SvrVEXk6tQoHb3whIt2zvxtSDA8ucit4qoL
h2RMCzDKzGQMHnLWtj/frP8V3gba7UzO6YJ/CV6LNpcM0iteoCpbrqtT32iy+ILmwsYByYrcY/0p
jGJzmgXbnGZ4OMrhRECTAe/pzH87fJjmslHcS26JkoEQPqQYPwHhvuJKbXZJq0hlHtcoDPJt3/ev
M8cEzHkD5g6anw1ohsz3UAfl96y+ickRrDdhk+bptEKunGHyRVUowaS40UGpZW8GuzwFVFiIsHEm
lyLhYB+ST5v433muXehi+VXH1hTP+IVXrUZN/v8VDZcHFqdpJuvZUjCMQYKsK1vrF0390y2lwWnu
XaPvWiWGpR98rHxXCGug7+MZ/ZFwOUCHkZdSKOc0ssaRCFFXe5YWCyLtmmuI0t0aMz7U+3Lg3R26
y1h9ALublIfJ+BWfeWND0osnlEvKG38ozaq4QcGG9ojpv7+VS2oq8Ocowmlw0z/YQ/nR3mnb2ShH
XrDJNFhS0IL7zfCq4hyv+tAgiOuPLfzUFOPP/UEtjwWahLinUndmYyP0gJx+B4+j60NNbjBBV6rn
l22O4eslHL/2/HgYaiuX84ulymXyXtl5211w8jORLWgSxbpgbjfPG70Q3DzEc/5q1cWIkI+0GH7M
2Qz1fQemYAZ1mxir4f0LtWe2w7HLLrrCrfuE2zQtRS0ivmewnoctdbu0CRmERRaDFtmR7986wkYu
iDQ+vaA8QrLPKrqLe0htHRKS5eISo+psQa6FKCRAEC4waYTwTuHuBxqowtu5UmrIHqH94uVs42zi
xns62bg++FgdJnfAkhRGCEQ5P6gUjsSE8RAvbwYySM+HnKnVZYfFZuSZngL94ak/38Qi8KWOyTXO
ymEaglNoXsmlslbU69YgrA5EZFahR9mgfnQ5pco1nF8h0BNGHAUW09IBrDtAasyPX1I07vhati38
orVCaLsK7USGysBzoab9MbSj2aIJJMIirJXT/CB+fO4+l128ipvILCqBUvOsQk8BWx+DIQpj7Asz
SbT+E8rstZl29vQwdy8ExDqoFQ7X3Hm7tQj3CecByyPC8ufK1eUzW5FoQgvtK1Z1/RbGcJVOcowZ
7QHEQOA/qnogcm7BSSiDWCkKrMV93oTC+AsKkm/zfqsYFlUjml9aBWUs+lWnOzlois0XNofAL4OJ
vKxq+LCkOyzXTWqEb4v/aJDQpb9h9ZOpxuDT4gx58ndE18mzZf/T3EYOPvj6+DwO/K38/do63Rn2
82IpjycRq4VFjY9v+Qvvv9FOFAFO4912kOvzARukQFqTfPbTliC9M6CRf6x6vvhK6K8VjmzTQiYp
pkQVqog+xoPCogIeNUkQ02faPenAMqVolRpGQIEKc0OM8ZqfC+qmWBaZP2nT70NNVoV3rxcCEq2b
xu3SCXQSlNEoeara3n/H7m8/Wb4515SmVcsFLUN7v5OirgBzfFpfLoIXp0tkaQXS6OJIMOAvCtf6
BXHhb5b+yIMUcS3JFUmEykx5A3cn983XEWvBwnHdSRajPGV7BdXB2tMPuzJchP06naiCFF8/pHR/
AoqkuN1Mm4OANchFjcqNL6CrfwB780zQZCZ+tx/1YWq/PL+/KbakawBvzkYJAG8Uq0aW0qUc+LK7
z2NrAwPvQncDL6414p3tXc3aFrhAlbXHXCvi6ECf7b0XOZqN8kpK9aAEgau44pgswxBwsi1QvMSq
TywkOU4UXePXYXbvmsIzTX25LQg77XKOuHXA1PmoVpEXrcbQzG2Eh+0eoPlv4uoSJn4Xau1nHxhQ
iCpmQE+IP5Yyr5Kj0KLOZ+ldSI7kUegOEpJ600CUheA023sDkzEJwho3AZlv9zdV1Ew4Yoi809dx
A0qfCc7NupPvW4+MxuElE6vfg6Q6oyNXvx6oX2MLEfaEWchuT9Evqt2ujBdAn0RSF1t58irK01Gd
QIU9WfNBMCmT1VoqgQAMraWplPn+IsF8+OrKg5tzBGUSA6MCliBiatQZvnNmnE8ysga2iS8VOAJd
UbvgXmJT89QiczYGG4OcezA60wCLIIQ7lnp+wgBMDGp4U1PNQmpOq7qw7dBkAWsKrA9UscQf4WeW
04WaQ2bvvf0JTGSa3CiR6vM1vdHWWE+9e6jhSfPUFwe+z1MFGiPx8lz2UqcVLc3ffQ/T+uQ8jKva
ygjzbqEvXjUOjLuE9NSczEewIAekRiRLGNGIH85k0kluphns/Fmj4Nlm4p5unYBCVii5b16B6Nn5
Ii0xwbKULdoaAzHgSv4KmmhKI4DHSAoBNmEV/5JpqhW/3+hn4bPXoN/KShvlW/26tsE9OZoubEUD
VZCYMKDz4oPy0648D371vCu3sTrCylvFR42VV0hyJCG4kf+E4fXfHpdFWVwon+KAGAfRFqs1JeCu
R6lGHWvopt07NNJ2QYiAuLD1o+fFIoiLDJKBXsyyWI4Lr9T6IspiVQnyeBuv0Nkl2aoUY82RMBC9
0haVt5tvXz3zlqRGmkvwitfIFoy1r/MkN8NwKQC4wVCDx4JUOwxTkGVLd2CVUSzy3NnFHp4/JtDT
nTc2F/839DkbrTjzgD99uCQBRiXh+DuqQui2jyko/sFbUdpxKDRI6nTRZzZILZ0YnM/EeOcE/r8+
AEJvvk51Ozm+UM0Vb/MAAv7W4H4hnNgmIcbWNH4SuuX/VPECMl8eOI22rW7QX3Zh8DJvZtAUV1WZ
rYZ8/bfAL+phpJQ1WQvr19QuNEWNJJsy/7lyp8iGSbFrH8xU/Eo1adra/oNqmit4Gl/Lq2TZeUtk
4TKaDaiZwskB020pD25qJSQtqXWnxShYpe7CEThcKLT8ZgDaDt5e1Y42DZLHOUhyhEsSifpbqDyw
9sQsNcxWn/nfLwyHSXSn0B2C4kNWzDqKZ9JRfTOMjXZm2AHMM4PJkAk8/CifKQ6bf1G7nOn1g1Qx
Y1kzpMVgPRwrT4yTqBocix4x5NTdGwe88eWmdgzJp8Mcv/XUYXz0xGfIsSH3hcZAa8PYIX5zaSsD
Tv5scIAUNgzTtTreQfQxy8fSoJNRAtEpRlUDcHRyplJQDRu16t4tPDoX+nrUOePsUVR3TrlkXuM7
xqycUGAKviMLeKqSastkfZPGThL6q7T+qeAflj4ZWpjDJOs3JJcZFlnE8r5GoZITEUO/I+jA+vuK
FUZfUyrc+owCMpt1e9T1jdDMzbM1S5vArhegT/2eMpn4krB9B05flAnA2KplxddhFUaxJEVcRFf6
QD6QT5ExYvM05ZRe0+se/nLq+RraTgpLGBMBKyAR1bODYBKEMrWRlbM0v53SXvgFTAVYBhondibb
4ZJewy4WV01b84iGTwHb6X13DG1XGlnRBH2HNMrAZ2G+DhPCSAHT5sQ5qbvsq/0Io6PRSZJ4vyUo
jFo0rlILAF4ZhO9TqPh6R40c7GlzpYr6o83A5JIvz3IqtX9yBLNV9hRYe5BgQzVDxJ8H29yWS8D6
YmQAJYVUQD2Ij95CyYRUGfsU7cZPwL+4Tsh0HhBci57i0askwhYKouCxIhbo1XHyRPesfZVUdw0x
bL/enAuZBDjVkVkLJmc3YbRoDttnjQOzmyexWRoBrKZzhWFomkbHll170rFq6fkPEeYA1GlzF1Md
+PAQbmMlfGG3c/lYU3dRyVwHM4wDkghRRLd3CuxIe89IcONRmTC4VOw6f4bK2HM8cegjdAK6+UkN
4C2VdT6Z8hkhiC580DysjTGimYaainxz5b2HN5DLM0vE9n6FCe8yLc/kfDO841Y48ZDRrn5vQTb3
GtBmvEij0vdXazBqJ2+ZtWCLDwmeMxkzR6Agybt+Rr/j5vAN8RoFPkGkhq86nMA1d+89HpoE5ffa
YDFjYXKC6kxBmrhBJG8V8duucpo4CwWUZEoqZh8VYIlY443qHcqvpJwmbY2XYOUZKlUE7JddCqU8
QfDFBuMcX9r0cNuuFBtoGHSEvcSvYusqkMlEcnA3G02VdY79dNgrEnUKtoeAQuFj53Y4EsejTMPR
JoPniZjtheKivnWnMl1XFsqaPU/MJo7aMu5KgqDnwzFTMcSOM+zjrVtcjy3nTMIwQ0eQbo6lfjkD
Mls5pbduaKsimKDuq+EHyma3Q/sI/uztCIVgTYmFtlxEhCT9yFA3riYM7Sa1sCcoTcCaHLYmGkOu
+OCAiRCoAbTqGzzLukF+02/0WOiYrmR4O0yg2AeB2gj3maM3EdQOX0Z0BYyxHQ7OzdLFjdwLoUZX
h0yR45ug3nHKuf35WbREaWS62SjHtq2HhcICxJbPabZCbJqRCuRiG0gFJZrHJOtl4NPOYNgD882+
mOCekjQoJZS7X0ScDAjZFQr8Dhi85/jfJe0TebcoIkhQnw9O/P8IazhoF9DGa4ns/JCS+OQGJOkz
qdfDAS6Vao3DwW86rKryS6OD61ZYkuU+pwbcYJu2EpuZr24NbCXQwT2tHtPD/G3+FxWRXVb15/+G
6Pg9sAMQeSzrPtaPr8PfPKybjFYjqwZ2pi4iAuMbFNrsDITfTrfW0i3tTM60Bews8R0mnjI+7Chv
8mBB9lnJ3HA6VLAJSOEF/g4+MDGA3PnIpyBEaPP0Mllu86eiwiCEByvgfCrUrQHlw6opa7C4dRMI
95Xc1n/FcKMRlVRRzlPLngEC7Eykp0l7yE1T3W76zr6oIXlAQ/hjsJBAtI0ixiYfUi6w/fPQba1L
eg6yVltGCnGSVEOvsMOfJqv8BGGDPVnepD/BfD0y3hvJnZFYX7pWFmo2Bhr5LMfSBQI9MFsxqEBx
JJJOJOHQSFCdwr0VAtiOjp7fDnqXRYVlrY2sNHjVLfscQLUmK6P0ytjXzU7sqv6SzeiN/1unWtDW
JyPTuF1EqYSN7nlQQrzRGCkRdlzXLgS+ygSkxI5X6MNFmoEfdgjSyd8fQ+LlhH+SwKDl0qDFcCKz
qFM6ko/GjaZjWjfWTOUVDDleHaf8wJj+vqs5K1zChP6nDBUyPHOD0/Ebgor+NfJXgBPH7dTQP4z6
1Ci3oZlLrYL9DsZN3aZVQWUgBZTe0BUTzSaAfHQNeL2+uzmvdJM/T8YmXI6VfNv/cG2+f5F1Weom
/9WNnkbD8p+aJSMZ4Mw6TrswHsL+UI6V53GN4iuUO6neFcvwsT59W0Zu1CheQdP5/X2IiERL/Ybh
RwqaeN2Dc7otCxBY6TSsl2NV2N0fmHOWKa1js1UjMtGtWxoXqzQXBj9jAYKrVSyhSUXabwfeTPoG
+JI3mUAeP+QZrmzcZb1YrN0SoZ/7CFH2lQqLaYs4zrrbYHN2XTCv/tIKyydvOH0jmYgFRBVsTlJs
MVKiGWHY8fPOzEGqYzCH1PkLViPUkG+dDz1Hx6eW7clIzvcTOO/ydHpiUVrUPNSKyHh05/844xBO
vLWzkXEZYTCHsqvy1bar43KoRnCfIFPUS8lLaz1eLcUQ6OdWq4OraqvnBumXabFaJ0yGlIVnNGUW
FIYBOp8rgPi5b3GzIO6CiWNbQ7ehp8jhQmv0INWieysj6YSGVbR/4Bv63nR8CHVDZsGsXT8M8Rmw
ZcadMr0UqdGpijaHN46s3yJMiKWtnnlPJdYfCEWBg9mJLT+dh9fx3VHdsm2Un22REjH4IMApr+if
uv8Qx2+aQaE/mKLuinKl164jxPki5bmKvqyQIergegT/EbEu9nRxuMW5ffRhksH/nLvweXZ0W5Up
6EcSSrIHmnoA7GcrV0oocxXlZTWADd87o1xLT+Sf87OEpQIJUb3G4kmxUYd6S1yzCeL3ZUWfDtd3
/8C1frMePoKMuIZbK1eP1uHfgJdq4OAg3B7EgQ8SwE/T42f+XXnGeKxw4e2T5olP8Aj4XLydqkjU
f3IivGyGivMdB6lxMCY74CpckK6L155PJi8O/c1+AmQnbrjW6/wJPBZP1EfeM+DrZx7sK+VGhxYo
rG+RInqJZGp3ogY5pjyimxkrv2qPy/cApbh2Zu+bojLsHYDnrkgfK+7174uCAXU4L0zqU85yEXRE
XTHjCLIPOFnlFzR0UdNpaN+xdsTAfoEDdhPGweBpdVNWVRa/ywmZsOAmaIY58HQqg4VFuuit6/Kk
bT5CC7thXaxGW4gkl1y1E0LX1NRvfUa8o1N3RukT5SdGsFHFYaEdTZd0kUwCUEfRaIH4v4xUrgpM
E4g2rcmT6l57GhtkIOfFheUPFZVQZnp29VwoJHukW9Aw/7KFTIr/4dLyLnVzRqLBziBPugcqgYh1
ieVb+t4hj2Wx2abSamPfyHJDJ4DYpvA1A7+DXGLqZjm+RjOkl14kTgEmsc076FoPJMyVkX078KAK
5KgsgUd2EvVmZPVWeD+WyyDjP3XZfGPq1T+V0r96C6qF9vNyBcP5DXN4KECW5Sp86bhYQddCg+5W
pC55UCGiKH+WfTygXSU+gnSo6oCkFBdc3BHGwZxXzSLjWmDzSFEyUbaPnyPCdtzuGcB/HBDhVDMh
Vvnx7YY2jT1tI1H9tBZDA+avS3ThqhFwLcciBbzufkKcDjMzDWHGAhD6ZDXJAtuqwMcUVKUW/WvX
hd0wI6rsoLQ+JyCXY+Z+kcb4hNEQ8N4lYtf36IuYPuqvQj6Y7Ug+qQ629TkAaOsUjrHPAvlMZA2N
uYD8+QM1Cz3fWh3HSn3uJyJ8wvKCyaWQqYrCxHK6KWxejSlOFMNSwVOvKkyCeS0twwSVAhButuZS
ah1pmcS8Pj0oqpr0NwCgeFF/jXtFNkyBIcx4i7+FaxHQa1SQSxQvVFawMHiS9MloevciT9Zpr/eR
VDEXOIYDCEuLvW6EpH2H8hHJBgmKdW1XIYrylMKcYFeYP9qBcyut4X/VRvX9ycEEuDf0KA3ChCE6
VjTScJRaAGQX+xtL72Dx3F0mRetnNJWQo5nWLDMij5Tn5UeOdQCCi1IouFwOP4A9rKd5kDJx+t5c
vYXBWE8VCzXTJ1xrOPeIFv+PdvTPmDSkOFsOLGJ1dTTRlvyr2FNNi1bgJbdoEX3NS1CwH4MbOfro
Oy+Z4ad8NznD0+X9RwvEAHJPc1gzMREa/V+sI2skhw==
`protect end_protected
