`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 70192)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aP0q4sFZj0a3bJC0chMkvhy3Re
Jt9hoQgLqVVRaxURct/2cRnyUrShRyjl68ubbSS/0XHSMfN+7dQa7ne7unS/L68SD61edFbIN8H1
WrfuQ4pXvLAuS2DiOCZCgbUV6OWrstraHt1jE0YwKNyoCIbxMwE12jQuX4aB/w6irdhHikUixRqC
oI1oDYY/SEOxhHF4sMiGWjsnpr0xR0bt3fAZuH0jUFYxH2lMHMVJCboQ1BhK1VYzFS2OS8n8/X2s
2M2i7m1W2rX9r+sEUlqvNjDiVVRXpFax6SQIpTZsp9YuJQGrHB6Om1iXL6ABIcik09bPraDbGrWe
ByvigjJy6b9H2p91dv2EIGBNstQ9MHZCNTXkQLOMDm1vA977BF+6lRN1gLAM1ZLvYcUTRDwiT7OL
pwcQBM3MsiOjP6lH80H9HEzAyxDwII6dIGTLjqG6VDI9HTE93zdkEhQC4KLh5wfrL1bNLHBCRW5P
eUOrkxIjvoJYozHg2dZu67Ms/WeuWWNU6qKRNCIfAQ+rXEqGGr9Atk1ipM74XkbJpiPVIERWx1fe
7ieyA8zJukUXKwtoeMYgWY7d8Rpc4bnZOTJU6JbfHsOos7XhscjgznPSPtStc9qEULMxTJYgmrjM
su7r9hTB2mPEH0Ovz9RHGfiIWXnppLdOvcmCe1Mmrp20XpLh+r+oQ37Xtsgkpo0ZZjFbsDYELFr2
cSvzaYofapVu2BlmiGcFhehb+3zdqrQBtmdZHGAvTYOyAEHEDFdYJCadeBv1IcTwPlPfbcPWqsz2
2wA0xZl+Nz6jnFI+VPFyfl2ib3A/C5l4EgFIvl4wJCB3rxuRyeeTUDn2xv5bbQpxD/t5zOlT45Zw
H6CCbKWC8m0C7gXTC5oUJSituburwfVGZWS9rwTfbtThLtOdejj32Vwhqfg+3Qg9R2fqbrevtOmh
yp7YHavxFC/Vr9TZrnTcv4IO+ULGBvWRyXLsKV0QADDCtx/koCRVLRc6VyF797eYs5RIN27qH8fN
YnuWiQGtmH/J1e+KbmXynsJYEAaGhpyjSJ4xtXIQQBHoWR8d0wLRjvWubkaD6SRJGdDn0MoLHjU2
oQ/PE5iIaQ2bRhmHpJK+xK2lUlKuXGB2SoMADbTrlzNgrRPJJoV/ON3+Tk9r4snBOtGHF3k+KOsb
d/VZdQSYXGFbeKNwnSicL2BsO210iXd0Yo4CHChi843TTCP2PiOqgv2EFxKZFAmyXtvUYakEbt7D
ofupBPx/gtBSwWbzHFz++T3y3e3A45eee2f38Ok4uq6oXRxsghk+LhZaU//6O3X72gZbkEBXvrM7
t5uh0YxlzpRrorRtroJ0Y60PDD635pinhaeEG4PIZTfxf7tB1YWtZvEDBtMVwvhUIH5fVHxCpYPI
BjisFTzrARXymIoaEj8x8xysLbyaZO/aZWdBabWAQufVXb5pefzDov4uLYc0j+6h19fnWeJBi0mS
IP1gw4UU55gOLWFmvDRGLcO1hWMXvXiUyCRcp4geVUIHySXI8AP12tiJJcwk0A9k0HG/3UlaPSAd
uQr/LEXA/xs/E1GFxjqKW8B/hfGyRF60yGEXLms8TZA0BoEvHEbxIg4xagbk7WORBZH17LNd+2MA
Ri8XFhjjwfCmrSG7yATqedWpa926XSakOKTpOTLJqNcnErRDyGB8IAqjRtjsRbdmrsEm4/Vug5gh
V8h/drCn2BspMY6xTYXzAbytVI647wxsUNDiFATJT0EtzYfWcXG5UZloMNeqEy462GqHcDznGa6p
Pr1siKAsccKPHQF+eH+PH0btC9wvExQKYnt0Xic2uNvRN5PnSMOJqkg8UvWYSy4W0n7jaP0fXp8k
pAdcIG7n95q8oAgGbty95dd9ymVaxGpMze5zIeML5z9TApoSGeOp3GImmKRP57U6V0L1wEnKDcSH
G4MuYiqkSgJbDrQn/slnlE2tM2DD3nt0wIP6RyBlk7b7ywmUzOxu07Q5YTs0B7GGQcKjmLQfpEAS
k6ogM0MGyYYth+SpRbotPmDGw8V+snddg11La6s7rpsnuiPX1GdfLHtKRaQI2xwceyT4BhnOIGbX
qdrGyZn3M2Et0ks/wkLfywjaqQaBYkQwXS4qaP54cBY7ioSOPMZKpnsrJeDqWJbch/pCkut+vjHV
JfBLOpVaA8ZnQbJJzUhygDaUXjDQe0pAcVQqAqMjnwiztWbUh8gFktqfwcUMQGfERtFVIxnxfRpL
sWHVXkeXRnHjrlNOO9/c2XiOju/sGdY1nojKA/wgtHlgNPgOXzKMYpA/i4a8slDuP5JcXdtJZLnH
oUtqNdTHhPSpidE4xEgzy/0raF3wr5rWag7KJwoEXsjed6HKLVGyuwV9aqtwHkIXdeIEQnTpzJhU
T6vgyZr2A4K8StXvxRh1ftMbay/kHFO+WL4kkuSi01rgH0uBxNv6M8Un50utyk1Yz+c5Rs9Nt3Wt
lQl9YmardVbIzbtcXnskFsIHDfHho/6G3bLG2eY8K3GMPq4OfRu/WsebgEetSjujp8+gVTO5lIBo
TS/sWfwQ1jDbXDkwrQtmsZhjR/taFjymJCCClkuidujpbAVq31FB0sByXM+YEDaDxa1JQ6UUVNuR
8ZKN8ZZkAZdLLUgMIlpDIcgXyp80GsPCoaHm621T0zToVjv/Q30MllxSNj2DokeakkrM5tepGo1J
pvJmlA934j7bSVunTbCth9kElkJmBwQZC7BCMxbXs0CbkGnQr7IJsYR/3EGstWwaPv/pWRzB4n1k
Hya0sgwqJzYWd1HUCzE43TzEoOg+eI9SNm1xqp0iFoUj50PAPsn0puHn7+YkuI4nrMkP7KwPnDfR
9QSWiu9S09zIihSzWjoJADMMCLUNPjve8GAO4OH/MFIX2Lz/E9B3X9y2uaJlUFyOoc7WHTyXTbIF
a4v3e7ykEaf/CDKn+sNweUk0oUzroxfxH3hSuXvJS1aKkSR3rDUaY/xBChmKmhiHumia/r/yPPDW
53/dd3r0sVUll2VN7rmNiDfNkbxNoKpjJKNRtkH7NUoQMd+cPcgHZW73xDIS0gBsAxXmeJjVcSKM
xUJ5R22ruH/sycNRPmnl6t6B5BBzhQLRcnxuhA6HAEClk7J5QotE+ZiTBzmApj5WslDT6RGi/N8y
8FYz0O255a3Izq0vDP2NcSYjIDmZ0NWH8WBYJOQQdgOSiPOyim+4S5skJILIYbiEp7KPX1QJ5Pum
oDW0CZnmLgi6ZDdIVNtb8TGSovLduI8cr+qZQIZRBndG+205Esn29F95w/dBO6gkp9bbjAfTeCgu
QgqiejfqMqrTMslXe9mf6fEq9gPpowhGxf10LQyOd8lTx+/ZT+NdMzdT2oQMfgaOatbTUPTJpaAX
I17pHVweLrno3cVux/DJv1pygNsbE6dw+cDDzgHaWUOzrNdSFk2K5aJGgQwdUqTQSKAy26Lw5UGZ
Tf8RZqkNb8xK5fWFSXc/x+/rXeNGBGT6JO8MpfgQlTUxCzIDRD3/N6Ew6Nw8ukCH0NMoRJBdrOAM
3w/XHwmv3a8CNTfT9EYj35nMWhNZuAoijifu1MF6nH7lWtF2Kfy1Ko3099RFewwznZuRBy6KbraK
8CJ/NHw22+cukO7Oo88VNuB0udlJmhkZZPu+9JV/58x/t3pj/5FEO6qgbEeqM1re5rWdT3gr60DD
PQz8D/aXFRsk8SkdJDCnu+o09I9prmeUYx/xl5uYtdjNwYJBO6dzVWTDSZe78iID9pbM+TSgsgM3
fUkCAnZKj2cvs/tjFzV9j57nQFJ7UzZnicGr550NDAQWTWTcXUTWA8yh5ZcWaSLvD6+X287ZG6Qw
q4HRTzwsq3Zx83/KwwxSqpxmH1VLu4ub5ruJuv6WGL4xD4scKlprI/RNYztbtBbJMmjzZhjYytqv
grMWx5f+A/beijGRqdlEiFP2mQu8r42L94TAVUkHFATMWa3/wbvyKb35ySFVYa2d/7QEhuFFS+Gf
7IJgD+vU1wQJfhvz5mcEkxigJcO6i3QSDWeHOdMdtJ6Q34/TyEI9KQgdTS3g+SDP4dOBPDhBAg0f
5ubM+GejwvHRZFpWVRd7Ccgd4iA8evWAJ8SEBeEip//FvXsSbv3Qy1dFkKa9etWwJVBBwkIuFH5u
T6/xmTnMhbnorFQEgDFBV2CTBDdsCIFK3la9W0rxl6Oc60JQy+vUcn3WSe7PNbO173isbtqIriiL
vtLFydYkUCh6SthdNrTQkffbP7/bVNQZg0TlYSEQYzIIUAKxDOHKRzlFXq+jzCB7rs3WPs35Elmb
W8CImi01ovP2KaVS3ASTAqM1RyI3gKwq5dZz/Z0a2q1rJAwsZOl+t/WT14hJLWIfMayThUGaby0m
GxAujRL4F7hnMoIDHbRYp/Nd3UZE97MC41fUPpmva695fBzkeeDPX8K+m3PcjyEwmuTJ7piCrSBa
P5wKX6PJlv1U+xtYqIMaED5Vuqonw9y7s0wP3jjsAicprzMEPgrn2guDL9B7QQ3tx2JPJ1RBDjUW
AZ9ornRzbjMDTLqGefbrZzNMqI++u1YzXh2c9DBMkUKdbdqWmJcuyrxlxAwO3IhJHnnXZ3aeMv5F
aPYYPODNq0xooJ2B3ftH4xAW46kAZyummaW6N8806wVdr+c1TwYDvB1e947fHT9xry5z5KOk4EtY
ex4p5IV3nY0XZyYcOJMdg5M/n5FP9IkSuUZEETu7vDdeThp6DMAAKjqcHEUFVy424y7O2jCF1CA0
LNE1DKT4x0yvl/sOCMJ4y5TkJ19d//mDz77vWfYPkWA7R50JEuqXdA/PdOlguIJL5j04znS+1kUT
xx1T5Ima/sw3F147shbeB1znMO2NQ0VANu1eLz/EGQFrJVqADVot2rBwSs6cwck1TzRvtaBOmN/a
/bIyFI4YwCbMeYMXu7x8L9ieQbBDEIa6+m8Z28IEk8Bmw2N5NVkjj4ChIwJfA8KSm93elTmfViJp
w2HVylQKzBo9iqVpGoKlaC+Kk5YERIsaxs2U2lTDVtKGtw3eET2JNTHeTwVfTWRRZU4ZiUOgrZDa
91KbVWebv/uMyHLElNfUYaJANteWzjaOEN4U9BPVc6zj4/F/Vkzp9xbo/xjw35wtanrZ8Tnq/Knt
knk22WOgMKH6laG7Ef3W8JQ2izuzj6cZBkl571t0BXIppvnk3QKpst+/0mYl/5pqB5mry1SOjNlK
+a9S8IqfVJY0Ut7356BeE2Eao6R45lOOwuZyBnziKVWdocjyOoJciuGR4t4vZPqkUmP7umF2BNo4
shH5bz7vziA4VWDSO+V7KWYsXGlyLcdTZn0QzjWhERijuZzET7PUpNQfXJRTzk454ceKFZqUI7rl
lqZ0jv4c/tnDXhR36S9U3VaYd1G3ZdfdpgP1zRSqTNoTBP8NFfgSRQ4+oYuZ+UuG5EXOkUo3Cxqf
de7eMQ/opZiv4W5a1xpg3nyQaJzbsgto9UlyVJw4mF6Ao8HkDKssFyazwM04PwQaavoPrdzJnAq2
7TnsF0CabdjAzxlo3CXqQLiNguVZr7xpMLaHp2xE5e6WVix/Meyso0qwRvORjCeAm7wFrYLegj3c
jKU8+3eXJ3gM/nTXyvkSTf7rkobWsXv50DJQG3p4dphSlL1mO6DW7pABCBtlsGq2+WZiOayAFmao
3s4NyR1m4XDm9v7tt5CU2SZSRtqDuyg2BgCJmaz36VW8lAKHid4y7BzMEtdILa7j26p2t4UoLInP
4soj5huUVoGqrUz08tkN5buG9BHB3Y0HatOOHg8tLnrtONw190kEbkAb1VlKr17DULum9o9kJA4C
fkXU6VhiUFpJXRKRj564xjldorULR0iaFXufHDyhHe+n2JYetAGS+dt70ZKYFMif+kpDWxdMRP+z
uijdwZZfMLoagdJHRkqAqQoY1iMPa/TYGZqh26uMhE9ncEFx/o2Q4JhPO2dxbmZviDS2sbvSjhYi
k3doyk5+YoDZX7afMeIv5fbEDbjjWb/aTJyCrHdJEzKVA+QNv8AnWNhwLWaRB04iezHvEf1y1FX6
NWMLd3NrffAawnoWLUy+gzMJ8sm8vV/JK/zw+66GTlheaWrvYiHrU8pThsXywoSx47tRVhDDwydh
nnhlcYbg2jQUd6/0XrJXpNOlj4YJCygSZ0Fzn/bJtXyHk4rk21KWypuVwh/6P/9me55I4JECuwHC
rEgdyD/6ABTDuEpy7pmUimyn9c05MTRoswt3Fm2ptPrSC18SA0SObb193iK7ZFG/ixDk2r7dJksw
hzHWD/wFA/WKJzRHiz+CB6VVENq24X/hQh/bMcL84OpHVIaLem0DjtoUD7MOpG3WKKaeoufFcIOp
73NY04KuRoTnkIVLeNamnUfEB8Ao/zg6W0OeO85R5nMBgosqZi5faXkYU8yXD6LtnZ+c5HSVTkpG
MtFaX4Qb8DtV8xVbXZPn70S1omQtXuFSkReVs+y0VLe7RQHaC+pQEQiX/vmilW+Vl49ow9rcPlUs
6ViWFsuJiVmWej/tMVAnieFj6as4I05aN7JwVso2OR3YJ11L/3BnkSKbyxQcCl3B3KDLGXmW0HSh
BQ9h+M7AHv4tqe9tPA3TmVGUkOs3fS7IQAtwl/D4/E0OsHBydoM0rye+lENcP0eG3vX8RRqhaJHi
I8LtcN+2vDmEfAvl1qQOLy+iTStCpoMBkiwtSbd+aLS6bB6z8YicG1hSk2kp//jac4P2ZtAzUbpc
VOzRq47gHMXZ9UMWGZgc2/A9RlBMPeBnzv/O+OAVdwypLOmXx6CTUNfroJGGLrjdS3qwC/9SgFAB
wjlK1wUv64VLAD5KSpFPF7Z4xMz/rROMFF6aSLehu4CJz8LJgzJa7mKVFG+ECh57glFWQwkEsQfi
WGnvoTU8i23n4B9G0vSfx9glxZyhck1bSWN1oTo91I0KGt6VGhsxHvJyXEDuYQ4gZ9TJ3JzFfAZ3
pOKn8Y8ulRTlD4pvP4kmL/Fa56iokAjfx1fHky0BVnr7X+xz73qQQTJJ9wdLvqraWu1ku1lbfmP/
NSYfMOyP3jD1Aw6/vPHecOERW6Wp4paaqL1Ez2TAZh3Njy1Lt6Jbkxkrq2va4wfHlqMwYnkIV8WG
/OZBS4lJIm66SVvlBztOS3WLuoCCZfyZf/7gFu3mTwRRLI4JKgwkTPZB/TmjKHt+PoSgd3UZRKPT
MO++DQxbH6C3E1W1yOuwi0W6mxIcvKRbbSbmSg0mZSacwvKhYDUZc3H4NPmZQTAeTwi7qxHqcDCs
WofxmV0rGVBVzWl+oIo89Bf8arXJ3Iq6ArF0+glxr7rvGHRbF0JlTlF/iHnlcyy8p7JpmORozg/t
wxfvSolELfQSAJCC4B1SSAzYRY/AWrL9p6XRy3M4CDT5VO6H4ssTY5jt7IWaH+p1gRuU+RAFnaKI
8IL8P2ZN/5r8UOhin3UhYqXbQlbxdUwdwjUAZCgmNbpVXngK1ZFUCZi2jPI9gBFU5r06HWIrem3u
+dQXfkDEPMGdw3BKY1FEg6WkNzSgfjHBz9e38LbPuOGtxRsr5QrKByEIaNgehpCrsUTwZRX0BYVK
HpGVypodoQYBgEQf2nPN6h9CtN7AdOo9sxct+is+D7NVw99jKZ4a4iWoTUBQCx974JjBNw7V42NB
qArTljByhAVmIuCpP0Yq+mboBjWO3aiJu8eX3MyHqrPc8F3sJXC1QGSwn8frpE0wlw4E3esbEd+s
IVD62qdoUeVNADqjj7kx+nxOTFxMfZQM4uHhmDCwgwlRtKVPK74ibtFQD0pWGvawKAC611h4YLI3
jTo6CrrDSxizKDdFf18NLf/YPHrxGwqTch3kl5r9tgxeG9/54AKOr9ho3ymDpTznFkx+5vKkH+m5
sPzrG5Tw3nPp1EVPLfTtaTOJLmK+T7CWcUBTVnB1MDa3UL1VQj/GP0uqgWhEWq0k5FnOgFuJMo9M
B5wmyLK0DJzlitCBPFouIFOPii/Ni1eUob/sxk5Ri4HzEy+rn3ghFoN5dcofsfp/QwagLD2wzZR7
X4y5wsn0WAWpU41udqI7P+jALZzMnmOFtVEOLbsiZaykaBXthApS/WNzIr/XL3s6I87v3e5bng+l
ESeHqhnt0p1GyN4V7yqbhr0vpHZhgi1V4XGw8UEwrBCLW60z/WrXjHsiqWsm2um5F9TOhoBgcBen
LQ6B16YvwojGOyfizKLJeD4hPDIerGQuJzR6UmQC9OhGZtByXFKmLn/eHoPUiwf3fDAhCnUHsu3u
b44opGN3opLyHJPdxk0XtbWFiKxGJc+OthO3IAXNCZjtdYbj8gv84zkcpsC30qEK2K6CfTF9hwA/
aM4LyCdirS8nCJf5dTUgs9QCBOiUDWJnmUx6d41YTLhzDeH0CEhygBPysiDUeeg/S3YlAdJVtjgX
C4Rzg3GEZyok6P03DinEmWIDuy2i1bz6zWZDlNNnCQ625BgC8Xmvg8lJUeZ/TehmlSIO6R1SbYM9
cAmLPl5TVKihGvbG7II1UW4KVETMxFNHHblgUJcPWPOSMkxELgfYEDPhykIM8MiHxFmp7nzV/Xp7
eOGEBMlxd/flxcTDJb4wTkA2l2Sjfpd71aroFaZt/dJAOfGFzjjW4sXSwqK13F3XtIeaAKQM5Ls2
Ynh9ZNjHl1w7S6+cJjHZ4FS948lrQe9m21G9/r0yrk+DZf964+2Bly4/R3YK3UTev2ujVNhe1D7J
bpucfjTcrWCY39AmiKB8R+vRHY+sQac44gyAX5DLABj1kcIdS9zZ7bAYlJHv8Jj3eeeaTboNKjGj
P6HtpYgda7ZH5+SpXv78aP8AP5xdbsqi46z1Cxx4TmPU8P9gEOj+JGMn8unkEwgS31/cqDM0AsJf
LLucl+czBem9KvBSWJF4tY9PJuyz1riSoDYZFAqZQ10+woqba6AfA8FrBDfzm7cWyFw65XQsYtt8
3jNtabBVKfHseT3knoeqYD2BY7mPZkbij+hBM4Mzrm8OAhsZxtMkJX9VSkFPMufQxbS+YFsgaYgz
CVVx3DVLXoWF1J8o4G1Epchb/UMU83WqjiNY6etFCim8sSX3w2ujTABIruWFahHSyck8+4+andjj
FQnC7VLBBPl4ymkiu/LrCsCI7u3yq8dF14KMPhOdlONAgR3/g2PBHax5GVeGiUoI84w3QXZA+Guf
49Z0e7aLRhKYP4EXT03wPgz9Oj0bxpv01xq+2Z8uJtWTACiyJoBomw/acWXsLortW/PgzAfWqN9c
fGRtxn6MqukmepUpWQKImndqaKMFalHBndOEGy3rVIL5jzEEXs1m8cRG9j9XrzdyOErJCjOquRCQ
7B8SISKEmKBECRzIRM5OfbK/1XjjSMjdHD/iXakRqPuF14p+g9XhTP0UIlMX0mWFKltJTsk4HWr+
xEhPmJR0P4lUNInnpEExke2tyPbA3Y0UF/In+VqLLNWztu3b+7IRQ35iqXif6j2orLC+Hjsi4GLo
PcFqXakkpv6HKva/3CS0GocEvM/LVPTya4EjCpiy1rfs9ApS7ffJiW7KxFAcUOlrKkiNoTwzOSO9
12tCB+IYlhX5ghpzKObRPUvbQkW5bDwwoxr9uub8L+exCTvUf6sy8JSmyzXp7JkbHy8hEdGTuHEM
+YhGd96JMidtLD3TD5zhqyvIl22OO78a75BkRIQ1dectPvLYYX/Jy6t1A9XjxbCC5iPefl4xfU/D
NnHHeGc3RKp3+JcI1kjPtXHS0JsR1APKN+yO21K9zXJlfgEzVs7QZQN8jb6hrtv/Vb+N/E7Cqw4Q
ht9dqp2kqlETFJCpsPhtdnz6PcKoOVL7kf9UJ7f3i5LAKaoCF1sQeYUyD4nMKH77/Av3CWSd0/zE
wBsqVwqhqvywF8Dk0kWbjYw7/Ut07zq3pab2qZgjcB9bqqZu+tS8OgwkJ0tWytux5/8LczgfcpUk
5blpsyvdKJzCObF3JZXwWH7LSrvyT7JtSAS/0tju+gUDwJHYz1OfvvyznQzKW96Uzs1SwH+hKyJb
FO96Y/lNcNHEF5/OgYm/FM/35BxtDhs2mBbSvBDzzibq8BSEKP2XBq85kOTY7wJWdu36j/nh2SxR
RZgcluclMq9kUHi1FNQGS8KFibIe43bVy4mbVOaqrAKu9Thi8i7mazVHbDU6pzWNS8VEYon0Lw/9
YkZOByWQnInpFr7JZjowksb+j1h3bL76PK6pKAZhhymtUcbKIHPa0f1uHqkXWswwO8qPmQw2rByE
kx9So5TC7JnRuZQhjTKMqN2qruJM+DYCxxd8Ca0es6fyJ+oTObhCJl4R70ktd9mL9TGxNUayv7mv
7NVvr+4DXPr2byy5w7q8YsB7UFylUsB8i1B3YfBXEgZmTe5UMpi0iM7V1u09fh63FVvduBWs1phH
r6UYz/XsCci1xpF00owUb8AvzuN5wvXm0qb4Fn28wF20cqjk9PpsXZoTnLYMekaMFqzmokSpoIM4
1uwEo4BWlYEr0qNwBe3ZCbiiIga8kLOTYaqGdXbRkfdzKzmc3WUCuJW8SUF4T936utcmnzqPPupS
XyBPLknd7kYYUbMvbkRa0YMKaVOeTXVHKhC+TItiUJaOxV5ngS9PTkKxE8FW1I0LFM7iZbieyrN0
HyBq0FWogy3qVlkmMHFo2GU+cJeHRHj1GdIHCwY40NjNBZeLJ9XT1L4G7hZYfrXaUZaa5eR2357H
ZTOF6p92MFboUSXF8YL7LlYuKLBMqm+nH/5IQV/r3rIRYqz26QUfUQ9KH99fzZ/RzUFUDJlJEvTh
hmeZpKLkGBaZkWDMA8/+FV2WSR6WzsbHTW+8ip7y/8qTHRAfM5OKXaUIluiOkbLT3a6g6UsRja1L
GTUcqB+wiG9ARiFbZpxybCDdig9vF934dJ0cf5yjYafObngN9OFaTeGa2tEEGvzTeM62nOMUuAbC
ckp0py1QmEHzMG9yUaiC5F1wdNzwsVc8o8nwYSPyEaPJpLNBONJeFN3Y8ZwJrZ6M+0RqzwK9a1sW
QDRwagcxvYzX+KM+0GtmS8sUIXZuvJk5P+PZnwX9tISlxIjg3Aak9O4TkLCHD734oYuDZK3iJHHJ
JoKOd0rZkSGLZmHQHUDFOSiOYTJ5kIfliT8aeasg4h6C7NlcP9zqRqQ92pt8iskHdCNEhYyNVX7y
Vand9HgWyXv3ku/QaN8ci6L6EYeKu+Fp5nvS92hziQW275BVF1nQJcWbRipbLUD7HrSHC/thBLgK
DgDpUT4Q0RWR/ZmdSoDrLLwsLVtQhuZpBu55g/TMpIO+Jg0R20hvXn71yi0YxdfPtzHdQpFRnGPV
n/6dMeKcWA5M7jrpS7t8U3toBvc48IHipMfo8EYrsE5Xc/B/U5AJ/1Cz2Use3COrS3T0vqw6CTt4
SHg78di2dyoW9OKejakWveUCt1eZPW5psAOi5MPTtvLdr0EMTKLeicQGlDEmeQCuODAkvDj9fA/5
SOf8SdH0jB4pWGS0IwWZNf2qU8TANNzTiuRy4l09zTdNWXuhjWeqF7OVx6zI84LtPxQuFJHBVwFz
a6XQ0PbHRywMbWMXY36cM5iaSX+ZrRGibXIVHgzNPiOxCgjSP7zRccBKntI9RokbXXECPEKrdEkF
qncESCe7M+eIkNusMHtcY/CE1PYYHmxkZJLpzRCoaZFDNPX5HpEzZ81Euk3xK0yyajAoHY5M+2pG
EWecZP46x88KwaQ6Jp2jFbIq49SdLNOiy0OHVY5lZUArPyp1B9wz8XJ6xYLcV/5mi8f39K8zn7L3
XHH9TCWzXJf1fCIXtO/C9SwZnzU9XqJ4FN4g/jQoVk+uEH4+6bQ2EcTXBK/v2TjqaCer+tX6WAP1
awxhyXk8lNGcH+LX/+rTa1f46AuYR1O1DudeM4q+9s4HmLwzUKgEAqMG3/4QYkqUKbyYWUGlGZ/V
xhgLFj2A+VQP13JCAdoEp7AnA5LujfyTqE2TVN1QmjiyY6HgTtiUmw3CEdmHsUg1CeGOCUqHraPg
RewTII8rip5cu+1nLdwTq7FkJupCoWOw2/f1zXSoGyeCfBtR7ERMR4QI3CcGzTa4jKZzlpKPPny6
goiCKKGUIKW9wdmc7mSrDndUIZylDa26H9AKVywHrZMKU4Lu3mpA6555+3DtXJrwNC/CXMz/gr2k
A+r15eIPX51/5gcj3wOqacnPNyaDGoymWJyhn3a6ei5sJ2XYkScTeWZH5vlKShJwKAjrD4yD5mIC
huE4/Ldbx5jdajWnNo/rUGw93pfkx9ZYyBpaIRBlVHPXlxspopKTT0oZD7t68fW3xnhKd27L8LcN
VsQ6IIkduDMtok5BUGupE+OLc/Vihg2ZJy5WrXQBDxKtnBoyQbA+eKAEP+cm/S0D0eNxyxdBO4+O
2+u1Odu6bMSFBQvFA8VKBQmNWQmYb33cR0YAjHfcp7LSavdqcChoTt9tOeg1lmJjTUNo+mw5kvPy
O9KnZb2ZTx8V6ZcG6YV6V444Vu1sMv2R5u7yoFnRDqaGRaJ6xDnnkpwG2CEQTch6sHJj86dp/gwu
FTGNe5VDCp5jFtBkW7Aa+Q0rVPHxczl6Xd/7rk3qoVrDrtu9areL7D67ADCSGaIOpXQeyh2yHuDh
OelKWhXZeW5Dg/tDsqv89obiBQGqrL5Mb9StFulkIiPnesBnjqSB1eb1c91zvGpl9dis1c0s8DyD
nJXFwjtGcA+uy8e7IJreTrP9V0zVxJDrB1aXBcfV88MFJegRoK7sPtGPOs51gEU3KltU/lVEYrOa
RtOHRkJKl0jhmIqiSTNq9eYyDsNODaRmewSZ/Qyu7RYnmCbJJdCiLuOyrTlwYyIxG7ValbCjsTUF
AdS9tbCJKLyME6Ttd9vc1MeZ+PQxeqNxVW/Vjyee0YX38XfApLQSwG+rUhcxd9jwNbJPZrvysj2z
GinwmYO8LiwKiS2L0V6j2goxiDj5mgsMBOraYY+ExNaOEboOjtAEwATcSsdH8dmT2xEjqrH0dH13
h3lAq0xrsi6KxsJn7pvrmLql4BWak/TKRe2dqmmpRHVKQxOBoivboHYsNCS6D4gdw1Sn864BznQT
YWkiGRZFzSe6jNP3qXPx5jZbP16H7GGE10WzKpRQ8gpdOmkXQs5jCnXhm6g0HuO8jCRJj0TkG4h+
z5+m++L/KMNrMixlFU5AxqPS6yGenAoBEkQxgIxUX5m83lWR3pGNo+Nl7N9KRM7MNviUeYb0n/uV
xcRlv49mrEWLnMp25hr6Itf2IdrZfqiIQ3lh99ByZtVTIFcyGfskTAWqW7Oli8OYizHsy3nPPOkb
KWnKts22JWyMioQDBucBP4uuNJrMHsg21vUZqm9R4QPgpeauvDyHhy1yaG+HnoiLqk71HFpGRbJ4
vB1shxIsaE7eGygOOsFGBoGMir5YL2yqBtVGRBwDJRr+9Ayxu/ePhe3uQYQvOztp1kfEG44LraJt
5M3KZiOvLvyo17GlXWzE8k6s0U+AbDxdhzNsXjax6Q8CE8PmaBYfHUbWgth5H/tTjXCzlAPNRR9G
mknUdoi/VoiVJv0M4tYPXYyBnetGmJUPsGUQDtHFpeBBBeDUCuLs0e4Vks3xXV2O9xgbU0kwTUYY
1X5jvZ7fs0tVBR/rUz8gP37lnw9BedIZOdemHuyMVw6Af7rL8FPtRMKNX3eQ5xhNI6QtJPOIE175
I750i4HnbHgiqGSu1xwxGbObtuCUz1mXwhGPy7dG0VfxQA5cAIJ95V03y3mMTHSS0nT2I8rYJFJ3
KLAvn0UAzd40MwCPFH40X5sJ+jsigDjsAcuL+M3oL72+CjOUE1kCxASClQ3RQg3EL8G1FGpHXKaq
lIszhES11mc2seGgl5K2CuSiwRe7jO/ry6xFCDMANSKifoxBD1gKl7C067DtzzCOkPhIW6GcUvQq
JUOsc8scJdLEH0SYlErVg+QlTowmeV2zDy/1OkaFV4bEl9TQWrzMeNtW3PJ/ID2NofoE5x7mcl1P
OQYH0aNVccCQ6tgLfzPuD4/ux7XRwt8nD/hNtUmR8j3AGzvLTKDLuollR8wJPQI2h6gnXg3t1RFq
j715UZV69vrgS0NwGGD0jlHCtAXviAG5oLqSQ2+du0ppArmrpjQmN1mGHWM932RJRRDMlfgQYbkT
HYnBz7hlm7zAPW6qAGzAP8Lzf1VqTXfSOtgmQjFYm8E0BB2YxOKbTckvxf1JhdhEcpZi8A1/iiRc
GFbsBlxQAvtmxBM25pmhmK2T6x/sn01UFHwKTQPnEhl/T3RdrK4GlSJfR/4SjTySFp69OxTdfyiE
JlcMD10oreE+Ex1V9jtLNQFx/g58tWuSdWIxWu6b7B0yUsu8R3WhUehP6Z3dxQ/N+jVD9GUUHOy3
FSDuEq3wVG98HARewtNzQwUHq7WLEGXq+1ZMyEmWeC1b1jQCeXj9sryVw5gEhjH2yhU8QlLkYJ0e
Dgn2C4cI51Y6Bh6BHXFmsXpObe7dC3KFL2WHVCpObR2w+EqNT/vwomj10673indmcm5+tgoydOAZ
Ix4zUk+juxXOPZeTaLTjvf8TeNtmqVQIAf+dOceEE2AMLqozSIHUG/lBYrFMI8CJ9mk+e982hDHW
lvh3lp0vpvqfMrjJZbOWutW04zXHy+xJL4lHFpeBh8KE4RH+iY+gOEPbW70/Q6Vxd455Fz3q4oU7
K0XPwi++5WOBKqtFLKiUlFEMFJsQo8TYhgQ9FHZP0B6vwa2rnPOTgIoLSH4kxZDFx2H+8bSRBUyQ
QPWUx3zcBYgJk1H8Mw5a0l28vJaj/2MoKpD1CWhaWZaEUAT7iONB64JOgw43Fj6Hdcn4yi4+TOt8
xgeRtJ6Pcbp9ESRXr8xT7HQ2aHx9GQhNrdhtt3hsDYFgyKjkI4WE2r0ccIM0+1iTz2rU59zooTC2
mTR1Z/60l2VG308WfaGFJ9SWwrd2zBHoRHJhz/fnD4kdnnWPPvCgH5Nq9RNRACT40vFgSjdBUMk9
jAn29p+AWR/JYGyPM8xrU4GqxRCxK/YNBOV4njfc8ofbx5smQNo/ZJFQJMECmlmukAk781q5ziDL
bGWektdSND7i6B6NQU3VsnTPMD9N1yocghov+xSX8mhuQj4gmbbHufv8bANlw24svhMQnXFbaFLJ
SY52x0REgBGIapsG+98StstOtPGv8PfMTatAETIBY/cKuW3CRtv7a5UWNJRWPByevLxkwMuu1yRv
LGyEjoc7/OFMMmzzIwsiTnhL06cl0dAahUrDkdtgCDWiZosW8kYFoNI0hoaUH0FF/XfCQ92u+ZiK
CkOpSNXb12sHn9RfqtAvEYTwC71s0c4So9XHPF3++8TPJj4HwTj1bT57wLvF7v6TJMVQ+TOWRV58
Ao9HnSsU7U9b+kBK0GkeA5Vhjlz/dkq98RhGWnLLXNvmZG1LNVXMgMERLqHOtNUJKxkhqMhXF5kn
QZSWkxTLCsUJtk+6Ubvx6mxY0uSrNWuoZu6iH3G1+dFtdC9P6MRzwVIIfNpAmLdETMtdrIauNF26
fFKM/SGfL9+KwKF6OMbRKmBbnP/5BgSVsCPI+ZAeybKJ609qChjhzpfB6dhqoLmVmbTO3qA8LFtm
1ufrIGcK/eUd3sO1J7e4ZQAeryNQ8wJ1Uq44WCY0vYVjMyUM0+7gI13DVFGOdMWtUKgoZVu5fA7t
62AmXPlTsafkqFVR+pFDz3h35bOwn0ZywFArTw98mKsgdMFviGJ4uC3YyJMBW2OBFGlGQ/G7o0pW
aPKJC9OqSvABusJhK8nnbchHkig8McpE6qBMrOza9/SYeWfyK/0Wizc+8C6nrNf0lJ8Gn/CYO9dr
Ydi+D6fgcVZVIszOSCATlhWEpMbwHWdyCC77c3NGmi6ewacvJ5TqURg9pSRheaJmjD2RfDrU70cW
dmf3jie1vm6HjR0zbEVx4hjLxNWfZlOaEriJRWq4M4peWji7zeZ8ZF19Ksdcwc8WbE0k5VoJ0OzV
+B5G9wJvEb45vGuF+laFajdD3r2+OhjyC7GCYweQn3IQsVGl5IxqfNThp7qoXgsiziika4ywJ5P2
ruPqDBo60p4UgUKpZSvHMFgDJNEocboGhlWjgKOn3XgWPRU8cZ6I7KYgYM1XrWA5F+hhS2tCweuG
6JssCPXoHsRs1ogVJ0gIlanBFD4fiZRDPfUHor4J83u4tPdtmcmWhDYeZQmoK4hvwnMZB3v8VqJC
2fFjmfkqyyDIA5enWLFEMYMo6WVZkBsIZG401Fy+Rmf7HesUnMUiNbEf5K9jRBBEQM/mAtO71dt8
J2cZX2bfpVkmJzGBiuq+wSieOs4iIR9CpEYXiItvPKj6VfKbT4SxQBFlYw0fCnmsJCQzsE+xRRDl
OFF8IXhyt74oQc0/KM2pKJ3Wpnq+3DZyjq2UZ8LdBd5jCjwTty4Vv1DkAQ5cnLHL/loR4icFPPrD
jo5FdD/q4yr7MQZYOVYH+63nDx1lSY8K+tUcBDfqfVh6LStT869+qYuo4+dNoLOiolH8LOapRNS0
Ks8dzScNmrx8FHzSKYq3pJwamJQS7xoo1YMaE7/5boFvPElH3UoAzxc9y97KHuH7/Vx2psz4Z9bw
J3Xq9UxQ0FkHtIYT8B88Bqw2ULLvsgXhh07AUoQbv5yYkyk1R/kJNp8cijE7v+zgzmDtiodZm4JG
x+wagHcCFuYoMsEcPQw8Lm2Z8KR+RFFV20vyBLcAJzPcZdQj44qaMJPszbvMZpEsdzcBIvPNRvNs
vdNh1/ZjKH7AlwyN6YucFP1ItgrkitnPFXwmaA7bei5qMVPsqGzU1rq2lRQmYlyIa//wUw1bXKP+
duKLR3bEfrm06pDG2wzKQ1SBMi/7BjlPbXPSx4pnUsvT+rCk5gfxlE0BoR9WgyTp/QwpTdU92upc
MPzoPKSPCogyIzq3nzDVLMCnBiL9IT7acQWm5p0fO+Py5AxZHoSCWybp6wpBdO8Vrah1Y6ffsYou
1317NNzwbEdR1g5h8k67JpjfjOJR7pRToBBThz8rDrNS7fPciznNYB3MENsfSdL2BPK4zT6zDjZ7
d3rN2Auxto83YP+zFi+94MGglj5Dg9o4bxZ3iNx8irLVJeb3uRMIAbtmjfgte49qotpenqdaSjPF
DJHsuNv0zpAuaGhbjJQN26JMecH9eASJtyO3kytS1UbnpWyTJkTl0dFWoV3GkHdNp+qpoiEyRvAI
x9oBBWZk7hcIjv+ewEbm/s9kHXHUWhucpr2W1arO38SSAYpB0NHgOJlR0JPWi6DpBa5O1pByk2oe
90HaDgX1wakdys9PhvOrNPHS4WIryBkFoHb+WTC2eMZ3tVtcqm+lJSbIh84SxsqFdhOOi5mjHvLX
gO7SXAVbRI230cn/qm61zTtnULjfyWNiepJAwkMktIRRJpvERG9jkxJ2WyqD6CUmGz4kYjpqJ/Rt
jhw5djGbIJs4thb8is3e2bxHiAKXr85ijG/MHJuqIxS1TfZ2Pp318+JmTDQAX3k1h+z164u7Vv5p
CGPDhNjL1Xgug9EBDOQ1lP5/M7sm9Qzcrelm3GCIPq/aliKwESSSG0H9mQxnnyoHin/2zG2xa+9q
Mnx4ePgOMN/C50oLnv4JHph2bass6XlD4uwlU0HllUlzkOfFWdUb/0HIlW0reg1n+WIrBTUvCSGm
IaJZeaQA9vd/CHuAhEm8CZdh3aaUFGoRpcPFRt43mIUFm9np8ZBrX/XfWPoazMSj9k942LtphYy2
gSKqqWzajDRgL+n0ehbYO6QFyujlksx91O7Atfe3YgHD5syTyJoVuNANo2tklp7BtoS6qEsZJ2Fp
R4uEb66InGQvnriVMeXvUWfIUDf23hfFNDMv7e+84MkRjcVWThEkwkKz+uFxnAtJvskf7RB/OYtB
8wr2cSQXhPAmEA/6jybIaockKwVd+ZSA6u2sISIPQY2EggJ50QwjvGYNKRj4ZXcnIo8P8BA7pSDn
9fsGoyvsdISx7S1aGvso7/cF+7EqB5mmIdV8AOf2VOypQKDqxx97iB2QEH4HRh2nphAtE85A5Wn/
wvMqN0YGpvFuBDSgtJm3Uch3w3plZhVwQ6dNejliMT2gznjV1KK9w8J3zZ6QaDg53oA30oRx5hL3
spblofp9tS0NY6eEvja3uXMahvGoVgvszHhvWTiha0Ye0zytc4s1q+FlxTvGWv8leL+IVcr+JxOt
bCFiCXDRydw3SbeGD+61eUXImFWq0XP/3HZt9QCXZS/7p3YsqpH95aPveUnLtmC0ef1QgPvbrwd+
YBqTqWmFE8XmPVdPEUPjlGq0vO+jAnNls34dsWzT5yjFf/L9Ib/P1Olj20dmlrksjwxM377g6pNM
Rxc0TyhuzDF+43iGXWmRem5MmcH0GtwkgifT+BIWCCEosgT0nNvlZWeZw6EphtcDOzvQo7MJhuAD
z3sBhfDwdHc/BySTcktXUFLK2EhV0u1B4dZkB4FSI+xA6In2h/R69Zc39DQngnjgEvqfX4wY8t9J
4UP4NIa0gCWADGAraYC7ShJbgBAZpuRSET5JqP65h1UBEFouVgLyUK9oNkZz6KZTgb8+5eZl4mQV
mzkf4UOBASJV5RVKrq0+o7Q8RTdgPxhUkJPy909fehprt8U6+U9kgsMeEec/v49c9/tD6aLXt31O
rTRytp0GfO8IEsoXRvrUuVXmC/vYPV2n7+oE8t56nXjgEVuQdk7veTI2QSubf4RzZYjan57TqqHm
mjMA1HyHvcYJDy4seeG9WvQ2CByoOJwwbuj+NXU7zkjwA29Ku0TPO1mNAGUTY0CNG+s8ISh7rft3
CQxsoNGjw1UzCxYSXTIFfNE3OBMLkavknIcb4DGPuHYWFyJ5mW9PJN+JuMSbgewqeu/8o4uxnVUh
i0zaqLMZXAHWKNxktAB7fFHz3tNd2Hb8+oz6kQmg2geqw+As+91NPTXcVSYGofnKBHMqpns+ruiF
Lcs69nfkD8l/FDbtU5HFSrxQoBSwMuDSl2KhxwfpQi1a4Ne8t9lWWINyiAGeKFc56LGnJSmOj6Di
O6VAkskG/K7THpaGI+b4vNGJQSh5sCtbplUpTOCX8Nwl+HnivPF9+I9dHqSIKh2Cbk5/l05un0+y
Xp3uGzjeY2Ta9x+FwzCdqRBF4vuTNMJ3jKRWqQE93x0aSQsnnLxV4QSR55eNH6xm3vpJ0EOFf1N/
0lybVB+29Z9+Q9dRA4s+vT/BH05tUYBaoMAACkjI1ub/5ZYC9wktxK9+e9iNhk06MwoBcsL70ou1
6D4k+x2nNKYx2AUfaS4OM3qFE1iiPZC/lceXnYKMw+7Ox8CCy2/mkTt27mHQd8EDJwNZu0FBiVN2
lABU3WU6MheplOpIK1Xrh+v6NHuoPQqXeidaOPujhqhLjdrYMRog3iunshmTLyA3BBS9mpfHLWx5
FhmhsKQ7s52EqxCeTUMNlTogMqUL/d5+r+YWOxZKBn4MFTzz+Ol0bQGzYNbOC339CtYuG8iZXKrd
W3Uk/1Q/5iQFnwFnr/WOjbrDHqm+qDPXy95btL2fPdIdekl016EFLNrVcdSsE0miQoiAe+vGeYtZ
XjgeuLqhMedHJ9RHuN5nCQJ9kk8nMKelHjE1deLMq5FjhATDAA0JZXsW4ZCdn30RJgdbiO/bjmB3
lMFj01Z7eZaDzd1dkb0Fi6B9gj2WX6ZZiA/QETfWF1cmeNBq55fDBqqCr4YkV2rvZZutvXYxCZy7
d1WtSYxbVd/2WKrvr28JNBpA7bZzvtM+tHedNTYu8ufU7K/N9bEm3xtX4nzCymkYiE9XBfE9imgA
QtPa2FXxCo/QIR3lmYledw45XAgGBa5IuqAYpytzMKeJ3ieJH2HWrCszrxsepkhH9dBYfYlCBvTx
GxpxvcG8Xarfe3dQ4Ne06KNDxfC4jlurGnjzhG3bsSv9GfJyYk0bolTOu33JXL5sHnPx3X31EV8p
Xm2gMeOJ30m1kLu0WNwWzmGG7LSVro6f9YSYxllVlOKGDyTjqzpzxsnW6SciHRblir2sDMeyBeV1
mJlcLTBEEhOmWfnZzuN9Wl8p/STyBE48GtCTIRw62ZLLbvE8G0fca0G2CRUV7g3FJzIdRLm9cOi0
+M3tdAWTLNL+ahVLzccUSV9FwGiUJ0E0D1EYqz8eAcr+qqRpTHlfBcjN+8OoQkIVUFuBpF+GCXxT
XeX2i4zc8z5qt8XA3lP2iLF1gjSRUW6p6FwwDmGUUvDJHCPj8F6k04AxEapR+tY7kxIiSVN5B60Q
Yp/2L7jBErjphAJu3L7qe5bI8VHPHZblZyh5y0NMBT+NG+dafZkyayyxv0+aGosjp6Ljz3F9oE2U
nB8dVySNjHejoxKZn3uJBS3xRK4lAIVn+p9c6UEIcBACveAYAwaEvRSsB8kxGxIw4DgpUgK23Gro
bmNFehwk4fmDXK6d/TasFpEhGNb/QLuq+HpXOV13e9VJ1rG3NhZ9ORr/H+uz0OmHFd8OWMr/RAzb
MMlWl5wA5xB+5WbZuj8yZQ7GZngiSTESHBcysTzO+ie57nZP+xpCAzM2UY40ZkANNMBYD61G6ZcT
bZTNKpGSY9IQQeEFpZIsskO0fljSxm5X7AZo3gnPrS4T8WuLdsicLzCT/MEw68fa+3NnkUYOMioH
EpAAEFhATHRpOjx2NfLscOLv8WCC240l7krhGpeEsNayn751FEihZwum1XVTE32rSEf6u09KDss3
2Hgm3BJrEzn94RTK67vkqoxKC3QuWtS7G5fksRxt9iJBYyUBh6wYgTXotTeQHNxfbrBxV4ZoWAtm
1ULk9sQW4Pb3scVzhDEDKYeCLNsLmwLExM7dYimDRcYKSkxj5ZyeZswe7X7h7AAv8CAlpZvviqs4
jtWDEPLmcSSzjd3k7d0V827PQyi5T3CshnZWF2JRVsH7W0w/lKE3M1yIncaXGAbLaVkGn5aoGYpl
1j9Cr0HssqvBXXKg5rqBnVsN5P1cnRNzei4FI2K4stUb0lEd53NBpAqlcpn/zzKw6GwQKndCd0MO
4FB0Y0lQcRv1yJkKeOXmHSTWHJSBnmpvDBcaFLfX0qWJGmkBa9I2X30wFY/vX3GS7hE1XC8n7NoP
nn4QxI+ii3r3jlM+d28/xERx2xF3jqKdU1RcOm+3CgVEZtQeWT9yPCbinBKD4f3bNo4zH/QORMoT
gGYqKqCaeM4v0xrEp2DMOdwiZB09CwVPynqndhYrHZGEhHo0LIe9u9OWbKZQ5lF6XhxbByfOKPgw
wD0cw+Wd4B7f+ba4qtnbXcsPMmea+iyRqy6K7E7aiYHgmIerYqsm5r8ZTxXTEhu7Yp554FLDPqFt
1Wqo32ovqJC84KI/VBPFzm5yTfwzxV6ODVohGzPYK65uTTEZ7lWMd3rrPy3EYzhv/IZdBCwJQzJS
4AVEuCF3N0EKXA6BqDOhJP3kPejVj9GjdmFgPqPIzn4DWKRVxLTlgFZOo6gU3jkacak9d/8Q0dn5
N6hEDVA5NVfKS/p2gwk+JnpqIh9R1LNAlTj1ouTL6L9Zp45cI+abv7i577MviQGdXOOWJSBdWV8P
+FUiBXfC9606rbHZqZmDSbM4YbMqEGuxARpEurF5zajjtts92z6/nfCzH+lN4EPYvWjZXiAiWPUz
0lmX7Lg+TA+mFaUdu+hVAkcf6uhqPdbHLpt9kATSikEE64TlzEbcUueTKNDxR/F0urkFjySzTIWu
xsQ/RTuIxEEHJpSxfoTjsrKKdVa4MCVLDpNzWeh0gJtkNmUtY96lG5zqs1u3O+MBMZ/kuZ1kwc0g
Xpq8ddviHnPHwq0eqsKP5JYj1xtSOsCJ/SmKcrCLJkLo2uRT+BPibN741D/vSEg27Z0kF+cxL8rb
iwc7cMhcolZ7HV//+4j2C+fuyXcNc1/sdsDP3m05HeiLlFgv6i1kY9l3ANPZsE6vaJRYNJpABgui
NNnS7eoAzMUfF7/s947B94z6fasIE2LssTZPDulhUuNWlCrd0ZFyXoO/APDM7IIfdglNTX/OEQA3
c1Juxt8xy71OTC0nEbEQ2xEc2qnsMVmeW82oR/pz7O73Eju7KCmT8brGPI40ZS1ldmBi8x2Yfm+X
W2edy0jZNqFF2xMpDYNSnQ2vbAbsN+RNOO5k5xoVhh+KRPquOaC76BiW/VCbvY/8FwYwSkIPMuyP
Mp+pgJkRE0o2CQUJdhDY57ac5G4O8xbCcr6Wvl0F5jyolwcRCYgcvHeSqOg/TL5EUkD2qJWA7Pb6
pCdZbFCXPzQT3cjb2lyUAY0o+ACxqPwJ4M/jD8C1h2zwvyv/MXvGs44kMkkn0H0jLBJD55tspcZE
BodtMlLuoyO+l9bcPMfUsC0FDnL+g+yP2ditCXvRGTZaX6i136UV+jXbc2RuZFqcCELP0RF1RIZo
2ku3vaV25t5L4Yxi+ia1bo23GR92zbOeLavPV+hAMrusAfGXfWkKz3AK3+PvMVlBQAduGWASbhq5
GCMAuM5jdhrqS4Oh/cCdBK3acOlgooswu1wzmTUd+gpD7sNFYoKSbizbbtvth7JxvmBpMKpZjVAp
U/mkRYePKzSx+8699wBBAw2KYDOFV2ug1pGdEoRrZZd4d1DjJuXT7GnOMtZ8oPOypdN06Vbr/BN6
3CEi4/BwLzDircqUpLOHaTlRFwL9idWP5ld4qBxXOJdqiPIXYHQummNf4R4xFcUURPouiQlRzOUm
Hs5vjIeIURum4kCHb1eH57TU59JRfx3XoaBzQJEMAzIMprhFMujoM0pyI2pxbeG5ef6nkWNEM8cy
CFd6uYluSOJk9fuE5gtojQ8mrJpw3djj1E6XLURn+lvdVeERwH88KzTUf474O5emb6HGZTRrbbsv
XL8ZSebb/6Y3yCaH0Fzi+8f1F8/G1THgDBrEKw381KLhoG+G48hqMd+d3PTaPfix1ZcAi+qY1rvX
2ioA1YFodN+kYB35yHa7rWYyihzEXUqzh1HtNk2+N3r4w1mPz+qiyZNrbxZmDvcIVEbBJOcLtRMa
ULj6YIdZnIQGt19Q/2Qp0pc0FfOiYm3GzoAd7IpCp2TGDe6sWaz+c3UCgoTrgzFhbyxV22ViQV+Z
6eKV57C+whCbHoHtoQHG8z5evnUNudKzimFbOQTQrg4KWyePHHc31Fpn+xdRHfZsNz80vGkebWtf
7EtQitMjwy7zsedGwnQQeKyUPAwQY/GsvYBEsErutEGH89Mjae8MzxlkshvsibPyz7gJFJ1YooOc
ObGSjmw7/X5zfGFP9L5GQWrnhOvCq0QQJvVINw+ypUtA2iU+1wctkCinIXw/RMz5cPFnAlUPfh2U
wxNq8Wy8Laar7WvuS1qRMIwlLNaocIVb5S0fw97zOFeVPLSwo51UP2rRZ8z+iFHfe+Hs3DGVAFsn
qOP6SBGKaT0begl6WSEg+3RpnH/DikMQSAh2QbOMNbWUQkDactag3UhZhALBN/QKDlv/T6I/ngHH
UmnIrZ9I2yYFfktf29xTPIP/P1ETt258XGD86BdPIYdrOt1IJQ5BF8ocgnAy5/DIMl1hLWNpmbfT
BoVW/b85eOHOlojfyo7zRaKJrl93PnvtYAeiM9LsOyPAO0o0gl3f3txMc4m7+1+HjLiHs48yJR8Q
Fvq6KobxBBIfLW7vNISPzrDf6s8c/O3iWowamAvoQoYB4gbLYnJzWNpAxzAV6VpwJ1ddKxOeFsMZ
iShmsIBM6eR6chXAeRiGH2GOeIv5e2c6rH1LMNrLMbuWGN92FNZDtJfSfGD2mu6PioHukXdEIZ8a
yUu9BGr/8OMBiXERpMN6WLbZj3pMquIZuvoDHX7pQCRSEsQx/5jIotpSzHNlycoS4e5x8Z3tQPFM
rmtaDPxMQea90ExJHAVD6oT11anTQuSKk7hQykiJH169fwcgVDFsS/gEiKBAxfBE1FFkrbHiWj3f
093V+dFrbJRFqLI9IYOljAfW7urEj3CpfSfNA/+VWp0aQIzWwfbhWRtdQMr/CwtTM/IjVFTWGL1Y
8E/oAf6wsQgixoCTEYQeVKrJxERCCK+9Sog9bJEV2v6bIjVPI6WXUwLyFpQm3RI4N+MR5O9Rg5Tq
5Agy+2JdX/JV284MQOFL1w7hdBjUwRZ7wfBfhBJoxwdSX21pezNbzZjk8rMtNWDnCJ0Cy1KVohHb
2h8ZmBZXbgsFQ4d7mx4N5JuHZkZqnyCCnetg5C7CZJxzh/ou/gYDTG58Y/7L5AKX0tg70kpnEIin
boHiBVaZVySYggjDI1v1m2tVyph/5+yKTmeaT+LPEEJ2gN8mrtf1v21UpKn72t7aIBhRZ0NII2Nm
40iOctXcaJwrz6kipRTXMazqA7JcKM0xXxDl9nbYX40LEBaOjMEGNyzvKLCw70bAyXSQUuSULh1Z
SDWnu9+HOfZtflB/BHr3wS+aj2FL3AITxqPnlPze7nyDk5KgB7Vn89kTrzPzBNV8ufb/euKrNJCp
6C5GUvIIl6pugzaE9onO03iWcLHlN+1P2164mft9Ph04bUSrzLSSGWZUtKiEUbXbgkrPqBvR3aki
ad+GPp46JciI2GHpCHEWv6kQGNL0zw707VmGapvod8dWY2D2WOhxQsQ3mEz0fWAmhCmhTfaVTluo
lMhXhnzILK7c8Erw3+4G2rvxVS53HPudR5mPDYwSllIUlg5aSefMwKZf8vQd1dcB+lP9cY+Uv5Vy
/8hkXxFt6bEkvYO6+woMu+ic/YIv0nimMboWMmIEXQoCAZexzWKs2PA4eivcuvB53VjpD/mqXPMZ
67lqUBlLVURcZqHCteBiGor2x3/ul//xOfXBJzEXb2Njl/Fz+0o3hjG5oM8GhVe7bHPRs4zBpSg8
2suNrwe3mfHp9dWabyjiLCgoii5H1mlWGksM0YURY7ivR9AZtkft8vPJNzLOwVmxN8IP1U0DNpIf
eV69kMWCb9wLiibTDOMkw7lKTg8TUzNrTg4T84T5hLpBr358YLDUaVZ/77c6nGp4CGeAf0tW1cFv
7m2776mUtEehdgCmUaGlMamn3E55YKKKzpQ+r3zaXY2HtrdvkQTgztZnvSJTzEMyYE1ExlJQJCXq
EQs37536crKoPTeDMgYkytMdL8IzL77W/ZuJ3NQf4cAAdTEADGtKxQKTSi50Sve0cAyZFI8tIlLa
fir53RIrRJepjp/M7gL6/ivJ/aZIuCnaX9w1kb3LlYf+U2JNiCpZjDa9n61TLCt1FarKFo0IKEmV
uCSAi0Mlye38FunlK+GO5mFHeh5xoTlqAmH7KE8iS2RafRvFNfma4+yqrqFlGeZBvH8EkoAynQ20
Qgg1Wqb6iNthJI/RgGHdMXI35XYtFPQ4R7e76SfhRK/5qJeFGChHWoOa0yvR14Mx2QXMkO362Eg6
XLxFgEtVRw6r7oVYUJwBJFhvytolC4AlXukt6QMg3XVNBrDPGGBK57MvflX4GWHC1y8Kp6jOk9YU
HP6fkUzsiCPYvFI5BayYjW4Ghp5yyQMMuhXd+GK61jercVNFI8NLVryWTQT5biUSUP8nkDlF37NI
sT82NVMSGcI23BCLdPSSrJZ3gnO9IwOULmihvOWUi3Yjd584kZx5CCQhQ/heUQryGXWfwocU2mrM
ewh8BZNyqq/WUtcEqgpQevlf884bsVqJe2aKNdvalhhRjp69QE12SiwuNMTrcl0MTuFWw5q9shtw
BEW7Hpp0HnGYL3vFDOgleRw9RfZqfKAvUVX4lV8iJqBLcBxiVhB0vLiSLrWVKCyHeL6nKC5OgKFO
j9RBN26Lj0qR6hSGcX6XXWuLkAbkoZzf9eHS8r441Xz9CQ7R6R2mqgn7V5eTV40FJQhsfmQisY6N
DhfRNGMJoIfyePurT0aTS6ScIn7BVsp1SOLSaBO2lP0957/1K2eejvZfFOUc8UcsVMt6585bmsDb
mHbYBZXB7Ulu6+XeK78EuenTWL0YyGw1DBotZQjoM4A6H2MP74gI3pW51sDV0BBuP4WZsOvsMeLN
7X+u9RpKKZUK1dnEtG21sGl5v2UPmYI6ARi6McTEm/0yDOUeHpQjrlQXDm7W0cMVdCnSkNwEvAv1
UrEFL/LN0/LICy1zrgv+QpQV5CXSnwdNAkc86//iKDW0fITG7rl++Ca/cKYsnLOGqhtmG2mhNzom
Wd9ZZNOBdHHsqr2YP7JyFYJu9OppE/CGjfZfwgv5bDZe56V10J/PEA5SG7TgYcPUNRkUvkoAWy6m
t0UzveOgi8V6ejwSawbC6FJpV6p0qICGREW/mBZha2iHWB0n/WpB5uUsOZOIOx3DDhgslyeq5PiZ
HpHLwqspncgxgX8dDSSXHDMhZhXvrE5YqiPJr1Frht50+VznJSsAdNpgUQb4T6UFqjrTOQFnpjfh
J4cvMFMs612PtFeWr5XHUjvk1ZIxyq7J/I32QgUTZgHfle5yR9UDEogjrDpRM0OrqKJGmOLPIc3w
klpdZJ0BvUpCsNwebkUvC/uq6t/HrJ8eL0r/ae6PSpXx0zLM0Q0lUXyhsjDY+AYTjUqsDvTl1fKF
/z0gW2unhdOHV7EdGAzWQh4UZmSRpq/AX0GRumZHstCGPkOCXT7lvO5GOsZiXmRux+fHIblOjMzM
kiROnzHpACy9aIU5GsTJVRDmk4hqNmoLMM3VQbNujKGgjAaemVVtwzuuH/GC/mGirxg+ruIr/JqD
s409d1sGyG6OAN7NcxLuCQrAVBDgxhF+awSqaOqztVJ/dZLQ/WIV4WKhDe1gwsBzuRhuhOZ59F7R
M3TXm7cR8AoVo47xP+4wGkV4oIlXJD0AbTgNXiKnLgKoWPinYZMULUEItukfLQ7nO7VWA6KN5PmA
G2MWhQjn/iNj515vPVX51WgzbwmSyvuJ0WT5+Yp2sqzH6WzIW/cxhzBpWB0paHggiRA972xjDfNl
Ew6jEyH5zQU8ftpG+F2E2Rp2FPgCyilbjbIX23d/dDblXR+xb+nzB4QC4GqhLY7PPuePLmKN5R0k
8Kpf2X1d3jGMPZ44uk/Y545tgNLeKX4H4IWcmljF9s6THzz/SWNZxM9zLG/RvI6VeBPdG7uOKDYq
mt+9N9nUVZL+7xys6vskdwcKctoWnc7uAZNG7gKfYsV42cjQNlThJQ/Oy8479YeG7gUzPv8k+OuS
Re0ztS8N+/Zk2pWSefdqgtATR5bVXmUcUoC12moqQtUYV3hnlx6D0j51kFjC/1yfgAEodCS+3TN3
72ELI5ImVL6U0Wtvhlq9+FXpiIYo8aXgvdBfS7n/ZJxU7V54c0+u7h1ujSgI5Jes8oU6PB6m/1R+
2lfMSnwz6T2lcinDyNgO3BBnAETiXBX+b3t/1BD5JT59INl3UlwqqBUpkVOtCsJunB6bKsCduKvP
2PlO1fuG7+xzgR6IudOOqyi4Q2c83HfUnrhQPFcBTlUbsbNAf4PcUfhhp0lobB5I95jdGnRBqaLu
NQZDoTI0zjEPVSHLmp1okrYrbJ9/mjqX6n06YXhYx8/MVkahzYQefapyPH4vYpiKi3Kp9Uo8YAP3
OVgBImCN4YwHyTQSuIycDTK7bzal/GOoL6y4ujVQ9b92zf0O9vuom3RQZUKZiuYvm2YbiSKIJ3FS
SslbBXKnAcNZ8aR9qsPhGI0gakyj+Pj6j/2Jz+sgtYKl5301ZvIU4PXke/hs0W3T6OYewFr03Q3K
ltUw5Fc8KyckH56AyJvgtHgyUZhOL+PkcxPNPZenSoaOtpyvhosuz8IfSiHri8GZe/ItC32UmP2r
c19jHE/zWwKVeLihjBKanul8En/lQa9+qtC72KlfyG55azZCeHVM/MJASc+GTy7ypXDtt1LmpHnK
YYORzyXrn3YeMwAwbuHlmK865aMPbfiKjz9wXZbys4IP+rDsnk9TAhqV8+OXlmggFpnTmJjfHvjD
qb3lYXp0c3yXwxhbMIUCllMW5008p01UZlOjU8yfwaILItuOhrnH5AdCskrmalSceGBFOj+KXNqm
D3wA+Qpi4vqSxfTZR1/HeEyi9+AV8i8CbdoIb4Kry9zfBpLsk1YqBHH773HMwIqLeshQVLIzCf0Y
+KlqoSrp7TXaNKf0K65/Bt4/gYWJB+H93n4Ka5nIXfdgn8zewhBcvlsnM74b8vvturxanImVdDbd
YxoW9T7zsTb+dn9wvlp5+JKFwtL4k4d1DuZTRUtu84dCoDkhgFd7PismInPN3YRGY6HSbbZ2R3NF
764Dg09e4EyHLXSLpNKQPAOj+rY+JMBqXog+02lu4svChKCyizgPy+XAJE5ZQT0TJ/tC1Ok3Vr3b
GwKAhzwSIDRuR/63nI6UizTvLuFes/voXzl4KtoanG4BODQ1BbN9mo5l6n3aDtLHlfnoacQhOnhS
G2bDN6iqbXtc2UBIUdzrKz9TubRvmqenNgoNlza8J6ks/bdCA19AAioiZRSGEgPUWsHb+0V73g4s
wI14NKigxTlK2jCT2a495t+OHSdJ1pOD8H04JMgFx+PTdS8ZyeBSbZh4i7XPMu+WrtyiwWZCJHO6
PHziCQ1E3SzF5Zx0y1ZdDWS/yeDcE5C/rscnZUdnPRrh+OWWnsecOIL8lt41Ddkweu+Oc/B82u9V
jP+7focEfPDmSzwiZzTpAksGOoIjysKdVd12+hhiB4neevNIwm7jBybpE1nHxhNRGPfubnViByae
RuN/jk0gU6TZIgQZO/3wA3WuKMGExDmA9q/1BxyJHzFoHWpQyJapNOXCI2jEaNg2QR9ph2wGwHV7
GnlnMr7Awu+g410tGyaUC11fKiQQTnaIZTnishHaat2T+LGECHSJeirIzvRrIzOh0/x4y0RBKnha
7QFOb3wPCecfemWP2pyTEOV/frSdw0Y0F3BI7BXF9DbKwh16Hs0IJqD+6DN0vskNiPammGjsd/oe
hgg7q/Q8Nxj7hA18F7IfpL5LIbPAgn2Fk0yzI8FYQQTUCAZ8gsRrORqN/1nPdcaMbgNkuNLs72uW
Ef9zfBr7z2q26/DG1QIq9TSp9+FBWfLMaWBpH4q1koFsjY7TzNb2wOyvOvfMhbz6PeIzCEWWPMqC
SQ1azwfdO4LrgwS8eZ2+4sVKkMMy9ixceYIn1ujYqhNjGmHWIp3/tRDVZEsh97HaaYIa08U/TmRM
WOfnbE5KbCxMIeLA+3ObbWVUAlnc9Y8LZlf+qHyjWtWnfi92lnBNZUE5gc1zviUr47jwi6u7Kk8A
o5JbGr9+ttJ5wlpQ60HD+wQd3O1nwBh+XkFhM0HetZ8wG7QMyoD6LVNIM6z7r7DqRW/ykZffA9WK
cDZS0Wlxb4R4n+Ot2Enx9GaahRIHJKijWHL2ewSv8JrWvo9W/VFqdirtFhhqpgUY0zZZeeOiRB1g
FrpUp9ty41EHhObIcobMWwXv/VHLBIaVQTLiYKSAsz1DEW0UQiq8WxeE5PXhUPMkyi4U4qhKtgE2
RXXRNynM3u38H56FWo7c/elPHREaveUpZ6DwfNhL0W2wPJ1QzR7U6LzW6kCj/D+docNFtP2lD4Tb
Y9kcZ4yAqr3UFvmnnVYhX7ot/438Wufj3UVy3jORGnRIqJ/wz4HT7JokdWqHP9TJobXwOINKByUS
QxAwfMYfuMmhbZ6QfyPnWTNFKtkgjdSXMvAUaVQYcusxIYxFmI1pKsgaHwvxY5u3gwKiyaVtpVgO
+1cUVRAkLEQGE3bGZOakSzrdCLX1950MH4LX6CS+aNpfuuJmM0PKKcfSWJ7d9MOVK6vSjOzstQYY
J1KUTu5PTvZG1ptKtMVPV4cW5la1KtauKWRXI4DNjGltJgb0HbBlIInPvXQunukvL8ThAMnZC3sS
cBg1P8euPvCvNC00ztzbbofxx9cyLcyiaVjXyV3RazGXy/D7NNGesNTriZo2hUBWc5armsUaz9Rv
mLsrPGI1BUp4nAWSCB9U1MlT7+19LmWUkBCKsj8pawJv/Gdz/eS+WxZXTllyx0+b+iqmsnmeerDO
afKcaEhgGa7KGiQcl/G+RAN9gycmixMMR+h1XteP28qzIDF3qvyCUgeh3B5VihnhFvGz7uP8Doaq
z8XJ6VBkgFtd6Jvwg+/XvwJuqEVAVb4s/7iAA2m4JOHZGYwfJS70N3xU2cVTVygOm77eCdz9jjmS
EPjYVqbzByoLREXpdGlLCvHL3zR1Tu7ZFYPixMoO7UyNqLrgeIc9/7cVPhwiQSSLLd+qN4iBm32T
j4EznJiIJM9DidMBiKBd/lAHBPNvm5cUazY16aL1yQsYQTqjmUNW6a/xowMZ2iieO6u3P7p+y57M
Zim5IbqJFnj6b5bHEK1ylOTxuClKB21UgkAm/Aaj/CcWZKAMgEzBKceouP2JAG+tDNP4ed7FfsD/
FRLuzpTcx2eCZA3Oo2GcMk2n0k9y8qDX5ouRsLYBILkutEwYqC990GFDCLOKLJwVblEaE2aEZiZ3
AP+VPojCCm2auQu5t0tjQkR0ue/YoDbfwjylXtZkvl8EDN/cJXVBgr3CHGHdvdE0bidcP0GMsk17
Nb8rkZrO/zGxAaJQGFCD1M84lKBWeTIOJcglNzMGGu7vUjW5tl3KZDySUAH08tlsbFjHB5MPZ+4E
+JMVOAe4y/Jh+OzuDCVK2rPwgw7bjsgKZCVRLFlT36jWKhwVsKZoh0LS5HpxjCzjZfrZV2shg1sh
9e7KrcC0S6rgpP+3cZTdyrEYY5WUh7DEC5JIpDg26e7IBg1yWFpZvwjqTf3Tl5AaaJB8Xsrl7API
5fULDz9fyyFGq2Z+pg817chvavCHoX/0HEaWkwgsjLs9HkQeUD0+Mt2KDpWUTaGxI0yrj8xjYXmn
DdYv7tnJgJvJ3FxI+N2FSl5ZynQDkDO6r7aKEWdX4MqdNn/pmdnZm7m4l2X9mVJXEXSgXa5z7AJD
RTC/O9naqW62a/Z4n3U94dXnbdaozAxrnWznq9hGJcFcuiCmD6vhG7Rch566+4dqPWJzW89iN8lk
JbCDuy3o23e9UdT9WCIZ8Ica/L/u7MJpEsq2nGFtQeR6AfTz0e5IaFtI1v5ls4H+tvkPKy29x6M9
y2RN7LnjAVjxQPDmjMWKCWTQHBmoclnwitSadwTh/q88lny1iDBcaErnC2Lcm0Tn9mOo9mXYWnEJ
K8sE8RcUViF7Zu5qRcHaO1X2kDZeqBTR4Jx2nBYab9xoQxdrybrGSgtAmFBnxD99KFDdM4EtO2oF
EardQoPyn33af+SH7AuhQP4nxZncOT1Ko83E1Ld/SNlAmeWapKcglxuDgWhiTJOgazEr5+vWif4j
RkWoW8pLLgMd/beWFM2D7WqNg6i1aCFscvMt37rox5THKIrmt4C/UoSv0+Dga1d+oYY7Z+sq4mzM
/jw1OEeSem62KCSPTFOu5gDzqtQE/z6+9Kwf53ohNHgUC2f02COm2wS6680WMrR4Js0rjLBz1+Yy
v/TGIYHISwfsRkuZavVpTqcOMWDsvl0zUYjgehXl+MLbgiGMLw7QfXAN85V5+Dnz1ZICuRmSTO/i
65jGurtohdxN4C9RNe5iI9KLdXxKj2+YHFsxFMOpxVDqpc/oevSDobTa5vPT5/hgfMDqQQTlM1Oh
0hOrgHaXLtp+bZI5y4MTjt5JRWBul9M7AyjD4UV6t+EQteYwIckYBpvwrrK3OFznbORq2lRNTpWP
Od2eBhKSXtDEcVoIttKYXOHtFQaJmFY0pYLDCd0SSdi0bl+pJYPYm7n5e9R6le8qPxxxPVJvozPe
sl/86EXQndu4TxZqa0iCT1XexcsJNfcQeaU1zxxGvyqNFb89Xy3Hc0Awi1Iwa4EE5Afh8axI80e3
ivj5rigyeF8nLbeeDgV14eN9l3CBiqz5EZOtHqb3EVIXIxcGT8n7MFJCC6ce1VEDm2KqmuuKWBY/
ASsY9G5NjgyBLqOKrmKGIOcqxpPlpxh6ASEge5Ym90Q5vWlYurbnrcbpeUJx//izEtOhL5YkfgcB
KQoWQJEm2Cdqp5kZCBYKd9lfcgMzx/R+ON/Jw31Q/fu592ghiT0wPtHVKeZ5FrqLPNL4/XKgzQzq
wS3z6u9ztXLNpOvLnm/aTYuOwT+vgqE64iEORlSpkBL4+iweda9J5Rqb3QLneGvJy2zFt25SrbIC
i05j3Dn+8a/Y6ANwTEgYj7ujSr1Aml6cROiQdvv5PeP87A84lsC1VJsU839tRERN/r59NfWTatqv
g1/1cFjJHKzoCw2FG16KHwDxVJxMGcONj4oZqeHxNB+1o7KdOEUEcklELoWRpG8G9ElHiHZRFFpI
6SFw58FMoierVwAbORZ7kD6s9F0gK2ULeCk4M3aQx2SFnVxcIfQWB1HrOhThIee7QGS2nqxi+uJC
1yEtvGaykgQSngv7MAfpC+c0SXkZ0yDHbTkfpWtBRVCC/BnzsZnH7VENSIKL0ti1Fnilk5vuaahz
w8HQ6QFyRTkverh15rsiANdv+vDZZAZg64dsVzNvr1UJN3PNA5sJ7iX1lubCvGB9WS62exmasTSL
tplqmC8K+GxPrwbTI4a0U7bTLVtk6mF6xW8RmaLnHajYdg0f0i0JqoTNs6ksy5L8UHVGwO9rMvqq
DhsGGVQMbi1qJ1ohQFMjc7wmf+Kd/Y5W7CNCr49Ork5GKfDlRwHznWs6QlonHF+iMw6JrIgrCBNt
MB/IEsF6Emex6qVwmOmaARV09RHODVSDXhKdl3XW8Y9NaT4nLZkg9iS5Us0uSQNq38M6HkRkZKBC
wDiuou1DaYeMSgU8nUvgc10qA0C5m4VPudjiX7+B3PotwHGYyZZOOJqmvQHar/gmcs7v48bh++9i
JcodJCpuSsglT+AWFmK4Q83DS5zIOWm9/nT4u65xzRuPlMjWNGGAWYhVFv30o1fk639N5i3WXrle
BfjYx8OHjR5LOGTRmwOy7V0hlCF6XwZQnCAT/Ne6xzwh7F0+YBR1L4iD/41VzCuUny/NxnpCT6Pb
QW83IBh+2ODM4ezSBfGuobZGTHmDmiCQQnJTp7kHqtNfXrlUv4cvWSOEJoaemZkaNTTxYieJ4g61
HaDYAkgPBBNgo/8mzJwROi0hQ7G914b/N5HNkU1RTP5CvR2iPPXGUdwGQ2zzveUmyloSII3Ysuic
zC/zUQdO/I2PkL0Pewe5RE1PFu6UcOxQYQlNu3qZwEJUevvpyqGYMYI0GXu7zQ3HkmNWJoe/06Dv
u9dXCKJ/UY9zV47NJwxlxIobXz9o5ksir0vVMLKvZbHtkYXqEImhWf2q3YL4HnU/jxetluPbf89c
V8WMrq1uiQTC+bytCj/1kKlHq2b9EbTxAqaFdNJhYh4NOQSw5f5/Gz9L1P7Fv7XHOHkSSUnA81mn
pLbafL74rlcQaN0zL+WSWZ8Me7uXQyxNK+RAIWiAhz5rcUbNbTdYgsrMUHjmYitR1vqeYQTrN0Jb
c5QXNdknrXsyYelh0h2dlvzhaimQBXn2iN7aeJC4UVoNNpPzZT8XHXs7T69GWhAUY3LxCLbqGBku
EN0ap1wFZoPyvH3raWduzzQE+o/sMlRG8o23DTYYejByYrt+twYOvySE1MAMv6GjIH9833Zm0PGY
FHvOFoY7n3WoMw7WMJ3it/unCdCh7L+i+HTyD/4Fp5ITUKml41RedayCxp/W3hobwBHaMpknNFj7
3WsW61IPwUxwSQvrBHbYSogNyh05n2Yc9L6c4MLaBUuzWxLQB8WB+Q31HJdg81ruBqfDm8vg2Jhd
b9s4HInzvgdoyGAIRt8s4t+j73SSq4uwm0ebKX1tclMiSbnGBFOFaAp9gw4sPG2FHp2AdTaonowC
yVQ/ScVzkdM/0ccKywp5K/azCSfN8LkRYwjd1OMqKnOyy3dmLxNGlSoWf+CrH3ylslA3ENKDzFrk
es1rKVBfQYyupNwL6cCLXy6jdS96Iy+fVHxKddOxPrKZanfnFoexmTez/VpgnRh9BHw2MPXT3yUL
caKFHbpGOx0sG3zHFW/6uQtOmpL2OyklhBwnYQC/y1D49Mpypa3tjBrJBohuMMp3HKO7+jlk4q4Z
SVCX5bEjBYs7n6qfY8V/vdsxxc2uYKxFept1EKw9IljrbfEuvXog+ALxnh/ZVXUWxK+707tMF3/C
mwci/Z13Z/o+wmBWAk6FEX2pNcBGpz+g3+RlM10iClB0gc7bbAXU1FbiK0qFqIy2Ghtnu0haX5Fj
3cmjavnq79Ps7kgICUMHBRiFENboa/iDaMP1ob8GofEa/bZfSiaTuVDoEDB9KyP/xz8aNCEvQ/OT
I/wjyH6bezRAGcg4WHPv+l3R4Lz65/Qpu+VNrrlaccJ39mDe5e75ErT053eK9Y7evo3SQIpMO2rb
EY1wxCo02ror5ewZOMZZLqL6QA4AufN8OtWXYqzFPji204cPmneoMgjvWlVNj/qdwyWklooWJI5Z
RP/GnB+2FOP+B+OesT3Qz3l7ryn7Orm7m2bSlT3OKNWIxr1pUsryWu24pJ7C7C4fjrH5R9hDwhz5
SIDL9ezehKRo9tWfO8VGraEWTrPbDd6YhsHVb5hHyh37bJg7QZHRCUOhFx/kDXB6MQnReAeZ/k9Y
0nwi7DMh74QHgKQHr+ikEqgYHywSPGyZk7TsKJzHBajsmbc0RxLuZunugiSxoL1AhQKfJI6o6tGQ
xaZml7ZMf1MhjcOLu29dEq8VmxtWqJkXW4CfrKJH31hKNR5LBOGaJfkiPh/wpwn6LjmRUG/pdM2B
VbUap8HvH6zAkyj3fTv3sgey/6jeWiITgMs0NGmYM8sGy2FEzy5Ad4EpbMWtKlwpwwn7c5j/2Rmm
I2aoJ1y2LbdP2nap8bfwZuIPqSUvXymifgKe0YFp8FvaNTBkVjFWq6b4Ll5oD2LChO/1r19ZbGbn
2xeHbbUtqg5tKmgsAsCgr8PzK5YyWwtyH4jiSXe2uzUk3gFYJTDSf6u4l6yX3PvPOKDAr5ej916+
5liq6b+2EUuglYINWC3Rh7m3NtoHWFSVIHl9UXBi9mcp6dK7xx/ma5tIIoqzLNh76Dzglc72isSH
Jnyz9EkCuUSX9FL76IuLGXob1tU5lUdEUvz/qUmPSj38PTDJy07XKddiWpdw1Z4vlBzIHrxFJNl/
mLzcPne7GUUb4dgV8lULtVIxUehRkFqzTenDrUzwAjrb+VUaT2e3aGOh0QPvhfRjk0wSoS5PIcHx
d72odp8WK4+QsTTE7g/304comXJuilMGef7xjN2sJdkcmXhh9gv4GA9hu38BQnqVlYKbJIn7HS5T
6tH1GeAmHUOgMUmwQepV+h2pVUgzg0sBsJT0wGUnLAA9++mF5qM4dGTbSl+K9w8F8rfl1EQSaxkE
45hL633FsJvUj+M7jIkZhuW/Wa3V0Drw0lOZpX+b8qPNr2o5niaAHkphVpPHR8O2XizJ3CXNE8hO
GS2E2vgWfDf2D0yFvC4tOuwyE5Xxd2ELhLMhXrWF4naEaW0/Hke2pR3Rq8gchOP8suPPEJYbUJX7
GM45dU3QYp5MQD2pv9ShpWNt7ZbXG8NgRElDhHlCu/5mSQ4Fp9zONd4DT0pmSEIsDL2wfh/w3xlF
4vAyYDmSD8LploJ/fLPiGPHvPx0ssfsp14Wl3TH4ZHL3lrTzCcUxkzaEYv0lAGfqQFVVj94899G0
zjkN3hBziGBhDBtIokiVDUI1YqkQHaP5uSWoiya0tdjWNdyceWdz6fJKtYQjAPvvG7WcLexuJVLg
OTunw9bNxm+X0ud6xLFnxR/as/u+RQZTLKDtB7TBAqTG9BE8K1XQ3pOAsrCxfasxulJsbTpDlMBt
do3f/tuHgn1MBMAiSGqAv/26remXb9xdcxivBok5Hl6hxJVfUtRIHtdYpDtOdJDIgJoOu+U8QP+p
ptXXn6vT/VPsWJduzJNOmqfFOrITgpeBYd37yW5r6sERRrFqD0zcmXJX8UUJLuVKXKHgLrzJHobV
RUqI8f0XJlS2YOYHo9+ustjQTut1fKr4ktVPO4V0C3PJ8yiCT2n44bzloRpFkGj4ICBk/okSsc2T
uC9jRB7rhzr52X4TIFZqfJ2zAISCmkz2KROAK+PYPCy29Ig2pI8kDJ9DCT8nE0ZnwF+Had1JDe+c
LZlF5DYpxjDVedrQN3COzgxU7r/QQa6g3PRTFwdUMy4/FkZnQ8rDztoFRdh1vNGpGVcU66bCKubp
XWF1LjqMnO9YqRlGpFl+F3PnyW6tgPYefKbhqbsK9Opc0/7k2W9qQUe/bLUeDpDcMOBzNNnoGrTY
HkSfIvaVA9dRfHkKoOV24hx0jWRymUhNmlcjJAzAGqp9zT1XJ52k/ayqiRCQvIYRJusFHpOIna1X
U8E2HQzoN/+S/aVc/jBjMdsHRMKJhW+QJpah+cob5t1BW6+eRnwX96HAaqM0tCkq4GxBIRIeXF1+
dHJH1gWgJb5mdlevMWGKKcP+TRYhTYbxWb7PI7Wd7gpv3+7QdJktd1M2TkLeCErX/JPoN7/nmPtg
PGF8nYnWcJC3ZMbTsqHqsbrqqIKpTTGfDnZJOGL9nSXhDk2BiQbwcwGnbnWA15Jejj1pg8pmsmSE
pl/wsiVfLTlFhXYGHPbEDgYx+jECO8HI60ZJoQLpQPnlQG3tcV+EJGMMx+s9EyoLcL0MHN+QOuCC
BlnWSfQDNOsjRvab571ohoJYardzZAMpCepPWQeUMNE4bQc3zXUp4/WJzqKYEcj93sbS15ylHNig
2BkQ8lESPATuTmnhqYzZsTVgUX1EduRU0/S2vCTClIn0o0ZmuxMM+i4c9aUHbhDhVlydZ7ud9jg5
qpUJqZ7utS1h0wmVO6XGNDLWhw0x6m39upp7CCuZd1wD69m01TkExdF0GqsLNhq/YphirKTbPqwm
GQy1Am7Uf82EbEJJKwiBBrVMdxaCzGMuJTOygqmJauYiN2Q3Gvkk8dVGLQv+OLOQGM+OGQ2ZRwSD
KnWvDew+0qLivA84KAgVB9THS5DCEtHs9c5V8l8RnrqG4f18DxqtAAwNiHAJik9jINPpbz4173uz
AmqEqlPnHmEbtN4gXZNFLKu47Swa8RKfhkGOcQW4ODC7F9gNnSbW2thdZDgjHdtrqqEPCL3XNqUy
3Z36pGKgFPjJz1QCMDJEKqR0jzgiiYYtzIfUh1CcKoiNWK49xvihMe8nK6CIeUmaA7SBX/SyvruK
2XvdkwpwR5weQMEgg5POHwy8XXfWWKGqQINXFsWutW6tg5XvetCQb/45pwnuvDTpzEffJfADI4Ck
rI1DKH3lu+G53+lO6AG1/aQPVlreI1t9SjmcDMPOz4wjuhs+krew7dcZcVwOkl+v8wR2oCEEyM+F
FiDpS7f9dcqJ1hxBuBs6CKG56sOoGg+D2/c4xvFcaq+kGkEy/XvakazB1/I9De01aSRnJBaCqO4H
nOCumZrJ6aUhWm5rRI6keq1nFxTDZ4bFzBgT6aymvRr59pnrljhx9/pKjHJNq5DcslXLBEyiq7Rj
Lijly7Fp9Y14tlQmT+ipOqViixJ6W/pXmD473dZY4gl3RBXJTXFeJ/3PRBBo+mIuMpaf2OcNFuFR
/sjVpTlvwEJxIT6QjliXxcVikaV5lStb85x2ZCUXe08J0hrkpeydHyDfRM2Nhls+HgKPrw0E9DFf
674iKdN9AiMMt97qO6LWO8vnFL2Jh4w09LU99Qq29hXvseypHDhTYoNG9PjOmCIc2xjwHtipk2k2
6uCt8ixPUti2Y+fRND6iI8Oe3VOVgC8KD946hxm2ENsR2CJKvHB/xWywyiMhHdfjFrFqhY1zIDim
/dPvEE5PmMY5O/sSmt26VwPQB7YjuFQsiyTb5zp0nJc4cYCaifWbPVSXtjpqUm0gGofXMHYnJx93
4eXCzgQ86kiOoqo+z9I0jcG7ZH7e8NCoPjYMcaG5PSrIPwFqPmatzPS4tBlqffjvCxhvf1jFHyu1
Ue6xZ8IN412TfqxAxyqMLHVIbYtuC98ioewglnyhbuYeq5t+khNH7M7i4F/OrLdq7RFb2oPYW4lG
in/iM4zKJjVrd6MsEffE/dqRpSj2vEJ4FI5yxyz1xJJA/IkHCzs0iaz/pvZPraupzWzRyYyRjyyc
Qcu/K2Cxa5XoQvuXqfJl7qutq0qV02HeH/9aXc3KcbXIAZm3+N/vWyG86EqVmHfE7yRRL1D+YZli
xgoGBVyg0lyGyi7NVi5vJDxh84jyh4+xXWOy8n2dx/ohSWJq3Xp0IuaCq3spiIbfKLEKQ8UqF0En
jzPwCuLd4jGYQUV6qH899EqcAwS8cZL7b8auumQ+BxGOLfAmCmr5A3CvuWVL2+ByP0xYs4hZGr6z
/HU7+MBs5FFm2h+vDVRW8wvilQnbAhUBQ6WMPNNKWzezxtJWeDaRk3PAXbprKy/XwwxwrlmjbXpZ
rOe+EO6Nb70WbBrG/Sn9PApkSkA53YlkrFys+Iyq03rp1rVyCw61FFUzCZtMBf2+zNBw+P0B3ldy
1nxHleYDXpSLHsExEAXsOIXFGFycNA5R/z5wLu/ZnPxoPCGDXzll9pnbo5s5egx6O9C1NOjL35Ig
VSnhcNduf9nA4GUCFovg9Tp2AbFW9UWnsdXAEKi81MEFH3rjpPiuKcJdBb78fMkcq9H+ZnAzZMrP
vP0wu9sQzcY3JGjNHSZQF++cwQFfVu+WTmZFzENkpRgqK+/MHdTHQ07vKh9TPSQZ1LyRPefGRSNp
wF37CDb0sHVVIvxAso9iot/GZ4mAT+gqdDCD2Y0+G0KyAgm3KFYlvynzWKC0EEI5nvq2glW7A98M
AmLdZlvR/BhqviK5qecaq3NoaCcgHr1v4b6jYayX2NsWs6NhwZm1iQ292/jf2XqzcHlEY1a4w95j
FY/WIK2yhHvLfFVFJpZ/M0GszWtOHWpMO3qXskcEb16de2ikVdc5Usd2652dL31hqJ/q4C6LMplb
rYYI5qaQN8kRUv1AYoDazlveRqEF08wUtn0kKWbDsc4VSPyiZXpI9J3vdii47AKf1CWpCjeNiGaQ
2js61Z7xA9ZEpzvTTK07MRbeSD1S6AeAvOIY+1kWzJDBGatjBqShcH17uOgYI1lg/bPKDJujGr1S
wXio0N/Kvroswb8uuCrzbK03AFoMlhqTpapO6s1LDlJ3nnlom9G30W2ONsgbrOnTQJWPjgCvNfaR
JT+sktM++fZfzRb2yxPWm40bqOvSq+knkCooM35/m+7zrFjzyFGEVyW1GNzGYyXoY55YcWg368AE
bSTg4y2GbXavdPyohpFsca2joPeE+MGQJcW6wQrXZreHWfurpEhHuCxGjkbOg8DyjlyMItfm5NhZ
k3bVAkZBM2yZyrcNCy2iGI2SLx93MjbXFakYSZm8DSUhAk8nmBv4lUXvYoCa09GUvUq3FposIkEf
XO1cpm/B28X8xf/pd20+8YSMcf6nURzesJxvMrBtr3pwIDZa4mqxLnkDpdcg8Tjs61DAfV68SdOe
hKAh3aH+LS+2HsQsWagyaR1KggoCGKLFB7GE31BCesE4qyj3oyxEXv+Di9UYQx9PksBlSuFc2vLR
EJ4CC7lmQcHSSrp7x1bdOR4LhSW9Vi3O2/sow3gRQGStshmbSceKvJ/y05SQlPqgoQ2EBu95r6n3
Ffvb1h63qBYN0B7U4kz1wMQrhzxkqUWzbJrIbL0nvqI5w2kvyKddfPoRlzLWnosbadpW9ivjXMBX
i0QXuoPlWAjRQZpA+zWCrJU3ABTvhLNB1+OMRU86RvKCEqkSQ0BwZ+4RmzKMwBK7MrqAy1EQt1Tt
oReAF6M1TnFvavtF7hYL9DKRXIZvt7oswlmkJeP45eOdcXdxFEgiMxHy2VQGzA9SdldpPq/hH8VJ
I0yPftfACbNXw1Ze41mF1GuKYv0eaBMTbtuAnvZ/hov/MqRiE0DjxXRcpUxsr77M36Qu0WyDoUJj
wryNzcFwYrxE3CQHcXnBdyPX8Myw1aaZdCL2fAH965x+TvmebJb1obucqimLgI1zqt6TGcsVZkpy
mZnLXj0Gtn7wEANuI6K62tSE5H0RfvO9VqvtmbcOAUlbKFZfnOuDZrjuSJVHrJxixQ4d2Uk/nroC
jF8sgOlcRhmuZo6WD1WZMsM84yXs+c+Gump2HXmuh707lNiTzuhiBl4MYz8aO1kMkiOJJv9S4YFa
hR8gPgd5wxTJKxgA/dnTvvKIofXNqX+eQ2KjOrsbn5vpxA4PL30lKVv3KrL6cCjuO9WsTtOR06WE
Z1VP7+IfFqed5Z8hytoWIONYlPbm32Ixrr3WZlz23DmqIb5+tvukg9RAbFT6+2r4iUH3PexSNPIQ
LMCLFAs5IM72OrVapxzf3zRpsWlMBlGWn5yK3SBg3dNtmij8TFzSzChEOyhoZ3ZphVnBtf3u0S5B
ISwsC5KaeNQK/r43zoDsYF5AQnlig4atoIRUEBjcsYMXzSgWeYtYx6vIq4wG2E0RcAXTlR4engZG
RpXhVExpjhJvky/8P8x2QNFg0MLg6ue1CLgMUwdLgkU6TzVsFdY8S1YOCaG0yiOlL7ob0ZfOUL1G
ZIYgiqD0XVBl9kJg3ouHpR0GyUZ6905ccRzCYWHjxuFFYGmlOzF64l/4IOXFip146Dg9FJ9gMr2w
7dLzjrsq3VTiqCZgO/rcwvElEnaoxSCvfMlXCAeU0ZLK5+J0Rgoaq/VyfQYEaPECLoEDEgu2C0yZ
R/iSbxF8FvddiaxMXKMI0PtcxJIJ4f4UDpJAgE0dkLFzlQou00ghN1BvwcIFHbzA8ZZ8Ghnf+8pz
rWhNnZNNUwG6gOnTusAn0ZLj9j7Q2ye4l5vp7a8WFa8NyqI1Q8xqXF0jOV4rt/NimNtEBgZl6DQi
8xyt2msodh5o5aryzVnV6CZ77Pb0mZLrrBeqgtHgnqAmZmvF6N1r5C9Wxb7DyFL+xUDF/V6cQoLC
h31NQAwFhL0gcS4vPZPxm/1H6Fo5XQeAcrMcuNvHcuDV9diSv+LDP1M2VxU37ELxVIr9uTD0gJOD
sInaWwEPUKTCi4xCmGz6GFurEfWK0JpKAe5SV7PVqUnSvuJRu+ND1bKpFEvhRN4fRMPzxpGc0CT3
FOJyTlmbRVJQwpvwYwM4vkCT+3QUzWeUcfikRBowV+FdiDjs8kSH4GasDNvSyQGR1ZJHto69e1qc
gUuvaDRKRbYFYeQhh1PeTVZNfjU2fEf6IrpqsrhZbq+bXqsmHhEa/6aa/Yt+fiFCvvrwek3/fJeB
Mws9wjdX8L7clXM9s/uyn2SYReLFSFkad5X/zFZjOgJSJGXUkKFpSNpEvwizovIeEiIMbUM4sBy/
YgnDKDaOglExEBTnJpL2QAANu8s0Orv4Buiu/z9856aUiB9dJHvCroyDkD0gLvn4cHgEGbiIBFLG
aD1EN+CnOXLvxU0xOJftdIELeTXEy5pm1FVfpvQ5hvkQ/2Sm+k2v7oYMWnhs704soWJrQ+26h/h/
05qo0U/CQB1KajkyPD7gqq9fs5d+APNdtYI+y2OSL4TZ0DLxrp5g/oXsri/Vd8PldNz5rZnHuSlL
IaTjjHKDamjfbZjC/T9YxXoz+vg3v9PNTWIanbNwRx44sOz+1nemjyYukmnx8cbPU/Peuon+7MKj
GxYM67xDtH0b9HKGxbdZbecmuhv5ybszKKlCHx7dWtbcl4uZulWS2jULfAG+No9ky5WDLuLxwpOQ
X8sns03c2gUeMe+SzStIUx31NSOCZm7m8vtOZeX4uATHsaup7GD2LGv2M9M1APMyf/ozmgUxvtmD
eVblj2gNJTiDgs9PoQJi5MI6hiiu0PJSX5vIFn1rBmUGFWWP0T22ifo0HllizsDBG+7aRzZXRSAQ
e6u3KDaLLgK+y/tbGfLBU1Xch4HlGjeBRjV+MEGi+J6bXb/hJOFrnhcai9Q8NDszMfQGwNA/rqNT
MKZe1p94UKUi3pwuk94hc2l/Jeuuwo9UupTWn3oNHtYOoUKgXFCm40XmrvtrOgAlr0QeZMI67yOV
VjQld7uUF4vyoK17Q2OX+V3/yeQEHiJ+NivdiWqe4+FPRADPzh7HjL7/UF+CKNWMnL57rpFJwPhu
PstkIunyOc5OhfX3iuRPgNOHaRryZ0trsiUxdff1kZmDQUe/9YQVr5pASco6lhwxM0d5oIMuteHu
QW+ZC+dM19K6MOvCgoo59xalvpCaPGPesphsz6I/HuanBbshB0wTlydiCn47l/paK0JsNmIGJORU
HJwoM6JPUQDukkQ9ol/K08DtEz2nKYCX+HpMtkRZ+whIUz61C5HMUMuguE7CqMEMabd9duz0SAvx
VYBrk+8MzCpOATEPDCOO7Y54IQBj15SGWDsBiYZl5Pv2p59pJA/xtL6DY/2R75SJsyizcx8vx9cR
Zh3JCbntbnrfhD0dT+1zj7fRuI3kT0McokHC47im9aAFwymegqF7Y+rPp/0GNTyCjSf4Fj/0H5ys
MAq2J/+A5mIHes0HUTT/cX4UH0eCGOj9M5wWi1RuPwlE+LwUZrIkXqVhH8yxR/rmFjnMpNWoc+Vw
gP9PLi+CfYTD1/PQpJANVWEC2KCO7ITGO3hJPEO0LPrcaKt4UOXvxjGhsObE8v/ZEsfzPPpDLSGo
tniz3tmDSckm0hCH8S7bKxsJZPoDr5BdzyJrRYoWvQoZyi7bY49Zu7Iv4DB5s+K/Ktug2L3uzEeP
M8ihR6xcNNCVI9UW95Po0AJo+yMjJAGfIkvS39o84VtXCsV0RTIavxkEBSg7loY8JIj6+zk21Vmz
SZRtkZ8Lh0sbmcSo13KNfWl3/gsvuDJcKUlcoWd6NVT7byaEbaCRRqBKUtHGjEdkR7sRX3RVgnvr
zMQVHUPxmOnAa2cY9nAH8RKs6qdb3KTVqVOYNWbdBfyorpY3KAp+oN836c0KkdToyFzAtKjOZwJb
nGcTwj1jU1fh9mPeN7GKAWHP43yTynqAjFhs0u5FL8d9+c1nLnF1b0h04l5ONN0tk9LdhPq9p/8f
Yo+A/tXP4a1RMCzrCVdHOyZUp5iFUmWsEd9z7Ue6SFH0tgzYvk1Mqy2rklekV5KywZex+6BRMCIK
YRVXRY+Uc2XiSuCiOfS5BAokxOzevRyONQTzYzk14mLrpF4kj1sipcT138GJwskYXRLSMSdgFSE1
2byhuDRZ0Pr8Si202vUAgSSts2aBfnfgvb/YsUXHZqitDtnH0Cw61dkPQ833M/0lcFUWfzpiKK61
vWcZvmHxwknCcie5NdaP/5FbK5cQzdaDxCYnExpprzdwXtsjC9uEyoMtzl4cQDHaDz9xUYAeN/4J
oLw7GRPtsc9XTfTugnJenRpg/X9jvonNv7IDZ9fkAInS5KnqNCHYnlJTyH63N5gdY+e3RO3thNwW
KRSWzfdU+hDcaUn4/SiqelNhx0R5uUE3VzR1F1+AqL1FYkL2agRyMgjh2WSIBDZr6EqsUdp1m2LV
x1YWgwteV1reD/haGucFq9nGbv+NBrjxaxI+/71DXOhN2Jh+kvuA56olsLROelzvIN3It+vo9WMB
yzuJ7thVTh0mW1V1R3Sp1gohNa8qYO7EI5mydCfosnAed+Ej4f8g824Q/GHddWSounhpxHYKqvMD
xkOcXQO8voqNCyqXLYxoyBdQQEjG7GtFJs5EWEc9PqfzdUR6ruR0blPBS/NA0ObFtLge9eXpyQd1
8C2myz77EDIeDhay7uzLaVp/FJnfezOofbkDIFtelOls8i6LN0VxT288bjZuJZBu+pWyViMoZssk
xsvyf8osWfJRGHze24JwACRuoHPy+/PbkVdk+9+BlaqM6l8PqKvhfjYRizJyz6EpuV2RrtZDypVU
F6jIQm93bZGHbheN/WcB9hk1yZ7WsBnTlTkVhhcxzIiGpn5Nhdcq+N/nz+loGWAYdoWibVrUnFOw
c2786M87fVzKaTGgOrhxJf2/uUb0gsr7Dn+4VGppCWcO1zuPjnGc9uaDvQ+XoRGOQiehOOJ8cTGz
K2HrHHyLpS3S+Ay6szMAsCbIer15JeQVgnbzp/r2MWuLc5X7JUJLpZe14Vo+7OsA9jI+l3ZTV76r
kHr/5nlmtlXjeI3fzXM4cMb9MaD5sYGvc2xKwo4dt6+Ej8DtvUAq/uFumVHWyKsSuPCLEIsjfFcl
QT64j0MYd0g48zOOKnoH13L2b5coOTKd6jsutAxlc/198OtJwEzEQ5bFnHrQ0Nwc9G4TLuUZ0+/y
D1mqbC4QeyHGg5rGf5IHFaMX5K/kyP6BN+lBt38KEMdPMICRbaGJHIL7ulkHTPEpaWj1zr3WXf9c
31WTQmVh+BevpZMyJUziT5WZOYybWnlxHIFyiNtuG+oQqSDV09yZoT5byoPY7kpChJ4Okk8tKdKE
CAX+FWYLP0pMDpPElR0q4CfIFbvszVBcAzXe6MMpCJswiYLdOt8bgKaltwCgCFxWAPYBruewJ6rN
3fXDbq9HCi2Hjia8PGJPChIo45YnaB/LjZZWUdEbJJDgob5BXD1e5MIamRT6oSelssq2RJDVsVYW
bxVSUDYyyJ8Ov2RidZTxLlqd9yuMRAmXL92LeorlUYeePOjsiV6OAM/dFU0GGQr6ciFb/a0VaUv9
k9D2MkJrNhjudDcAYq4VyDKFbsXmoIDeFPkUc31Ilra8FUCEiCUxex1eA7E6oozakM+/7m2cuihp
PMf8ESRNN0Ff3PlbReMygbEHiIFCn+Vak6KX3yPTjMmLBLZTuODYDqb7COY85mPqofJ2ippVuaXG
p0iOLedl1VDyA1ABDrDK2ccQAv2cPLuABRn2EQxPk7rrvW1WU2B4KCne0qrh3OwLnFy/fEP/BHRo
JJqun4VqKuZhWxdSZ0Baj3oi99aTVXrX//lK2T7s6rEeFDaDC4AgULByI+5y34700eSWWtIPPLzr
HyMKazfO02QCZr8N5oLpDUEu2MwXKvqeeTJadQnm9gYTMa7PyN5+CPvn47j2NGv9eEQD7KKRQ9nV
U8/a6N0Wlt6sUhn2x9C9qegzrUUKhLikHz0dwYL8HrHIdrbDcrBY4nqTSygcEU22x9eSZtN+OcL4
A+R8nXICF7O7Derfs1L7mYkm1CV7GN8ircGtRaZjT7h+5B5B9ettgpsFTM1VfUrp1sQiP0oonmsM
hb0Tdo5uHn1LVY5ocuaOb/QOoXOgnULEAHFa0DkhiOyuZYsm/FMydzIWLui+i5A/VYBJLano9LSZ
V4KMCZe5vRa6FUcPTF6/ybLAn8KXmPzpnQXolQ4fn9DFzHSFTlupV0ZqsPyejO3zBdd2k8ecKah5
m14y53GWtlSLUJH7dF+mzFrCs3CIau6RsdNGhFDm7uAwHNM0U6/d4VrfaoEEk+7RLKZGhMuwUXiI
fM0Eexl6EeCufHQIvjXQMrZbgk51eNGikfUCOUWNBwgDuh1jN5Z5xAAcPw7DKG2dAFz2U3AFDcWi
lpQfguTPorJfWvKHQeRocI+43vIiI+RAbb9cj8ldbiDcOd69t6Hfsjaaa+Rld68J7y1O+UjVb83Z
/iz8GUJQgVSJ3R7wB3BTis+Iqx7/t/ia+C2BzNGJOXeXqZmB+am0mksLlgg/6acXkyeTEDV7Q2mL
dJz8aQNqsvH77JJLvM/UlvqFrbgMTsPDxKJNIPA9gAXYSZ4xoOXtoBwk6eW8Vlx5J12YqOGqv9AK
1W+4cd3shl2zdY7qb6aTc2EbJ7okjZ7MQh10wUD+kk+pJT9DkV1SvBT1AuNQhBpMOqU9PXSRcMPL
7FASrnjN+2tp9ovSrkbcZ3FjcbYDQfDEp3PEqHF1Sh/cXqire97H7RDN97VQ9vW8LuzvSt0Ckd8k
HTbZBU7bdvDN5Magh0+27Ff+ggDboE+tzhg5KXRt0W1GfQ5DbSh/DZDbmc0kJW7GdGirDGI6Kcgg
D6UeaOWQwzm+tCgZ6BpHA4mhZ4Pnd7H+IppCYHD1JJgatQcjC/Hu0/90wYP7pxfAs5tBT8QzLekl
7cIaN54jjAr589WaZwnxQ08/dqCylorCWCrwtePBg3GeMka4xJDL5t3DQN09AGkQmPy1cib2gxVK
MCJYRT63OtzQu8SdlF3c9b0w3C9pNzir8SeI5DeF8vO3ViDWwESAjBh9zrRzHh+ANH7KUb1/tvq3
193DgsH4H9c54NNiOoRY3ziVtMyzK93gENjZD2Lt8Piq4FxNRLQ4K7SPht/XT/OtjRW5pBh9TU9x
j6oPoaabXlcMUEtOQRWSGWzZGryk5nKlvCDUhUNMxPYnDeVFPgMDgxIEHSa23SCbbg/NTK2oNn5N
/eMSiW2erpKDjpNOYPzppTc+lzEVeGXLZ1ifEpBUlixjD1jXagKWh3POYiTJpCDgub/tg6ISoCHZ
mySZWJZJsgQCBRjkzAOXgnZLDwA5ZkpL3oFiWw4B7Wy0OACzQtZOlr66YpZ1NTBgY2awYl5dqXWg
NWxB0SPVQ6TdNs7YoAff9UckDGfkJX4JCNlp3TK90a1GfjSZ+XQG9USMdY3XWkEbTo2nISAemlGe
/WT9NvLd/7qsPMwPLunowbTJ4qwKW9RqM/ptlNsY4Qf14FT0ISboC+mfs+VGTR4is01v/QlGXDe9
gtJmjJfbhuBucBDTtMOWJ25ADl1yPtzfnEAh+UB1SnvgpsDrcVyY+ueU00fW3HRLzt147ouSo2VF
9T87XKak2ZInWh2pLfg05DdGIariP29VT2eVl2O2z/2hpMpEJKcubhBgVeHNX40uPdacTc19g0wa
GnqogLACM12UE0KfY9jpSUEZ/6UaK5mRHEGslv1m4f3cjcOO4q5BXNHh/43GGezA3PrHH3jZaN16
knvkyK3kwVfsOryNCXH+tzqR4voAobt5Ckyv29X3R1gZeAf1NxGy5nhxk65h9rMNrv70Olipa7u7
TIRwyR2oro0kANRR60j/cXlU1JSXBZYFZZyZ5SU+gQ2qggaEALBsx6AVcaTeJ1UNU0wLkZEeC3i6
LKs1RJNApCVFFWVNFAIYftdpYwjwtJkiQcf5uChY33e+nX8M3XybVQsaGG/yufFqY0630pw6JRV3
6RD4VNXE6hDlvSmyvKEjLSY7DbdR+eIDDkivJGVzm5Z0y+5LLyb8hA8O6OiOjYkXZHM9jqgUukaT
cbGcRUJlasftwHCHyERp0wDffkPskV8qcvKey2x1aznvOvP4/xNVjHxGy8tNtIPrnANaPmCBW7gg
ecXBwD8LgUpoB32c6h8o3xDaVIq6WkjpXkXkF500DmplKFRASqeWVmKQ1QqrBFILbxnMcN+qdQ+L
uQtoq3gotZqTLFZf1c2bD+oC9aVdjzA3y32eqENJIKhie5wflxEPjQA4pBqQwRrDItl28ttkBPKg
uTvsSsVmEyCG2R/xhdvxDj7wJgReT+e8Oey9gIQhFcba5BjUZ7P6lt12vK9eqIwEgpUccjopvDkf
BMir2UKIBnHqe3suwsjy26smtBCVP4r0YT51LoXnMzNhvepwb8YKwhBNiLWyjkYFigEXRrYuxh9C
MBfyQzEwjd9Tzxkv31ITJiwiCuWX50+HVOURWAXTK5IHlvr5bhp3ef1oNRNiV7KEOhRyEGdAIOtB
DeX8i7UoIGmBo4Fc7Q9WCBgl+aL0w+NIwY9AY/MFZV4HF64eZGX8fofxiIGI6IaFes92s0+0BHnt
w8Yzzk42m4KAncxoghfo8zheXJOqfADxd0V0jXPbUkfkuxfmFBtlwPH33r4XUxEH9nwy2MUHbtFg
2kRf627zi0uzE+In/DfI1NLl5ICpdtk2FHuIu8FYpknXmfTt/y9vHljjWWWy5Zq27d2PyeoOC0pH
ubEgkhmvA7JkT+Fdu2uIxKdyYMb7vkXSQ0VtGXeIctl7H3rIFc+JB+rm+PwA+v85X1aiLlhD0iQH
xaAgpbWcfVZmZyV+Hcq4XQWqJV/OqQW/LIGj5t1gbYkVjWg3t5B3b1Qkw5U/gPuug4I2E+ztzuTp
yUxH6Yly7/ff45K38U6Aw9aVZKQHdAaLi8dUa/Z/r57iV+D3YGUWsAdD5tKITkgW3RqWi0rVYo02
Q/qogWjjijDkoxtBvRlOC24fWFl6N0mxgvtzcFgK+nY8xOoy8DfOlbgki3oCTdkDlzQJq+PENzgY
zrOOooBvqIKJfc2wF3Z3ALMRT1K71VAPneiu1dbB89nFrQwpwaKKvqLzMDo7Gw553hVOviooCrvx
7oeyLHwmSPTrazmAGfh6+ezWIgo8c9alP6v/pJ3fPfPCTBVk5Qoupn6PfdaJ581wtv4MfmwYEfal
+NqJn5Cq+sxtmI1sJnL1s7iGRPmdslD5TmpXNeCEuCj1c2msLHbFZjKriaTztivHWYt83EdKnaV3
AOgxbjRGFVZKibyhyBBA6ObHmx6f9ZNc2lUE6+1kkXpcbrxWDcXwI06mWt2Vx5u3yeShZogIe/nu
zJ9pAzEyBVl10tr5dYOaEN7Uw/qqUFa2VATLtaeacmjaoxW9nGci52FgNZIDYCSD0rj6OLVyZyds
jAJqcSfSYHQbGqQ59SLwYseeJknQvX/8XPOFLD8MLM7K7tt1KfWjrEWJio1Y98ni0SF3rfW4iW8z
MwZwl9HOhUnW8v/DUaW4gvoDoJnF/SfmoxBN+GYbBJcnfQAczraFdTRV+4ZdXPUnl1KYKA5y8wpn
g5/k9ZdpLfC5tXd8cTepHvb8M4sJkNde4KJRp1JjYbzN3k/AnQu+NClrUqArWb3eMGSB86srA8ae
pa4MmUDDXeChQCCxzLhpwZD5S1hjSCg2z69s/MvnfoGlMFVhldCV8u92dbvNIq7tuOlXrCrVDAY1
3SkQPd3v8XoiJ9D3/7CQdNAax73GM2a5koI+Xq1Q61XNPCIjvhNiiotcurbitw88V733M5ToasFx
JEV1upBeh7i9AzapVGRfAQzwoLTxobtv0KxTUvgXsDQ0Jm4MJwhaR2NONDLEb+gHYCDAXd64Ey5v
HIDq/0T+AULtG8l9JjxiPoLBaJpUSFXs65MVEUAkgWoDYwUFaM5C7+26wjId/y7HONnJj2a1zEpJ
gXuR0faaNFM6UT62DwDJMpFyiTVZbc7EEJbECgZp+GRdB75sjM1rv5yjYTYfyKIgEcyTArdxp+Em
J3ajhvBelpKVdglIhRdotFUFn0R3xcWOoEtYePJx9UPVzyHCRw3vPSUfvan7SzMeN8pawPaWo2NN
KAMr1eewqMzxrLmkAC2cbV3fL5WYxACbFle52CKHFrd+QqMoXaHHW9BKZXpVp+GCdBCKiYNeVnjd
HQijuCv1kMpojYHIVNBpD1XHXPjNoumPjYPV5JAKpyqeGeKWgKwGS5c3DzL9LkM7voO1G2I9rLK6
SwP3JTYHIqHvf9ZIqDzIElVyxNxhRB06u+F2f3uvcf/o5K8Es4KWp/TRyK5NMOO2Ps0wSUJnM5rI
dPZ0iIpL2+Z/tiz0yMpMxv6U3/pkftId7k0iTIN+UqynYukvz+GtVUGZygZEe8lhlMMYgmhj7qm+
8oyud4MUncvBQGTc8fbnntYA6X1Jg6VwVL0Ckpmsm4pckhVYMAva/bXyk2u/M4Uprx+yus2WahLu
iLOlon8xOdf1Z2krKVTMVuxwSzaHyWRIlpBxRnVumbCk4L/xYHD0zrAUGBNdDrrXLHsOtwVU8kPM
+XgCtswVPaBxg1BbSQRddwOTI6/vkVKjZF4CJNEqiLf6+tP1EHf1AfxqBG48zIpFiC/5c36XubVK
L0+6LF+O/XDSG3qhRXN7By0uCpZmQAEgAZ+rAZX4YYKh9jWPunVzVMkSkjW4w11GfFzOKljw8V5q
S0Nip5iRAkyzwfwyc3F71qBUQI88+UIJu93/sjbXcOzcpEZ8eb9Z7+Yk7yBPUiihty6xoRTy+57c
rWMlZM+m3u8FWUienBvNyBeOBnf/0e7UfQp79ETgxeOvxcRjruQqxwieGAi7h1UvAHQbGSoSkPFL
7N22zrdhbZKm47N1UKd5BdnMpkg9RWzy3vezYhsB3adqEDsA7voGW46OJ4Ncu3k6rUA8TLWPhJ4I
qIyyDTgZx8rqGHqqIsbKfgh2b/vrOMofEH6pkrr/5cAqlDN3SQUnpZd/tkJVJtG/ZEv4tAVBm8To
umTp9ucaxBm5hb3A0vqtB//2DLJ4LAwsFMt3s1/ljxHVFln70aXKId9ySUVSDAEtJzI+gVM9GTUn
CXzY6EEFMp0cLz/4QbEdA1iXoTpczkg5LaoR+1QChHB2Q2raRAbHzzR9oJItgl1rztJwHO9jlFw+
e7lVo/zMLu7sIvyshf5zQTsrXx38xxS7kmLEOPBroqOGchX2FbrU1mMOlGZ9y2+o8OFV2Lf5/NXz
Nnk+2fC8Y9e8f8B1+LKBRHydHEXYCQ7lQROjFY30Hm4aFiWee/3FB/rTFgEfEkvhe4MSAnvCWdFM
/fKhqtxhYmfX9nMc1Gem6jMt3Xu6jLNILcbKEbRFxrxc2muD1LvlpVyKyOySbi0XQhonjGNanXAV
1ZGUCoF3lmcdbd9sUP9rvqCKv0h+blLQXK9T7KjNpWN2+/KhAAxP4uU2lhuwyRXMJy65FH8TbE+1
IO54gKuOoR3JRk6y5/KmHKSKXG/QQ2hOOnlxwmMnEFfNRf8gNkHHSzTUOq5ILNkMLkrB8HHjFl+p
SCN99N0biAuFHv2AnlG9p/VxBHlMCElbn+WjyOYFkEzaRqH5qnE+IFdS2NnfY+4taMDbj3UtYYal
EJD02MjwwqqbHd98OrhaOk2dHeTEEv8YK7LdAauDEJXGBDu0sFiPX8tlI1A5cZQPy6P5C8sqgtEm
ME5YckPhRHDYzoN6M1hIUwgCxF0jNovlJ1FUklwDzIhVxeDk6i5kr4FpeiWEYj/Y2U4+ztagprzp
8CF5k+bGBx3AmbR2OeYX8A3rf9pXb9CyRMzOISoOB9AVbv2jsBHslmt3hP3nUePTm1DBcTm44dkh
X4e5WBWG4BJeAHBOyPmiMt+SIgHc2E362Rz70FBWcBQaOuYBqOClG5OIcIzIyl/qGYryIuUb3yqM
kenswW+OP8QIa8x5Bn4R5T4Gu72AMJi871bla65odJyjbrU5pfWD7MqeLX9fIYQfuJx7IMmS4ocd
KEXKDKaAy4i+YS5PX+rFpkjCH3DJ6m2jvIyt2vIxu4ARH0DfFBpGJM03QYWgpNUWmnUQsWpAaEfq
HiKZ4GL9U30PzntGwClhUi6r7en/zO7lRDC/hHHhWnPHWRf/SjMNq1AoGgYf7y+nuK6OOOZhbTIG
MGT0+xPzhglfYuzDEf5YAZM+CIEsoVqZmFN7biyuhWJRRGcaIpRbae/yTb5eHpEmt9gYHgQeXr/M
lDa78LOiEV3KaNj1XpEhFVsplmXG7o61WBYx4A7uRbi1/N1H/Ll/yMLWeLXQKDgqmiVHNVLjUC3L
YjkNdL8Uv1w1qNKkYLkHUsyBkNUOguLjqi7ufJKXF0ZpYRFhvCO8Xod5QGXH+mHwd/aJBg5XCGcA
2zm2dfGIWl0XN+1SpHj6Kc7XROPhQzRV2g5mAv1nJ11Ph3kavm8mk7y22TJez1BjyS5/JjB7EYsR
/IxzeYj13azKwXyJ3CIs3FlJs/g71znkVMS6GfzYdqbWHaax78AAKp2mvi5BlwQeZv2kZQLPUL+b
NdR6kiXin4l6hy676WwGksUqh2LB6pkKvXt0fOM47bzncN3W6GGRbHlqtni1r53+HKbhs1aWTWr4
ZLLBCEQ8sUh8BTRNDgiTQe3wid0GZSw+BdUilWzdBk2AL1967b/q1RRp3EELVEupkkItn+5fdNo4
ftkulfJEVvhbGHNX9lh9quLbOqVIHzaf59uuNKxqbCZcVZyU6mkzCSaCLlykFsoWup97XgIjbGLV
QMRy9ZUM8uN5KbL37k8djgLJT7008s03iPabXPl/N3lwHNJIX3tSQn15CprxNVoJ7y/x78DeLgTw
yaFqCmAaD0E7GbIAx/VoTclKx+wNj8W6HfsQoedPB7RZ0CxR7KTprhJD8cWT3NlzwGi/Tmca0Tme
ZwLPk5mKnQb2VMTm7zdcWH7o5+gfiqJeyAXZ17WQ5CdG0MLxvVCkxFyv6vucAf5rq8vF37SJ1ApC
WZ6kvPfUI3y9U0hZAarf2rJJWD/7wdYzHTEqM9sXYXsG4WSmTnYpBMXjFrtnw9YEch8cKAKw8Vns
7zfr/vSmh120M97ZfUIeTxZnl7Dz4POJJoHtx7IAUzjifSlj5+kH0uaenw8iw7l38ytGT1RykWgm
dpGndvUD1I37vQWEbWsXH3qEQi4yAAEo5vN65Ep3yIwgKFKHSdQ/+Bma1rqpbf6wkZ9aEla62Y2q
pXbu1XLFpwOYWfTRwe5vSFw5khOm653zv59dXIp7thOO032FarlssWIQ995yTFRyJsSm2ViQhQcx
C8wLZSuQHFI2cQS2gK0k/9FNBH4eiR1qCvXjcDcJGbRMFMnFGZlDeRXLQVHaQZwflGZAqw0z5Unj
yAHtsLPIYYyS/D+eqb0nOsQKR+7gYnHCXup2zv3eodtsZaezmn5plUdha5H4n9K9Li0cdm3lDOAi
xBB81MutZYxSsY0UZFFobpBhrdi1D5DWbkJ6USmGc8pc/jSYrjpyGBiRDsrgk4BbIpqyr7qLwDEy
b0iTnOP4kjpjxpfLl2AZWldR63Uc7yfZECe1eho9RKjHAvfIzIrraaGCYacbyQaLffnFwbOdYA9I
+tGtCgqu+X8bOVTg9WGFU8+rq9/8yshNiKOVGp4LDThz9bjnuLwuKpw50d7Qps5OZDB+kjG7yJRD
k+SssssZsfOix5d0bzHGH+c9FGWb254+WrvLX13A5kzTOuAs++lbNiZ69cu4XuGh3mJkxZDnPBZC
dryctHAFyJBvZ6XZyEzJhKW1vlWRr7kUm041Q5mKvDnWFVXZozqHeOOdMaOoVVBXFPa7NbqlzNe4
qF5LLtC7fLh1p/cyHTY+XnWGEip7yn/XlQrxyMGS+sen0V+lTs7gF7o1HTIPDy4lpRNcYrxGXtgr
Qt0KtGqciMS8U545IINhDUgOXChjZ8NqWn/uDTj3BltmQbhzm5jbUBXKOfQk97mz96uw8epV3vxV
Os3rPkOlcqBGieFF0n9sUFrjiEe8S5hXEczs9hWLL6HsPTzTcwSZVsSOavjvMJ4G9+v+oKDzuceJ
U/BrpiEj7s7GWm0UI0F2Ba3qYLwO9gcyto5K097VdhNI9UaPFD4kxkrPQfFDO4F1mFD2yfWXAq+2
g/WQLwW5X0Hki/MVvUTtmYVXvrodvsfCwj+Afx8JFyElo6Y6U9qES+daNi8E6Q8WnrUTed4EJIA/
a5rCEAJabAhY2gbDjJHmjrQ/xybdDsHEQHB3DDKVqjmi3c1rC/PjoQdBA3xpOMMbL1OhGqbHYm/R
PpkMDzCdtrsdFH165Z+U6V/SBQbQZLDZ3BS6YVzvBuHT6UfewMsOxYX76Jj/UdftAHiURIWOF8Fz
KO9WDSU6GLQzeIG3+uQcZxWr8qYH/k4x4kACuQsqlC1U/ubtqDF9dTdqMdQ4mWe6UINzfr9F4FGL
/UgF0K6YUgIQ4uoPHZxWb/FQtNWn17LWoMApDa3OpzWF/UzDpIm0KWoDz11qVcnwQZLIcLSR5EKl
zWlZMPE5UgK/2jtfYx5mQUxUiy8OfwB6gewV9tBSobLQYpF/7ZuIJrRLb7eXwb+xOKeIl76EsVgE
nLrfTX/fDNZUfDTF8DYVVu8Klr//aBCGNr3LL4r2x+Y1VumJ/3H4MTuXloCBIxhXMlBNMiuWerDl
7CUYa88MqmBYQ7+X3AA5kOXZ5MISzySAvLzHqzIKf3MvvXkrrfzqG726748GnApSEDLTIgzr/MPi
D5YgeOx/kQ76nue3GLm/fjF/80aj9i9436hQNiij9vKenyxmLI2gSJ6qKXpTjd00ZkMquEN9OlJ5
Z7e6Mh5DochOK46xT9JEGsTTLUFDFUkIyAiyFToI7wltKWvN+VfNQp4mAr7kCZWG4mUec3jADHpo
X3K2tSs18hL3dbGt6PAIuVa0dvOtdDz1vUMH9LQmiBzZCIQvWtuaLyb2Z0ebzOFaXvlWaFkO5f1u
xNQHChmV8d2abm1oClVusVVDDAt2T41VrhcHoKGL+/kBht663ruMeR3NzJIJTg8tgAC0Zdues3sy
Vwhgo29s0nu5HNsLnkaKuJr7T0GbB6IcqLe1xpkF3IVWQkEuzDa8FhIuqJUKuvEuhO0zUwxpmcrZ
HuBW2WD6+VFfR9BsVt18T9oPnH3MBizSE/6b328tHz0Og9oiDiAp6nxZMKJYdATO2YXKbdh/A7W4
SakT2LjcjiUoWjgHUEayVHxHEeJZ0gDPzy+PUI0xq9wbCOeYDS1ZlmY35L2KzketpFuRa8f5a7Tq
l1hZPDKal8zk72ILCjcxNB6cvmfAhJsZxHOxk2XxWTvjLB+davPu5yoz0czkeJA0vB79uW9b5Tei
lfo7FuYnRrRqjx9dNUNKtgyaiB5L157ooE+D3oIttc1LRr7Ama+s6vjNZekW8X3tutNJVtONdU5m
/3fEMW+/bmNpmapbFzQEKTeKMufGvqQZ0fHLGV8MO613LgBKHdpCteCCPGl01h0def5Y3A8ngZKc
oQvTTjCLWH4XwhsDU6lB9rvyRjkhaizS8q6iMlklKsD7fxrILcFD6emk/Ml4F+l7D9JttKa3Rm9f
jvQbzlETc/M1GUaFQ8NhSR8eUNCIwkd6HNNx+6n4ZdHQXEaK9W1unMw5nS5U6GPe1Q//fQnQo308
rBfMfFtzAt71xWjS23Z5s9UnvQVDtVPJnjLvBnRx7KfhszulgXZW4obfhqdp51W+FU3b2CfIiyNZ
WHVn4nsjnJ+3YriTJTfFPlvDjVeH6O81O7tTMVev+RA8P6YFpSvrLWl58bge0vDz/Aiq2hxdu7S0
OzbBif2RDXMC7kkCEo5p+mR7JdILcaDMjT0GCjrFdxMWISI456Pn1TwLWfbz9UW7ebjN7i08j9pA
F0eAJVENIPbdoeGnM2JhXrCW3o4wx1QObTKRvGUUsEuvyxPlD80qVmKvpLPjkD1xqsOjqoBpFoiQ
ju6uR1HtIO5+q0J+FpG+vxxfq49H2rhkXUEpXJgiwGFH98VLknLm9dKIN/Pw+XqmdC3C5YVI2h8c
Y3uol2pMKGjCv5uhnS2Xf5elm7xzYTDKHQUwpLb5Qa/GzyTN+XyBGAoBw4TEgE3hBm4eyk57Yoe/
uAYMe2spNrj+S6PT9WuqWbMEo707+J5NeKd+MZsT2J8VCEtmpAnms+Z0Eus1podPi0J9wNcwjsMe
krRmCqFnDM0ddw+ukIxydFMJBbVBGGnK8UCCChw6RiDylxn/72yFat9abD3KFcmVpg0VkygFviPQ
TYXzmHiYghitiu8maZEYoq8IbGAah3wFzgSlq13+KpZsCVx2t93QorxP1TF3K1JNWHIL+cUFjdWf
iXBwq5z76+cw4MksTteK3neB7Cg1v0Nq82+1qL19qlFAgBJf3BfZvDA+1wBYxqqbV6afQ/dxtIcS
uZRExjOXmPE4KdGSXnQsXKrdmOWvjR9e12ueC4I7g3hzWJPwRPVpDLvU0DY3h719/R9bbSEnHV6Q
3hXU9w6sRwJtHD7L2lgFSIFg7nqptU0eARfE5fsU/Ys7y6Dr+KdLFUs4AAlszLVOtP6zf3kpCKI9
YYqmIyzjG0+lvXhqBJHogjKWBQD3K3sHiTGz9RTeDG1YldUhcAqmKLxpKx8XqbGfDbLpVlw2YbfH
EIdkUiIVxD1sg/e8N9neTl9WNHYvgOomTGd9CSeFqIsCrbVdaAVb+tbdw2rprg4EHIlQROl2N1NG
wzsRFf33tELd+XVHChr+/AFL47rbye3mE/La26VGhpRu1bMFCWienWgZX5ludveJsuf9/aU/vF77
69u/WzL0stdZTvdeHAacP81pRosgRCooqlnLB6SPyqmgpwQMtFbwiQVIhDdm5xZBKVBtVBTbqeZ9
PDhu8aGYyOENdffJfZ3b3+ql/rkTQlhl34hD9sYfI/5AcLKDPwrId60HrEbVkkrhmtAmFDBfndr6
5GMmrGLrhQej+B4T/oSzBW5rxBNa3ID8SwHLvpNf2x5yVrC4jCBH3n/x+UDFOKfqIGR6YEDnVyuq
VXnrqWB3OLRUyqhqNm7z5Z8zyK1O7cOgezYsZLTgATi7rUBz2DtNybew84Vpqo2WyejKpZH8naZq
6ZMm5DibnBoeKo0R0sZ/ntuOGVU+JIqd04SWFO78UpquqgUMuWGuaJ1LHD/wZwkV8a8Ovn0ey7EP
BbfQznLadF7wZfDwH9r+9iVQGK69mlLhFFwxBf6lESWdJeXrqrSLYj6YNru0s5PqXBWcFORlSYiw
EzEBSu6NE97vGufzTF4+YJxysk8QqwTP7qqzhTeglPKDc7VRgbo/E9lUerGfeFhQMlhw9PPvJeI+
HCqTcu+2Wqhtu6QSuV4HhJ82OyBQesmanE9PvDOjXQ112gug2u5o1ec6tZpYe78r8qNfB/ExLVyU
mYiItI0296zug7vTHGJReHO+2MX2rkrxvxK0uTzmAYQF8rEIlCrdTs63bCrwbSFgYYHDqc3UyuvJ
i4A1pnwlxOxH5umUlJq/AGR5iP0Wav14ox+nxCaFiNaBpfrS6YBu1iU/Nv+Io2Tub4VxV+qwBjXZ
ouLvh14HtsjKYFbmT6AZch74IVbJQm8m9CExYXGj8Hij/KY+XVoGTFh0t+N7/O2iHEyxVEaZdmte
qSZ4dlArFpfkevZYJkYBeYHpvPgQ6kzFozDfVygpm/HJ1lMFmZwVxvn5NStmHRdkJEPxgoj7L8P2
v2cLgIzP5C2tUaWE78yYG7YWgYOTsr6DJCx88CP0ojFdT198J1x66gAGA6PT7g3Or73hofCxf4Xd
/tF47Uz63x2KOvj42EKBQZojO+++HUG91U+Y6yAWOK07Yh/8saJHn4kOksUi8gG5GfCVBfa5YLS6
DpgYui2S0a8yb/y6hL8T+J4zfqNofRdAgV6Xsa7EgR39Z0nZeHDZ1zXfPUipqRZkm08+DgT02+qx
56W1zx2n8Oy2+lfRpwwDfgZ8++L34TgQeOI7TA2UWsFGZR1OaoVaU5tE+NLsTabwP6rbHL34qrLy
m5WxahOYaFIEkQf8VYmLblqV+oom8wRZ2YaHKr3j2zjlymP3PBQVjZfhmt/gmgzLAVUf4sN4P2N5
1Zvm18YqCmwNmmSWCD1rakTpejBVTvOcM5S7DsT3ib5Yjvkp659oSERYw3jpMj6B+i3305yNf1Bw
gX57vXe/d8x23/2Z+nR7UTRwQxDMqzqZcxblXsabkFnxtAHuPlwKkr3cadDBCfTOUYF/M7MH64rK
VzgDIGcNTaw/8O/K23MOZ9tZQ/cNbpcLSQXzWxNclYSG5OLQMCFNdhtHnVgS+31YBcKd8g4XSCGH
KMhs92enCkpl6m1RBoGME5rOuLiG04kyXRYGSkNBt3P+FWG85esKNFsMfarm982WZvA1xsSG+tK2
ppDbZX493pRrCvmQFRzrgCnftnRzOIqhuOFa+w/OQCgjtnSWPsfH9DW603PSwmcpBT+Q6vuFgbOM
onXWmsoUeAaw3ne56DC4rXUsnW6p+8v8foXnjdxW6YvgvWnmrRsosYIHyBO1lmZTONpUIm/P01/e
8aEQKD2wsHDsnFzQRfyKyDPhGemE/HUjRBScAMLk07wOQMTJil1RWePW7b1L+3V9qWD//nJhGBwa
uZZRXE2B0Z+Bz+KAQrWHQFSJVr0dLAGDQWxhAW7KE+AUZE5w1DTo8PVnAD2q5Wxhz2+i3KGnb0q2
iDWtLLJD5212I8OnKI17RMVDVEFMQMdLu+jlfcd42IGvdrCyt+maDwCeXvmwlAT5H4+VwMW8oPJq
QiMy3LfVY5GLFXA4Bxfur9BkH8TeEAYsYVWmOiMEkvK9n09VsLDZxXRQ1M5BVUh1Ky2e9zH1LTeK
t3hzkcCr3T6qWUpsk3SEj+pCcgl4eJ32EFRcUsKWXB5AWjp7d8tovEpbJF8XSdCI0T75Mjl2wzPp
JgR6qXryh62QTgBtLtfr59mychGVLa2F1O40hTaqboOkQY/DYOzVybWFoBQrT7I2RYv+raRdfMZN
+n+2gVehHf/lxjk534KWA5Qc86/w6SM9AyaTOAVqtIQqRtWLd2lXuiLWL6RXz7T/1OS93qBQqyRq
mbLdvIX37mkZj9R+Gw16MYlWOMkZhJBHHsZM7ZmGErSNgfLszM26mIs9HQ7PT2Z9Hz2N9CfHu9w1
/vV2xZeEOiCk++Nym1AjlwtzZMPK1S/0N42w4xVd5R9qLEoS6BYY3SCYucK9QnNvUpcgJdTZ8xB3
Uty/h9Qpq7+lXIlqW6XKsSyBdDOXK7QOHC7niv79MdaqEbUZDgPM/0e0eL3FW51LexI1lJ3tGrNq
1e61y5zaqTF/VA+IgNbzsJbIVLG1tw1Sq5YpWOIC3KZebZaP+6KBg9aGRKcTuv3B6B7oEOXmNEgH
ylRIdAzEtCjkdYXNw1vlwRob3tqfVe/GXAZISGfR+9M9KGHbi+Z42d2007vI64mnPoMbKP7ieFal
DcEDmNZFu7acE/EdIn7VRQb9lIovOw0Xo1yUhwuWWFyEe/rBfjNqtr59ETVEcMhF3k12jPDLQS/M
f2Rtq3Krbn7TatqGUdrMTRFs2X3wKxhM7xaf4hTHjff2sAquXfQMBySn4lvVaLA5eecqqxF1fPZ7
c8MSCUuy2WXdOW646ix1PaiKAvKiWy60h4ih6UlBVwvYrI2N1figqK9eP/ubmPFonYov+oWu7c6t
e8JoP9P7V2jtr/6d0ZNjZdUkH2jazzHnFxt7C4hZQdrW2nrzC9taD4yXqjcsGWl/tOFkWJD6lpHG
exCj7agI7yZIKdWrtjK8qvgXmACl7f2HAFWNrFDIC/o5H1Fv4HNBrSqM+gAhAQsMrANqNqOZ2S9y
I4CIYNp/dwfdf4ysBolXUFaTqgBUMfUuJWtH0LpmIP/y6ziPNADAOvXyTd4/BAdyyvDf1v53bXo7
lfaXWKitDkRMb4TI/iKXUpo/Eh+B+bXqVtPStfoxyqhtMrStX7EIcEF2DbxEo+5ISoWOkf86DR1q
4TmBp52bmdADbHoVJwjRi+1fR7jL01wDMvqix/RycRCKHvJxDxQB16oQS+jhVAiJt+Xt9K0DVJJl
9CXgc19SdaLSmXjK5QRCj9nOZZJNT/gC4Q/VFxsZc+DO4arBlk5dWQ4ipDvRKEEMraCnn9Sx4WIK
1jfkGQpkMZPY03F0I8c7vjn82NOkhSEqqdWM8O680Z+YowNNw0sXMUcHzjs8KGDb9RBHyi7W6Uye
mV6N3ipuKOHZbgYYCeJPn0j1hSsZAUqNvDGgqTDIVatQ9LimchrAQfwEF1eVDf0cFbp6djUEK4B4
STYqOlyKvy5fsT7dCN1FrjggfeXIMBLaTFYSm4uiZ8XcfykhHWPuhX+D+s1ziB7W6kWcChAj6Dta
+Vs3C2JRRqgzqxOCweauS6eIeAPZDwZAqZe11KwNG4DvgCDXxTn2to+T7FwwbXIwVrWLhumDsp23
eBUHWYwe5HebQB+yQuyQx681Q99+K82qVxBbDFFu3IYq43w9wK37GGzORWZoMWBlwfD974x/rizp
varl9ztt7kv5TkpfAlsCOVP6p5uX2pPjP5ssL9+a3B68bp5o9vI4amBjKl3SyVNPLKUyf0Ac3KXR
/8bFnTIByCibzyBUrsvRtmKGye4+1qGUmbcj5mmrFKHF2Hd7l3vORvqHmxaXdVUo+GQ2T/W4exVH
kpG98mEhig5C2y0Z/tbiqZE9Iauc99CF4/zqxqasr1cCrOT0IxGUwrva5RklEGzPTQBqtf4VxFyA
TVoluiB2++2323bVZL3qcEFapljxx8ifeHnOFG6S0Nn5cHipkGA0kBmEXyv2QCkBO7L0bZy9hTfS
YxsgN+TzjwZBYErg1mp7U0WecNsXGEXaqqX8sXGPwXdh0cWJ9Jhie6/tGUrKbvzqgJivewelOUqS
Dpu28BXSkcn2+8qT6vFAqIZS+sdWDZePPpKL4CMO+R9XyMLA48llDJd8qnU18ybZl/G4JGe6A+MO
EEhJ15hxCnjAG+iOOINAvs8DwQc7BCXIo5nkCwVE4eGmg1Cxe/TQg0XOh2SGZ3a4ykHCz8X8FFpq
ZQWrIqrA8g1NnvdzjVuJVHIMWLF9Iw+heszQPMcyfKDTHYbvEHuhkvqC142D8cQBEVN6TQOuDSql
j3EGZdIM3foiF2+BFRwy3JDe5SoQmhzqBvD3wtv5DlH/E+UcEDLxzvBGz/cgrPH6NiKBZi2W0XmR
caBdFQRwnO8a1Lr59qvBgdjFh+SB4w3orE+ot0rd4e+MJFFOXB/2hIURK9yZf1PA+jJIbc70bItn
24EFSkHeIMi+1WipfjNybfualphp3ZHj3v+cZiuBN5Rk3t3EJcNxlJ/LV2VW5y61UXk7/FK5GDCW
Hujb6yG1WaOCAOZ3hO5jSFzyQx0IedREpwoBQOOdZbj2V7+Ey06nyJpk69gohl1BzOszAzLdDi+b
8wVXpCidB3KhR/NI/Y0ebYc0B1dL5tmxS6BaUfObjw39G6xLeSePD/z/kkdz4352Co82FRGB5Y+/
BZqWN0i8dS6wCSiIx4rdC98aZVEz1EEJxse99Ak3wMBt7U74r6BTojRa9STCGQk073QloYfkPDNU
SeEgA4NV+JPvT5meZOSjZgrW6BEFRHgwK93YR9VnGHjcOaTpGlN3qvILiFnA+AKcAdcVLUvXTZCH
KQiifmJIcndVX0kagf0ywfIvhc77R3yW7gfpi0ZTnLtDhztNu1X+Q1Rw7JKEypsaBVwBl6x5Thqz
W95Ouq7H6G7EmqjS4qgiwKGFtENDtlAkpqB3IZyqntfbRncSTR7RghEr53gubwfzyQlc3wZxBiKp
CfiaRTBxsjZoZx+gkV6ufcgDvjyC23cTwZHe0H3dPoKAq5agRWqNvMvss/3Ao+7+VT6JCT9LeL7b
NB4w6msuKpLQcDF8vOXB1x2R1HKj9m7GxYOOcvxalq0NQeJcsp/JoY5lJ4Ern4dVovucfHmOgxZ/
UTSTkrFlds3qz6Ky4jCoBIozpOeXi6D/rszaUIcwyEYSna2xueyq/RDHZjrWMUWpmPLf9mZLkq9R
w+yevaTd4nt9Ldu7usMHu4Thv3VpaECwqqwTVohYrog5jKUrn+Qibiyu7o3YrOvKXCuYwHgCNUEc
1X5r/lChk4V6TqYp17sknYIIVSPN/8mXcqSrG8viXjFLH9hAngQC9yD7eq7WUAJfifmotyl6e8i7
NtG0nivzPvoQ1sXpi/CmaOTa9DvAKuy222E5Ky71sIyFZGAQ1KfE2p2MO8+9yXvqS3VpkEFg+7z5
ahSmmj8bZm98i80ceLqOdkzwZ1HD9xhX2ywHdnid3YQPm8CLa37SsV52+H3MnPlmiWXvDKmm5OWt
gDgT1umOrdt93WSTuY+cyn9+n6hKSdsWMQXZ/zeTeAt9YRSod0V3JBcE4peLNpbUc30qvgE4cFQH
+YkeroFSo3PZelgYcM02ueOPTUvm4wIDazWHuIFFbr7erFeeLOmuEms8AOWdgvc48EDBQZsT3Con
6OBMiLTgfohPhNL3fq0iRIKUcSOKcsEFyenqRnMMWnp/Yn7mpuZGWEp/WIXAdblcviuQQKG6SyK0
vK0dYTJa5lHbev6X5hK2XCbn4f/9wIRNyWMmBewLX8ApoBDgxJlVsi3VNvVVxm2OIFIGxjmOhbd1
i8U6ruq+He1xYqI3sUFFk4Vw1gHzfAOmg6XpFYZN32A2+YubCh5rZhqpqyhmPoxJE4Qm5ZiM6+cA
Ac0FeYWe5m6ffSTNqvHwiT1ksBxO0XrAXxIFxYxp3zci2uBMubOJMHeFdNG6tNV0CA2IFr14Gnrm
DqcwKN2H77T8gFNRDefo2NP+4eIroeRM1Q9wAX9LzJMf6V68Ny2E042a5SUBS9iC6VzUH9dN79ZO
DcN06YO+Dii8f5pf6by7jhmk9cJmab5m5cwBx3VRoBMYVBlJCIJJQ9WvsrNyLBtZ9n3mfj1UB7Re
9eaFlsYZp2RhzGlE4yWvvY6GwU4/6QcYslax8YJsjpV4Wyy3yEiy5Wk34g1F7I5Sgju9jK93NQI4
3VFzKeQF48n9FOGmIooCRmdYMiy0APLd+hq75gvRpUBN+VTjE+kkkwq5KW1kVakxZcVZR4tgQT8t
NF2qYHzcxLGFZygpIQy4vhdX20AXHoo39PVvrHkFN+AzLvMLAu0LwH3YVj0u9rxmtv86UrF5OGWI
GpzJKOjLjfMUCl6iifNYoLeOL7kA06pTBqcxA2EoVupg066gRWduwB2RTEAFQn7ImA/OF5g7oVpO
iw5dFQLXc8+zrTpzIdKwSQy5hfEkW/zxvb0U4XZpoUNPkRYE9jVscMVyv2yyAPhW5Dk7/0X9CmEP
lrQe5k+ve2BfRI6DLhJ71TNg+9WRoK2siz/1ilSjLGh26R/P55zY0FUS+Udteyhj3knxnTLn1QrL
9yCoeoAAxLqZif3c2CFjWia3Za5EHm6Equ3A4lsQ6kzSTpQ80Ue+wPGUltiNMIuOipzg4WAr5xBO
6A2nv+PW0VuHMPs8Xqn5pkqQIFznvbr8ky4mqa79VczRXF7N35sKSEe+Poq92diHpoqiNd2vKKdL
TruDD0cT4eSjw3PAQBxTESz0JK7yGDkNe7U/jLKTzJn9QM9HZyVvPGyLuqb9J3TmO56qw2Pf7qj1
ipAJiCCIA7hjWMXNjs+iN5yebf2OW/cZVStCtpNziCEHV9ECeuauSoRcRAcM6nJbdfxrFDxziupV
wV2izJ9pOiLt7rWaQP34kmT67BWWkuFSBETDUbVXzzG0fDaJzS59ow2A1p4iCZqq5Q8wtaKNrscj
vylnTskmL0lTJGrEULkfD9b9VFnMHrk9mLmReBHmaA2zLDrt9LfDSFFtfCLIBXXDdHf6ddZ48nXJ
bcrTWi5TehORUPzTZam25LNJPs7Egw9f0uE9TYHYPIEzopZGNG28Dk5VbLTODAsXj6CkqhGq1CoN
hGoemCFLTGUUoclNu8kQ2HjerZMetyZ0ePft1ov2HGC/wfPrbLHvW8l0bZNu/+ymu0Y5pOidDdsr
AKSwpJ8A+m2YinNbzSu1EAb6T8WCqIVPMujr9ct/yr8jGks9IxLOduvZs7vb8psr8hJhmXBdIQIQ
PGQpxafUOrvJ6+1XVitklM/PCnsdW55q3baCToet9/hh5mCCA1DJsTZY+5JUa2U6fwdzu7xCEIn3
8BWapAqhylC+9weIQoTDTBufYAg3SZ/1ZqPE2zXfMqTcg/jt5a8zOjKNj0Km+WNL6y14Ems+05cY
jOJdyNU27nlZeIOjlI/+G+e0tR9vMXXFoqVNFgjUYqfv610Fj72vtVb17/FSb5cFBrIEmDU88K4M
aOeO0HrsXtlNDmAn8m4F6DkyEMBCidhQLPeGABwVXG1nJur8LHkziqEQCUIvNN62b8Q6lKJDph4p
sUQ4vJfhACSKV0K9XjOxg5N9pg+2qVsPXu1kYpot9OrNl4jwsSEisSV+sVywhY2MAJTD6P+Q/phE
ETiWFpX8Hg3N6/mL1DABWnm+QrYXtWW6ULk1ILY++viNQnCgKdg5yeDyKHM6dlxyhYptVqePvS5a
06Xp+fAXlB7cu4J0bFZjWaqWUbd8G6E2K5gnywx5GSYp92XvYtWvO1zN62JlfB1PkrtfbjGwD7TO
MczSv6WVzAwOms0j2F0d5TT9nA6xafs/d3UpjsgudMD/sfKv2e+SF5VaQudNV1Pn7Bfq0+gIHNWT
OsUETsfPdUzx3qSBzEHoGP8FakIcDx/I9osTEkHDlSb6tDRGF//WpjY6CQmxQAL7vxfdd9jSQnQ1
td+FZ0Xt15WX73TbeRJUizlp+eaXcMMHdk9J1gfKjO/IyQPAqid6Q3t0e1Z0nRl2KYQxSvfPa75H
PjAq3Wo4OKwvnBNHbpnHHJ0bwa5Qf8YngFi1Xpk7H0o09V69Ionga7lyMrwnyrJCMBTOFjKyYgbZ
GqIWRUrtwCyaY/BrK+LokZjmVPTCYlRG5wDyZyuFC8IyIL9dsjXFSxmnmMfLYrucqwA70+eAuqJV
WXKts1o2Zx0ypM/oQWS4id6NHGmgCwJ9BIGwiU3rXsPpTGhVtKMHRhpa8G/CU/vhmuDNri7xNLlN
OY9sNMMCcY3ZVZSKF3wVhvGHyOJf4nFCNw7w7yVHbbhpxCLNL9j8RAEI7PF6T5miVqx/GFOx3/ZT
fAq8uWJZFFyrr2T27E4OQpwcYZIEAxijhafGOddMdzhzqIip/7jfPyiTufDOlEtMVHgcIucHdEw7
e+0FhR1M6pSmY8wMYVVGHSE0Mbs0I0XI3fdK6bGQp4A0Px1zRBEEw+ivgXGl4tVXq4hd62kfP5Zb
de1VlnQ9NYphuCmDdaRHvPPxFRcFm/P57p1yofzdVfWbyOm4rsZfzMsV/UmuWK0HCTSngoublZxH
Nc4pQ2+LBo3QWLD6ucgXIIYKlkV9vKHjAY42eaRBrRKqoN+NLwe6xwVtda1kzqPDxiR3ynYYlt7C
an0K0QbsVYtZwrB9WvKbB7dNe17PG1ONmSLJ9pzXV0wFnECSVzza1luXbn9lDCB6eSFEHJq17NIY
RHPCvFjr59U1Pss2s1AUFAJFR6kHnZAt6E4V/7BYE+f64f/OSvX2mT9izOgiiwExB7V8isDnje6f
Czcn8nb0eqtMzuh8C+ILxS1dCHh012sPDAqIIjef96KnPSa1Do4Qt2L8LsFbsktt4lE6thlknrvv
EtjYJ1jNNnANKFYln3MVO15HqugWBQE8PfNnDS9af2p/09KI7rY3W97gTXeZ0/gOymBQavLZCuQi
PWms7YhFsWZRCpyi+UH1fa3u1Ru5qSThZ6jM4xcYVnQWpeUcjekuBZAnEmr/PFwUJJFC0nLAs1Zh
FDZKF6E9NsL+H9wQZqC+KSE5e0CQWjdfNLDdRa6iGj0zWrC055TtrdNoeDPe7MqrCdX/116+p7Et
aUsNftcQaKXfiLqMHYLkFLO+19mMZEj8c8CiNoNTBvP27/68qt7CgjWvv1fg+gwKeDk2ZMfiAUJi
/oFe1G4p9wuwHLwBMeueZjFJRq3H57UvA58vIRJ/dApUoCY00XNhLf8ZFZnWNUunChfBIfhcjhjh
+S6s5hzX4tNpp0+h2jt6Zke110LZR5b4pk4lLTKXXaFqAd+Hp6HwShysSAHn3jvs/+FPknktKdAW
Qv5vHEJ7BL+i/R/c/5czwWHKCmPtBAnhgkR41xBNNuLkhwDdUmRP4e/r6ZFMsfypTObBM22frtFQ
a7RftnoEGMxlw4E0v6xfzUP2pWq3PQzcriZu+B9kx+O7Sp9fMxDwgFy1IWJhvnp6BYDD5byM6kf2
R2BIjPw/0cG8344Zl2O4ct32+35vFUJl2UV00ALQ+VXJgEna4/LAg2Y99wdp99DcBYEUD5imkYRT
gJzHnsfqJY6CkEjWCK6ArU6m8rQC0NFJADpt61oEQFOqa8fNFPAvPgl1D+BGH/ic0JwiXB/9IrQJ
sLDd++uGqllwtPrPSG8n2ocK7QF0KQEYS5zG9rs509MbySXD3H6MZElHJmv4ApFWV0pb4w/AYvVu
TBw2beY01Rv6Cte1FReakP1M5WS6mdFN3oSIH+SH7QZn+6nrBCMTZ9gL5fPR6Ie1Jw5iwYKg9wNb
tgp/BQ/i7CAovH7p5ArOC2sPE53PGVRSClKOj5F2miP3dqbuFvK6xRl9zC1gUxCZO1f2fJyrtt65
UxTFZoVMmNP2FCbieF9yKrgfrdWBNzW+5dr9ApNtpgzb3IFLtT+pDOF1+82BQUPysAnYFYs096Xy
n4MrAIGZCKJmlLM07XeDuHAfa3AwH/F50fSdXcVD0n3sJ4xEbzK5757N6jfYCkXG8MAGuoMHkig4
uc7P1J3TEp7IhtgQMFkUvIXP4LyLLTTtDB3gc/G+ilxjLNHBygl3KigJDYeJHIquQ+9ctade0Ofi
d6gEG38lZ2b8gGWwoxgEtm/doWRt7WJIQEB4zEMyL5tKlXM9+cKWeFzpUf11p7N5PXmLbnNlmKhH
BnhTDQj1GouPHY6nhmPq03x6rBW79xrOSkodujGduvA1+xXNw5CiGMxdEivFWoRBMnVHpaf1hpI9
o+4u5jBhvTltXxkErMPp4HzfkHOdGpB6FkmAFLv2wYTwSwCnh5MeGNGDrAKFCrvodqL6sAEAU+mG
phxtdfxCGdmng1VK1UC+ay0KFYzUOmNUdvsMxyWcPgB4XDUtUCWeL0u7O11p6i1gNLc5pub5xseI
en2m+0mR/FQPE6ANsO07HGOzXfvknu87HmYEDWUI/zpf0okj6j0g+kTnCrpcLFcw3wR9sMY4eT05
4n7MOq+54HEGDaXi89CHoZRtXRTQyhf3ZFsgosNurYi33n0mELMkh6FUDG0jPOOf32uUeI36cq2Y
YpKPkPWydG97xKg20Lu0EZc0GelQ4zhi5Tsc/F4zPup/c27P+Fcdou4pCIj1/DBycfpB2mURLriz
zl4Yrm5ChJHz0N7Qsm15XrgoelPriGkRi3NZPnTemUmdvXgzvrFuYZPoHAAThfMbr/BLtIOBkkfJ
idE4V8LT9vZKkWAqTtzMgVXIpReEDynNa0l2VVkuxvntVldV9QmZSWbCE1Q8AxUtH8SD7egAcYU+
UQFoYCbC+pZQPXMuE0yYSc898700p0a6UjtP7f1ceafZWU2HPmYbjND2GU+CM0nr+OyTFtACQqQW
hNVU2aNUdwniqHHmQGeERjHwbPLP7MjLbNSLuTZ3mL8HVZNnzlHyPX9lCgBvLOSBheh0iS2McPKL
87I3rTtROSpYFl/+8rA0rfVZsXbdlIxajsMmhn+oOUUlxKbo+nO4ja/JgoWG1Vh5CIFxeuHUy/Ol
KNptdIml9+ZycGmvplq5X9/TiI3B4DlrovWsc4KRjHZs/mExV3d4yY1doEU6q8IaddA8IWPyTvO3
8+mhFZySio5eRc09aMRZJyWl2WFUbh9YqXzKE4RTmA1C1r0eUOF1YGnyRMP+NpcdOLLJCQ6kPMxF
kyes4nmLeCo7ep6PanBjs4WpdjhUDW1hRFvnWKncu95NyS2OkXxzyMDaVKZRE/bFTByszAdRSJbs
nf32Qn55FOja6xfWPp3feR5tOIQ3pCyONUdRbKup9PCdP0AmB0Wmkz9Hqd+LTVQN9YkM7Fcrmlv9
SIh9qjRrwyIrMzCzmEsNXn6NGhJqhmYXYuy6It0cIrnxhBeFJln9u7ZAjFMifSTLhMl25rXIMxqM
Acr5wYysRu1hpCy7/PdXTeRtlFwZ318LXX7+pivrWaJmkgbvi9XX5trilLtZn8jo0feClrc3wT+D
3L4lPF0Y5rA+bN/9PBXQ7brzJ+gMIDDw0NoY6/WexA85xjaRYW+ks3pgk0ESgHRxQ6+TzWfvtwAa
ozlh5LRn7+5XP/S5AHffDxoCLoYxGFeLnUql9uJKMy25H/t3rHQzG/HPiBCdLPZw/iVvnDEoOxf2
/LkRXdFA0Gb6U8IJ6J4hhwi5Zyz3ph/ta3nw9HJyTJs4kCeDA9gCh7cMQ9JgLNlWBZzS18wSI8xG
MT5I6vJoEMYoWgkk3phmEQIivplz0T5UtGd92040AGFh7666OiWkrjvgKJEoSMYAoIlv6Oew1LiL
15QY9h+EoXUOt5l1P17FA5imzpjjiSqgd/ZEFgRClu3PPLOdcccms2rJHqPO6dzr/T9rnO3HT8cp
Mgu54cc39Os7YCRZITb/dKuNJIjjFdbwPABsvqZrjOxVVmSV9T+EODK1feDJ48Ens5ODSjjSdoVN
L59AipHRXNMRrYeWtuPXsoIbYoSe18tOZzZxY+7W9hlzYjpZWx3saHSA6scAAI/wyKbIS+O+lmdG
hiIfF6S9KbZA3/blwLigmipCJmmLSqN7ABfk5KX8j+qMHa4n6q9XGpB+XHK4SywiAtPMv7XM/BNU
lExQ1abgpSz6ztRGQ2OnGLsfWySsRmgb7u6Xc0ndsNFFOM1lG7DanWvX2qFW/qKv7U4s+Bwoo6ZW
M6oy9DmFcZpSM+aF+Qkg2bL4IUvlI1IbLfI+Xun4TNoZzCvrTvZohkaA4yl9GPvJ5qJWmFSTcgmV
JdDc/snGb+ZTxT4f7368lCWlywz7ek4hbO/5FlFfRNHiIsrd+KNStLzgl2STU8dCE5ZPDtbTNmMo
/BniO5VGblV1dns0vn5MnxloXiWxWMVkNpADbxremOxWO702OHVswGgSqftBV/2HdNNnqEupzF2H
7UxDkSG6lf2uvcjhPH+jjqHNYXA1xRfFbRWWPHYmhTbUt3RhCoPj+8dKgXatR4yc+ctZ4taGe01Z
STzYNq4lNdYUjNR/dOLILu9SaHf7kVlz5qMcFdFAbiAKAzSJxyES8DFWAfNM7hKoFcdyhGyekQUN
t1x571CGEG2fANaRwA8dCcksnOO4xqlIiNeOCM4T4/r6ADRN27TuZWC7GJrVBTkkfFqd9Vj3NjyI
7RsePQ0bXI1U5c49FZB4Q3mX/3fmraxRBO9LID9TbIKW/jZB34AfzS4pi+1f+3JsrcjqC7XbZFf8
Tx1uRQPlz/MwKY39y0KdlVRlxq6ISYNuPuWz3SfYWkNpTI7P3FvCmu9XOJmXHcuJLUXSCqbDTfvx
pzrhmyRC56utVnt7EUFjQHXEsLhsNyL0J6j3ZYSrraOy0DVywsNPIt/LAN4zJJifKJ/97LD9C9g0
6j6uc58s53ZWSlrLe3hr6ZoGRIuVSBq6bgyO/bkWxH8wZBK0y9kiqWbz2izYdhD6Ic7Xo/yD1dCf
Na2s99uBLEE1Dch2Yb6U/ggjPstuxJOtW098adntxuBTmOJZ+H9ObDVghY1wLnfnSGm0SBR09M0d
FqLIkDu5zjKiIUsL8brV/EnHgnrsBa1nF9Y3YvqytKKn9UqFxsCp+nsQ0ZfSO3aLuC0fOker5anQ
wR4Mv1TNdQF/MFYGB/IiqyG67JmTtUrNK33G1Ip54LM9JtpbC+qmGBbSKwG1LF5F/Q1Mp+v/AVGp
9RzOMYzz2Z1DcoXIghtK/GwqvXUh73YRxzCRvxR3LvBfpH83DJaE+YySBqrlZu72C1PoD8l4vova
OpmTLpMNBjRto4tAejayudnaWE+1Tf7AeJkWa/9p3WLvdIFaKaY7qOxqq8+KqaVe+EHcluupzEKh
9tDLjYArevTklpG8gu/wj3LVR9GP3xQe6p16rev0tbaUEAJPz/vmZY9BKPm4FuRkwKnM7BDoW4u/
EMvw20i2JjdBMKpj7D7BCXPA57/D1pG+RmdioMAYuTNj5iB7q9jnGsFgJFWm2o9MdtZCCJs6nAlR
gWoJu/Sq61Un4Tq2vQUrz7RIerFOydjaXLIRx/c7f0PbEPXdBY6etC7bUtlkjUBkioo0W8n2tJQf
pGSxzrHoU4TBLK9a1mKitRFl6AMgERcs7chPurkHP26jC4N28N3sF0H/+JWKxwmbNwPJla35HYAq
ouy8mLDIMJC6ReObwy5LYdnK+Y6HOA7YNxJ4HfQnTJPECniKmtxGEkfZ0XnpOVrhM//BbEDTSIQl
cmL2u+RqWKp86+6wIyJJMJXXhK5HwVw4GlDgD8EdrgoS8EtCujdnjLGqkjBwVq2PQkdbpSiVvIIP
7t6XLNz7ZE5I20JLPBIEKdOVE45NHTIFbxB1fJvV26G1do8ypQrC6NqGfwPnFcQbrNXzO6kCRS9F
ReFDCl0rCEz7e1PxprxD2ZGqgXGw/RmBSDRc+Bs7PF4X0SoHPQp2EWPB3G2LQH1lhFuzKdq4//16
UQ6+IPuQ3hQ3VPHSK9RKFyWqkNPJbWOD2e1kmC6gi8equ2jXuzNlCdkONrARwENnAG1kthFrrF93
KrHym8VNaNlEOn9TS/sAA9E0JaAGTyhUvG6qLWkNi1rOA2F5+lXTx1axLtm7Mtcms92v9WCB4qwy
tP23KYI2n58Me2NSVxQYmRpenfMFUC5dN0lnSnJoMIgsiokAz26R747zpX1IFi/wgyuUitPjvbX7
R+2SRB3hpUlSNypQa8flhaM7wl4jQboQeQCKlf5ZLzCVGhmTSgOR9sM8D++lLegsy4PL9e7VQUgt
vNMv3KPdadXEzBf9DyGC/jKk5mSdti0LTfZgmr9sAW0QmXsWPeO27tD4a3O/aU+YYqtHkJa6sLcI
rFfEbMi/WCgM0GgOjbqohCTLyGUeisjB3pOTUbukL3MS7DolgzOOR+ZnKLGibmXuMo3tufBn7l++
qbg0DbW1m/uyobU7ggPYKTYmYzuiVwhjG40sPd8gJaj40gFWRIBc7RS4758TStKhb/Nkyf3fgyC4
g/cIoyKEmxd06K/7A+iFg8+lPgK6utLscZt+UhkExL1W10bpalVXWtDk5HpFl8xuLEfmSIJj50Zb
vfVkwHIgE5AJoJjb3ZYS9nOIGNYvOqMvGukJmc+Mdvgxx6agLJ5PlwcOK2MMXLchGB09tIs++i0S
Nb9lemA7IaX0jr/OxodhfDgD7HEp1GX9JzWnSxU3EXpmBkG1LOAaacUZhhndgFLc8z2J/Dr5yySJ
cf39Zoi+thO/miyNllh7oJCWr7XLBKgcfPMWwrkNHn4ebq1oTfyVsWvgyArVJOmuna30mzLi8wtZ
0OUlkMWvfdFmIrnF0AN+S90cyrCdsScUkghJMTG/WioriDipywyITIWa9K+8tGKJmqoYlayttR+v
g/qQU65Zj89jNfjLOlDDblGOhQPtmdPBG8w5O7lhC5K+bnu+SqclmsadJltYjCT9VKPY3G+wGH0z
snfWP2TVlm2cqvKzBe7kkcuZ0BvB/uOk0kIxte/U+GTZiJ5mhMQcBV9bZUgi4I+r6Xuvv5IsEYoS
gPNBqF/Aw2DEK6qH/8ZafH97JR7rQnEOtPNVB4o7vfeW+gEETqktkVlcMYDJ9Jqyj3e/tgxmpz+R
s7VSI+lny3pjaI9AS9knHgI6Dcj6JZXY9gYsJ0HzIvg2P/SBx5RJmzNbvfUqg4BY3e12s4Lkr1S4
y0vGdT2g1G4bRCkJahZi8aU4Hv+ydE4nHAqDrouxLTopgqhuh7j7Zk4ttGoAlR4xU8svkSl7I+z2
cHXIG3rxRIpm0qtAETEhm8WbF5Cb1C71j6fhH7/kSSceN45J3svQIgWN6sTiEP8lNjtUNwaXCcWE
4emwO/CMBFb6LRSs+2I8pHjRaXvJSYMwjiv/Q4t0Nzra7UeyEFWq9AwbocHZQphFIKMCCvMafJz/
7RN7c2flmUOzppkt8FuMX9I4v0eAcXiqk3tdge63A3Jjo+IHw34UnBI9a+FcI1MMVroV+d+k41gK
fcxsrkujvFeO31mr16HullwTPC+4b6BVhX0MZmbKNdiLGjYb9A/YCkSJmpDJhamd9eYyazm3NqjT
J5FWai7MKME7U8k2OQveP418Ygd1Tm2mNi7S+eZff899Dee8P0H65ZYgxjYQGaQ5Fx77UGnz0CrI
LH2KTj9Cz2Kvx8gow72Uy9phdmP+68WKJM1p0XMrtV6GpxbCXddXHx2ww4dvgqS4BHZ7RMCFM+tq
1OQDJq8imrV7NZHpoRB78MtEtKOJR5C+xEf+ineVEUYilcUj9pM8kSFu0Om9LA4a6O+zurdYV2wS
KQDcdN8Gf9JJCOioa0Ra5c9DH7rU3zuh0pQdjAB9DaLgxx5ZlK1hxXTPlvXhpsjsnhVhSVBMQhsR
/Zd64G569Dwx5CqV/GElOSl7HSiOSSbQZ1JMXcpzyHBwxVGvIOLloL9hwlTjIQPP6H6w/WTwBrsI
+JFHu+6D/3OeQ5QxHr09DddFQj0peVEWLXKHVS0W6tL+XrRx+RcWo1lR/PwYO2hXLYCtn4MJQXHt
2+b0oTKbLARngpznKuWZQVMFv7c0AzQ+QcXUq9CV9ThowtsciuorQlsKLUaGfox/sWoa8zfAQF5g
xNtTUnTXkVl4OaqXULqBTTmTCfWamXbmwxVc0/DjDGTqPC8B+7eD8MiBznLrPKkwuH4VOfoTsOf0
iyT+A2inS2QJDmV3jXjIet2WAvp971UP4ArqSHmmqHWK1UgvZ/dee3wGec17tYtOQ2x3RfKD7cz4
Nr6wR9dxC6UqRfT0A0xNWbASeYqPNOJBtOX0eT42IDokRSL06jQrWOU+vLBMBGhaldmrpoOOKJuA
SKD5IrpJeffTKchEVn7Zza6xMryhfkcPZHBxXxVWmSXUdP0z24YQKo1m+0CyQGnVu3WZrLn7td1I
esHn1Lzn7WyFb83Q111PIv5rpQ130CNiaoT4RpCG3KULg/7tkfY3INquj9UqaJ5+UE8wYH6R/0At
3Jsb84cHWwlPWEkr3+tk2YXQVGvhOtxY8PO3jDZl93SEvSFSLE+VMh2TfWS3/c1n1UC21Jivzcwz
fTdQvO8QXPvfRTGFNjJGYGjICtPEc4+s+vdHaVqnMYWwXWwZM93RMsWYYPfV7y5p3GDxM9lGLS7p
mPvGLcBwyiOApNkXnm+X6u8BVMv6WO2uZDK7s/BLxviaaoA0AzB3iEWem7A2utSZ8FKFH6PEq3gx
zysc4Zer9m/X2PAA9tEQ90LBDKsXDMx11bKiuEPcViodHcVEWrda3rbsUgBuLy05uCb0u7ZkZ7EP
i0dudYJ8qXEJoimrwfft0jsgRPTF+63N3H+pFrbK3IyAZWiuaD9xQioy2swE0cYrxAbMQxhbfGBX
0ywuBxyVPqBR5mM4TlqaxjxhRfm5u6QxfnIzgnp8LmPLqFBZRnx9UClRw71w72lZwcOv8oLpU5WN
ZkOR151/eXoaiQDyrn1UrUKriepuF17AHCDDh9mkYIDPzdXaYT4u0uSPSW1WQwIH36Iv0XJc+l2C
UDVMBQdq+II6OIEb9l77h8LdtBVPtc1lgxmQF7zz7JSi7HLsxjuEp32CcHs5c+yhabhXrPCz9/jZ
7PvvUp/40ERppjz5v0/gADoqoKVLJyb8yQGHZxq3ju9aS+uhuXEWJHFCS+5EkEFB1qUWBYKyHP2C
pydPz+sLKcYpAB3hEW7bLObF/RrxMQy2oiUHp8rnSJ14Esyoj+oJ/0wPHhF/OVwc7pU79nUjG1Ks
wW/SBeRbQV+zITD8lQ8KBwLMQ47iZ9tTOMC3ThwshOLzIINQuj7JgmMeThkGBCe3DDfZZQ/N0lKA
ws8Z0ryGHkOiW6pJHRitbfY0V1/B/LnNhLsQejDPwOSgKJP44iBDNM5vOdUs8CilE4dYh7Q7QUzC
o6U0aDvApofCJc14aGCi2ny3Js0Wwq/b5c1gwS283LcZeLm+Dqq6tWvEevzHvxhOnmNMXriX1936
G3sQ37fwW07usZMKBTd40nnBalj95yHiD6z7bVPjYltknnD/CkXjrF4LaBgTwXi1rXw+LwEbKzYR
qeIx3YrJap5L0jEq0XqUKa6mkQgozX6xxJyE+gH8O0mf8ar2+6Zoc5kLZTqoWSIMNhFlCPFEuV7B
kTyFIMbhnldyLudokiQiHf64TC4+FbCangMKAKMkc0s4jkLv8IXysvFIgSM+9fdn+26NhYbaMN/5
mlGcKSfaKxasAwZ2976+3MP49/ttGx4wJugYW3ZAxdKKU79lBiPu1ZMjZb4HJqTl1Rfdc30mp2K5
OPLomfbQEg559mgOMQ9Q+KZoTxs9pZKr8GJEyKmFIFVRSpv7crcAT7b0LumccXbOZAPjHhXF0isQ
2zDH7eo9aKJgI14WS8GFftPUVt35HXasj4ZjbJm/ra0EE4AuZ94Qa2mhZ9SfjGLQVubU79fQc+V1
7aWmPse8twLy2Y28Lz8/zWg6B71DojiWKfiSL0WQrwBoH8xSzyG5/aVlJegX0pcpkvstwCsiCVbh
CBUpk/5FoQ4E/5s9DQ6h3Km2QFEyxAA+OrEgx49EMzzxveW9syDqYljrz8q+eNkIaBIRqfrJsyeQ
IvrxaoAzCR2WLm7ZyBGto7Xl/6ZAfJB0zaUzj7IZXSmlxI2y+luns5dDJssTE/RytoOQa+wxkuFF
q3+2rmCELzMKmjQahp2WRjRQMT399S166tdoJFeLkzSGcY1Ix7aivf5Wys+1aLwkNAIvsWpHGQyN
uxU8LmM3HdYP8JUop2rlYyx635Ht6x7QJpr72sgO7VUOFQRdzkSWcsW0swzBmHR7BLolky+MIW74
paV8n/huAdJ4TmRG2Tq5fg37KnHwOp4rl3JLt8cazXRAILDbjQ90xAKpJP93uyoPIpsH2r7dVYJN
1fbCQ634oVscsaeuqbdg/gFLwxLdz9+a5suTLB+3HMrihA7Wv7g4/dEqQ7pg/SINX3FvTdmQdI6Y
oTVoDrI6WCSVjeHiOtH9nXwaw+EUml8ao7t8xYtXSYh0YCPRA3n4pPMIPun9DU11H2n/fE/Ktukf
ncpoEIRFppAN8zSA336z6+iq+VbzvagTZ0cyQeJ3Y8JIwzwcG00TraQsHrJ2jew2L9P55wlwGthl
ezzVxeT6XAORSBoCgXVi50Fp8NeJsYJdT74SRSFuzGUX5zPr+DPyV6OvjmiveoAyFdpozgjhksQv
LQ/RXJj5aHTFjjnCt1TaCxQmjshgy80A50hoGCjVgi5ckfyyDqsH/vUlRvs1aivD71kMvn+UM78e
eLt3jVBuDJddcUGeq/NUb/W0VTv0502SD4nPqUG5av5SI/90zUj8ZCoCJI/wGT4rmhPcb5bgiZQV
ozAD6vtZFdm5mL6SqDy9mOeH0GWKKVmcYUT4ksR3D/a/Z3UaA4xqlTCawDcdKZ+wcOvRiFSA5xwb
YCQlttNOUV/0wMAnDeq3q5m5mO8Yj4v4Dom0+DPI3i8fyaRFjRfp7Kcgq3/jBvGdA6/bF5mVnRoE
olwxWYvfL1cNK/8ePfZ0bXyT1kskt36H/tDxqXulFbR7hjj7diumWPlIb2cMkuVBVShoiJvydc/T
Qgt5IkDdTd/GuzaWoVV8GZjwPeq9/otq8eFut+g2jH7hREsTUFdKAUuGTca2RDbj795PgvD0CgjG
RpIuXDGh1thyUWrAMuMVJKtMNDO4EgFU4RmujWZfxTR0d5u0v3ImYBLmuj0o/Ozb+T6woODs0Xcs
oRDNXd9WyQ56sizfcBxsLUQrv0KRYUWDOWaO4z4alnsOQxUPm4OHUBl9fSfGjIuPqbPEEs8lKX2G
1Ohrie0o3eUQO6hY4BWIv8AsViAcLbseMNLrJmpgGguMm7/BnQMpfogaefQOEnUm7IOEGozjNyNp
n4BcqyPlYNsWBZ2s9/Gw6/Traxokv98LftLcowZ/EM30BCJvNI103X7aXf0eFb39qrtOPRhrROz7
0MOVBB7qa0I9BX2aUPKMAqlfcLz0OhBaPnnG8JOrYSEid678Nvg3+FHFOzKzu3X+HTCfMs0rmis/
pe66f1FS3mFXPj5Fp9Io8Hpde2DaPQA36sxxRgPH7NPe/VixWNDjrkWLVkp+v+ol5HOoJJG5nvhP
cZ4zAsnhHTiJ0wvBL5VPkFGsW1FRo1gbxhoReyE93x8IgG4tXVzVaxzx3EEV64/DlMKaE32IdtVi
1MhftUPs3cll/WPTMoR2QIjOiBxPCvg9HEQIeVKZUwZUV5L3Spb+OEaLRVJd5kMTzsmFSEJGdOF/
hQaKp44AYFrnvG4vbMAeXqI04b0TE297vfYE2FuBrIVf8wgGuTRyGuD/Q1ol6Ba9EEnuWkTPz6WI
aNhyZp8FVHi1obudsDzjt6bcevF6FE93tS2p/xbjOmo9CYapErJLX29RatyvT3l1AKu1s9e5nCrT
iC19U9ZjN0CfZ0uN3u9t886Cvc2882CEimUnZoyNczGDk/8VuqmGLNrRuKrzsPBNrbL6cPJp+amy
PEHya/mm9/Q4XUblj0NSc8IGiMERLzcy121g9pCHsUEVnYFKEBQ+8bHW1DY5J/0jlxm1ozuhIBip
k/90rCc3vlXnG37pt3E+QtC/URvNkTX3YKeiJwLdBtJAN9c92kQ3F1A0+HrDiAZKkId5oQkUq5+e
ncqi3ON/L58JCFyMpFC1fjrv4ct+iQOrwzVrDYhFesQ4jMlMX54XZh2MSh3hgLfMlu/X+8CvcFsi
RIOLFER5t8S1bYwQndFh25dow4Oq98IfvfPhy+MnWRFTNgNk6fWEcAUOr4AAVKutHDRgGBB1BV0c
L36TvATlLEMhej3xE06h0bzrMeHY0j1cMfq1/9tauT4hNvAEhTQwNRGOWM7OwlAr89ak/Sz1A/XG
cRJzcKJqu58qL0est+zhOJW560hUewLqXAfmzw50w1wlq/F5l6YCBiT5G+v6dMRfUpHCIQfJAoB8
0qU7TP+/1Z9Z4KcEC6kTyQG2GwEUbCkX9zkYc1Vkoh24eH2vY20o3aQqYPqPW+foTsm+kqLZlvKQ
v5MsIq1RsASGrpIl6lYYiPrMflZUHJq8zb4OmyxrSFK0L0wGU7lK5Ax5ba6BeRbi93QQypFEPz0s
JuMKphdye+rjAdY1jfQyrNX1SfOALlKOwbWaf9SiizjPT8RwL6nXVcXNy+VRxZQvtL29GyliBwCj
s3aMCLX4CPHU636gXRPhgGh8ev5JNfwu1qdi1JKm+jg+IdqYOgwkmx1DHVQpvO3+cPuEFnShq2FM
Fb6bFDdgDnHq7Uke2xzFFCU6Ki4sT5jLBYbKf/ZnxPd2J1UDS+5JHQxVqqcrBOyFyVGld+RtmNhs
pV6qDyCfG5Sd+q/lkKpOjiC2i1djaoe8kZKN5woHFa1Tl8pwD4ir1woUgkVaM3sncZqwm453yH2v
OmhfZ3aaIgpjF6rbd1Xr9YuZd9jPH3bVysSw4HI/MO1hBpFNdmPr/sEGcYO+DuE5uJuldehqX6kC
oAqObcBTptiPpa27vhDQ3xD6rjZiQ7ofvf6c2m9jt50Ld9G0lbS3rw0WHQeCRL4QWxeNJsaM5ZFL
TtDJHzmmETuTK/jBHv0N2UpsMJg1kRxXCEBkyi05Z1hhiNkhp5G7g6ZcOuJhMte1cPir0P9QzpZh
qwPVhvknRe6PwND9DKU+Sd9DyqNUrVVmuB/En5lB6G5v67hv963UngOFIW3Z+I3vMsJ6/rlu3GQG
5Jb26H1VXRGzW6AZicyuX+Tcp1PFakRasmVAHIA2JmEqirKRxllvEj4mfGo9RVRSiBI6KHo1a4/Z
Bwhjycare5CvreaFlBd5l/uBLcOlYeh51+/uTOf8rawNj2+tX4V0JWlhAAOVBy5xUkZFZW4HpHmH
hxhQjM7kokvzMqnX5m+l0CyF33cAmAe69yjObizsOJuniYzsE7uwENE0D4cYDkddusxoakvbXeL5
uv4YivIYVnZtvX2U8gD+6Sk71Rjg2j/+0B0LABdikB+XgOrGdY7TX2Xy7dp2FagwfiGYAkqjAI9D
7IOQq41p+OOBlHVTM9ct4Xe21f0xDTxjJjUvicWLKOGZxwsVtjd22hUPL7Tsogoub5uBXVccbCZu
MrD0/S23R4pKmLLHuoF6ypxapHwORpC2txB5wJsnGdeP7E6kGGrGSzG+llderTQHBipskWx1oxjA
8yvNoVar7vwYp7j4IcCmc9uf0FyXveAz8ZkaCBohZfuaSk+sSiKsV+Rgxyd+b+LWflhMzz3QZUQ4
83c1iPlnRi8BBDq/E1tLmJYIIyUpmXsgbt6WuhBrKz956+TEp5WPZKu2i/c9ufe1wFaZyAp60rhF
KIc1w9gKWFTSJqDRLi5DWb6fiL74YuG2+VI5N+Lsho9BTvIxJH7zT2k4rgJ44sx6zokcTTnDhEch
uMILqmcm3GoDTD/wnMSquS3fVBshW4y3w6mbfrC54uK7WuZezQWvCfnW/govZxPPGDc0MBN3Cjgz
VBHWljJT3HPcS6yQNqyrMCgYEp25bcMDSc0Jd3Pypu6WWWVLNjpcEozma3XJQw44Yoelp3r0ZkCL
htlHCIv5Gqa6nl6MtEeaNwLryy1ZOpjj/A5BQgr3UNP6wjl7LgXsiafAvAVZS5m4DQrQTZeyzqTz
XdR+BrTpm5IwohG1o2nxXd6HnVj1a7Zak+iPMU/UoA5kO2ADfwdpoxfhQEAwhOCWOs4nwEO3tWZX
1h/0jvhDOCPAgSUn4dkNtbtR9fAzCdVkOB7pU3JGZ0zy4KPAe0CPvymp47DAPmOiLVbv6fGTd4hF
gdZHCV0OU1eY+LtOwSug99Rf9/dopg4VAfeg9aJqVfHsM00BjZ5z4jza/Yz54OKSGIWSYX+tStdo
nK26Az8TEyHez5LLt0LHukE1XIlyzWeWCXfjY8EGqlVbjg2kiHoRZj+F4qgjvKtJa79KToq26qk5
615cq6opyP3F6e3SCW1HrtSIMU7Nti5C1TWuErfOZbkrFyyOrUYSgHTxWmHUj+d3PlzWyffI4TQt
b3DA1C77qGXj6No0FcQhphGP48VZ6+INTrJkbei31Fje0W+Wzxz4AomIuNnHcZ9f3YDtAWxK1tqv
SNNLzzmmJtF3VtFe489j1Aji7ShFb+W607wH2B3HJFPSnxCCvX+DvXvze5M5HQu5CWU+6pOYs40d
mXj+NVoCUrxc4vJwQIqjtNFoI+Dot4WGy7EBWD0eb+nqX/gAPqdLF0IL9G+OVeeI4iFJno5QJZId
wRkBVmaakBuh38scmTTG34hft9qkAENyfG2WFaeM6Y3YhaQ5Yqo5f1drOUtPYAVjwvx30feze8/C
P7sfbPN3ramCsS47F8Q/hFMF29N2fG7tqZeTeRUjDAMX7L/X10r/cH5EWXI9TLBdrQqM9i/4doR2
251rS0ZKKRbNbXhhjUH6mJQ1U8VJaLnjbJPI3aRol2ypkh9sOiXxTGu1FDNBUNVv3Cl4FFzovhhS
Spdg1kBHTeCH+4ljJlscZuTR/98gnKqujsISoJv3iOTzoq55tkUxC5vWmbonDiYfoobm1sg/iS1B
TOZsuQH2Vs2Lmmu57deakoRv+b7ZSoUDlvxdxzd7oIUMXUWsqYc1FXdRVOHV09B2iXwB1uRmXuoP
MdmbeTC5J9dgCMA2Re0DScXnf8bDq8PjeHp4+0Jh5YKJ8DeTmNlEifXgivjVMHrjrW+ezgg95LWc
f5W2QfWzSUf2GWDc3t69dKuCLMwmd3FOkaVYUz1lpWVbTPr0y91RXRUuLCZK1MtMg0uuzg+YKJxv
2ntLuHCLXbKZdgKJAi+g8JRn0p4JVcPcLHHsdnLd3hD6BtMtvGzpRu7Sl0zkGdAkoZQ0rO5MRoWq
cR5thxmKhGiKn+suSD58GrgBQzVf1UAXsKX4iYu3Kz6gmDGYa6+Kpw3+/Xbjm3ar+cG+tCSjJaLm
XCOpF2VB0OMDrFsZ8z/U2DwzILQMAzvssvRM5MBR6gcHAFlEk7NMu69E46PcCSU1qS+5FR+HCa/J
ChZsy6kQY1jYAA/O8MM9Lz0C4tlL8BJ57VWUUrdeVsELfjkhjwyKL1T0eJOO5z4nhR0HlNxzxNTa
YSlP0jXz6GCEP+oXPRjTkjMAPwktZWMZaBf8koucg62Y3QpUFcZx61N6aALp6KahrkX30+b/S/3J
Yys//YBiZvSQ4DebiKHlcVpDv7MAhp563I09N4C2JL0Aw6LxhYOJPh6d9YK0YPYxo58aBXBpl5Ah
B24+n/Hz7I3UqMOiFhZTMcN5HX668OK3HAqjvIYezrVnDca9tQn8ZonFzWPwymfZq3+TJCtAnbUY
5D+IX1cqQ2dgaHJAPnaMrqxZp2RaWXJW5JQUEZk+NWU0jO903IQ10XGb/shU5h1apbbAlNbqZVDF
/vx/zuDVMSp6Qki8pzuEgqwJU466pkQPv52LlUbiKusY11LEAELoic1L3Lk2sAtRTqzMcORCbBRU
+4GzjoZT+on+vfwy95R9h4IPdakQObFE1qmegkq9YkW7ubYfIJVUtm07O4ZLfXRqEYbWYolEOVxW
m7uwh0aWcv/gZq8IWvHLh2pAmVFAUOT6Ogje36YYih5t/rP28OlaAIPJtJOcbnRjFxWfg31K8w4L
BcMSh0pAyjhHR+AZVpJ2sjXzsBh9c9YsvYI9ek5sg7ApvjEVblivHy/vvIgF3TwZPa2mkaliIIzh
BqepXCj3SLWLTVMzcUjN+WsXoyIYW/U5z5pBIuayZGqT9vHiCEL71rL/uxwTq/6rQOebPdLqy7dZ
iYuyrUCTV8nXi1XKtYBQmeiQ4YCndALIwJ9hKl/M3H6nsaw3mGdPgD/bYMsFZFYqwg3jDyI+17ud
rHQcil6BdndGRsi0EyQiyGEafLPgRJIs52sWvdKbF5o2qyo/Jd5K/FE7RhIyahfoXJJSfGVarLsI
YANB7P/o7aXYYpHvKlB3HePOMp66A3W1crEiqDx2T8WLBI/KrzkZF/rnY8KJWr/xd+EuwyvHr6Zi
UwciEiWVYmCXRQbLrPfHW1bcDB7euYC9PyVwHthooy8pDsRPDNh9n46id1H/DPiFM8QnY6qo14FL
7s5ud295cjSkAOIRsga3qw1Og/OvpWc3n7MLUlYNt4SNDSv9zO2jkFKXqwkOdUsDjnctQ+I4uyQI
j71oRx2lcz7r5ht/JEZNqzJZur1al+l+udiv8qbM/miII0wL95OqbBbtf3L5ELf81YxqKMvI0rTl
BKcZyzE1uSQUYmSun+1fUlAVz6I9I+f5l6LgdyDUTzhkpUIrshKiSMO1h8FYT622WADA9MzDDGPu
KOKVDohtWo9XKl7ugTj5thdAoSq0L/z7Z0QErjVUIQKcPfWdzDXzqYkoUN0BkiMSWSz1hk7zTIjE
21S4MTeQiyUSv08hGUGEF/jqO6KHYQHNzf4wpeJwobFqH6/vpCqgu7GMmBL23Aiwj3IaHNhvT7lN
1E4OCZj4IW53iwz0VkPKT9HYBp1voB7ydPayJgfA3YZA+8hP/VsZ2d/hhXy1X4i0kAmi+xHn5NMD
OmCojLNjSkB9eSsDPumryrbNM2p8cHNzolbmDsSPOgogHHJ61hUzwN9KiY6PZLYTgmWoPPzGtNGq
3ymGAziyJgbSOSYXJ8efjNKw7SwI7jz3let8EJtgcMyosPJ8cHF35qSUGhjbKGH9qMLmA+ToR0gi
Y2C/qRzsS4ZFO3jDWUCaaIYP1Z3It6qk/72IYMN5XYEq4/+FtwMpIOx9w7Ki1LK30Df7ELDwc1P5
2d8MHDVHenRQebP/s4RgKvz1JWzpm+bsNtHPXxPDpmbrCDV0nXHu9/fUjzshtzoRPdvNmPNUqVqe
7K9nC/YbQDPgqf4ROovF0MNw31KFoMw72WdZV48sy/DuHZ0K4sJ5MMVxvvBh2BG0PNBqn7MbhtCT
p4DySUQHohbVujY01iKIzM/GFvVM7uTLVfeGrokzAugfwgdSWtOzmH908ZFGOb35T/m9hozH3kZE
bS/FWA3HQRkcuwhgW6IhVTDWSWVbL1XVzAAK2EpdXQUz1RPHzJvb9fSD4EwDtfFKdQst6aW0Vf6g
gW98i5IKJpwMxTnKt1xxq048+X4kauXoP4/YYkDuBtKBx2NvxJud5XyLCtGtvS+kre3gy3NjkbzM
lSf8z36kdtWi2JXVeJhy60GuBF5x9eZHO+ukMCG9axxIGePi4rFRgeX3fWJI0Jtn4VUQhqBylm9Y
UcPqYYfstviFgQyQ3NhAyyzuT4WfPfauOQychgLcFsxWH9J/R3gTfiCPxYSmnYKqBBkloyfrXCJA
RcBEQuF7fpCR7vXFERqhf2eGLi/P2ZzSUbKkAlZkN/gRIU/G15Z2zpsWnC0VfOwLcI73rew+y5xC
JMOXRWS5L5aHQ2ngSCFsZ8MxyuPPVnwdB4jGmYOG/8H28VWEQ+hO4LAX/PtklH24Uj2dL81MQPmN
zJxiLY6OD14SW0IGSTVUv3yKttYOLRgmigB3FwKVjReHee5tFohS/v9wGEvAkzn6OfK/HBDRDI6T
qf+lhVYei9Hq5Q8+8pagsiJ9B56OFTLO2QraJnojZZOn1n1wsdXxLwPezoLDT1Nl1yVK01LOH9MS
WoqEcKTD4s7+580aOJ3FPmYaQVl6CR47ReN77naycrRPEeU8yMtBkJqeK/GlWafVpuX4867Kt4ci
LBNFE9IcD5R9Kf7qR3hCqJn/9hGtAjuzzh+qGdLuNqCvsS3aPutlOcmm3+qvhpnSJM7RhxhY4+IZ
4x6nh+2beLkN0xWIBcGhmuqo0de/5tR1BlbUa4lqCSI5SPUb6QOgqUdagKXTk2kM+dTt8uu6Sbsd
PolBDp9MQLdnB8BxFBF/w4FXuWtAwvc0hTXXjB1Au/WHqLc8r5oh1gyXXKDKocM+rfDjFip0O1SM
BjiLo75BJXukbeLkO6lvbJGKJ8EIkb9hb/NC9HIJUHsAz06qBkiBVqXAU0+SKUG2ierxOAAxRSmd
XS10sEiOyKUNHIFhrF5sHaew3DL4MMjGYxu21Xx3XWL17Z6YlNoNwypggpVGZe+F/Ki09s4MXLgb
Ru90wyEuCzJiyRR0wJIBTrtziT1Md5p7uohHy4Weaw3Muc/RlpKhEJB9ALIbiHnq4Nd3FI3yojTZ
QEovnZt3WeJr7WmMuVKGWaYjpRpBDG4Bxry6spsRnKCRLVmDx2RT+0BvW1GOJ22b64EI93UOuCsG
1FTgbZkmB05Qst+StXajMdlxXZRjnH3HLtamOdZU7iYq44v2vkhZbrp8jfb717Ixv944L5SSEAoh
JCsBRhp3DL72b6yUdjy7FwsGHyF61Dj0wuE4b8CXjoWf1FwtPmtDboB0uI9J+jecgTfNpvksjkV6
Fc5Tveaj1ucKipBOuReL9VTpeTdyT5BUcMT2Sp9MGi2a9Ns3wSr51M5wduCnLvxh0GNuDvDJ3ISb
v6S/BiOUC5sZ+apS7DfybRb2JLJscsY2mETyUYHUQ1jegoyohL9QK8Ul1Qu/V70QCh7GGd52220w
/qxDpY+4vPyYljFNXnnwH8LXllaBsGKnFNtGRo2sd5rBrjMIa3MyIDRW3zf/e439yanUxDPXr8HH
LDYvSUvMm32zlo+sA6b/Ez8jG19ItOVmkqxYL52EZQ7feBgR/xcSs2TIdpZzjrSlVJBB/bk3Npaa
NTWadAWGKfvJH8Ep6okVs1W2gUlh0d4bXi0yU1liB88ugp6wcCuyGPT7pnK4O/wnmK2vWFjDAJS1
ZU3n1V8llRfHdYI+mhkJLQkWo09WDp6I4RhevtCMTqTyf63cj47Gf2QIWwFeL2Yf9o6kLw3lOkEY
ZasEDxue6oVRd0132ICkFqEH5enbx3FdsvOPaCmfXLFTdFuCOIM6bAvO0VYq61E5oOQADSjzjoO7
CF58fSqWKU3R1J6o4zK1DAH531TZzt0+7onJaOOcW2ioCe8j1wm94mHjsQzh6MhUtuBJSDShKI5q
h5rdbIJetqVYbGukCrFuhI/2EZUdI3/cBJ3JgrkjtuZiEeJhfAR2dsteGHyzqRCE1CHYDP2mKAnR
H9mRykmHhYtYic/o9GyEjWd7+bJE/6LOtueRCXPLKbsafMJvj2qljF0gYhgcXbSh69jgApU89n80
pkIasn+O+2m40BxXMvwUj+wanxPxkoNnM5vVkSrOR6cVzFhqUSd+0MmYjbLBiK08ykWK4oW32Qxy
Qxbit9Uw/e058NFOkvncTxEw11p5+QV8K09jkjd88leRQ1ONVQfum+SucdLKM7EjGU39z03O7mzj
Y1gIJGlhcp/Z8SBCegOGNtd7k8Igd+DAI8UHubKEvPyU8xHVqaXCeKp1Ehxpd2v6vq0ZBp84AGK4
OiJ5kMQ4VmSiFPUaV2W5MHeAj1Kx0NGdW3uZN/DoaHcSmpQMEUvc4wkmV6jVGrCSTjJvuzMgQSRt
hMrgbX/FGSGdRPLdYThtG3V5mxLBRyHx9kJtOwKmUItNSckE17XJAoA/85FhMffcn7rSOv4/9Hcj
Y6W/8cGZPk8OiIFxi+ANrf1rT1xE6mW6MXP7pCMi2J0o+sr/hcdqv2Qd8VsCridJbWpEF06n5UqE
AtL4sUEDBYGWpUSXrdyBTCPzSvinpJeM7NL5qkDKp3GaXNBspOPL2fmQeCIPav9gKgbsI+zMt+/Z
cGm6eposa4ZxXcjUAp0UCpYZ0/u40BWqbKK42kZgRQCHxTFGa8QfpT4Uup6FtGI10GEZMBblM+jQ
aaenQ9yPtguHOadl+e++MPKFXDbl41k7pVgCZDGAVn42PHGdT0vNvGgEOUsk2NG6faBucHRqATu7
1QBfBq3GIRX9ZwCkIeA4fAsG5bN7RhggarvRJRw1oLRJKK3+jQvAFlcAVHgGVoWwNMTM3RicqZtW
ZkiIehifFOqTHHBSYj+1OjVCgwsO/QiAKhprssX6NzO7MiLZshJf61FqWOauSe0WJA5DD70uo65q
eY76PK46kPcnLJutq+DFAgSTGXhwSS8AgIZGg/ZP/v8s5jEOoTYSEv3CHTOw7jBQw+f4Y4VtT+Lg
7juWhOjXTxBPbytq9zCCCnSsfrBH7o9bh8bMDSqcpMzyicLGYlYnVeBH0o5SXmNV9DZx8jZAmIgt
SwT/MjA7OjIfX15GBJiL1Y3hFrxLBlPxgBjsMhX+1lCElEHzNj4AgyGLKYNjoj0k2qDeOgfXJHeA
gOplMc6LSRSjf44d9PTXZmLyNG7WEr77DeVN7vv44BdIDH97bIg2lBoOJ0Ehv9Gvir6ZAH1gXiau
VIixGWMzZugBU1OwWjyfb8WyJPcfcedra+CS4lywyPk5FumJ+G/3Aw94VfA8auSehrpDI7B6uC8h
tC8KNbRrEtVjkjoyVAn++ZcJTFf3lq00W45AVmrtFv0Ihj27SIx7Fcqg1dM1Oe+O/j4qwK/5/sku
/Q2M2lb6ZFA892MfMLttf1tBB+udBh8v8B69P2pnSb7FB1eo4fhPM2vKT44dWo0QG/PlxkNYa2n+
qi5SCXQ0pChwbkZLVPXF+VUaNb8JfPMXvZO/V9Ecruj5X6nLg8gJTRMoo0kKha4zcj0phMnToqO9
6RwOB7XGFqXqhopNNu1q0SaptY69YzmrcjDdE1slLQe+iTmTfH+dYjpVcLBSD9fdP1XSrVrIS4rt
BLRsbtsZYdCvHEKacZ57C389mVEVf2mIl3buzRi0kSnjvs6jf54t0L+y2C1IrP6B43yUmXZuVn50
0hKT7pQbWI8zoV/Tb7dm2mMWBFQQn2MiqTNrvtHIkwAVy1dl6dDzam3p4uTJlC5DoNBIceFOKk7A
vcB+HCSbvC+LDRlbXyg3Mj0zGeyeBNQ8tezn8U+Td+WvNnzyPR7lMkRl/gyHNJwQmUbiSjOYBdS9
p4M6j9RRkijmV1zPaRWQYKYlYo5OSTicZEDCY6H8FBQXVFBDgxPsYnyT6YnTF/3sDMGE1rpsz089
MR3KG4wMQXoaKQ0c/rBXY9Lr0tLKoAu+GvIMI3GVuBNunQFxhj55gfu4Q6i4VoCbh3pyyCQ5YX1i
i90m7tZPC+pP11HPbxRmg23gzUgNw1BcVVFqPD6hO+xX2iX/IdZpJs80VuB81cNbk3empxUkz/Up
NdtZoCx3Xr7TGJ+OGPvQ+UGWhhmXzBn5F4K6G6a0AqTsjcgXtNcXLX1jFPA/FKcOQJXlPIrqRPDa
3h5NIEA7XvAdhK+Oj4pbAuJppQKWFitSAkPC6gcWjPNnz48k4RulF+vPr3M5u9zkZtUyINJLIr0i
MxEnemgYB9tgYJ71A3At0RHc5jl8MguYhahB+HaelnIZ0fI8hzEXDUISdnUZ7h9Qg1qMrrYWVtqo
rb/RMnyUzcAgxfwEdrP+p4UtHG14cfI4dUOi2FWMJTmAUsOo6Mf5VYauBjhGoHEipFsK8blE6WF9
I5zGzU15/m84elmF2Uuv74ltnx9hLwE5rCqLqOLnVbMdrcZv/sz3X6vO5Xvh/0bJW1VfqQqJ5vYI
b9XHGVxiVbxWyuBJNfdRPNjgHJ3f25pgnahMpW3DsRtPkidWhhR4fTxHncCzLf3QalVrmRRGNBsx
1tip+D1CpemujPRtWG9cBpidUsY195yhOpOkLPhQRpoXNy2Znt2RPNikkDCMkbtbk2LHWDr331WJ
Oxi6mjYHNJXI5tYWIDgqx0x3PI3WzoQsARdFOBDe9XG5w0gE9DTJWVMUcpG73qEC1AZNZGa+l3zo
RQX/3HGx0TukAHGSW7q3p3nfcUVzWZ4pDCpe/6YI2BKwcHdiB7aoF46ty2Itq2TQsXFDYU55w7Fv
P2+iVdFiBh2w4+iHVEppE03/ZmERFzprHEc2380ozCTPvnmrxKY5GGzk3fTdR8DvqJ9pkQbQykMr
XjXIYo81MQ1pT/kFNUcCd6aE5VQPhI6es4jLmn7pR+CdlFrAXJvYUiMx6RZ1xwpjU5IlZZou4v7w
NKbfocjlpQOIQE/JPl7LoPppk4XtoAEMryGvyFhX6ra5CrymnyZzUt9PS2nt1cqgxRPUKnkeDw0u
F8bI22G1zkZ1J2GNQclf4b+svh0YUyT3+83BTJNVBO4zXtEypbk/FITnw6hkiX9Q0qf2S2oTXTqc
27pDkUTC3zXDu4137d1XhjnqRlrJC0WsKddkRn93cO19q5CLukjwfJAP1DHR5Zh4tG+234wL0tpP
dZ+6nOZw03vQPp7O19mWg1B6AzutJNm7vC1gAMUmZ4VaG2F5wdYIo14cgCOgvF3+WlHpEyY38Wrv
F7lP4Yrh/YOFcZgsB0gjqk7k9I6DtRi4Af7AlXaPpbeL4+qOxOHzsuncfbnrQJQXxcaTbOS1wktr
1khlTMMcqofHPNZ2IeNSiE1TsEGpFOFaf4Se6LWT+ooGGYWhTH6EAeBW4MjXgCtTnMS/99vgEsHT
gWZuuQ9pZn/nisYb5PnNMkzY4kRikD8gDbT7dE82vWtRXd3m2BrLgWRU1L38eQelByN4d5l8kaHr
zEbbGL7ejel9oSIq8JnikeJ/prGDsXeo52EIIVCx/EipQAtsBcDVGGT/TEA6FqgAZ7nQXSN8l3rF
96IlC55DJVMWNvve8z85BQg5s18sEWeWtATiji+V6QTgzMwShU+TfNVx1sdakzYnnwGKRdIdxmq5
MF+ahcYCBpmRu/VHpjPXjj7HZgLMZUraEwjcelGeURv+Wlyu2F0FLi8e2gU2tpqF4OGAhQCknirv
KKyIbqntjk9v+7obeI6/3X4q4AlB62h80aRYhy40sB+5I+mhb79kfLrXNhcO14Qiy/JRYfYzuhVJ
iYnmWH54y72qHL19zUW8Rt7cVM98U0/jhDQ3HOzZcY5wI5LkGOA6brcrrDICSGwKUiCrkUE8M3aX
DCsXL0AnD114FLsHkdEm+7CWvG19B0FzVx+Z4YTSBu2TfN+R4/RNHQO8jPNAZFOC2jwNISB/bGeX
TltrgReKlAi6IrP3qMsUMMu+02cpdVnSpo21UIbP+L3FzEWd9dMC7zdbrmQtT/95bc+CeXW7MAaE
2t5jvtkJCMXDPgURNvad0HPZm86rHlDMJOUC56c7nrhuub1H7HYlrr9aAMIDc0b3BeHTvipSk9Qq
HAZKUIovJPIb2CwAg6FqNbseocRUXdL2xcS9qPncg14TWdK9Cj3moqvutmvGwphWs8gUMpRuk1K6
0qZoVV65/Jo2pZBVoimIIDmVqDd0nzzUYRzTKUd9dDdVPKzmicaSYORsd8y4US3TstduigIIOrkA
uaI9G2EOGQ5juiQtFY2Li00voEqAysIcehRNyhIH2+46mYNYk9Q68ALZPsuHC4lWaKRCEIaf9itb
pb6qoiqFG4oL8vce7QAGzUAZ7YlqMrpNr2MvQlD6jjxpnOYZZ4v+uINfWNrEcC5ElGdWGdFOM02I
6EjggxkR9RCIAm3GkKnbmlOtGp8jYAuN/g+HXtv9LODmf66Vhcv6SLkmMhkQvn6vdZXkXIN+t+Ts
teSeu9M83O+nMAD2PK53NhVV3AmQLa02tuWsYeoTVuHT3RlFMeiwWBuUUZI0AYwO9EbXSmIsEC6l
D0vYNNyiv7eM3yBzlrTFem4t6RYewzykHgIDCRcpf+o5vlZcq1MpN0o7K9aeY8F7+sUFgGifkmKc
NwjeVtIwjjGcQXITuG7tKfoTtQGY6BGq675H/OAHP5XKEaZ8acoxhWupBG3BdjH4chcy+qqNaCd6
lTlNJkyTKD1tsB7RfnccCrCaNMQ2jQbt4McWnsYjPNbyBiLuGQO5vK74L72+v7iob32c9ZSmwkQO
YFBXBcYrKekBc768fFpOfaA1+GUiQrskUsmPS+SLjkclRTQa/lffZv4qUxAap9argnTD2TqTK4Tl
pC8Eqm0udsS4zsHoAhdVBu3tg6nbtbwerZYOKWMT2mWrH0xT6sfxb6O22gFF02u9r6ydamHVRApU
ly2DNMFlvdJ6NXMJBxsaV6A3uQIWoP3Ic+rp2CR5qisFERlSwHj+ETqcGLF32t5lu1jgXkpxyIbN
K8jwNfNaE2J9VOQo8HydhX1M3/IuvtcaY79zbT/vRhBEM1LrYqCTAh7fslaBRslqWwA3V4nBs4X4
tXCixZj8MrIODMJGsWAkKO7yFMqikqyHx90Tez381g5TA8NCLDcLQmdJ2F+Oaemq1BQ5a25z0nwJ
FiV2WQYB+/mf9kkfzQEqYqGPgsB6ZYX5JL/zczGE07WWNRJeYkXI6HaeGwLWJLzfKtUKOiyZ9Da2
bM2iI4gayfca90fhtUcA/nEHOGDXFU1z5DaziTICHBMyBdE6XasJZ5dkVDMl7+79Q8+vahqUJ0Id
z/KxCznHer95DqJgrWzINR7MawEFSMUFwnZxQxcC1w518H2X2C+KhfK0uwcCjwfjcd6e52BwRqJi
hzmMTbxDeCid5QlfvXSgycRCn4McQK/BgApQnSqcGiuSZvL41nmRMbvwOlClSY2498yRXRp5f1r8
b7XpwDLT2vnjXvCjxCBg2P3uaiPZq8xePMSebtWsZ0fFs5RBd2yVU6aLLJrXagYWUp1E0VeNPVz7
CbZ5wAqSvIVzhnPrgv3Smaj8orfBZLo4pYbMgK7VSWySNZVNlo1gcJcuh81DhkKGijs7ScxR60N8
X+7trGqM4B9xL/bowPphG5EfE9cjLj+ZRGkERctIk7vAMkGhVMByK3AS/6lYuhWuBj6oQYEoVgpt
n6SAbAGbS2lXfm8J5RnsFIu6hLfOQI08yjgyWeNo9NJtXb3PF8i42X5JpM2LDEPTBuBoG2rQ29jr
FFO3I+6WNN/TFe8vQM7iNbQ9uWoJ7qy8a43+vlGpp7Ec1mORpBY5w3N9sT5xnMf3tc730u94pl8O
hTUf/54KHjmwffeQ8favPi9vdhG3Wm9OtGEmdgPXidzyfZbcE6Xd8oSoP/KXhp0f+staSGmiRA7C
/4oA/epOP9MmZUTERX8jpXCsTOvfingUebKF43AHmaoUfuuQ7rgQCh9HFmmbYwUcTsJI7GBIz/9Z
lepbXpKG7jNL/B9cZn5Tbc6NP2gyZYbPeg0rppgjzLPIa5OcAX4Enpb4SwpOi0eLyhbTvRX6vkE9
Tw8xb3FgpHd40JmAmYNfJvCrQN3fcx0Y5IADUQQRpAfMwzKwlSmc9OHh2C6xOVaAAqAenjbojiwG
9rNPHg3UbmSF6p9Zxe5tgsrTmv8ES51qmPLo7kYgyOYzCl4zfkGQaB0Rd2Mp6KDBh9kxehEfDAOD
RnZmzpkfOZWenWxQvPdQ5SMn2L7J9N/dHpV3leiDBXFiD3xFHriKhErYj9EgzVtKelY7VTBT25Jn
iXakMdYK8a4keNnBtyW2FkkqlmxOcH7fct9aQybZfV79JlN4JyasjUmB5TG9lIQZb66o4iF0Ld2b
IlFXhGZOf4KTqkmAEWFv0bmi4hHkpFJc+vkjwu3Y8sfTw1o3GIwSF/zqQBddQEyOElxXgZDvrr2P
ZLSt6wbC8VCbSYTwXw7z+msUOeZT+udE3hgeJ2jHZz9RfeklvzVFGonhjlBenhBUjBzgX8d8OW0y
L+dQJF3aLi5VL5g7JCGXYx6TsunLWskgfni8hZL9cVGmKauKsNiGnU58O405QuLgSkxL+UertuTK
JaQ9xtzR5Fgk5hzs9VHUFfRsZa0yAlY94djCWpupidpFiXhlVDZ5etPhgPkmLYvJjgL6lq8/qPU1
nh6isuXq+IlXTbmF4ELG/oyxD1WP/gN0ZoN+u2fqbv0SvTTsiTcdpSyPo0zJv/lp1lRs5vOmxMKX
6NKQO8UrUpNY9EEnKeMs9kYc932OWj3eNVcBpNqNYKz6TCNw5wHj0Y+FxABApxlM3WXUfrHHNKq6
JuhTdcRFdVTUjH9Ly0dpz8vGQp0rPhxBLc6RnVPRmTLf7ZlbK+bPBdKlsT9qvWhBNJbytqDiiCb9
4kMJ4kx0Q86WbUANXsdG1wd88C/0VI0w15BigGSTViHbCimh9xjn7xaJAj1f+tQ4dYvc0mI6pEsf
4DvS2aEPVFW7RbJGowk2xMrGsp/XJ2ODPDcGfjW3iJ2fe/4mhLkXR9kFrYBdsdLDRu9QXYyPvlLr
kq6xrI+21ZayDnGpicORWcGHCpFR9jtlxjLO1pc8IBmpYipkCcQga/02yej5OqhVpBztH/TwMEgS
Wmj404NPLDi1o6yU42ic0oi2XQ+kofODXMOUWx6eOdKTqYdPx9rrC+UBbqCuwcZnMwbwtpXr+OZm
Pp0Xl3kitYX17/Gws69m983tikytH7t+O8vjgc+J2emFP34UsH1k4PdvLgvvjqyVdpQW01GR4E3l
fDjtFDNkIj0ff7J/b0N9e8a0iwFP6acapOOUJqmHrK+OpiWwmjrUIF1XFRmsw+V/OnUgOwBcRx1V
wQJp1Xs4pRaaaWs0Mt8gjxtjSrI+icxCEZSoykiGkx1zsTjb53vAhDC6km0q3G7Q87SqHF1Sxx0/
L6vICbGppHB/Voml5zEoVG3/OLHqRI5kGOvbJRafjPLHaQ+pE82eX9qaJvicIM8RvwJkQseBMrv3
rCkk+ZjgFWKUxrRg+Vhp9PLKQZFO1Ofw2fYL1+ihuK+4lY1cXJARhjKnnobua0A47MxGDlfPfA7o
bvOxeJSPRaKZv9W4sgArrWoJMdYOuiYU39JHRz1voP5ucipBU5es77NXfs/2+oMXHTCWwo3na99s
3JzzgZoANuQEGnoKxevDi8ZjGKUBTxTV/Uns6pVAEmGGUje0n4/BPO5I46Dh7bfHnL0m4TogN3My
/pXEQZ/dpIUNHM9jvLdj/BAvqsmomGEPf22FrEhD6RjAK4sDu6g5OwZ1t+LsVW17EbotA0MbcOsL
kK6zO9+XjtwyUygYem+SGwoBQQUfc4JbzNvVss9dLqLCZL8NHKKs73Y/ZCriJTyKUFa+bBlmXXoK
mKKPwM9bWTRObU9/8hNwLBEhoGJ9u2/XMw265uVNNjFdyrQmOw9B2xJ6CZE0LKd60zO1ZVVFgowU
hyL8UlG7xlTxYHbxELrhnO8pSdigJk0PZvpitqRy1IhM/Y463wGac5LAcoh/Fi+s8uj+HtbBzw9H
X7+hjhAHdp89NFnQ35xqvkidGkUnmFOw4KmSYzTJmpm7ufe+6fII2OlMMgm32sw1RlSQVFq/E/Ub
SJCxR0Z49UZW9vPQ2RzN0MDjamCi8MU324fecnapp1SUeqoyLm3rDKae532iW10QaDXTzvQ04g/0
ty57369VDfjZMh84TNRUTVG06jBV2qEuxQeMv5LQ2dAO1gCEDrYgBQKYjpGJoL2gB75Qzorq77er
5QRrAHf3cUA36CWsLvUqEI0y0pwP+vWbXdyTyqL82yLRaJRRtuMSl9axxt5hXVfL2xSsr/oRrSvB
JCvIR5F9lyjz67ZVn68M6CpKixYHLeUl0ONEPcTmyYcPx2cZwBSH9zcNCq3lF1ZdpDYh2uIlFE6+
2L7+xxQu0t52OvosxIp4nwCF2V63SBo1UzprRLZbi2qqO8B+En3pNqCcXDULi/XJOeP77N+a97Mw
8bEcks6yGUjIJD5Za9diWJhUhxpZUp0iQZQtQfUu4qX2LPIJ4S7V7VPa6WnF0SMkLkXk3dcCUOyl
1sSxtj2dqmgaLytHCrgAHZYBc0sV2wTmlpbIHexiCH3+3HqsA2cHsDweZEwGY2+0QLVTlM1EpOD6
MEuFkreWZndcLgs3wFdL1aXh8y3R0tuSJjuB6rPfIJJpkjd20DJhTmPWT9mPh/NPfr5g0WpRfURk
UFXqxRrb4Iahd9apNA34Oypppk/24GKf4hp7eRNMEUAJsiOjudUcfP2vD/8bQuPhNAbn1unvXPPa
ea96f6wxrh4w0EW5jpVPf2MTVe2TdPHrD513sLLxN63u0DowGR9j/2U5XOn7bF+qljrx7H7loO0f
mVCNCS4Zk4HF+lJrXCzh3oh1o6efOZs675iRj+NvVxqY+bX6wmjji2fp0UfolU8jqFPyA/u3curc
nliX29NX7x5m5CXCifEgiywP52ybBVVoNRJEg5B44K8mJHbEZFylRGndCgpbjClr7E1ijogRiU6u
Mc0uIYiCnHLopxEpLTQ1FKG9z/NC8FpopcGV0pSUPJQaolB0+V1J7Os1Z62PKGHhXjq/IeDJCZ6T
OEgEcrnQ46CLyId+hdKtLnQnHPlS2ECejrGwsr+AIduYC4clGfxCbNDU3Dz4HPWciN9TEoSa+Xa1
cxl3mw7orxaM+kd111ri0LK4WFz0wwuNzZ3QcHoUTxxDHSz0aVuqMrkuK6E8PPAtWZ7sPJFWQkNr
JbePX8tChaea6TJBhMUyZNdlDz8sOSHNjolfzSKMo9vxa7V7nTPQvqORW52CSfwluQw7oROwqY0+
yMUm+cWkPQM0V+cs0wHhRvfOyq0BXOUvaz0D/nVTnHnBGX657tudHAb521gpd84cuTRYtYeT6G4y
zTpxQ2oDAtWqmlke0Oebv+v/ZZB1nONeicv2sCBNBppTWF7Qjsy7QBxO3Vgp5SiLqPTmcaeLi/Yl
NZU3wMEBlLAYSAcB5WT1pRZcX+xvnUrolekOv/HAdcIR8wuP3iWrNgCSTZIqvwfqLaVzMAFQt/rK
0KDMIdGFZAAN/gA/st/3uKg8KRJwQiyJkjMwFC9+YYGZBmVk9zDhR3Srddx9NfoYpnlIVF4PgLb+
lUvhnugZUwxwxTcPwmCC80NQmlBbgHoAdjGn2+zdUAtIkQTpimwBK2k9sPKACwiYBbFPIUo20Opu
cfqvfwdqF/fuJlE8W9efNNDIQCME64ueszFcfrlv3x/l405ppljd1EQhhEeK8TpZCs4Tipa3w0Vf
AkEldKNlt755ojy26GNujU+tZ8p9PEkOOcn5lSOSG9k4rkrgIfBgBGRn+v/Jznxh1bnQsPTcBJ8s
2xhmEmkaDvGTF57IDKIeRaj87ZJb/Ww3bfwbH2ltpbTdieAB6daZGAG0fUHYuXbyd54m2kothmaX
IlpGXWuHQLdnwoyrFTS3iiGhsSaDUxbCrKIz5XeeLK8i9B7oYt//4cB1Q5UQgM4D73nvU1PcqxFM
3U4qzFJQaHPUhAwC2nV8in4CcxZE5uDZEOviFE8Ik14DkENkwf0HBIICHBcmErqyC8lojgPbEDC3
PDnT/I/qm75tfmwkAwKIz6lz6v/WXY7BzrfTIK3MxtdrZCo/CyERGh3rUPYzKleGIzsnJ/rAeX0u
nN/FBqk4PELcON6Y503ermMPA1b12+zCCW+Ky2Bq9KB+U8lh7WnXr9eIV4sEM3QOdUOW+nZiIyoo
qKnhP9yGmsSO0qH73ppnFooT/1jIwmvshCJoQGIAtsw/k5VsmkbwQsNZ9Tcyvij3SMDSPSoXPK8d
N9b2+yP8n8alqwNDP3aQWc4+i3WBRTaj45bP30KilfPEnwc9P68LT43HgpaSxkmKpaHMmqsUjt3w
JnBC+wd3WNhGOImnlSXaUXMwgUqPTxhNCGrh7bZSvyVtQDU7c1rIKXSR0a3vMnne8udRRqWhYa+/
S2QILamQk8fZg6aWFopq0OYI4Hdv/rIu+A==
`protect end_protected
