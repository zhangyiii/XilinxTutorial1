`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cI66OANCJw8fIIQbdpCG1eUZiUrVUYlTNQ823416CUh5RU0Z0lUSscJg0VdsbyeOG0GIlqnKKDcJ
g+441OyZKQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UgqPJ9i9WiJwgzx9hA1QFTAyJQbYygHQhueZLDtbtfbgNYIe9Vf6qQf08t96mKA1gKActJ7BeV+K
6uNMiJfx/3aUXCSX1zJ6wf3n++OQDmqvxVVq3gnHpb+740+sx3yxZnt+NIQn5YfqgmEXSODHM65H
T6IlCQG0Rk76FUmssyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JffVUoJGoNenA9JkXMLk3KS8XcomfWAzcMGUl6pS4bKWUvYmY13D3pemGWR5ICLizj6/IEASX4qM
MrcOHNOZ78VNNGbrwydnmhep2T8HUJ/34A8F6RlIg3EPqaoJseDBIuA+1YYmvMYUPXWmDmWnG1uq
4OVHNHuSMmViCS9G0XZMw9OZMd079W0WWlGjxgCIsCbTxgr5NySjw/l7QR6gLw2PWlOAIibLSL/6
FYbf9Pq748eBFOa73RMaFJULQdNMNcUKu7XbHElWwAbBAEQETSA5PY/T0Ovuh5VWjxfKceXk9gE2
s16k5nL5jvgzFecQSuS2lSlURIB4qY5hje3ZOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6n3r5uCHMurGEnMpYNf4UX/MkeElsrXqvd4MQdfthvZDOuXHZxcs4tSf3laM+WPFVbsOKpN2K9r
vOlcg4pO3R/XBxH8buk6fx/j1Txb83yD004eikrbAzhD/XMeJoB+vwnOXVjryL4Tq7ewJGiuFj3j
3aajz5Netn79SPqpagQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ux6EQpdIiEpdxg0F62ecUw7+0Os42ovKYC5a4J5nt6L0NXwWYNruQn6thnH20HG3CkZMjYPVsVdV
6fsAhKiqralBKaBG/Ej9eLWDO0kqJYBDBHDr1KxCmmsfP7tgcSeensV8aAfsf43ITwJDMIO8VHys
LbnRxuW/uncBTBd8BpuuF6FOlCwImGuVwEh0SYaZjLlAA/zvuQGePlYAraOXp22pKz1CICW9YEbL
RHIga+6SQ98q3/eoFGq1j3ZXVJuLYcvW94K/kJlph+VD6UU5Kix62jbW5vyq5E8KMpqmJr9NNRFn
j81j5XKXBOZlfp+VVqMs7Hlviysaj593wan5HQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24384)
`protect data_block
td5QFuuLITbKOtkE3oI0mLzB/U3OEn5lA8+gSvm4NzDgr1xoKZ6KXCYimdZuYcgLb1Oo/1ycim8W
PFfdiPDalf8RhWG8Bm3Uye1fGmokMIeViJJFpudOlf2QwkH2Q9nSjhByWCvm5V/7FzruOcyzJZl8
uis+1q6Ca3nhUQR21H8IcHbv6Xy9XdyKOtDQhDkDGI8SOYvdtcIlVOvSvgg1PlHx6usdcjRT0U4H
P6/B+j6sbCmxYTaRSW+MrSFDCMABIOsqlOFl9PQ33XhNbwlnmPJJi74RG+LcTuZO3a+NNoNNaXCV
QhABenvGupCPr1zW9oEkPZiPmlL5bJ/hsRsgM6x8Xwa9Hpq/uA0gzr+9k6QCatYnkV1uffMfk+AB
tHrrOjWxg70EKI2/v+20j9bZDx7FvPJyBx4QbbJq5yyVnB1rulubesFQ9KK8yaLZwjAxSUj5t5hI
0l4yC+sfeXOFNnQChxkDiHzVvVEZ2ZDI1EqnbwvfWRsy4F4zYlvoNCRclytBjwQ0SNA56jzoo2pi
ibgPJl6O2vJkDEU/mqUOIjLBt4kX/zhQrtJg2imknPMYFFMgL+cX1RJB5qR622+ir5MwqoH8pNrM
MKR0DlvuT6NFrmdcNJxgc0X0UcoQlX5lLClp0ARhGIIaPIp2BBcnnQyDrmL3BGJCllWiKBn/8koE
IretlINJ2i24k15Ckl99bWLwRUtB8E8uu0QBmD6dPPijp36ElyHzVnNwvk5fAhv+ewOf/T6Wv9GQ
jtxdf+SfuJ/kyTvdPV/ktcIFT09VIsUkzpUADFZofq/oWNWh3OksJnVOLBKMMt6F6Q9DoaBmRogs
nHO8+7reweUYfqt9Pkd68Ho0peIwVti90VYbyohmaRni5f4UwxIB8j5EDDb2rQ3ZvOs4WU8AHatF
L9cdJc4OCUpYrop+QXOr8ndfwRgu3YA1ejE3j19WjwJt2XyXG46Irpt/+v8q9yQKawk054ywesn2
HxJ/5CQbbiZjC9PRw0Z97Qd3ZVDNGFOPLvlzAW0lb1T5fuECYJPYZNxt7r7YA7VS1rzha+Wr2+ie
MsNYtZ0rJLR+SNttgb9AWbjsDst5mMroXIj4bxGBN37Mf3O8jadEo5VlW+BRKN6hACMJO/kEIoLg
yHFS7Urh4W0pcXuEvqTTOjhI06W3mX9dIKA4odWxzGZXdWbBQ2XdsUCrIZWtceu8KQ2afp4vxO5Z
tTOxABNjUALSuubC4hvapzfA4Whg7qlww3VBYamoGqxsTWiut22HfYdkopSx62VFK0tGH3q4ok0K
iJNVl6cn38JbG6oXLCWuL0pDRfjjZsJ4IkBTYth538/zPSbbgBSrl1mlN4NGff0Y3C3amXvfL62J
78DkWy/o+w57JqJoOEUbVt/HQ5lBXjiHhLsxOWz6GzIrqRh9NsLeHRFqjF++toOOqzOeydsNtQe5
Wc4LQjYZ8qMVN7f01z3jik9EsaOZLMDBlDGdUQtWFw+EDXjnuwUPq/goVUdAQK0aBH9fhTyWiCzf
KOPBEB0m7y7P1FDZKhnXaWh0HgfjGDVq/5vMP7F6filhYmy72+X5JDJJFrnEINtnKQI3npB/R2gF
g0sH3PoOQgNYLkifERYPN4+qeRyFh3m+aOJpYpfQe1HMRfS46MdNBwfRxkbKTvCF3dosm9wJbPZ9
DP90iF1AAkPz1HfSsJYon96F/1N3B9GiaPDFAeyKXPLn0yuMyTQV5zYYASTW6E5o86TCvJFtph85
bkuKScqoeiv/LPtVv886DjEPcch6dMsYMNqQ7O3Z7bp08Y2sfuYijqFhRFOeWE2k7JGZUe28dhps
MJibZ82VPeR4SCjjwBdvWwpLhsJES617eGWPiaJ6xEHj8ze2LrrOaxtp8TgzQU0gMnUzGiJsiSmY
Cw1E/9eQIwS8yhNt7CXapbrLxCyqmnSiGpBL5Fut1OBKRrD2TP513liBX8XJ6XQHXonT7H81RZMJ
cyEyyuyJ8frN6ovB3w/mCbDgbAjKt5iunbp98yP5NcGOM0psBlOf4qcmRSC3baK1tl0GxV7sHR78
QIVYdLFjPTFIS74W8F7jutZGcgmik28xj/UOTKeDPqtfPqm5tGJqq+uQpm+myhD5NGvpKjqleAeQ
1e6tAkq7vxVNLDuZVyLJI0mGw97MecUYvkQf/EDuoFSC9hseM9TVH1kWmIb9nsrtuqoVv4h1iRHK
AIwceWluUcGfnj7el/e4rh/FLrIxdhd5R089iDFElWUcNdDGXnFfBEDh0FFqjt4JVv7rj/37zxff
7wZRD3eqMIzka5HGR7M+EwUYK97UKyMtvV4MslhYc8QR4YH5N0bC0qIYH3GG3aDd0fwWR0zprEvs
pD+XV69s2ray+kraY7fBGuYkclqoLM8RbXwfh2mCDeajW6q7tuAYiC7nYUZuQtIIU3go2JIpET4E
cvxjybwB9QvPcA2cGpt1ycz5K948fIH2boe8J0jaFU2uI8bkawJEA6XwaWJ7bpTmevaGUX+N27z/
N03A0FPFLrK++pWZtG/91o8cfkGwXGTnRJa/hhWYvX7szqVXuvMxbbD6Y5/YfOd0hwco1nZxntAu
tWfmVWeK4vVVD5AhgWG3xZKBKt+QdZ9491YA5at+4c79d98hbxHiM8LrGdLEEJQ10s0WR6lTovtb
b1cHYwmr5ievuTw31VxZN0MUxCyXlqGDkyS1a8ASCnQiQTL93pTaSxtuX3Bhuyb4vjk1H+OYLt0o
UkCmn5g5dQydbHLcNCnNanbMgi+VsQgs5luGPyPV0BE+kSXEQX+Oyi0EuvYLkZTHTolTQHRfeSJN
hjt5Nw0reHF4MtFjzQkC9HlmXnF2eE7iBDDBYjcecrlPCtPWXXfv5Z8AQC5OU/+mqqw/hKhllnDM
rZ9s8gfQoVqhn7uaQZ9Z8jlhemnnV8N8B+3XK0RBaoJqtbtyZn1Nfdcv0mLKgt5oNo/Rb9TDE2Qf
B7AVmaaYePvmZKPrq19PeMRKACDY4N9bGAMBoAj0e5EvFZ0qNvHBT8LpenEFXAsayPqEmZUROjZw
Pf4tjic7N4bMQktVUXmLtHIzb5oc75haMuTZ1b/djWlMfzfR5OIVVftN34Ajri/aiL8zDUwG6wK+
Y/0j8Xj/qEeVPfyUG3pTDTYEgSwA6GQ3AlqUV4Dl+DmMUeOAonsomczmM13CWd2lPpOBBSOm8S7i
0nyGXB7JjiLG8sDrTVVxVLVqY9/z8JLEuu/w8cEogqB6weaUFxJkjEBQwYxWKWT92ceKzfgItIWg
KVNuRuPXdwrX0e/MpiPvM3YhpQm241w+XILJxSPKupGBCU7cBaQj3kCLwosmrVh1vAHuju4GbHM6
++QUfKhjPQWyb8gtKjzuvjE0O22sYXN2uwMU0CVAbuprBy/yo9jkWyJlRA5yTnQLzGnnAbBtFUZ7
d/MjEiFQZOkzYP5vNVqlBlXOdCFX5GaVy8gR+q5qbBv0KW3YaUPpuMclX153sTP98g5NWTwVdnDl
0PXiLEdM9RnrYvhnOLS+6cyUzf46627NjIpXTXharI+3XG0OJuk4Lpy5UDb6ghkjsFZc3t7s8dDH
iJoZ6Oy/4IOxyhg7fchmNZhU7HmR+7+olPpBSXqIh8rWdL5vtYBNyUs5UGfBPgzxsqGQfpGqO8DE
EhiFJ79CkdIAug8GP4qo//FErPuINsUSg0qIas1698IutD6p3f8MAQSCYeZid7fS8VGRHEs4Xr7n
M+oVFpxyuFHpXYYI4cTFrzUWboqM6O76TUFDLhXXOEm2eoe0mztw2OiT3FCFNky5L/aSd0ISasPA
pfp9H7CR4El+sb6Qrj7+dGdRRjT4CclaPXbhh1W9fWqCsSv6kskD2LUmBvhm0VlJIOdkaOZi1Np5
6Wf7+DO363ViqW25EpoQDcGcwJgKE1Blx5X/QlXpp/bMeduYkuq+LaFzAdXcrxly1yYmu7JV5uC9
s1DuugPZsK/uUPSPHXQovhs/UeRj2p8VTBmQYbTg5kv3kVDEcosOKr7lC7cuwjMtLyojdOjYjudM
++aWQmoI0++gFM+KWWcPkxiLG43GlI1moCtECoQZ3/I4eOc7oVlA05moSEoqZlevLo97AFF+/m/y
8Wsv1mrscEDugwM+zk7i4RVOacbC2qf4rbe+zRrv1K5InwX18ceqg3+/pEyJZqbyLhpxmCOD/TUp
LtuJ2/0BvhesZjtW1m6EfbIbTLejn6gkt0GoL5rxNofP+4A+sTXeEDJO9cV2Txxuh2Fr75wNcD0y
P4GrO7tDp2ZrvS3THgjUKCo4mDXQ4jUVACBHDsbLfM+xQnowi+ldprgzB8A4P5HNdSzL+fTJhPW7
kPHeroIYJf7iSStyErs+X8wNSGh/2Cot0Er3KMd1jCt4TxBz52K41VXIHUXSVgUEC7ngLNegankx
JpFUFWm8CTpln4YS8B8DmbR+2pI/vtRgUJT3R4dvNbSRoCvCVBzoKZH+TWe9YNwwzb0Q8SjpLmm1
lizUWutqo7Bc/O7jRxdqVpQzdlMXZqzRIkohsTKnJJltCHqVk09/e2Thpb8BSsfCcnrAS5YGnyuK
j5SYlwSuTqtXONMpADYOh9U6FqJOMbS1mU4ysXFH6uTSEHqjmAXhFpIxbAw687xiQXXljIIg/0jE
4FuKuXa7INcxRSNF+eHCdiu5/vA9QuP8VllYsQXM7Y8x5z29zdxYy0Nnnn6umpxP5HiMrzRhk/Yc
wkVORPaXSAdPwYDsHaQ+fATU4x99778tbDF1DXH1x+aVcWElVc3Msi9oFCsJovYMqLZiqk326uo2
nkrIE8exzAso+ViEY9GggMohil3RduRlnGhheF48VNY487ljK7xxfXUsX7Jv53vWpustu/G7VlJU
zgi6YsM1N8BQmu1CmNrlvzC9Z3g7EnWdLdd//3Yfj78Mp5OUCHoJ+ZDCi31yjOfUdyRUqfbsi1WQ
gi6t2N2yx2EMhYtfoYMHNLAHwmYHpgTw3Y88UdzDkbY+5EtZPFMJQHAHroVeigBuYixWAziWabCG
kKM/IPqqIkRG07gNP5ns/S98M39FpHd2rJxKasBm1TGwdE8CXtFJIoL5Klx7qRZ2UAExoY1spJyH
rdymxSO3v7+450IA3mInnnPMnLoTsSFhm/xEnEi8T67GXg09eM8qUfZkL3Oz8cmOgBLOylM+tkOV
f/J8gMH3ygyfQ42RshBqzMkd5iyenJGJWxGy6rCtOZ3xOuL2/EpdR1flRKLGf045+W4o/LhNylRB
adECvXwZFfG3E11Eq2jjF/fKE7dTQ/o9uzfO5MGXutTl/ijAnFDpCxZmP9j/h3DQM4LisA6fhRUM
uC2vq1EMwRMkrFjKnsNRGW0sQ+VNGQ8bU4t1Kxv921GAHkwsHOjmKZ0BBNfcDEZOsCy34PZY3oBu
AgLwZBPIIHSiIM6KZTTaSeoeR3L1b43ykoDZXsN6sFdKBk0tfYXZUdylUbx/6faMe5SLosLw2yII
1RchmszCmZXav/AbQNmBw9TCvGBXxyJvx08rvCXwnKX8QJsPQgbLPxf5JoX8gJeqPvzs7iwUAATs
s2tEYTalWjpzW6+3lUcr4+t8Kd4uJPhwtU8W1XbK4U0/x4IPCSAQiHrHP+VIz5hd3AwXMmiV8wCn
/f/d0Wo7JFJTzkhIrzEmIZw4DYgEo2bHMXeMLVA+i2Dvsn+0OYlCgIK/+BEKjlI/zVkIegZLjBPK
n7j3z+XbyzsEa0CUdPLF5/EuoovTdyEA+h9TOcommOhwFnNqvwO/FyEnh5ycstRIzcdNgncqIq1b
qHoNF7Dp/uq/GE5TSVE0KQW5INwTzo1fe4LAcG+1ZWGlKJll0bVhhf3FTh1REzfxVax1F5TUisVM
zrBoTmI9j+igSxyFVVbbIa+s+K7a3ZsFYu+TrJHmHpQ8rf+pUe8ppA7SsowynZp1LI60cwI4L+PU
x/jKOHskm0olNjVQ86bkEKgmXDV/w3OpcYkMZngcGE67gEWzfNJSUlkahCrOqKXpuYa2m+QxgXmy
lop4MT40yfH/PysTsI0BymoDHLVX7BpncCIWWbGO7/vWPjt4nZYO5gfOjNxXa8LhUR4Iyn9P3uur
hXK93lLYryuwz612H9Ok9fNRJQsh86i8NqNphkqd8YUtInfhWQHftSEsl6fNnQSnN0T3/pMAZF3U
BO4idUuvgqgzfAveMOWigA0BBK155GJ2p9uKSBpHUh5GziRI8xvLtN4Zr//3/OvlEnEcsnFd9coF
OxNRNpx3quBPrl7D+XSI+jS6d88z+EmSbcwg+zt7ouYj6W/BnYHR9SWIsZ2DiY2gYKgyqfllLfdi
guUV6OWw32RPcWT/xojE3CtQOFiVL2sVHTA7lqlOQ8ai/pZVeM4AcrlQfnoZC8wb93KeHN1c02FS
WOO1xOwj10MtGwZjiSoT2fsGAJcaHHg5MfMta6X40YciIm+3xUtO/rleE4t+ABkq73vQAoTPvc6V
AJUyReSc3eZ3p/0gnF56FHB/cqT50p/4y4P1KpsGtS2v8hJbun9RqghhpA6xBP5xPWfhLXAjwI3/
cVOsoB8tJxmB5zdW+/9g5tjHtgGQvLVTTEdlc7Z1C1ZIjPbb0WrV4wSR8ixZe8Jv5DmISJUHxvnT
tq9jKnnbzri6Uqtf3mXGmisIJq1RevKfabRWnHQSpNrhfrtrgXxcieMmk6NKnhmS9E+yPxe2OZlS
ILkflfLKIApKXtIeIb/ZMjhraUnjTp4LAVplHZ2owmtk27DxJTQTsI+sq5Xy6dXPvEriu9qyiR7o
qF/ow8BqIk8DZQYbMbgwcAlpEbi4dOzzibGcOMxIPY1xaUMN1DxdkrP1DGrdg7gYE1wFaqjphLph
yXOtdeWHaMCZVfo0/kg3Q7vCEakQ5sy+fBX1njktGfn7jDoCKxQ5Z09Bgu1xtH9fXSgVXMePWDFi
XsSowwoLoS6hRaA9q6SuPItR1iwQ2s7HoBuB++7vLZZczuaovvu4Y81sWSlRejrY2Te510uGgdN0
6fFxTEzLet4NmXnFt8kDUaBmmeHsE3DusnTfnUFd6ehgFBzRJZ6Ok4eCSVBsZ0mg8mCjDOJYaB7f
DLbQHWpaIrJtPO6JvuGh8NOTDezmCYTq9hIDtAfh7uXNihOQ5j7RKFgKMbNDHlPjjxvDrGuAJVHs
nWnVo4zOt9hCMWP8qMpTahjzMN+xONh8HN0U4SjfuUQfFr32mlSkg8hqBYGJt3QsvPlz1gDeADRr
WdmRfUFmEWdewA09/Ejf7kxhvW6Qn13/HODW2nBF3desGjVE0oRazIltqkFnRkyKTt1G85yjB3c4
Uk+MytRPimfMp0b8ihfNkdafxiuwhWbfVom8cxUM2YfENAljn3UqeKfg6WaecJ7HHzSK7bRK3LrA
oXuaNGqgEEFAfsLznxtwLAsJEAp26F9/e3XrnGM3P2eu20wjlzS+ht0y9hUijSqAbTCkD2Ngoycw
UqGJKzRWuZbKPY31CMSuBwFgj+1QVDus7h/fJYVOpq24btIKFEgdGFTUKG4QlHqPqhhbUQyVWRpa
N+uoXZTxAN/DM8TifvBw5GH/B1/2sW0l1dq5OwP1pvTTwXv78ukXvZV/s66oC1yG8vKuZRteMhh/
2dka/IO4/xQVV4pk8tdyUMNBeADz6UbivDikUqmX+EkpkbIXJkx7k7EcBPjaBxlnjwXT+5j0PRF7
Tq/tDoYv1F+i3EtLyU5od7jYqkTmlFLsZrj+uWcOrB+LO/BjkdS8WqLfzg5JzXe/6wJGNxKcZD9Q
AS+tkoJS28aGbz4B7s8iZGmMdqSgFZWRb8Kwhi1GuBMYTM76hrNZubIjFRv4oPiXvh8WYezM+qpc
cgVI7C19QZcmX61P1J+z583FoPu9CCsPEXWfD8thhPn171z66mIcCADA1ldcRR+43XytzijCYhkL
oYpyydYyav9hglbCE1vUu8k/4v/CeYsIUpHgCptZ5kpnb+T5IBv89oBetplpfLQPWeL6/9XAk5J4
R54sdUxWh3ihTxJ3BRhq+73A47iKdIqqioUEjSmIweunNCWKk15nAUtUJfsmfIbM26Vda+MeJnns
QDbkA3w43M25XK25NMGpUUvoeKs7+z9nPypeSAHANDUWFm8ugEnruL9X+4PdakW/97MjzrtI91Ls
S8YyK22G5iRD4vDUyAzq7hdOKNjjMt8aUFHr3Q2Dt9HcWUTUUYCCV+wiiI+nMrDrtaii0xevrlGy
CWSeH+h31EFF9qotuFYHh50bAAlD16zx+2zLsQY1waXRFWjRQ1V99RnMw0LyhjJWddKpTmuxMti0
eY4MXjX6BRRECy0E/gXL7gODBFGzPrDYlUV9ZYUY12zZr1v14COfBytX+g7Qi4mcJnWSIFQjiZui
/DyDyRfx4k9wWWj8C4/NPzveQd+fWS5OSpbv/9DzukjJLPtMsT+uzBOx6LfbvvMUChyNnqBMudor
Rkq5xjOvLMCiRvqK3in0DjSAtvzg20Rs+K6aBm5uysY4aKJpMKos7ySrcR7fN9Mv+IBX7aPuqcMV
sX5tx6r2dpj0NdBYrKil5eJomaZHewE7Ht3cy1fnmvf3S2QYGF/OGUt31NEfUxHjZTpWeDeaWXIL
SSxgKW57kmepVoBH1BXjHDcabdx5KKTcuzWqOfEohEJ/M4JMhOgNGUoJeCrIcdNbhi9dCRC6JGr6
1mPNDR8c5LonfdId1s64B6EXyeurjFPexuBdjgeC8jhiR6BGKdmcfWSxV2C9WYwDBGUBus1Iduzl
noZzVPYFtLPHhMDXvdvhQdj8mG79x4G7ioaI7wKw3XGSKG6+W3POkSzkHAcvsaoSEe5847Q3EQo4
IJo3Czdvdfh0pkKfNbWClqy2fpob2H4qrQ+6cGhGAp7GFpZj2YHinVu2aYVHOTcQ9wR8p6b65SE8
NELXnfBfNs87XNW9kL+96DpsNga0JeGMxxVu7wnnv9TlAeiboss5OEX5eY6A7rnbEnjbCAqn733Q
SbSzDCcOFedEj/oW8NViioxXV+IXVehciVtghasBLLgVYSY58sphsMXq8ISK2mB//88i2CamxZAW
XK+Qob3erVDmJ6ztt0wXG23D9NE/9nHOfahIEbu3Yri+mqYM1XqRXJCaCbXXlP4ZtFSfGBXxmH7Q
OYSmraeM5HeGbWRfiO467OIn3861mlyGmNYd0krelA9pb1iYqkLsHHJlli5vCPZAeBQExWXkqV9G
Nc4l7O0BhObT8I/W/6pAEzGzVUqMsZLOd2V+7Vc0Au5X9laMrB3tnZECfldD19OUggkifv+QGOBt
SZvpmeYhCfJWVU+sUmki7DCbAvHwUcVuMK6+E79eZn3yTlyd7dtshcOKEVAheU+BJRhQAnfFPGiG
FtaBio7FxdyQCkv5Cq+MxgWdKwjWitW4MWzYRCMVvKkdbezhEa1n0FoHVMbnH441CSn/9/SYp+Gf
HQAR0Xw+mXo+EcQyfiOHxprZO3c6sJJOuvwFYhwFFfWJg86eCcI0j8C4N7D0tQbOZpb10sBEd3rG
rVLDOu4AqMaQ+17VNimV5I27XwsHoqBym4LeLm1Qf1Rl7GG+hs+QBfwSHv9uygK7nT8M+n8G/Jz5
2AFFJiDwheRnL8qMgA/PR7GQuJ/3Qkgj+wTctwMWSPRkfROrOQlJDmPmhWxWedBxmGPUwdyL7GpA
tz3lXuCB+PZNr/X/4KekI88yOdMRJwNVflwBstCDXzIdYRGxU4qnW35Yth2rk8J24wJXjaUQeWNO
3GpDxOCw1vAb1Z7h3vnvtcad2CUReqy34M+O1Q+iUnnwFdc/kERWLzmJtuKGPTY4+9iC9Th+k5kc
zyShio6esQmhSbTtpVovJY9JaYW61JUxkwZNDiLVM71rjmT0yw4gGZNGYKiyY6/UXzVGp1OW4cHV
7eyvUq+ftlwzt4rMSkdMRHQttf6vOH5zRQtjUmLNtNTUD2Rc258My3A384K+7BTcItgzF7AM/qRN
cu5bC9qmKaA9oybgTQ4HJW7T15fiLdodHmCXZVGcJU2eoZ9+20q9NYNM1HWCM3E7Q2MKhkjfh8Y7
PHLo6aqKYq0GT5dt6djZEL5OrkR1R3hgVOYWjrpMXkq8DpEqfKhj3zNfeBt4XLo9z077Jv+IAqB+
8ifDA307R5xDdcXBAek9Vi8CR4yqZLYVU7UkfWEmTwDn/nN9/sv76dNHkApiwab4lXTokdon8e/e
pLABXIcsOUTKs2MxFvcKqGVd06AYtU8bF1O601IaMJ8K8ylUqb18Jj6Tabs1ACGD+Dtikf/4aLrV
IcIJio4xgTYstEwfGZhXVFOnrNN82CERr+xYRHvs+e8OZyrVqlK1uAai3DRrbRDXmlYheePHh7Js
4ybOX45qerbacJvzXOl5F2SM/QP6c3s2M8SS+26pdF4It+URbrYspTwPdJZMjBcSZZscvuvcR+7q
2TBIbqHgJq3yrBCOSbbwLaaDgNNN6ppJ0xPJTFKdLiuJwYD8bRk6ONRYazVWWgyXoM/0klltRvdZ
Nl8AaQJVQs2m80MGlUXa3ugTwo32dm5oZ9HKOxMtxq+PkAN8EcrxXsl/C1qotrgm30V3bvNhLa5N
Zk3Q7e8P1E2McrLKkBE5W+r5E/duLWErGPrGy9irhUeBG0/EilQ3VIpwWZJIsqdbJwJCNuvp8c2K
eFju9ynOgkt3oLHLcfxrbCcAAzoS/IWPoUic2Ofkvxt5bAsow6Ml5T0w+KWZBfCt+QWOg2dfpinc
KK7RQnSOC0x9SxNbnTgZxS7klzQwAxFeOEPU9Nun07vBnBVmMbIOLcx5N5/obXK4u5cZN6S/cWkZ
0JhmR85GIR5l5JMy49cqKhnQZpV1OJ7LOTCL0Yh0N7pJ+WAFO7Hkq5L9dr6hcD2dyi1prnwjKmBy
aSVocMLXnn8ceNTEXrJkFQrEW+WtuCd3xowgBJdgehnEAkBLjZ8LwZwwtouVM8rZRKHSZOcMdYm0
gN/r+KZr6JwuKLLDxZqxJoGx/s0I5DSelKxpGBuv7MSNsDSX2v99rkpqqR7vCpUX+SWAOw60GTI6
Fg70BNAfVf2gnroLJmO0Oje/3vSIf70jXb2mQLRg5ZTDO7IHJJ70MmJsPzPmKvQeHF7vunSPGwUH
gw6z8qkv2/j4VPMQHIIP62bRYHj4KK0LxJobU/E6d1iUfZ5gFIe7kq0iSk2bhiFvY3YQHpje2VTF
JBwU0zLk63so/5P/J53XReQoq1IYrq/EqiGF3dV2rWKcqSyY9osxsCRcFy3vLEY21sp3blF405Zb
TmESOFAOLanshQnV5OBNdWbM04fg5EWNAZY20EjFijtH82HzUFjiKJzGpMhVcliPzk5rHoKPGB/Y
FK+JuAzEkobINVX4kQeMZ1PhSKSp88aBfvxKNGmjnBUdHo3ihTAL6wbcCTIWia3Q7dqANr/VBoET
pnW4Xee/hQgrHUJvGYYsJWoiqu0f9M1QWGE68lYnO/5ezNbp7e1bYokOtGP7eVrC5tBSCijkxaku
0mUJrRnMZkpPlLnCo42KVfPsDBp+ls26Jb1mHyyptkMl4lga9MKo1wFthhf9/oKJ8Ts0cRu8CaiK
38ewW8RD3ID7SyKHfaSZ9vkyUqHctS091pwYuUKZydy22FLn8tADha3+V9j5j0P+6Equ7FRj1Y8G
vOGutm7FWs0ABY68fixCwmJsmvmZz7BHYQoCZsq7nFIdGtEyzV3/RKLMHSPAXnpnw4KBbrqbKHQp
9Zedp5Cq8RBHXJGeEKOjTJKc07TsQoIYo62S0JFDogRKuglMQaayo6gfkUUZ3uETzRSqtHuoFsfz
1GtZFLrqiQ5roI68gLHYt78mcCH7TuPLAzLn+Lq92zGg51g/a5EbMzu/YMYCexVjl3N2/U6jScSv
s6mBsuZzNF4wArT75BsX6X4jtrPALHakzsrv9LFXQg9ylnNG/Hx785sq8mcRmhsT5Pp9K5rRfHak
/7umBrID5oIaS9Ny8Jzg5Kzs8eqHmxfmlujxH/8O88Qstxefx3kqIwZnvQTSgoNszPF/V1JXX5WU
53W1xFyMcvk1woznK9B13CinBQd8uwYaX0hnftZvmN1qKCjSSORtWKDnH+8uXcRdap6MTqPtbqqi
7mawTYouofgYvMo63VfRFNQMSEiE6wHPJiwlNppecwGleuXsWGC11IDqmOBHRDemn2thH405g6QP
R4UdfcN+Ab9tSjB+/JM63XNS0DT6XyGEH06kjidohG3aoGMkr/gb0wyqfa1ULv9aJNPXFubrsRz8
K9FfAVjaUUxtuUwnhPYuYCUwfSX/LPIBeYnNI4QAL61ir8axsM3Ev6evCuPktuTVbZJeI5B4aprx
NY9UrspuG6PHCWn1s9lNEAo/aVOSsxKhKXevfyk9xwY25oKv3O+lsZ3Fwg4HC8fSL9u7g7Jir9Vw
2LAknAzJMQj6HyKPy6u29nrvy36ReIzTu64qLUrD6SVF/6wqkwYRFyTPFevQrsa6KvzT68PuC/cz
rGwE1SVfwfnavw6N2zxepEUaOfKMZvTAKnnrB5Bsj7zUa+Hu3NKMVvD+7R64eIHCvBYpcMhcX8K1
htxOhxKHH0G9+WV4Fu7KgN8kArftGla4XR9ihsY36qwmzHHb9S2LwIyLydMIFFdKzeX128bgHWfd
0Sg7YOj0crGmKY5wojEAz6Oexyl+RBZR6QNsm66XSntCXdowxCQhpA8+R4jrW00ZYEw9As5p5fsd
/9RJULIQO5cjiffDSwLFLBq9ojwKszc8kHZDayBHicjdCTkSVdWyWKdhVqiNWRq4V+wvM21n1ePf
LNE9YKSpqIf2rPrRhJ0f5KVDaKUpPB9HYLfYUy4G2u5q/Td2uTyHvEEsk7yut8bHymLs+TyqK7Wb
zXDDlfDYPr9xNyNMvWCc9QMQXEZpzXshJURA2wTj6b4Hslt/FDf8YxRF8DHN2tfFXeT7Q6H6KAGd
TeGh5CfXxfJAl2XuguYzg5xruc7jlNntwDzgx8jHHh67naA4Bt1VuuEIpDU+yJJmE2K8IA5eY41O
2YY+U2LoVpuq+NmvSSRhD43f4Ru+npvvm40MKDgyHfZflNKr68I6ckiVDhLNXuo6OYeHmqlFp+sI
vCKY03ThKmYF5FHckG6XUAI+lLwFFNwAH/K472VtFfLuqL6eRqkfQ03s6sl6ftYCPz8VzSVrNvqs
3ZnE+K/6VKmwITfo0ww40pPsQ2HfWYHWnpdP+kbOdwN4JDMgQWMf+rE0RaMQ6cNehE3mw72qLIht
cwoz2DNti2qaObcWwPUKgwm/4MNxlQ/EefsJFkmGmps0asAOC2n7EZ28Zb7N1maT2RWcR6oj9ksl
sUvEOhHZ4VKnZSnBhrRXFPPQFzzLWkqQKZyLD8uIaI3/GWrer72pYVn6eIFpVZDqQcpCKZvStTjp
EZLiPdt3PGGEpdQFpCmWQHTl0ZAfClJa4hzekpnnbOglCLQ69gl1fRjewMW4Ges2o1pARPlvurDY
czRAR+B0XmFOruJVat1JkxyOIPNJ9GLOQyf4jmz60RQ2WWZnRfBg+o7anJmHwp1vbi4QAr62tAyD
BSYCk4Ou1UXcES5zvlSOp2rk4+Q28U8Hz0cJYG2Y+u9hglSIjshplYPGGM1rM2h+Gfb1gXQD5NfV
xXLgYYKgUFUjLWBDuVSgTvrZQuOmsx9KqixL8uHARXWMGJvLFu2By+x3BTTHlU72r7Sg/OEGgMBp
hHdezg11Yxd0zXdOJDKKMTcJFnPtzl+zI8+S7Zv39PxS3t19i9koBD7xAu7YoU8z+od3hSBCZp6B
u/7pFyjspPOZRg59T6HFf4XPJZ8/R0mmcSg5wD6zQf9nWiwyMtqTRVMRY36cvBjFLAIHHum61Z1Q
MLO4AsIMmKcY4PFtOJjoaece0u2h63TG3pSH4jXtMANmHJTMt7Lr39DSfh7uRm+NWExYAlmI/+yk
RFFvGIfF5N9/K1ihUyo8q9LNUOvfKF+80yJa7HyAkDB7PAKMKd8iKJk0i07Pf4ynFlBs7bLc3m2Y
4QqVldeJIxPrCFxZFHYaFNoFZ3x/Mp3OPj2UqPq2+/HdCYV/cVVT/UHY5URIRdrkZGRf8uZKNS2z
FkYs4CU1IjV+itZdcbHKerNoYfIyBE1MRQE/6AfYMqJPEeIsSVg/sF6xvFrM7+5g+u/nzb3za4Yn
a93x8KfX/L0X1eGr3kc5tWdiGzCs+grgnHzryZNzdvtK5DeOd03lBUPHfdmGtjGNM1pX2R9uv+3o
pziW9IKVceIomPM1jkuSub3fSE2L5Lv518wyUP/OFC9vA2HVWesH/azPmsxa9kAIxRDJruLlPJTz
x6bCln6cB3W0PjSCetw3YdZU5mkHeg/URWWkEUgHi8YXmv446+lvJYaYNhgtDrOXLlkQKhDwwTNu
dCMjCnQ44KzZEbJyFIN88Zd74Ue7aYZACSimic1XmoL5/iyQzgUBu0eSeKqgyqcq6FENtftrd1Gd
Ao+cWfUV7AtflqooyKowRUsLvG3IJajuPx3MhUql54Q2KFseUhw9Fi5znVUBfuKBQ2DW5KRXl9v5
MXkqlayvjWNgC1Sd2D/dJJ76T08XGKRVgLPcD9mx4tmrcUznMOdwSImU6nRTcWQ2qxR1zsWRwtAh
egwqbmd5J2/hM7cWujLH5a0C3HcXMNfF7YNyZwmoqGLDVAoreYSJvd6j9EnZyY0xfJdVQZpiIPfN
eq3ULwN/1GuqF9KxGDW6WdOTU8XuW/zwM/Y15flNZ1/UJpAjBGj3zlUQfFVtI8+UnkvuAWdJcrot
Vy8vRPx7/IF311eZDo6Cb+4yifQv94qJ6ygy9J+szaH0feq0CmFoENEUwgr5laClFofoxC6C6nLw
Km4E5syk88MogIT7XXfEsTLvfrKGLTM9JlIcIq0CU+7OWSFOyiwnSmH6dvqbRYo2y+uWLgv3TCRD
nbid+qYdVsYBkUUtmoydqVydhMzmKz2J7JW1YVUoGzKbVOsLVHXW7VlR8Kog+BM8YeE/I/M25DIT
sFaBAIPlWBx3Lbge3f3Ic+K5NFEqaq5YnkYH1fW9DZcI6JkglLBXlH/Om0PMfGL2TH4cfvKXSxNu
o8B1VnpmHdk2SVjoKVCFM/afQHwubQXauHGj1VN2WSeHekZxeVO+w54e8qCRCHqd4iGpR+YQOFHC
Qpj+QKcxARQ6NRLxfzH5t3JFYS4UD9AmOQJnQ14AoC8TWvEPMwXOXepeR+g+d45HYr0nxwNyYdZf
2t/9zXlnYf784F54Q1vRvX0dsjrUlfbs/wSpSn7xMuVgb7sEOhPJa0e+lrSVDFI8UsSQ54ecQrfq
Gjv3AooQrNOlnG/6esufcEJukUnQAkrqscSH7KBt5riqM2hYqq31GoTIBklCjT3FhNftbm7BlP3u
32rLLqZmRVW4ROiFcwvIMnsbzP6c1R/76CZ1bR+23+GuXbt5OmvBzRc16fjb+XcmeMZhd1vrU9E/
RvZBUrwFocSNDaU49Yb6UkRnnB2UpdOIAyYJu7+O/E0bMD6Ud6cJrFVRncqV7hKo1pl9GFUiRdRK
l+fT0ssYLCpJcxSeFIHkseKu3mUJfBQyVCRj9ytnFmneiyBysRi3ZepwP39S1/GDrvCNyGdPUGrs
NKIiUf+WdDkq6atcsOxu/j/0gCxpihPPMtNlBbw0dtyLT5JTXPeM571Nvo6sztbwY+Z3jPRxGWWd
p+AVW5ikWYCigIbqP2vCOJsoQocAGXtlMHJOn2WCCDaMcltHwqPCM+JYm61kRFZBRzYAQLo85oVA
NYSl/cSg0OzAuAxWDf+yDAjPdUZEHJBqPl1ZgO9I5LkDfdcibX64TiS7kJT2TFdSigAi61R3FySv
ii09zdZW/92Ts4VEVJ7cRjcvJor8cg/rOrBeFuFWaklK4DkGnIJ1pzRIfhoMG1bFoGYm0bckv9V3
htsN7iioRj/f+N0l5U7S35Khl6EGUc+YxhwqLPeZ54YfvGyKfCvxU/I8vXrT2MLGSTFJUTdGOegj
+jKpsdPZ2CORem9CrHcmj7JyYInS8PRlcu+vaC1u5Nm/0kE4kTCpfYay9uR4jvSRj630UikMSV40
91bSoTWrt1UrIFk+KQrW1vvEEzeud8LuoJF+hjTZfwMutNNb+XvVXCybvIwys0AQ10zjSXCjz3et
Za+qksi180P68YVUnKhP+DYaJIch+iyVmHqRlyoLSfHYrHknoApGHDmUdhDbbJaYjqqQxKaMKK1W
fWtNXRLhIIsvdYPDwdUnss9gsc81EqYE4RbTal7vKr9gAAhh3+K2SxFAKW2f5JSLtftvrwXYZwaL
rn/YveJaaKtsoT5C7oCFqCTi6kC3AhPI5TSQpr4iutmlI2PvdaLapcK/E56A6dh8GqgkrupJuM3p
6sTK0+osG5Fb3vtI7h+nu2+4OlLw/cYTXDjbceVwiF09lUTuCH3WvH75e+wxHx/xWgY+SxH+urUz
2RXMItXMz1h437/qwZUGC5x9MYYipyVF7hSCrrys1TBXV0PCxksMmyCPBe2JjxAZtJ5KcWcfQahe
71seAA1+aTU/AvF3wVX0YZVuZQgiHnrL5qESIk/GxemNR9XX/3ejBi787n/WiA080mWnj2JKBCWu
IG7jccXBvnYIzmPem6K2+V4mdBpdQN9ptHtoothHvX+4ff1rPqgxPYasR4B5cVFVhlpFS5MLnX1d
oA5EcyBu68XznytS8RhPpivkb4V02IHqcS2cUe2wWPF/88neh/9SU0PIcnuZg9QpqPqrG14MrR9E
PmO/KH3LSqhzV77spfNuvZcBJA1lnQ0HcvG/EynsdAilZAzGUhUX2YMAyJcYUD1PRW1GRMIhtY2P
qsBBVgTrrpRVd5gVl9GBGf/4nIDtU/RdZl7JfvpsE6i6tdISMGpMSRrYOivjyM4+gRrGVfBb1CDf
Azv6Drbh91x/FH9ZMZV7i6xi9W8XnTGDuU9eUAYUmId04JS98vJQDeQ3wuLWUgGDf/FGPEBNC0zk
c/bXyTYooyMEOwYU8qE4zWGGajl6eGisjYDdlZsFDE3m5iAoXFWovUXjJH2trCcZEdNcMvDM0oVl
MfdjvXDp2W3+ICfMLGYCDADrvuuBN7SmE93OKlCCm0Dx/3r4QQIlxB0xTkE6rUnFDKq1yKeNv2X4
BkNhr1oCaMUk6CBpL7N1435MTY7NTjEd7dseeuKuZuhm2NGTF7Xsqiy9D/Xd7Ac9RTZJJwN6cWHm
3DfcwVvty2VLN2I3dty9ZoUanHFKmg6D6tDs6IOT7IoFPz2unO/giNmHhygf/2PZk9XPDwpuNB3r
nM1Y+dB1CmPAkQ/IE68Y9WCakZvfibJHTmvfb/njav9GOdO5uzP+2xozCWOWZnok7xiJ/pi0HlxF
Kxq/3RJQiKIy823sIUoH5pOZWNf5nlQ6h18lHddcTuBkjxFzAW97gqb+UXRYFHZRHTmoV9LzeZtN
B4ZW2bKsqZUBoz3lEfgdBj6QgRzsGm54GOaUki7kSSqxk11X+frbZiGKXtl2h9DkC102V1MS0XRk
H3jTsWEr8GhiWiwtbPBlW3PwqCqpPHpPnXhsEJbsnWt4uQt3OJ7xm8cKcMx/TrAAFAjQcmovBI86
1XnF7sNgC8PF4nh4gGo+khLRyJnHewXrQzPiWsa1+nBWmpETbDG6qEGipUDPymw5O43YVrIUng+4
/ocN9TuFIwxs7gSBvfiwSJSCW6Jt+uK2S9Oi/219xEwc6g9xv6MtoIDZO+IjwpObD0naAsWaCkyC
R0tLCQLqj+6lHTmpOUiXBX5UCv3E0Ow+G9SP9yefamW7RcBGGHnslikRcMDN5ucvje3U76FuVOU7
efjRRKkMVN19PWEDflgZYekp2l3MfwhYmhbl0nGvAZtA1ZjNxVejj18CEjslCip6McHqB5+7IIUx
vMWyjg4+lGQW9xjhOVaSeIob/hVH1GfheR1LDPfcrGL9Xnrd0eVMxKhoktBgD5QOpC4jCURsx4+Y
2LhDIQEY7EmNIEZ4OetOPna83EJ1W1Y/fGK/X2u7Sa3tm9e7hexbwRa+EMjk8kd7zeJXT9oCLybm
yrc+gszrb7qFUDw8lphi6LAypfh92IskI/qON1Hf1lM323MbEZ8owI3qud1HUMJ7xmPHeNlCak3u
OnBQxZjRpqJlaNXQHAInohNPoD2efCu++xzO8QNcJsve6H2UopdC8jpFq+adNNH24rypWERKp3ov
yQSdUgbwbWqEa0A/FiIBoRRk4j2GkJk7kZzMb9y/5J++DNj1sKPbjxjJSqES0hpN0WGToFVfmEGs
F2dKBwudPcLGcgf+8IUI59HpC7wnjw86p+8M8xTG0dT5O7e7x8gAiAgmfhIzeQ9JSz/SD/K6iCZ/
OXKOopB+5zVvBQKWN2MdWREio8w0XwGusEzgz7LjHGoeInbRjOv8WIeSL+I5dSpOmb4rmtL8NX3h
UoHdL5lpy9KyjlJ+BkQ0tfEE1zxR9v+vBpY7Z65ACJlZBbkZ5uTiANI9r/Ca1HsYx/rmsKR0alnP
R8hrsREeFI8WNRd+OBV2iP5x+PvLtZBNNb+1Ff7ce5HGEbbKKqoyt17HT9C1axHEXgkDfdRZuQDo
xLcbX3KiL2/38SY2ldBUU3o+KdfKbwHxSVs/gwYXpCQanVCrUKzEkw0jaeeTgyNyORqDF6VEwd5Q
EkTodS6lIBRzhCsXIaj6adNDml1PyyOyO+BqVdILh6R0nK0UxocBFcWyqWWce+4yORr53jMRX0tw
xQgLIqH2tMDmjzIw/KZ1KNLDaPl+9gT00Xlyr0KTe9ek1ypm/y8BJVLBzyj8crF8Tnd3RBi9SBc5
IioNcUIu/jU5BiQQRxz/5/et1Zazqzn1QlIxk9KJOoCXqLXXDD2z++7ZQY/Ssz9D1b8OZMTr03sV
7cJPRNjd8Z2StL1PLrKeOqWTQfsHReqb5OhzZTnlSaHMZoEBOWpf0S5VZq7C7XzsdQLohBAABHy4
L7nLQWmDUUjv9+V9tAHqhxLmm0RU+ye8dWRjmaIB0MViiKQxaJb+CdpcVo5bxLN6PD1JDzA9PEjt
xyZ4zKbJ3lsPMxflUFMVZuzjhmjE/nOvwHODBLc4y7/gkvi0/OI2M+VlUSW2vzWd1M/SvEqjEpqv
zvEeymgNthKpmcFxJw2v2Xv+kKX1VrkCaLQFE1SDnd2QuwCAdy9GsuB919VcMCtsm2WptMpUBlsW
OqxhnfGwYSjs7FWJk3ZNXW9z0t1mk6p1V3ahkwUg3c081Xoevnpcw+zv4HCWkyO4h48OQs1b1Yns
ONn3wZZmO0LMspvxc43JMpD5HTGzZ7R8q2FON8nr6WhNxpykgXMmzXi639tgxTWf+fM9dSlwOeqo
G6MI94+SosUxDF6BFyyrtNyqg5Ib+YQCiCUOfvezf5fJuVQiEUT+z+6od1dWw/ui1jukw+nEzgV+
VHw5v/ZTtROZf7BGWpATO9UqxJpaoumGixz4BJHC+ToyoBUh2smkM6aFtIax+z2Wf4C3Po1mwnrK
95ujYF/yVCXtkzjH37v41GhyD4q4P68U0v3kpn1tIXSfc0xa67NvHxKPMau/Vemop+G7GK84xiQ3
EF9NsCNNZTmSb5gX4X4I8OQeEMHz04feQS99jz/9hiirUzoih39AzxUDXj8HVc8mWlm8TVUIg5Tx
zZPQGsuNDYY3dj8QOzWF3saxiWpC+Xj3Ye9F7a5mI6MKeMKE0TOj2rTHVbT4MBoEP4VswGMz8MND
zDA4KGhbBb19P+UUT+Yo+ik4Kn000WqobJXNA9q9EfUH7es08/dne5bugLgrSMY+rCeS+rjz/hIO
Zc2F0yefqaMrEGfy1Tl8jRSWk09d6tBe8OwJMpveEXAr1XliAkjAz5PCqFnGracG0qpf2Jw4tTW2
+D+gARpvlZWihPYobwu2eKASe34utpZU4V1oUIa3CP/3MyJs7J/fl0e6CyjqoSRry1Sp15l9ZH9S
AjQZzXe4He8xVIl9kQKirv3nYFNhACvh4chgb70jCrv7Cf5VXuEcYiLQFpl46fSVXIHme6Afqe6t
1QpUFkHHXkxzjt4TmohNjY2a8bXRPMURN4sEH9h6z1LhV8jki+v9IpRgqXPYDsXWzYGDD4iOXJmf
Bu2Lj/BNDFPVtSMaN9S0E1EDIFYvq64bcZ+filJNtIrR0PjMoCTzzoXob9iTaT2CvgGdohPSCyUf
7Q8Dif04eUwRVk4P7eMLYPn6KFFWLyHYIBip3+r5693jbqJYu16sdfyovNwr35DdV37ODQchkQEs
biHMvz0ivPCwTR1Bc1pxUb9EjHk464IvTu3ebt7/gFN75cBhDR99vdGpnT/N8OmgwDAMuaWiDBcn
8DhcRExYvQiylDVPgTIczR/+YHZsthHASzaFibYS05FmPF+Tv8bWLgY1BmzploDLFKeqw+wRolAj
yCD/w2Kc0q/R7n8OdZUS6hgNN7khherlOna6YsFrzphW6/ZcU+n6dfHwTmLEgZO+Qvxj8mqOdeS9
skOVdCiu8IO5TvZcAaEfmPVSn42Tn6WgaG3u3dA2KxkLmgkf4bZAuyCGWcq/KNvdAc27QhaeyCAx
CsuFjhAKLmylGz/L9LMXsjH3ccNuqB6jFo1ZWxm2ND3BW0urf75V7CADBVocNzSb/XSIHpc0eOjE
aTDJKKS9GsqQ6IIefx5QIFozZwGn/qKawPQ1eBmCBOzA6rSLFxAF3B59MUPytUlg/UHQyT48RmE8
SBUPjevW42guZkVpyDcf8o4XoIpV8RGDaF1+DFsd7qqSkHzCJGHPx0UMvZYU7T0oSG09keN98eV/
6/7rWHG/SVo1mMP8MlIJ1FCbgP97ZSyfHTLEnbn5gkI7tZbx5rSn4rN2mg7NxUK/cjkhEd3DWu8/
hcLzC2YKNTAS4NaexFIiZBuF2yxqEUf1GjONTdu5BgNK4pyr3BZ4shL2uo9HCydiXcO4fI31QWEK
M0uHxN1iKuNgX9lf4oetKnFJiaYqLgooBQr/5GyrH0AC8IUGhgJx4LFsECtTu/F3+liDI3w0vwhF
5zmrHQ8YDnUu6/4tEVY0tNyKWgV3DYUMb369CShRsya2cQiTSSvtBxAqTp0zOBatRJAR7AFn3lO8
mfGEXhitlHz56ZLK2sMPBBNJNUZKW1FjOiXww9lZmR2NC3ySDzyC5yDbkX+lZqHtduPxbJ5pB0oL
7GN1KtG/89XjGWR0fBz5Ovkvk+s3fxZFz+36pqiUi19I9OuMQAJsJikg44eWMhdevWOBWepSRyFQ
fuhMKEs81R2N7C89j8wL0wtVZ4xoiq3V88NFoKairqjnCRWisY+5/o40jGlzrk27WwBcJnVnwV+6
Y7VUElOVWJ5FtpzEPygDodeSYjMwnZg48QREU18evjm2xpgqmiB22KbB30nFn8xPOlhMO9pTHIap
OmHeU11nLulsNEqs925D97FjpJGYCyMASpKurf4SwxwlKaSRjtQ1VIqZBILoxtD+Tz975DwSFQ/Y
gdwigI6M+aSkiTO1OI7EL3dHqOslEYW4b1+2lqGeYyT3abFpETaupW7eO8tf2RUwK7Hb1HxvN7Tg
e5WmPHq8w2VPOFiX3bxcCSMiRofN7OlYbaWH10NF8yie4lBz0o0bzI0P3meHPofU29uiLpVH60ZZ
M+sNriQ5r0f3h2n5hbCKyZZse+L3ncU6wfFz98hToY4swfTbSyVpTlvh/3/vtwxYp9KbSHLeje+y
fZGWOBbyRH/eMGUn7RmpRs6lVhFIq7Zi/H84tZI+YCt7nVRYOraXvA2lSUtrRiVddOJBco4ApM5x
MCijH+n65C5JRSzUP0QoJtGcuSWSnW4YzbpBbAETd29gBrzREZ1327mT9YeqIWcBIKV2sGcPvljf
oZDf4KwMMVJyA/+Th3dDLjFn0nqR2IbgAEyxcbDP3yCKNNL/qKj3T/ohVfmSMDWh6w7VxvJOsQAp
udSPHHVvM50ZZsJH/J92ANun3L7UhAkIsvXBcafVEKSU8CP+0EFcADsSOvpVKZITsIAEH+jQtmel
6Qg8Lzjz8KpIrHSuCMjeK41BUnynx0dEEvicEaGIewpxskbkOSQOftCXDbyWnQaGf59eCBEDBeI8
quMaiMT2VOHltz7w7CRyQVDQf8uya7qf/vGaGEhuZnVo7GRjyRweJBYvVO9fT1pe4A+B/i2bCOUU
QPXVmYB9D5i/6N+box3ym1FTANXw3CO7LvyP1yT5fmI2IXBsdAVkv3zcLKBi8V/b3mjK3U5TsSu6
sQ2UT2vRg+o3lSbQ40QouThi3rF6emwNdAttQyths3xynJSj77IOUNwBLjThm1CDVvIByD+U9p7x
y1l93nkVI4mjt9JLxOo94mQ/M9GfHkHcd76SNXMNIFS7rzmNoF20im7topRMglKH0ozNVVOpc51m
L7HsiytoSaIBdG4gEfViCr9d3IK+h0Na/8/4753GE+OVy66J9cz6pZ91M62NXWmJwL75fDdsXKV2
C1L0ANQFcWlyUmhUJFAuwS9ER5KtH13lFjJM24lLSAxzujjdhU7paIlcB99mxT1Qilt8kdGHzHo0
5leIJMuDYkVnt8XMG/9pWr6ikHRjBoMsQy9JX/EgsY2clolIM0QO0cltlxDpym64ieFCFDxP9Bw5
rl3i8Eq8q65p6YJTDSPeHEGw0ujbc5yuysZSYVim44UbG7ROlbPzAAY6dLgJUYvUk6hqYf6ILfxl
UtjPx3cHCkUaregNgGuXohvGhyot992YddOAmSRAhIm/Hmw8q/Q68Ieiav+Wy18gjRfB9IjSMXWo
7ejwNVJXXUKpHOggY0SFFHh9m41QG05vR/KguI0qMPRz+fni5Hyl7jn4d/r2tMRe2TvcbqGoinkS
t6f3i583f1s3wbPO9+pSEWoS9sv9fh8aVlxV4O07Fh6f7ebh3kARTzcioqqL6K6HGPFFfjeDVpgH
njKp5NqIwhs0bpggVQZq3mjDyNCxLN6jKwkA/TiJLgzOdXA5+FxQJewEMcZ0e1zZbIJZlt8N4Oid
KBiU1LPPhyrLaVkSpdTcBQ2NryP5gikJvitkSFsYHNxedzbH8Z8KLxrA4OJoNauWzZX0f4iM8nC7
d9IigxetcwQXynu564Ow8KW3KtaTma3N/MjROQyW0rYw49Cu78gBnaZkzLMIln6Bvm5IsGburoxl
vBr48+tEXFvBNy9ntBywSLng13hdGVUPKqRD5fRO4rPt0Zz4Y34mUZ5ErjF6i/AbSAiVxxOxEGC/
hRaPc6xv5q7ZXWaErDlalo8WXrABwaJwGm5NKsFn4KnyGOxyw5KuzsXGyuXVGh6FNn0La1HWuZRA
708D0/1YUCsLGEHodzb0e+88wp5TeUpTto8XwV/OjEmeGuXch773AU5GgdYGD5KhEKJYjN642L0+
IBqWjPQAUpWQDPuyBsH1k6goZIyKQmFlqtQYyA3rvw0PQMN4Od2IGgTWdvigYykaKw5ArU0N+ggM
7Yfl2zeVVTU5umvVTh2haP+WR/sSlHLbDsPNu+l4wI/pVoGwE28fdwzcKCC4Io4j5vifj/j6ZlaJ
2WejUbidrWsBNqMFk5ltBcw1mPVSqeaETue2PTaSTIdoz51mKA650e0uwNyKwO1Q8ZFSjMjYyRED
Fz3vJPXfcVAAVESuISmTkflkqJYASVFdKWQ8OjNemrf9B7LesNzhoZ9PNwIbdNM4L0Afe/a5GG3j
VIBuR4eqqP+GJH3AFzFMOnJ3Gf5IGx7uNFpl0A8fhC27SAKiUmWNEvNVyW15C+8TzRuf93295nMH
pKakHq/EZT7D4PZN5RmgCxzbkh/WonJddXGz2zSi5yJSya3vwIauOhHezsoMKPBb8+ubwfRZYcUe
GMlGD4dsnYEAd6tKt/4VlD+CSgi51wWUU8spREkE39r4tFZ7xOspEQwuxJ8unUpi/asakyY/ayJw
WlabQM342UGc34aDphy3+yy//o123rAlGJ5z42kRxLzPAkwMqHXK/Iz8OhJYr7P6GuKkmZu24RdV
NpfpdX6jV0pQSlJoNajm8kkGoBqON4ZgwNDGHzD81EpFS5QbC1htTqpkxhYnFwvAuJlHCHGnCf21
SSta9YWFMcFZH84gZDdlaOhFHERGlgIuSrhslz3eBanwWWMY9CUPaKWKZ7N8ZeNA73mAa0Qn5N9Q
1X3IXQwWAomUUBFwYYrSzxjwHbB/7dl4sHXgaQWSV6wbr8xRjfZQTDEC7McNlrfogfv/RrvpCGox
hORTtYyYUb/RUvaetenNNf3VR+eGoAsXUuTM8B1f3tLnxHF9gk6T0dajcFOUwOZihnySN0RYY7R4
tVKd++i8Jox/gvvDIKY2a83paU5+XLLw7ahFLlGw1aTrXBYJp3sS6HUgBNDomZHNBsHp9K5tU5jO
GGXpDkg4QGvGT+spEsp7QhPJnug0bV8rR7+uiXKAimnGdw6iBtMgnKUM7MfT+2K/Vj69PYyNVTt+
tsP4QXRQSMfPZ77pJB+GBizXdXeJVdZ3XMx2deWU4sRI5duq/8PsCgeyhSm4j4AYi+bqeMOqDdIR
ZOpei7EFsfuR0978AQZ3gfi7PPd2HZmUYYGYHKljrhuT8ONmTAJnRF/zom9uGpUjHPVjz66aI9ix
z02txGukf/vlOE5Z5EYsjTSb1k6VrlZcIFEBgTOrFu48NgGCMg+KHYd4ihjc/ZG1teyXk9pk3exv
kL2FhBQqx4y087LDDLAG6/1qrUVFWqvHEIeeBvFmRZ4RXJtQ02jtY4qPBzjvcadxv6uB4PFJkEP/
Zgvg1lBLZPHiNe0BWSqfsABWKHNYXIQsBQZrpPL9+jLdaObdeVSTYLiU34kEVYsqQU/Zt2EyDslO
DY2JdRczJXx88NpPbs/lvG0ylSid5NltxQ3DUpOitga0nFRDul7Y6dkuyWzOAMxT1RPYLbXEYpCh
nqJu0mxFSOY+qC3QCvPgFbFfyB+NJpVCuM9imVgojtNS4aWhQU/bCoX88eRE1N7U8bt0VOTnIoed
UwGP/QrQAc1CHgjrcQpr1+mBRymRfFo84H6tewraH0AvZejKfkGr4vNJZbTu/d2GLjOtLgJP9xoR
X4vYBHvTYd368Nm+LqOuBvqfVP53GYZgq97xRHCk5IvUmbRClar5nppTwJcI3+uPx9x+BV/jgdz1
GQH9yI+VXrS1imC1UW6YT6AvFdaXvz9zNPmZaklFHBIARBWGSgl2zrdC3A0t04PsXahW0M39tb0n
0CJAEL6ri0Ldz2wiePYtxLtBLW8vtVXRK8hweXUw+cGBvFkoFrZJN+IYRrzjIYOh1R2srh0lSXBV
J9k1dYnMD+Oapei6bHkGhN6LTO2oNlNihgZrDCb6LD5v4N1gFzbzChMylv2dfKX+MSVTAVaGNyBv
+Vxe+2sw9eAOKr54Mu2WnSK+85luwNCBec8XIoyfqs9ckwu4kZ/KWcGNXC9xKwi5hwPfLOvrFRiW
QDQ8OfLj0007SdkPAcd1dmd/0Ku/1v0p8F5uhpv0UPCalLWgIMiAkIUn60B1G5zgay4ka4GnXZxx
s66JLAf7VYXJPoV7OF7pNhDBJCVfpDC5cibp+KGR6iEWFxGHjOvMqO/6pknmXXnfTNIPITt9Ybip
6iIN8bWGFBXDsNQByTFdNNb5heGFrauTwC69fNoU/ffyxIM9ctjntKe7oomd3B7CCSvSUBAk75ZF
17s5UuT1zn/V22XAjhDWzkeGDf48eVvgPKw8XG1x2f9IiL/XL3rYE/TlNior2kJPdhoA+dZbPiaJ
IajqOqEeGqOJeHPOIFfrMEKlwhsA0eJE+cJ8PV1SuJz/gGO+zxqKM+xq5qe4cOrsaxKXlWBm9bS7
FSMPpFATr629z/8f/NTXfTnrNMUeN1KBo6R2mhbol1kQr+wsJZ2gRTphlhl2XZihVCqX7X19KMt8
4agAW9WJAvZg9j+Q2Uw+orb+45xbV7pD7yLSBJmY7qAc89IZW5qb0kC0UbNywvXYvW61oMP5O81F
ripPMskAp+H4neO4l0l7+cFs/ttHERwKzu6WjXTAq/6s5X1E1BRWLqei+SxyY/b2syxQXCVsTw4G
AqQuMaO59V/Arz5LHYW9JxxGGMCjuDUQAXzHsAu3bSkTPkDzIluvbq6EwPhtFdc+wZpsCPqZ7ouZ
dUBB2RXRIxI69L6N+s5MdeP3TeEK5ggKg6e+vViRcrqP3PelM0JO+LH9Z6v153paE4O1p5gPmviE
HlfoicwU3b9uMZNM251owrSSd4napXXQ5eLJE05FQlMqbeFNEx6GfKRxy2kExCe0GlioZnNPk1M6
QiMnM4B8MPFEbSZQbhgNoNdV5txtFxrG+E8UrKwBwb4IpgnTwTOZAQZ+hpa15qj+/lxZeTOILiV2
/pSINtBNQduaoJ8k4gzS1Bm2TrxPMXTG7MkLP2CFLAozBO5nutRF9qV5a3Tmu0LTLFEgko0k36Lf
kfxgoF5rvtchcO+JWBB0LYUEXX64SjfoRHnGotbDkg8c+epwsNibMhaCaSbMvFG6m0R0XsZRYfJq
bRGcO7BBbAiFdSy3GZlhMY1vEN8dSHyrwI2XA/ejgeqoO2H9kZWGZb7Fo4K57bEYr0tSMlcQ3xZj
cxt3Sxl2o9l4X7YzJLGNpKc4B/NN9mAHIIqdnvfsccLAFHD1Ztg+4HqxvxOpgILFljX1mKJzWbKB
+3zkeCF2r+S2o8ejixp9ULkdtHYgI38Wmc3nJL/5r325FAiFWHNS8ubM/FxnetZMhZutS3fnBEYX
xivWn0Fojj8Tdw6sfhe7k1kosZU5gVKorAjwJKpnzh/0ys7qrtsrEYdFmHJaMZ1sQyLept9I0JaW
plPFqTLXf3ojCsEU1mOyyYklhBm6vEKvSMizSYlAnXf3D9klGjqR4CR/ZazVmhZykfkEj1hjiQQf
5q0D/gMN3a+a67EydmV7PlZYyn5wSYrLCu7kOAZbOj1CCnKxkAgYF1AQBI4Igv6VT4kWsF3ysm3r
LyKj/kEEM/YUu5M+yabDuTJCX7YvBOow64z0hDUVfEI32PnOjcK/u008WUuzOEtzjx35Jld/4Rc/
ll2AfHvkxsAe0kKoewzGaLf0S+iwjk07nCobxn18T69N/bE7x1FhdPX1nyclGaD7E3iM06N/JvGg
aEA6YYXXjLdhnyiLORyefBJWc01zkq5PWcfmiCgUrmadprKin/FKP67sFsTqbMbpUqJF8BBCJArR
gaRv0jlvt9JAtO3ZPeYurRdj6srWp8HES99lU+Ef6HehWTGFX/ipdVy3tBHA9+KbNxVDcFk0OhRC
Ok3E0CbvOIeOgvl3SHYVloH84XqmFsSaC9KnosyHRXPyCm6rfHxmouWHEWom77lsJGHow9rJG9fN
bkaCbx0m13ojylKwVYAj8p7GuW8iGABQGWW/PAOMBjMl+gdU/xJ7FeBjcKdAkCSBqTw7/AtKGyNI
OEziaXtIpS1WPZaalEmzOp7PqrEMGf2YG64mgtmty9fWV1H/200J45U4v708+2UQv0LWbn3BgnPd
9vrmLiUy/3fB7RGeALYvmLmUSZndmNGlmMRMhTptkWGtVc5DQ2IUG+L9TDfpffi+XM6QegIs56kP
Zzs3huNEzD2OQBu0y5z3CUzeS9GcEWKRBRTqm3e0RN2dc1ZxROUO//77iRF0A6QA6kfSo+eMK30l
SO3AKHZGviqJkRmPTcBT1YfOrP1JRsdcYI/tOC15dR8es6ETeH1qm+tYenv23i/97V4sdodB2vVv
gU9BqkonV5RQAJosfH2UI6E+9LwhfLyWxx/5ZP10/BCJXSjKos8jA1248Ybxs7Ld+RsxnOFWhxv2
9P037OYJfogxl2SbjFSpnEgaBICOycsaWHYJYrDmFF0vRfhL6vLbDYHsqqf14Z7+VEreKrE67Hmy
dkpzINyiwLnAYIz9VMJhv9OYF6/kk6HY0/JS3xUoeUvD7mUuj/4gLWbezPSz4AJ3qIK9F89V+ier
eUCB5aOhhuTZygEEnDL+J9WexC54eq438c/XGF/ISF6qj81J9DQB4Wx/05edJL9M04QRbrSIPAJm
D29LCx1jmrbSSMxaujoYSDnPbJ642BMG40dsW9+fA1IaQf9c+gEfoJoVg7IkqP1zVL9TLAy0neNH
e3L4KxhMiF66Q9tbgrhgf0KV9AUoI7fsCp2vuRgxnkgdCHclj8vxnWBQ6POmYlKg70O2Ido3kSNd
K/x+M+jNSm1I4+Mi3kBfcEAwRRW75OYOEeT2Gq0a/2nRKmV3G99qeCZDWdSOwHELUvkOOClTQ0qt
iqgMdXyhD8cub+SDkk5NKljFxGszbv1drwlnSiUufv8pSV3d/I2ul8cqS3qBsMLWGSR+PeYpo8df
o6ISmRbdlzaELRB95sZPkip9cjV9ERfQDeQJCnUQsJPo/OVtUSst3bpYM35+d3mWPFKZ2a3qNBPI
kHs7hi2k4SeyBqdgt5HqsOM28JhnhFskBlJkYwb8NuBlVO8+vgChF3Vb8SlojFU0fgaUIUwlW2Zn
uxw4E4GMGgma5bX8/zN3Lm35dIuhA9X98of6oTWck93Blg1hY1ed/QeE2WjMttbYAkdb4KPpy9Cu
BXt9Z5zIXwpGxpmRq8P4O9g/T1R/Q4FhD/CLXXPKrzTvB0U0flQnHorONBbxUFEZMHxRgxv7gpXJ
B07mxPWwTg2el+DOZ3ZKGsWrueJY5xCEGMUV8Vxe+O7hS7w5SwB+OIO5T12bnG5QaMg5Kb26HPHe
8qTym8A8AOmaWs7m17r9JJ3Ffg7oYYSxU5U4Ew19GRW5o1+gQjJ3EL2Msa6obA4d/o3UujPWlbDm
4aG7iMztUK1U3cjEoZegLbmiJLQ9I7PlYAoydDI+ayMBFGaJ3kBLKZib+D6H9KzW8cmWumNBdWcb
ZCzGQXChGyr/DyPuuo9Az+Oglg3yohgrkn2I5gkQDbXutzLXNwN7PiyfenPcEV5d3GeQ6UR/wt/e
eyR2x0wtzhve6fxsKeuqi4OgbFLbuR0y9w2UvfJiH1fpscqzMB4CHW/c2MQjDLvQGZU3jMH+7sqb
1VGbznPTRHloZf1/bduQUMtUGA4r4S7h/BJCKQnCaXpxCMJnhtZMfc/iIM6v+u+rpelIhwHgjDBv
vs3n4nhOChCanStCiz8jW9spcPWm4e7ftQ6eG9/lqODMwW0JibbC0JG+y9VMpbk5FgitZa0/dAmx
oUFiVTCg4rbabG6sAtUGS9v5qFNjaNAZGiqHPlzFekceqlgpskgJgQXZSH+uVDRP486jme4yL1al
Lkf5PQxgirtWBGFETxMtI5oq9PABiDESTZJ/ysXLq8SHR2B/fFhqrgPeeBXQXwx19fBOhcNx6BfQ
S0omTzTjFJvbuILFaV2rFUChpUmR/O4W2fngu27JmGhGI7qBTUaSlU3RVtCzSZU9jAVYI0Uq0bz/
ByrefOvIujeZ5kaou3aqAJ1mGTSidpecqFUlwMOipHXItPxMo26mgS9JTOreJg1PvbHWs017mhie
einvA3W/PyzIawgSCj84AgbpV43+eKU9BwEJF2AxXG42Ism8TM0QlYNzhHZh4yXkVPtUQ3365pk3
piP8Z3xllpEJ/AALj+C1FQyOeXHbEI7uZXK7HwPI//ctiqUc3pHpSV6ClhsUc3KW3Rysp1+E4C82
IgHCEYwZB31MDQhcZirjuDiLl3zE6TMKh6hfyVohTd9ap402K2zdC6oa1cU2WxhiDAsjEp5qtXIZ
9s0uQgi7MsDT0YWqbuzKJs8mFE28MIWKTcmjja/wYVokp4l7pM2U0PZHBTNT15OLVscgfLH3KAOU
VlKbJkjKdEy8fd0Dhb7Lpu/ujcFdbujAaKppX8FmGELV1l9b6fPkv53SzDxB5n1xMSQR8R4keAE8
yQ6E+/93xODyoIWHt+GSjDDbHgb7AQmtRHTWEERO555sBy5fJas4ijvdOoC4J2IeiLVPxUv4rXNc
4fUuYGg5de3/qWR+tLpxecydFu1qJgL0j0Bhd1YtX0AuEmYl6lSZlENxRXi9Tr5NGodwjDe+3+eU
PQcE+XHWcj0NulBeIuIggCTnYzGpbX9m/gyU5Fy4n7/ZY91wOANRA4oo+Bmq2k5lRKlBH0LV/KYV
Hrzp3vBswezAssDLAQC8U2wdyuQEIr2BxEfuW7SkuCm10I6RPnjxWLHvrgvJh76ctAbM/IR4a2T7
gFNYe6/wTDbpUVq8h8zjtou2WlUcMiFUWt47o6Ss4Ts2u0wACjJ8AxbEVabJai1Cw/0erq6hi8N6
LWBFUtQl04A/SfY0Tznx7hNzC2gs3+UrdDGQZ0xeqM0SOsCfuI2dJnyq6mR/8E0kL+P2Xg2If2Um
fgtKjdi9g/KHapDGbMQEIQutldHcrzyiibJfi5oF4hl6mt8uxPcWKn7tddQmZ0rlKosa7DnhZ3tR
6sPELS1ueE9MpK1Ng+UW8jMu1aHo/2/jrzdWkyS+/jb/1AcuyLiTsuqshfznqz9qWmOnGQcMii9Q
CcXr4FCOFMZwN8MLMYCvsMHYOe3V23MKuATzhYyE2K4tf1rJNJQ+9GfXCxKJbaxdAMtzPmNCPh+J
5H+2yPcJt/GfP2G3JzOU7bYHnLkFo34rdluuBL8TaxOuHCzrHxxmf962WK/4zBfdEzIyJAIZUPH2
dBHtz0vnj16ENUXy9nXbkkn8/M4Y2NRYEbSjoccl5dKgFe5eRvUHZXr/AUc0IpE3G7HnLxjTd3fu
LshCjY5TcemL+UKavII3W9UGB/OaRj45lsWDZV0SxNmK8khS55GRefLSSCN1TsxmBIqnBqiGLoAc
RlTLBje5+UPdpF12+WRM+oJ8iF+k1GofetF55onif9cKgTEb2BwkzMlByeUR8AEwfvCIhmERc/t0
rGPQIeHItUsOxJZljfUoHai+0wHCCQ8LUjs3WHM1r1y0x4CVmWu+7nN4PbgIFXBj1koQv6TjAYBz
EknKhxRJ+r/vIoYDF8PGme6ntTclZLHKl1x7NtBdr5BRU5DXhMl9mVoDzL+ksNwitL0rIyAbXAmz
XcInnyHq+YTQa3lb52RbF0/erYac8MkeTGGZD55RDzfqTdPBvCRyV5XJS12cxMblnZCQU4KShu3z
agfmHXnoeYIugeEnDDXB4yzxgv3iANNHVlOA6rotssKY0LO5cz1RKRG822LIAKLnjxCF6PYMSV+8
07CCJhvaTSK5rkqcSsDZ9W/CKd2ZhxOO7NJfckEZtk2Y2NZXXgln2bszSAhvR9Onk1wcJeJCO7BW
OAd6uX7WygXDtqRLwku5xwZABiF4VBEzTQcKLg9od4Ep7bikTjUoPaSiJ3oA4pJOs9pln0GhXnr2
YWWMlh/9tcFldxmfOtTDD9XmxdVyQrSP+aE9fHN1xynEpATASQDCLxvdvoKYLqoMNFg19AQzFXGB
MDhdtTrYPTDSy1Nr3+ScsIvZHOAJAt2auBc+dqfta+mSRxXRRJ3B6+ofH6fCdXXRUimHRW191ehb
bncmmxIlVkiiYHkmPDKKlWhMiQUi5lmXRnWdUo8oxcZrzBYJuqrkRNFcblTojuAmr3CGxo4TDjMe
1/TrnEjd+B0JijRsig1xCtlUVf4fadfFkuVRfXbavNJake4zKrFRqBdJygLsrKCZG/fF9j13Oges
xAb3bVFLQA7WMkmfkFAwzecFPVAW+z0d6+SazD/l2V/NlD4w/5QHx0BG4ExZEypb7mAQSihZJIpO
7EzXjxY+LbKtzucCvLgWsPSAHaqMrSyc+0cEqaUQh1tw0UQI++ivGIa/cRiMU4sbgOBd2cTKgZ5r
Y6PV/DfnCdlHo/B+9wf/qy02550O74ItsBmSZhbtAPAu5ckoCF3i4V9QgqgSu2NRroHV3cMnF31G
CsCCWbvL10+Ga+YOq2pg3kvBYVjcmPJY4jqZMI9nDd0XCVeZ2orvpQAgTTdIMXH81YOTpGlcH9Yi
jwsD5+caaJ0WQA7g7FdIc7Y0ZgDOf0WaVdmoY8JXfye8v4Iqm/mGGvWTEqw8LZzPADUmOlfoKy6S
g0OymgSOkqPvlebY2wXpO+MEoKwgVWOqNFwAzZ+ET9Ih/GFEoURjgG8qp8gwjUndWjNQeDch1aVh
Qekl491diYofI8zV52tj6UgzTk3YsoNvBG11ZUJEaklzhaeUuXsvq84n2Ne6iSTQoQhUd8nbaEkz
mWPNOAd39opIC43XC1mewC9D3T6wbLpnlw0/DPzHl8bnfuWRw4Lhn6aWhTdx+0ZCLycys1XMN8zH
9ZLGh6Uf5ZNg7hPWr/bElnWNCsxUuqIRoKHevpTBYzSj4H8BJAfpY5Ozz4AAC/rAWYEx4kbTlKir
TS8e6dXZDyUKpRu4VwAXj/bq8Im51TyNYVrM1W6At3ZztaUl1Hor5FafIEi5UjDRe6kYhF80lZoz
wXHpFCezsIGXkSsqONoWAVY8L/KQWnUz6Jc+XgW9kN6pcWfI7YRw5qWjlxlX0wNA4RvWglkapkwU
XhF7IKEIqQnS8Y0eASrE8dyMAdDdw8QRKlnfXKE0pGerCQybMRN1Wd6+iYkhFYUhVRcyaZRIP+iM
3JelcldAJXFDowt1tf/7F7VpqXEjKFLyGWMyEOUPxrFvJ9b+g21G3rnAWSUa
`protect end_protected
