`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 123680)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf+kF
201k+6QR2npVEY+494p8x3Y/iVMzNwQUtTTNrheBLY9h8bbdcsKyZaY7KuUU5K6Dirm5yCA5/cKy
fVLBS9aoQtd0++VTEa8JiZ53ivfBgt7O4dPUrWryf2eOg6vahaqyDuI7QijBHrtM0mffeC4icvET
5KSC073iVZMgw0Z2so1EQzosT66HOudBmWfbcElxS81rk1QZh5OjzgLSlSqxFjzcvu5rHGpQcO1w
qnaGuoQFnWjNoSBKSrzae7L5Ftf920LUqRwwTBzn5W+l+2DkbVEJZz+vOcY+z2jFD7aZSVSIIL1O
wK252YqFpZjDOVCgaCNjmWl+wBEtjhptK5mkqHrYNArkesBAdxwMDfhRCjabFv1GWh70PaPBrtHy
xtLHhcUEyGt7Uj8Fmi1Mn8xu3J5AduHH4kLys8MzyD4ej8sIYC5BhdMOlb3/CzY98m/4CPoSQwyu
sjIOavnwCGYLV7tPkxqjoNPcVUVBnlzeyaty8mR4fTzgT7pn8Wxz+qWAsToBbfvrc6yc3ULGX4ku
9dE8qpMOurf+tzHgL53mUigT6wTpjyH7LRseYHKs/I+f4A64mNXBs+C+wg33fvDl3yxwqkT2ylHS
f+8vkTjh4OjxEX5/khVWDowb9+oeSWkSBf4yBU+yZl1lgHPXI1ZIZFq/JuAqi0csPmmmU0/RT7BQ
su8VulrppPO/YlAIDcVi3KwVtCkmaV09z+FEup4VbeRipyEVpAB9DUNaFCyjAUcVbbvJfBU2hA8w
HKD59tiRvlwDA3gepVbAXFmrkujLlH+Nnk9ev18QubE6mC6zPq5jlIseDA0AissvrVnHro3KFS2v
ILX2Knnz2mrAqF+/AuP+pK4wC5wObPpcPfDhW9v+4Qh/+NZ3GaxrSNtd1aIP5WeTh5n/KNnyzEdq
JvW8IbWoCTAtpP72fQ5ubQmM+3KfXOWRsb5Xu7TDPcqv98ppvoHv65QPJE3xuZo+GzG88l5+rwzY
E2XAaZTXdlPaRovahkaex4mC4sueHo80tLZsZ1tHoxfyfLMWvexPlKcMrUozBrZguFUFFh1H8JmW
z1TQVNjaFSbB2iUtYLi6+jAmgI46p02Td7f9qHQ5mLtxNTVRDsm7xin92m3Zuw7FssYfS3C5CeVJ
7JWLzWONg3oX3DvDQTDMciBVFD/eXOQaLRSWHGlUcAClcE3sRjGND5xHwdAjY2dn9ZfSds6CMCpp
aHMRUs7bR+Y5x3bYi5TKR5XRBJZWQ0oYN6fvPU44XM1m9b/TiTjmDDgMPcpEs5NHbvThp5RTBTFF
fyxRkc3sBJ8sQmnDvexsmuqMF+YOcYItTvRQbUQ7InN8lFxYOBgrqCCcw4pQ/tgilsEvLlp0NUH8
lzyIqDiO11W6qDj+0TG65cgOIp5J6WDm0wh9lRHAez61adh+TsBGO34N+Wa0eULto2Bi9S8cP7iV
KzghSp41zR0YAxhhP39z5N0TEgC3bPkARRPcm9KNf8YhvMZ33qzUb65iGTTNiH429Bdg3+7W44YY
JUsGdF/N0qh76zCkeOItivpfI3qRuK64rYBQhJs5qpWKC1qhfgemW9wpuLZiO2ISTipGXEi1DtsD
BZGzbv+0eG3Hhu+BhVG+ueDD7ssTYjddtmu28zMhuPAPSGdff9v+fwDBAW4jktWT+BWp6+F1MnZi
0zUrt1GZJzUHb6T0BTKaaJS8GoASN63u7d3ceXypFY/BWQfC9G0y3j0AgC6eODj5OdkMlf/HwCDE
QrEGgBOY3qDVkwLNKIkqElL9ECuoTDqOsrCf71a5gYiyVPBVv8w3d415XWHlIg3mSyCbnMrR7ZcM
EIvNSIWsDlbbrLA47zF6C/JwQIJeZjsns+yf9HZQE41iFnhB9XOOTP3iUeP6U1IpO+AYBRhFRTif
ih6P2IqINzPQ4AkVcpJ04F8fgcRJ3j6b00Ts9jVOF1hwDeEWN4EvTDk8Wn3xGOpTDFATHiotto+R
2J4nAQFAJqUY9GF/zah0t8zAecoPynXYV1hDZ540oC0Go/Ohl2fYhLi1ONmJjKbZ+6SIGzwj4+pw
+ULkBGGKQT3NbktDjus7X1kWFzMA89LH6uSwFnqSL2o3r6nAlj4rPKvwzgl2x6uLdZnE/aT2DgLX
yWe9P8AdsgXhOQWdqlf3I40K+2/bnxLT/T41QVADtaeHw2h8sq4FYkOb4l7hqjwLik1eVW4ypnaF
x+iN/m3AcHvoiUoTR3RIfwfx9YukCYBnW15YMKn6/+0BIc5gzoAFryIayPpuNOIueIDTJNrUoerE
NhwjENn2KmulgrzcNP/DU8U2zUq83AkE3Pief3wL0mcIYb2WVKC4wgRAR1E5H0CIFy2q6Cj3tb8F
xx1cV+8hRwH6Tsu3oHaBXs2boydZf2Gp9jisG3qH2i69+p5ffs4aM6JVlu86aICxso4qcTbrxaIH
iG9zSm61JOEU/D0wiZUmIAx3wcBIsyDBoIX06XbsYmgCZnlv0w4MrBG2g4nIOyW3qRSBzryOo9xy
3f3rTjnb43onJ0z4J7TfcPCg+LWv2KA1SOQOa1Lnj2/HkAFpeeW5Xh3B65m0D4o5PCUYZwfKPYLm
x/7uucCYzenRnlPVRoSD+5YVU6VRxOd3pgMLdv0nGgfGxW3/PE3yrMdT/PuZBw5rV5l7zXog4ZCQ
tKlm1okizwuS5r3Ni20wp2MgtTE5Bbql/UErzda3ClTEHn/atSfu8OZbib3IhhLMqgsoNdvXPbXn
tT6lRL4nj3pOry6uqHJWRRquoDzUo9apJgiM7+/CG4yaJieQ9NeyI/0QpcQHzvykvD6Up0J3xPOR
uGXKX7FpVzNgH3P5hHjsW6JjKgKXKviLzLcntIaTb4plmXfXuH18oMrG1QbppJxboG+rbp8KzO6I
+UpmQ1WcvYPI0yB/5PcQ2VWpZrS3kUVRpdCJc/v+csn7fAXzl3ckdieC5ci20tPa7Er5PncqVi7f
2fD8wm0OezWs+veTNzzbqO2SOpgMp4QKZPKVsS05k5YhEY2uXPGe7bN470go0n0leFbQqyjN9vL3
Ba/0Kbi/VwQ3MSLXr9BR66apvnqF1M7+SVzxCs/slP+4ILqzCWV336TqJAU2wt0DyvbiPwZgViy/
ROTa7nUxJUyLyDw3zAVjR5HGPST5eiDZZc9KeQeDGtonnBoRFaFreqDHFd5hyhtE0u7Cdg/ZIDxo
EAqb3Subz7E0d51KhixfA/Xvd4xnuuImH+Xg/tbJHsamdC4K5WJ7iALxx0QEgkNR8TZZ/lDBr6RE
iSsD+s+6kGXCJsQu6CmvGDp8qf23sHl4H0WJEKnjpq+YlV5+SRJA+COOcsUXpC40dajJcS9lneIg
c8ofcvmWYiNnPTCIIlMUGIOpTpGZ8RvTbjeNDA8bAolY2bl4lWPPwcQ7mYVMcJqz/2VLPTbjWxWJ
XatKGhvFtYHGxTWbXrr1QrBV8+FkBvMn27WVQsgcfkcVNhEgTuS93lTECwkAETpW2ewDSjRXeC6N
2NDaDAjPCfasSzRAKbz6XJNvPXu4OcK+Yv01VAkV/tbM8G9bjMNJUX44J2R+DuKCk0W7QUot2DD/
d6eEktcFDalDUVWKq7ffubMN+Dk9UJhPkpizuHlo2QX+tg1mgl9dRII+tMduFenjHgkfUgw9g7vP
2+pn7VkIuGmgpZNyxd8/ZmJk3nutzfWKzl7xRp43KnFHC64RW+4I7Fctglb3db9xVTajTxRmOl/K
PwH2dLo2m0qBkW7oQkKw+y18iQ+bVlXzMJG3SlWmfVuLUKGP3y43sHrCPU6SGIGdCalXm8L/qOSk
1AofYqiWcS1YlmnyVTCmyet2rHzFtUdCn2sSRUEO8wL1gVWxSTofLPo+ipewNXuYUoV3jQVos+bw
iDG5UB8gLaaTQXsHUyWkz9iBMQkgC0Brs9pwxdrHkXJUbookD+PocaXu3VBJOo6PcpXCR4qs9M6w
ilxL+LP6uSRdJbUGsxypNj83/8+f+8Qlfe8ylH/WvNOZczP8dj/Kx1hxaRTleT2TV8nEh6jBrBJT
yMuGEsuwWC+Z9wdkmvroSBDGR5FG/Pves+uulyD40wg4/ViSv0t18ChjC5134DRvODB+RHn5K4Ny
ztce1Tj5XOfVoonb1cmYqjVaaduhHUQnLoIkWP4GiopbowE8puMSKAn2Lnws0N8NdLfd1ZyDh9DM
LX2ScYlU2W8rJEkflt8osA2HebkM8LEtSWUkO4QQSeebZm+uyoWuvPmaSIGqSreXMdSCTIL9sYFa
dbpNpuh243X8v7dORSz8rlDTo6n0vyu7Ds7sGpbMFdlb6GMZYpp4M5DCn4j51EXg6yU2dcrUXwxF
xdLA4QPxDte2Ygo9XF7xjmdDZs7R4OCU7YdTspbXJ8ufALqmQ4+3RVSP9ShGzYZuivy22C0HlWx0
Gad5vyy4J2L/qWcunN0yYjKJrknw25ZVTLTVcObo/MNNfanmyqoitBGP82d/brSn4pOp5hsgiwEe
/czDKUZJ1FSkEhT9iOsTovFvHRS0Kj3K72R4T0gndqkaSp553CkuEJ3eyzchmOo+qijfunw7QIXA
BLeyfR3qBc2tz7Qz2F36mpiqKN4wzDoPfzMAeYfLR3qMB5EOMvAnXwEzLZEBsW71wja66ctxhiiY
/NwtBU3bbeU/hyD2Nu3FEsnjrTC9Itj5VH91ceHCajTwj+RTokjjs9Wu8xHpTFflRMOU3puFV2Ua
Hsa+/IDQawQncifo/J10auJYVcBLJJncAIXwInLQKRCCbOZPvXnGXhCj/sYHkKcx5l+8pLWvx5IQ
lW6OWI6nDxyTZ8Cs4hKO37rSZa7GyDtKrrdMgTV45wxqpCXBroiHxjvfbqqLk+jZ2tsqmhW2dzp4
YiV7+jZeBW42BspzntLgpkgvHX7d3MtpWn0BmuI/rH/IM9x+CPV0igDLkCCxlIld1xOl4CKT/NYQ
uopYPOe1cXpZJ80eZHaZ09JYX4nEboyrI7MH6NdARGdDzOpg/g3QMh4TZlKQU9p8fR8M5AVRkwTU
eSjFm/jPCq3CsvM0fef7DO2zKVNu4zwlzT946V2TulKAp3cKa+luFKCpVkwFZLquxpXDLMMkslbZ
FAnHBgZFEBZPhTEoxNW5AjVsX5eg70r+KuWLfJ6ARIe7Gm9a50PEM6n6LfJDZdOrxdbFr9gWtisZ
v3uGlig27kPEwCWrmYunyeIock1EDUrnJOlVbD1yThkDfMIOgVjeSWKtUnvJ6FwwHYaCIbihxrK9
Nua9+1TdX3Dw1OqkeS81C7oe6zumFPDJwzvBocZ8nmswjpdvjOkodMydqVV1qMMp4B26Pk0/+JNA
JhNDQV4didONJhgVM+xb3Cn51E5tzXmuoOwE7Fzn9EqoWEZaE/ameQDWPhTkAjL7mQzeXuCsqcQY
rZq13nHTnZmeQ3/V90NBF7c3Ihz1V4bdAbKFyRUK3WvO6t27oD9UMEBymQftkTO/IUObhmRaZpHU
x+FdAivCWi8579KWCemYF8mTCRlVYGv7thbM3HZZacLln4lneG6zRXNDzTbEiBmsshhQE57aUT+h
EZRZA3Lm1ehrwyQZPpy2zw09EAU7sFdMd06LhRWQ08+R6I4omjJ0NwsA6OL3iwgt1qryvV7dMyix
hqzPtl/uS8owx/agFLNA0Xij2Vr2vE22ByDf2dOpTEiF0GcS41w3Q2wtwld/R1h1RPs/W9F/7+59
7dAc0Y2IrOZTDiEtb9wOBKyjQSUmAI1j3eqaR9ryvbKoxxRgu/61Degs2MVIf53IYOoCSY4KiDCP
8U81M5/NjKMZvThabQbSxLJxBUJGSpLX1rHwxpOdSmauUMe31GSl2A2WJHB5XRgODve6qI2+vTAF
GDfWcwo2wCmQZ2TmG9ZN8hSuFlC9oCLSpsrECTawzjJ86f4vNE/gF8o45vVz5Dtvv3ZCkog0Fyvn
utyEq7rpZ+cYoKay1z9BiuFheIswf/7//7hUqEm8AMWxEx1qGp4RVkzMH/kt17WlqrPYWW3D38tX
oXO4/wCKC9lWJibAqjyTB/6KN/YUplISB57ThZmL3nICw9gxiSuuEl8INPkR7bnjtEMChEfSvXPP
q1breAxllXEMtJFxFFm1FP+6mPoxeDsYQE9IEhhmFaTGZ4v6C8oJsaRhyMpn7a5EPjKIoSR3Fewf
u98zwTLAkLonw3ymRBf6ZJ7OvAYsjg8jdWKFtPHO5dFSgkk0CG0gsjNpCa5wsEiUYzt48idmPBNg
SH3UhT3/XIpqkvP6kkGQNwQKt42D/s0be14CvcIG+lvXhErWyHGFNApJ0dWu6bjwfKN35AuyD3Sn
7p32K30DyuioIIuMBFPknnfrH1NZD1eI8db1RvrqcYN3FFjz2hdSer3J8Iz5hE0BznTisJScup09
9XDjY9kvYHqEsdtYI9dCTCNCEo3CEUThqKEW2DM372C1XQZwREVfMhtw7vCIzWtgDa9YekjaTq/O
LLg9mniA5h2SargK8FKqbVEAfkm8wbu7afyvCzrVYL9tY3eDfbv9hm5F6GTyYB6oQPmZfoxISiyz
PIOgf7lat9Mt9MXegEyE88spQXA+Cl3A8i7V26hXRzB8ZU8QXngi8ZKhIKaGBrZpjuKDEHPcgzRm
yZypvSExHs7TEfBsU0l/vUn9yaH2cfagGXY+FYM4LFtRYngs3U9vJLElVuW6kpT/SwHTcnNpaPvZ
3MGgVeS6FwdgdNOyePj3sC/IEVfjGxUxd7jLMQWvcG2yfFELOH5K2F2mM87EKpPkYVcujzwTVQyo
5cbK3VqTqJ0KkhliiAciL7DREdCLwXvh9ROQnmmtjnpLd6akXe8D1rVU3DJQURxhtEx7AV18PgwD
lv31FRsbjUIQperoZLlnxhbs+F++weXYIMyCchobisBN2Xn7oO+JU6thqgbNhvOXBicpbSah0sx7
czAxhxlWXjteYB2qj0KpSPjy3se5LAqk9KGLxHy8kVujgokxmrwGhsJGS6CwunF0H3yLqxjZbeaV
i8bWyxV6AgFWSxf9izuaEl9VEjZWkcFFxNoozxjIWwIk0EaeV3XGZFWT5dBqOFkv5YqDyKoesxti
0R6beVzV9tUmEzYI/xh47BWgFmHmp4CLcqlgBXcm0Wfy81Xxr4/9Z3vZZl4oqk0Z2DvG3qG/+XY5
dHrZC8VBuEK48iYayktpnEAfTjjycro97SV5i9t0s+CZLY45G1n7Y0CrSNxmOqrM3xnMLM9MHnVA
CcuiaB3KXT6MwEqB/wbT8LAQHlLrss9wBznncOsUSKC/q+BBkkY1Ky7oCkyIWO+MjqqmRcZ1ZygI
r+0dytxVaxnqAd7IbcZyAVVM35a3Um2aDLv7AtRZyL9bzkejtGMZSmmhnbL6A5cB2wzOd5W3SIMK
7y6hEd0MFpaoASLA7U+ldZYkE6TuL+1xxCmV4h7bJ6hQc/dvc0EfFdzwbMDRH/jlr9x77b0E87Rz
N5QZ0db201gJ9BNj+lUbESnzRHI1UpTbpnwBORhclRpjOCVWuSRk6u++qfgW7A836i0fioNtx8cS
AkrKes8yf2IdN1RdcW75wGoeeLucM2WiF9itYTz+GUuWWPzJYEs/pVMr3gO53rPO5r/NMKbRzXVk
kFxSfyxyjJfh1i4krmMmnzJpjZvXUy7fennjlKGG0YbFbMulvgoKvQPUIlivW3o42LZw69uc4h9i
/m9eoRM+pZ87W5aCs18+xzl+5U0yO1ZhjyZJqyoUkUpNdB/fEVBvorffgU6XdOT2TmjAmCNXeG5Y
mK9OBA39aLeyxNeRWrbk+HVZQRPgLOvLe/BhwViXte2sFWR9DmxYiEQ5NwnD+Z5kvpdKyC13LB1H
6cPFji2rqRTD1nS7O+oUDsqtTO0DBSPmPF97sSM9XG8XD3X5q3xFnfu5Ep+jg571Bc2ikdndLbCE
bpQqh3gb0Ln8KQcPzR1IPzpA4vxYn6sXL2Avi5YnDXOUceDNKIvpHOq4UWT1t4D3HeZObDPgo9B2
mrafd27CqG78r2Q4ymiFprcLYI+93xFnB2cNxAfMAOBLhrb6/JhceX+P/M+Bg2YX9/PAawHX0AnC
iPILdZNSdQ0XvW1RoS/pb7NGdBT+xrRRGm4oOcayBmJIYR2dlcmRuzB2jZOJVFc9DA7JM7mNTczJ
/Kvx3C1cyeMu719QoFEcaNsA0X1oGLAj/WPQcSAeSwQTwFKBQTNGY+12zLeI0+6IEroy3C3Xr1az
QbvDIlvD2Igee11YtqEjos00+r8KVSlOV1ioL76BU83FxQsKOVHyY8yTVpFnC6gbAjy7EFCPoEQq
YWn+N7ITGiufvN9SWDUeBEVzotQ6d5NIaeKWSXF3Krdlw2EFG0NdBxdOwB0p9hmFaHD68g5mF8gH
qOfLMSqqzH8GhqAuN5Cx31IwZVg0Lwdf8SQmSnA9VKrLuVdfPxedhkpapphnwrzemTnZakMprouN
cQgnne8AUhUa8Hq+kg3UNjW1ZvCcwUwSERVhltYqeVJyhUXmh6Xq+8qynJEG1jOV5F27OKSSEOQ1
YX4yepcrsBwoWQUNGDLDrY+nnpQQhWQzIjbXyYQ2j1ThTGO4AC2kEN84zwbuosap9XNuwknlB6RP
NtxfDcW3erz5h0Jdp7U0gq0E3u+y4wq9Qmms9BZ8gi/caqJisgqI/nrf8lxsO6f4DHUNxFVWFNvs
jWBrzyDIGgKah3b+rQu03MrxrIkxl6eAHbBWMEoGihYa3tf2JiRdzD8fGIWPBtuPG8EdcEm4kPaX
AKWLlcUVI1bQowxjKXOBHuEQSJKb5ILCxK+h3KtEtl4zPqmXEcxSDvoCTcJA3uJABWVF6/1zRk80
aehXkrEHIfP+s1SDuRESxaF+n9h667Ax3MXjEjLt0ujg1sT1XGCOcfrhMGwIksJa8uIKjs2dDcyP
bPQTHPCq8Wb4PYGgzqlFmWQONAxIjGl7wBZs/bRa32CuwO3MiVG4+HGuOzHLuSRKSeVyUXZm2lMe
2V6FFSAvOcFFy/4+rD7ILCBGWHN69/gqL0P0eJjgAaxUXf9magju3zQTVEJAGXBH5o16boF5gFfx
R29BDo8lVEvcfTwPXZaq6keMcArUITAI9yDmyBpj45BxXxnstEZy1OoNuZmteWD3AScX1Zgp89J9
l8dNph2Q3jFGFF7N6/tOe1yVo4JZ2Fhj5vUhm3yarJzzOJrUDQH7SguRKWNzyQeH/Jgslk2vFHlP
KJvWgAI5tdR6JzgD1XAjFrhHSit5qiQAL7ilkS/wGMqd5RcOUihA4eIFtzQyDh8aIa8xZQyY7kgy
nmxXcG5U8mDXS1mzsXH+8IxrmMJtKQRypPBdNX2GPuOVk4k/V2R6dmkjpSveffpKKm3i0Z5Ct2FE
7CxD6R/ICF7vzAyMTNKt80tQMFBFgtmT3UOICNzXP8SVuCJDRpKvZ2k+2u3NalLWJOk93UBPfXC3
eTx+rrTWeb4GCMmbUNLTGD39azdhOA3Wt0AMirg16UfFIsMC8gYu1CbcOyn5+Q7+UahtAAa4XC05
z1Q2aFzyQDdTndUB6HfXi6LCmiqYCvSTlPEdtbsN+1FNl6KKjSpjSyT1mgfM7bA7W0Aqrlg1L2LH
SD4JVbOUIRy3PAvdTUGcIRso0hNEhMqF4VcGM07dyTMdSytyvIAlEq2njcp5kPoMCM3OCCVj49Pp
JkBX6KS48+7Fhk1eBQAucVrhte+SZ3rv//BDNy/qTIevWIWyG3JdinUtFW+gPKDnkG3lfL4HpI1X
XS95ujxGu93JTzm3Ruu7yOymT8ptaHQOosXYP3qgRT6u7f3SjZuYYZvhkc6sNTFz9X3kfBjUSVBL
Pawsc7clzPeDIz60l00O+Ckl3ifNvNfkUn/bilxbgETXdcLZHr82au8E+qmCZRgq1ZBaDvBSxtuL
od6x8ah7Ybet414ukjhVig7jQSck22d5XcVMuzXKW2IN7Z2dt8JzPI0IvOsLUWhFOZTigJkiMwwo
Ig+ns2j7wRWGu1Vgdrkmy/XjA+vZQWLofL0B71mzW6ZJdRgcz0ELLYLPELvQEBY4n6wrUUMzcVqw
U+WpyrNUeQXORfRJQRtCFY2KO4oX8o2K7VK8mDXWzErQUz8pcNU7hPuZCPw9/WTko/VF05KstwgF
05QrKPRZRTSaKacYXgwpqYbNftACuUDX8xEpVuAGj5DuNHdiPiTbBg1/D7+06sOlAXJwhxbwaCJL
h8vnikfB87RTlAT5s4sPiOsz6psIYkCgaKsRcNqoPo28bOGFZGvI2v1zatjIz5V0V2BhP4OLlriD
ZL+kIXT4jYDnqyCZdQjjDHv9i3qqTS9kn8sy2fF5zfcii1GAdvV3pv4Mh6qCtylY24XaI32uNkqY
X5C3i0JEE6pKw1laSDuxUvZx1zB0NR4ZZY2BA67M8mP/FgIAH/CKGkgk024+BWwx/ImwJ7p9rf0s
JDcrmsCNbYJJSzwfXQ+i9esn0Y82iWRr4zh6looOH0VR3pgXCVc/LTsfPpnmliZuNa7NNrAs/iIU
2RCsuKxaBTr+12b4RS+lyNXX7U/Xddn3U8dmiUZ5IfLtOBATlLsKKgCn4S4bzThcOJOJhT+it9hp
VYZduHBdsl/FHu9HrJ89ihcEnP8szBSV+s4241brB7u/O78moc/DLkMV3qTj3embT/Ygalb7e6Is
207MFAsyGuIbQEX+A9zuDgAbmhcXHhEGHOvBmUrRMrBM66RnSwmE7/+XzLlCJrbN16Z5mLttMOu3
M7+SHCmMARamjsnVA0yTe9EEl0x/f57err2MmHADPD7FP3ZX6aJbQm0Y2ECFTNkcX4gm5L7tG0T/
VygfhepeYHnOLk1VP6IRy6elaR8b6PytUfABuKmHTrDqNY6KwVVZYMTi8Y2I3UFZXPm0XZZA6fYh
JmWabglW+SIoYQ/6vp6nQwbZmutEXP/ydK1ewqrQiEQnWTvEE5ojXTcSISgQIUA7y4lDTOnwPFRH
Xl/kzpDhiCIGKZj6COqwfEAX4Y1Ee3qpGy9Ush18pxXENfGLmFLS65ufQVo7gl6QmBx//CZ0mzR0
iJowRUksEtFgZby0SM0HglGXBvYzNX3WJan8Tda46Q9ix2gwuAF2KOP+NcYtmHDsM7wbvokmbx/J
qM536PtCZ9d2nwb3E1JF2Hgoe7l1IPF/u1hsc0b83cZq9YX+StByk39xCQ/cOsn48v89RwDf+mfy
6FkXGueSIzNhnuzkeLvMkNkC4KHXbXNTRjds+jeOAIA0Y3ef9zFEqjZExTQWbiXsA4Y9j451jqtZ
zcYS6VlaXK4iJI7EU+dxvDD6dC+UjZEMy1486D0JkKZjCE/cdC8biB8uj0Syresn1T9e9pXIl9NP
f1yOOw8uj/NStHisbJE3wTVbZbiASa3ONPuYpS0V1ADCBWLI1fyLnJszhIqRbr7l1bxZeU58eB8v
T0I2hmSUZtnDE0Hp+d9rwBKXuRMR200aUNDGaYqPQ3lNe4JoL+cqTAuERXnYkdBrWEUtSE1dTc3O
2oGaKpPegkPcSUKbiBN4Xwxmc75J6jm77vRmAcE5E0lKmc/oLVzUgTV1n3Po7oBo6nMIgUlE45jb
3vWrQaRzY5GVERV/CmeVWmf/yt4iCvdoffvYV6kpm4N3XK+GaN67+zhXC4Geh9/dwPgCTozMEKr/
1eO73F1PXD3/5saWtvdVdKGRCKoRobv7n1IzeTgr7HO9VJLseX57CCWm+tkyQs4STfj+Tr2y57Sb
IV1CcAacCfBhQnsl3+wDeaEc+ZKy1Uh6SNOurt8hcExEA6hLC1PHvb3fxefOfWi7C70LKlKmqyry
HqMHj1slljLQDmn5VYUSqixK5Dk5zeRXkocopEne52wnb55qM0P13hKohc8TwMeMmjcX/gfim+iy
dUn/1p109Nn7rtNz0ia2zBx8Y5vqw69wgoBZyJIE9GZWUOfiszjxIlbI2t0gq8xkEMSelzpMeaKI
H6TlGrnWj0lq7zycFWxPdjmQxyf1CV4ulhwARkEAmGVJGfPge1BgvznTcVXEMkzv+atxXEA6e3n8
ghnxRn+w69rvLgsNWeV4QcLh5CFXKYzkv8U2vbN157Sm3gFcg8EqZFp26B6geZyOrJbRhAj7Axvh
0WzD+6Z7uEyxE5jVJEc9D6PJvss+V+plO6goaF44Ka6GAzrTbDOBoPMeCFObQKB45Qy0PsEFwcp7
EJOmhEWU6uovojJrw/cJfgafQQ0Q75lHFXp9EEYY7g74YTnQLImcrWvkA5B4Vn2OYe+itKYRJLNm
aQ3DeBZyrCryqSPTJSJig72ClTrtFHsnrHa6bk7SOoUIjBnYAeYS9J9eKKMC+lzHpfiFVaPLdnGa
bqQaLlXrX6JHyWSXZIq246phQvrc/9hFpAfXYvblgOF4bfkvviGtoOOJn/RCKLLAkYIsf4oKI3DR
tEWd/UrihPcLkUGOCZUJyeWuFSIy1EyVsDvL135F7lTxl17NsRFrHjkXocPE0dF42dSdiW4pbGD6
kVnpvz+pEcqMLFbyCYNVCcChuy/42ukZQWpQ7vmOs2WDQidVsZBv8QFw+RI9dssGi0tkxqjzZyPk
gH8c/Az1Pxgu8TpTr6NeHLooEPPdtD1a8nJ6n/mgIOp1c5hr20wwssCnpZpqAwInZ7yihjpzrWd9
TjzaQ3dFwP3vG+valWCeJSfP9rxrok8mDcswoZUBYktnsuxn9vC9y2cVcmG0JNBvDr5b/CZVuYZE
RS4DU5nEoTOUTqlo/RjXsmZbJpic4zSMyFdvhxZ+KbAYgrNWloOCR8mWLb5FK0Sc/+XBmM1JnMLG
pS2lAE5qt/thn4ZClSHrjulR0UCh0DYu2IswtOE/h2KvIC8H4p2u3u2uUD0TlZGQbTt5qYxyQks/
BzyUQQuomPYg3Yu/J4z3Gbzny7ZCmH4Ubh94lSCJC2yhPN9gx6TUCV/m0wVtzCakeRN267qDSVZ0
NwlyrMrSC7KKUxioXcR5y7MMnL6ZX0fIIRJMuL4k3ys3eSa585RYO96Jf0WcqrHdbCxArB2vr+I1
9LcSuW+rDrwHX2qi6niSyoT46DU6YywJ15lkCCCmULOcRji68HIZVRcHaL7SWhjRqBubF1wIQix6
fDuedY18CJ0AnNLPZT2fMToFfFaVCmEIiRy/QyWor7j5SPFrqJM+g2wBSFDoPHWn1ww89PeyqiPL
Vm+T8P+NEgtLESn3EKNuMLUDfwW7ktGjERlcmu5YxShDrQEIvqlYssVfdpS2ejVRxX/l9ab/e2o1
7Bkt/ySKRP77ZU1ejkFXhQsP10252htb2+UbsuvQWA/sHA7Hpdmd6eUzX1rl3atIfHuiEBx+T3NP
gAUOr6snFO7DFUdQoRPRCwLHqHE9LUKcuqlPbi/E409mlOFz3W5WxMluPpjrcHKiSZUhqpKXrK1p
L7SjEFdikiCiNuG+xIY9gVpDJ22ASpSBKNIuYnfeeS0nIWZd4h1IzsGRPF/3WfUcqeRTdjkxiXb7
J6rdmmDlBA5u74XfzBd5AD0LDSbMmgafRY5KBtIOuDrQuc4r7QGFUy2GMAuhGQpqC71nVkpCWYIh
t26vgSQkq9LTQVMNuWWEwQQl6IB/UUsow4dnfxvxylFXNa1c4Ms5ifSyy92hRWnMuNhC3oDhBknc
imWbU7LDOBwTiOlivwqMGHppAR+cbcbBCu67BE6wvK4Zly7sjWJ33vd1MKOLuPOCBg2P/b6j6rDX
ED7GTE0wmMsm2djmD7S8xqrFq+oNiAUSuU15vnd2t2TLHmZiG3qOYZVsN7CBppd+dWyZ84N1z8zu
iqYMP0ghzQAgEdgSaVTomlRsaKIZD6qnXjyvw0Xh72IVAnu/qsXS0qrs1S3Uh45rjOOiRlR/dNQG
9Hpe4h8SQoS9LrWFupLgAFjNs3ZdDa+Dl7spznVCrwJ12lt/x6q7ELrS8u/pIklpQeq066MFJKrV
cbPx7Hh0uSf9qBDe1VZbaQ/ock9sPo3XxS+C+4YFZbTARDSAEnJ9m8FIueL7SheON1awmgi/CeGk
4Wg9ASCikpXKsD7T4aQ+06Wq196Sc0mzwGRny4i/kHj74tsVGOP8OQ5MUysHmbDmV27nUwOD8Jxb
gO7rvwjx1RSY4d10BoBv0/X1LZ8fUqLeD7+QLdwU75jcVu0TrvMQrVx56C49AdNVGe9ZlWGSxths
a7MihiMBzkOgdhG+y+kHoeW0qnfGAxIXPKSTpvXCITz9FbqZso6Xic8ihgjZVo3UFaV9Ox7f1w+e
zcF12mPOKTMeURoxyrqidEgeP58jCOZ0Ktl6SQeJoPk14lNIYqUHArSzJiti9Cymz4qK5dph7aHK
iRKFCSCPeNBDieFw4IqwGBcQrsWrmh4a3yVL+NNsL5E0tjM3HlenzKNQ6v72ynFTDURfY7h1v+H1
ade+vP/7v7C21jO0MSdZK8rwfWjgRiJ89uYpuBbHa+NygPc/IQab3y4o3iEzpO9rWmC4/gqJe7jO
0z4FGmHNXAdfpKcS2YnBfsKuyzrUxkV1NB5T2f2O+ClTsBPwI5LzhQJiZVeXIzVU0O8OdccTCwN8
V43TgH0jI9tKWbvx+33VkeQd4pyahvoLvvrKRC0pNlpbi3kibqA3PtfkpQAqREMi97Y+TYZw4y06
Q96zNBUBM4Jr30RfKsflK8uLOPENAOYapRtB81P3eK2640PS0/8b9eSQxgH0CqVC67iaZXuSGV/B
vCREzhwC7dZaE73B2frEtteU4FfPqpsj1t7Bfk4USLU0FfXXtJPjp9VhYpbanmfNNvi2fKdsgSvI
D/nOBxWz6Z8Kho+nMiPAdZGVLlh8jsE7NiA1A/quJJ/g2nljhQDyYhD/HYlXEU0MUph0GlosqFe+
YZi5SWQ+MKupo4ulkr0pPKPcpuXBAVPKzo8KYwK/GxpgYW5YDyUPbg2dOSXmgpK1eVsNju2Cz+4p
qkoUts1xJuYaFPxKuH4KSAW34ZTlQaxvmLb/Yfd8KEfo6BsHEHnjv9aWPjKB6aOPUN1Td6GJC8mS
kcBLXTN14B4cVpB8c3D6wVdoCduS8+c1cI46Xgi857N27s1VNHQkOK9ekALlZ+7yFcRapNJ9fm3z
Ra9n2bBBCznn8e7E7n5kWy/lSUhiCZ3jBRIB961w7BMC2viDk4ErKhQ5mXRoNT+F4WYTo9yP/YLx
hE3KS9MgPXbIYgnMapqlpw/O9er49qGLSwkSmkFhIiU/5DYoxCNqcN09hCfS2Ftfhesyu5Csdqyk
lHIobiNKK3JTqJMO7dhbwmiCQVKtnFEgEdJs+E8QJ55q+zqHIs22SoSuqm6fEq4pM1fuslffdnX5
1szJfFoKgHBjzjKldFsJinLVMGteqOa3JDyeid3XvLLHAY1ght+/ORJFOXgWGU0x1Knn1l0pdn8+
04e79jyBNYBrCAZlAeMiXMl+s9+XGbUMIdMQetzYwum3bMUvIdaYRa6vCQuypWGPRwek1Sp7sVIV
STB3Tp5cJgeOT2VDGoEaDwUEDn0OdP32xkiI5wuPUswXaVYvGDvFrzHG3DVnTmu4CPyuKaB28usm
84+C4Q6nniPH0q+eSr59pi5xds3kvS8bPSnKhqv5NNmTZ/fhZVwQTREj/1f6/7ozoVsWF7QBlaAA
DbjZx8DVyIQov2AcQXbRdrupSDbF8U22mEwM/POsv0n7jvZx4AxEkbe+wfNByS6aWtEVdGHymRBr
wdmC1zxfUG503vgnfIZdoiR0HoBW/M67terLqOfKcjnoX5aibw9n9ie5xcUn0gW2J42Qs9GQNwT/
9IG3ggLm4vkg0b/h5451ZcsOdCRQc4A4Q70No8Ju9RxHFIiVkvLAoEs+k48Y5BNshc2YBkd3OUPs
WWdUKKcy7V3SOeStBAu9oObzOcXcvUplwXCEgf3tfw5XEbvfFyxCV4eI/uU1IT4kSH+5RP8SOIZ5
vhj/i48xb07elye52t0qMCWRM8zrtp4XJ4V36I3AxoACNX3ffShTwrBNi4KNrq2uimCD9Dg+tkTR
uU+xWDsdfyJHlVsifwRLwQxVBBJrZIqBHeNirAZoMIpWzscjQqsc69DEzkslw9MMmPZGkYhhq34b
R/yp3noW9KiDzndeOjWfBQpOTYrD8ensl10/x9kNx1aOt20n34Q0Nwtda4+ohnuefcGdcJyJ5lva
tJmb72hxtRPFXeO2fuVjHn3JX7cBrkr/NRgIwKTYsygG6V7SuHsJVfVblSN6Hptd2njlKnCLvz32
+lL3k/UXWb0OXTJaOS+Hlr2JCPY40hSv0R+CL/6fYK4mY+X9nKznYKazglnAUNRkIg0IHOooN/y2
3S+F8GxHk9C1i2xbZ3wd750TfNVkiwb1sMeB7bCbRf5rce6cdn4Au3+srpLFQRGw+5on0hDR/FHM
Sw7i0BPY/8KnyrqOhwhiQcPXbSRl6pv3YrhOck2IymP9fHXU93uPT46a1gattFEQgs/9+n5cnY9s
MqzcZCweJrohSiUvT2C9A0N4oVjI5YWdb1QVNbbAipRmqUwWcfKfPAvbpqr23bWiX29yrvRXbbhV
0EcXcMHw5aJONKlyiD/oP40bpAO45nmChS8FxkslVlmyADCuH7K9aUE0hl4NQVbAasC2Q0Y+BGHI
n0UjL0Ugb3jejsY/EmTjeiYqvAPR54fgZy8Awh1G+/VyKyPydzLt3vgTI9w3lRHFWugTJusN+vxd
iEFHxNDPz+WnHYWl/NsFmO0ZL8+XIBzJpopX7ZvrKcx6At++7WZSdHErPDIkXB08NJnRoaaKvJQ3
Nno2Lv4RhtC+cIq3BLcIy3px4GyhBb/xe5ASRJaOnMdJgea+XjOa38zs76mkplOmfskTOu8IdJ8o
YGKe5D+TxatSxYXmBH6SI4QEQ3k8s70ijI5vE2ETLOtx0cjw+Vw3PX2wmgog2qayJo4PfEULINFl
eGSacpiPHugIpvl5n9pHEsAquaWZZ5lJtnlbvYt2bmGHE6Lkbjugc2rMBTx8V/Mzzr0eIL1dernI
xIbB2E2I+qfCL6Kiae6NriBKlS99DF9uDKQWNMCr3GqFOu3j9M73QSE52nmlKOXLnGfZ08W5CZy0
1iZvRGUq68ASA7pyZbVHHcS6NDPpkqme9+Mf2dsUQsY6e3bG5mqk/RHUECgNzkXDVvJLIh94n9K4
6K3oLAL56/5xz6O7A+A038mpYHZaQZranLkJbL7IRV0A6vecnksWRD7OmEEJ1oh+7qkLxvzFrPp4
fwrEStRIJRSRAC5asmsJku8nbBVkHBNEnnuYrLGD/lctFeJuAIcpMf7p87AWrvfmLFQvBTIr2+as
pdvrIy4qiL9khMRQEOiwCiytcn2dehIl+jNPpdnkh6oJSq8qzH2BQDN247aDC/LqlBVEZChSG/lZ
CSs1goYOaj/4DuWfZfjMtQEJwQ31XJrSi/I9g0l54mJCq0FcDc3gN6iQ+Z2+3Je0IjaSEERzc+5k
uLB8Phsdmfwc5n9MCeIevUrbS6TuBvrrUa6PWknznIjP00XOIY16rIu4MQTZXOxTF79uVqdGw9ME
tzxH1QtYKJVGgAIqz3y9V+VUQXqK/QbCQ9DrUuljD8MZln8krHmq3bX4JYC6JvHQ5eIkRAETN7nL
g8wRJA50KH1WIVaDKmqHJU2e0pZwbarv6GOnHIHAchuCyl1g0CHqbEcwsZYQqKaXxxyVKNFUKfOZ
5T3ZYzYqGGJJjqrYCdS5sxGkED0SWxWw6Dt3RDwR7HwVr5CHlXrHpa79StzXKxxiDRFlRaxiWGR9
L4gpClnPsTwGRAxnJ19i/sA7SF9rQnYK1ZiV2I+dJv13fLoMD+V/ekEFt1LBuOQVk8V0mEpb3vbP
b8t04k4V9o7OIdI1Df9+FarSf86O3wh3cKGoMwkUBQWnMAhaZkx7nuOZTAtPfc6ydH3OeVctTiOV
bPoQEy1y4jxWGISNUvJ+ZWIOsCC+pc5SJK/N1pwMFIym+bUwsYJr6hsw3rqqxJaNIT0SSRuzYah/
4vjMth8vqSKwVtct5knG6i/T+jx/B/MLLzSq+eYDwJk87KhTmWY2jwnt70/TZQkW5AUvqxFbkMRb
43CW99D9+MF46fV0DGx3tnCqZEpb5A6TLZKDrw7svrmXRnefezmcUmGZvA7845CIDIAmZuhUHBcM
Ll+JmP5xtdsYAnHb+PE+iTZbqo1PGDfNIDg4Jj3dews1Vb+BznwIuaO0InKHWmwaEiXuW6qJpMDB
vui+j5n8lYexV4UpytbfQIG+Bm+p3wLDvuz0j4rgT12Sf8K2UOYrWupfSqI8LmL+WpJl1yX8ZtGa
zEhck2X1wBoleLBspqyJwkQKUpPRaDfp2OSY9nQZUiQi0CgQuPtKUuXcKs/0KHengTdnH7tZ3Rgn
JoTULDt6h9b7qPQn40IdmSVZSE8p1Qlbx5pLqF2MDe/1yOsIRlngd+XTxap7/mx+ejcWymrOyEAu
wtlfF4rG0dBM9R3PNunDshRVu+D3XVTtWrBnHtH1PDTlTT851f2ND4z7ls23GrRalA1MmoePb/pk
r7qxW48M3xyKEptG2gxyQz3KITTkyjdZjVkmURokHWh1rzCl6JgPz5yTYJIK2HLhg4X8YPNhiuQd
bIf8VqjTHgd+bYA/O/aDRPxz9PbJWhfxs3Zr5L4o16TNFl22k1VK2QcLDgEMHp5YHnfP8kPJvhVQ
EHnRcVIRzxrFjb/m0oxjzjtocrCR93vBDCAtgaZd2je+i97hNIrFlmTDQYmeBj5LxABBPF6Cv0OQ
V6jkYtRWdQnFnuKW//SFGcjSryW8KOce+ZAHg/DPciY29fWII5YO9HTqMEoQtnneA4uQ+fE8DG9k
IS0boc0m3cycovckZbBhOV79Xw/Ao8hNM+pjqCDJpqV1FzAxiRBIbKEf7fp753rMJqVl+CLZnvQh
KHHPstuXm5ZPm32vNxhYwyJK7jUnN70woZ3DCjo1ZrM52APGrm6EiVs1etcfcEH8OZlbnhKlJYlN
EYTYnD37w4niha7mD93iNMnNCqIWuiKkVC0n53guOVtFRRAbwnm0Kx13q/puZKaspL4gYvBi+j77
U37KMqIHI6xLZRlUKYF4BeqZNJZjAjxTBWRF3hf2RTCEp+1y1NLGlUODKdiNb/egMMGC4utBynnY
Tk26GQUejf1aGTpe9oXbYlbB3A7Rl8jUGgEUWHoB+3gtFMJXuJ/GhNWKValEQM9nIvN84SqWgIV4
0YBuv/BFlKYA1hoEg8+5b9ANBaSo3BxaoqnCSZx4usPfkK0Zp2wocstv5lYe+2/Hh1f5pSjiSswz
ClPeGS8QCFKARXQtwhfJxSSMnJnVcIGZVBL8uxruRZPYBOkW7VHba0uR6+zbZg6ty8ZlLNg/az6J
lRJ1YNpiqUS7CnIblZUTPoRUHLtV8blwb9u4kOyNw0/URgpMiLP3lxbD58+lPlYSXWLvcacYtx3F
ZWbtzx5OsscOcxFlqYiDID/xq09EFCtjSp6O7OBYRY9k+F8EK7XNOoJ03U2lx/PQnbgO/KDMC4p6
7DKkUz0jFOukgFTxZGfJKISGYb+2vG8V4y5B24XoPuf6NKApv8Rc1ZyBNDX3FbXQOgSUdu+tk/4N
GDAOiriuTrKbHvUjJXarOR0h/RFSArBwREuzlOcZaunJko0KQBBirfibpDYGsq6j13EBCEuuMe3L
qrsMAUPSSWIDMuHDl0NoZHRxC0/phz1uqEMFlugn3ajb1ndpBpOgD0i4qJ4emcBQtPsKd8mrBiPb
/BF9jFziEPL3zq9JKT6ad3cXXmV/VFAqFT7o00U+Md1q6EiyedDyTXfpxOK4dtfgmEpou/n7rTpo
DmNPjz17NPf3Va6xntN/HYDQEwxOkx3U35yqTSGwmlGbqtj+OSujFmXxDrPKqP9Vc+/3EQeJOWZH
gFK0ookkHAY6MpkjjOaf/LtgyH7x9qpH0nFiUXlsmUyhychzmpkzfr45OxKFyL94UChKESv1KlFS
AoujrRXp8etBOYyVi5hm/UuIdzhu2phS2MRdwzDdvU0JUIh11cj8SwFL44Zk9gfOpPtbxKbi9HVC
jcHO1XSzRAwonKv3cIoCtHs60AkwITrHTRfQVrKEQUzo9lz6Y+T6plNOv6RilPO3/hgANeT930U0
qaOHpWmx16nToIQpqRyAR0t8EKSjHULXAM3yfMGIisXc79tWg7XZqCywvlnKq0OBUpxrM+vZm9bT
ugHYBKTMNfyfcSSI5GbRrU4YlFdVbz+3sENColejujDAGkTh48EoHWm+g6bBzUhncF+q4EzGsGj5
eN+wS0GU9gXWp6JxNFfLBHw7zmJAfExiYdrEtmuaRhkkW3EFdsyQ+NXPPWm3n9Pvv0WuWUGL7eiu
DZfQLSepk0tKQmgcaDrSIaUkeVa1wpZKtZ96lhiwiAFJpaQa4wkpEbPE3pUWCde8I854NgknnGZ2
NwYynfveNj2gMnFpcJxuwAXzfgBW6PpIFzTmkLkob/QKBg6xugJK9zjHa70TZynewuR4MI6WCi7z
gGJHYu1qVBf7AdWeZT7G2IwMQYVAERSjwic+SkhBsvoISJ4h3Xcq7qOiMXH4UN2qamlttF+300XD
1FkSOilZ1+qvdbJM5ExBqKyi/DUCpCMLH2WeKqnCbhp3yAXI1vEBTuU0F3WPY9ketN2yspTbCI2/
3eAoc2D6E22ymTMPa6htm1nsL/koIGvnQXrCgO3jDDIGiHEI+cQh0FC2gyfPc0VSnvgByqAV6mK8
QmIXCb6toEf5HaEye8NBOmLpQu1YBkh3yn55ilOOJgBScVzvUyn7xcKM8xX13K5zy/SkGwSDTQ3Y
LMYi9ONC1bJPN0BUd6D1XaIvk0/sJEDeaDAGNt15d/aI6MEpiietvulAhLn5R9FhTKz3rqQQpQa4
OdyKUYAPS0tKJyWvxDbDgiXe78YM4doDJD2MtOv6k48gtXHYc6M0iFr7gL69pt8tFqk4cX2cb2Qz
f03Vl27VxixFMBc0ehI8q2GKuzjw+DKzupUf2LuzL+EtoLYsVn1RKHIJL2NTHf1qAk5Y2YVv+6gN
IT19nnl1ERYfxuTAwl12Ghd7BxgWjpXhkAVELQhIeuaRMM2aAl3Q36k/kqF8LlE9b2902+se7nW9
/61n5W+P97wWx2+lAdk2vs1cJuX4hbEMn5xcs0LXpNpJl2DqfIi56tG8JWfl8QRdnBlxpSgqZSXM
VwEIFDzDbc9E5yxt0hnOiwERbXAfSZYvaw3Z7PpUO/9RcD+mBai48fG12jYNzA+IoZI9qHGETkMU
L/9UBrlNt+gkGKHge+T7tn6sIGh6+Rf1rzyZdU6FC697km3w21/oV/eXmN8B+R2wpl4KDhY7bvWR
vjYVRNx0jrgLT9jdtd4kr+3bOclw3R0gJQqhEkKkJdnZrK5cH2Ghir7QzaY82DtFVpZjfgfX/oms
zmovLnF40ijAMKKr4LZgAwO8BWFsHZuZptSSzd7i/NL1lvRjx3cQeeP1E0XgSPLR3+4wAJjl4/Ux
zmb39nd1Cf4RpH0KlZBZilKuriqwGvXFpOXMHZvDQaIPZyDG9aTP8KCQ3wmsZa5zBEC0Dgn1pwdn
Ua9sTdp7Oh7yjH1T+Hgkn0HEQJxV7rWk+dJ6IjKnpHGiBp9ADUMn/qxAqxd0DPbqmgN9X/PbHS2+
rZwPE/RFRTT6JxC7LW6ys/maS06qxiMfEc2rjPllt13NoH3CmeYvm4w4Ak9QeKGDKWl+xcBJeqPY
TeNgxq5OPDco/iMbUOTf6PDft3Sv1NBYaIHL0T+gIOtZWw1Hl9fyYj9MGoVb71T6VWYbl/3GmH6Y
DlXA4E1XFPiX0OsuzD9/81Qe8sYZjyxJklsey7PgnA2P6BXQuqdvTaK7tU3EUgP0nSlhs272kvtY
zQ/g1yn3vijP8kImtthIhw724sGWFhzQaChmOxoM5sSc3rChEDJ3ueK40QTIy844ShdYde44x3uJ
O1JN+nw/+XJ12qsNXZl89RAfGtGyL1CZk2VQujcfUmsGH/ITMJ25KBcBTpkaErClk/ZUq449D4N7
wpdSQzz9pzXi/8zY+OSDtn8MaShrD4im3486vtYtUXvf7wSCaRcF8upipTcw7L4oVIal9NuTCmgQ
GbPDurUcmaJbj3ZBYvB8W/VGZZvJoNZF8fW5tBPCpjbb9tLHTgiCt5tsd/fZzmTWI8gGYncU28uV
cCGeHdI75shp4tKm3/SIXf4YpZ6EFF+xPhbaRu+/xl8t+XL6oOaeNpZcdE6mo0vH9rn8DkRClg6g
NDgfhx61rYQ35CGuweMqX2jtsrMx4glx4jfYyah/4UTufXblIngVtxPbmm0J8BRL8Zs+jYqQrysK
dVd7n423dMgb6vuEsUGbwz9Ty+dnSB/+5EGuIpSCGKtrueO7Ko8/dl+DgZLWC2TIDOEC44vb5csK
ztyJpW81UAdvJjNu7kbeqDPg4UVSiRcPUz5+SERMoAaYqPUtSaW3fR7JHDOOf7r4zvrpXChdYbyF
XvqnRJ9VT3SvO7kA2TPB7lKLZkCiyQ04CPQMeZK0+3VawezJzCXF2UzkzHT+CC3EoxNgRNWozPSk
ow2RizFq2zIfhubqHDH9lrUYd5aOAX6iuBIkyEO2YKcV+fnw+F5Z3mO8dO0mmZghtm8kNA2NFN3Z
VoVmmW3HOHWlrTtTEyhK/rQo4PanTG2c0SBQPKRh4/tL/cev2tEtMrjlNNZvXW/Zuw+fm/PV8MWE
O5+geqfuLqSageoOth7e9iCYshK8+ZTyWPdlZ6fG2wivZAJ/6BZ/ZyaLJNq1B3J4rnUBI3iFZXiM
oenCBve/9iQ402/l4MWNyficEhI0d9iXGUHRz23qeqp0bwcgJYeQmjkX8RRGvTcSq4FMrNGyAtVJ
M+J18sPon4TVyIlPIqJIK0px0Lwf6qQ+qIaD3rOWuUrhyfA4y0MhB/ofFtDqBmQehLElVmF9LcZP
ZJC41RVUsrV7fawkJN4lzf5vFZsHSMfiuDN7vTGN52p5Sa0l5W6NV4ARD48ZEgATW/oQBHeljmUV
F58SMkgc9/RZIALEBgOIIBGks+BxDJkuIPmTzcTOns2SAmWh2VZTv0k1nkcdFP242ZuLRYxdI3gf
UP8KXBE3FN3sqhsDeMtNCERGFZgTQnvzJct5zF6gWMbFRJrbxS1pycy5bkfg1Iw/iG1hFvFWlQ/p
+CaHMjJ8H1g7sI1xfvArq3fQrTEo/9zQvYOYYWCU5lLxECwAvTyGgfPsB3AWbTVpCwAiZRGfMoNi
NDhYpRMAO/owwFvGRX+IFvMwTGy5mJftOICkcEHTJHIT+oQMfinE1zDh3/YhroRxCtsP1czeK1Ez
Mc+JhXYUZLHWAKFMSVTE3e8wmVH5uv5nIwK8Aw6GtoLpOaOxXdDHTqjTatHZGcmNsRrT9sJi9D9M
8NHpbHFWlp0WKTzSfFYleHjc+W/aOgwZQ7pn+1xbKho0E9xHYOpinv3WdFj1QDvPnUGvJIhjevZQ
pgJz6fbqX/0Hxq45q5ZJkXk3FjnfY3PdJxR7S5kG7MjZV1BbV8v2lmmnnQRG93GKyi3m90FQeYXF
ocp9ig3BKRIMqMc6tfUatCbLTbKgwayq3w2eqIYS4627s6UejEIgdnEB3xZdHq5pFZzwvYzllDJV
yr6NOlD3HmVE1odLY+CPZXCLM0+UYvDikHR1I871StXtaL92GTcPsAqdJq/XM9d6j1PFvkyQAZ0j
fyVkc7nnS3nPXFgkn1UhJJuqV38qjYdNIPdDaLB9iXN/QkhUR9qjcOZE2TmphfIyuLHK25dSEHz+
5n3gTDQXhjIlLMWRxwyJdJRXPFcTf952xPJCPYu06zYQGwbjLGPgfmpeikOiKHjutexnXJEkyDwY
wZ0R07sTesC4t15OPrRBv487xdbcD3ryLplpzzsOShJV5xggCFeP7+73ZY6v+PIME2GXeXcmPb4m
dp9VEqLXp6OCQiSZn3oD7/xCU4g3TD14xyAKDSsCdHEpW4KR3f9P2uyPF+sSlIfcN7b9nFnZRnhq
TS5+bvrMJgqpKj90szjA+UQz74Ypxr2p1soeB+E0+Zj446FPrEhhp418dTi6Dc1O8w9CesXGb3s5
q6xUKLza87oS+AhVo+AQy7iHPKHb0dbpxWf8LNkTxfqikTyg2uXCT9U4uANZ1KQe8efpvu6RTY3e
l6cWQfTCVXrog6ko7g6V0XNsM378xNgHDxoIRy+2cZEoQsxAWmN4i6DuOVcbgM/qZ3HM5Y/z360Z
Qn4VI/S1Um/yrMkiesIgtpFtbKAvxrjLMx9EI+j9376NMYb6Om34ZA78A0BBJZJGoT2O68yXGkXo
fXGPmGku0n1CNocjjDJWB6dwmJwnER+g9LMYpxeXCcEEvgFYE7kYwVI93P349GJskRcQUBpKk2AS
pPRe9nLeoWTwo6dgLhOl/Qk1DgHZYwzecrReuLMZ7ZuHZ0OOIjNub+kGiCJbM++6hb3NmZyjVhU/
eeR8j9IZqfYhs8T3VXYwRztDBQjNZF1d0i0kDBQO8i581n01x6VsV4AV+lo7QNherzbazzB398Mk
1aZvVk55w7ryzetNMEpmRDHnJV10tcuuk8GwJIBP2nK4vHXzMq9t+JQVZaXfR3H3ckoQaCmIwljY
2QPuRFCbwi5XFElcD4UalcJEQ/E4oCD3IUn2KA+8wN67ECe1KHg3YV4vI3+9GwB9UdSo/Ah8e7i6
lK37L62IyBPFQL37edQKB2659QZGW4jcYmOquvEGoySd+pBrglPJivNLQsbFqqt2QoL7IZXU8xHx
1YyB1FZYjQ6IrFPRNT4fdUOyHLWbf/WppSoZRGuTNo2EnXuh6M/ro8wif0LdZfkus+5IuSKSADab
bwi14MQGrVsiXn5cZp5zUUi8e7o8DVRd72K39fqNurFkDc13b3QwjcMTEaQAKmUqPo+K+CJGjHlv
1n1ThxAYklnZYnyjhn+47NHlL2AFhTxWeW8pjh6b4yKfvbA7UrM5sTMaRdAyV9fAdalXINQ3+8TT
vLr4s/+YF6HNmRsAO75/aZaO1LjDuPJ7AUoyGrM+6KRPpVxo24LNVGV/Ew2JMOz1LPRWaC1gP+VR
91//gLIkyPQr/CS45UoBRXJjmz8TxwRlyXsQEQemFWOR/GJ1I5kP0raxUuVKioy1vtlVnyM2vO2/
DwQvotG/H/Ec41ZMSLig3dJ84FK9pTErtfCWDQyvo281VVmE8aK/TQmPF0xt79yS0gClyTNmmTcn
S4FPoMSroLtrJV+dQ0/4EzpKMvCS2hIV0atcfa7p4G0TZQXARtnuP5p/drXnJz4ZaWfm2ezziEQ1
UuzrlZE+c7VtsVYRB+77irpuZG+dPm+c0LN24iUO7OsZcBK/Y7fZ8FyKYrQpUIp5UzHSDDB+4hMm
ZFBCh/bEKbqMXx7GFnyBBDfbYe3SaxTkHjJZomNq7uMUJdswKxF4PhuC3Wsl2WiT3TyU7O0Cz7xJ
5O54BZM3k35uRjYpusaD1PgdbOSwVWReId8660mjuPsWzOx6PvQwY9oSkbYRgpEqNq0tjxCK+PED
gxgarKcynF/vE8Qv14xQqVm23p2sXtnCoGw9U1C/ZRfOoD9cC3EZXYFSNVyWJpWXqsZ5HJxT6CjD
1jAPbLJnzxw3N83Mx33PCZmjOhEPOH2oPb9p7KW/TV0b0IvbYfijJVCpeUeypkctcqPYOAouIpgQ
gNcXZ27Ediu9Bkg0MjHyNCBioyKVj9CU/Eu1nk/Jz7xul/I9LNmutyYqDYfIoDIlY8Wh20l09+92
efU7QprWp0fQRDRF6Gs/qvO4CvwdXlOPtdL9XGvGVsbTZ9DaDdsus2Bsz3nrQcMgcSCZu3rEl6sl
9oJ0n+bbQ62rsq5SRYyb4hBvtR+nYqy8Rvq7E1pSr9UXyAhb6GIbe+yiWfJ0BZGAY6B/Orka8Zo3
cXHQMa1t0VE3eBuaYkQCaGtHSrxFDANTROsZFEm2tSUWz6C4HbEinwbLY/XWMG6C3qzeWA3R45pF
jFWPJdU6xhBG7DrRXlUPsbAMKf7OQOy7OH3wqEgMDoXdR3YGJFnHsSnQ0d1XQTqWAgGqc/xTtO6h
jXKfbWKNJKPVvjThbw2GJ59d/Evw1FU3NjOYblcp0cHMSmQiZuci1QgiEC9bB7GHdZWrk0hS8KbH
k3H3h9DCKokU7K/mBry+nDmQz+2JlhTlcJPX1j/p101UDQf4o0Z6giAe8wT6Qpkk+SHa3B2QOpUn
vRCjXzNehZ9Oz6/e4avp7lB3rZ1qPlfabBuIzCHBBhqb+3JnvtEfgHHRXolpzyybeF4gem2kQ2aq
HfYvUCGqSVcOXt4lHSi47n+6FQvkiRAisICnm3AFnq1h7W0GFvQlHi1+ZmpytBtXNXdX3ywA3S+M
76m/jXCj0rBe27TOrYvmVftpBD4J+FqhVwMKAlDI1apaleb5xCCazG/rO8I4L6ZVeELtCUlluDlp
zEsBui0e4FzVAkqgokxUE+gzIgTTPKMBdUSyHaUBGtj5/oOVxkX86en8pQQaKVjmApPBDLHmawS+
OR3fAt4Viyh6HkPIHfLaJanvhgvpSFdqv2G1lqyYHno6hvgoOTpa0g7LUig8AfycRtNNft0L0d5u
2GxvOP4mRHaNpWr6XUA6ZXcfID4odXMu66+LM+z2hkZe/MhkcLIpuUGNU1Hccb2kllcmHsu6ZAYP
0ztwWDDN5XyadOypPG9FGWV/Um1cTi/mt0roCDWetp2jn8KhCTPpOTfMfmvTFrXMd1YL/ReJ3CRx
B0cyfpIFZjY5dFtm9joSEyLXs49sBTUQSTRQ12hwjnFbxIPvgMcQq/+Am9Sqx3FbWI6FUtr2gk+W
lCUnSF47jRlkeOzOnmhrsBsx/O5wNNzd/fANfReK/WbOrz4FcdvnPCRqIIecFUYViYv2Q8tU/Id6
J52PiIIgZ3fz/ot858fk/fpRAkekGbF3rgM7ZE3EnzimorW3p1LGnh/mSjYjuKrXMECPuTHPo8WI
DgnjZSk2+lNMGE273cIqQwgiN5KSQnhrj2f04y37E8GEmrcFlcr+C1dL0eoP0uqHwAjejsM8wxvf
QWL2W4+ZYtAvfQNdeXKK6Geek4Yyhi5uJ7SqPQEKZvO2LWkdC651Cr13C7lkPDrVOW3W/pcruAbX
9rdhA4/T8dp/N6AkM8qlEaEuNX3YcabyS1SxMhZX11ynce6Rt0xo6RaqVRr00nJ6cONnMCtKUF1N
no5r18x668mcE0G4a3Ves00l6yjcaBNI19skDe/sEt8YO2s81Rv4bCiK7IzLv+MaGfOybkR2X3FP
ttqzzdicvkXWzd+OkOqixfUwtrWroN8ywo3o8SpqrxBr8lqw/J956q4PLzz6iKCODdYNj9p3sJq3
1gqqwu7IAeUlRm3H0gQhK3AM5nn+kslbN9GZr3RhVbO23b8uJ6P+l/MxWI7vn3X8bN/fgh5Zhiq0
Oh0WKLGRQobx+NMnBudD9zFxHQnmcsaKfFoLSqSw+dByflHHO4x++r6yPHFLsBaLW3YbeG4NgWRf
QOyURARDJI5TZHmS7Sir5MzymCxkqm8dUljmUg11dcdRManVL0BTJ7czb60X32hehrjOrXmKarVh
+eGlTbkLPOmLckG+2NU7WKMOBk6yA+4pnvaM32+JZrUn74VTXreaxF9n5PiS2MeqRW0BAw8Ja9VD
WlJnMuKX4B/KgLOAW810oW7BSivxQCSyiQtZ/JX2bb01ji0QCyUlm11kkxHwZSJ6idK82uV1Z3Os
Dk/ERt/2U63yl7lwWddmR/AmV4D6+MObUqtVbRZWaUH/JgFNE41WG7xjZDXiG0bcca/9JtG6hQ7t
in8WQIYv8YQGsbCHWRsGCseYiwc7LlnDX72QeM/WHppQXvinNikeM+S+fr6ARRxUkohV+KcMXFML
1+UfifH3sNGGcGMoKaqH0iPrx03doCEfQmZsHrHkCqSxXK7d9M9IcqXwsvS7/tLHzoSBwGcplNYr
hTE60Xm2N1ZzJz53jw+eLU0p6mghmwj/OKGZFeQ9N1JxGBa+r3VR5H7bKfKCIYREUBytRZI8P/s7
uMIvFe4gLBUqnaKBNh5DFCrh+9Vuw4ZmOOAwKXcd26SXoHUqQG8Ui5QbBRdUe906ciZRfVHwJjfr
G45ALOTdvIBoZoVBuhu++2M/cDLRx8l6CHj58JJqIDYrmNv16LaomKZuKPGGb+V+4u5HsjnsrKP2
4bVyB/epwSd71bUf99QhwJsuYwnCYhnhOFkpU3/7FdqPJ0dXk1kpIWxVlGD4vsncsWndyI4ESJsk
kpuzvoc1w/ztVEGx6CwSCU2yBXwiDJAuOjTcWLzj5st4kQf0TTMosiDsUHEQRl9F1v3B75uNXbUC
hipwItfCbY7P6/PbLF9LRlWQChOlPjlAAh424160yJf6goXlPPiUkyFp9l+oeVoWHRb8b4UzU32Y
BDLg4sI4/ONMK1k17h/oNVa+AVt/TLKodOeydvt4oaQrZZIPjSWA2zVjZGekcKyo3ZPEmVMOhw+N
t9ypIShuRT0PuvCWy5tAgxjJ92QdGo7ODTBbK7H1vfN2cgxOj1x6rlUHd5mOBFT2kI7yu7tlprS4
0JClK/0+PW4aMy/RQ+Mmb27lkhLu3yiRELuAoyfegeS6yhoHTfRTTemduAcjiTMtEvHZSUnAS0OQ
jFd8zLeCS5kA35QjHIgdC6gTipjKPxqPbi2CTiD0ZE++pfiwvrl5ndpRfLytzeWsIo2J6rS7lwNz
NXPPpjl2uRy05NDhTJvG6MlW8yXobwdN6+fVCKUTQYCAwqs7bt5wol0XmpyPUlgEqssc+2Z/+fMD
fpXuJ1tGTXit7WGX32OZRCsa6vWRorTjGqQ7Ii5ejc6AH1ixsZJXpXhlzP3BuJNiNN/WqKR9fmje
17hLxgfU7NFb/4zYiWoWnn5PMhDkDUn0BoMEcjrIwKeXGUtyGdceO42cf21g0zux0ws7lqrtAiE+
pOdfy07cJwK7e+mCEPM65NJ7QY4+OejjTZ5CSYejk26hM0QYJj6QaWUEKLVpl24DLv//8Ltz0NGS
0r25GFG4HyMj0UkGRUs2Rjh9AYusTaT/Z5sP7oV4FS3wxmmGbCrwuF5yceb7rEA9WjEmAcL8mu6v
UpEWKj+cC/8ZorkxLXTmfv+sFJXN6swflEP7u7b8VyVwIV8+OHJl6Nj05MnHaPkQpdaVBSWkcCnN
Jtqm/IGgfa068QKyh6zZUA7ZXuLFe4hCgq3uhiVJxhIQ/j3ONO/nhgxs8I1MNLlElTtAeFkaAXg3
bslvtUPtuhx+pQzBW7M0wX+XtOArfpYwD0gImikzPDyXlBZ7kIL2NJTbMc8nBcEaaTaENo0KtSsN
cdfoNqxBNTnffTsy8uMPxLkKvBqLJu+M1jZAHohIJNf+GCHL6LgiufqSvsGugQ59pVX3ZjYHIiOe
yCaVRVX0OJGkIF78PqjdSrAwucxAfWofFLZrm0rGCdwRND+2mK+8Q/rufBfWmjIv7AGwLWprDdQ4
vwO+CyHSoRYU4Pb853upgb5cbrFoJcVSFvRpSpucaCOlH7+EvOkxLNAsBUw1CEdvl+pE0iYHqqv9
4Ar3aSyUt+XjzKC5Rvj7QFg7oq9w3FYRUpNOxbEbRjcXXz8by2CkBTjBzAb8Z0pYsV3z1RHpPoRE
//kSBsYkSl4aPMu5SnHfsfH0chC5xO+6lbrQcw+KX2vosDhnxSPHRd0HDLH4eVCcZYT2H+qHuVjh
skdxU1T6/IcZoJROVvpyf7u3ytnKXTCAlc1niA6l8BAB7EEV/4Xv5WeV9fdMHxUS0/5s9378WbDI
NcW+V3StQvKo4Vf31uH3aJWFWANr86EHCi9MvUzv0HyLtV5UjW/Jqm2ikeY68tTpUdrcEqluhOBu
I+0KrH86X4GgF4hOWFm1aKTgRMNTjD4u3cIfQCug216C+NjnNsngE8LHIOu/jujmUXSsgtYsqVwC
JGfO01RtoaG0zrmgNdf1DTqFbQFVHIKbuDcF+vRP6tD1VBtWUB0kpO/j9OEG82n7vo6itshmYw0z
tTHr7uRXxbVcu862z+nEOgNPezsnKFM2nfPD43blydViiHkOcDzqkT7YuBiSYvGYBZooobqOiZgP
adJCkIAHnXqWAr8XOfHDxzb3F3yFWlJhT3OENYskjbx/2QAnnd/WtwMxmisF86bYXxwDNfeSe6zz
2uZnxTrVVhUuLeNVts5gpjVP9adrtKxqX1GhyXzv1jAYcD9NRHcPSLTFWnmBcP5XGe1MY3D4gZ/9
X1sW+ToHpgMtl0kxSSHxT1/HIixvVOlGj4LhfJY+ORL6dPNdU85Rd5nWPmWc4lYoidFpZ5nwIf4K
7MwjdC+ZE9Kdf7BiZyEHMMBv7uIvqT1YQH1YOFSG9QrGuO0iTjHEgpgIETdYoUht0/qKip1tZ2R9
A1I1K3768JebldfDXNvst2pmdyH2V8ps8PvpDEbVJG/58kH+Kd28cxMyOwB2vGgNQ7YzXm/M22Ys
h7UADcYZiKV2/8iQKAPKRE7zN0gghal6CRZc7cqnypa049cB8thXIiwZAfzeerFb9iFIpVcRYmEG
vSw8oOTIboTYNaLTp2oD2/6DiETr5YCSEsK1oCr3q0DeqDWdrhDFGOz4kcCrHh6FoaxgUxn9TH+3
WMY+EyvczXUeFSHyjyIM/BzmQ6Nwlh4C9c+i4GoMUnXRbqqmlObB5PQybZgKiREitSRwa24u5Sno
JCv5jVBBH9nzID1ZCxdrFaUawZ2S7+s6dcKfSpKBbwI0RlHZqU+Vuek5uAqvjZ4I95odSc2dppQU
T0jnxmQRRXd5qwsFdovi815WWhWzainnA6ZMnxCmFvA757v13o2pZoj2nut7B0z1pQftIuiJSvBh
Mlpj0GTamoaIiFhqVwWdYuTlTE+71kQPAxgid2oPsWxxCfUT8E1OqEeMevRzH2A5Bnjh4CTDEKJ4
ud0OzjTTo4vf/ysqC/Qkvbj0c2RvPtMr7FNJ79DWikTWu5YxOkSwkg+dPtEMQT0cMe7QjZ+R9lVA
IO+H0QlylZpDGkenGKwFmmCB2zyysZroQ4gvSnJXMYYHZ2lNixAiCfSyQKj87wZWlKaatvoI+ucV
uu/UFgDxkz/2Cv+E4RzLoRa1RDpSZv76FbhwYEZQIIpfqHBDg/UAuQBWfMcrqJzMjeZr43Oo0H/3
HucViRPVioe2LBvCBOvds02qaJavty/eobSCahhuflN9SBm8bLcZVf5BKAjsPEzMXbkq5e97++fS
fi1nfsj0EY3zuEiIVnsjQwJD2oLFYcm3+ZPGpq+yK5r3k7ykWT5jWvS5T0ZqBf4ZqWCQg6PpBVvR
84nrC23RJ4EugDD4pxITgYhJOO74HMIy2SHY7oYEVQIzHq58oPpnCLje7yssu8u3te8eBUTTv7e5
Ca9bXfLrrDjJi4n8qziWW+PbBkYMAacA3fhJayHPV/i+GTfO2HVOu0sF9cZG9AAa9oLd4PYIFgVE
NuEN6pvdHWK2tyI8FM52bd61G6yCJoNJqj1TDpYvDnUjaZP8wWjhScjaDiJQ0S/4CLX4T4JwwAsV
DSBubq7hjhqZVWuR03/cQyTROKCASYkt1zsTCH5OxHAo9SC2ucoUti8Zcae8BrjQrlgFehGeVxBd
aD1oynfFE+q5bmouUkwC/9VGYv+WS3cE/ZDmHlI7Xg5ffHBJKaM2IdaeLkztgt1UWEXgdA3xDCHR
Leg+oIt4+bh1TvKNNy75Gyz2iYd20HotwuOjxldxHK6TOVVmBUQWE4gSY/yYxdnsgQLH7DQVlgjF
RN96GFKmea8+6X/bsEI1KDlPOPTn4VMMKQvQE7epVwk1+qFUCaJzIX/BgvAH58c2qD2biHV7c9O/
uw8jDJIrMVnZhd5J/kfb8AxgonaEOTY0OWGPbPYR3YJGQEiz6u0tTJXf9qK3CSnOS7gd/vRygfn7
zmA67kVbvyrnRpaq53yJeQcEBVqP3Kw0QiCk6NxzBgrp3X/52vbt64wxxASaf61PwgX8hXBtJxSr
9U5viuZ9TbFAgNAKMGGo0CEBAIMrJIkOWhTEFlSNrHIwGbsE3drUxq874/jwKVrQ3ELgOTIl1Yb3
iGD7DecYhRfnEJSUcZyWZytBZEY0hVZBC3E30iBKvtaBeMUMD9oGMGG4aO08zqCwW/2sTHnuZTCL
2VvLaWyzrJyDqrPPm5z2wCV421gVjISaaLtLzp8qUzqDFAG7LLEiLu/8D6BtDt6ov2aVayOkqhR9
2BsrLRmYuWXsYJRrIP+Gn6H4GnQSX7j5hN5tBHATnJEFyZ+MGPjBvLOCGIVJke2wSgQJ8Afp0x/P
b9z6l06A3LCbbdWonKk7zAIZeANORwOzSgN7/zUjsnOzCCZVKYGDkvjGIpwiLlkIrs2VRR2oPAu6
5u2GcvWM+mT5FliFQqWmODVkcWhaJZ6cjB8w7IBhkEbdlb2XU1suJ7DDSc4f/oAjVRJ9ytpsXIe/
1tUDWoTS4oB1Qy9CRizaFB8ag+BR0CD+MrWIyzQKmivV2Pgl5eY0sS9BlCRNsJr+7m/IvVQBFFd2
4zxDUJdc43OVMJgRnvxM7Y9Sf47za1pxEDlP42bVJU5YHAvHJW1b2nVYceVtstwlyh6UDOyBrYEe
9Bt2ZEBP+A4vr9akk02oVfvA8r/9vgh0QHiF58ZtVDRR1jpxxdqukIn1YRRM1yDuT1aluBXuiAKr
iiCK2BZlinJhhlpm39dxrMPjHTTQ9iBJ5TYNP+XvpyGobtSrgmOfKDbzaBM00mSz7htH8Svc0hgT
9fJRV17fGNJa8JRq1PIvJrq8b4FdIufhaD6pyD7bsgkeFg/EfU1yjpQlauan5vaLjz/MxaTEWJlq
aYUyIkS2idCMu88X3tfHdyJiKWH/7Z4RLU1SKjO0k7sX1Mtaz8lk1jNZkmp0ltNGz2cC8wt4x3Zt
aq58BuUd/gKsDEEdeq0xPTdbifD8MI9eEmuQ4SfclMSXADlu5pLBPKFJqDS7bp2XXVpbRUScuLF6
YkyVoOAlnCuHbC5+9/BGAYX/7i+y3Nzj7KMGvu/dw6vStt3rQLblg2dQLhN3Ka0Fz2BxT3A9x8s6
wmpDFnIXgqx8y1/hykAneCbUWVBtXdBcfzITyWytAvVBeupFNKjrzkvh/EjghbVd/8OdOY5GsYlI
RnEp44K25YWg6UktAbXhQhdnoROt93PDSBNTLKT+Myod8Ba14mOqIBY7FjfBjcZVzHXj+cEUYeEh
WKZN/jwZitdpZ8nztkYjZZJVKGyX2Kq9QYOlfbq2YPStKPcLKXYmDnEKz+lczNxwqZg0j8uGTis8
U4JNTaDcF8KKK59ydjM0HwKf9GVbIrBZibiFMO+FzEkfWGw/tCAmi9132KMwl+g++5unv8tlDU1O
TrW8x/b4HunJh7jpnmHzvH7HD6W7WDsJzwF1tm7Zi3iFRTXXi5Ipw3nLGWXISyOfPaxNMWLokASE
TSJ2eXZiXAHsRkkRT+lYljs9x6LwkXWgXZwApLhKey9IC1/zJq25u36muTM73N8pyfHyNDfNfLuD
NJMuajue+nxI6ufdlG6wkaOJ8soAFub/+0ROvIdbUG9/va2W90n53n8j2wV354+atD4spNkXiNWL
/ymNLfEurAJhtta/myW9JKnt2ROTNaNbX6rhVwbrlzScQ9m3PqtfLIrT/w4/F+GdDK08sAU8zUp3
IsBHee3/WrSLf/7FpWM98pv40Ze/xrkVEg8mhfnLZENZvuDRoPaqeNSWl1xzhc2IwZ6Df9gGzNU5
dc4D9gM5J7KoqYQMxA9sl78W1k/eNK4Vz69IOuMSAfO03/IV4rqQMbsmS8z2l3IAGuWNtk1RT/8X
CgTl2EcJ79jVjzuEykBdqni8tWZl7atDby7u+iiVoijAJlt6xUtZ3VRRoocGDj4LpvdJ5uPPcZbG
VT8JNZZbdD1smFw5jSylQC6OaDMKUZtnzMZnkHXg9gBmad1ZX0/R4+zJzqGBDrlUWOXVdcwkk6lX
gg3zEFQFqwSuqx+E050chrItdfvP3jZxiIZbE6kGZRhXouzJjIy6Ut7RTJyoqsGzFfkZlymp+Wq+
4fVDK2Pd+oUTRtZwQ1w0WbJEN/ez8Cc93Ivnnt7XJZD1e8vCS2hsalFwuMCmdU1HVoVkn3l24u4Z
iWgVUeq0X7SgX07e9NphAAciGIHzkMstx8oyOUbcDKP3LZkTybdXvhEi6dULbHbaUOGppemla7RH
04Xe87uRjMz8y1pZsyd3/hIYCyvIWQIK0zoGhcYeQZrfrtg893HsInDc5oXtd0NsAAeI1ZbL9avB
SSHxFjDRz1llsj4ZzjPFQLdoYzQwPabmf04yaRYDtRA6DfYbbpEP+dpXG198Kn/jWukj4x38cmPG
JU6ZazUTkaZZA1Uu/kb2fIQSMOeIt+FfJWfPwI4heZNGBzPvmwEeyKK47H6Cfb3UM7Gqxx+7ZXOU
XuITqFVsc/CXhlJxBApDRKaqIv03ltOID68q3rJq/Z5bYw7cj7X8sbYNy6xdq3oHjNgi4DWVTRcD
iVAiSUbSQCjG8cgEizUfOJokgk0eDhhmKwnPr4jjSaypeB/Yph3VhRaW1fkgEN+EvMjkBQZN21en
z3Ri/8QOfyzHiljWduGeZY8feMDI5KPcQMpGgQqTfx7LK0v44nddtBrTpTYS9KHQLjLcFl/oHL9j
Jsic1fyfZ0HKlzjQnspddPvQRelBDokbv2AfqDIF8j3TtDtCkWAO60/BnXqMlOnsQmyC+ck9+Vn0
Kluhq3GhdsG66ZOyxl/2ExiLr5wuABM8+GKmlM0m05+HBHy6agvEAnQiWjvZdHLt9rw3QeQHdLfg
nJ7KMlIMM6VdhwZ+9knIVrSaU/ueX5o2Ceu02W9c7xorsF69UCkiDuRYkRfqp69MPxpmmOqwZqOZ
WnIRNr2zeWsxVZuhf2i1HbMYZNa9LbIGeHb9Zx0dRVcY3LaAyefTf3OiQT+q7RLgMGQju2nA/Pr3
dxdj7mWALig/agzJjWwfYdYW8+k8Sowp8hBkNoeI1cMEuAnzxP+23LiDD/hYh4VTapRJyNLZ/aFS
Wa9zZxfNzIw7UMWNO7GPkjPpgGgD0HpiOWV3GhiKs8zJnsM7FGIiosDGg7Mxo/o3XqAH1fofNiVt
Pb01MOWiCGsvr/qkp7JwGJzw6hjSkh5OpGMFpvHWbwuKmHdDCoPw0kPu73kIMe4gke0biC0wVJyh
HN/Ya2Tivm07LI1bjIzvR194zek0mXj2aoi/dW/xDxb9feBXD/hqZilBftWXjSirVGIHet7U83fn
3gqUtIG2h/Zrd6yZyJZ8zWaF1CsRYT5oDX9KGvBD/fERbfVVDY6XpQ8eUyecAEAgUzrwnAZrpkap
65z4mF5wt/FO8wdTVNVngJBnpmvW+Qcp2HSZwZu8LYfpTqKY5xBuYHfSE0yd2U8heL8P8asn0L3N
fhnLwgy84PIhihuwAgIrEl5zVRKPFgxIlHg9gD5PBQkQWWfZ//Rx5GBhMQ28rCD1u0Lx/USBDupF
Zyj+CSFwDp0C8V1afYb2uohFSs2OZLNHLelA4CLRIXD6keK1Q7pO/pBxtzZSnrxyKSs6uJSpMjAz
cxiy+875uv3Cyv05REqE4RSzMYESyyjX8nprMuxyrasVdqzl2uPV0RGL0jGcujsYrQyY5A6hIlXs
0+QVd2hYBaElcRpTPKZlKCNWrkPSQO5EW4ems7dXrh9/9hAk73s7dOvfGPc4jODRabM/1IQ6VouJ
SUaBde1DTUAvPv0MVY6dN3yfwFxRrVwisiGMzaGrvEKHfHjThn6jwJajD0nYKYFoJNVJaPeT1sFD
xAS9c/xY5ZQgUKML4DEknK8cpsc5HxIMyAZPTZWnFNgTw9UKPrkAN72yXf5zd4dctZMAMzxnP0zL
rSxxuKyNq3tenXdGRLlb/4YychoOOLZcYEJzslQibkp/9gkuc30rWCUNnOrx2lLaaBxDuka+K7HB
5qPKIrVJfY1qiGuRkKgdNSeQf4cOv6rXfQFLP3Fi6p2hXyfFVvQjwpD5x0pHLcFNtJXysKE7LVmR
NfR6/NG0oNp16S1scIXmjNYdd7DtGbAGP1H7U9WFhtMECLvIoU5ZdqnWaWrupvLkIEZgF5PVHi7u
/r1hhV3ww86D3cO9CErmIklxdiPVwiNQK5DPyX4iepq0CEXS1X5TirtI4mwCJU9OCPriLYMksk0K
K8og1zgtxgnVu/F4R76doTNH45kQzxZYIvDodxRXxn/bNNlXTrysVB2JM+6zYarxAZ6fe1ucmHox
cGjilTTWq9fIjRydEjnQKlOWZATVxmWK2a6k8/kT6qJn6PdOleC2shMCddzj4UCjjL6xAfDW3EEr
EpJaDxOnGbcscfKKfmEp8sBLyEWObJY3lmze/rovTVA8D7G9txxprqFnOomVj4sIGTBF/6+XXp3C
0XKvyKBgBnBV97tB4NpW2k4jCVIAEqZoZ8ul+MnQ6H63nn/T+9k28SCk2JSW8cG4EViqLDvuT4Gk
rMWUjfKlApRknnG1gkTs24FYUfrHdzIZm1DAvgjM1E63NmUHDHwmtbLRskTdG2bhWlN7GdOZFPbo
xC7wo8f5I94ttpdbrNHFvpIDbSvN7vhMCdPByU9pj407f7Xs658x9CknOv8tSRn2kSA5VyX1mzb0
QNqx/iNbg7mHCfeAYeCfQsfTMgyXgWswLovU2vmHISg/Rdu8Bef9snU7NxPf0etcagK0i24OrtVi
+EaROEi6Z9p/D1FMaRpilqvIAnzq1jdqLWxBLfdEWcb/VrY1ofrRcpMEovhWG2W/Zu55jPalZgQX
dnhqqy0GHD7aQuIpS5CMsPkU5O3+eJsHAWnRb51Vea0fEVKl8uSsDovfRtcNZXPjql2tlNjiTXa+
xGGWa2OotEBWc1EzA+5RwPbLw9GBut03Yb1CYR1i1dAJypFYLUcTDCkOadeCUaw3J9xZTy9Ne4Ao
7sWS+CQz1DFJmkG3Qx0FgNhLLZFXYX95ZgUeUOhCDLrW91mBcrL2/tDqWSDC9q/nGjKFJu+Pa33J
QOzNmtDmlT7OsGdru9NIQgPwTkximF9z6ByDPCr8qAf8EF+HeTMay55F0bNmMy5t3Kq3svDIodsF
yFo+x8VYVruQqljJs845+m+M2x082lnoqmXfAcDcWQMAgUpSv8Dfurs+ogyuBEFXYO5klnsJ6e9O
Bub+sIs1qYcGiVYjsl1IggIQ+Aipo5+T5TyzB3+kP4W7YSk7qyQ/Ma8PFxTcGtzRL813ESJIXp/k
TseEk/m7AeSqdfWjumzA4B16vkrKq6u8I+C5qajusb86Aye4C8s2tYSYjQ0G9+nNJjHUA/ngxhxA
md2b9heuhmdDDOV0my7VJLcB2PUddB15McWbFp06kTifT9+8JRSHyiLzpz080TIt62Z6i+0JyAHi
amLOUtILK82w7tzSHE1TdWz9f0rYjkY9tk6eHgnoQtXi7a1jvdnYRgEsEj9qvqse2s/gWUFQsa9O
fglVm/uY1SxEIi5yV3KG6BFz/PKNTSJ44ZocS517NGZiwsl+JQPgxKJupYjNHVJeZZ4Q4x0q740j
fRWe0o8SyW7fbB+ccaOtj/sKNWj8GeJLeHPlbhYqoKp/Q7R8xBnDtVWvlvT58LEZmK9vpVgumtuV
1P0LQr/XT/xadGxHnJe7bPK0pokbGByN0SEBYZeQVdXXOt/4YSJTwg1zK4g/Cl7buSXFEYrIOJJr
MIiWYQJPIKk80JQM756Pr5Cn3F5F4UFI1RBJKN8ANHqcpCLOqG06Dq4U1cjZTCr5odR440S3hBHU
RAltjd3BoJyeWAdfuGQXo5pbUPnPYnLjaye2A7HQsuwP9/i3F8AW3NuQSRkZdG8UWsG22pSavMIT
zWuBNo9tTlAy80CQLV1errO7jLW4cl4JhTMqxjUcoKsZUm3rJCoXFzDKgnzAhIe9FjTCHjQkPhjZ
PcuntZLV/bMQkyZmsITjtvt2hy+RV0XsesF6QkfEovZCeeusndDmENLkjD0l/20Qp0VhcxbdIrcE
RtXc8TwQ2L0wq+KexseJxFvf6Vg+ErpCjPRQ6g48PFrnvDfLRszchs2mkaIJPkRr8ne64dUDprGW
2PyKZ171zO9wQHn5lSPDZHoqXlbhiscBWErxcHy3SLYX31PA9/LaiN87gwa5d/liku1MD/rFE7w4
wCPqd1qSOfxULWKX/xH1/Kt2GKqw9Pkt06/QVRNxbXs9mZMQt4UCJyp3AwBbKd5dYsbsYZOkfwK+
AigFbxbcbbvPVppukXUNi0iZB1/r5l/e+Z4W5BzxMTgc32sWmYhftkVaOMCb8eBAvVTGO9iAhXBa
VC7Vm8xTfb0E/lnNE3cAUXeo88X+kSmk8Na4/dXCkz08NHMs/JG1THYd4zZ9CRDO8Gu8l6aVRd/6
BZqh/fDZbpmspspBB1z9RktLFLl0A/tEIFTO3xeHuS8XYcf35JZAh7xYWGhr7tg126JzwD7J71Zd
txc/fXW3+OsNVjtuAifdoz5SgUHonw3zu8Uwf3Tgp+tmSAaOSFaGxLWJa7DsumK+i+PgXWBBSsW8
lRcM+PaeN+qIx/zXFUjAANha9qRdxdIPZjX0zPSpopCdpRJJUxzvuLslfh+3D3IBJYAc5DwCoB2V
GIrpiB3TYb48eh7T8/QW8nYwAcVYRnyS5d3cf4LkkirQmmeL2m3SVIABjt9ZgUF8exuNlcg9WRP3
TjHdhDfg2YfV6wihjaBWKJaQw/YcM53Ejshmkv7Z5FmTliJYnLZbdWOWoGyvxe15lSTYl74/0ix1
XWlCqExqCf8pYUU+Qoqo0twwvNciCkoSoxeCp2rM7cnez/3LSTg5a2PU4iS3AoQHzv6dm1UX6kcj
BdS3fToeIQpg8KSkzuuRN+BB9WwlCCLNHqKCF+E51PCdCSx0Fb4g4IGFFnQcD7y1lfrglHZAeogj
H+wxmFRYXFy8CmlH5V4Mbpes9G8Gur2FBFcHwH0hyir9I9enwUuBIsCJG2Sp1oHBehaTr9YQttBl
1NyRmJEaiBOPyBQ10nz84SKK3xy+b4QAHeEmPdCvAANhtsbCOUlrjTT0rFRxQKvzJAvK5XSUOk2O
x3D+VgOwXlj60le715nUyZPZLSbxxw90yWqSXmLfdsgTP3KGckMLBOkoU7Pud6OC9EwIKPZNUeuM
3QuDlAkqxlH0pWekkd+j0dE9xac/THgkTUeQ37pGgqb/wLNjZletueJZ6BkjIrwdv1/hwfTa88GF
gG33ps65JmLfSKCVTD6mBN5EvG5Fieyby9se8nIoR+D10i7i+4OwMyv+aTkR0VoN5ogwQperCVOo
oBIJqYs9uEXwOWaycEjdeBJYz0U7+QXTGPBeql82kHS8/L1y4mA9+waUse6ZVGxua4f3o2s8wDO4
SGFV/5hpg03eVw4dMyx3kbiKk+tG9xY/6HH4x2Teh3FMZNMtA0TZmM3NqM4rLtnbJcK/IyrdDsox
c3WhbrWb3jXG/KWPvUsHm6xnYyI0iZxu396ewUVOUlJvY5acZsD0vtES+Taa+YYfh+p5jLDZ+EfV
YS6imklN8WuGiw7oPsVhs/pZSkp3M15DezvRWryid5moaviEzvzEMXdtNvBsekKyQus8NnOIOoYZ
jSPZLRtjSw8tnt9yQVWNsWavp8fy3sAYL1Z8gxt2SmcuCPjLMmXjbsaXHA7DYT6m7yQct0mSbBzs
kRhfD9LIf1lfAlaCCh0u6Gt8EiikxjX6JijYMMuJINFjTdSGfQjQvrdl5mwpykixifkw/5ZxuH9A
VUZQrw2BaIOpoDhl4h0SH9pbj3mrftt/a9J1uWq92McfopBOVJXb4Lpb6bZGScazgMWTtWJNS85P
DxwNyvWNwDIdmXUFXt9Kz42W3QlE61im+Je+25aHZZolLA8uVMH8NPqYBgrK5SKAlm2KEGjS6hgD
khSsCSwNHIDQx/O3tHmp26YpHQZSvDuOxg67FDh+JkOSFnuodGJGb5XBNw34CliETaG3JygL7X40
/fCAumh/yqYgpzj56RL49OlcFE77Q6iI2nK+H+KHqB1XLFfemqWv3mr0DHweKK/Yy8QMLhy3XGHa
M8ZhMp6cIYB8iK0+jh5amrcOluq98AUv1c5niwGiEGIjQhodqo/3Q27v0cjC0hUSIkdCkptfHQXG
QPndlbxBRbUFbAm+3tRG6H/2XAz5REsUsl408JT03CEmiSEkqf7jC2+KkWl0O7okQ0LtIsz562vX
p2INB/FI/jQx9sCnn4YZ0DdywgvzmvkKt5SJiYvpU8cbtqkkaFFbloTzGXL63Bj6x6G5bfvQfh5z
HdtizhIPJsc37TTO2CaLLopx6Kc6pa0XYd2nrI7oDrF5COiW33D8sjWgvEvgeScBDDEanp2a+mWr
IoA27ps+/kB+ahlFRkYi6clCy3bNxQScLUhFHiO1taAynL/30tp/aUFmHJfuzl6QXr1XnMg03VIG
vCKq6vBlkwvxn7YMLFsf+DLz3zJ+RL7yugIik4Rh995rZTYZEjJKzedzqG1U3KZHuEcCW5j22t+8
Kis3Kh6FXsCt3+xE5T7n9qCJtPIF6+NtOlD8QZEom+aMUG6yuaLcujc+qpJp4zoGIXGXnNviLXPN
jGnJxQ3txRTuZUKE0svPXjvoKBMEhrxG8JgfFddJMkr2sfoBu4zXhM7I61MMK4GYjMSFIgTyLD9b
vFIeeBcYQPsfQ/kxVpeACjhjUjm0MdhPraFrO3BDjh0IHni+hz+qW7VxwEe1quc+IM80RFWu5rK4
G3sc1cqEMRjQoo9WjMfGzGmlsfaPN76yaqxu/pQzh27T1G0pMS+qaZ82rput0lx+NHPyXJUPk13W
LQq+MoW1EPDfDWaYtj2cvuThOuydlxFx95EJYEmbEIqL8NggeYDzlw7n5cU45PXQfPFQ7cO/tuty
bYVVkt9bles8kISdXGWw4fxPYCnk1zPMPMQUIt4iZmsIUPaorZvvpDOJz+e6zBlcZsmgsO9IENjk
621uPFkETga/1B6w0sbQf1Bph6g01VsDnLKSs46vZxtWlTzNFVcFvm8RB1m1C1GY499hu3ldZ/n9
51TC74VDhjgaQk+e/LpkFoguMxTpLC/ej+dO5DZ7tapvsmJ+HoaCdT+kv+d0WvQOo40E5JVlfp8S
zbB7VdboPdr5PSiBF/JwkKOq1YDKMRhWXCu1neaRKzXeWeOsh1lwZFBUgFT5TGE4m0eplv0/qggR
GavRLEfkmLxpA8TNBgO1PJ7l8I7d579qNUkVg7TlNvwmim7a+5KMKwUaF3LXX8Z/mvhfkg0ilLV0
i7hkoDqZOYcR5k3ZP1d8ILD/IZ0jEPchpgbBKhtq/17z/5HwL42x0keeEKF5r6PIUhlSRSh4UwJp
sWLkfDFFT33qIuwMm8Mg3K+0rjSSZjGkTIWOUr0gTYTMaD0KWizbvSM/efJNR7Q4yas9jvCcMXqH
Ww1cKOlMyNe7Qp5XEiXe84WOsAJ1JM3CXtirF9rTxflCSvoDn3y87673U7q2S/Yxmi+u/cl5dRsM
Hqrq4CRo7Fn35hQ/V/SvLHQmswkpV3xJA1/hZ7mqUxo3OyH8+W68A95l3ds/6p1+C2U/fwN3CDjj
aLvt4fvKnuIr/mXeZle4GOCGy6PpO8CRXXtO1SN/Pasr0k74ZNGAZnLRUCN5e/rQbDvQ65gMmQyr
RoZ+AYPoySOBR5NjVjO024lvm1Lz73HCPbb+GAm5kKK8qkoaklm7qdw2X2ka4lihwrxoHrHe2v8C
fbINkyTp86nD2gTJ3iYF6HzTcOYg7R2ogs+8OWWe5Ea7Uy3CEbm/RDiTf9Un+jLSuC06vj5/nCW+
zsckQUh+0zyRdqa+ls5H1RSnaKj/x1Mhy7sq23KZmsufSGXqVXC1UHDKWaN41sUmvwJo/81V9bUV
hNgCsNfqmJPbsPwwpl6lCD1NJp0gDAyRrI04rhZG+Qbt9/ObzF9gpcwTb+AjbXkqbI1IbxisBHd1
YdhSWcTeYYGLG0bXt4Je6ORAhQcS9E2dZemTF41doKJivSlv2I8qEI1Xd7KewZErEuvHJtz6IkZ3
Bks4F7vvN1bBtLPbe8QY7oUhkeuhEGL63QaCiWGAw98K90bm9CAUvKGJvUjXQkOJrm9bC3YIASYe
5BRq7nPhKVgrA+sazmHpU5N+y0XKBH7v6ZO+e4LBJAh4tj0m4Y75Cae/6V6LE1K8VrgZYbAH/GXg
IbIPOEY8h3nNMvmsKqCUivb+5mDWv0KOziTz/a7jtDO9usjGQIs03b6bkq0OpCFkuAZLswHtP43S
ztJezGaWxxzpSmr4AuEyi13tlt/sMPLtZCsCeB1RKieQLJ6M40FmLZ/9Gd87iZqTgnXtVHO6EiZI
QK/89Fq24wwEb2/dmOak0jfOKw4AP4qSpfxLB59QVd2p6JlT7kKr9ZdDViSoqk5FVYmuiNt8vXQm
nuUWstFTiNrYtr5pqysVwl4QSckJTEuwJllGEyc0g5GyfH+YbrSTR04fneYBYhZH1QqP6kPA+8x3
/apMEXW98wnTWaqkUrUyzMTWHg/8hMay1PB63rwq74zsnTvKo7dGByBf02ViCxgtIsEaEyZlyrfW
WfNYy7Tl17jmLPEThGoEQsrCC+yfxyrlL2whzcB5QD8+VtHvNySfrYK94kwOq9XMnabGb3GS3g78
IgqI6VNzGY/PCWOIiJLfKHPkn//SNC5eEMiVmXwmrwKH9LdTHtco2/e7wXbF/fiRxdBxmF1AMC66
Ria0vTV7Qx5DwrmrHsNTG//eZQgK4F2zKOjsXnzR7oP02EEuncIiMGm5Vk0flWkT21OZKi4sklwg
1AeNAjOFJm6cxZ3i9jLO3/VjFmNPLyN0T0KJYXyDKGWJFHIjzh/Zy2+N5+22QHJrWQ2hITABfQ9S
AWmodIvfZAAT9coytzycfx3RoTw/grWCYHoKZ6XGXXUMcyNgmfHB5ErcmWRQB6k3SS95+Si/buYe
eOrusMTkpwf2lHWSEqiwOlhWgTwLA5IvVz356acIXPNH9Bi+pez45XuJJ6B7VNhNL7o0KnOWxsA2
RYibIbQFgAwgt/MsQSsiytBN07+DwMOQGQCiuuKxqRMJGOELzakvVQwhJhRY8naxwB+J+ZbNpbBM
tjaGacBXOTOL0UVD5Ile1sQ6pVV7ecRM4myUHHqoHahPLvQymrWAhbJFVI6ImWDrILgDlTdLOyZ+
PafwUzkW6YMvIi+o/DzS9xcRWC8Wikv9CuR3uKOLxwaHgXSXHC4dKVlCno35TWw6b3byMmbXi5yG
lJ7yh8KVIAea0QkP7Z1xGuEIe7rxwmaOhVMm/Cd7D/w4UugHytpepDoB3ef6U4xt4Pwe1f0O2VHG
ACGKCYJ07mlKNhfY9VWWJ/5RieYbNfCi7CDIvQfs3XTUHx9T8EORDk46q0aOFNA+mMZseVHAVv3D
uU/bFvIYmyz4DeTnbezIx6jqdZ/VdoqgjCn1HSJ8D2yGiUxlwYQFcAKjyr0QUEs4zjJbFKgy5kMW
XPJ2VHCZg9KID0hwwEDAr3f3YHE40v61VXnkbJLXHOcqXh4TrIubArXlLpBA3fX1obhbJvXzXQTU
kwt7cNP63LVdFip7MwjfbGoSipdEv1z7IZZ3bD4OyZNvoWmWne5KqvO+7p8kWl858n2wue98kF+X
Q5KWCKqWmClY5qbBVW2PvhRLzusmT2+7yQ7DPhu3vHiqxXhpJ7IQJ/e/nQBo+7g1BCot50EQq8oa
hpefaFEmsKjMHwnS6w/Af1c9BmzXhcREDlGiJ2XN6csW7Sx76AEsZIHGHv+Qi8r2jPXNiJAmCOQ/
44tVwf0fa5wUGJVjdzkIhiqKVvsrkvHkccdsyArcc5G895Co/dD46p/pJprzPy8me6ZMQ1mHrP4n
hDyNFU+yN9E3cHLl1QzpB3tzooQJkoRYHNXSg4yTzmQWI4WFBDeQK8CHOHF3b/NcYw7UMzuJWD0X
etTGzcrI1yLx1Kabr8bjdBoVtploZ3rIHSrrWfEk0wy/ypjBn5bjDD7d1EwAkhBJxvmPCgBmJEGq
X6zNopYxPD+oiBmuud8SlquReilWsou7TjMNTerEnsV0rJLrEsG7+DmsFrik7gf2nmCgwSaF3GKe
SGNBCh7M6gZof9cXcy7xiPbr9zvTRF1eFyvcG3XVlaVO5BnK4rakBni7++061Gamu/F71U9CTCzi
BEkwTlhW2Mf8BpPp1x+cHxpwFeWjlZQm+XYowxiYrMm3+dk/QCXbBaOTaN4TopO/8XS7MMZKhEGr
aNxyYF1fyGB7PeM64arw+58qvQ7OXdS6PKYvMY5FSKLOB5kZlvdFTPDjW+aW5/OIqvgyKT9ex9a1
5o8anzemvqgUEDRtrW0hDGQyZ5tWmPCDJeh1JPd1D94VY1AIDfSUnQRA7oj45wGZ8k3Z96CeI51w
Rqp061fZvYQgd64sVMUFkO6S40olGW93wCnd+xBUsGZqHNkcp3UWwd21htBjqAn6/IVWvNlv/y0n
ruvVJvm0THv00GPVggBwlH0lynyuMwJa8UcbvlNITKeW7t32vt+U5fHLGaAGuDt7ONT2khJtL0Ss
myN9ZDoX0AyGzYKtPS9ULgCpDnFdBKexJInro2IlnFdfI7r1q5tOz7RDNRkYPfoG3iURpaVMhyub
gepKxbtzv8kwscbsZw/0wbnIaKiX1MKZGqRGqHpXZ6ifpIi159D2DLwMtp5zOSjrPzPRkDPZeHQO
gYOOvJIlvpj8xfgVNlSPSpPXhlK4CcXvd1gKLn2U9NOhtRbaXHYrMxES6JNRtuvE60k3LKC+j8Vr
kOfUjCj272EFibgeK9qnd2M+WzbLdgYz2B3MVXicfn+7rDKR8RcZx51/iOtDsJCKmpAA4D3TtN3I
v+xmZ3zzYbSuVY7aVhSkOe10tN/mVfmddDc/66v9WMnVmitF6uRE5OZr16FtZ16JPnIm/TsTZqGy
27Ugyp12uk/RZRBC32kqZ81XRuDMPOtwMeCWXPwMnmb1qQf5L+Y0+EaohdEIaRAeR7rRLVus7qZ9
aydlDYSGvPHmEI5jIbv2Ts6dhls0Ug9MfXTPmlcUYQ8HVmTmfUhkIGrPCVCnXQTa2UintqzD6Af5
Jzy2TYFbUxSJkAuL0Vt9PGCtDsGpyWV6Nx47L+WFMoIFkAAcku0qKlta5jPTgMyqdUaXpEUGJTrU
uK+DTlHpQjrfm9c7WMMDkvH2pwEYusR1unv4rdbos2H5pl1zKDY5WpBeer9Bu5TVBIS93zDUn75R
qrUkFIGu5QJOheFbUIHOvzJ+iTklz1hLjTM8Ufwcmka0Qhp2Vgcr/4LwKGh5gy5G4oRcp+ZAExyJ
kn45EpRISNsyqwRQX/TyHkAESwmYDGDxNs9MLAv49Z2+cO4nytTDZ1yqlU5fYc/xBZctRwgNX4fL
BMkDytF7h3H7sYjtJiN0BIndMTfoaXYpqA9XIi77ImE8Xg4MmOt9k11Ooh3JvME4NpJ4vHth3nWN
2ZKlDytOjLuDxaV6Zf3VLM4xbeVBlAOhBykZnEKwviL2Jun2RGzc550O0UNaTLhAJgjZdfwZHIgu
ZYEj85uIi2Lhufyc74ASutVzzS0iHyEDQIv3fuJyCfU6qe/vmknaO1UUb3sQgwYppnTCTKFp/Y0y
EnuXVejPcTW/XtyZzrGreMsLueSKE655dHoT/zv0Mg3z2W8kcwvfyCYDtIMgGuVqWj6dvu4eBxvb
Vi5NHu6s0NbnedXHboAy6Kb2a5TZzE+GNgzyeWJ53fXcqfYEmHvuTY9U/hRM0CTh9icPD78f1+J6
G51jfxA6RjiouLLpsf+LF/ZHVnmqwtAFljInSjouZaEvPM9yATrlJ9wXDnfZnLx9Dj49nT1tkZmh
pxPJa04SWdv8RFloPLHwwXZK9ef7fxtl2caCAdIaI2b/6bd+p3mvb0u1jIRGP/c6Gtj0s0Hyl4Ke
+R1QBKHP7PNcKyL3aRXXVQ1pmsvxGr6XudJveS7r9I2ZMbx8y27L3SEXZyjQ8b8gy8B46cZw04Qr
1l8Erg7T2DYeec8EScEgT749Edce0rexl9zqR4onSYH8uEjwqcl+oCopcWqLijcR44OipetBFgCF
EvHATB7StiZ/gh9W0QFCipMoU8buUTgXrWoIXX74HAu4uvgzbpVQm7SxqXTxEhBt5qOIJTU/VLxv
uKGKbwsZPMGgBHqu2IFswt0JYcxOQ7dKgPW5v8Dfg6dqSjwPmWobPUwSREFtmrxhlfnpaHrBguKy
1shYtpkU5/eEKSv6bkrXZc2pHQGonQfGAjJBP8XjHVm2hlOZDe3A/az8f+8HsSNUgBJ6HCb0hEWY
BVj16eHvwb32RP7sywY6rePlEMHblbx43cthQxXcCtm9AlMt3GT1dqfeR3aBmZoXGXJkKf7fOlsy
JqD40j88EWJaEQKiRq+2X/wM2OLGB8I4NhIy4Zc/4lbtNZp7M7UCbgHcE7jMh0IMNjiprte+0IKL
Vmep1Xp7ZHtPBXQ3K9zZAptvZGOLnNW5A9KytRIavakecZxFkGfJvWm+DpDN60xj0RAnowudkWs2
onN/agJdGxwNp7IDjqrhhOAIx43QOhaz7Uetua5rSzkoCuadlOpfWJIdw3iDMakoM8IzHu1BxBgD
s1kCBkV3AgusscpnIGWa0Y8aSUGJn7nkG1dLJwoHSr1G0S/8NvDInn4HemS+o7J+XCUhzGTX4H+E
1Y1CJMXYDyWc0CbtpzHZRwg9mXpojIiGV0ThOxmFG1eQVCg5T3XAwz3v90d3NRv8jmc7yeDTqZkF
bf7RAQ5Swe+Cryoc3eWwWcq258FgWSTWu6IZzpo1UB7FnVoapj1Se4Cf5iVY34AsEqwcTVjR4+CB
c7Uhjr/usOamxbMl3xL/Pd6CxmBAL7lU+QunrLIv02PR1xt+Cmev6vGZgMINu45HIy694OMaeZG0
6fvWYuedg1IiWcZ5kLtan0kqBUmyyImB574Q3esvRN+Knxr/ul2YuV3XyCOo1GeaKEAqPSsbwRiG
j30mYINJTCXkm7JGrxrQ7uY4690uqxRCymH1RC6mVsObRo9m9rs8veeLESi7Y3sLRIIjCh+RKxLQ
VLSEFRZ5uuhJPY7gzlfwd3QvBMfbBJ70KpC4JFK5URGnq2wZarr7MG/xFee5c7j2tiqIlGZu9ELD
51pkxtTDX3L9s56zBF3AEjnlkZ+5LNg1z+i7KJeADpnBQ9MehFKPhyUtFfIn2orHjJ9g+Uq88UyT
3bWui+hnfNCY1+G0JBgxb1ajpVhbG5J4f6GOVwJtWoxRdtN8Z8eat7tmTmrIdqMW2w/OyQ7oqlLX
qvztn3obPAHQFJWgvykTd1waHb95626NXGao+eS6BBbR0PAjmQlE89UwCE1sN9+6HFrvXingPJWd
PE2+B4vEuS0CgJpBe6U8rlclnPsIhPCELsx0dP8h8uZyXzozWtuSM4oYUR7gEaubL64PtMO0n4J7
x2aNxdCWGo8gYxppB2lg4pNSHBruo/SzSi/gj4Da6Pa0SOeS3iVTGcWbBLL0+8vaXS2wutGBVjNa
CaH2lhpt5tYAje8UDBUtRnMuqlWu5AL+c6YPUrNFc8+xb9iYjposhEd4mG1zH7rwX2Sho9bsBQTz
Oxp5lXDLjn14eHOoIOuM+mGeVpkA0yIArezE84N/ddoTOtcgbR87hJAwJnqQgtXv9TOufgc4/ny5
wNpp/eNnDGgIQkNQ1QBUlYeFPIq9rxskU/SBmDoakeYRO87jsjnugDoitrFFX9xDnQf4xOQGiBwF
HXb/LWnK8UQmh/yix2yTglmtWg3OzMOYvF2hZd4rdnrQeX3to8px5937UitjTnMtNzhCwTpUwD/D
Vx06PW4duygHXlIHeY7Onz56pv8YA5BX3RCnDp8zFs25Gt6SDs7tRODIeZNI3onW7SnhJIIjBEhF
YluSMGI1TV4q7sEjJhKkEVkRIZXdBfFTeYqtQN8rCQGi5bFmLwSjqMM75GcTlFO4qoJRa00XyQ5b
kkb7q9J3fnBpu7rB+p/JI5CvjkLrxMQuSjL3lIERJ7ZX5SQEKKupP8dSGQmyUjDfjCqu5we3ATjB
kDe2BUuSeiTykkPoj2k+RQbHpfTfHmO2xORkosSvfzQmEuD7xX7QeHkaO7dvKrOHqef/dvgAS41Z
VQtO5OZ2XXBw5R6gyZ6qvtb1rLA/6++7bBSp91S7BW148zVna4BRSZUh95BRLcRhXg58KoRZoSPi
Pc7NkrHvc0ZHbsi4iBXxICbGlDKkMYiawuB3JiK7d70PQB4JBuHC0Gb3Lz0Ju7obLz43XP7uPTa4
B0jEck/TMTaX7GVeVZAUdvGyaEF06jzlQYTNUjuTcosE6lmT+9K0TVZqAVFqW4ZivvMuMCut+VT5
MErBhUnEaLhUtyp8YFzs+BO7lq44v9rexPRSlh4KKm6wrSzZnUqUrn32ZSTqZg0uLqC8HRD1LFk7
GF/8cxahngRZ8i4gSfqF09yfDtS/HuGX3ZD+vICReOoIEGr9wfxCBMWGfkm1DStlW5ntg1otPCWV
mVoV3b/Y3N2DLakiILNSy1O1Y8+inUkgVxCSW2+tkOdHL18wTPs8tIaWNRwPaD1zJF/JzkFC2CCK
3nJnqYaW97NJnhLLz266m8bul2tS8SIT9+OGhBqKlRidh5ae54PicjIsSSmKM29zi9ek4cNF/t4D
ZgkcBW3JjqJ/lV1SXj9cWetMp/l4XynQA+bzsOWLIw+EKFbxa3YZwtnYiDYhKXsdns2rM7/ru9k/
v1urDP7+WiOapT+EcVZ8iQibKcL3wYOm3NV0Uk/VxQBXFalpJULxkLqpKUXK8GHZ2KnGkshc9ZWm
+wO31NDgPbjceLSm0QPbq7fVg8pfyVQVWtNWoz2f+uKdaBcz6RhMg7BLz84mb2S2thUEbVbvmOQy
vpmoi4AZEmUt1IzUVSb3PVFaecfQFpBNtkSM3gIoH23BuLEwCJ2Gu5uVALuCqANkZZc0oGCGJBTL
B+4FGc49rKkxyHXKFF8nQBhp9ng1ThmxUqkEPAlx+2Sz0NssqvC5E17DwrRRc7wlDohNOwNj9y6F
opmBJnK5cA73nhSwLqQ2FFeLrNpOmzyWA4qyOA3tUeYwKo/Hjq4L/SSN9pHpPRk5iy/yJIRFq9Az
JWw7zbSrpWWL6vQydOxcg+nfJgp2UyOm1bpxMRwdyDEOgMQXHCTuXgFivVxCR0ejq2gubqzIovEv
RB0hZQQBr45eb8y8rzH2CB9oTdO4kKDfP0eURE52s+Bfq0j0HGeg44vUmZwJ4gHyx75y49ee/GaH
yL/+E6uC0bPoKXhh0ffIkH5ny1uR9o8gNEI/m/ZFVHfSPT75qPPC48TdboHTTmSKB61BXXRXgWMh
5dUL5+eO8VeBBTdjagK++Njf2M1iBppE8MZWVml70pRZlvJc0uBTvlEVENltUGqyj6FZuIIu3djs
TwoJvE7CPkh+r3cTvFrxsewoBy6TT6K9gtjK5cI6Ws35o1mTkVRbxBP7Ec4P9jV0Ner5JpiYYZen
HHqGZV+wKjXE9J0r2V9VTSAippQuFOCHM2YJ4JWkMXvntsWkKk/x5ZLMfj9RwaUw3fUBdlCySq1D
KAZHgmQKtHz5NcNkJldpF0OGe2HBWD9XRHN2HmfXS/ItO+KtGQLqA889xAsnce6o6l2wjSoXqgfn
XPBEI+cvT0UVvzY5+mA7I8VKDaRUKyUbEdX5i1DNvzhquvGQuDeAhKrTB+F/75NCusUN42GAAPn3
Bwj92h/BvJA0B4urxLP60ykiAGlg7myAnp2Qtt0BBLJcnMVPnA76JvqzT3QkgcezayRYUpjf1eIg
vb61QzVFrWHCmGUV4bcZzclEILv68MjCI/2oZFkNwBYE6HPe9ByJfsWdy9Sg8LszG/Pto1bpGklb
HMwyuyRfwH7vdCoxYLwwY1L8A5MOg3mokt+s5fmkIayiE44qHs82US9xo9/Q7jGzk+ofzyo1q1yD
kHH70WfxB46FEJctom7y0ZViCUHp3VrbV2zId/up9LhBucQXd42LhPuuq35NWVIy5tRdC+r6V/Oj
ghLeF2ThYBZ6KvhjcPKof+tfmYyZXTgQocBpHt3u0DPiYMe2XOBBnYgYJo0FAyqkxE2lZBDaR9oj
SOegYkO2O7iPvYXqzay/GEqgngItlLH+OJ9siwMRkGgqHwVlE0psVZkkWjDa/BGfYt+YBbmlY+BG
b14kaJf1AHvAE/35w96MK9M2FAZZP92X9qaH0fWtL/9TLFpJ07gkhHXNd1+JOycp3JjSwjTv6ziz
0hTmFuo+sTwb99yv05JMyx1W6WFMtDMLuTFlBSMs8TDPEEsmymc7veEeJOhR14gdhIJtxv2luRxH
skEM2RNU7HGYuOUwg1jJLML6RMTHg7Lb+OSUpvV1N3avnk6b+UWrh08csKSYdhO4mMWI15WpbuwD
EXaSythGsAzIif6dq9Z7G+XFNd6t94xLtYgcVkXSKC61jSob/Yf8PRdGH5gs/ZnR0ZK7hAhFC36Y
DYPRM5l9GNaDBYwWHkU8aik6p8kZrNyXkqeH9Gvv0QuMqp4NhsteiLFFx7ix4GlL4NzNKwEXEdoo
HP8uE+J0RiflhP279IdcHzM+og9EYxR1SoYkVA/+HwMFdaN6TRcxNjaVScfQ+HnZ+I1dbhU1OrNy
24yM/XyGFZ5VtY/8DOsrsp3s0BesMa7nIke8STzeERPMwlMIJH0EY6hdfFR1tbHjry7P61X/lEZW
12QMtdQkoHuUM4HyoC0atbNKgUEkbjbP4mqj6fqSz/eoeTeRmvMUzJF40pvgp/IVAPq0YbhQjTh5
2bsPFkhMfZbVGoSIP5JceezjbGB7N49H7LVQPOGSDasY4ITCc01ryVKFv9MtraVDv5CJRHY8sUTD
h3zcUyTbRwfnSjdo+1ZSNpx8SG5Qs2a6MBKO0J/uNt/AdkGbW6SzwJgrhJBY/AnAkQCf3WWWjOUh
fmm98gygDRj1iy+8IEmdSZy/YJyhm62pimgaIrhKG+iSmpc++3KqfrTa+qgBE/W6o3Nqky4LuU4r
lKoOx0Pak0ulIUt4D6WtG2eXZuwRhQ5XX7oLdM5Fg1TZ3u7WtwYru9Ui7UkN4EyWoQr9FisdKUsk
K4M7+6eBAdeO12DQnQ2fOFEioxzSdFn4gXcVC8QLU8rQDJEQAIQnJyulGNUKd8Z4Cz1f4TjvCFvp
BC/DNeKifRB2vYBgvHYe0SFFmMkHk3/3SrS0F2Y1TD7wmIe6SNdcVN69QFhwByjwXK1EMe56PuBx
+fCpGV9T1zd2al/TDp83CQiKBeypc88EDf91TL3xRpsaKTlFY1PvGO6F1FNQ6FQkjIjIUI2eF62A
aC9dzOkCFOdSwaqeU0SesLSm69zRg6a5oH8hlFT+1RQXldfoup5dHGD/HoLIanAMhyKdU0y5d924
7WqknMve0R2pb4o/giglLWOcCs4AYeeSUotV4CBW/+KZCd4T1w2vxsBxw/AtVTIpEbDQFbPD74Cm
Sjfe6DjkQ+GpAjMWZ8vwVxO56EgYcnn9WSA7mJ5f2/6/kTpV0DK2QIrJiQPmluDWGFvJjkh89IzZ
nHM2dGUqIkWMS8C4hO3N+rPRVlrQvYnNigHdz3i6WHE5yKUr2ezK/bYw5unPMEZ9WwN+yvfdk79w
zVst1Lvm2YujCmr/z7tjP8J97qFrLvAWmDRUDH/qSTrHixxqojWhvwNoOQf1w1r+x2mndTPLHz0k
xcfDFzuQelB8ZgENmunyBxLmRPRAD9m0uMuiWP1npq7xnucRfcKfgLiZbmn5AD+4etkMoAlvCxed
YXKUvme81RbvCLsaImTMdKqG9hgiFvTnHPfDFkU8sZCpoDQX0/D+FcS3JPu5qKB8KYRZ9OqYmgzU
i5JVOIJm+/bYAXRn1WBvf1L9C6o5WGVNd+koF/bRK4fWlnvcIWHvgzXg5crr9RU1nbUfxkFdm1ct
AU5aScQppoUW9vXI5yZH/tftBCbDBscZ9tKkKljKPTdPXiadECLEVArBrXkrvsiHjnrTn+1xhvLl
6jRV7HCJr31fJX8kFK9I5dGj/JMSX13n8h429mQmiaaMzDtEwd2ZM5IwiIgxWhkiza7Hh03ynfW3
f51QkEIC1qYAfIEwO0MGdRVYGNwnG/25t08FIVXuHTK/t1+nd/UB51m2g3VbjGbHaMlbKV1GTGut
XgPvJQRbCcf30R8WGIoxNQKYPRI0eM2o8PaMjGdS6MEiQhmfT6oKZDmMLMfZsacjyZxGIjFZvy/K
JV2F4a+oXe9dvoq3jmQa28BoABwRIpiZlzrU/1SR9SrHJK+8C60cyp/2KMYie1EV3HDvxBBPG0LP
kFluJ7xGZVAEsGVh+WeYBKB/DyDMhplZLBGAlJEXAW5TDZbq/+jbj83K1dhv253jLu46rUWsBQ2m
2qnnAKhArmH5pVakwx67+i8lOUOQmySdT8p8ul8evxf+jjSm00K0So6Rt+fo7F/gnZc3G/xVnFPk
ltycB3LMjHra+K1Vy+/xn/39BXDB0C6ozsd7JC5h958qDzLFgvsVAqHl11/Jgxgw0VMdvaM8Lo9N
tU9+Iobf+KI4AL01ZJP7TZClwqTIp7TZuVqBgzc9v8Hr2khG2aUkhOy/r4ap0elKSCrKNhNj8+MB
YkueGKwctQOFzQUIeVnNUh5Lmf9KdGXrexCjHD+x5x7oPAVXDM9mstYo5hsilBkuLUbPNsKo1dly
chWCRumQwPKxDwtXG4ZLPURB7gOiz0lzpul5fXzUYgj1IsA4N7Q/56FECdB5RinUyoCTsEXE3l9g
dqcR1Dxr9Xh91Oifo7QlqD7o0W1FzIOaKbEkixHaYOzB+ed05glQo5WuYoIb9SHQ/in67/BD5S/F
GnNnzj7klUzSEM+ard3GTFbnpkmSAqkoJ5i7ciLbxfzAB68JaySvnZlADETmTT/P6vqv5R9R1uPc
zrrnTAtFU2F0hoKzb+WCET37sA6IGqGeY7mw0CbK4i3FXL9tVxSHlS9M5FWq52yP7eTlDwU2w8f1
mbJVsgkJcfDrHIztkK+xT4QUyi1E0PRtcp0OqV8avnCrlI8WILK+U/4hGNqtsXyV9cJ0uggN36jv
RxuByzreaOQ0G+VxR7yJN2FqmIiiom/7Ne9A+NZfSjvAppVPH3zbH8GG87J180VgOxlw9zMIfPKI
I9C6UWVNgPxfBm6oRw511/uFcQyv6jgmAYNDe+81DIptUn4AC1jHbxKUzY+Wk63fJQYZP+s2b25o
ciPQbvUmZXcbL789naNzedCYMThQmF6pIoE4c1aK++ArrJ0FxqR5+mLW7jTkfEi3ZZ7VHkIoi/GY
gXaI6iobHKg2uSYfLUph/y8Kz/jDbNjY8PXlQOp5DghVO2kkVrxEJi/qLzZpho3a582WZ1deN6GL
R6FXV57nJjI3bZLPbrdXGwHbXzHLUC4yGNBXozGkvmepF1gGZkz/eGJ5F0WORjhi6MVhxczVzl3a
j+qCgKVztHF2z9U8X+gzksn9E2f9BCA8NQGr66XGmAPSTgoYuFwwci3waEQar9asec4VyaMHCCvn
VmJuymHhD+3ELJiPsaPRYDU0K6xymKR+9KaJIVFFcnvRZ5x85YfbvJR1Y79f3G6L+k69gcZXX2To
1r8cHiBNyK5W14uncoZXxitfG3/9vQHA0k9TSA8miM3LCPZGSJT3h7hDn/gj3hVEBz82xakHrFqM
9tlTyM1NHq247nOzqNcE9aTDJVAvpZ6L3DmMfaAftBmjVjWyf6UXbwFytJeAoTckG1MAfOJReboB
mK/nBz4IubSvnioZ1qNuz60H0Y4TWC/mqN20FW/vCvkia6Ray/9hSaZWqiRlRKjdOkRQp2yagLrj
/V4RSpkoV0eogsArxVJ9RpTelh281heyBQJ2eDBumjd++pAQatA/hh8vRyZ2samOOJJmtNHDChkL
ETtEUzyjk9WbL5krVU40P1SboifgAUMHXsMpgGoguYviwcm42jd9Uur4/6BylDkwcpxKMiKk10ka
lB3JJPZRGfPffHbjNIjrlG/rRcpQ/yw7JuuPJrZoRmv6HeodifuYPlxkY7r/Zu/Psuqc7Ofslt0f
TC659iur14xXSwD3SdlwRcjXXTMShtBVwtYJ37fXnVya/U9rNkTmEDTh4rC2+4jwfY7Wm9pJ/XzB
cfvw/1p21EShC4XAneEtStdogyWErJo9liomXMCR6T5BTUcLLpJGeAtew1aashGI3GlDEfaearJ5
kYf4GQatbWUn7ux96dGWTByFsXsU50LMi0FKv4Wqu/0N4dqAY8ujeUcDV0Z4QdEU+CMcJd62KGYS
bDbgX5u4MbTg3Q0U90cMtXFPxxJfmW/T0A4zolIVi31U1CcYyPApVbnDrTLJAsK1EK/HtBI6KPDd
cpVbJxh3xTQV4LZxnr2/5fA9EJP9pGbCMP2GJs95pDBrbsTcvP4aq38yOqMN6eljVWUN1HCbbfbI
ZDxWivHWV62EKmh1IB1hAKGbwu00r2AyOKKdXfKxY1svM9oh3ek4Rn+3duRfTQkFg/ZcSjY9KZyH
yA/Mw51U2gyLQYXMwlvplcJeFee0EcZmGUH9JdywvzoUt8H0iJwT2Y6vIPKV1UsMiHCxZzofQKWT
D0EnhC1uNYjIdDAMagT+tVwRRAbEW3WlEe1rgQf8UPVH6abja5iUrJdfo7TaEpAW5tJrkFAkOTt/
DR9hZZfOIVuP7urcMvz4UbgWPP3Xe5MyKROeHSg4dVD8JRsrRJx2ADE3wzCs9vNyfiO0/QT9oQVy
0e2LwBihGCEBAgNLxSncFayt/KXzRwLvHvcJB57vxYun/FMBwJoIL+dj6bPyzxhJpHUiG3sTIIAl
gb/Sij69aQFIeDiliPU0ujpjT49hY/YM12X5uvbxSTiOG2Fp3LvSGqfdXPPjVvLqaHq6CWGaj2VE
VO1hLIKYSfIjSCLVrR4CIZDzIYiKOucrifz+Jqd6htPUMSMgzxHq8EFRS/USOLpBbXRN+h/oEpcq
lMFQziXqx6/Kz07yyGNW9eWwOn3vy2I9dsk9dVq0ifA8vQ6a8wBWqOIJ/9b65oPFdsIvOejeFL73
pxyjGdM21dUOMFcDzaZ+qnr+0Bo7f9gUgkIrvXL3aSxJEBidkKfHUQEdmNC/dyFW4p1gmqtXGyTG
qCEhvm3ZDUm3Y3kd9E4YdZJOpkhb5+dLXjFWMzw3fO3d1I1zZbHnX53iwCebaA7sziN8/SAoabeG
e57boRHsSqv9+/1k6v6lia/WNwJV8D26yCIRXkLdh3vbgMuaWAlCVJmb5QUpNxxlmOWJW3Y3uMEq
PgE1aNXkFsUTZNRZLBPY+3Ahr/Axl8wsU6V25epKN7QXNb0Pv9Pp3aaIZt2Wu6gn9FVpXnfPCl0/
W5StGdF4XMqYFvjibX3eajx0nJkIV6xWg0Ts2fORnO6KXW86Pr1/EIUsIJDrAHvMQcY619z4PrtX
2c2/DykmUkShVdGbejiXiLprWh3eHgSMVlM0w32gdKJ0a3aRMw2mNXgzfRnBnxCIt9TTxClyWpuV
xt4PcfZguCJOjLTKDHe3oOGXWIXleRTXDAgCMCK+U3vLNhCHUya9woogsEtiemOmnJSY1Jf6UyJk
aQ7S6iBXkaeo5IKapX6G7B3S+8u++PON7m4Id5+iMs8J8OHl+dEteHJS56EalFGOy5HClDq/8ZNg
webzZhCRyF5N2x4d4lrvFzHCQnNq04V3NvIKGqINng9iAxnwEioPqTaQIG/xhsAR9+6hEOXMYGs7
Oj2rgKglf8SpNWelshDOC1ZR/dAs7XwgeMQPbvG++EMBnDu0mA7fftddE/Cj9QEercKg9J3sTn/Z
F3hIzZErqZLPOX+WF+G0PtsoSrTUP7Qk5C5J5NWr+u/oX8FqarHopbwDTaScnwQ0B1TVPciZAize
+q2JaQonGFFJ5Tj4MixAF2QzLVcNYquF4fwRIp0YdTwa961b+RdC7nq5FJG2WK7skyaePC5/gS5H
xOIzQWVEAbENdWqLjuzXfU1S7afjga4c+ihY4xZx5lFKSSeG5bpjG23XO1BsUQ28N6o264zg3f/u
uJ2PA1+i2G9q0iHrrRjqjmiGV5xrdNhfpcPKhT9cedmXzy8xmmVOa26g8F4jieKvyOcnHK22WDr0
wX5jkquc9FCW14AOln4yMJXyGk5XpakHmjuyKn+KMIavXnvTOnbQW7P86eEoCTuk/Ez92lbTi6bS
DT4S41+5VsUd5bpe+UQs2c5IWAxG1Lz93Xq0ystnqqoTb3OW1Zlxep7BJlXmn2T54nd5waqJzPQu
8cdKA1IWHpvL9dgEsgkINiT7vhIhLSUjPDNj3d1u5jnLxHh7fnHKFCgrE1qAAuotA1/0QP5Igkjx
fjipy6JzymtX50h3GbS9y8lEHxw0tf7e4TdC018cbHRVS5bQpxbfcR0jUWF+t1kycQPaXBxdJoIZ
8ZhRwVFTln4xuoIiIgZ+YIYwQo4f2wqZbupBZ7jmU6VIZ3lr3m5guledGgLMmVetV9Y5RtugNj8Q
lnkJpYIl6cEQpK74zC8W1IdCrtVP7WdlLzEMLj81AOYuJ1V2mu5FDdnRdzGVgSR2DjYTClQxmQRD
FvfC6s7Ak62wr65SLhVcRt+rcipY546h4xmf7wQGKoVfIj+M0tvi8K+4y21+Nhw+Y/4WbsyXK0kW
ZQ2dUaz7KJPNLN+nPz76XR6yr3FozOz47Ge+6BHj1v3xmwTMhbGKfVq5EPFMAP+bZ+KeK9y0VHTt
qTsTYMfoFflMJUjbLN/NxG8w65Gk87/6bRe6uTxhTrFSEUnWJmyYINK0QrEQQd5C/HDmJAw+ineE
MXRUG0L7LE8fjzNkt3g2k0lLZVH8Kx1dW8zZykRW4NvkJ7+VZx3pwftuFp2TqLvce32fmwIR3Prx
FFPTZMAUHCIRysBxZoCotKjqkXs9MJRAdF5Opvn6HUXp/fqIaZD3/WSvzvT28D++yq4w5qY5hZlB
jpf3hKG6W1lNB/Fp9YqE3RriZn85UmENBTHUrZXNhRrq3DAZKyKLZnz+O4D5QvlYnM9x+sXyBzuW
NPzxBL3v8nsGwMUeuSCayiVE6bHjLOsqskfZhvgQA4unSdHC69eLLPEL2+3O31IE2Gi4+JebrFLX
/qAoY8CBjkaPXM0CzRQ9TQJW4duhhGJinnDwD3MKk9O/HqC9zOFMk/qTXUim/6UER8i2q1pnwYhc
6iI84Zn3nJ9PhJ+CXP2W2r2ft5lS54S9OJGBG30kgMd6ZQ75aRqdYqtUrQa7FQ2Sx1LKpF7G28X9
SSbusMN4Zjd+iNQdw1Yw20oUmQF4G1EtAialoQK8GwcEhzZILXqQiScB1Gyx1VCyVyIpeN25uHzm
DFvkRDptAuQRmBbCJNLNzr7VBD9XskgBNSkcvrT0XMRA8JZss8gTmHb/geGmBODzN2/47huWn90b
2L3gfODcvvMOUaYP23sP3H7WKGw9Prx7IMCX/DGxAUEnWccyOhUEdzH4uH3zbDkv1akvu/LIVKNF
0qTykw+AJeeEjWmn2ZNTEjuKWNz5NpN11jWrSjhbFvEZYYedaUbmA/1NKLpgdyQ+JNuGkfESE6rL
qW0obOsaB2c4BxxdzI1X6zDW1xPBJzGVaooTYesh/B2Yv3ID8ImFsKaPeJV/xd7JMiOO1d7nLIbN
beKzxnRze55pMhBss3GXl1I/nQmGwuQ1RZuGB3ljlU8AiDJ7Dzlqq1J1w+n32R5j5EL4kMZvwb2L
O9BbJGPubTCFXfPw94v5yyuG5DTMJtvUGZ8m/DkT8j4W5CXPHMPae0svSyEh/MWrU2pBBfG/xDSQ
a7E09cxDO9VhzgwpCURvrYTDHEf0pWtik086krCGZpn3O/GcJu+Gfp7bLyAPsQwdNQ8tcYihJuE+
8iUoSC3B71SzT+CQjvpOhwsyYJhXYIVQnXtGKejITgEHP4b9DqgMOmYYLr91/irjiZpSkMGKWolc
yNyBTWmDYK2pWhDYsKSWT3lZE97F34xiu39eG5VmWL5FC/CzJl2BJ9pVznjxMs6lYvszZwMCmYpd
V5HJXrFdXOa//nf4+VEC2tjL6y749b9E9AY5CkzhCEJf5BcaqyDsNZS56I6xYYc7d+mbjpqc7WO/
B9ZZN+k3xM9RcME8RpBdiUwJbTksbWXxkQp9ptPlgqNIb6F21MtUY6KBFafHF/FB/PWqBFuGudw/
w2AgHEgp6gOhLjVn+E5CVX3NXOcg9OqAoiuEOGF6C7E8lza/W7KTwrFrsIZM2ZXYW40o9WppznWh
V9uufo75EJYd9282iLywNbu/bUskfncmvbLmKfQm8SRob+lTNp6a5OwXP4QZohyXQXZl7Y3BNJRi
1OclluwP+km9HRP6ch7VZ0BdJEK3xQedsR8bsyn7R9Lq8YBZPMHMxD4xSp8cxhwoElSBCWADSBm0
CrDzJGWAVp0boYyCzXxhY2xfW64hXeH0ZZV4iQ6chdtZ4/x4QIENM8sB7pV+RLYFuvvu3NtsaGok
6GG7FaR4fHIh5mL+w9YTpY//RLe9ueUh40CtebhSZ0GT5yPgkxyMY/ylXtH51tLYLG7V4TfZAHj6
HJWvJBIdRRYA2248TJpatIooD32o8HhreOYwFuEOrOstetEOrDVnsvwJkE8d2mofrbOemrKptiiW
GPDeaXiGIYyruqhKpmZeWmOiu9zjjFJlu1E1ob+yvQOL4AFFY6RNzlgHy1si5OtUKN+v8QmKkwmY
G8e8xEhtFF091MiCBl/xw33ldrc6PYk7sUeaBlkKtXBEb7ac8UVAnCQVhtr6bMJUWoaaev4Nx+/B
6Gq4OtrNYjWYpPG9NHijURO5sC0nY2v+Q4JShZPAZtB9tMfybdODh/17A2dsE9/lXxwKcbhWy8FM
J7b8XIZeihPU1Y9Q4y6g39Jx92s39R85M7rHBY5tnB4nJuZMBjv2BCYZgeRMc0qpBV7df3KqKt14
PhOXVY2kXWShakBPUcNsDTWHbK5KFooAPV63tArvw+TFT29xNTG17oQJQtO02MXAFMbXV0Jmrp+E
83WCgzcSngt9lONpmYmITB8YeHv5s1HutfhHt1qpgpY157THhEFvalSnqkz6oBc8m5ZoOvFXwB47
LRokv8qCR0UzQ+IjpMYBeSNicxCHZmH1gFgUnzwqxWncnmRAPHxWPtbUED0xXaLoVfNW+XdMoJbZ
OefKHtjZGPBzmyg8OlOXnxsBdsqupYmmNtKEbEf+aCDBQwrSkEP4uFt1TTIIGi4O3F/ph4jTKwcg
nA36Yw4H1b6zEmOWiayIepeoNRLalfEh+IYuW1P5iVWlcr0cmAWahi4igq3BOmC53I96iXBGScQC
wTxi//jTzPW6MTEo8N1vxKa44H9k8i4YL0FiWg9i8k6H5EJxkO03GxX7DFtqb5v5yc2Xj5dQMlGy
LrLG+zahv5oux7sJmqgdUo7G6m06s9e14zlx+Q9e5GL51Onzv/zsdH+ycM/SVFij/CKz7mmXmVdu
8GFkPACN6qnwhzY2WydsAxIxDX/9Ad8buwQsW3+c4jpiJ7ZLJaxkUmerbf6q48V5OI1w09383Wcu
dQnilePf3vnjvvMGG2lQ/ILzVCGRpkqfbvcA6YHRzSCM0EGOuBHp2YfWCRf6EBffWwz89lkJxKUD
kyFedzJ8IBXzkI/TJxytx3RqJJzWwoFNMIBdTRgcWzaY+ZYS88uslEcLUD2fq+r2lW/lclhavLGF
BJRPDIX8z1ulhBvYDRIvZE4JQbvBX9hC15dsdZfDq+vxliYxUmSvVKEQVuoaZ6FdDUlicCMcmuCM
mDBKoWZcGK4Hf9OFPUgiGhXwZ8zvlvx/Xp6PuQG2v7HO8BtMwdzLE2OaUFyfFzFx4fuWooLE/TLx
Ji6izhdN1JD6ivyisfO8dDW8xK80JwzxauBZzHgAqwi86i4Z1lJaew+KKIIob7YY+bY+adTwcHhk
L/b63gz2WNckwQArt+6YU75p9DZyFVPUOptHB2StejHE2uEYfZq/oWByXKrWVgiwClhiWsXbVo2O
3d2z2t1ebZSqXUJhxLDWKUc/dNJTqKbgKMI706ixojdlWWS/F78So8hQfVAJmtHu5KpdsTAneqWm
IxHvHeKNzYZK72V+yAHCHLUgvalGEqiNu/D1gRvmMprsBoIBcCCussosoufTsZaFcEQQToHegRXT
c6l3Hn5qJMpbfvmGbjQwA7x0/v5aIHYJ5dKLh+bXcQZRPWtOZIZ50FS44JGE0mnnVGtCs4d2HlK0
o+9Pib0jBA5oEokgpgz2e5vBzS6476pC2q1Lb1gAUVbRqei1hhIO6iVhStxBBZ9FFfqvbBo92btP
0TBgA7/phE52QuzDF0EwJoiYz3XJ7/XJATeGu8MCRU6/4n0m0swnXVDeUbdOvskhQlEqywYGbwon
0/7tWc+XOCw37gXH/vEy8hrr6L57HKGQ9izSqGIQQj4X4XlhP9Mg4tNbqDDmfGUMZQljGjZU+uuX
fzV2WCrDrfPHQhdARsl/ucWYMAZZOBGtkktlIlEs/3NwGN1bMQL6tqBqnCP+z2iUDR0d+2uiGLve
riwoRA7lkTeQs7CA5vsIsDxBGtpBi437scAebffC/x2VMbHbsWwAOZArCHqN0R+9B2MHsMNLknFE
AWqf203/czWwb3ZjBVkvAwe/nmfzUabf1YHlaOFcd8csjDanf1EOQ2rH7MZOnHjbkhdHt3ZTA09r
M2bTSzGscXESHH5cI0Wbv11jaby1GiuJlNPca/gAArLlwAfZl3tII4Up1+9fF3WDNLOEGfL8BydG
4XpzhPNaBCznUGXngOkSkBfJmGwLZncDRLVh4StAtL3vR1qJ6apm8TpX5hsm+JoeAfXpaHoGeEoB
PlsK6R1+Dbf0tY5yRVd3Or+sxXqLgf1zgubQ0IKfWuF4INIRB/ehRV4F9MpNNMDpz52baXRZKlPI
o5Bmcf/PoflIay4+FCOO98E+vm7+jf7SJ8DjnLYi3sznAwB15MsmWBDapcrgR89bFq2aitecOMmw
ACGx+RIPO2dqA4FfNZ6Sil66MnF0fZlj1wTCD/AvDMUMJNo49QCDxnqnSuv+UzZEbVXvN5omBEP2
/rT4qhhtupOy2MGjCUXbTo78Odzjszhfk+tn44bYaSayjhx/3F+BtDtyn/EhftceOqT18tqoePvN
efUkphCdmE93wL3vPnHxrxlx5slWA+xoMICKUI+x7IhBplB/XfFoIamapTOiPOYaQDgG5bzmTIMl
wpSjJoH/MSzeU5VXYARYqcRJ90LZ4SjqxV0FeSwVxC54M1E5ui18G/RkAuuMY8H0XdEuSklQY1HM
GiZb7lNNVYC9HRB91OmQgR/1Soh5xkUW+ajpdvniUYfhw/vmS/FqiuqdJV0G4zvqlsBrC7bXeA7k
AuCSeLqWuzx5rCzvaRJmOcfq4NsLC6AZJzp52AfHMfl4nLo8qPUfIGnXlQUqvp6i6vOAEsiVC+i1
WfILQFuBY1urJOfdl27XGiepxb8zmgE6OV2tQFD4ydQKKR3FjNVAtiSnKKssHWu5f85tWQfVgRkI
LhiOpIqTWdZyh4Ken23r27ergKyO41hFaxGbnk8ZiAtjqmLm4vA4jxGNqARf3YilpHrsGpItvP5W
R46YU+gyTZUDiMg2D9JloWZFd8RLrtzLTAWLRweXqHV0srW0BVP1/WyQNvv2/u62LWePZ27ARiC2
GqfE2C8FPSvLn5MApzQuaQ257ykJclHPMECKU4J4EvYRhhPNoE6ilTbnHG+M4f8diykFkGrSz04n
HyDZcKeAevLiSvjvqKok790YgP9sY6E+t/hBCocPjPLODLEOrQBAPYzgf1qrzmDO9oOZFfr82IGg
8mWpjwmz54kmfVKPdg1Nfba7nieGbg700MvDYK+PuGi9FDiamDPCF/E7Nn92nnkzda123nMsu9Xi
KltN0Eyt4RxS9wgos7gha8DfjQ0frJTGsjl1Y8hsY8D5sjD54cfM/jfEaLM5rvLIgFI4KiczrDst
VqhN3xcNZUCcbiLsgYe+3i8Gz7JeuvV2rk1wv5zSva8PzEmnzL8Sj6TKdhMCAOF2RZNDQu1STEUU
jW9pQwpBaJlKLruL5P6A2xtThC0dYcnh/iYzaQuxrVIxbS3szCZ5SP77bsSoRKsyGxMRSh8wVDib
aCoAsxEaLBIu6u08KLdd/Z3aFoT/Wdmiap2tZOgZR5R6lp2/FvxzIT+Ko2Rje1Gw2FKl74z8kqrk
QhPDPDW2ftDXg2VBW09/Hk4C5XhG9aHRv6aAMxZrIo/wCuzjUy3zQ6gyl63/rky+mY7LUZXjGMhw
ViIw//3a83oF8qdkkhzhkkHNdv+QqyZtdGdk2VGkOOvwjlPJ0mAzM8ojY0RSvvoIPVCOSt0iwjfd
adMiIaFueM2CtNLJUJ5duPwLJHH0+FH1fwNjTK33TCykxKd3Yq27ZJS3j7AIIUkbYu1UCEGDC6vT
oUpVOeV+Ej4tBYnKs/ujXPNh3EETTgl0+xtBfNIMQKvnpPdaU83vpjAEdTw8a1Dwoe50ubCQtSQ7
nEaWv7Lm5Wth10nkU1JRuC/L7DOpmA+bV4doDJM/N0uxwauocL4nVGKiXpQfmaXmttp5yBycJooH
c7zSebAbBP+5T0VY1jLX+GvCR4P1VdcGkxga/grasDXDFXgucNgLkNcJaciMWzOThl1x7JrK82Ph
DFxaebcseEvtY5kt0VCHbI5HElyWOYIA/chXBhDdhBLNhi9cT3AuZjFSNm6beL9Bm6qcSOlhLyGY
okHaAOetNL3jLvzmOTqkoO3WcSN1XVZIJD3FwoQkc8PGIGMYFvbDiiHPqpo/SzrKIPMF1w0H3KFj
i06s3rgZX/MrnmzLsXHpKPhMejOzmmyoWhlFIvdiL5hd4JPB1iPCcU8jHNU7wVVg+Sh3Ga67QxwI
QhXX+XWuUdc0T+vvY0oVbPPGxovoIzBAj8mm96XBpXEYvO1Xg6oST73VtLULVes1thMp3w7MBPfB
jrD09Nu6q3c2YUY9dUaFqXaFpC/PcicxMTAPYC3G57XEZ35VjRttZcwQu27+UFyWNns7Eyalg8xb
gs51gITpolgbDI0yqSVc02t6YxiXCLCFlO14RyrQ70kef3FZRxaWdqhI1uZxvE7xee+FrSB+dSah
Z2BCX3e1wJ1dh+dFUXI66/35OebZd9mquyM3WnbZpXsliiLyGPBDIton7L/v/AP2Tpn8nS+85ORb
FFXhUAHC2S0DGLN4bRPiIQszUjlS7w5MMriDQwRdZQdRupI7eWHotV5hOcKZfHiytnMhWZ1ec0Ku
2IhaEulmJrvI6EOJelfldAvXk1A60N7NAP8eJgZH0ddU5kUG0Y3aVB6PCffTmS54h41CjLOqYJ7i
5v4PmkhNHcgREtRM014Mdhs4z11int0cgVbNOeqzzPXXfMHR/f+ldM5fxIfbyaAM7zMBC0DQYd7E
h2eUpYrNr/M2TEEXNKSs5SE0oYsMkDSKCuy3v429b8YhMSkbbyeJY7Y8m9w6pBbBKf44REsw/r2z
w9OXgcwSN2lWOnaxz3jDLaoK4Ko7nPOm5LtbnTHEKhB8SruEliHgFubm4RLKTLST8pt4g/Qw15pi
oYOvpZgZ4QPXP+AGZrDRGDWTCbzDD8OPAXMpl3ZJ4QBKqxfb3reoSTN79DEUseFQgq/nnF86gJtZ
GqRiEUViuohiX/xuxwiBucnoRo6vFuMyKbG/GvMKNsRfEL0pproP+FOG8YYetEEvEjnI7CG2XA+N
ugcEMNhacSRaiQDicZ1b3gohw+YlaMpSsAYtTzD9FhVZr1vx63Kd2x38mN/ZutiP4Cd7rHi72E1t
0cokxjJhPl4vAYX38DObc7AW7m7kd4SbRVFWatv2mL4aafGM3yObMVwChrsAoY68Enf1DSv4ZgtF
gpXw2lETu+ZKbDod68NoIJ2mbyaVTSxaLbGc7LDHCwwZKcYvmiTCSNNIqlbxS3OCTV2bnC+iQHlx
f0piTUAdjNHOi4dTIGjR8w6oVVgwkHJjbjTfBJbWEB+PYiXF5skB/4azuwsHQs6g2sO6o3fh9ZGX
SYIcs2FakdiHNFpBXBH9+yhUAexorhKlm60Nq2x4hfmhHliiy8KhmW0qRxtXCDAlm1OYKa6yOkyJ
yesZgqWpf/VGl3gHjT++0qoOHdskdjyKH8guRu9cWFKZsfH1rLU1iqJz7tZn6SzrUmZRRR+yXyMh
1XgNf+YZX2lMDQWXDO3Qon8NVedD/CLQe/Q/ylTBNAbWO40sKEATgj5er4lqoWZ1t98UOmV7qVCJ
aYefw+9TEsKzQr6yYANsc+pUrWxkzW5gMQSDmJOMb2Kjdg2hneABRoJirkyvJwXndzDDDWbCxOEg
hF01JUvDGaiOv1TfnHLihTSnmF4njuSED5NGac2PmChEUJtRuGpfJtEWorptyAaQ8s6vUBzZDy5B
uYQtl/UjSd6IjbRcOU1c4T3GpexsObNbWeDYfEJzvALi3W/eL/hEcD2BdOOYr4Ga8euNw63BnI1L
owadBd+9FtDOBBkAq4WEm5D4anVNPVrpc0vcmPNbT9SX70hdxgy3KWF8aaC0mP/rKun21lkLZsdv
J3TEE2PARUEMn+RA8V/W2nBd3awjCC0+9PWHdFwSJkHrp5KnwvGVqzhJitC2jx1ZUmgbsWdMTXgx
m46QkXMLkIcsVqYQ3V/Ncz7riZAmb4c0rNq77YzY6cKATaV1NIBdRKXdJFVAROv0XsN1f/9DA/II
spxROvZbd5dWXehyCoUNaTmQdJMDy0dCh/2VabVaFqDqREtwXrt6+vOj46ddDSqMfIdDtisuko0t
oWSTbMsu60NjW4MQz7pRqOoJHg2uJwn0dyqSgAiZb5hOrv2+VRka+GUP0Jj1iQjESu0L8eIsLpgM
uocC9mOALpq60KgDpLN7VTOWOrXwt0dQyLIF/W5FXwZCsNF2ZKiS9Miu+JWT3NTuMCb94pTyVO/b
tu5lts6NWm/LL8huSxajra5SUZTHCveeM/WPPkGhwo/Wj7+XYVAd6QUQIY2EbD29Th8D/T731j2z
K71HGMzMF3ebpHPtz0/b3OPWCBiU+a387oFHwQjlaobI+pLmp44a5rI77iY0a8n/7HjoHY7/hmKn
/fu3DaZikhoKWbabn0qYfcqexa4KvjZsMPFYS/qEjI5t4EZ1+hLXZd8o4dWTKatRM+bR5JqlEij2
oybykxVa1ddqoIFb6kIBgx3RoePcwDH7IoD3IwQ9zs1VPWD/7vtvAjYf5rfJMbKrPar9DZksLO11
YixtboYLlaAWwhLpYJhukvNWr2b8j4naS64wW8MQIb0PDVYT2oJ4h2ItR9LEspnKsGCTSZX9fh6+
WAalfc0PmbbZ/AOASs6gZyGRRtio4wSUHFZrsgf59nVWyiEarGdH7F+SIlhchP//rCrq79RaVEGR
XLVC21Ilw4OEOWP2ZMQJBScQnsEvNuMPePG1KT2wVmZUNLPd4pU1DKvkJmwNB4zk79g+cK1VtJpL
7vZgzzYlj5NPIiS7w+4b7e4OUi8b7V0UGVLGkbgaDIadc7kM9QVp7uuW8WAuc7HXvbV8bUTMZyD8
9wyq6b+giiS5u9fpTwBqrqmp/RREH21p/JwiUi1PeId9Uc8uWsN3bSkJONP8RzCewIX0v6rvZEuX
N+wo90PLbi/m1YsrhgfWjjtLyISxHS4LKnAuHQq6eF9xWiT742s95nalzzEG9v04OFBlOuwZKChv
Qm0mUTFRWPESp+766t2MZxmE3MWArRiXQOp11+BwekGTbbQGrwFvcjpaweadGyb7avNmdpuZl03d
ZtSmwckH0cZ5rc68RoIv7BS/cXHX1dIwhf9YCdg7MZNwg+IQzjq2BOcLs6PCiq6e7NGzkMBfjK/+
v72vSF1385i9Esclg3DsTk4sB7ybUYJNu13gL1Tw7mb1b9SLq4JaiKZGs77OfXrKgrv45aXGQN/a
7Ynu7AC4IdDnnChKUDuWZqlR6+3ny/7gtrmmDLW7CII44IYUkjsnKSjY6mk6i7dIm+8RKfxTl3l+
g4SG4rD7UDvfLU9dRHRNhOnAgAoMzltY2+2eYEa3w4BruWFweXUYIIE+wX/eZvWaAN/dNBAy9jmb
pi86LTpzlpb9ywT+TVFmogTTw4sws+okE6yodaHCErqBlDw7t5VsJmrVDgg7zSHA0t/kDJ70tmhH
DxeEekJIwYhzb7O0+cUlZ4bMat9ixOnUZCXpnrVu+jyU2h/nNcq1Tb8uXR2vyn0VdOmJJ194KJ/r
qHI2OmxBujzh+HL0skUwRP0bQjaSFFV9Jfl6Y1wa1t7riu6G+ZN1df1OAaKsqUqf9J5CrfhN22l8
ftVoAKoWeAMtDkpzsE1m/buScjMJcfIKiEDku4FTxXvT0UJOQ+8Iz1crWBG4BaIVgANbzctlIcNK
2Gz2XYKMAOTAkA54cilumz3a3HJ6u7l2FqMXGIG3mj3h1qFT0YkDD7mTy7qbb3auz27fhayINuu0
hoTMGUeYSYGhPVNUZr/pXpfNARBpg97WiO+HqQ4d5EUt+4QtVcu2kPMdCMu+IlFRzaJbxZkiStkW
g3gyHLj3D3TvgCKjDDgz63olFnlt5OFP0xHLH6cXsWWvWD2YseAANzldD10m/3s8fznQ5BZd4Gfs
ur3RykvKmfBZOT1UpChnMmcsIF/9LmuNuIxz4TGPZhZjfhSJEYXmLmmAAscBHAu1e3/5MMzrv/J4
/Yfh5YYS1fjG97DOLsorh+Rvqg3PyM284Tw8cUsPt76hgLqVNsjKTA327L5GivFvRrFvLHfsxY58
sFOi1RSD6VrJyXmBuTFcsrAhgpKBVwOff9TziTmfusY3zQdA89zyqVSXrf9HTIaPNmOvLZR+isg0
1YA+h71hsJsJItc4QBSgw8Oz4fH/F97evoiMLJsDAHhOx7dwZNJP6RGTGMvaFAkr+gODXtWcDpLQ
EQyDe3uf+Qc8YzqfZRukkq+QXRzGPrdeeJDpYWGsFvYVcwxSH2I9+2bnhccOeJ78qkuQ/i5EW0bq
5U6GSY4ta3R7TZ5ZOwqPxQzZ2sImHU0NNa32G8pnRFkoFR05pmX1rjFaDVF6KLkssFWrTtF1ZdvG
iFzzBx0UzuAvgqiNixKmuJfMgWazMb3Va2fFuxP9BsxVk79/RIMuxrdKdbTxB4A+UQaA0Q+HVpd8
97R5WGwFXsG4+Nfz1I4tJFMswG4Y7/TJmz4QPl0YjUuhTS6+d22xe9D5qvNX4R6hU+SK2yx7YZc8
83b7opDUId9pwozD4ozFYneZwG75Lg1NFOlxnLxL66Alpupf2y5N6yN1XfOOduSRzvtS7veD7181
NyDSPpyNRk+kZlXoMdrbbMIOeJ/8eGFMb3RHBR9dbp6wWB8/OmuZtUOvv2DESxJKyPoIfgK/Ke9Y
ZKaXc4esOKx6EK7c2e5/FGYvEOF7Ps5gqOrYdsLsozkZrinFLhTcibrzJE81Ydish/Zr2D1pm/1t
cR8zFYh2IywBq6t1ObXJaM61h+SXgEK/ShBa1F64oBFnbBmgItPopUKCg68lfN9X3DDLgpXywXG/
ojIzRCWpOmubdhkp3AbJ6jpxwTGcr8YHnYYy5kdrFdBVqZP1MixDDM5muIp5C/nFVSCBe3rEKwbt
deZAy08rvAIxmmOtoRvDeefDuAMp18BzUA24SkA7PhwGLx317Luj1xeQ0zFOXCbhDyunMpB8Xq8N
ww7fKvkry1pYo2yi9U76WCuU1AsqmldCjFSYi/sO050htwvUEIar+slpkUW2wfYTX4VQ77wbFaQR
8gkuHPTkE17LC5bcOZuiEHGraSpV/NRnuyIbuyGJpaAO7i7aL1Ob26iC7V1lydZCm51XCXqheueg
NNQmYEA86GgKHNAaralZSgibrHEOPZOsgAPIBM5Vbt5MiIjkmG4e6oMEQzQE/yzeCNl5ProYhe+8
wWsbK8blUwaZWYZFfVki6srjdM3nEMEeZSY3u+VN0VPXC0VclewUGDe7+CfjWSMe33vmedQ4uJvf
NUPwpLyX+CiIpI9gDuVX07+9KJ+XsYuEtHzFHNchc6lFIEQ+s4cdtpADrs8F0RfbAc9tXvMxL50U
bQJk1DxZjxxnESWg70LYh2yy2dNbo1fcA6Kw77p/9lpcsA5N8Na0O8teVQIvpYkdvZz/n5BJW3g9
T39gd4s6AFxe/dDxx6TzWCNM9jCUdsrMnEg7cvSikvKtmR/ozuB4+8FoaQRfG19t7fTN33J4gHzx
4JTk40k6O8n6BdCP2hcamVofjihw0AZm23TdqTmplOPmL+zA1IP694qsKmw1qGDMqW/PTP4Pn1sL
YRBjFQ1FtHET81IYvyq9gTVNQU2ca/S1KTG5HbJGyfXiImS0G2v9F96jWwdHh/K8JdGq8hJD9hoE
eamWjsbxd/GgiFI0yVY3aLi3Q27WhIl2TyFGV9puVVUq8v66ec4d+9+CcHS7vo7IQ/Da8FSkkeQX
ehgdcB6p2Tvykw5uJ7Hum6bXFVYNBRmQCA/dwXZ1ffSIilVrBz5RJ542hqQhWQE9Rz6QXjQWHFAk
o1iunQA8og0Ftuh425QuKnDSnQUcmH6m45x+XLKMAgbOo5WfE4SphLC2/I8dA2fQzAa9F27oTNcU
UZtutRYFZlXHIXIFiwvFeW/RpjNObQT+A6F2v3EnHJ/n94JROBTwAbcB6VUI/3KXCSgSmGZh1Im6
J+Rdusk60FHt7J0VDm89+6F6o/ZM25ppcHs0bgPr/WhqfkiQ/qZ2rOLnrP3i9qTRJU8z4UAjc+BS
hzPtLv3IeVJqundN2eZVv8CjwuR8NY6PXwXlTuYh3gqzfwKTQO/Cc1oICd1JJzTBE+KC/KMbNtfF
8ddgrisAnS+NUsilFf+U8GxGWpLSTLHgfOUOK162ffDX+bKihnrVxMt9tOtThGZJMC01Pqv2owD/
IpuTc+Mp9/kt6ulEJqHcHmdrvmlcFlKatsayF+Nwx5N3zvIpj4i5g695gp5R5qR/nhgStEr3ivlC
Ec+vja2MPaNxDMO+NPAsJuzuGsZk4pfWizeIssdQ8BQ2vGAzuJPOc5aUGmyKsUQzpTKh7eswHOfa
u3yJ4c1Pe4ct1h0x/n01v7B5uL3uXGavxnz/iZZbd/C/StrUmcvThCK2i4pcXBvEOvDJmjdzNUO0
z47FG9gHBm4h+7z3Kqxb/qm3Ihik7r1tq06swJc7rj5QDOhNSsvBEL6H08oBgyhXOVfL3PsFn1J8
fwF7WuHc2CD528fK3soU8MxCmrIR1tzefo9S54dRoZM4wZROdnYmFaPY77Qug+DYePjpS9PG9eLT
mSOCrufjy1ZN8DXajI/Np04fSGppuwOeaH1vdIwgQWgJkdTZt0/8EgPwW1q/L9zkXRMr58GL5oD1
TxDrm0taKoDr63bamw90rrsm/VIuyQJ0CdXBBeI+J8KtYwEhWbamnhfgBLml8F9MQgl/+BwKMFPU
Mn3Yd9CFrb5yAjC4aoXVstdN8gvmQWeImGUhlmOU1Z4WiPp84ZqejqyDfnc/4RJoba/Ho/Jsi7Tm
iz2dgQHDSf13CT+CnpzJJ5YVVEkOs2PyfmQqQZcfyX5WzhNzJGTd5vxdEO+oYhHNU3ZseK0MiW15
hiR8YZGJTh1L9ZclHGUM/cq81jauhBYEnrSoTDFLTQsSB6mO4aKZWD8BmVxuO5g+Q0PIfAzWAxyN
2u8vXKMSNPbGXTSBDkrAkMsHN5HlLxLbJvL8bDun78qA0Cahb0j0SnJo/ZnpZotZrCM0nI1tMO9l
P+sPvBkmAbeSDPh2+mAt9TKAq0I3NtQfwgF225blMj32ZvkMf2J5Y/PSgauHDabMWm28Y/0AzhjQ
W0sCxIuwvlboo/vZxp9cEZm5xDBu0jrDaaUQO2MfGCTzCwKTBap4PBtGyXruo/e2jn9Lsj9Yggzd
H0bUyfv5o7cAFub/tQS7VEidjkbwNlQ3PYpFsJHgsi/hmEDHhywGiiYTE0JG4JpxdjB9x9RJrCS3
Tn2a3bPs0ZkG9+6f8IU4qjO5qUiNqPfrQQVWGsDGrvmUiS/LYfxBApkTc4ORZKw1GbKnbN/N4y+f
sqb0jbrl+VBxh8K+4tKGbaB6lGzfIy8jBsoxhvcOP3txKlVTd/8G7xJQNxw77Gn7bbcGckiwu4KD
HGDblnvNdosOBIgeoSfS6hqTb3HIYMbMJ4Jw/lIXms/+Gwdh3OThae8Fy9x020JhHEVanYcsCv6r
/mzk6vyUGqg+Tbjd8ZD8Se70YiNNWox5ype1SkZMeYVqh1waAKudRlLX7cs2kPC/kW85FGWTPDvq
y0a9rI/1DC/of42niJ4EQI8Rm2DgYhKUHQeTOn21YYGkPCrQ5lHH0NT8TvkNnX0kWeFXingmbxwk
kqaJWpcyBjjehF+m5FZG6hNyYt99HQusc2zTMfLA1auFfTDw7QjIk7qNbc5lNOdraymDc7RSFmpl
SNCaSm2IW/FLHe1qLb3DsF8n+GDDvbeHX9f6hPs7BXEih/vjhq5WGnUlb0K+GL08ZtdZIygBg/WA
LGqfBSjaAuPmqL1DrBvuxVtfV1g2b6xYUJX1MF6Y47dWQCxQtxbMic0lOn4+cCK3MipVrD+tS9Bd
e6E9vsIRmZ3sGv90YZjH977hAz12T3ZgInJ0Ian4O2essn6Dugjbn0qo/LEDKwUTmmmRSHk8XO4K
ghcNaHtR1XB1+HefHcSYDZksDkjyclx79N5EybYaqjVZwU9JptBnAnngYLXUglmwufZd7lrWy8cH
vf8CzdEANPLYJpKD9VZtTcWdAGsFO2hgYZHNZbJBYi5vv/NursHjHtAWFyuMG9huTw4mi1tV6mP2
JKM7TsuF6JlUlhrqh1mbMgX3jGUEpUxxejCV/9Tv8xoBrHJVkdcPqKzu/GBr45aAVbjH4tA6KVm7
dBHjMDGncroWEctxQXZCRI0V0rCdkuyyt0PZOPEjlh+2TlBGSa984JEPfXCQwxF+SnwQ3sOL10wo
COFe4nZiZM3Paw3gCKZ+IGbo50kBTRMClwRm9Gwi1TeHUh2C5ICemy/FB3bEdyQW2kUQo0D0hBJa
lruD40PJEzqKN22ezJ8s+d82Fgnkd3iHBfGtKJFwSkPSxbfMoPFF0qLxC5Ty/5TYKJoOKYdJfZhF
WpeTGgkY56+AN+kddYU2j/RfUFudGcJl9ADt9kUVaYaxixdZ0fP2rCs3+hFdZ2nc6GvgXyt+RLos
f1Eo/gG+taIibzOG5QTrz+uxY0+cHHSfYSYHHnz6V0zfoE6mQTIV+iuQhi9GUybbKHjUlba+ZzV7
MLagd+GCxN2eNFEkaUuDS7+ALu+hKvgWEynwW5+xBmM5RV6BR2Mmi9sHm+8Lb+0mffuDwwzohosF
+bnjOPjxxQCZlIHhwnF6qsacHCm1Dafm01Yf3LKwKzOYR8qhNd9zMXbKki5x2JIwGHlv74GEPqeP
qnfc3gnUosgTuXmUkQeUAEKrr+c3f9J0yxUtncLU/0mPSFYCee+pCglJyEyLCKYYVeUpzbBxXzf7
ZofrWPPcWHK0wymvHfqIaoHbERujvAWCjNIlXvxa19i3DIZ8HfyWh4Nl1wOXU/mWOCPMxBfiNzZE
pCuXYXbDliwLvRb8lHYqsNnrB/yUd9zXUUhz5QZbpy9qCO48Kmc5/K2Owyb0K/Dnv17UU5mvrrSk
PWskd2nZw6ZdsEbTuLYsvK5wmWrBG7khrMaXfGY2hRaZFA8JC9uVn0ZwhZVY5OQXl0KB//TRw6IE
TU6li3cSkDN+yV+9rOqXFDYaEbWBpD+Pmy4MTBiIGTPYqjwewq30CyksAoyxLUGo+Jievlhoa7KQ
tVh9OmeuSOIQGUQTpSv9dF1o46K5LfWxYkbM8a4zQg6TpEdXqOs8+rXld1P1OjVdmn2O4c+YRfeX
9GfDE01GZYSJKxOOAyO2aAVPVbLm8L/keZdMwtoqarPksVnlB24proPKIoCCD8Aajz4n4K1t2J/C
k2tUlA5h2wSTP4FvbMhS0129q0pc2HMjH4Wt1MuEjSJl0ZmiLS3sSd1yCPAOLWpUgIrowd0Vd6iB
5+tbSMwIwbPoVRk+b9OJJB/RlBuoTNWupSRkcS7BhZviR5a9SOMTE8UH9BEQzujf/05kW49LoUjV
79ufISh9T/UJzrNRz2KGAjEyU8JsUFAiiDSk37CLT7ZeSygIGLMOO8RqY5/CgNzcgZbHpYfy9C7q
imgBwC74RCNTbKpEOEJjlR21tQfG7U7HFzfEGv3d6VUwiLQN6bKnkEwfnGUmJ0fAVIe6iaeDeXep
4HYGNjPCNtB/8yu3HhYwRoH3fJF1eu/mptcWApt4FBi/SRdTKP8FhfohamWjKQBnffFNyAR6fpjT
71Xdckfr+zvqDXACtGFX1dx0vKQ6hNf021wUosVey1T4XIlRR1MYOdnMEYVd7hUvprH1A/arDPPY
fsRfcpVJCiUUn6aGd36/rDtJ0dWQBWjYBE5r/gGyLLLbiY/kRg+XGdscWa4IpwVW9I0IRCdssdr/
0yKotGzVGCO7wgJKqleBZD+/hkDP5KhSR/n/nTdiA/dpJtr08IJfnUkezu/SXGhowTYSXmzDh51+
a8SnRWvOKq6YO56zsPdgJdHx+PCu418V4t1jOa5xbp0tzIigEuV5D3RuSSX9dVZnoutF9g5wNn5r
jnXSDLh/kJWwe2wL6OUU7rNfzO6fRSrFn1gEGD2AKgQD938k0M0H5gfHHlgj/Xvah5mgAYaUcGHl
Sx8lO3wJxx6Go7wc+/Oeg2h2eJ0VDPf7R1ec79s+gzJ22H56/J3OrlYblHGwficfbcuPavZmuUn2
WJweat7NbeNsqvshN6oKOZQoVrA1fjxIr6FMUcr0fZ1bDUCf3vikMAGSQPmXjAy5xUouI62h9AgI
E5rSpqdxJF0mEyao1Ng+Ql0jCTX7q5E/Kb7+wphPRftI5eV10+lM2DJD3mzraszlEHxahpDQ1LK6
3jgxRTQsQdpWiYaMkDwTnaVqMZcuVF56hQ95AvtBVZ85AlqDwxeLzaJn1Xr2cN0LUaGRd8Kv/kqh
IipkSmmnzcoC8jLuyzjXnmOyR8NVxF5jdOQnyrckVx9XiylmKqw3R2FW9GT71os1xIsbqwWEvkEF
i6JiFZoxq0MwLjCcbquPH+UoZUefi4Ib6jcAxOVH3QIIrDg+WbkWoN7jx0j4q0SYhpS5ptL5ePKk
02p93KE4JQVaXXMeYCSB4ff+CN5Iay52Y+XDVCpSj8vNZdzluIeYzoj73pK/FptrYc9whZw59g1e
NUCH8sRvYUWws/bHjFN3E9Azs0grx4UGwMPeCPb42raCJ+UtL2tD4nSZcyk3vmbjbDXaDlX+ZUI8
XvEAPJFlBadbnHlIUC2SpdsaCOt8Mtknj+5tP4dhxR7FToL+IfHNyn2Jn6ZYnHATGao30zqLLzAv
n7TA4bUoDi414ZBFDqnycQk+/NHVRtpKNeuHLCzKvRp4dyQCrpGtfHE9OWibEpUYUmmOPAb8bSn1
gmPWvWofI4iiGPmhG18QpaLwUHXrb566voud0WEZO4eTnkc611lWCxsL+Nd1tQngL8yMRESrTk0/
bmA+ukZLIipfE/Rk3QQvlw/Px56nVDHsSatBUuSKjf8eSg7a+hwKTzG19B0hO+HEY1EWdaPatyeE
x8w1WXJ5skf3JYxinNakepPvRr1PMjpQds8l05STI3C5nbgq91mSkGUFiuiOCYQnYAD3Ea7uFVN7
KktFRwBlLMYAO8d/J6rqyus1sk4DR+TbQtaV7ghJySddDSVkEWWit/GJYJ2qnfBj4Xb8zAgtR/OV
HWjr45E7ECQ/9RS8hifjcwQGvWQUxFL/qBmbcZAeFFHOE3mh2cPJp+3ux09hdh22DOJ1QaZY6IXg
skZ6plIov1GHVT4LvRd1yJG+s6kCY2DfupXCPbYbRuRsMLHWfbGMZNWwUS2zKB7M5UA32dKqc/sE
fDIK+0e82By7qaTE7lo7NNRAzxQ8W4i3jAHv6uhMCSfPd7JDBsUjn69vf9qj1IxBJFlb7JJfNsWE
gLCd3CZnoVx3h0HyFKd+pgeOwJpcF4xiwnLBBfa+LVg5ZV0yAcrXxJrhEwNKSL5f7X26qU+ScYG9
5kN/FTbiZ+xers2zDOzlPofoi1Zf+K5qLagp1JsGZf/H4gXO2iuUxtFmaqgAR+s/1ZC9wMLPfAo5
3Li9ObEsEoCOL+Up5eEZVWCUhOb/7qtKWOVpgm0TV9dVbIw6NFp8hfVPiDlRIC+OGSY0Av7Q36C3
7lWs2SGLkZoXto3RyH5sb9fd0WjSJp/eTZBnQuyAyndNEYI4BEFVs+TxVE6ZqtDI5bn0r4sVY8Qk
N9vvtlGVGiv1Ld3Kkg0QVEd2giY2b9QzdoYlHQ0ooIKdTITM+ttvLXNYSlGfNVBX/FAkfgW0jvY7
QNa1uVUEIRqkthr8z6ShKPs9ywH9YNkRcVf/NG5mfitFUSwfnH/U/HE7JO0Y5tQDgGGgKr+U7VOU
g7huK4zb7KgyAdzPHTWC9uE4dzxJyz320E642pKm8o1kofhsR04s8ghyYUrFy10BK09Muwti2apx
seTPFSUV7Zn5/Lb9Gzhck1pSN/GSubGsciKhfJtLjaMTJaph3Wn+/mT6zdE1ExvIcEc8bxSfuFBd
AbusO0ODtHBsabKMNYB9YYoYCe+R6RNydiB6QFSbSnytFYl7NPEPavaKtdnL6JZbyiADInJzqCyA
iXY1Ee728zNd0BQP8ZgGbc8ZYNouZePWEq/xgOdoABU1YEZpQTwTdvuJ49a9M8yLdP3ENlRjSoMl
m/QIcfFukBvwy1Ba1r0IrxVmsbid1rE2LE2Zx4JiiYwQBjGK9sC7YVpZgUnrMpRukRavlmKIt1BI
HN1DZ7A9Iz/yFBE6R4YSlyVaWdKKttPv3v/LGEfHJlerp/Y5anjyPkvW5iPYSw4gFudLsGdmPmK3
ibAboNwWPKeX8a/43qwk0vx4Z5DEDBB1ZBOdOCRp9hW5JzoNi1AWzh+009oukkM1hiRyL/yhruRt
YLYb90qTBb8cYxvfCCzy0Ek3HMKQudcJap0TWDm8dlygnBiM67jGI7cOrXSMaSky7ZUzsnOaDWzm
5IWeB2NfhcXCMFeU2wGFQ2+kLesQyyVmQCktq2taiVvOVWWbHEB/8QQeiZpmbmz2o9DezPMig9/i
W7qGiAOGzz6fRg9N0AgaOCn1/T23wIxBQUCsM8zGfGaKvy5qgJv9l4brD6dyKl4sfw0LpLDNm+lM
5yRy6Cb50+4ZrSas4qVhLdDUe3t77xEn1piaB+24K+T5oO8WHUtSb8Q89mT6BIiCcSHMq0CtebpE
hh2m0BoBjuhrRrNYjfmha8na/FQBw367h5r1vtiX0Jk6TxNfWe+ruG/jBBUBxrJdmRyHi1WlE7ur
ZI4vS8avsoXDXUCIV2rL6bQTv92PMnyTqKjz1hWUzGAn9uiwAozemgpEL3g+hBcELeQX4uea0b7M
9qBCARDoRiP6i2ysEZQR/VBWCpYwdMPahi8xwDN6xwydRdI3maekxLtdfqBq+ETFQ43QA/lRyUUt
yehQ0VwrFlMTSyIx/9M0ZZxF0kQYLdbImET5wd2NcMbNQOLGfUTy9azgj8f6pUcXU9BrN8GULOEq
rVdSQEYZdPqvb2HjsmwtD52wSvt4nmYb3Yd0umSf/76o+mPozf0ewGqcXewg7Et+W8XELEpHzGY0
E1tLkSlsTTAeMkPI5VF2tzCVVgiW+OESzSjYexVLSIb5FgWIsObGuDUjJR/sTYt+s5ZlzGRqxNL/
LVOP+pLHv6C/oShNHhpL7PIowL5RL8L1OAnsfdFdHKtwkMmPfKjYNpYIgP3O2CBkc7VnM7e2n8qG
udjzPS1++jEjWZtilT8n6wZFQES3eoj/KH4P6TAndUz/2XXG7c171MiINa0bl/UE+8UYPHQG5hFI
a9DHmzDH/sJiiDHZNWy6n5wYy5V7jRCeEoRnRxAkLuJ3hgokMzHWmKrBCDYXdOXB+JmX7Bgo1nea
cYvLvE3HSBbzp1uqM/PckKk0Llepc8SdhAL0VTY+aZsUIWlmoq1G7xQkQK1wAvjubFOA28utF2RR
5e/ZwzQWMLv9sxg68vdEP9ZyaNSwcoiUd9+xxvVpvabGTafTCXHslcUOJuotbhYOWwet2uu7kMgs
0XUgKEYoBidl+03ajaPBkEhl/03FhJ5m6+/KfNEGKjtm1G2Kl8AGBXByfTJipbVDYxRQKNlpKmSG
B1QgW0STv+h6Z+qPEjOPQQ7MXBdqo88RzsdTzNYwXRltBwNSfwHjhM9FaEw7BgomRQ4OFVlyrOEG
bx0BU5+zoKg+GOBvjcmo8g9nnF9ffT4P+mHPZIUATE3qO7VwaQn076rjM6GDo1+mSb2GurYT6nGk
DM1b3Vb3YkiRArUzyuz4/kt7VX+hlHMYARSIT52q6chOVyhWl16JAZQmo9qodWQ4OTboOvjVvCH/
/gLQO79WJl/IT3Ukr+yEY6k+0durpKnRy8VVziH/zSbGNfnUm388svUrOj6uCWGSW6f6tztOa4AN
YM9L66FYe6tBqWs0LdQuMJ26zWzG/uspawpB4S+QPVgZNhXHk5JsgLo9eUn4sTUmdLbvlvd6KD6w
Hq3TpfxDTMXSjCIYXDKcKGWKkyvVzIhONzNQ+gteMAd9Nsghu7qhx9RPTAa+Ds/GdQT9GAOLoA4P
uCWHKOY8BXa+aE79p4XLTJ5pFkcGWAxJn5H67cNhWmfNi1gMfJxVRbmYdoC8GkWaHtS3m7JW2vGt
4s9eYg3Z//1S92+qJfFWXkzfY/hJxF6YYkw3TRwNQiPE4lGNKwLPf2E4AThnLpCzuoH+3SrfNy51
36W+ZOgEgEPlcZ39CTtSzSHwtIFZHu5SbI/DZyA6DFL2n1rj+LCjBpAtJBTTqB7XQKGmq175FSUP
Bp73JvT7lujQrAT4stveyP8QqlXYI518frSTnGwzAMfrt2hZXsa8Eftkj2+49y5ypEL4ZmdgFy9k
Hn0t6FW0EXeGuoJ/DmMj1Rc685t83iVWnAseMqSQ/xVcVogAeE99yCs7HT+NecETnsMBDP3+rs5M
yly39oTN8j9txH3naeO5XURu9CvJwQC2crufzK+ZE6+phQulAfHlUIAMadXwhpmAsxN1Ckhoutiy
kMpKfLBg0jxXw0CTpDqotWyxteMk3cG2exI/U+FYrnypW+Qkfy7MrK3OopcyyA0tShUzW25jblzn
rdCR0B5V4ecynp7F9TAK93XbSqahpXlTmv3SsDg5b3ZvYEQkdlnaKvUd0/Ps2NuQ3ebCtLla2w0B
1NxdX6fN4JarBYHppuMOya/ilxvpdxECF2547KgeHmePuetzztNUH4BygycSA4wUGgF9l7AQUbVV
puuUZuxDGbaDVBfAySeKgkLZGUzIWqDOP1Yqy8D65IZzmahBuzbrh9D2QN9mFVMoZaGCNWEvqSKj
9g+oj/TKrSZr/71pudUtBPRygyWD/2ITSs8Kvyvkbnh/CaR4DxsIcGWO5YXcTeQLUkW61RXwh3QY
DzJyynTCKekEZWHb5PzCUXrBDtsPg+ru9nwvRiSeiDmbaJt570CoCG1uwif1JEQERonB7GjLQFxD
i3j6Z32XpEiSShFFGM82OuvI7jq3i8rdTWQnt/6x9IxBXn1NQGGrkK5rbmt6+XV+Javm3Hh3yXxC
L2bT75s0VLGersyZmT087/zKfe+/KxZIjTIO2N1k6LJPSfxEoZrotQyiZB6XWDXiE0O5scoMziV8
1bym74mnfLxZfAfx9LeumwkHEL/Jw4Z+WImOe0WIXcNgS2B9AoyknOQu5vJG2O3JscLK9qQYB2KM
6rhTOxUmj0MyQ2dZhS/Uz5AJtZBbRU8mkI2LWLmu0IKFjBeE+nPMfEJbQ+mR8svi2WVwiGB4ttX2
qipJeZpIqmewcnajk64LySJs6yL/GPb13XcH8D2DsaUH6uhgT9opvhC4YrCKeOHqtbndZ7AHaxGK
0+xF1iLPIXAFd3VnKKRktfXeLM8XgvrqLSXxGXYGY+Q2aH5VxsO4yo1mJQfmM+8CUo7NEtIz//GC
EbewnInGOqy3fcqSC1/qVOPvNXdKi0csLsQdit5xOIEPMacehUqo3LJTZYnaI+LQI3mZ4AuSdGpS
D/fa4anbpgzAgzsvLz4RHQ/b01L+XZTmalyjXOeAwDDkeA+eJ5WIHxdmO1f0jCxljIkD+rwXJlvu
jF/nrCO6x/ecpb7cf23kNe+JgWzGz+E4WAxnD1LJsQvbEs3RgmfThitel4vg8ShcmAkPdunwnS1Y
Xc5KFQUBcd4x5YQZ2a+eQ/g78FKGgfHrxjif9GDKbOsgwmiygqKAQ/fnq08/KGMKA1LlsdjsJ0VJ
siSHkHAzsdCXQdu9XisTgOSoX+vYki2/DsI+3Xu4ohboWQxX27DwsdYj26msA9kq/PTk1L0ttYHA
yxWccfXhE4finflK6eozty+LFgsZWDFsO9dy6E7lDsWSGFiQDQcLRG45KLpUBIcuevIlIDuQaecG
CRKKH/qR7khhgAqJ+GrIk785HMp1Hsr/QM+pVhmt0cjIQassLUIXQJVFLW79fy2TEViE2GlXmcq9
/QLIWBuITN5k/DQzAv5WYE+fNPROVwr7FZzVFP27/ZXvX/pw08XSc6X+SWSY90b3mNZT0CBtU/7q
vln2S0/QRF6t9XTnJcZnf0nFxvwKeBQTnYKBUcuOSwrkei0frcTUgbqEnM5cNZS2R3JkX/SIjyWe
sktBUKa9fpWdQZWgY+Cg4WVD+gegPSHgVPRW7j9nUrcX8ebqfe1zh29R7vV9qU96AWL+DmviHJOO
mLpk/3o5NVr55S0/CV+fAtxrjRRMhMBtwxW4qqhlK9qHaL48xcMHWxrEeHT0/psp8hrNnA4XZwsJ
ZSfByFCZPXqiHZJWByiuyz0tCSHxzOWp/LYMJiYH03HUoVSKzG7tleyl6XLhAOXrUe40veLYei9q
+lFTMPwRfl+37m5npSUdsz99EoJD71C7G7yc2lIosHqhkvQJ2Aa3gap+4MW6kpSHjQfHb2jdtVkv
hQRWxxKhwJ25OpgD7ON+QB+hKXjnwgIKx5gl19vHfmzAEkMipSgACIzw+YUlnmwawJ7Wc6mScvtj
cjY3sKq04LmEWPnM47hJEc1oBEJ+hQ+ctsxWJb0eO7hUrIKtHcAuRIDgqxn1zCCH3HlZgfabvkpt
C1B3noONrnDX1v/GdfZp/lcS1TZwtyfjvPPQ0d/I0GT4l4hWz+Grh1t1z3XwwpaYL8Q9fL8i/zA1
pKnfYLZQJPSpKlg3Zza3CCbyJDM/saq4OJj8gX+/7Dr9n63ZQbyp3ZYXEZDZ7LgKRbFSlF+ajDbl
psS9e+TfZNYko5xtWtQf7gJ+WqFR1A3JE+BjPiuIRpoKMBHP8iZwv80ul/oD3wRRt0iGlBzbdffy
h9M6ptoN+M+SF0B4wj4f//nz2+UryJPBDP3+GsTk4PgBVNmlKrxA8z/12D3L27VFrWLIJsApEHfm
Sqkkb6zh5wDINRtRYfssInMfh1Q9DtvaF9sLEuNuNONal4C94QFLN2YRxhCUxx32flrjOfXeC7Ry
aT9DUhmBfxtL7csOgrQgnqvFaVDOtMgSOSFSCeQqPf2gL3CC2DLDMUyXVfvRw0XjqCIcnSTYSc6i
uk1jxsgjm1mEl9ZpGhaapi7iexo7NALQ90KPNxuZDEcrA36nnMqkrrUAsmrVgomgOrGpr4HKbKFq
QbTKXXbw62v+ibxZUkfkWK3u7Euu1s1MwAw4ZMYTFBj6Qmd1ODZn6owKEf1NlV07X4K+4moDFo+k
zroGWLchzLZt51bUZ5xPzE725rU2O2lGed2OlP1FfesfUfZbsyzK4GRKxtOARMOmMAwWgtKJyIuM
khrvl6ePYA47h3LUPYKhLW44SMSC4WtChMfnrroRkD3rgcj6VYuuc9UShyVhzzOOdbN9nWcCeShw
tenJbq/Xw74DrwXUrg6QRSMriU4thFFcb25DcdU0f8goqiGCaxM3/utPZr81jAcJu9AF/evz9WDV
YheBdR8YzfaTGL5uP0szXmq7/8X9n7031p/ih/XP8ysnoTCwKvitSQhl1c69kjmNSr5HlPj9kGnb
ly2Ta5lT7S+bpNilvy35/B2VmJSv/UNetc7Y3g9UAwWo8/7awtyAaiZcWPdmzff0efmyknTKz3TJ
95oArXon87zIwUqSkoVOgOa/th1nJirWmFAvQ/4q7Hd9KGpOeUYjcMskiqYScs9uMBFs751UK0xG
2eqVnXsteetq8Ls3cE8vDEjP9kCSaTV3txH6AtdhblBZcFSluQm2NupXqNz96AkF0ghoLPgFvMxp
+LFYuZ4dJKS9wfxSLt1E2OWZ44Phnybui4wYhnP1tm1ntSb3opfhhCCQB2MPUJC/ylTqaeoSIM2g
/1C0fq3+Yqg1qDP19PUYok9mim7inNAEdOL+3SUlBtz1DvmDUpR0eGK85nPxEUQmtvTLNCaFBgWE
sXxMxYWM/7x3d9GvTaJiFMWBtiOV+BccffZrGS7DQnhI4L/hU2cIzEfgujl33gpS1P+KNbAOWdAg
awRfrT93yIccOQORhXuBavfZ+bU32amHuxGK2BfhN0w+98ICig8P3aaNZq6fmZ2JuL/pMqAySQNX
25xPTCHX2G89c+AY5iEUtiQgJuVIhqprpORpUo34q7jANEdRr2kJgJIP1GZLMkKlxvmSoulYtnXN
VspsHE+/iq6d4zZfCcdDjJeZb74qhlJTFbTblWst0o//nDxhRLIoPcafyXp/TZesUywCcHLxRfGP
1nZvBzpmyVKaIpZQSjW6/mjXY0MusVpqSucflzZqSIVtfBgH2dLfQGB0XXvvqJx13lmDTtYDVgXY
fV3ZZEamtfMBtuR8K34zH/sH4QOKX7Exfe7In7Ru1sx2Rex0WP03kILkVjDFb6QE9kIwMTyPtlKR
1U0WO20DMzHhDCN40GlMIJ6P7QOoFVKS1dci90cJEgOjiBUDs6XiTgRII3v6sGSwDvVvRAitEUjs
Resn2XH68rST6B32guYzppZy/3XUjLoAbj5bMnrAka2HrDIJEllPkzUykKej6nvnOkLNr/Nb/JnX
6YCvqrtPUkyZJiQLXdOXwfwJusD4X/0mlojY1IB9rBWnxqVgTRGhwASRhNlRgho+/KjqJ0djwWLX
D3Jo9Zc+ay7FrX5Xj3EGhurRYQQZ8hF/R67cl5cWTk2kb0B8OAu+F7+PtLjCTIV0QNpmfAnkR6i5
vYZFPqspjQrhSsCzGKgP+YnlbY7tlV0xKdguWyvL3bIYh7wayPcRZl52r3oSvs+UekshTT116751
AtGDGOKUFDYVfhdwvjsYPeTpkJgB6iCAEmdj+NhbQQUUsELxxDGvGALLnWx5gMSgSjZBGHhoGU8K
FcqWOWOdIWlZaJc5GdvX3Tiq+ekTVXvJ0hB6BgGx6ACIdAPWXQfq34tQPxvK6ea2YQa27PaaDhpf
L0xfXRDK/W7ilwHmBLTAAquSGCsttUCqCMtT3Ez9zc4QKFB6im48Yqf28SeotCoGz1dcAvY8I4DF
lGeABs/0upGJ3H58DZLTUgGgF4ZTtABnR/AXzKWKlJm4J/Czc4t11eP1WVEfroDPq8NuR7eRYNDN
mmUj7Ej1RNHFlvyVDWYd6uZZZjS+A66BRfhhyS0TmNdWUk064aVfqvNpYVil0z4vf/7h16fw/HDR
ncRVkVw++EE7KGVIzSmojR5NmijHAtj4Mq0sbJr1QDqOfDea3zp0YQRgOK8nIg1pQyK7XeMJUamv
7C66bNedRLJt4pJc8x1nq/+1wLk/+j25dfOGOQrewVj3OhkjjAifxO1gVrul66uPsNyRDCQ1TB/R
xW/QjBWchR7Hi8lOmriXIiiO71eq8PdVDpbJ2ZCOYZlcg+WsWRy/gczI2Nfk0oRxzlaWYMFZP3yO
9yn4qgEL80n736+iBln3E/XknKrkNXPQdR1jgngJXssdpm1fjyT4WfEST6wfjHLXlT+mScbmHssk
bT9GVv8M64VQhrVDvxlANxv6gJ/hIUsA5dnbO2leRX5hnlYeUhArmqNEGNHLHphFiwuew8PlWIjL
g53zrncFzxDR7vcEPA4rrzWirTr7lgmo8YVjGsU10ZofcycyiZqwOBYXSfsaQV8d0Nqov1hdU6Br
0nhK8B1MCSO6L1bWDHdFBxUwLrT1BvR8lCmgUUKMnNFZcKiUWdR8mea2372jj1nYpsywULJYM2qu
iInxyDyjaV9fENxqzfwiGDU+WU23uEXnosRmNSUZcZh9osAwGi6t0S3z+RHnSxuKukoOgg1MEckS
rMm3oYlm9RFIIsvz5p/1lxS+Z90J4szjdQ7uzk6JiOGDaDhU2cp5ldV+zu/M0D1vNp4YO1G8IxLP
kdMEG/rjNx9/7a90eaFMRmnXCZDacNlBfCA5iIlNTcwW+umBg0ZRzUHUcvrIw9OemhhixH2eliQ0
++HlS3ucq5QwfuebQOmohx2ZgzdJtcc1PsL7jTo2fv9NAt/tG53UR4YIph7Mf0HMObst5CD7xXXL
aFOCtR4kAwl7Rtm9MXb/+m6okQ7qvdJy+ZGwwDifpvwb22/MR0v1/k0+TLrDL03uUpJBUU+dXPI5
p/DQAtfPkFcTYKBbr6ImV59DiuCEsZXyrIB6YwoGPeoxhy2s8eHfCd8e4OPSBDXbCmyOx4ANrZUK
yUc7odVq3+/GzPL8Ve4QSKSsEUgLg4HBu7rTE8XRjf/wrmQ3Oi7g7mQLra5W5gKNQ/TimqmZjyx3
apARSpVe7WzH9+EES3O0+geQAsiOUhf2YrwHQjqccwbSvPzrx+kK4Sr6IxwQMwUjTDT/KH6CN46o
qn0VW0TiZKLqGG7Rj4IC8LvhU0doy1izkmZ+I+6GoXId4qTRIGxZgS9mrSmnd+YkyUxMKdPcf3tL
8z9lmIL3Q+2CqktXJHSl+ODRoDMdsyDO4871PvAitFpjmgEnyMWE2p7+m78GQecP3NVljpQVovqz
/1a25N2A/T/2es53zW0BlpLdEs7S5kglOkE2dfucLwHGOyAT/vxFzv5RY71rqXNHo7+5kfWiq9Wi
EMzVIj8mrGYknDsvo52yPANJhCC/KkqnviPNEYwCfzzYvHkr1WtZPnu5Z3mJpYZ/rap+k5elEzOY
SQy7Vc2dJS81iMVouWmZgtlcpUnJP9DNm0c++JLPmvcduzB11x6r+EXR9oQ8rDVlDSaCvpNBUlAU
r6t/1qjEQcaHLYvLTzWR2cbiO7XfnyzKOV/rt6BmACxczAiaVcozasdA6hR/CYd09XNQJs5HEUmZ
GKOMLFx06586Y0EiA0DpQDA2U8kzOIE0JYtwR5dRRu0BQzB63lm2vP5BdX7cEN25Jbv1EadobVQf
pZWcFpYu5EsdWzbK9/GIgTQve79tWG+KOBpWaRpq3eXOGJFEn6pIbolp/dZ95/b8IcfOcVsz+12j
wfQoKOgj633tMPHorLdJz8FxpLNl9BgOgIsSW39hk2bQFno2e7ahY7Eexdn8oudWpaL5BOY1twNV
vWj1x/A4RiuhD8wsrx17xQxls9CNlKIEkF6xBmcQwlpQitIlHhFVkQgsqFeXkXLwb05IOp9mBHM6
P3QS4YlAxk46fTELcatA0lpsJwB/zr6tRDXBlspuNf0JNtoOE2b5iIYu8+ymq6qexxXFR8ibCPlc
flmP4ZYiRkPy6TdKnkL7Se+F6P3wyEOIiWaxrm6fQeGQoKarBtsec3Z48m4OEPnrC52FwqySl2ce
Vso9mrk/CwhtDdPEfh+1IicQUJoTwgkxo6wVNwfZvzuLXoaHdq+oyiI44tswwVi3S4vhypkXzaUt
lwnDJ4qczlnrwo5wAnr0facSJ+/I3TxVdn0BqoDPFF4gX74IhYSWRR+Xre9GyBpPUv4SBWRxXq+o
xtNWOK6uu/JZ1JGQ7VH4Umkxj95xAIZ9gq7rOlgVamoD5EaDzOcwtB7vIrKT/gC0um6hkxeqnu28
PL4/3FuIdsErsZbiB/Lv4VnOx/1S1G2Fc4E0SjkAJJmwbzqPyzi+JRZW7pjLIQh6mnIqOz44Vadx
zu7m8jSpc1fphW9z9Tu8G/jI28P3ubcCB2Tcy3goZH2YOw2hw7bp/eANoRkA+F/4Y7gR//mB11od
pg92L5K2huqhgHoR1h6N4bVn7i3ZY+KSzoOBaR4x5xYPKW4G9E7gbDwL6TM8+aNmaHPPUhKxJLY6
/oujUMF0JUTw1h8DZBKPHt4YXog7H4p7sxL1trDdFba4X4+rILmDq+pWb5GF/Vi4Y3auGF21jKHL
fKTGVdBD7TV0d7PLzodygTWO5PbMGsVEHG3FyxnbNMcaAXeHKqPUY/oKPj0oGOMrdMKnwhCPFVxV
veYWiPiNVA13Y7ju5ifZe75Ex/rUDj6dk/bq9O2Csxz9b5CbbrSaoVcA+yHZfonV0mFAvU3fStKt
DUViVKkmMvH6zNfb+mETMlsza0x7tNpuCYwwFnJZAhxOt8k79Q2sJiHJEideqqgFnVyChVgu8h8x
cVoPicJhydosL1FJWT1xQCDjrtjOs9hdz0AgAa0xtCEgkq0gWbpkhhjFIfwJfCXDAgoZQuXvT06+
cpacuM02BdTGsawu+h0j5xgZ6KGD39xhV6uBTztDKfogUVK/Bhkmqsc+vmZXsGJPUSWJfOpzaUZs
drUC8tyU2QIgwMFle0fb/lGyZ9G6xaBXh/1SVxn/3yZpL6XXDRVtxyJZweEmqIlBwGEKI+a8AQMT
my0duJgQuAYekL6sZAtosgxA8KUwAx7/a+IOEeRnoT3IaAge57yh1i/+zhKDEs+NoJCX73Z/8XTX
T/jMz7DlWZijHmyJB2BKcSBoCcICyFWXf4gnW7LRSw4Oe8z0xBlyCQ/lizy6bkgzeGazjJChWYAp
CFzWecDsGnGqSIjWO91dOz0np0RrERDR6KgCeoXZDIaCOIPpXHbfGNzkMK+FarUzcl9eSt9dnmE0
GjlguKJuhYBYsU2K/2/g4sZ/ZaABoyuntm6qTRC+BSXZTm2slW7cRu/5vBoQsVC887vztf2ezQZB
lcvIYqvYU9+la4WQ0yufOw1hxbXNYwMecjO621xIfX1GT8V5KHHWAn/QHqEzvceb6KeV7LWD4NO5
98VBcsQ5ML4hrSsWmB0STN84Zwgo5xh8sBBEgeZA+hkyiOiR36QMZTBCgLfAcNckxmzzsjayVN4h
etUcYiEqPqwgp5DbC0PPOtr3TL6Lr8TUFT/NGgDXDuE1zTcyUjbPIxm1axJhuwAT78WUKssIJ+uK
acQwqcCWyk8k9p7Dn2MvJASl3X1jILI5Oq7CTjU5X3gx3j8bKA5rQhuh2Ua3tfH94gVh/AQAVyGf
4ODWUHwPLvZPxDTGxMlwvTS1YdWp7tQe0TMpCITodI/PM4WFWVe2lhqerBZ9tk1NLKKm7zCq2Xx/
vvS+rkkr7NHmJGnF2M2oW/6zdvZL+XedcBfwY1COE8Mf0SmfKUgzVmxdQjXYsSNp6trRYOPFqXXE
mY1F8w1MpF46cy7cQKl7kKUMXBYXXTnv7kepHWJEq8bfHI7rwMcw3+Cpw1JeidCWZplNWc0nQub1
HVzmSMMzQ4Gpt6W8DBokdzflv6mANJyRmbkqR6HodU2ckThdh6dZW2tfn2tojB7HqosUGJOtJprt
dXV2WLmHbs1yKFWNZ8YqgtldNam1a1lp7mPOPds+B64zu8xRY2UK5gxOW4iHtuvXVX3PT6wLQDE2
VK4VvNQSmduVHwIMlv2dIAPqaAoNr0UT2fybr/eAAAN44t7s/bnU9O+J9oEvwUdakRYaCoUQMzr6
qhLr2DmQxRkl2fVm4Js2m6lns7avvv3I5hviBFDwJNtRe2YJCAnoM4m82fDs6ZmgpxAPQ/jprG4f
QlIa5HnCGsTCvSH358aBQRIDBhuZi7Bt6xuo74YpEj1I0lf+ZhtXYHYSaCH3v1tyN64XVlw2p/Mk
m62GMsscD1eFYwMJrUTw6aWQbx18rvRUXGG82M0e05hoCPQfZWcMK2pEjNHWRH+pLMxcvqGOs5ho
rvksbi9PbEF1WbbLEG7gxiWg/AODaKsElAe2jlhx7tNUK/SK48TGwIK51mmeScrtGgG/Y1Eb2GIA
dkGm/KsPKd5D0Nja9PGP4rXn10oH1qB5riNzlARjbX0VTnOa1G/e3HmIWLS2nMLHz9dnW8qJ8Vtd
+OkV3MFEHK4R65Xgl4RqXVN2Hkdais+kfNvy+6MgU2GUI9MaTg+95SmrQJibj4lKwMG/C+ZZxefO
A+dYE62IjsZTU9N+Vk04vmQ7bY8qNN1z+8tXT7d5tj/t9ighmMfkw2zhvajs/EuMnNL48DtJd/PH
57ToFUirINa1Qr39Om0CqEUaG2oQ0/qjPWFhSDkODE9d9ZrJN0EDrtIyw/IPDmP/612zoDPTO4rs
AhO6BmvT1nWZWVNQIP1n37PHFn8HKDOEROcVzM+0x2mL2Ah7+ZerAJE5as5sAl+7v/RLzqdLiuyg
e3av6spLEDkxaI5/+RVbbMJwi7ZlIId/mCmGy/uDq40HVCOpPbsAXIY57PLzI5RMyGose7fyq4eA
M2jZepVpBi5XaqefPOKs9KwtbFTonm77ySgCfXHd9SjXGo1wzVf7h0vpDxF8MaG6jLUu6qfcCCfQ
OKS7uLlSZ9pnQL9Vu61B0n3NRYxpqsvfYYrPPsepd8GQBNCX4G4s0F1y9etHHhehqaHiZ4LMQNSs
0W223Gmdt2DvDDTjEdPVq3MMxqD0xUztLeJdXEsmzVUF9lYznjALhOAQNN+UEFzrpkZIoutlg8F1
XDDzpi+4MyBBCNnGEf3R5Ad70azF+cv0IL12d7T8N3wuGUtjYHN9Bp5xmlvL49CnE//xDZOJwjxI
M3pePBVMX0oRWmO13ZdPMNu2ypjkkHsaMZwjQYt2S6woZKhCWFgIOIK5pg/oNqDbGrYWyuM3Ly3M
ljyNQycft7GyrnBG7G/C3BbueXJHusbVgPlm1S0fASYv/+RVr9YY5hwNpjzEIZPIeIoUUzlQbItj
FIgaCTLFpY+IzwZfROuk4upGSb9AB2LNcBUXyJnSYbdd/qraoQvsW2fUU4Uj0Y/3sTapA06ElIwi
ltY/5DiuG5YOck9Wv/OocQqLOjtzrfIVBAJ7LoGQSdhOGfXH1fXNi9zE0SblHNYsA+we/VCcveov
CsV+XIlvp0pulUPjCAovLzD1W5eVyuCV7IUA5b6Xu7zM7I3bu2L7X5/MfrpXwN+HRiVHSTV13nQh
kA92z6lZqDTXZUsBVMgSirddy+iRfEy872blmPuFbFKsxTqVotgxTfdSXqiKeG8MqsyErbStT5CM
D6zADZvtzKYyRgDFD6RmXnDh1vxx+Dx0/X3zsMTtm7W/o3Ig9YhmLTiKsSJ9oswgmHKh97bpOisI
aCPKuyNqS1B49r9PV0JzXBXucGXe6uWNdTAv81MBcDQkMJpEUwad6eL5GAfwDhJ7qOoU+4BY/x32
PgXuFtpZHniVlhY9xF8pMro8TvkE1WsLQQ7OlQqv9ULlJGXfjIV2q17SPIPcVJmQtLMpDJGTXODJ
W/awUayAZRmMGwlF33zs+NE4lus69kehUCCabTdMFRmJ4goxc/Gcrs+rGH8NwU/TDDnfGw/FGVx1
PhP8ehsc1brcP7IR6lE7CXeRNTUA8Xr8d+nlIBf+HS9k7H/mgxk/9IP8u4gS4O90g9t2jVRGo+ZL
1B65UTtFme+FBd0762A9xN8jTFvzQ+HKQ0stvAcPEEomHKClVIySjfDqHJrjX2sLyeMVVtqDHArN
oYKUoc9gdYhpNzT55jK7brHrXI7pWKpS5LeNnYwk0/vdaicoBEZkwWKjcRxaal9RXXG5Ads4+zFj
tnzg9qX6sGMXIS8kS71ZdqeizQWIt9tnl++EhIK1xeiCPN5ZpperfxusuOSPZsDDkFy+5hvVMB48
xFIpmANUS8tyuIFc7mPKEqvrfEBXoLUZy0DLSiJ3kipqhRXr/U41M1Z7A5X2lhTzldbou0wUmMDL
5vsbI8DUVC8Xxna9HUpfTJLBwBuh10tWWgJOZbN9JWHNA+n3/KiSaq3uQOo/bqzMQjFvilWxNFP4
IGC1a/tLlIgbwCi5AxC2G7jxInBdGFw4cUs9sz1B4aGhcnimg9LsYv8mC/5sf2kpY3+l40vYlPhc
aialjQjTwFu1RB4QvAr6+BdPIkx2coOPT23rHkjwxEL+Q3B8msNYcfaSC/LAsu6piHwmBCndTYEx
X4ppXuOF2YS2VYzN5GB/YB/7r2MkC/mwwqGx1MM9LU9PiTs+3sTDlKxltiO8x468iCR0r8PZDQuq
A56187PO/WXtbOzPrkBH6mMaNbsa2QcutdTW2fV7EjDf/GtbVfON8CahZFIcV+0ojhCJNlZjt85a
yUaHR50x2RrHg4fOa1lapEQUX8rw/V7taq3ZsRnUu92apqRL9ptQpSzmoDg06qHoYRKFEnEKHVZl
+w3oe2LZ3C+AtljWiHwfmGpSagVJ1YPGvFrVbEFgSC5urAJd92oDfqPZiBadPoAloU+5Ob8fQxg5
G/nOf3nLLh1J+LnHIMPapmVJdDcwD12MMym1MoIXFO6AsKp9LHfCCjIekfIqqO91x8dQ8/Tqzc/d
YsyUViEiPbNhw8zeGnzKMhDj1vnzxw0zUVGDYPLZUPZUabJgDpQJgSwfGN9FgTJPqq4CjvkcQwBn
TTBJcCxPwSnb5CI4YwpAoS6YjCkmG0hpfeN1hVOhGNsr9Q9M3+F7HopFSFhkyerVtPFL84y90wUX
D11cD6OPi5gRYf8vQDqLc0YJsEDxFBqXsRnCD5KrMZSWrTUo1d/McYmkK965knspVNhIDqCjqoxf
+YsAFuUSjhereRKDWRvkT3e+SKP/Yv6pWlMN2o4ZeeLfwl4oGdcACHCA5vILWQeKkknp5ClKii5Y
ahG05VIrP5CbBxl4Nk463g8wlULswj/INxNJzkITdhEgnsJDA1oMfBGuUKi3xz9uydWGs1VlCMfR
uzSRnjUyA0pSKSGRypODGcyQVqROm0C7HaFsapMplhI2s8QLZmsWSRJgpyDFX+Oub+4V82AZrRjN
ZCAmhcQ1F91udxViWKWrtJfCciz4Hb6MmMUiAjXxRxovFXTNvjMXKBZnf4V4oVhKAMkP06rQLf6u
g4aE9UI8v92ttHV78TSgcF0tvqY6EPmj3rMtX0dhpOunNH4J/Pc1+QM2mMyUGoc9nhLVlM1Xcw0V
5wcLsH0crkofC0WH3GEBVPN9Ro2lnfe/AZe5lnvqdHaoTNF7i8sfuIWheH9nUZMsqRRt65CzChPE
sqi4RdxIIWNaSnNpi+yko3rdg4RZhMVoYdhk8cWEijMIz3xfHxJ2oHk+qF2i3/NT0X4pNBt9lqK0
h8G26VSwcICNESW1gdC/ORxd9ff/jZY6JOEsbAey7n34UqkMu05/YICHx7mSKeZhaMYC6+Byc0E+
Q/r0DPEQButBn5YJAkrdy4rafTPmyBHH3gJtbXch6wOs0p4Zz/XstTH/Vr98WxQ8gba6AvIuWz1v
L9rZrZVnaVsnMtQl/iHOosopx6UGpNZ7rqoQYzukO/XMmL19/7twQ7lN+FTgnhC4M08unLpJHry7
0JKOhuujgls/xWHr5HPOmH7HN/cRYp2psdgabRJCri/di/06++kzNc139Ig9aUkAIcOgBeHE8Tdl
2JC+pZfnj047+HnuHo58nFQgd+2gBWLMXrwG3ZaJk4s9tg9pGEEp40jsiRnVkY0ApY1qjVVvrvRv
ZpgZZqYc0yN7VVyFyJ3XR3Z6KucAC0Rty++ZtgTMF1ya67m1+bWDO8WfQ8KLJ+xk6g+M5cUjxbaX
9VZu+/2OozQsrUuQm4fuqgTGwCsDR8qhnY86f/M0RSEuwOtn6X5fGVRnOaOqw7RZdhqyIIMIGBYO
32xh9s/LU/TA2dau2oGeDSswI8dVLNV7JjPqjFJM1mkOT7XptrgvWmaWSXN4qkLTnOxxbkZa1cc5
W8NN+v3RajtTojo1c5LOVifnvn3WGRNJM2PyzdJNXJLA3VBnNV61srweuJt155Gp9dux7eUwmkv3
h3M1rFNtGDRmmfsxhzI+lvqQNfsjFF/DFXgn6YZk4pW8sz6/YH2tFvkxvswSwbCE5RK5ec9mHYxi
/39rmYu5IauDpYqL9MJL2ejzB9jtNLIRRzHEFaCoUvnXDqQFuCp16ovKbFWMC1LRaJvkgFkMmu7B
yoXMkESjbndcWIL+cM1nORXTMCVu6eAjbOrL+L/iTw8Ssa4iczPyzbmMLJUU/P88sciTcizvON/V
TEYD3d4dfLmtPjnRynY62Z6hDFtyQyxWByC/z+aRPweGuCHnlNXsT0kFJ1lsR/PW6tAXOsvcrIjt
fKAZ0L5E3OFdtcvNpSC4lsRPUGew+15vZfaHSrP2Hx9AC7ooOVI9ZkcoU7S9rLpxYwjv//KwFLWm
bk91A0Tx9O15vBZ1KPHmNPh72BrSM4QE8aYZfYC2KexFYDMxHhaVA4+NYQtLJ+BpVYnfgEjAgCob
Bk70Ydd/TK3SzYsU/rN/APxpmjUVd1RiWnLc7DxSuQIQC/DklfA3lH78GADXsIcvt77rvENhq5Pg
ZOY1xkXDq92qN8rtdcNOLcOpfNsXSlKPKOXWiWZ6A4r1JdcgPx6ZZF+X+q/B7wyLIZWwt7NlrTgh
QkU3mjgXbKM4bSb3rWZqYjEUBPLkDh3u5L8kqHVoeMf6gQG3lNDmo2sYS93TaRBf6G6jqcaUp3gY
ldo4pJSydK6v+3//fnXNYk5Qciufb/uHVDCpRKEBe+3/250yQGRAjJlOg8SvrQTaPGGzHy26Ef/5
iC9HCMB/ej+Gnvs+BuZKnzciL4Istc7srlBvFXEvpmCI3eh3KAMw7xkAnQrMdsLYMm0Akj4w03Um
8BIA8YSt1uDjkDaaG8AUak8Cqzoq1dVS5ELC7981Bh/RDqcBvsXZ2grKFaA51QVvtKjpQ3yPBBDJ
rhd76OkwlBrJUTStphv9o6aLbFjrRG/UmEYVT/q0h3OPAVc9QPdFZAfGLJUIdYWUbTk4fri2U12z
UhcQhqC2AZp7/C+9oK9esSyo1ikkQyNLnYnyvb85vCQBtJOBdDU4bgVX/l81gsOZ05DvZyOhG6In
OuP8lRbByjoW2bZ9OvqJmYjkp+GjaLfh6mtuRLRF2cfOTyj1EXuz4IO1ZXSEbFBVpAvmGsp9FZ9B
3gSn7sskM1oBetxoOwaDaYjwrF6X955J/oNgzp3+pxCRAQajM1lbtSO+as5MolMPcmYlUQV01/xw
ZHZJd9svwi/Txrz7WMStRWLDtcGKeQ4u3hF4oox6RjB6H3XezzLro7tFbz26PBHOSoM/wIzztLc9
QkWibjCTvI/p1ccvfH/ys9tj55PXv0G3RS3F9cPmR7fPihPZB9Fm4L2rmW14+duVtpS5dcwPCReL
aKrclk5hM4qBsftKfjzxf3SFk7tM/A4q47jm0RBS4l2useFGxRmKSiF0RyJ3zFoAKYIZU9PJX6zH
aF8ev/NGVfYl5RBJ+pcu/GtR+ZT4UNs64E/osykQIn7nXnv4T3dclJLd43NIa2b87CRxrp3guzgS
W7JcFgkUodofjCHCRUEqttFBmvsQkMfgQGq+ZaupLKCyEADrc4czO8Q0gVRDgKOWrCduN8+dC0I7
4OirsamS4ddfnZF6iww9dDoi0If6e9tKLYeNZYhtO1R7ebXBJHQSwxyYqY1EdmrQc658pY3/0lmT
rl2UdxEVUq9TgEeWfiw5i7NnW9bu9BT7jfBMc282C/1RJu6rGUZXzO4ZCCPhOV4exADGgTrpu33+
2mJSEX36gYrRpznKPcOqr2XYgrJ/XYje3dwj0841d3CaTbRYYuozlB2/r671t87AWsyoxdfw8MvP
3OkxC/oAuYJIJeF/7xykygAcZHfEUJj6WwE5re4kzJqEIiLHrXtSuHVCpm98n5igTdheDXSPgeBW
zBlPdspqTwjliMhVgbMoi7JShx3BeTvLN53wf6DHEvog2chdc2jWFN9x6OObsEiE4JPlSgCu5u1V
CocLA1ZNgv/63rMX6FNYc2Vf9kH4pEQRFMOZ/sYaWowWa3Z0fSV/oQvrVUBsYU0AqE1TltL6lVMX
+7y57IpCaCjf8/TiQYkubZmNwmK4EKfp4jXi66PSbQu0YAjOqC1MGilv8CQACSlleH7vHiYEHW0V
Q6ZwwkjkgvUYxU60hHOkKirhficFH2GjhOw/PzYtXdrFv8b5OFCmh1s/GJzN1q0i5ULo4qp1VwMw
4+wqTebh4cgRmVjVlKF9Lfs+FwL0C1C8I5WGwFimlbjPhpmTOV3zWSEKDlEH6B4ukiN7XnYKLgZI
jZNyiQOmOFKAecBKh7JzKz+xxL85P3w+pyOg10Y9bh2y8LUlLhbbH7RoGpshJvB+Ov87U4C3Ydzr
wqLzfk6hr8Aw2CpCxFh9h0TLbGLieNfM6re8J/KZp4hmoimB7Vg2Olt3X+Il1E5rWHjFVzoeyELt
X1EhTwop8mL5QKhAMdof9jJIMk/MCmgME4lJoMEBcxl9jzRQ4gF50fvZdwPmqwJCUNxJBasAZDBw
7wXWe2hrmSKthV7sVc25nFeqlwA3bzD/gRe2Es77rL+WfBDsCKPgpS0++WbehdMRY+uzQAx560tp
xFxs0Kdunn2l/DKl/ss0pujBAGGP/tL2nDWH9P/uhAVNPyln+wkZkI5izLjjK1Os790QF8Xw/CYH
gquRyW9s3Zv+hiboIsYQgzrhFgi/oF3zldTz2DI9NB5oYrUPA1vyuhVNAoGlhzOMon4bnWWYto73
TjKpLc1VS6rZaukZhcIGw1DmBPvbCtAkkNvxA6J+RMqflNLboCQDArY/fSsy8h+x8HxAL5NYAX9S
FyH0si8ccZEXv40Okt6DZX/ap0ZJMAbL+uOYSSK2vBu8aN/6YsqJWe1HuwHHkloOpodbdPI6hBm4
+WPvc5HSh8jhQ/lbfLCxGAysx4AA2qhb9gSsRO040Dy7mia+ehfs3jdjiIKODOIZb0unqS89VJAO
w9SnXap1C6paYABY7lEYVKB1DlrSsJXxFD3PseFtJDsCEpq2/KDrwL2586J9KgyxbTmG7reqn7bY
QAzCKv2EhSaw+QvTOzYKxgoG0sj78VbIvvENDt72wkPRKCIVE2p07N6Y9VrR8rxKBvvQ9cs92hJu
5FAIZwow/LsqHp3yskYLC6gdZMr/1Q3BPGfEIaZOJysXHA1b1qbBheKJHKrHwSUmXmykAUbVx4Iq
k9MNuAM2ah0lW6ugmj2BNRyrS0b8OZXOtq3JNm24CYD2OBbcTezzf4NCGwW2bxIpmm+QautIj068
X+X/FRZy24ls3mdgW2Lc9l8deFRtoVx1VxwnOgKdLg37LIKxyswHRa3m6k+DyOtGAXEplm29Y1tD
S8fMderLibarYwZopkTN78HuKvPPJOUSzP369MmoLFcuwQO3+0wPXCAkpKGbq6dwEkKN77AA+eUh
K3yFa0kDUsD4ZItVCbijapsLF5v6DUsNtK50B3t60stKXdF4Il8ax2Xu3q86necL0i0FVoQt71z9
UXhjTXp3+d3b4q0vuiLICAuFYn4ldEJ1XHmk4j72cXeS6fyMs48i4jBHoUheX6ScG1CFfNUQD1cy
Tc4Pgz6Dpx45+mrmYnN0IWPiAh6dMXhKBz0Ek7KSnYcUrcJpLoLhupwouktV08u7vLo5f4HoAzzG
4xIpjgzglNl9wqfyZu01Go44wN4kACoFJwRyTIh+rttVAuxdJf8wULz3XSH/mv2UVzO5qZUz+cBb
hpfX2/m+F8UivXAr30Ohqhh6bikT5KAjUrkT+R12xpEgYs5fUvcD5uo5A+/JnDej/8152eeLKwCx
2NzvILNfNdPL0eXhHu9zGA8Ip0NX9L8+dPgE7n09DJgt+/xmfSK5oCl9Ki5rHnqdmqqEo7y6auWB
2NNtJNmdiSY7XW0dVKGpus2qpI8UMghu2KQpEQu6GOJj6k2SyemfqKU2J5XwmFAn5xnj1b9ZoUTx
d1K+cdQjJ+GY3EloYK2SSwZWFCtOzrv6i0Te7jyKp/9OwTzDFnZUczIP8qAu+YkkfBcp1znLicE+
zUoHVpTsk+lLH2Zd0qLKndfGeDt9CJp2XIUZxWEatXvYR3hIqI8qDzn59C0VR4WeOOGTP/0jMOrL
fwpMRBtuM8zJKUeFAlClG/YCx9odfjhBs1TiRMeqH4w4aOOM2uczkPJBVhYCsMc957y/oWWCkvrC
IhX3J8IypNU8g76r737T2V/7p6Vwcjvj6YAEY2CAuFsAvGZk4lFFgQdR5G6ATtLwJUV6FzQyBmp6
UzYwx5LGIgarKdMPwxwPajeMz8ym0XEhAZNstCmfdk99wzL3ZQwmdU3Q2JCERfF0zPYDFBJFlS3v
REtoXVuCZ34LBUSFHVWTt72+7j7s5hCXV3jtqO+OwxGNjcxN+Kx9l8Hx0MhREKuZltHaRIPqt1xG
kNsf9LSVmydJrsDvvBRNBC+/jgaBnP8aD4UKtAJuFpEb0zxcQavSvKSkcQa71w6wu/GjC1istXJR
sDrYDRs5r+gxkc5dxSLtOAUlCwUPNwcsqtKKYfIj9JJJ8RukfCCZjR43J6VazaNq118s3oDP4v5g
C0t3F3zkdPGLX4RJF8cKMckb/fgNwxK8iRiFh2A+yESbWhIZET8wcwZfJz2q4wrLVP+GzV7u5ehi
PMlZwIDmuDHLQmlYH6qsWddKHY9kvnJnu0/amXlF7bnfbrkYQh+RkmtB4vZ9Y7YLqh1MMMm+s3PG
lx2ZwpY7mzSrhQ+Y6LVuYp5Ou6qHzUKf9mmStgtDMGUhsEd02CesoC5BXQIDh+xK3zGqgglkBkrW
8+dhotZoGgX20gKSLbmnu+X3FK+NJ9ceGngnp9mt8xeoSytbOi2t5qEyyWOyhPMSKswOCYYXdnxY
AyZvscdMIHcaTzHjuaPz+aPPod+sv6//VrFF3pufPI9WtOkl/lZDpkvghdHxhWPYPm9Vhdd1Awax
MrwG/vsCvrDNER6FSylJ69+aBNdS+T5MZ57WDNPvz9iQjhgwpA1R0KddlglnlxvzGQ4KwVZ1ihnm
yu9ThSimHz+8K99Mvt5Xr+qWVlvpqyiG5Ms6tSPed8+TDHzGIlJsZgSQigMjnvXrgxnum5WDhcTR
881chrRcKtHUFEEisfYcl2AH8g4U5jWxs8sbaNWGY8qopn2HUah+xyGNdxQgTbbFms+PgjMW0XEF
SF18mTBMEKEn6sLDUh32FAIFk1nUrSLjTF2x1SBXBGs33C9u2C3+1jvUY2BY7AYRiDsnNcauuBtS
+zAB+7tAXnIbcsYQJK5JiytKF+W9u2xa1v9sTMum161AhStgf5xZwQecmaBGoJS69Oie3UIvWZkS
UcnEov+M26RO2iLPcf5nJbtOvvmMray6X8k6NaDq202AY4hZbrVeN4Ji84rWS4V8jw05s7llMA/u
bPHaNnYd2UTa05/pCU8tvIm/mR7S8h+T+RvZAnZyhKclw9+LrMqWihsJ2VonlRIv1cL3mduAD3mC
mRxuj9KURyi3tpxgXQLSDY0v9pHgrAh3jaJYMEkrbWyuU8HO4IQRM6U5EsYaDd+N2m4lyywYE3kM
5tKJkw76E0nj7w4gSUFPDWniOWXwSclqz376tTtoO1+A+QZJJiz/BHtfOvkniWOm6FdcBRscgHFg
8BSEomANOQaglBYll/UQBXk8CoZfG7BG1UDssxDHjtzBjD/cnTFCkomxorbuc3JtI62rW2DWXO1+
cR+WqSy0MPfs/MZfn3oqlALTQtmZVtAnm454XTEXvqw+Yx/yKP2TSy7BTgyMqPs/IltQH/2jcZVW
dWfo8JNBpuWhFY5HvCfCVAVBvG9ua/z/fjt0RVusfSmHGJajyd+jlKtCWwNlJr31H3wdzol+56F6
DYNqH5xtwwinU/3EsUCV/VVY/MrPQrYmvKkAd69oRj2qBq8pvox0z5onVS65Yd1F9af8KM02ztiW
M9uTQFSVSgQhDW3X+78TDnA/luynXApczQZ+1r6mLC0ASM2CUJdPaCpEZWn9wEENt6OrwfqAXeE4
9jYpwgAqdv/xoWqNDeFudVutDB/Ku7GbmEWwIkrGgidU6cb6dOlhuNWh5LspAK/aX6fYJRo7+rYq
ePEGk/RH2wkNZOEIw2e4J0i07WB3eMRYLp6YjMyk7nDhLWPUY1+j2tI5EqhmrLlSkkEvH3Hz+o1d
F0BtmU1kh2M8T296a1yJsY+MPuY8/qkF0xyXJS6hrX20QEkiIphdVyrxInxMZc78GFrG3qUZakVE
x73IAZdJZq7kzcmHSi3CE4hK+l19d9BEmp2Py2cjqNhoEWTRxjhGGKescU8O70bqJJSf2nEhYFf9
BuR8U4TUy4vqcohmQeaQO5vjPCJHIdgTVt55n8/Vcx63cSdv8tvXFUzJhgePZguj5od8iCr5Obhs
0xnRb5vCgrx+37Rh4rBgEY2I76NaUeTQL3lsRwY6H0G85XqWFMcGyFYsOQY2i3M40bkKEXMgPGVf
9IY5vuMmw5jPwjfpqrfxi/gnF1Cs6SoF+C23Egk38PFlV2RedFZtsS4xxK3RPhww6dnwb+aI1X+Z
tUS8LczEU5OYyAAZ98AVBjHMZsNB1y5yRGycLS4XhURnsrhOYCPo594aqsdRKl4tIOfV/ifC2F44
A9st+eqNplYwzp3vz1N1h0DSSAIsw53DdF4Ma5M1cnt+G1lf4JuDi1XXo513X4bsjRacBylC/XvH
lmg+YERxTCzj7h3awUO1abyZgONzgSft9oLJCTln+jXiFOTJUCuGfG44ZOG5OdgdBcYcQBLDtuZB
dbIV0Pp8j1VS+5OADOpvD4tJgamBcKfFhumoW2EPegc1FAfyXqpqfQK4hRnkQbkcgKpUXXu2cJFT
u0kXZ4B8OcHDss20B0ye4lbJPG6g/dCyIBTB6TyIKAaoWmFCNsz542v+2cF8HRqerKfNAPae71j6
mHQZwG4udVQu3R7h3EO+gj9YI10DBIcFTrK5PHA5MLg1KKrQ1UMZYKaTl6rUBREzaa6GwGaLVgcp
FJFpHEKidTDN9wYKIR/WaWpjnDjZYzkrhp98powHMUpqEPG6qC7zDPI0mGnF+e4vHXmuDIdnI1NJ
nvu8KuDXxclzXcoKNo79K2lZEfw/w1fWJsRVgxAf3hDld3hJllvhYU6X/u7LAvCGMmb0h2eyg7zJ
MjyWtBzy9EjGaOo+VjoVRtksQOFQ8wrZvCZL9fPmVKbu+eb+LryGw7tVV5ks7cUrsc1f41QJDUOx
YnKECpIUCHc8Pv9uaToUSirumZuC9MOVrYGgRABK8bDeu6Jk3S5tj4S8Pi/LH9OZsPeZ71YFEJuk
08RyXzDqHwu3lopgsuW/Z2oes/vFAP4E/p+c/xolmJZNDZSWJkN3LVpHSd4SiTi6fAk0ceg6kcmI
4/UhJMXWOlwWoXxt49+eKIcdqKbDUY9/CrKxPKv38GcpXU5BgL7bVh2XcG5hL7ur27SwoAnWbwEw
rAsucPeaLwQq2EhPzivqNo2PWNI7ZNb9ig1snfXByeK/uHiaTv85kkm9xy31mxCQp5uxA9le5bll
jTRz1NxgxQd3Y2bMizloulZDeL3ffPOEMK/OBlj6YcoXaA6wOkOUwUcfwIR0+RiMx61gVy/smZto
NAQlSqlPMJWzX710WvMYkFZnoDGEY5oAhjMmyrAaxrAjhmpGfClXf6tgsgD58lT3cLciFvCG2sI9
AuA8LY4QfcmdizAzV7MIK67ab0sBSs2eMZOIeOhpIUx0N3JUs57GhCxlsuqyoW8yF5EALzd//4Mw
UbmVaqDt6MvUDfL6BA9GJEN4D+eBoQtVkUwkXjbgdanGoZVydQJMViDLGoLuKk9wCZfmMth5lvhL
+0cKN80ivvpMyLtybbQ6OOppheGN4w6UpDurTPgtq4Z1+oHaJRL6DIFMFYiAX4SuQT3bk8I9tSF2
mZhI2NU6DLxd7i/K5QAOxlSbUryvqsUjNbfBqQcn+3719qiBz9yhXyU3YEj2TTFdqDRQZ9nDU6MI
ZddicFdIpaI5Je1MgBW3VUegdOXXKyWozJK4MqIrjyZcBuFBZ6AVDrjb0dHJfOrQ0yCdDAbHgO2J
J8m75kKPLTliFrGeWjft/VBMqL3fJ0hWDAtvF4ZLkdA1186DRj1ZUDWbEth7mzQsiCjlo9ti2zv9
bpyCXHcrmoDi65v4gyyvOloFJ35fAcXjudxPtIiMCJra693iFTf+/8ghMUY+XwW5+MjcwVWq5QLf
vtodfd31AIQxSZw5yYQVN2YodEK5GAhf3mJVznCyb3o6j7tlkQwwrngybjeZFBufW3UvtcbCEWtE
0v/n86Jq5MgX/K6u9oVTxfrb+d3bc6NmIFFQFWPfj+QUGGpNa+udh/gZEWXfHn2hOgFqlsJoHwvT
kDvxAymonhptf1TkvNFhCxBJoMXYtq6i6KKmaoUEOLn2soAtE0bssSuqsudGHisLPYZJJ0a/CFOm
ofYuijPlOsyOX5knlYxmw3iBnnoXKaqS3SGLfUefQgOcULgY38pJfz/bicFoGdbkw7BWYmEIbrFU
vErZd7bzgoXLgMr3zHVa0sbc6UQtGQRqc6tjEdaWEKiYj7pG3qWGVVHtu4Cm6cAmd+qZRJsl4JcX
rGV2h+TonulqXu4rvRlwdZNg11HaG9SnxNOqOeFGDQS+daeXonCxbGZc3Ly//58gyyQLsaDSLt4p
OW5b8DaDXRjjCdNE8waKuRGs7Xw7lN3q9SaHUCt12geswHsy4ZDiD4mHrCQ36Wd/q99QuKZtchX5
NDlZmSEEMS9/UoHJUncU3ydRKxJikgeqr8HVO9tcbSXxQ7BUBJUPUFvPG7Zq6k6GrlFmGMDh8lXk
v8mCbayiyOIcUSaUprE9aHgOv7L2wR+SkJjYo47Tf6eN5L4GNscvfSEV9hbkiRlS2rligyXhNmEH
AL/+5bvgHutXlxHcliMOpSZnTvwulvQH7K2r/A03DKQqj3KQyp019iAvcQwzXF667/cmx7oysIuw
A8UjJ+jTrF4l1ceiCN7rQIefrrkMdrJEg11XdVZ8mXHDBPY4jlxe0BKjDp4dYwnoCjHzRutXylc2
v7RVFFiwGisON+Og1yjZTkAZeww9gAhl2LudhbyFn/6GQDwyp8xDvSHPw6uYh4gqieV7sHNm74O7
9JZ1TO3zQtEcvMr13TFCdeSXnzWIYYa2IrQBSMS4vXtFv3/WzQfd3TP4bgf11u38xotSM9PUPAWI
YZPng7heBzd0WPYDi8YKxzfzuIl0EeaPZTDehdgvqFy9k+gXlLEcpcj83cEsRBXP+sPviMWnnK/5
cwp6kNjXNzCFZDpnDuQoFJnOwGudpFBngv4gouefj5RnYsUpWT7c+v0ac9nY8WgNDn4eMp1iQD9l
O97/v7X9DMyzOnEkY3vjJL5t4B8EpPLW//CKVHlxRv7cH12hpbm7pHK/VlicQJku5DkGH2vre2GR
chrF9kQgP72+R9C9GzWaKofYo5TMGl3SPqwaq8sTQmwjHcf6EwIFQ1mwiUAdS0UhsqyhUMDpLVlQ
ecsv1+sKyPhqboliqx4GJly6Ch0/4CATKW11sPRUGEm6lzSldYsRg7FmyOSzXKITp5Yr17hCOujy
7N7Q3iTdQiDAi+JmWXx1Hc3nrC5OBeuS8g4jHpY/PExpBgVJdx3x1hDFiWtZjdujsxwEbkXwot1S
4TsPhMaSeKIFOl6atLC4gnUHu2eSnyan55cKFZdEvFQnOx/3Ocl+vV0CnVAgOI/Oz1LSH3uojhXA
pWxxfLAL3Wm6RwC4YLgCTc6xV9MicIhqPEsG/MgCwBiHqe3uICPsi677+Xy0IMH/lngn6Yt2l4uO
Jc5yMaT1s+eGZ4pB68k7rgPKZeTWNB45w5Mm+oNxdNxUxKupLcgjs6sfbqnFjW5KrVUla/wL7IOE
dTUMAg3oonV4IsDlTJpkGdEi/5J0sjHpA5y39Ijfbdy3orrWudfA4Ycdjo2/7tlKWRC045k0c7Mw
GELZkXTfnU6HYIGkzeNm0q3Y5an6YF2smjdFj5R66yirv8B+PjJzY6oagFFhHvne6qijUx+d0IfE
cean4wR875nXSIWI3HZAJc3Mjo077bvrInutTdRPo3o5rEdfq35P8AKWU8x66hibuuQbq06eVdAr
RwstMPuJj5hB3CH2wFBprZ5+Ms9fje8vj/Ikh96Bluz3k6TuepafatahHNP165keFfI9K4CEHxgA
P5qB3Z42Jkd0a5SmFW6AkKzbtZfa8ATnf86girdmeK55A6MQ0tKfBxrR0oci9v6kn7Zz9m2jZ/0k
w8utfPtwC0MiDKQvhchwjSV7y7F/D8TjFUd3aWz2+uLw1k4KPcD4XDiH5mzY3nzv+wfDMWzmbWB1
DHvxW+ZHUdarcDHEtDVwiWnqlc4wNGr3+Q1mDYHF+AFboDX8H63Wl0ycyXNEFjf8CCu2NtNbJJq1
4dSgNbs2ZcLX4qFfDKTgw9r//G1wGMHcqNAY92OlV/BRnwtMcQLLfe9HErJelNVG3RJPkZ+cYb+2
S+xlXoMGYNZXrsFnxfIRrfVGhqHiBgIX/Mn9eZdD6LDMQj69inb0IKiJAIlhQYRv2I7BReizcxA/
uhySShj2HzCjGQYXH2sksid7EnHKm1IKgOSut/QqmcUUkIQgOOaS3xuW3p4gN4MKhj169kvUSeaW
yniilcs0fvNZHBtKM0rehZIXwnnyQKX3fxh5DzNUjvJi3lxaJbhFvrX9FetOZs3fvm+PpvVwEIxq
HEmU/DlCs+7Q4nMffMTzN3cBNH+cTYtFxdh9VUk8jdfkkIY1JIauFaXZOwfi9RfFIIZ1AJTNgXK5
RJpLF1ClyHLWC1+n/qhPS1n2YGC4wDz4sMLeM1dkOFHqmoCMVZrV1RtXZu2RV440jLMDU4BPGlD5
zv+NTnNCTljN5wK8weprArGaC5m/Z0MgsfU+6a4IgoScvXNfqaiH7OLQBrBeElsR0ugW3LJQsCln
2RKZmPZTQTq8VG6TP2x3oaA0kogH0xvqLaWLYl0dewc8bcmt0/6pAHxKkl3eK0bi/mqAVWNofKLA
g4uds+XPDDiU6UwNgyOLATpE3tAyWnhQhpUh4OHtaW5ngj4fniqipIafKgqoJalr8FpHOI75AYZ8
Itut+JKFsuLr8vMJ8s4Z01uNThmz8yjp8WcYdIaph+GtodBXXorYlyXPaZYbmr/WnMkYMhw4Z+/K
IqpQERwoPUCq/yBf+hBht2hVBuDazKLn4dM45L24qiR20AvKhu4BrBVPUBSvpeDUgdb9L9zCUyWE
cRK/6Lp+Rlgjixzg095wok8mndcTEP0P1VZPbqjeoULlyc4ec4lxl+ZZ8JA5YOLt0/Lxr9z/mBYi
jti27U1oXZZ1UkMpUVfMyjoqiiH8TNx6bNO95+RfGbrzFCFlYaEvaluI9/zAMuOiZS8E9S+Y+1G8
DSsuCR/F4rmloGNOK/oQqY4mavN9wuZ1NtPtNUG+H1pQN0MXjuvTjGLELXKnlsSSe13VsKaGLRHJ
xV4VZ/NSZZr1X2ksEZNJIH3K3KmoysNf4Ez/MTI+huIPwaYKhQq0/rzrYc1JpA4Twi9GU06Pxu76
/GHkKBSWyZJY2418uJnSWp3L8z0xTIKRzLL6IKbYP31J0IFPjxDxhWSL1pnl7zBSiSeroULneft5
lCy+jWATySYYQDCT8ckCabIUhhsDjdo2yg0IA3a2emEjfe328N79xRN4aVdOZdQRk0i8Hya8BAjp
OXcdOAKILO9MRv1BYTiQs7j8HoR9rT6SIUiXzuqO3ngw0+LJWvKB8UHm5Y21t9h1gbZwodvOhT/4
aPBkKS+z+7zkAwYe/4oUVb+8XzBxaMXgeHs/yIjKU9bF7cRXKjbuIAVs5T4TOqjWZDpU4GdGXslT
0MxEd18xjqjj22rMkD8T868Vj7Qhc7wHbcxsLi1N8ylVki7kig22eovqg6K/VbSrhxw3x+zIFh3m
Zkp5W5QkdgH7raS6XjT8b8XTm8EOCZ9qJj01mXwMCM/oiOZMtYWRzyQtgHc0l878iHGc4CvrvDSZ
/QdBN008GV80dluqsblyD9VIaaU5fZlF1tR6UFJPIIrH4AkbQWSVw5w2bCrwlBOlUiHVha4jR+y4
thW8iizo0CleiO6EEmd9DwJBOUOCH6J1RNUVj4bQ69HqLoJNKKSdDyGmNJ+IWSHcw4hPOS5At6Lr
xv8wl6BijBfWAZ+FxAbKIgjMnMUmZELY/r5K8CHPFPAO3ntIajirByegUpUzfDsYs6cGZ+OvXc4z
ZnBNb0bIfKjq1N0WSxDs7C7VGdlVm8wiDVC5bBnuD3C4m2nvAObJLg5M7dVvjlJ3fr79AdikqCwY
NoCd7n+JINAFl2KCrfvvffncyWamHwHmA+FF0Zu2oaOpvz6rM2pxdcv7izHAbhQbqb94EFq3asWi
X9RqZj+b5Z5ZG9Zx/z1omQ87qSbum/xroO6M5BkLRUt4feLO1gsQI1+b8eVDpUhS7sR+DUY5cFCA
oCt4r+KwFqLflPpZZIAjSJGRdgmD6R1CjNiKpCv5vI1Tp7NGfyeWMGpfprB7sd9SFvA7XINdCl3S
i07JFb1D4GqbCpQ4diweiuJVDzYj1NUOEzAAjJca12SUJ7bmWCep1bKk1LqAo+J1LSdWAg4YNwNL
kT7XSYN8btnhDL0ck+C5qKG8PJrFzbpJdL29VFxC5gdfZ3rMtcCOxzYi9QCxI7DKSry5i/nnp+Cd
gmBSxMYJwpyDxRQ4oCc08mYGkPnQhkit/ZxZMWDzAFkA6EgxVTUdHdr84eZA9/If2S9ogimvaoTd
C/WTKHUohPBv1PLjfR8a59XOYKKsKjazxhN/Png1eDXl68h5XxIZ9LhlJqY4O+T5aerXkgGxeVPv
owiP4zp1z1ZagmX3PgPBjUJSNx7R6HAA2aVnYKqOpSNVi1RBo85OJ3dRLdvYbYjDFl+m6CSj/ATy
noq2gwRLTkXQyz0m8CaJ8STF9ai3qFoJtwz1R3O+IA0IEZ47WzMBICWjnmImmpYmZ35OoBUJGnhU
mqclFTg/9LpWERZL9J5wLDoNW2geLt6SM0Jw7lGm/iBXK2KxPsjKM5SAAKApN+2T4C53U8CfzHUg
y4kPqkdqIZkZb9kpPbaJPW3SaGHy4WbIfxsmwAr45YYTTJS/9NvZOtk/pno18CrbfadTFDzgH+uA
HWI60b1/jpM+kAUb8hpEp6hVny3GO/8eyxIrw0+rotiCwNkrle/z0aLkVPc1xoKVuM0vkRhhChFG
wYJO3ufew5+QJTRP7KSfHwQ/Eclc8x+1VsCXsBkPEuUK9IKmJsrFIt5FYNY2u64DUaytRIwYYx8Q
MX34SkmgBoaGMUDpxv8DukP3qMg0ZMXpH8BaUxtcOaJT+oxP5Xtycdg+Mx7AUXCwEog5bM74z/vC
8CF0H2E9blpfqCK5IE289sxfPz037nLP61sgNz2JZKGvGmXGdySggyeBwJtebgjte2nMjjVb25RI
L++SewkEqp/it3JgF1bKdqkJr1lKaJ+yvxH0l5GhPiz+9wSsXeI1kzM8fD9IGTIpbrQYnEVad20o
FUG7PLAxTiqrmQ8D03b5flKtXS2bFmbscc1EMquAzLyioJTWVUv65PyDBPAacTUyvjy5biq0hrUS
1AeBYGI/diZAVwSi25uJSlpLJZiar76q36G5lupAFmqq+A6wl/prEtSAcFtWYMY+8ouBvSvgfkMq
ZoqbZheilr1RAZtTmWAso9VVrT5HbxWp2pHk8I1d4KbjibINrwe2z7/3QQjAyf/XwWtFeGWzBxr8
J7lupTDqsa9WoA53JbqJp5k0aGYlsI+arLGIfVoFFFejTNxZ443+ylEsAQh9ryeowNbTHGzWu+Bv
kwccFm7E2L5Tbf/T8H+93PVU9v2IcCFbthiuXOhoNzjEvGRpCiUKEKJsBt9CbGIPOxAkJxo5ayBr
WCTnn1zfr+w7oYZBv0eMnwQxtUjnPJ4vHOi9YNPrtWJHaTG80aH8VI4vuDblqvq+0O66mZf/fqVb
xwG/sZzkTdbsk/RO9AqA32jRZSuDdFG4djOYyyJY+qP53/l0K0+3ris2XuK0LFt4X0HUpNtEk6hk
W/IxqGPcb6wFYhFzraKyAqmh28XZKEn6pzSza1HutqE3hrV7bPjhVXJkXZ0fnHLiv8RUQKjY2S8x
RJA7OQ98Oef6w6N/gESwitkcTjALOtEQQ7wTRn4QQHiqXgsz9BDysPRvTO/DRrWUhtl3RQsKTAZk
rag0QnpDnKpO/+U+I1ijKMAzPu8DLCGtrfxLEFod/Xy+MBk3bjrK2iA+bT09YxqSQV5wHdUp91Qh
eT81+LKp4D2ULPqA7jXubCz23XJ/Y7aVfEEdVLxUo3keJ9ig4vuEvC8/7Aj7JrU2Gjm6qtZ49oPC
sploPqaLAzweuWbm2JCf5HIvjvL6TjecTa2JNI767KfYSSRQ9KTkKtQZcISh7jQIrclUKsoD07IO
9QIzFHntPvTb4TIMMkk6FIWS09UrTmzovV77iJPf+j5Q7IXUxOVe9I/p6eztniILIFGQdBCYFk81
Wa9SJJ+hfbbvvEALSCx7bUB6mXyyey72mGKIYkpVUCfj+bH/BeFlXdMQZ2b+PTjoIR2kjuaXdB0K
mxyLSndYy/QLKRheh57OS6n7PJc1uHnS8b+dTnBYRUhnugEmb4tEOycPTQ60+qJO6Rb4uNgvmazr
+u5J76ZEZ6CppGN4rejoUo3muGhJTwbVR/lJNr3Sv38leVl1lwvodbG3CvSblZlM4f0KsaiNPiv4
KEr1y860Q+Kfw+M9FEQA77n1fQ3h+SktN59DrLHsPqLku+pM4ou/85jghb/px9OeI45QvE6lNpAn
l9l+ylZMgIKu5NDOLmM2jOkMpx9FSIL4WuWK7iI1cNjliSE2hwXbvpsx7WGjWagm1d16l3O73W9b
N6ntf2773hAzDR3+KBJeBT3uxemd3TopUxHtpw+ybWBBWtdlCx+q+WVF5snt/npEpZ+qL4jPs4oL
1wZjo0NUnZyD1zs0ZarDRgavvB3wBQJ66WtQDgyRLMFpC5+4GkIdDTUFKhLJIj1RdfGOtJLqRSzz
StWnFuS3ooEJDHImWJoIfXt3JWLhUM5qGDP1fKu2VrSbGBMT5Wl1AOga4dxcKknjp6w80MAu4mO+
ZU0dLJj6ZpsGwbtCX/1XTZDNz4dKPJ22qOxBjDI0SaNqueIAcjmAmaOIEeAquGMDuKE2+TZKElPI
1ZCFfS2jlXBe0+DF5Fxug2Eq3zWEhPDaH/1n5e5DvSX0pDpj4EX5D90sP8KVTexQXIUwwBpWysES
8g+SP6B/vpyNC8SrpkqcCqWpCwxxZVXB0AZMgszQ1wU8/Lv/TrowZTRETTF9uqlm1Q/ohDfmE6Tm
bJoYkBWUSHqbyOPAEnHrwErc6Hzjqxscw8Alt6wUcdkjKqq+Pt7xG9QK3eu3N4hKL7LgY/pV92jp
f+JKCmpfL9BPe07Ohl0wDHxPckzavWscUc6FPDr+YVLusXlA1jN7JTnhk7Izzu9mrSoEgyKi2NeR
eSdNGDPZpA5MOAfTPgdACHcJbcXNvHm8s9BNowpGGH7OcQbYrjD4vNy6o8+kaX9l1ulJmKM60rcv
lqdYqjVT5vtx6XkGOJrKq+rysCOq+Jvalv4PxP4t60RXI7iETP84xp1JsnkwXl5NL/4buGf5yKKL
Pobg4BeCGo4LpBc46G6+QnD4baFbh2TKltvno5ZiiJqL5XYffiCM+NsjKWMsymIIXjQSo46n+rGX
RBYCR89bwa6cQNn1x9KT01fOkf3vzi7vIrr35o2XVfTPHp+Ca+aTxx/mxMefGcZDT0xzPSHsmqMO
Ywe3EnT8Lj+thcZ3/WVGqu+ggx2kkgGbiJtiuEGRshF5zZuAR6cLb1aFILYXWMs1gvuI5uTtpcpu
I2O4t3UsHSiqDxtWgRYwjYgI4rrxka3E8dqaVdm3fjGE16bas2ubmR9u74HcIKDJapRz3+6wIDhY
1VHgP5lssbkKWeR1Ml5sSqiMHIfU+4WOX5xU8waR7uAFAe4GBKPn4h7atNkc91pV5IhmeYCJQjyc
OdwF9sg8I/3X6rvugENkp0Z4B1xBcrmvFwJ8kEOw6kEZzGgxjV+igE5cJMPJRm+8qtr3JGYKXFlL
lGPX5PD5ciJP8wvfcj9CMxI4fel1YsgN0DIi2wYPYtXgHtnN0ibSSI0f+M9URwhMbJxQU5Wbh23w
6Gi2XzSPMvQC3NKW8cf+AxguItK2mPMSYqoJfTsdAjdDM9xMMx0/aOhPBItrMdQMwuyZJ8SelE+8
pxOLTlGebnKXp3iK491uQQYy8IfJFwpcsSDF8sl1QoNtWqu/BjO8BnIRyTrpILDJ4UWom2m/5lrI
S77ofWRM+m42ZNQlfxkFP3H6ZfJu4KZ0WkvonO/ac9wZHdOSXIH+CZXQy90XOPxtqwpwLf04pdWv
r+RQ/mCxLSkuRhuNmNwajY4r0jt9PjN3pUUzaBzWnjn8E133oS0GcQOJ6165qYuEgjTsAQIR2ykl
GTNAHrkStzNRxiNFYJmhCPZKFadnYgzgFvldWvxs1ontfq1lXi5FDNK9dK+S6Ih2aFilROVk0+gK
T9z8zMAnUxWdpLdpNQvusA3OoR6Ib7TMMy5w5MDkdfU05zZOqNyesuu1OTomtRcSx/3fckRmi5I3
vguW7AOO5iOCI22zIVyu4GCp31fX9Rhyq8Z1nJPpDjiYSK9xLbsljhlmt2ZuGtIXiBSc/eLZXhZz
T2iTpvnVfw4fEDw2OrFmcYxv7NNt645wmLXYgrEewcJ7CpNEIejitfEF19aAho6BVcjbIY+yxo69
lrEthRWFkyPIz/kAB15TYS+scLm6rJ7Of7fedaDdQY6zPIvE+u38+bfAG7efyrokCYwr4Yw8+llh
CO0TEzauXXvfOOvCs1ERQMSW1JBJLy/Fwe86o3Wh+UPsEx4c9+uZBcdaQZTdiSgVwabnka4P5mEK
fb9TyMqp1riz9P2kKO8NoLmwVDBQb5ruFEwCczEzRDqsfQ0e7nqgpV2iMgTTpXIEowNlfIAeF0sM
06gO7NQGCfc/u9uph0XLvkrJX5KjYS6rLYhCWo4txfBzi7ofQ6y1IhzqW5+l8/+6NjEzlAC7vfgQ
n9sybkHwgAAhZld74dVbBl2gtCWYPYxQ/MVpd9Ugihe7xy/ZpsuLhTF1ngRbgXMKxXRV9XX2tE5d
TnATnnY1VhdNmOgVqia0SKyqbgZJwMVWSgBKCqorCI+4jgPoCq9yH74Nj/UXfzIWiDCLygQGboCF
BOPYrWYn0ir3sutE3dKjEdCPdwsxrizGi8QzxIip868hE2sFODCQ9bVRb/9lwxuQfRpcmwFmWgPP
hW2tQBoiaWftd9KUrj1BfVoW+y6imolhS828dSf6MMi8J/xyhLzc6M6q0FV3x/wbUSXbXw217okM
EseyuA6YbA+5QGelyqglhDrXFp3eYPLKCRP2KHDhALvN/MpRsZuY+AvuijJ95y+zjZU6QOc0c54I
Fa/6AJSvnANgJg2JlcNSRs2kEY2gLEWbV6zR46ZGJ/Y+V5tC1pllYB0VBNJXIuiIR+X7XTnpu6jE
ncv4wc5HnBi/eM7KsAWBUQs3P0YI99C+hE4LMFVZ60DPZ/U8BZ0KU4URE8aib9mxqtnnLumUwzFK
XmXzx2uoEFguohXKV7zUCxZ5hKWA7tJDqk4tuI6btj7HN+IfahSaC8kyVAsuNqq4xCdj95FuZJwW
MyivURJ3zeiIrIOsQ3tVySNG5SbzzWc4Pj0fKoUyNvGpjpSACNl97srZIfly9PU81uBcZzLT5eSy
EpxoSR3HxBCEi0un590ZEEdyizTl7OgNlNWkkz5dEJO9YcC35EO1wxn2sH8FzVATSlBYHQmniVBt
nuz+0ZZzgkSuJAwRY3y9Ph7yCLQMeBso0Kn0iUYJwIJr20gDcsZBXk38lsbKEVs70CcutDhKl09Y
0cZPfJPUqoDbWPe8K5Jl63jOWzYZg/fwFYwRDMs6g0lw3w3Nu8gtYgiRTqM4x7hAyK2JvaHqFaL8
C8t7N6bcn+mBzBuhMXBuWbNZnR4/Th7IZrCX+NI3aB2wiwS2UFadJvoP4BQDvMQilf77rD+xxZ2P
EJsj+dtFYyq6V2LBPLIUVEMtDuZ/z/yOg2puWiS/WckkHa9SODUeH4QtgrVK/H4dguwHxYLnst9P
6BvMl1y5vpRk7jSKtsj98YVy4s/IV/Zrb5t1DJ29ZhSy2M3fSPk3GqbZczlkLidCNhIRBe11fiPT
55sw7Ep0QTemWEAKm1N7+bCMs90jFWaeyVpG+jmhrJr4Ribq0zn2cTl9iKkHqUf6E2IlrYI3b35d
EiEtgOE315fK9POzx3wugzN9EV0m3sovGXHLB1O8Zc8cn3D8R4dcNchk25DNPVhuQ/dAayDlWmJK
HuPvh+0wyGHf4KyUNJBJWsOuo1Jh3oxsH8Z1Btderk98XWcvoZ84iIN/YxUNyrCG+iggqB3LZ+PS
hB80vXgp2B7Th6N2KS/kEaxNu3yHTcpjrgVde2OILE0oUMZsY8EyLwLfRKIaqPcVMxP4JqpvpxEn
Bn7YXLKBl4hBDKaF/BEVRJeUIEK68VxamYk1wM5iAaTEouAEdxNcSbAgMakb+kZgyKjpZxlpYXrb
HAejXHKG8Ww7u8RUKW9zsSY/X3KeVUGtz3W7+x36p0pclmyenSYHbujL6FgtAaDSWJeR6oB54GJZ
FZWGAR3w6Ca47qit6cC6xHvR+A75GDlc7lEXBZ85O3rEVggwp83a15AK2AVoTSn7HPgcbcNpLj9a
/dn0ikFgKFlYLSAPg1u34d9yuhFRm1OvMqU2ZCXB+Z/Vcyj2OL46i4JDPY2AW0OGbml+gfSQ3m/W
loE26NQBxSELigy1Oy2yVvWpIozn2uOqB9xzBXuE2MotYWrzpToL8o4MPAGlqCeCP8GHxJ4ZaNLE
+YiLe3YQhVnK0D2cM2DaXEb9R/Foadhw60rQrcBz6z97y9yJL8hpEhthZr4DV6Z8HK+MVHR0IiXO
8aWprTrLsNIBpivjiEU+yNH7g8ieUdyok8sW1mXicsLdBW/j5EmxNLop/m5gAI4R0IKdyg9BQA/Y
2/PZi7k5OTD/aqkDpGKo5vS8RE3B6HUVX6k4NEm7AANqnp/mEwcxDZuH4UdPSUZyK/Rwt6ITn7C7
Gws/rfadsWWE9LbH2khA6Dw4TG8fI1G1fGi/CVX6a0B2ax7aaUZW3XucJODWUkHSoiaFZvlSZJ2o
HaqCQnKp1hYPOLqFnOuo2bAZg66P5j9KkcOhQbzpsBiXI0153PGz3XhzmL2eaxtjre+aaudSTSy3
MAmCLC3oOt+/QbSoUomE82pTd0+0Kqsxvq/w4M+o+KMeXNqwWV2p2pr8O+5Yml1vosSDD6OajeYF
o537Z+QsOlnRUADV9HYYneivc+o7Z2orXswoq8XpKWy9UCDlelXE2i25RIMVT9r3888Fzoif2YOo
WggSXhfwH8YEJz6FLeppZj2nF8VRrk6tjRbUvo8imaWmWgxYCH0M4IDry7+nIicFglHF7kJHEjPP
SE2SxPr6mY1ppeqqbzsmUTYxdzYaCVaKGNzgx1TYFykdSd9Irkdw1uSDzdf8LQKyBKJhqHGzbyyo
2krk1yvEQtE8sDByx9h0UUKTlpQNicmdiJiQDfPIa7mlA7DATGWxmNuRGnzN2sL6HHLl8HAC4l8S
SA2O/yvpGqUuOxSJZAP92NYMLvOfsWF21jl+kRKNh7su6+Xzad9wdif3pu+B2pPVeY/30IhN6xu6
XLOVyj8xv5US3gODZc0ZKty6wwjtJEI+J6mU4cdU3/U4LYfq9iiqVsoEKboPAZRqVELPK4POpkcg
fszoUhkEpcn6600gjdgrVA/pfqQXk2nxU9gEwTwi60QeI41H0UggUUXPo2juaraAGPJgwBUeJwEs
MD1vbrEmdUV5uYEXNzrovPYUYdx4BrKyISRtSqlqiTxrv/LKkSid7n3wl6RTMH7AWXNIJfyQAeEx
y+00hBc5ST1yZzEfGoEgRJu15kq/qVV6qveAH50uzMBhS3KpD2+UkLaCu0FsBINAo5Q8FRHcbGU0
P3jsjh7SCfSDYA7ALYOxG0yJOqFew7vUwlIuqcLGE1WgE5FmNgadA2UTjvwXop96fG9FFv/Wlnsb
3Ap3g98cNQVPs2MdBrVsgy5d3zMY0bLhjQL+ThGc2gwcfNVFartyJy6kPuYvtrDDGNQITjszKg3K
NvB7u9WanpS55jCNInu6gjH6+B/Ro7JK2pFrZlJPEoyeV2S+A7rhJ8igGxkKyPObEkEWscdDQOJV
iG7+WW8Arx+t8pH+lI0Y9l0UktQJkv1uLcaFUWACLDuSzSWVEfbv5POm4rNpdMb6L0i4NFEoMWom
LZXU4Ry4GbLL6u+mC2JzEiKKY4upSBdN5tvW0CSwHhNPff6UcYAfcdsDJsoJHkFPjTjYdto/6wGu
jovxBcPusItPwXJ2fERolyLMsNF0Ntrnt5XPf8HKq6btv+qAp4BLJqxBkj7G+jPeUQoOHdiYuk/6
EWfF4F3FUoLIlYTakSiGh+vcr1WIK25xmgZbMr7Fcmywuc0CHX2Go/oz96viCfuja4i+igxZwcvC
PqbTSFhtnMi6vfFcNaR0Xp4SFE3JctNB2fKCeKBltgnLEXl3EAx3P3hpDabRm8YhWegTGixnEdHl
QFZ0R8gKsW/Uw6JPzLJs7n7bmKWi0iyhNY3KnU4Tyi6hAHnORxXOKsKI/E0X4nchGzb0B+KU4VLT
IBgXj+leK+BLKDiV3ENjq843UDDG+8zkPYT1b8XgMtMyaCDIslR0DjmDolrfwPqFXGJthhNQ0IKM
PpkrldKbdRyvQpx27VXyX+PY0A7yO8SVSQj/feyBMqPSvXq0O7lx249Ias/BL0xSW129COZet+FG
fqNCrvhgxeEukmCy2Y3Hz4t762ll5oR7yLsOAZCuLjnijBZV5xRqTxKNlKGg4AldVg8ba1LuJAiJ
p/g/Zl/AXpxQIXOPYBJ2DWtIXEeVs0Emj1XgyeKgLnZRBL3kcriwRHEds8rpq13dQFZ+c45t3OQ8
/DP32qbN5RG6J2R3zytqQYhF+Wv9yZOG13XWEzt5TKsikU6yYLi/AeZLe5n2iaaWJYknhUO1GYTz
RzrxjsTtfZIX220mB9Jb4xj0BxXUUXATGeAS0oMakGj9yvFDoMHYPg0+/fk3Y4glhD6avRPD7iPW
EsbcK3eMUYeYEvt9wspDW2qz62oCCPwIORkab57ITUmdiTKf4xF3cOEw8ZxLFNYdFqp6gdn0XAC4
Ib91B2lO/4B4zmvR5PJ5vQJdr0y9nmFI1C9PPnLzaROVNEr2VIHaATvJ+UZR38RrI/bK8et+IIK/
pa2Cgf9nTPRPjDdzs/7Udvr4AN+54oT046qXQQwvSTHy1tEqmvIfmC/nrO0clUk/dXFBpN12wxcl
8RMSSYudtOMA4opBwUBCwPinokKejhOY3Zci9HQIRIHdxMc3WSrQ3cI1IYA4P4z7muAfrMdf4kcy
6WMsfCy6vh+i+PBUijHRwM/sJAfUBBeTS48Ry4y0LS/ldpFfnEkmrsmjshPokiqGG5L1J3yTg8ww
bOxujJ4c/QT90iDIpw4ZgwVFjKRZaiK8uGq1YS49AnsWYXOorbHNytUEDy9usHaaBPXLdQi24/Vh
cUwtnXK2pxyEFtEcll0sD0n/+QOiq7BICn4fnPE6nnoRnlNLuecLmT7INl8A4ZIDMtzDQE1Hysfx
+uEiTZ9xOpXaTEBnzOtHuDHqaYCZUMbttVESTuGIFwIGIScshg3YA7UTgE03ppQlsgOmBAUPbm+L
dKj0e2DNq2KnC6L9OnNxlbr2DOZTFa6KkqyEkoOB2PlcLKND+SxP8xEgVmGG+RXPJSO26/yBVEUV
Rc08kLqnUL5LsV/F4OfItjOGVAuUtqgo9SSQU9+KP98q/HcF3Hf5HrOy26gjJxoIznJ6zh+TdLSs
riF/qYEV5UJ1VNKxlYlljOCZpa23LeHp7n1yh4it+4BXTgf+FIKbSxwOO3+4G5z4CI50LfgCiOi1
qUjaBHP//VFQVNGXBVDhjktq6se3CJexH5llMQyotVZTN232aSMNEf4yw/cz8VxsS8I3IzD+LKC8
DSyIPt7KEeUQY4tkAaPAtZdPzKTV4wKT1d4vWnaP13G+TahUOg/LlLC7vU73u5cMiiikdx4puisP
aMr7TwYpHpV9UTKpBVpY7TaQl7FDL9o+WPj1HhQoh/JBCIpREQxeHccjiPerZ/lsGXt3T0f6s8ul
6rXtt12xKhK622Fluc3NTfEk76V6WQFM32sm8m1n1HJ2JdwvUlkW63DVxHThiYzDnmViA2oAf5K3
I8sQBq8DRbRnYi1kepR+WkYeC+E0pK/XCt4BhKi/l0PTyjqoHpg4vMBFDe907RT4jgFjE6OPYvPn
dn3G+LL6z2VvFOf7jwpMkExD3GBbpbH8UvB4487jflKJUrEF9NwBq9lxB7Uk58oe8pAFte4vxB5U
lHO7otoUjjCv0I4hZST6hqXEFvWjHnyFIoKuiAFxj7dnA+rjLrMEqmfAh9/FopSmByn0dT+37YD5
g1Y/mB0fH/DBT9yW3gFWaLVetbLsB+OLl4/tlbQSvkzVI4gHcIF8LXO7TCcVHb9YWwoieMDYdx3o
jvEbwZhlqCcpgZtmPz4SIdyzqzs7vGRYQWD7xQo9vXJxC0Ub5CyPJYNCJznpWZOGsG8HDKIqczSw
IgE/h2k+CLn6s+sj8QEfHkwDrPLpIYUbQOrmQ4UwRnKJxAeNf3VHHoxAlOhvfiNGGHTTh9JAnf22
rsHCikAg71nTt2z39V6eT3KNAUNV2RoeO3lLYvQ6E0sZ8dg2G2igaFKQSHCq65XOCvgPzPwUna7M
BSH4tXo0139l74sibi7l/rxwxQF9im1AaooQyFZFC1nxWwxXa20TQsOYilfC8zvvbQw73XNOOcag
WQkdkr/xoiXJFaQOH0cmcGiprK4rrMm7N1ZXA8rEgaeIrK5fXs/XtSXsaZ3ud3RRz8bnlkMRgOKC
h2BQsNggTBfRpai+5Vuq4nXTQ6FBJJi9KJWiDYKkJGjX5LQvJP8sgpQQQNnAV4VdLaQPrSh4NJhw
80HWaldEXyo2Bzm05uSLqIfyJiIrlKjB2HpgRojUfadeTW4Aa7bBtD57ZM4Jx3+L4Ulroe1f+y7g
ZqfABZY3EMbY6/DLycDtJ9qJiyYj+Rc2hEz/zg7kwmaSL/BfT+4jb7ElzpiJIOuk+XTjAjXL9poB
e0iumCCkGxnjbQHLx3Cl4MpSaBkNdnHDK4qR31aOz+yFCLl6psaRrGocvB2f8snKhaqq0YHub6/w
RtYCtTys+kzgo5DUDMBEG6lg7xFemqURwwi13H2hFnqIqOlkdPQATLs0BTZhZfixHhVkgIbsmYoW
jWQWj65SBYh71mwpBZR44HoglOLuRJJwQAIsdWMpU2yOeR5+xxasP+sLRufsyPYAM2kujxOFX/pS
nBKwhz3BI9M169DoCQp9pgfBSH96SBIQl9aPPqJaRItU7Sf/YuDLhjIWT+zajlCfjrYiTQmTMd4I
VG1PsjgknvaYtIBfU9vcUJe3G6Cf7MoGPLTq1Vwhfkl+cRR4JRw6rtFdtLlwxa5oL0SNj/eDn2DF
AM8a+4QbErCuTtJseCEBDBOYGairdcZl44ePZf/Dz49U7bgSFJQGsjby4GqcfXLWYPR5Xzghbx8Q
sKkYgqHATSJXCTzi98KggXKdwo6t2hpGeiTsVvhg17ubKJ9UN8FayrfkDTmklFnRnAQkA0WXTGvX
mDZx9Ncfdp1tjZYJxh1n5mJG6StgT1KN2NEuXpnkjaFj/6ahFND1mGrHstzXs6XAOmhI9W0Ns1nL
sTmk+cBZZc4EJ5vL7kwtOEH73sl9g39R8uLGq6p2bD59ewyZmNUhxRIapsg5XJEvP+m21G30HNRD
XlMScz+TiuaBK9LO4I7M5C0XwudxuNlyfzl+9JfDhMW9BtT+Y/lFUtc88PMcC6jc3RF+128WjkzX
KNXKf4ZF/ZaOCvkonHlnX1x6Vyh9/fytaVM+Xd91uoG8Xpa6XtzLIsn/FH6a2nK8/TPNXFquHXjy
a1ZxwOCC/WcZoR8W+6UfHL89Ai+zA56L2iJzUKM2ihMqI6geAXR2H55mpXFfRasxuCUiJNWCCUwI
ISmYPadN4Hs8aIOiIAvrexQrtGrlLbYeZ02qsHQ1n/qihV9GKP9nQok5h8KFq7vyxtgHeyoCw3NZ
SauFUtGhbex2PT1qrHC835iNdAJu2DnwUt3bqAEqzGIV/+NUjG/3qm3vNBHrzTHhdx7nugIxdeQQ
uYP1Yp84EYhM2/RpA+K5fsWBYzjpDsrqNodr+wI+1sT/uQFmCN+wpF5EWhPCAVavzLxbN/5pGcTK
1+kqvp+ipcjtwlrfAUHxuX4kFC4H9vK0dsh8/R63esFkrmW+DcFjKR9Mxh7keW9ei6vawLWMJ72/
M2evjrNaY4CO0oT+mhrDGPvLXYxkyosZESaQX0vxUU2D8LWUAC/J3T6BdY0frc65f/3jWXdfPT/m
6drfxUP+Jt+DH+DaMpGUMngmVPmg7ake7gOhCNtu9HjI/EP9VvZm3mo7uFaGVwTqlXpeXbJ/aq76
FIo1CAM6py873jnCwoqNoURayaGXWqeaeqfbV/6191XjXHXxCLwajDi2m78di6/bSC+3p1LhqvJO
KqswBE4Co7x0oJGR6/0xGQ6Feb+OXucGpM1Hw/cH8JHs9RX7XBhklNiR4s88e4699ipKqto82YZl
8yLpQjsl4wWVd1oH6hM0DXfFKLLjUFSXmdGODuBw83d5zHFCulM7PwTRCDn53oVCG/sFIhT4EuZG
27zQHzDb6WVZ1xuWRa/IKAXw3RnOj+Wo4l3XUjDHJmeg65a8MOVyNjVpIOa4AQENkr+rkTqKfONI
dSW5JhXbU0LK+O9mFRK5Codb2w139Munocjv7mkJ1ejuD04ePoeMqJ5tzE2ppgLOkYTkrUDB+PVe
RLoWanxw4WBX76mqn5VhXiILsqTj+ZC9G02bw9IfqmpCfodUknzpgpEQzZn51tnUCzjuGpmo07Fq
9AWaeePqWRlh6VX633Kjf+59Himx1Vq4dtSFSw4uhxEEXRhOrk2oXKcXow0Dy3JVnfzfPChPDXa4
iUv6kEgtSnttvY7yR9D1LGoyuL1R4Vhn0ufaK3FIspfG1QaMuhitTPMUZvZVOH63nm/ORnbgSeCJ
bWNpf+exQK8dVpGS2yhj+2io1VRHpp0cRczdDBIMwjha+IZpidLrRsUmkfUDiPYze7eOjFnzDy7+
Nv3PaPtCs677VCjg5SFsHBG1QObgmKe5D/IO38Cq940ZGWf/0OCUorNRPzeeFctx129+ufbNT1CC
vdQKG48j8e7JEi+zD1A/SFetr4udRjUhCPFCzVIYMZPbTiE07+arWrQj3dx08G1u9PlH5wgzq1fV
cZKeFtIa6PDwJ84ZAjjLumdNj3rgmpSoXMEaO0ZlFTiHBJMUUiSkRL8XyvCryM1uiXMamoab4eae
PhnxVHGfXPks/lSGwU9XeIfahj6ObmXttEbdMCw7CegWweCmmYQqCQHtRt8BP4sF2MMfIRqA97un
W0Mef8ZOVhFp3VnUrSN/2LSVSy4pRs6jcRXU2gwl5hTDXWgRiinV7TCUFIGntJpjHGhnqnMZJqUL
C0enFO7wyoxJETblGeIWZmrV+6rVzfjfBgw6oahXosTTVX9VrlEdOC74dldilzyFsibDrgvC3cLd
1yTnfeuwd4hiJwTEQV3NX4aCgu3U8zZIQ/z8SZlYz97anO/3oh9KuRs6ViIcQmq8RpzOln1gtTkC
e3nasoVmv6CFPAQUxcyqdxRgQwpNi4mpKEs9oTqcLeGO/Ghffyht506aE/HbhfclVFnNWWDmIjPo
NJ01VXyvFnSa67BvfBb9FPTMCyrvhVyhrtXpswuNoGNbP/wkJocx4D/6jtYi9Qv5Rt9fY5r6lMui
gb7RBKAgnxusLkBmL7nLnElJLksk6etDx6MqRk1k/46CV1qv2Ex7Q+hkc/Y3iUsV9xjQL+jE8l/3
nql6qVqrz3mD1qc3acEZDrY68ZC+Js4jfuraRXkNAl6HkBdGRnixiv5AniCXwnFqf5ADkZFx1ecl
Uj4g0pvtsNLoU16+IsdV40beNu3ZZNewILfge+gSslYOciviBKFubQN0HM7PsC30Y9Zzmy5H4LiB
HA4FFjhIeMxcIYJUX0ENfQhFJ7/X/xNyBz+5ZEGnlC7yiiYOJyfu7ENLyHVgUpgpbTpllAYasinF
dToMidNFTUA0n2n7L/QP8iXGOpLzbiZsguFk7lewofn+1S78vYHweA27EY644qP/HfzFMktv2On3
rkDsGqrrVfE+Pcsk0XoPn9sj8MtfrGn9Cn2l3cyznZPX9PRdMRv88Vo2rVV9b7Fme1VafDGKqW1N
Uk+4XA31MU/Q6lX7SGKqpyAR4gxhMRcCF+JXX5ukflTZXvXXJ5lKdsW4i5mumz3DCyj45JhVWwSj
SNzZu2w1Lxa09MimoDhZ97KS6Dj6Bp56QWAfRjv/tfdYY92bVnd0ErFjaVRlKAZOl9cmWMbWa+xY
Wv58OohCdMQFfj8976zgFGFH6ZaD/o/m4NPBH0hb5YaSMYqO+yxSgVQHekLGrQ1kcYxSbtCLmScK
KVEsnEUFEi0LIqjkYpNNOc4qPBqx8Uc6rD6JZr+gv2k+nNdC9YmnFVTTym3qJhdpq62LafLRmjQl
cxRlVwgczdNJVNo+B1h61LKY68bNLS68TISSFTfMRbeiF+NQvHiqsICbiPqpE20/2FaQZD8p7sWo
PUu+fRLnEiitQLTt+Qxe29FRDG9DVHQrloQa4/4MNjoTCOzsm0/SHX+D9L02RDE7jRtxJU4TFvjx
I9zTqC3o9Sn1j3AZ1cyBm+aiSo4znMLYH9y8oDwyqHRWwaIaFA9NIUmn15GG4by32vlafgwpwGQ0
if0DDZ5BOOHNoAA+xY2p1emWyWtjm+oUAHQRQ1Y3YhdSX2Ub4aUMPP1u5Zn+umT36Ia/YUZY+sbO
Ph5O5B+eZHzLFSRKcU3vTUvpR1WoxZcxdm6FHUYs8bykH/e7o3Sw42iLiI77drZAkTOZVhTxJTrn
5uIzXrB7QY5p/ufmPZ630YbHF1otNpdLy2z+Jm2V4/SFvYw3NEMEfc5TpLtgh3k0SJtMA5mcMpzz
zG84Kx4iQJvX4zn3KHS+BC+qHXN1UDdM6c2WoLkyW0VIqGdL6/sdqG8mMTwNTaloft2qZSvvVZwH
B1CxXYtgooCQ02QGySLjG2Idxoj2BxQ1dE4FYqGW2kY2AZ7TZR/UifiEz52wp2+ty3HJRxMxkII4
wxU1WZEkJXSWMLzeD5CWonkDn37z30EkJnWBwlch1vMsHcI8RP7NkzZLsUGM5VYbOBYODVCt/svU
01Knop4orAvNQvq7K1r0nEcUHSzTjCeQhvp+af8+c5F9CnEg8wF99EUfkp85nHpiQKaiLZTTPA97
6X02YkTN0piCP7K32SlOy+3N5Pkg6Q3sI1OhHhfz3p8WyMYEQsIXV5vS0x0axo4q7YrsXalLB81E
sr+/0JR1c6cv1UzOcNdVLBgblf8eeutCQRaY9pa3KsrR2DUe766SXF+xLt5cavlrQXuFDN+sVmgv
BmqZmME3axxElSlxQkJa83Aon65crh3Udt1jop2Ht/iZ5uWbuZ4fBsHaAD6rxKTq/FFenQwCclWi
vwx1hZ/YbeBDDvDFKnzukD6IZod7l1ewhlOKGKBHstpjXnErE2WtE4BkIbhUR932Eh2+cWH7q2TG
l8r02yEZd+M2vUhIkYi/u3B3CAFgGr6Jl62gAxbdaEnFqGXBiCohpjyEvrWUozSHhot9b2gUy6AI
Gf41hZiljt2oY5HCo4Tl0aHzmXPo1N3y1iNUK+Ys5rn0JmejRlASogv+flF26PSsGUUupj3XcHvW
WQxcpOugB9JXw3EkbPJU9uDGzdfnoNtnb9QqqKAg9UElxS6xRSfihjbh4E60rLcuOelF9jNOrGwh
51VKyUXZsoj0UPXNVJcYxjxH2VTHmLzHiWicZeS4MK8iY9pqlYJkOdnlPFFQxP9BBZWhumc+MvhI
mes/pBwckH4OZrN1hm6fvyxF+qNolFj8xyfW5c8bqd4KvLzwuUqr/92XFXWdYli0W70NPk3sRSt6
Os5R6vL8KigqJXEoq5OQ/wK+sN3dtdQvEyw0/p1EyEbfX2Sjm/Y4Q9p+WQmgV3Pdzpg2+bOXLV0E
IRho1ZZ58i+gPAgrCb9nn6lRhc9P0EcXE0r3C7puCfHcBfKOGbY2/8ifNhucraVLzpbW+Xjdu/rM
uBStvhQtkGWjxklDv/BUcs+q8xIFp+rQ34gA1Upx5bVdP8oekZNfRNG0cQGKc0blhjOiXKwqCVp2
CPaU8QDTCx2pBddwYnMN3JQOMJscW41LTAsJdUgVsAGek7GUGI9cWNvlq3prz71ZkdL/mA8n5sLg
hoTv3PuX+3lbeWN2iTfHjFNpB0grLBx/9QkK9JWpGKaq1dNDSjkspPYq/wXvDrviMCC4gBxYKqII
b0pytRKUFBraMWU9B3kkTiongbtl1QlXdPQxqcjzMq8d9F6EQQ78nabOyUK/2aG+NNlvA0ECqrAy
io059ZxH1Q0MGK9IlDUNoLwVCb1+E+D0WBdoaTRh5sbd0bEfxKS8tFgPqMWTwtCXuVoi8uneblJq
RHEDrhAjvUeMGF9fCwdNsuQscq81CKrkqTSkhHEpz67SLhG1rfGmKh7qNJm/OSiZXnd8rEsAzYBJ
6pfEamc2S/e6RwnNpfwfhWsh62FPV8720Uz04V2OnOLVJYt5nEXXV0L6qgTHKom8EFEb4eUr5XJk
9VEr0/zoyTh24N2CVpOoTNnzvCYjeHUyHBqH1S7yOkb92N54P3smXfb6O+oVWMHi1Uj5DmH6uOwu
izLqiSYX9SliuNAzufCNygAdDHgpc8G8Wtv2o0NXbVtrI5eTwdJrOIRwqASvTrcKrKHHHMZyxslr
9G9QRizU4+ciPIoREhOSTvC+ZAvvnZNvRgKLsal4/8cQHmlbm3pXv1AIzxh02Q7agokIidvSUvvo
9WmQopJByMft9oNxl9SQL9G6IAwbGLsb3za+qKwHzxq3oOMwzOhX/NoZW8dGlYGi+5O/QBfi4Jnn
yXYyz2z1u9ClWpVVUdAnvmME07aad5QCiSM7jHx8goD0k1L2/Fy+t/hqFLN7IHLgVcsQwKQkW/Q9
qe6rLSauqeFfpa1Lz3bCv+o0WUahG0J4bJu8vEVBnKn2NDI6bgot5i3a79padwhMyri79p0IQmSb
noQ3/MLsroDBktC/cHYtJGjaTxfcDcG6m/z5tfIukzXIdgxDsOSYIkBZNfumxH89FCzbA49CVVcz
0bJ1+qt1wdjc1A1JS6m/ItnnNAIQJeE9lirATckrnfhQdfP14X81rc8OSvZoYzw4cBu7424L3P3D
/ZTX+AN0iKoPVLz1I785H6w3K44uCWEuU5A+yjJtWkeV59Mev3ASp/iZz11B/b8GIa3AriPtGwq8
UstVNlTQnlWAK2tuN5XXHJPiHSHdbLaNNmkFRq059Ub4eRVxRIUXdPcevvA8eceijPc39uc6ocoF
60S91ZzpXe8w84fTq/41pSbXuumqrCXgzxADzg/mVsbDp1ymxihU2hjKBMdWeSBsW/t2J62PtU0I
kcfncb+Tryer2jz5uBMggFFItas6cZIj4zQsGoHS+1uS+cIGyTO1eRdLYDS0gWTODI1zQcaS3lTI
8BULqviwdyv1g5fsFbKhmDZGnmDPmIb0qbhV6c0zRWRaus6TIwjTAU0babvR70ER3MoM0dY/h7qj
9vUwcIE0Q7WlfRJXgGzAxlEeSFdWb7/hIctLmjzYsAkG6n8k+NsDkBtwOZx6jMZR8CPtvlGJuTDG
AVRU8G1KlO8VRlUVVG0I8NFQ/KM4mM8cWLCVVoc7T7GiJS+fCmrNeuFk25wsuFAV8Gg063YeFQ9a
LHh7dPnsMQ/TKkOIDuthz3Tqru6CHiKk4VH7qY3uiAncKZPwemmlV5IQNxpvmYiYrp8FHFywX8Si
OS52wLB6MUk1DfD0OADSD7qr53VwkU95VRUThCbU+yIcRhOHBmYno1Mr0UOD9bNAfGVUbp2pYSij
aqamXK3x6ECPdcCXrirXQOHlj4JFDkq+o2pdhl8oU3pN4KJravTuSPqiMbUrH0YBZ5vfjg4L3/Pl
z9zOb8yud4IpcIjYMihlY7aUkR7lnbyd/DpcSKcGB7xKHkifwdKpXWkyibFGjQ8XZmsaK4AV8GsV
5TakyA8kRmGqOkfI8J99Z0Hi4/UK7Ay4r9S4nH9DGnve2tg2/vYkwpSxhyoX2wDdhT0ZXQbeh5ee
pISFcIxcr7BV2bOd1oamZrewlZPyKVuYFvo8hCfQ4zXl37kgv2vl/seYoBx6ORLo5uivg25ks0/1
qbYPkd2FL38v3F/c5L/oV1MlpacCoAuwZcbvGkIiYBTu7HpxyvpJMPo4nDQz1ylFPFJUagGdMUke
yLN+GAQmMALNU3pnkGN8O3mEBECjbbeq2sTDtmmdM9BBJ3iMrvgDzYW76pLbxFAVeDvb0mF7w/Hq
biG5PkRUHLpIGnDBZjkqeY5Z2TVIz8L4gqb4/sByxPHl8/YqF+RaV1jzLahOMzn6m/S3PUOMkj5G
Az0c5w4rTSh2/LtweJjjorJTOarF0fIybqDz7oMYaNoN+W6wxhwKYOSyQ3l1apYma0BOy/r8SE2E
tRa1BHylMnX9Ot/627QJwFpfAflQW1AkcvC+ODAq/t1SpMnRtqiblzr94IBaSWf6BhGkJvsV6Hpq
XQ8ABax9TqDY2myh3kZDl6gY71ZA+nN4wX8dB3nQM55pFfBwjSXYvWKjQB+fXV6TcTAH0FKuGca8
duAtDtXlDSYk62dqO5QXbP6L+NNPoADm1XD8mFbJ4cR2k/RdeVqWmO9F0O9Wbyhy8mW5BPK/UlXX
7RulIPZCFerDJy/mx0lWr8z76JsLuugFRbncD0eBIqUnOI62mFIOdoq7CsDQHdXOBkZqfgRFiCXN
4YfB6qGqurwEocDy9pkB2qGm9mZvaUgnAbETfL+SJegEvOqxkJXxYk5qu+Il2LdzejBrbLdZbw4D
0YRIaYRVbxg7+5sTHRl/p4yKLz+qAaS4pHVuSwY0NLpcTKiXhV1yQFBpUQbw/wLZtaAY5Tm9yX1V
3V10mP5ub1ED/dJhxcdTd2Ypl+HxsdvYAaYskzbN1CxfKu5F4rIPrfWT9PnkrCrANPSD5YY1XXiy
EugJLUy9vvGSUEconTFKKfkULCbBhD4JJDgRwh8dxDFilNFf9yNM+XtMahlPmZHke89evQhZw1hW
cT0vQR5EjAAv+ASZggeX37QUzqZvOLiGHsQTmwZK4l9QAmNgN8uKF1Bej61DZa6FJ+bgzk4oBiUc
Jt/zsRX03YwZIsEmv9rzNNPrQcZU22r+ZAMAV5Y0+Nj952rTldjsXCBzgiCoz4IJmAyNjv8khXjQ
bfTUi+fM04aGWNHuaz/iLrtxJwSppfX5Kn4rA762cDkgmpmPRFG7W6ydTB2MkAwa8hCysQ3jIoeF
uVaZGqXY6ldPtP6ELkiKgRR9bCVLZRD7TtionO1Fx2FGyHHzWZZy7AiF+zhwmZ9mD3T5leOpTDp0
+98fCSl8mpwPm4ZpUcN9GyO1sf1X8z4w4jprjNBE+wgbXNptqZXjhV3g0qerXTkwLrjXfNJPicZ7
Y7wG/eTclYXGyYrD3+iRtLgmV9VweCZv7b8l6ML7fjW2U5nZ6VU8UaBGBTWBYWLGSkUO+pL+KpLF
L4RTpqnvXVet8aaIIo0c1zFrNKYCZGdUJNqU6K3qrXjMU98SgRSpoiXl2DnxYWTqJ2b8WdfQn9zy
WHGIJYwSWBp7rcC+KrAvyCuFyOfrRmHyxqzcTJmt3/obtU6ZnY7S894gfwh2ZFRM23bpkoYPzKYX
NlT+5cgMKby6DsFmseeHLCsmpxXgM+PakbT3tAqEeC2o8/HlJZdp9YxDfvMsxcziayDtCAlnufo9
IPqQe9vy6K7BJtHWhk46Y4ndsm1PVrGy0rcwfIPfKYbj/K7n0PSKU+wwsxERNCb4jrN7yS9RFFnb
H4L5jHn/zDWnaD0dOqwMlj/KN1YGJ8LGJV0cCM7RZweq+C7auvuKNmYeD6d/FlkQ1mX1YHnhrByw
b6AnfFq8xqmLumIqQ+0uoTz+pV1PpWyfJLuFSopmjOcmGiDSZj5R+mkX9XEqD3lW/PE2COEdC/V7
mnqnXZKE1qUW/Av2M8QFo4Kex1YVLL+m7DW5aU4cS/MeOOq/wBBoA3EKrvykLhbwU2rgbCNLEfWj
AgXFDna0LrLqeFDjV1S0SSk+SldRt7pEz9W+4mBgyDMnSOecKQgopHx+tAnoBm6oif8fsUv8uE6y
44+Bpdz05lG9SigHW0DclgR9ScB89LBmWiL6Usil3Bp3iDl5HsI0RXsdz+xaoGZ4LjSpYW/robzw
0vwrq5xw4IeGvL7gVB0j61rMQGuL6oLSCozm/36BFABWx/sBer82fFdsQ3wEL9rsa2wXaM1Jel/i
BigKBD8YkN2l4iUal0wkWg6fLBBOpyvhv0nZWAgejDjIlgEPS8Yxty4VRKrv2ufDOdnm9mDOJUdS
5z8l72pbg6wanQlRK7YUNEkxcx6ahkNwzvVUYS65Kt/3dC7iE/h0Lskb7sjAKBC0kMZvbsGliHYC
+sfjGnS6qppC7ynK+EnuRcTd221ht3vaZTlrFW91ZmSSk9AEZ6IedktpnOzkplQXFH7fxp79ElYd
9NirqujfuhFZKu/I0t55mzBUowCzD/auDq09zZtFwJCBYdR6dGL9BHbS19olR0LjPLSIvBie0mUK
6dlolIkgp6sod6Bqe451pOygU/oRslrWZZvXzLK0DA6Xv0RsrdHYMR8EKkdE0s8BKNjjlquZazVu
53rh8jFHV3XbZWa2/T0pfd4ufakphxl+X1qpIv0ceghEx+f3n+Y0GgDcIw5mFzY0mm2SalKKE+zq
3Qww6jNREMk1ImQcXroXDbtcAqLIdw7ziwfb7H1ppK3ft8p/R70iI2DQhvOWDA9KsSmO9FhlXDI/
BZBXRM+KOa2Vaix/TG8W4mKDR3Ht5Y5R5RVoja4mnmZv0Mk0nwDU5ofFnU6ZEYl+OtD4LURZTaes
P/d49CDJyrlAG7joWNVdd472/9i2O1PIiKhd/SEWZc8CCraA0WrscF9NdIZD0zvIS2s0WAtH5ffg
5w2LKV8O9NVf2Q3u8HLRpXbdmcioIWaPyqEGJ7u4FBWEShI8aR2YEp9FNXlEAhz13AbuuS03JUFj
uPew7Of7JF8KKzt/ADCoRI4Ds3dUu91KbDJ0CR2+Un9W1wJJ1Qgs+vpBswI2QYZZPth/if6cQybi
VZeVkTi3fge6nGKDdrbA6bWey7h5IS2nyRqkvXBsCcoY/H7CDqcUCV369c6fyMRMHdODZkguleNS
BX4U8DqFBq1j6JD46cLbBgiNfzUP3XNGGtwrwURMlwvMYBmBZ/P+NVE6kCwTU5OTtLYfbgnkpf4b
De4GXXXWr+Ze5qx+A7uoX4nOwcmFLnAwdGrZQoikqbmIYKPcSKmE63HPBoBvvHWgnHYSA7TxmyL7
TTxIG+t2cPZwhNxh/+agJQ5dB2cvKbifb2hNf2BaXzqWG7nDx25HbPUOoK8/WibRDYmm5/EO8ikm
G6pewUgFY9scGSCLfycpFUGmZnntPe0DSqtV165F5/klyLTRos3AG1HiXoin4yb0UKOm/WQ4Y0dt
P0zcboXRIcMWHcxqn/5mQKjnxkXSG+Oh5ZMIihsXdi7iJLi6eeAgmoOvD6TS8cWvdYMjJ7Hr0EWT
psybjdeh+R8lD+CsDqvSBbPN2f+Wapi3XdhxQ6/ytWzLtVzYlWAL7JKlDSiBrkaqTHpEpNK6bfvj
L5XnSi008amqn8EqWItdJsen/AftSozQ6WnyWMk60EtQjKVnEpWIVIQDIQNDZhldgQqyBbNC/iWN
kpuCb2imqyIKjg2qraYD0VK+wD0KA96wsKn6T9BGlTkB38Z7/YdjV7C89ykIMnKGqxdT2VHsvYDP
FWSdGufmsBR/zkRRWxFmjHtIbQqkfu0y/Y+hoJ1UmE0S1hTwz3PF5ZvDt4UW/sA3ED6CsAnDMYiS
kCOZiYyJjNgal5yK5fuWMuVwnyFbgtKMoU6Y0RH96JzKEyuExfahSkgzFD43QTYOX9OsPLOz0Kzs
ubnQbUfSe1Lm3dh+m/8nitizi3P2nZJkvKxoySm+tuytz0afmzAxs3MJ0eQ2KidIBv+HC1ASPfVS
Koj31LxXkOwBCVHsxtW/OuRqnln/2CiUOrNZOv4p7IttIS68j/jx6/tp0QmQJR3u1B2AmSfE7v4i
5jyLlEpbjeet9Ffga/x8/IH8vnHSmKWrmWkPPu+Bny7giUXU1N6bT+wIrv8ez/XnfHTQDIi+uztX
5sgOQxSSqvtdDBCfofhQ9lBpzp0B3Yh6PhxSmthTGmhPJhW7nymNcF7YeFRiLW1JXLgAOENEdte6
C/tSDP/vlSAGEPC/Phb2V+0hYjAP2ZJMpYHFy9ZUeN2QrfUEsHatcJbStJ3fj3uIU760km4Pp3kz
VqTOCkxFoE4TRsI1nF3KHY8Nue5BHnW2QFrZ4ASGvyw5E91661vQl1sCqJcpJ3qb5ErG1zFF+vvl
X+LHP+zDuW+B8qSwjtKBeW7QgMdy9OHSh6siIaUkbBvgbOSDpmTR0Tm2FgO+zMsmO8zYL0gLJ4Kc
9G/4VpQpJYI3+JZyxgm/JjFllEnhXSBHRRsmxvn63VLNYCU9BnI3o8mE6jvnzntnECNIrlFzRyNa
Zv8KOJZkM76xQXg9qNN8F69/HXp4I62moRsahziU37wFA5eFUa18DNjYQufuQ078955lp7Qp9vCQ
XHaJvQgddu+8G9xya3R9gGMhz8Gq7XY+0g6F/CCq4JPVRhG9ASnrHF1BjX1tob/0k51u96gWofa+
7nHfSdVCuEd+82Nflh4aAZlsNnSZPz5RSqe3paObg/UOKLE6erDwFg1TAtI+4u3edj55ZkhnJeWk
NZG2IOgmm0nUoxZkIgRmKm/JPoLGB7WDlceFwJh/rRj6xStEjQe2BBw19ZT+KVJGLJ/QbjcQqcOF
gZKWMvKWz/Mw/+nGJIHZjumm+TW4QBK/SXav/LUalBf3le5dKJDlOV5Ug6M7WSr+ExOCP/Je+xgv
jdM92n7H+DDtwzlxXTNkexjNklzXJ27o2K5olbmM1EQhiSyOjJv2oX4EYFbuXqo5ypFAB4vVTk3t
8Bata1pOiNEOPBefr+6LEmwB47UK4m7xTlv6cEeGH0tfMZTjhoUMlKR9vQJL2g5vmvcFkqZVBcHj
G+8b5ZiwxD9Tw5Hn2T6QJEqvmz1lroxYj3/nxJstobaY9MQU1T2sQRAAXHFoTkmEsHFNSZhXOzMO
cNkQnfxOILsLIaru29OoxEiMIZTh5VQ+ZUTF9tGzpmsbD2QIKeBeakFwybP31nqxSnyzm6IJTNbF
ZFE59gBNHYj3kccCSLoo6Ml+z+oEp6ftTmHKDX2DqJ41VEbX6v9eveG2dH/V8uIi8uLQeGcfa9nT
s/2BKp8lyf/oxRq0zXTLufcysCVx7tUe3HPNQ5SRGFl5TPEVh3UeWyFQSv8dY+Yp+UDwdkdI2FRU
4GdDu2+2sd6QQhZIeALzFDvnq+IwXy6hRX/paic/yh92clDLsJ1PLT28kIWsSx4ZlZno393EkwYH
PiTdHNZCqUQwJpCEKUPXRKcvQCVrvr5mLw4sBjVlEzXKvp4y+/RHUwNfM3isSbTUCgN5jIJMCZnI
Ta3eiBPX+MHWtrS9VRhmXcw69j1RsdaO7/tF8K9TD4ed57M8L+v5uSHavW8WxfhoGO+SQNnAlomi
hgNXBzxBLDXCYnU1ZL7CxcXcKvbRSheR0pudcGimlvvsTiGSfOIqGRTz12Z+gqI7UGM2du5wpxgr
FRyzc673mHZ/npR+tzDjxHGuzePP+QoRiNiig1Ek1ndAQDqSKC1AVWof5PgTknlAMu9PZcAuFDCW
DGvz64I/QVWoF1pgRhQhY14CBJhUEX4lxOMIgNBqPlievW7SWDKNFpoqNM24WrGE/DGJeZEJ44jU
0cDimy6/LlfwXYkElcKme7b/62rCOTOVuGa3XvQkn18U7Aai+vB5ehk9tBqDrDuOVBUOgSrIPKOX
083gGdSHJBkYL7yWY9Se6qwt9hvDKeCQ/SeXIxbnOukc6ASUbJ3PXDbgarC7Tq//PlTCYtmIemQ0
J8jE7gsYDqsxCSnuWKy0jNVtpI6ae+Yx4L/bqZLd+zS6ogdt1TT5WhkPDTsY6wOPpF/TE8jZiTNn
fxRqNKIgWa5sR7PaHqhRnn5ezeraw3Eam2JkHNPSyzGO4uDXFpViWlQhoTYxFvURIqEyDj3xNseV
qTm0CtMPcMuDj3y3823y9gd4Jwa3kXtj9KFNOeEQawo34cCgVbxVHF3ugw7XKxWZ+3wQOK69xedW
ARz6iCoyT+5ociOynKUlrAn1b0VYEBEQJb719z8KDvFROHje1tP0ZWyL3f4mNI/FpcrS6nl2R93x
/NK8vV7HL+qCS47DEba/XzZ+ODGxv3zvTSlYDSe4SUZXCyBQ2/RC2JgwIUNqSiR8ljw5qDkXC2U1
j35F9xtNf0y3B69u0tR2luU7x3Kd55QbwREONlYBKBCUpKmWkhFr+qu3UJGHtNxtMdmPp+O8N2gr
pVVYVJOP8n4c7AAfla1RTfCFbtqg29MzG6s5vml8RbZjMAHzuWZsyUYGGxPP4LJAaPec+jmGU636
gx4vp9IhGBdHklpXHDJOFp+96KQThieElD9U40vYy8VnWUGg4V6xPlqWY2I+zQJYGbFdVWc7cKSZ
cyOnkSBcCogehngvzZ5yZmwSz1tsdHwXg7/IfhtM37Twm9pMnsjS9Lzs6oa1BXXzGov268JQboPy
uy3RQ/Qn8rZC4JYeN/fwD4jJ4ulh2DSkdBKfCy8teOeIaLZutj9As60sKZp7xM9M3HdR2LzLyFwu
B2UQGUIY7f/jOJ44tkUEAz4UiwQuaL8bzJz4gVt5GJG5co+582ehEg2lnT8qNV0Bpm4bZaiOIh0A
R+H2xMjUKumYU2tORsvFIDYUhUZhV/vAAdpHpMx/jtL0U2OvoH69inRfQ4yk5WY4irrM/vY1dv2r
LJ+MBcW9b5bV2qlLEY3c3OlGkNrH+us5wSrilixzrZ1UfmTioF3mw/RIurtXS/rX/r9UAQxEFYrH
Hy/CIGWbwN6Duc7Sz/ICL8f2T5lnLAatrDV4imFYVGnvsGPCtS//EO2Es5Dj/PGnTJEuJpPXbsmr
N5FAek1px9Pybyed5XORH9F0ptZ6ov1cCb6QxKmSJsFRt6vRPGiXUYqJ5gFIb11MmW0b5V0vpb2U
6u+68zPz3P3bdpzK5/0yD4iyTKcvYKfrn4viVS9ZeTY672yaEXfatL9sGZd3YTSf3qn+O8BMmL+Y
p8kZdd0fV+JLk5gl7YOCZcFuFrSnCBwGZVBfUcnyXdOaqh9ore//7a8j+DlCJhykSLvAmMzUGG9f
1kHJqmmrD5fREdEZquf46FB0GJ9AbYqItgC/8LR+rgffb/TyC3bwSwPxjpu8r095yjQZ3POaHmT4
nC5fuZqHCHgo06blJ4OJjhHDxwSrE7Gw+CCY2j8apFiLqrpGrZo2zykPeveAQBH9adRjrdzK6V1i
V2T/uIXFPzxkGoT8fLQYkVzqanGdWWIiC3Qlm7wU/Lt7MspvkFpfNhf20cy2uiG6M9wCshymSaFG
lurAGObR7zANgjUDFkXM7W0DUj9xjerIsZwxGEx0FTAA8w+2pbNXfFUUG0O7Nm61fMxjy5/VHHms
7FV0vEf2TrvI6VwEcAaQI1N11EwJ9EzIiTvRXkPVtmtWOdpli2IY+KBA3YukWTwp64QKHBi0w4aB
PH20k6CY/RjZFa6iKlcHdoWyyVMVEWZ9QEkva6Q18AzANriJ8GL4yeFtC0qEJ20k08HMhasnrGtS
mylDoP4QZ3PyR+cYYD164rgnhqApxmM3QCdJ/9Qb0hNdWq8hPsCzJR4DhfgcuqjWkBVA74uBwHHj
VbqZoEutEw3U2EJSnMAkk7fO/mt9GZQ6ui6lwaP9OANCzyCmgTTgLIgUZ8KwD96f4rWQhBKCSOEc
U+Df7gvnA2urem/zfAgB53Be79/mL0oMYOAS/oEjzbvon3U6zOxVndHogetSBGOizJ90oszKgdYf
8sPKhChIbEWD9malO2JpSG7ZNeHshugUJvdNQbGkSYJwc6379LXGXJf9yf3pBRmW2SN68b3Vmihw
EhOP9DGAusoaAE33pN1ODu1Q5rEvHAdTshubSr65J+8qE2Bv3cSidlYWZWcSbBgHT2n3bH9fxX7R
sfdj3cN3q9a6LuT1WCXEpSJMuRDsNq6R1aeUrx7Ba0SbjGOUCSCwkE/g50GsgyAYsb+BBrx+mfdt
BRaPan9Xsxc1sHIXuBNjiwsjv08epUOKDoH3bUDbfMG55kb9RdU50m18mhVb/sQsJQLlLFv7OH1U
QA6WX7Z36nQnqzrlQ38WOwsqXMPsGsf6ZECzbqwwa6m6Fr9IWPtR6s3IPLreeeiohu7OGmi/ktME
YyPJ85OXNSjZMeCseDLuFD3UA0EI/lj2XxXwEz2WFWzf/43PoFz7DdkYdrWIwZC5Y8XovXBB/9DB
OvSx+JNW7O5zHmsxbPXXjBSHu1ppJO8TryJa/EVwfgHMN/RzXW1E6BPl7DLhIx3f7hLLLLne72Kd
R1mTaeSM5AKCCjeOInckcqkJtJMW18pVZNv6mghCG9KO6+6bLcQRAJJAQPd6OpwzCPuWl5Z/zt2N
QE5OP1ea7sifSxgsLoAkztESrJNLiIUj2QrklxnwMu+0tL0AICWMlPtMbyhXRzWmJghSOTpK8fJg
csvUCUrS/lCJsE6FsFCYIKgYDhS9SCIZMKx018o9YIO/Or8L7OpDGSS3tPdWPNCgJMfDP983V6aH
KpFdWCNBQddi1oXa9GE1YRVWCmu+wo+sEVX8GM91CAREQFjgmiFv+7t2js6uuPToEJq1p9n/DR42
Y1brlSViAv9/uOdYBA/o3AUiLQaesgzJ8ihn57Zse8eIOGp6UIiEuunl8TttAXx/EU/Z9u0ee6Jy
AJrm03ZPV4dZZRUMm/7Mexg+MtypLe1UngbQad7en0ag3z1vuKmxDaovoNi/XVXgtd0TS1G4aE1f
q3rugTaN8L6Vabz7Rf0wOx2FyLy/oD0F1HBikMCZn0Al3zqOMm2aGyzjQgWh7ff+p0pgl8+eZDRc
lc24Ck10YVh4Qy4HJSELeSqu3BuSZ3SVqvta6Dz9Fhkgb/4z03t4njwfMW0y6arvhJPXac9oXxHg
7jK013YXWsDE0pGkffu7y3lhAaSaRCsVIPfW+9ktF90N7oLANfQHvpzindsBDxS5+l6zZN2Sngwm
c9OyzBl5TrXvRhGhtst4+grbtx/YudRP+2OLYr7Wix5rIMHTuqjQbWhVvhAEw4BS6KP0HFweJ4+p
lJZlq2yIDU1mCQi5B988uMerjWOoDXRLN68695G3ltsa4qJpwk2wPl3/3TvM8ubRvaVfwLfu87Yu
PSRzJbUgzz3ijfS5kfrTINbEwjQgRcRduIl66Mb44FkH0x/RPf9i67UGMFDaYedzdczdfyFu9gPy
VjSiP5UbqYClhSkFDZ7ISxYZyvGhGBBChvbqiQgrNxw9oe/eUR86yK+IRaFyHWt2tYRUTyaiYM/L
y0NVcN2vZc1fKVEQ1Zgq01jJsHlceBarAuoAOrJ96DANWTe58Owlm5qCdCl+63i6czuEncUjXifv
MxlesZ5bI0STsRiXtja6n45T/n9ulHl/qfaodpXveEbOHiFI3KRficKnwDliJDx5/3dt4RWdLJV8
E2ZmHnKMJYcJdOqPyFksd0FoTCwi/fgLJPelbf7P+G9Q1uZBOF+4Z3AU8T7M0atc2alWy2G0Ptrk
NrkXLxygYwye+e20+FrCjkQD0Pz+tgskvoqesQM0DjiQq+8dmCSWG5CO8sOWathfrspJhDdHkU+V
Q9jBeSGUyV3HxlarFF0pM3Wa4TPsWkqXWP9g8+StWRyCoonOO27L3dqJGCmsFrXQdDr/Fjg3ywUb
gM2/UFMl0XjkdPIdv3D79Gw0I6dYBfzcJwWDzTmDP2mkwdA/jrlb4rll5a7K20CzELRtfPx1CykU
GB8Be2aZg14xpccnU0ApmUYUm3pt6ucGEg7xOCFKtVbT7QEvc1rzp9YriWlQTfb1hIge5FwLG75V
Sxu4SUqGMvGXaY6gu+PwYNEkryS9lLq/Z8MbTqYtWFDAg68B6khZpT8Y2EjVC2vHMJ4vdWnzzCtR
Ka1xjvFKhxnH0uCjFD8UJe2RV/9We/Xabgdb4tlWuEnLZkO6y6cJLkEHz0j8wxmtK27SPNjFGTzj
+uhN94xm0zKm/M4noFhI8aQWclnXDZYzqQmulPd7PIW2cO8TS/xCjP9PYxubD/AmhONjSxVzEVa9
5QiWf8QC4+YdkaJlBOvCwxUEcSHg5YeIDZc9cvAfe8G387o2djdpIB/8JqxgPtg8Drwv32+hsDJA
oF9QHOXP1ZaDg9dTxfV/F1zyoR1nTpitj/CdT17jXqGGyaE/wymmMnS2U34HYfA4EJl8NGlYQz3W
+V43iUC840v9ZJH9ycqc/BTJnPHXqnUqI6gufEyVwTLk3yTDQ+qrwutJeb00+8dgGaITWhSbwTPG
y57Ry5CsG4XRp/MNkBEjW+OrfGGK6skIGNUG2ViK0b020VdPiFuZCuOBooMvC1+VrhlUMSukTjb8
9RehUAxESBvzlCcyRiMnRbqTOeFF2sG4DqcUMgDI6WZf0RA1V9/pkBiALLm/cCSi4EKPe6U5MYGr
Ebwj/6mzUiM1xKcae7dfGsu9Eqa1ThCrmiTZKIaTd0aVEXh4eHgMr9uIs+QHgBNE7PNY68C9BOFV
N1XUNPiYqLgXCzT4UnS2H6Xmm7fQ0Cp/thisS6cGnvqoU5dXz5299HLhzz8W1DppNMlogDM8q5z3
2w89ln69rgIfJj243B0k9aH1T2E8xYm4rAXFIZZZ3WW5Qh9ERtVeX2HCrrM8TaaXzS+3VIMmkTKS
TSFh3FJd3nGxsTizgY37M1IfCsnqHOrIvdKAr/kAonUGo/XFlJ/B0sPe5RAGYgIvOimxfUOu8xOy
V9NkHnjw39ER6IiTdeb9XdRHtU4UDp8gfOY1tiwdoqxPFesqWgver6cnGo9R6MU1+8Xt+hZuYHn+
OONFlSod7Ztyi8fR/T/VtSHNr3KODBlsq04DZlm9CRbIobg4lmWO99wZOW2Qi4qRH5Q25QC1OKYu
V/veeC7R4yIld9tZGCnn4Vj5XVvxO2bB8aLPq6444FfxrOIB+UiGp+IYlQIONd6In9ZDyj4hpznx
U1azM15GKwFpjIeqkTVw8jLrVZ79SY19Nk8jdGyQpoAkMxN1ekWdUsbdkQTchcQzQFPsr48Ph3Iv
EwUf0tCkBLlriYGCfCR0ILl3RH0EJ1VN3HupTaNOBUe0MO+bD6PCafTHHl278kmKHiXyUl9MyM81
bNN+5g3vwPTQLiga5X87mbyaLlLpaRpH4GXaTN7bX/5wSgzNcffu8y4KDpQBUyfg7ZOPPpNOEuGc
XVpGBwwHdOsMkBnxv/Uhbhv3aoKo5zT0EbXthQwwo4VtnQLI7ulQ7vdoGNJqK8EpwyUmP/xL0tXG
9ZohB3sH12EHpw8ZgfM4K7lz/x/yJzc3W9qUpJIi7xE/dpd6eIe6kx/f6Wli9L0Gb8Ol2PpSt3sL
UCjCJzJYjWzlYf5NSzRlFCN9oP9bgPcJh0Sfo0tTF3m50HuCr4faphqFKp1dIjODR5w57Cm4aWqc
lLOF0IlJW/sF0qysHdB4+A5xbH2nztnCnrwt4O1qKnsoSlny9pGGQWUcdgO1Xzlky9cBokkRzEy6
L5veQ1M9djYkNH+qgsXt8rjCjgC8Jv67XrJ7lhmvoG1U+MIwelNf8x32I6UtnsFPEoQNfDoCjreI
fzsa0npgu2cTgFIikH2J1NTHjFMCbTXdmE3P+AJnpM746IyGStyt1YKOGh2a4MxEBlnGckNUiTuX
YSEymNMQukI/PX6bXtQtARsDM9Es5Ke4iMJwwed8ZkWdGHSlQ/wnaOH+PfhZCxhzljmnXmgcwt13
6IkPdWToywpwyPDdSOEbVgrGecW6rcj22zBEZcDTmN9crqs5ghEFLxES6rlXpzcjO1cRf4AUu07a
5DdGu+oSiLBvevjWfMOM8Tx1ep9Fz3NKrH1vHp1h3kRWnClBBqPISlVqLqG01p9h631vHBHw/jV0
AFIgWD52ABVVkMDZdqxJDIwiTF2QGtnh/zQAhenwg4n7fgKHnQwFci7fswXloQuad2FmOztf0NAJ
0kQJhJl9RbM6ZEVMUbfvfvU4vD35JIqa81Eq5HQah0fxD5pBmCb5/4UpQnb4AXx5rc5SWuNkNRVI
3UjJ/7MO1pFFa56SXzvPPLnyaObaYqDXnCeq/rm42jA64HYyjc8ojt6lLDkcNbxmw6nPb5JcGv5q
qLlkjbbSTZ8Hckil5qpUKnVbxz/P8/yk1GS6FA17qq4y6swKkrF1PbcWwmkWYxEZHsKFj3GLpMdP
2sIuCbE9lMYlU1H2m9mt5UbnjVdojUuE2Ng0RQFMRul2a3axooGoRfsqDda/EHYwapJyBlEdeIUf
gCzOCLnaTnFj1hRTamcOR7UJ7JRbkuwqr6cApG+3WDmM2v0kbFgRDw3JnpJAXDU9WpOuyETjgQVr
1Q178HMYxH7sfCxifK4iWd9MgYtJWMXqQ4wbeczWMxvm0RYKuehQOqnvAU5qOUDI+UFHO3RPShay
PMY001LhY/+pord2Se+EgMXgf/fUwfY38ypxPa0fEIfcgkCv+tWLK6/iypnwhi9u4fA+6+G9AY5A
Ft5oZ7Qpc/xd37asK02ezHJfuhBUv2JFXYGQBhPime6FgKf6DkbSlMKUDZrzW+OOmXZ/cDNJWjcW
LvbqmrRodc0AKOzF/yKlKpa8ey1yZa5BiV4mcHqhmdqyFxQ3WOgN2zoBU932jWFMm2J/psa5STko
i5vvLtGwl/tocBCy83sbQGQcQsRxGHFsk6K7I//W3yn6XRHI+jC13hJ7Noi/Y0PBiJ8YYUfURlUX
hQpk/SPDLG5mNPEwXFmxEbPoXJ1RJsKvXo30/0UFaABIin5/F6hgXdeJtsZmnm9zvjRXYn8yYXI2
qNUbRFILBwgDi2fuZ7cMdEl5YGQWRi5dxfnadDb23CU6Lx2wxEtDxjggvOo7FWhgAwcaZgUqrlpV
adw77RhcUQyVDZyjJraOsGRtfhflI5o9gk3YXqGIDv8mcziK4PrRmVEkoaiWcpxwm6eKwXg0D8bB
oMA4drS+gIBVV/cYhL0tBPkWqvwS4HqmlRAYxisEsesrltAE52+qvoAGWtwBh0xxrHgP+CMr4CAn
eKxKoW8ih9R6ZnUmj0KhOGj4YFADg1HUQJMvRHCW30zT/3wCDwHBskU0bx5hGiUyL9Qy9X3GbCyn
kFGEVMv4HFl2rORqCRTIoxp6MtVJJ4PZLQHhdiR44Xhl9ciNpLd8Xh7mOzbP/P3UPAp+51kbxMrl
p4lJBIVGPlLBkxCAVKGkui3IbuqUT8l8ISWP5bG2q6NlH1YlopRbs3X+VE4OmUQkGqmIENU522oD
kPrTkx8zkeK3LyTaVY0NMsibrqR7utIHVQPT2N4LCZQI7eyewvYbw3+yYRJ60w2WQdctvEW/NMtp
MwDm9KoNHPMGfPFJbcbHHlvc6uGuwASj5V82AOw7a49Am53Ev8UHQ+qGBCdHTg0mkjyNHsFN2Xba
0/LKXYDOkZnisayCjEysfraZCDoYn1DgH+MU7hptQpIjXxe06VIfCc6lCX09weEIQ0LijfrfBbWO
rvrqYFEhU5g74DxIv/1x3HCpBDoBh1+Fzc6mQGuRfnSCQWQHV2GtUMqAslPl/6DNf6D5aH4HPWkC
GBXmxJoJGwY48tFWXLnl+Xv//S0CsryggkUsWjyAMuTUz+kwWFnVBKqoHFEAUZh/7VmjFa8Cw7f+
MvuXh1dHbFVoSf+R4bWb7KZV0KoMBXoRPvkqkqGYAxz02e//tssq+AKl54ZCI29QGtVUd5NJ+ZeP
3frXN9eYSrhsbqbkEmXh1qXjaSxgIDlHDoHFDNQSOOSG7wAL2OxfIeGM7WefEQV/scwcEOT8YaXT
KnWajL+lkyIscYFUqGamIM9G1as+A6RTGLjMqU+XxC8iA4yJMxJN9L5Oye4/dAJiKrUoO7bDNTIW
3VO2S5zkPEECo364UW7rdJZRGAXG/BYgYB7CdPlkK5B/iz5Vlm0THVwrL8REGWgQcxHZLKEvDzAE
Cysu1VVfVpWDzUQIfxmZErJ56kIYjLl/Tgo/o9IZO7CZlkcz0HI1m2cx2aWsTgaceOKJFrh9Ln5l
oub0YpKlOefFVq8PcfGEPn47rWFidJnEN2ZJKY8MJUYtwsUcgpIAT3BRbgE7FQzM2RAPQZJG9xnE
KxFqqd4xN5dnLSBLCtAUitJCR8iN3cF9FTGUuVb+yfbuwcsbbVGf3iXC+/dF2hBA4rHL0LiLRbvz
vit99T/WN40vL0c3zk0Nrk8KZHDovEAzmtRZE36CIVKPF2E/CnuGRLj3AeXPpSKoLKxmFryM72vj
6iehS1LpOXXg2nSddA1JZcgyXZBTg6SJx88tJwnLBLGdCkSgazXlTVimzNhtptsv95OehDVC7nqK
eiWLvVCllUk6Iu4qjQZMt2+bbK+2SdLtCOx04OEtCqJRmZ6/ORScJjykjo24/rqFSPrsMxDmJdN5
OFu2+MgNcYCR95h+rDBTblLMl2pZsHQSwxr85V2qKOuyasGmxnBO2EGVioNcZrG8ODiSbmbsyVBI
mVlzE3gyPNM0jkig8Lvhc5asePTEKUUB2b3SStfD6hVOsstC7WCFyQw9aUaXGsv0WspDwWTGJrul
NSpm2K+a2BR7yQP16ty+5xEFcVJJm8QKUFo74rud6W0OdZksvZCZOVj0FfWNP/bHtQ8ZtZWYgU7z
GzFLAzwlZyvanhQcxdzgPlDBIv0lQCIfMT/LRfLDmsHalFSl/c3z9qjQg8X6nIE43o0WotlnzYg3
6a6IqqRtNnIdkf/6+wf/9hPCNiWZXJQl029Ec/kseg75ZT5mCtTCApfSk9F9W239aon1phgBFW/u
57zB1SbrBJdaqUEyhlliY0LBfDhWY9/sRAuTIAfSNejtb0XUEjjDqyLmiaGEw6H44Y++s+7Fcdfm
XlHuZnZrVO/oejO7RoT1HMi+9el/5v51NPOMrfJGu/0cX6jwIotrWvtXoiuY486+9xyHMGbdSz5P
uuzvGL7twF2DHfFHfqeiLAT1MJoTL3lHeevVaxC/OPp3o5Awt6mwfThCpgJayUEd0kLQ+BB/CrU0
CG8ql9xvNLahaBY6FAGGyxlE9J0slep44Oah26KUWOA5wrcXAthdqnjF7ed6jIHlzNN9UzOXx27P
7XIckRZxXEuEFUrYyXngXuaVKDNLUkAo5UJJdI+fPBYvswjA9U5vn7MECKksGBp+5A2kETvE/7cj
iQJXRuUNkL/BVHkGJz8uVHRmozbOUVVM1RNomQZ3PGoWpNBoGllZGFdzD3woUoDEGOu1HrpSiF7C
8vYAyVRrOHAIickfOr4PedgnRfy3/BayjIG5kq063l4KTnp6aMg15hu7jkWux8iO23yx4noWvQQn
w40oB5A2/kEBu7sNIMfkvxL4OuCnzHyS3FtDVXBCenHEJiS1swspqxV1HJTJ6BGyF2KqJDfbRi0N
0mqomq8U2VHylPAnyZvwKCeeY+v9m++B7dH9IGjRR3FrfhPkmomlpGIZpF48JhRIjf1TXF2qaxNZ
qkAp+H3ehWXxv46wksLklCIHDIqcHdEtPUYIpq1JHb3zwx/8z7aJHuMRFAHzlDx5fygblKx50aeA
OL+iqAQDtf1b/aqHH1xWHW9qhnSw6Wx9KhV+rr0t2XS1OC10FGvA7RkNYq5ZQzCXf2/L5gwKHyMj
mYVwTGmgjfn2YJlrE4Q2/5pUdYT1MUlIGbO0g1z2ri0T62q8aYZsC2uy+Lr9KeK2nTeKcMVl5pdC
uDCgkAu2dsSJK/wTItPNMzaQZvK0aR2fct25YXyVsup+tmpIvBohG/T8qLKNqillxiYBjuXJ1ZJn
gZ/fk5BlrVQUuWb/Q+LL9ECghVYP46DMkuKWz+OnpeXpuFQNOje6v8PcUkwGMjefTavwMM1Mk2rH
MsUpnH5YaJYjHiWEcooR3FFatdsiTTGe9q9IYwFrBkmISm1Zm6W1xrjhCvTZB7D8Ndnwzvibo1k/
cRn5Rn/os2jZOFzvdnrX6MgJboDzfdXJ+M0Sf7XLKlHcWQQbExBIoa8EWAGmNSgvudnNMfyEMpoz
Sid965PZhOgbJvJRI8EmwuSaROPe2iROz1GICvnd5kg2Pc/Hfm/Ixsag3dd243T+afz4xSciwYUe
cgqAt1fsw1x4oG2QbkR35X3gypKD9NcFjXQgkWh6MT7zm512Q22hc9rABv+7XyudmFCErp/pkIQn
JP6Wz2yAtKm2pLSHXICFd0oTHy78EoZBnODKqMpRVuiLcN9kV6aXM4tXZG+n2QzIVmTWe0cbRCxa
vUSyC3ySlLEJcW6qdyaoB22cM9x+2lDUY18HoFtBPPW4VU4BF01WIBwMtsheQPzBqssTPai9W48p
6YMrCRhKOGJUGeSXWCZfZsWfgU+JpuoWDv0MLuLNcvPXTRKWrmjMbWz2DPd8HfqEoPFIRtyc0eL6
VAIqjKIc4ufFhbgma82xgoV0NuGH53NDEYSaA2vYFayu6yCPMcpo+bAvIycGz4gmBUG2PEoP7Kdo
wNEu4WOb91k5Q+lX9WGDYm22O1uK2glTUFIEm7NwaD/dc18ysUgYLCEWGQky7KTp90h3KZyTDNs5
Qrs3u2d9IFAo2oZUj5n0Te/Crrdf+N330hLiuzanXnmdpHyCRcPVoTv2EAq1fXk2mKFXb7kdC2Xe
UfQaaIwEZsRObP9aasWT7g3yabTaKhuvmT+DDlUHhwiytLfEmMcwSkhXDSBcOkqNFx+gc2dttsa7
mZ1YNMmIEfrnlOHwm3+QeSYm5ciieLVdipJdMt6dQrySfsdo/cwHAkTjU94ynvo7mG5RXh9R/Vmp
fVK/O0zgnA4iu8KR8UjF59yCuSREY5tR5qyvXHvpy7KlSX7J41BZOykRzG4r4qsARRNuzjfVK2Qy
J/cjY5ZULYA9wTIc/GRP2awiDb6xZAwEGuJMDdocueN4qeMZwug63DFEHOAoorHSa8Z8PDuhponH
Bj8tZM50Exyw9RW05dIkRQsIvrxXjNPs2zPovOhaPdxKd04HsxazjadEHpiY96/4ZP9kJertuyM9
/6jw29BNhACx7UTgnZflEup9m4SuAXYK6b6CwednH/5jChfnhGeVn3f/ZdV0lzVXL0ZAIhNToXzr
gDX6sR/z6bH/gMGpk4X+FrL5ASmVyFiAZOWBV2LhGwKCaB0326njB+zTYLfa6Ht+7YwHpiG77ttm
sOI/3tcc1d25ycc/YuynnOEgEZ1o+AaOZUdcWzxDBxLb9FANfGIl5Jz4Ca/YekE3Mow3cBi5SFdx
VwDr6bxay5FBGDzE6Ip5pZqouRDyC8gaAyzlDNnj6yyp3AAuAKwdLXo7JpkGbvQpZyO8VJajpDWR
beXi1fBK6PWUdRCaJHJzsfWHqptE1dhCqryMD7zfj7XwU+qMqS1/7jqrxHUjFAmWg7Z5w2bmpkbW
BfJ8jqt3AsxOoMzxYbGEroa01iRn29UbQY3MhkA0H24ZIfdJBTRLiskRRLKChG580LDHKfb3NAdj
zJtQhm02jEzHL9nUB0UboGaJ2w2qb2PnTJKzrAL5KGdXdFJsjIfS2fLhrflj1BOM39l49XETE2Hf
dSa7ymbDj6kqtUmkJXEBTgyB4U/ECgXzESzzoEyBYXulkA1QLBwMMFKgDQW+IX0YganBbRUXN0YC
hmNsTzzg/UePwPIShfVBuLAF+UKWXS+H3GOh16f2Kg9vJ3/QpOR11HzL7Janl8sUKgqOp7K+gVh/
aRSiYzAdunXkaaMPOIRKi67HHey8KkJzTNtBVqgN8ehTWRqc5z4rpzigtIJm8MTFgiYwObd3eK5r
edoirp9FBC8XU6eG/7F3uvepQOOQW5ADPZyp5J54z4m+L3/fSJyjaZiUw3mJbZqe7UUm5qUww0O2
5dc85wXpaLRbeUP8hnWmzNEl1rGcXpgZDJ/vT83TzFIiDbV69x0SGj4SbXd0/O3ff9rzIJNOU7Fq
bmQv92SN2Nu9O2Pr+pzTg5wJeSWQdEaKJhO3saeKxSJ7YKNGkDwg4ErAU+WMQNePT0xjvNZWN80K
UCbkZ/KYuHiCbDw6tvTVp80FoZSIQMexrwZ5PsteeM89yo/8VIxxtPuZyugmB1nnu6i1EOZ7Y1Vw
bOafbiQcszKjmBy4nQW//aoNgOprIrkOxFGCo5GM68zLp/g3pP8cf2YNeiBRL265aa+loHD+MBxs
gX2jZIjyEeT9TmZrdi0yUzz4MjeHkJbJ7C9cOsJJhno1IUCSkD60XGI1IaJBOup7MiaDLdSGN489
0npoq7lobWo1yLQO8t67ODNapLdmHCv8eENpensyRDhkdaBYpn4Fb/Rt+DcznceWbPPvazdduado
NIoGjo7vItB/ZlphObZICyfDd7E/dUJgCa5Z+GU97U8A4v+9CaPUvY9D6XZ9TChaYJ1kqP/L3ffp
+gJtdZq0YfKJAaAkEKNG7nfXZ+b8nc9G5LV+qUqsG6e3gwCGD6H7n7TvyqAwdTgC/9fDEy9uZuQo
I+D2vMpBoYkwD2aM7PeoXuQH65CQE9F+HOOP5r9TywcfzwfcNgv3DsXs5icGN+MhfbTFFIIyvjCW
iC3zPyjsgf2Aiuz8hQyssLbFa11sS4iiexFjXY1leNHbyujcFxNgFNcaPHYEUTNYTtG7YWtbvC6c
Ea6osUdWrYTqjhOm8XpMSz9xRKni35NPBJzd7jm77Mzo83uBpEy5CiSPvewBZQWx3cIE8TTRKGR/
YYq+sxdKKQOFdxZzK9oiBYV8AJfQYawEJHHXFQelNe5g0zvT5HpbcCONsW0aGokGoJDhrotk914F
XXzlIXS/uS4jCgHN37IakOd3IRLE7X5grUWQYm3mFqUt2o3nIC8tPjD9b/VnNmKMH/ct4ReLzGYb
pNDbyLdBqKbBd4/Rdsu1gISHb2Vz1XBguGAOm1g0ldFIGE9CekSkQiDatyjJdcYkaNMnPVymdOdt
1prmCsc8J3bDiY4/nsXvPtzGl6+fbM28N5y/cNAkgrPsKaM+a6CT7iinES0D9Jd6tW72T7o0rN8f
BEZO5F2ApIbLV5ygg6ay2jmaGD72u5iihEFm7MQy3OUunVLFTEKeIDTmvWrEtOOY9J70YL/nU0IL
6+FfdbsrlxJigwqZHStZM6tS51hsi5pEQGmOcEQcZ87jZi8ZrJgC/H/Y8JzV+3zYA7XsIOwcv9sC
w7yDVWwf38pdoHwhRXtXjSD3K+e3aE2RD69xAEesdZpOP4pLvrUGKx/XNskB5F1r+g10H21f5GuI
Og27RUV1fVq57LpUq6XsY8FNRXuG42Tow2MRglCOljv/YtQOJA2tj3ETBqYSVvGK30ELdO6beERo
1HSn75qU9GSdnujoY3ZczAPyfC3NDZlw6DaX9RgBBEIq7R3hhLBiYliKD+SdknsNhvPse0WqC8gq
XzDpQqcriSMTZm8DB9xjV3Yk4SBGEvLJFnhrjIZ/hDGprOLn7cAFh7rwtNUgohv5zYTmuDPi9XVy
599w+SX8vnEWoXe9lYtEXIgYoD7aioKnw0GK9n5iJ9wsd146WejeB7+bY4wkunYMuYaubMyYwwfZ
Nu0LEtfvrro+lFWwtYXSlRyTpBFfry5jcckBOjiI8lRCcFHuY404W2yWooGey8mt82EnN3oGimKD
tLxLcT2sG24oid3Y96y8Vga1znl3VnBjui9YZTNzonxf9IH98uY+j87jbiuODwVEoTV1zCPO+LYj
IpHkjWqn+uopn5+JkRtjsFLoNKersbo/Lbb+mt+f3HujyjDsaYSQozImfyu8XdjcsS+h8L089XVh
6Auj2SvGhr2T4Vb8wdSUXcfs1IHyqdfn9Q3kUNLEcq1AdSFrWmYiEkPb+w0mrWrYtAdTKiIKvpFo
LktFLLzxJMF/X78SjQC56ewEBkQ/BE80tXQoA//N6Rv91rQAIaBB5KXiD4lplDrER8OlsmDt5dsv
poo8UAu4jSMLBvQB3knF0TiD9UgmzceUskT1GfWz25f9LtPYOxxugbgoqqWqlKEKZI9XB7VaiS4o
4BRDXoTFDPv8FlYtP2MJGDOS5vv4jMb4lAm+0crqn/57Al8UWYEtevivFkp+4jRUiVyoz1m7XBsA
4cZIuw8A7ducguSwiBKN0lofslNcNNbTy3JapOa0tjvCvZRh3STNx2DWRJZrki7Ypbpy8djmgIp3
l4V9L0DqdqyY1hfEiR0N0dTP2g1bAInIzy7JygM+erhvkVfEZ4tVUK0wbqvds5Lyk3XazwG6C+s7
77FZUoQ754g6Tz/M6pPJnfRsLz3pI+UoneZ2JjAKzrUx23jHuu3y8kEL/JTR0qc5wYkAzUzpYtW2
wRwfMDJWOi/K68orLLmorYEPNhXEMcRZJTzEIEWxz+jwtACB0LraZFvPxB8GpjlYO2L5J50cBP75
PPEIfycolmzNQLItLo4Enz96lgVOtdm9UIsbCa6Q7DG0OcrhJ8DgP+cOR21i3KT2guQ+F1XBetkU
aUOSN2oEQ/Zh2dznqhhxNh4M8hS1qIGTK1ynpujsWhjJFYFtPIR/2J6fkkwnfWaRXK5tcKtMSDBm
uckST/1cRua78Qw2qvxEKHOmpJSM3i8gOcb2kkckWEwLA6CX0PHnDg2tZvRaRDnib04KpRjbWHnn
VpkSi3mYo27KmYc75G4N3tKE5Hj/KNUAeWuF+A3GCjL/jkZmcAF677cH1yLxoHMiCLc5wHMXbZtG
JW+iEgA0/1kfpfZs5FiJ6stpVw7I/9ieBDy6H1aeoR+xNTGOQLPhTY/HAve8BVpUE49te2T3imE0
MJx8GcZoUxkgzJ1YhqVNKlJKciEtcL5XsxNvkydz7Dg6ytFz9JNDit/CfdbEeD86f/rBNgZA3stY
5RTcTYnBp6Vm7AXn0sWkEYbHtK9fg6ztJdxapQz48b9BP+qvuklpqDbVFb5absmSCVVMI8IF6Oxm
5usIE2aLPhw55lzUmHf8DyyKgc6fYm2AZ1UKa3WDIaZSbGnU4JqIPfZMwsIUX4Ex+jMFi1IukJ9g
V8WEpOrKCV26tu5I+RWl3OxncQkRPf9g78zu/m3p3epuW/mJD2BxDG5qsNg4MiIpAl4v9ysNU1h2
7wtlPAMyfOtJFOojnCsVAL7nIfl9oTajZSK55lDnDqW0hHXijoc1VHWz/CSDe9IBMEDV3LioVnEO
NhPqjkrdyEnInCxbbQ2N3yNwJP0x/EiQ7PWeGnY8njtMDfekLd4dqTlM/ni6KIUOd6xR2FbYW9TZ
uomraCKa1vLkF0QLbzyPBHKAEdE1vNGS7lg0qISxnd0F1iag/WH1jiyxESx80plQxbKBS8i4AJo/
n+JdkulKxndFh+o4/BPpMAtmBoYMgr4WXvdVFHOrIUUSndo+KT2+g3HUyFwAEf05RHk4IBHjgp2M
oOLr5qKYXFzxGYVHamn3WqoFf3sLh2eVFooMmXchnX2EBCVxehlXB0pyDYAAwR4yWYm53MMEtXko
33aHnJB50Ab2Vq77V6LiJgWH/d05LDtxuu499LwIefdJ3npYFCHO49TMGy89Pn8V2He84QrAZqm1
PEh7wHSsad8MRgd/8vq1S2zUUbr+cUXD6qLUDXwmAM1+soApOujQ7dgj9UBBukIG6/S763NqL+Mp
/z3vEAi/1mx7TKbB3e5zhQW9BTwijrWFNNDJlMBsp+LtSf48bQFi3jXXca/R1Ccz2E/DrDc9DkKt
cMYXMr71dW1oZ0fMXvId+lA6j4+DqbImX0ZZdXuj8D0OgeWPtrGYTiqUuYl9SEMwBUbMvYGHEulw
jDGozqAPy/6Eh2Ot+yNNZCqref97J2ZihaufMrEeFtejiQWRaOP0dreIF6lm/xw17rzbdbj3hFDn
4eaJXxS54XZbo9dvnc5TK6qBCVdTIzqmpaKvxv+qlS6e8ScKsT98BQyMmDLT7lw9C8nSpUOEgtGf
2R1w0VItavSjsJ2MtA3k8rtBzzufa4tR0nPnb9pKvlMo+MvlZAM89paTdyfWq5C8FRUz2qxbxVnl
gukzHnV2bTQT9OQNlZiW2CaOOFWvlC9Bnymobcjx8CFI6J11jMKAKRo7sHGP1kxb+5E4ncCZtU/w
dtSzmioJfdipD5lkwJgKhw/HK1lZ0S/fshfxt5zpDha7bJtMJRLsi0v49jSmqoGbDtkzL72qCdNj
CFOZgLl7YaQxmNnvSti6xT5WEIr4Gg9wlWI4fFHBzhJfbSvtziHwP0Skp6S5EHrJ9ow4bndFcjGq
VvK6XhH36FzZZFvilSTi8+EJJIIuxIIt+0s2h6YdfSwGq5MpGHIZBOBDntIMbdqTR5GYhNDM2DI6
nnJL57K6FV8daaBuk3wYm/UjH/+A+pk+4vtnyny+adpt3HH2ioYzRufbjrAwpfgkCzcJCH9JZuvf
PNOaZv9l5AhcZOcntTVUZYPHeeMJN90iWpZCqbJ5TejQzdko8MiAv43jRlIv0C8Ap+LubO8Nas6K
owjBSiHfcci4uFMEq1P3mjz8RWl6WTh8O5gyv7Uzyv3NLseWS0gOr9rcXk3Fp4ep/EGRHtSOftEi
Fjla3Nn2XSF3w6gHLsa2nc5k40Zvp7oY4z/yW87k+yopK3jizeQ+Zy32KDuXnX8NSf4zBmQlzN6v
y39XigbMvnqnBvM8CuhQ7KAw4kqBE5Jp4y5rg8+oMDX1Hgiz71Ms68G7+D1wZPf7Pp8oEr7kZ2Df
Ux5CSWz4OBbpXm/7/tX7LVO+ZWmw848hM26N/aLdF/Pv1Od7YITPvw6yNZl4UOEOMS3wzOMQy4iv
/EPPFPbsFY5B0HN0UIWwhYPWm8pbo9JNCQAJS8AaolK7Zx9MDjs0LrTigiMRZyV+hvTYU+Eqn6HX
kI77pHWLtWnx/suSN405fuea2Ts7jogCTzud5IdgswKqIiSycKAjUs/eIBIq5o2Uc+iL3ku7W1PA
GIGUqybDg76WzwM+59cD8O4LeyOxWSPZAS913ufTITQswsiPSOGGJvXiV2jQ4XKSaCyOFqaM/5SQ
3t1ExaFDy6p0U2eUDvmpxpnl5YpXfO+qyd4ROMhQHOYgzf33Vsb1lW5IzACJW1pQV/idmys3/c4T
Mr9G7q9BokyCewOpz59vdIxPSIWhwO/Zyno4pMbYKphJdk/3NH7xqjRu6sSmiQDR/bZWphDVA9gc
UtclhCExtRCjDrgKUgNy/ba57YzWMsAP646Droy6Y5uduVWkhbn9KtpYPbPdsc62vBsdvnbEqcyH
Nuk/1J4NPf/mIcRrRtB7je5tXLdRPfwGsapcOLnrkQGWdhEOkSQmXgvandkQ4Lu9kjk2x8MGsnxX
J1W8aN00wzbcuktsTcegNWfFLtq+YgbXJvUoCGkOq7DmQFtcuLkRlcvT6hlhFEDAjdA5iB9b/4ZE
t8XNSWsg5UNTXHsbeQC6ghjHjhJczbkmtCRlCH9PljeULHGt+YK/zqJGbm5wpV+cK9Zbuir4Ddgx
4ovVNaVEXAQGj9/0trpTrN51TjYRLCn/5JrHd3/jKF1oTCTTipM3rz7pKP8OWDXSCWC+4imQ672d
h47gqIg8TGu7w8We8PcisdJu4VDwp7o/n3F+o7YGvBiB1X22/Toe37ouCofkFJytoWYyR0W5zpXW
RYN8zfb7NXYpp2KEWq2WMwFNAGXWbfZBkZ76UDFsOonwoThjjrT8NTiTNkXXJ9m9dSGPeWZW8r1x
H7QjfXw6EWWl2snW+zYEld6AKvyB0dwcjyjZDfbrMNqqbOONeyx9p8xRBkhov5UpfADdbIAOqdtz
eSvyrkGmIAXv7e16o4hDEEh3UtV/tQj2oKuQbsHPby/mD0z3It3QKjsermM+4u7WdOFDETm0wnYi
kb5sNmsWlp5nfhO5D2gh1NDLRsmtXYUqoqdFR1l5SQZY3mxd/NjEZIAR+Cph5cPlWrfSFGgMrAn/
dd2nCTeLZbxgiQyn2bKaD4DwaD4qNsC3CPOtSNUY1P7Ts+a55gvH6noPfb5EHYHm4QD2TF79UpuF
x+XlO9nSrPZm6xJ7AFKZCwHFcMOR8VGDWe1tXTGxTlxXD8Xs2uzKfg8dglJTYnofaC+U3Xl1GQKX
W0zB9vJ4HwFY5drSWmENbjpFuRFJs+2+psEYyoShPxlyl2E09sa1Fo61SkQsejE1tjSk/7w4wUX5
uQGJBC3qv27h1BGAe9haq27db77jSwsyE9c+so5DTs8SfuCvrI9PaEVDUCt6HkeGq9dG4YIX+Mde
E1ZLp1NCIkPXDDsFpd4ebWInz/It4guiWFgVmUPoykaTgbLjKq9dfSIPzohaF3butBBhf9HBoBAf
fMeGXNtt9BAU/+jS6qHXCSjBNMUCVAMkvsJhOf1Bk6uTCPLyTbU66uZgAcaypDUHgm27wZbZ+b4z
r0XiGLhB/lLANHwpIaj9P/dXA4RY/dfKwhgr3mrBPUIb8Yrgb9MnwBwC5Wxm52lwhNeq1jYGpEfQ
l4lJC2KcwiRCxfqfQO84V+qkWJVojd8bpba26J2UtYDUBKYBb/uSp5V/vjjAsUXTZS8/83HAy7EB
qdi9hP3spHOiAF/r7U/2y5nqTbDFgRQ+DNuQ5M7Cs29Di44g/YNiv5L5OMioyuD+TK4ikl2RG6Wx
h4YxmsmrAgMlcPd8GfWj5R1K5qghvzFU0GUBQMRnyB7mmOgCzKoupYKVW/1sRSFeHevKD/MCU8W4
MVWNtszWoRXKc6Bj/wAsus2ODSUDgvOOt1GLKBbebDcMlZDdePYet2+TxHXEsEvKEL5P17qHswb/
FQfWYNfHx3C1LQJDDiip1WvPlEZ/0CNMeZQ7qWDCqIy3/40qWYCDt/A8NPfYuH/ABpCA07Nc33yd
0wil41jp4i0MTrWFDIn+FUQu7ku66fyWOGtoaJGb/8GNJJ4kmcov9uSQhW+w3ie1uMr+UcpaB0jR
185ZNZ2w/pWI+Xul/Vm3Vk3Pi2+3aVvwPks5WO18NzXzc2NIvh+2fmkvXMb5USTUzlPd0z3gYaUy
dmej4R5U6941kVsY0s2zwXaxuvxGaLf99jsrFGM6iv5Ga1gaVDaS0S/jlWCVP7UB+P/DK3EqjLsM
6QOTaoK3AwzlQt4pDI/lsCt+IVkri0yml5HtVKOa5yIt0saRSgZSZISUzX6YWyyb+4+CfpNqlmER
KR/iWlt2kQXBGhOYY9GYrcOIt6CU5EsfBimE+NmFsHx9nC1zd3t+sjjf67sVD/jgNgNsyj+ziwtN
Djm54hLxRdLSvkbFyLJEseE8DoJOGZ8xochFf34kk4eb5tg65ncTCeQEE/QYuxn3y6OHOFueBzly
9CDcsmGuHhK4j21lORw/ocxdZviXa01xy3IU0FHwPQSaz+wBgr7XZ9xJEVg/CFYpTrSv2yrV6z5r
bEVjOLIc82FEzX3p/ir7iaQ5jKZaoiZ3j09FQRHcphg5zeB7c/6txd0gmJxlVyIvSZeGVpiSt+kp
/PBzTY+jiPYjxCqZUpL9671nx/NNdbiElQSjp4sYlxDGv89xxGOb3lqMsMJxgLnVlqbfKRlzqbWD
6rwpfhSpr1WcVsgKmmdxXt+H3dB1ftTFCLunzrkI7K5ed5fbXepCcrkGpTTDlN0Q46wZwOJ3YM/D
YhWzDu+kFzE9cnQFwKj+FhCULX/Rqa2lmBwNVlWAnhPvG2sqZjK0HdJJLqUPBwtpqc5YOy/OdWfx
0hutDvN50cKz26N3o8TA7VRH2pm8I/Ivjmo09FRJHy5b5Z4Zr3L4X00I3wgzfkYk4JltODHLWjTQ
JO4xFhwRCm7EIZG+CTdzkRYE8CjFPloYL3HJCEkSxYp3or3KUDK5iDxXkWXnmeUb9+8HC276vGbh
F7+juDniV6R+UxZvkf3CNkkQG9Fnr99duFngxB26EmZrYqTf4ogrTPB2us8oTIsxdlpAtJmUl/PV
R4oxJpjtTdduo0q71SKzEOwlWfaXzm3jMwMK8771GUL1hQdrbxh8hI0GW48iutJZabhHTWra7kXu
Ojr7VwaXGE2+dOozF6a8KHJVCvsXKIzgOvWAC9strIXNUI0cgg612JxIwdpqe5kzetMuKIEITUtS
tlH53nB4ToOYY3l1nnL+klTmjT9pxLfNJV/Tfk9OaNA9Hj1jlLYRKhk9ZnxLdyQ/MTovXJpZaY8R
XVSGCs+qOFI4ROi8oqMtzAfb71E5gxzLqZoXmqm0tbGBDbJsKNDm85FBSXMhiToL1cPv8yjtP4ok
mo8ZKch+5ovXlXBObyphZ9nhPbDx+7EbSzugCeMM5+zZHqqytfcrySiuoOP+8qd4q10gpbDLd1v9
8l5v3qvtPIFX1ijC03GvhkoJ3jhKjCqbRpXQOB5Sm96hDYkEP5qXfzTP+1vFZqd1ncs6m79ebuQB
qC0gkZ488w3GhLLzL1R2vS2jex9QFFMuUXN83sowZLjrWe4JqmKD0GsWIFva69VOLEDLu1dIYsXy
Dwtd2RR1hIsrriM4yy4BCQv7K795hcjViTsTk4ElI+7wPYv7rdU+t3rMqi27rJTFRKaUbSV7BbMt
UwnuzDUhCKJLnEs0HlOg6CnZIBlsJ1v9IGruRL4x2QGceztiH81wXog1LU1zsn//EtQhvZMuiAtS
sV9zOeRaAZ2OGQ+zRf+hXtwLAhqfVbHwOBSeqbrWJrarqD0ApRL2MoNGmpqIKjO2sbeAOrQXs6d1
kziPp6BO7nv9CdOB6BxjP6BXW1GctkfTw3HPyb+YQWGJLFKzz/yFszDI7d0ZHZeeOAwDj9HWsKIL
aJkzyuWbH2qtdHnB5jsNiKAHb2lbyAdjCf5FFwuW2Hql7Oc+QZE6U9KvfALZCxOHIx1TB/mVyszq
YPxXSWvk4yPJEizT8akmgWUxGEzkry4Fgp/qWvClJHlcH8UsTxAUTny/jz8aAAWgekSG74k5mk4a
ox7CAKRSH07WqKlAZjcgOZA8pK0viFVfz3EUYwXw+WPWxpuOlrPxHp7LnQqGV0p5xm0zf5Hf1h8n
TfTlPxCsIAVKCgENOceUXUk7/g8+zkcsjx/LeqGcOmnX6mY+DxOMjOnZ21WZOk/wUwyo/KvSJleP
4ROGg5h4neXhJdboECHHkbIoZIWoyPi6s2eRgiEzAV919sdw6OfF12kSjrrRbuVgvWIH3vd088lD
BeW/TYMaJ3ePtQr4ZwfOioydDNmZyYsd+W+rz92F9mMU+is5o6zKdEIhlTWXd0/mTsbcRILg3Jk3
GCR42CFfaqtgq8d/dmAeddzC04RVux2aO0s57D/XNjiJEttu6jkFT8lsHxevppxL62Wucl88L6/X
GN8XFDAUKYn8TYj+l/v5DFFgRYsKhL2esyeaEZR9nwzCzOe6guTSq4g6TnPU/7yrFz3morgIFSMw
PiRFU5y4IzGC3Z3ztwJKLFSK70HkJCOO8UwesXv3Ocnvb94i9wByCxhW89mirP3+pJh8KdKuGEkL
vDItkJrjKoX/GZurlGZv4wBkOx9bRwLyo+SD/G1SAk1Yj8XlJt7YVfCh/lj/ssgxryDrWLt0soFD
JAe6HjNoxhchJMerzhQqrB36pYm6No+4+3FaP1TQLUOHyORFw4h2MMVLBerZNtWF4AQdM/IQt0+t
pRbAtEpMIKOIVqE/N4PR9tWRztwY95uN2+GiWAC9aDb2BDr4LudkNyg3Xn4E6ZjYkqJuUHnA7B2u
rW7x0RW5qN4e4jq8cc+bU6lLld/jrvIIcGsXGZppLhsNyn44226bAbUNx15PbYZZ6h8h4StsySda
Ly9JfDzQlI63aXd8RmpLOEIK+hLkHrJ4M4swq3M0kyb2LhRLfYrA9Z/5z8GQmm2odPxhUKlHQzHR
oUAkrKeWdZ+qIDMDDS8HauZ9zVIxTtp0JzlureH/YGqtM0XeZUhIPwYR58QpGQucOoxLBCInpkXy
13WfCr55dZyF9FclViMq8abYCPjlBGTcq5uVvxEp1zOtdZeLj0pvgLkqTJpiP3MWJtvp3z+LfeMK
tvsbKnw7YqovcknBoSjEIzoQuts44cfXop8dZf5XE5PDjk7KOn6Ts0Wpg8BhIfrpvhn+ZNV2CDiD
fGtaBoB9qwTQJWe/pJDGoOKQNvuuV8dryDXwbfrKCfy1oPZl9nQPOBTQP84x7QY+/KwRFQbtghlC
+gpSuQhv7NJ8UFzdUilLc702LGp7oV1RW8KRYF/DE/zsqVJ2BnF7s40nnNyTgkthCLReIz85YzoO
Hhc/PZFA6lrNOACWh59jAKb4s/CMsA4xYw1ASLRZ9EgkfMDgUw4shICaNER87yu7nlmRq4yx3qPb
JpWmMr7dPhhuNIlyHcpglLuz0sYTT562foGx4nhcZuw75P6vkjf52mWX+2hCZGpCiguX7+0m903P
Hkw1KqqFMjHuTrPie4Xqo/5ojffgExN+d6EZQQn1mmmN77XOepwtKpgaYaGWr9CWmm7BzTmB3VDq
gkmHiNqGG2AvT7XFlsMaqKKd2++Lr54WK+4JYMk5fafwAZFbQLEfJkBvZmJDIEEu++6mtVEyhRcK
ljZuu7n9oUUiDwg51h4Jj3RXoj2nWZovgsgx8taw6LD3WcRlpHKKHgNzCgQutOl/0oXjQhO4Ucem
3RVg2dqp5QOxBganl4fvphG3HL8CVapgyAH6CoH96d9tgqYNvH/Hc0g0BEVFlivwZDIJtC9HcP6a
RLMfCL6gEVAzJLVc6IHnHUhDv5uYsjxNlpaEDc6ds31d6CXpaRulpFSc5c55a0gyVEJeoNBXxZFp
krpaBF+bpbzqc7FMusgzS4MFnh+QPwNQtBvBlQ5pEKwl3UfvDBgoAias/f13/N+Kqge3OxOwbeTr
Waghmt8ldBAfMZtzijwXeq3Wav4x95ayp41SuCWhUTQDZDD6sfGdLE7E65hXy6XmCqLdsLe0DObz
wO7r2sAKLamHkWTYKdACHxa52fFFWb7QAFaj8RBjQB/4QS64g6w2xVl00Hc+03ilG0GlegdNEcdF
fru5NQgLgZxVp2KybZwzffLyea34II+ihF2HtngF6hi06iKCm57TwV1kOsqyaoxMITbUnyrLyBKE
6CBRNbqMuAoG1o0GD2X5KMyiMb3UELQ1z4eNHZ5gpPOg+xrACkA49dk5a2w02LQDthLQwPd/Ct2u
tCMjJpqdvUQnf1wvcMggiXAeOyciZxKoanlEwPTu4BeylSrNecv/AkEwoWFQ6zFjyzrdn2WYnr94
3faHEM/UTGnv9p+0TkypCA/Qlx6TWeCItdVmHv9BRSiRoffCm0MTcvdukDH+kPQoMkDpM95wHJar
9hVyfvoF/4DTslhot9nNGVhFC7MZJGs2Knn3p+4ld3sPVg/Wq2h4U+SF0vLnWARfhYKNqfrdk0T0
0LCfrW9CPp6XWDFQXltDTo6wXwas5A0zXydEiER5BDEt8eH/jLs7RXK9Xoyeq68uWbYV+5Y4utqZ
mnlTTip/VKdtTPBd43aICAhUzQh9M2RSa4iiXOMdyeZ0xK3kLYKru653WLHvtZsjsQ0ot/YjTvLH
PJThIFk7a6SCFHDgZFn3Lv4HVrAm+yKOTVQIQ1CY+xCHEd1EgJ9HVJio1dwKUgM4Fw4rIXxTKmIr
f19cUc7LPxaLd0bLi4sC+zoEu5J8ubQgu3VhvvVi7R4JsXJt1+FJhbEWgn5hyysRSwz/CA3lef0G
J8Let7rldIbg9Wpqr/xsszW6mplBk4rvrA6bCdAshyRXyClDPYuQLj8wqRj9l1bkYO8xePKsg7CT
QrTy1+oonCxnZjjl2jiVilXKpfdVLawShn3kzQlkS7nbWp8jKhRK/+BDq1K3imCtimZISlWuYLey
+y1jR4cyXtH0t/HrCrU+eFcgxY2qPEorpo5RJREbzcfkBIpBhFHMF4cIZX/jjBZZLpkNTLPc+HS0
HBnPChIWDMwxYErndK2A6Exmzz+65hxpmoRCywACb/O0q6R0rvXd0LfXvi+CaJZd0YV7pwh+uMYT
dN1Od9ZJLEmDELmEHTGGScG8j4HOVDfRH41qyjGU+ilPSOyZtse36EMB0Jf1Tg4MghnuY9d4s6ad
igKZSX6+sEyUMp0BmillTQ0oUrAcREz3xOgGO7TK3csyvZopAfWRw00xpz47CewfAuClPczJ8h4Y
w0A967dSA3ihVQO5ZdiNAG0qGg4A2g389w9ZtrO5kJdJ4RjlmaRQwMeRjoGvPs5Vy2eqZBnhnWGw
xkGy7+2XQpTnARRG1QKHO9ry6pCN+PjnyXEIGGF/1agUXs3fJKSCDHSYarVy+WF9GTyi0N9xt8a9
2nENk7apGNLsmF6r370+Qpm0yO6eCmRZ4l2stVPhSQSgH/7PyaooO+g+234kKwbyoD4nbX+ivx8B
xn99rDiRS8onKYEM2iOR/vXIgFGv/CoMEtt0znTYKgJ0FxwUBQuxZ2NlkA+1QvBKbv81wFv0/JD9
CWkmpRcdJklgPiiRUnmLu36u60Gg6cEjIdIG5J1a7l+IZpUERFUR0D7JhO6bf+c36ueJP9HJKu/v
oZCj4hBJ+Kv5KOCt29DLHgdGZfP/gsTZMvIbk/B29rnT0rvdp2e9BdYnIevT4U909qxgQD5EARuj
Iyl/+Uztw3kvJp4EqDI+CUP4N2ROW6gsV8kOmaQ2gE8LTTn7T5KqYA4yfcCW7Ht20UslFY8K6EdK
39WKmCV9eVgQHCj4sTmDzGZyM4FaW1eVggsxwQpoehUq2x+qheoJb4UTdESK9vblBataGzz+qUIm
ePseWlS9joaMRdtV4mv0LlXrUtXwNzpHG88QjCU9UjAwKFd8vQDkUyAKYWxKrB2AL1HfSRYeZHT2
R4imfUR3zuvURnKVqvE8Z/oGBpSe6BfsHuNnV+Svwc65Gm3AiM37bhkLeRRFpwcsNH8Leg4W0khT
TtVpUIz+nuE4+3QuZr3dKR9UqBIkOdOdg6jAoosEcNbFfrAdkBIX93FsjyyMuofGenSfcJTCELNo
TsEiqGMZShkGyLq7n6kp2uEUGvKADwTZnERwqHJ6GdfoF29nBK5pRuL4TDcdtl9dPGVd4fR9/nEK
v8/fWeTjdYI3plPrQQL3U+nnZDIRm5C1dRJfAVwmMb+PZELTisQWjS+sJm5cm+L5rUHmhR0rrsbp
Ntv5ZkISwailIhsx0b86Ih8UgIHPgdS8tSCV2Tjflu55YgmWozQGIuc5Ciy7DdekeiHKaRLXdYNE
3B7mQ0lIeQPKLzTuVit8He7HGtjCQ+wJZrgpIOKwFQj1dOwgYxvvBWU3dK6t7Cv8+G5NIRfVb+GN
pLVS+1lNJOcVzFDxernd+66T3rmK5/xeNYt7bt1CQ/wHj4oGmzEuO30k+MT3kw2Fdl51iotAKZxr
rwC8w1zlHaQxEbsgQZP++XvsUAwebH1rcxHo2CWYkq/BEhbgRsVPLmeprOMGemMsIBDCFI5voEO9
G4yr+tLGIGnvbCn0hdBRae0+rIpQ2F40dpslSyPSX00zRDgC0iAlcVFu7+4pt420XS0toSvY2Tak
tYFFtwiaw6nJDP1zrxmGsxHis9wB2QR+ffP6zw3bzqQ5FuDDBLYdB4s8fLnTcFFRfNcoKFCcRS5X
aM0Q+/cgrc2oOMT2q7fkJfOTJ+e+UaQNNZ1ICgN2dF/Z++cVffTWKrtCqZIQuj1hkfA6C0HpYxmd
unhKU8PxTeD9EVBfb0R+WwZXA/cuw9QjuwwCiV/7HSBacqAYONiScMBlv0Qg6A2zJ/ouT5u4WBrz
Yq037HAZVc+Vv+6Gbv0DiykkbJLdk0OvZkFkolyrWkM3T+xSwSu/wrXUBsM7IoyBzF7q1CyLzLip
Q4f8MdTMIY5GoI8+wY+JGDLKNculyrRHUoGBGvHoRrMwxmKFQs9lw0+/K+ZjUUP1+lZ10vd79KBK
D0bJmzV3qCcJjxx0j3wMaf7aChJRxg8klplmN2ByREmEUr+luz7jSvnFDW4moQP7qzNMSyZVWeTG
dnfqH/Sr4tH+enfF5ys5MSktDo7V08yn/28a5nDmOR25TncOfGzNt7KcW3N7XpxdtuuaqDKjxBpf
RMyzYTDVvI13fJNVLSNbtYNNnIThcpcg9K1eZF1zfb72wphKH50DCJxff8rmlGITo3Bx004wq06X
pI4lreM0xf96Oec7XMK2A+EQB0oTTkldRi+bgxAYeT/gE12xy1BxdPcKvjW41FCp8Oj4pGsBrNQ6
TWV9VpqlGTfD384NjeX5QX9tjyb2A5dguCWgMA3pBGK5yhx+DKJ8dcALt1Ym+ZGLfinJOJI84OJp
QVjGq0bw/vsM5KZF5CgjVy3vjw6wWl/UbD8BrAPpdoCapuF35DjpNRvKrL3P2EFx78Qa/WGJoeWe
oqwuMh1LnNx8/6T6rwO26uMTguprqefoXuDDaXE704cW4PJgWHZRhcw7U+7a4yokxFrdDKcSdW0i
UkOP5ikWIRVArVNQudgSxQMQLq7VLzV97Mgs83a/UOEE3fwAWSMDkMvN8HM2VV4WgdqbNypaQZ1s
pNazPjWBq/IHmbc+kITDdSHm2c7hUexB4zKIxIZx6O4OVcJzNZ8qO20AIYLwlHiE0v6hILAYb+Xu
nPWlLVOqQXcv1S7Dv6GS1zL7BsH+miNG07LK39VErfxj719tzPSW8r7grbrRo2vjJvJhEwYbpHCX
s8D+GuI6Ct2h44JBsd33mgiooQ5Pm9DVjYMmcfGuV4J0dlCHXxXjrM24M1bKAdCdB9nz1KmMxke+
P8WOdei+5Ckp780caiVztvAPsMXll+3KHTG5Zz2qEC2vkiS9PfuTKIRalBYvlJU22FHzcBE6awh6
iBbIIEQCTN+4OWM+rIWEobDLjoXDkkw918QDFoqLnyv0LV868ygDnEgGPiDGXhwRvIwaKj0S2gIo
Cld7iqFKI5ZRjPwcsF8oB/muMFg4emzgeVxg13OsoB8x+Tq+/2InhfL/CUTs7obF8uxfzsgP/kxg
jSu4xyPikOwHj9IPB7alpekzv54nGH3kG5aoZ5CTW6K0t+MDNRayCU2RInWEzBDWVfG39SUmUmuw
jnWXpwleTQWqF3pX5hIjIAKgBZxZSckKvDdP9bArQz/HneZs0EqVEGliefImiHxNLPA9FBeH8+hv
gF4WwPQ8umVIcE1vCkT6MF4jVNKKlKCBjIxso+a/b11hZtjIshUO5ElS3WIIizZKfRWuS9RaMm2x
bx2uUNlq8mkiG6nhPmebxC1AmP49Y6iq683WImXmC1YT1pkL7nnc0ceisTJrr8tmSHE5Oua1LzPR
24mLkO213bxc7l3qUBCZQDkdrqF1kXM9Lgt++2uV42CB8OH+qysSe7Aikjzt/0ANg1funcf/xzvx
EJI81cLlAGpy10NImu1/yjSIZ1qlSyCcrL/sQTlNUC/QKZLAZh+cT++SMCp2xw/jZI/LXcHKHyDC
JnqD75BX2VifHM6XweGiVC4ftb2uzynsrp+7YbeFOK1x0uGqjcf5z7F1n9U8OLdKbNxIi/PNpnxU
oVxD6qlTTdga7z0dAxTj1d/p/F4DvCjT/4AE0qcK28YMs+Jz6c3zg/ObyN6vxC34gTirLpTgzOLS
a5McGNkQ+JpKNhD/MjBAJsQiHeF+Bhc2g/cL257cC1nNHkAsNjc6k7mr9zQjWjU4/HQ9X+TB8Lcy
KoPe7LbroAPsw1rmoDnsj0fHfoDRMeC9UWyTX65bTiRgf8C/Mr4dNu3loJR0eE8nHQMF7O6Swt4q
OJHP8+UEPeIj8FaIytKB4Y8tiiPTjfAipJKbB6M7GQGv79y54rE6cujkeECL3Pjtl+To9/16M9nA
1id1tfTsTrAMyv7BLlrDCn3+x7d1zFPi8aNOX00jDL/cdMRFPjHW7xXkm4d5FcmPcermg9UDlu9s
gVLzodDBIuh3au2rDyc/LRSBSUoxxO/4d/pojn4FeujxagZ+M+8OEzj1FoJUhKhTtesuKMDaXQ01
hhPaBj0SV4zF7FomLzcmRpe/04pfYaEFFNv8kG8fyhA91ikUgMeN4U5Yt9xqCGXJSM08wjCkyCaC
N5vkHReNYNF4dkfWvKp570RlCJf97peWEurj/HBD3xe7KJ6MIprK5vljigFm6DOJvaiPKN9hFOAF
DAJDPu3TyOvZHFnpzTTzMBFsGRz3om5YY7lKwcfzpaJSwcJdZ5cSXcfSOHROg9epXXMc7D4C6mZw
Mir2a6qwQdXtvh9D5x1M2iW/13yad/e3ssISuEjCj+bXNCU1cE/VmDbYTp9uVKoP/m37om0GJBEE
hf5yRHug65b8qxeVkcFedDH5Ncat3oUx8DbGndVkyIzbH+6jNmpcUm/j5FQjHb5DMjhtLFjzyW7f
1/gUcX9dSl9BhdnWNADuPv395TTuxcE/0zFELEcPnh1Nv2jDX4ppRTOORM9FwaXilBl7Dj7Ir2xa
Xce+HALnbYj/QZPaTkFBBhzbbI1t958m0jJkYPidkXfVOWNVNjhxJNMIbAqxyJr5aF4oN9qA/0bd
Dn5d99GSyC354SenCdQRseCCHnRbIJFieaBWGHkizMyWpH2HGfsIAx2HyGD1SZH29Z51i+MbOgV4
PW89vTfZMBxO+/PJWXnHtUXLrCaZdc8ARJQ8C48n+5HsuwhpJrHwsVYoRAcAGTPJYCT+t5vpgtjc
217LliK9ooJPaWB9U151zCP1OQswreqjNpi/BVjb07LUNbNlVNXk0EdzBXILC0Re1hFl2zlI4rWz
kryorqhtTS7UHYZiZbTQiX7/C2/G4m6mc2HNgoPrzdROkM545wctnoGTAg72uf7GJOPHOtaPmekM
ookkeGdSSM15EeoEv/tnmSTrpvGjjSINFCNgTCmqBPikJIo2JD6dhtJCTh+bvyRlLRwKhGWEhUhW
0oIdXS6S2miupRu7kLpVcghFvGGrLfrphx/delmFF/pZaZZNSFDUzb40FgWaPo28z/TcOjeXeP3n
/BZcLTgej/qmWLFgcouCfWhdU07OsZSqe/0XoK/xVpo696oSQTC35gZFNa0kcp45kZY6oiboXExU
rJzeuK/9A9dz8rlmf52E6vn91PR/9/d71/HL56hzawfFhCNF7Mu4cHaKHVZdsLbcmjsNR1aisj/9
S4TV/Pjuay5VhFPAvf+7IgxdlgyS8X9RWsWmrbgENAjTaavaAwmGC7vlf73p0MtlbuzBmtfR+A4o
KtA5urAlR5oBW+RuL10OeOxOdgQYXY1OMovBghtiqUzc484xzKCY7OGH5Haq2iklhU3QCAoXv1v1
8EUhoYgePvalx3Obnhp9ANZLUhgz7cc5ZGuBSkgx07vRm/vttA8gQZ+x6fuNU6wZJi2gMX5kwry7
2jD4L0iic6deUo7DV0+2tz1YOD2ND5mIbMco36zzRYtRFXdGN++ueUt0bA/nxTbKldZrR8QURdjD
DNOPQNDYmgrVqw9aX/vnd/v5sf2QO3RAa1Iqdy+T4RHdmZS7skBoc5mPoHz8UhIYKA3R/GBnSl01
axAeFlmUybVHhUa062CosrjWXJClvvDbfB+VIG+rJshpr68aJeLBL9ykNMgcNSER+nByw6zOEVXv
cQoWWn8lAhmYmjbZFjNG8zL4nRvkUkum7fU51sMG+95/AndopNbr6jZgLtZkMLfgr9lrSjeuDE84
6pkUgICudHi99jTwJb6E5CrtL9WtK7LeReZTi3jpfYTq7/4AQN5dNoc6aM/tsZ40PfhZEiHlicbK
/k4YSOsYyZ/nh/442z8bmHOOUh3dMmwrSKL0gmaFCxrI6EGV8M7fDc9O8BmI5+qpF2Cu1LN7ikxa
WepduW71eK2diBLI8czuVGDbZNOUYZHA8/vZa6u2LaLxJ7xtUWsHKtFT6g97os+KDlhB14L5Y3QU
+8jPelyFKcHv46wROcnfNTwKrL+47/2lJyKD3DWAdMi+fLCwEerlsCNLChooHuZnn9u2/Kc1EtlW
lxk5INOh/Zje0y1Q16EKiHdhFPKm/zrbe7GQiahoHCJNwmKmFNpHCm6Uw7SBKFxceJUtTYF6n8Qb
Hogr6hZ93FRBopKEOlJunCWSaQrkK5xrFduMGlhne2jEMmklBz+L+kNxR5GnJ/oT0QPriVEO4MII
SH3jvgPpLumgka4xErmSLb2cGqpivD1zQ5et2z3tMRkTVP5QM8r4BZPQVTNQ6bBH7bcKajJ8rDY3
cIycR9vptj679RC262eq/eQfRh7Q7GxiqtfubP48cnqY5zg+EinCLxQwr9Ust5pqr1RmP6z7mDEq
cIBMWdtSbzLSnuIchH6g40HA0YQfFyGh1RnMUYL2mIWmlLERxYxTFgby9XUnWYS2iBpcq4MHMtOK
/MBHC/5BmG1mxfyX8bdcMlpyKNtEG22qWz9W4ZnVdZo2PMssI2/hHbZrslCH/6i5/FelutyZwz5i
BFZf3RAJVh2HeBDHqlyjdolZggyCAWryMIzmqAsB9FAj18PGlDgrfQC888ZsSP6KmFAFWeb//qqy
lcMEvVroucfpbjH7XIw/ej10GRMYUedB/nCmob+o4PD21WUGGQ4jKIYNN/s5RQPs4eJnaWtPyDbR
/pUHCASJAfm8YiF8aZ4Yr/gBfKQpZbD1prGdLwyQ150eVvFCtTPRZNMMQvP1NSUlYHUhKLAAPRdW
N7DVjG92u65xdjeL31szav3+UEMWWeprNOAJHzhDZvqsbIpSIMbQUbfAI/BBf5uMZOL+B6AEbpdq
ausIilA+WsymNWzDIi7FsC/RoPZflXxvk5ijKe+Q3rWV3tSm446vsmrjfNUwTCt8aS553NXZAsM1
x3nFbjNY1+TeiPKh5fcxtiXINr1kg5/bZeDeMW71/01idd23rYLehOlu4JOOIHdUmPGCsKRiyasV
p2RJS3YLnFKwaIUuU/rySjMfglDz+4colOWAjKKNL4n2h3i+iObcIxNQAoRLuu4zrJp5YaFUQIPM
QGoyPeAKRjW/tnhpZkR5YReVpKpIw2aRczh80UKQqGv4tck0oPRWpXy13kahgJ9I9jv7BBFGzpfY
Nr1g6jCU06015LdhZqXDn4QsPFetb0k6j/LetGwk2Vi7MeHgxBYoF36f+0WshIK85I2p7doB0sMS
BDzT0I+yk5/epHcuhltkw95oNWG9qsOl7Un1oyZKaK0nsli+JMzsntupq1smbXm40xv1HbvEq/Os
d/VmhGlSPBA6d9lK3mJeUyEm0PZPjqJu1JsKCkqgx6TVGpQ41EEMEcOhhIFkYy/0FT0AXM9lOZEK
eR69IbJzoxFMQgV1NdCh1WwIT8cwl5dZzUjx2WnMs+4FMW8uYwdikrJKmkIlTU7z6t1nt7DaMqzR
xeVdVa4fbSer86wIYpn7IWcnGP3Z8eVBLHDdd46tvXJzS15IGpXHgISv7+NLXHWWLTsZanN6YW2p
qQK9r9ESaxGvsf+4f2g5vN+ulNWJbyCCsN2qJN2i7sa0cwBELgCTSegU2g0fCQW83YtHwsMsC+4X
2fP7vufasj51RBt718hMEbNn61a2uL52C4I1Gr2TOSJJ1J9ML+cmlGE+6rG2hFuIJmunmEDqD7EY
NQ2El2p2LqpDvcUCP+H3M8jI6W6aCDGlf743blKMFsbvxtLXtccxxoRK8tS8agL7DlL/X+j3RbgN
d7LZhMDb0qQ738VW8kJMNnUgqcJa9f12hl2NtWJGP+u8nATmNetrNn1x3HI+3D8uJGOmyJ6gmje/
iv+XVV8IL4Xon7JRVb0QvaU1GlNjdyWRD8CJB4o/O9cm+OR/lZSGP16Vzg9WUxEzVc21c1NZaMdr
qg37sOkyJKdNSo/XzmNJupnbKKZBf24ptTJdpuNCQTzs+NqAMVnINJXGYYWkENvoxa6i8Kw6vCl2
cDfQTFXVmZEktHeRAPNXW3VSBow6mUXWz9rntvF6iG8+8HbSaMqAkPPzBi8vn3btyPV9lOTLVZ55
jOTLw7hFwoLXVXwB+8y14QZXJX0RFkPhgRGf5nh7mS6gp7MvBrfSUMizx43DCiFsZQSZ+/7rF/hg
xCgNCvMB4xlNf6rB5WT/UAEUtTi1R+QD39A/ZidpP4dcm2vOaWWSRKkOkycauhDYFwsg2H9xgyJe
cAu8CrFSv7BD8Mg45bMCfjueIfSdgjRv8ATAkzLO51DMhVCKYu0kkPAhHKKwlgs40JY6sLDSkil/
MTa3SjQ8wIEfKh+A7/WVzBTT44RomZ8Z4RNJUxJBsaCKxQCiNNK/L5ikSB85DF1VE51IchrCLTHY
4RdlpVbcli8aQTQ9IHg6D/PZRYN7WizYzKUPSic6GtM+3+E3OnkSwmY9sGsakG+WvZcQ9D8XMFt4
YDzYnLmljX0M2sKe/BuzSwX3HAtiJgSm6Fvb85nPJPH64OQ6UuL89c5T5wvfjHVonyBYaPMfus7L
ckEZOzr5zQvRTy+IW+s+UVRzCR1p29vQX9v63b6kibpCluZcTEGpagXBnlNA/fRnPCIHF/PfqMZ7
e5As2m60YnPE06r+X8+9RcJXcf/Wg7qeTl0IEwAvpY9BKG7u3i7RVyTiITZ88wdwcNHavHUhsaaG
n6+hvVBd8hL5htCF0RiHJD0pC4x0afh9aqLnDBePGJiAPCr8K9+B8tXzZxqHRa4TaY7Or6ypK6XQ
W/DlHlYqjEbdC+w3wxWkTJOwRLR+5DX4wNlgzTAkg/bdkTYiKgxzYCB6AN1PNc7jEuzvcZqJ5h4X
nzL/ib8NsFaGEKzlCTJNnAZN3t9EuUiQ6GBFwjJDOTxJhiVJBzJkJNjyJbVQYhvgIZX1cNfUnxBi
dexqZrM3mroq49WvzXr/svK/kHIOx8THJBF6sgEPDRs4GFyOT1riyYenmORa6jz0MdJaf9iXnvnA
7UyXZv7w3/VYgSTf4q5fO0YlWquz34D+b89Hz/FJqrE/lBQjABVVz19o00T4RFMgLv2nTRcnRjcL
DcNxE5xqR66tWEfnU3swEETXpDuXKbVvA38m56E7bS2N4JHm7lA9eowgKbt3CMfLflVYj1H5fuw6
neGG/UUuRDx28eLV/iyIL3LSN8gkEjpv1sO41OYEswR5JE0VUX1tyCnh99m4+NbwFn8/hXShAVlt
xd1Eal/L/nSKLIkFFe30UcU4jy02DRt//Ki93g+OjgGHaVJ8sabGnznCASmBtSal+dfna0YXc8Pb
OQezr7QTYw54ST9NSFtFoSIclSSEH1zfOLmBt7ZwygUkhNxhbrxO696nZ2VgMfbsKIGrR4eLQBos
9dXzZ/4n292LApWNdzBod1W5y1/u4vkNsTqTfDyFuh8vgi8WLjEiUFUzDaoXc6480z0GCMbsDyKt
A3dfA2slCNtA1Q0nsubf+ime6m2mSD4006imMPFowuCvD4vKFwTGOQovMlUjj/Z9sVYA9p9FvtMy
uPO76hA44G90O/+USSIv8TOdFaSlqrFRAZuSBBQrLoaJ7Wft2SegqQEhkZpRLvvpyhoN2qhRg1rs
Ns0B5UM24JsVqfwiYhs3IKXyAn6GD3Lfl4vz1Ys+gxoDMwUg/rWtdqIMtJtQewjN1lpe/WiwEM1S
STAZ6YqWiuho8G7UWuH1+sdm2xpHS6qh03PlntAGpDIGagYCZtgQ/s/B3ZjOEkePbr2XwrZlgqwI
++fXcv0gcuThg9jalWfwChicYhSKjmqRhBm9YVdrfpMuo2+E03UvVJ99VXwGR0XoIqE56j6bFz8T
uwLmUbQUYItNk7bQRcuBwHr/LZXXrsmQIwUTEpx+tXUIaIdbxzgKShV2FQx6hf70S2KCFKmH8fzm
d+5FVsRRphV+0O9ysG2V9hQsz+s0hY/VZgiSu9+9RiLbRUNn9rfBThrbSX4z+z+PdAgrywQwwpts
8bpHU4rLWd++XKITjnzR0eJogEY/fyn8uqVy8Br/YboiSqJKGV/+ZuPfsXu7bLcDe3Izka6Dpurw
E61Mx8axNoC/zNk3VLqfFVmbIV5xd4Aug9V0PUUEkfmoZFCW5Z7m1IUWPuplyjObO7Ysmv0BJ2U7
2CtInYsCwvVVxNCodhILwDCLnX+DGV0S5zIkFPTw8g63+2rkFksE8vls5ysAklxbkCYnaYnVlT3D
IenqJQB4OBfXs0HtQhD8as1YAKwVEuK6miTWzVv2w699KuOgECTt72rlSZg+Jq3L4ZOT/klfBdo6
Ww0IfahzqDGk9Z+7+e7QkeJKRiA+9rNgN0cA/Af+Jeu7sfHVXx597QNY52rrMhdREQTsoscAL7l+
qIc9xGcWi0t+pTUuhu1rRrwogCso3aMRTOA+VUPtPjh66RtSWU+0pHoanb+V0Mk+kwCYuCWslyPw
R1Tr/j+HMUI5kfh0Sfzy6XoArzKf1CBd6f346aMyHQKRu3WahjsVUeB0AXm8LptQwx7NKamSojSM
iNf3NfLQs46qz7D9j1wcoCmvxdisGhJ2xhNBZU8vADHAjC74naAbNxjJcmFtS5JdTkeoguUfPwST
MY0xj7hGzquvHeOZRlnUgfrhurpQ0/4wdXhzqn9bCUNMDA/tK9aQ2DBYH7XjFcbOYAOrsbplk7ej
Lxq02wc/TLQLdnOyjqn1M2uGbSP36EJe1Y4nldj+CIOIKH7uxWMyMe8InMunadRI79yhOVJgzU92
+TSDdaxkrfnb33A1PfYivTuQ/5rOubaqQjV0qP21eETGtDo4r7EBdIi8R9x1dnJmX+QOBWuxwZFR
tsV8x64QUM04jH+I/C1Wm0HOvMAT+OPOjz3+iBtyXI0ff1sRlmWwuY4cConPFKmyUsio+JCm0XQI
T7xK7M2GjokvMaowlqm7Zmp5o5zt1dZHdgeQuuUibr4gT9u8+4dG8t4Bs6YOC0LnBvIzs3mM55bC
OIlCBy2psJiNxQJwBd+xuXHpqUk+tEm+sYPXvWTZKYJSgvISeYj6riTEDitpeCjnO3GMUzawOWS6
ZCVnkLl74DKh2SJj+WQQ5Bnoz0CPkN2xtAFssb7c3tufUdt0OtVuEtAVMadvbIUfFPjNiAldUq+H
FuSbHS2Vgp1TC5W384IdJQDgOGTHvf3nPEV8ykHDDGVzdvVSrhOqQGAv8STmKh/TBEq9HLhxcvX6
UT3h39BwqxGBku8H8r05GBR43sD6ZQ+REgiVqn2kTRepqE66chtOGgi6nSfPE0Vy+hN5m8tVnIuh
cFQ811VGkkhxgGmNNNdTNravFiRalAT6rpcnmgTihdxTh1UWGlaUDDZldF8B7hjVLcn7a1gONU93
aGl9YNHCkBPf8P07Ni8jCkaisCeTtpGACLpegDiphaRtbAtgj1soM3h8XV9hjiLwco00/l29/Bq0
Dw1wAWYsqZrGpyRfabQroKmO9DujtzIJ/Bh+/msU4FMWlVG1PAIN97mHcazoH66CuJ4EpgbS2x6P
ICXOyeXqKmggzuSLdRmri0kTjwi5PAdyFdAqhHuWXFEhH68OTro+PFGQ2mF32HUljgt9Y+CfrBFk
o7ZgA6q/z/SGOqTdXhR0MxwR2qoxUgEafv0enDd8jBe/3lK5sz33t8kGaAVRxbWw6VuS8t2HUHF4
flCD/2vAyoAvq+qe1ti5lyrxJ1Tz1xVfQBuWxF26V+/YqatkzJ7oJMLhiueu0FH2H6ZdIZo85FKd
KDd79AJkf9oTbU8zPbLsq+12vDZb79li6Ce6YlgPJon7gL9+MaQLDQoLI/ke4iAGRXoRxngQFYpn
LAzONukYgoXgZkafkwKTm3oNjKwujEJ5V/ZY0hyfa+0XKYwkbxR3F8umGyQLhj2/Zt/D7pXG0SY/
VGI9HGD4FxHwJtcET+aqfMaV/CXSAxinhyZD3GfgAZxRmH+/vnrVoqxCvOIwjVsJPyZNvyuHhv1e
Tw3hJP9N+EIrJ6OmqhIm5FC3ODha2Hog9637XGrmKGCMfLHA+QsaC5pTssKbUtit/dtRoEXuUDcn
4+ewqdjf2FKxkDiRFw0QWMleF41AYH2YDs1CuETTAQZvr+K+EtTdlKWylIOza27eit+nyPkO4s3E
0+qvXywoVoHClZQJu8eTiUeAl/kPZADj6iMhZKD4GUVo1mqAlGc2sWTnZOXJGmMmBM+XklOK+Yop
Wibv9lSXcOzjacOGLxWtR/vDoXXqkEisAYaFfcCyjJ3kP4ULpratkTe3zZHRbPOzWsW55FsKA8Z2
heruvxNl2PVqAQgRwxCHU8Nw/rmGSZm5/C28+lTQsucTdRpDHpOjp+x1Mi7ginLP1kFM8mheICc7
jJVdav80/jr1LCowA7GNAb8Ejl1uh+aiDyrj1jMOQPhaIRUe5AbQUQg3Z5/LpiuuuBPHfX6X8rua
YmqgCoG1FUos1zBiodNPMtnH3JawvUsMkT8pxAjJamvPX3kUBB7vFrNzTF6nuctdXGM+b/gpC6Po
v1FQq43jDM8+EuUGUQ2TAoI8X0BW0IWAZk3Efl4Qst5BzyySEnajlrXLmaduKmT9c1e4ghBh5Wtf
4Kp+C73DHiR8Fm3UvIqdytNX8cKsUpZCqFk4AcZLnjPO8KXvYi8Q2fJvaU2AlQ5bxqPq9DgS6Kny
lqiODQjBDoMkbkRPZTFwK4gvi0figHD/tMftF9KwHSlftlfl3AkiFykJAygXdnk8hOeaWP8UXOhi
LmLPe2YQ1bAYjNMUz1h35kFG9iHk+JAvwZAYl8qBhtj6UxgQlyin8CDb6wJc0BUIF1HFnEIp75t4
RVhymP/Unz5cjWTaVoRNTk+h/yv7Fob8eGYV2fF+UCgMb5Ru8SHn6fbmx4EYcHKAxZ/pdILxNk/U
TEEp52xIGNJUPBu514bjPRJICGzvWbrQU6JjmAYLnuxYLYUGg4JfNXGWcc65NLYVOmLVxzv7cB79
NtLdnvdG2usR73LGOaR/Kg3vE7G0KlH9i/KbsH4y4NK6T7iY64A0DEcLQ63r05Qy539xAEnzeosU
p140kT+OvZLSDUK9UErHlsjg2atCTbjbxIciUYqijX+seQeTaXR2olM/7G0HF1wErEQ0eVuK8bOg
qjSvSIq/zCS8L3+60cWcHa0Ym/JCmbW+0SqpO9z9TLBWAu9myoOmtvsjvGmznerby5KGQK9XrEn7
OQzCbam4ITn8XDPxG54jOr3+lB5deo44+PRpH7kzlVFk89OnMCq+srismuhuVli4h+/TkNnV01Ww
gj6Ufadj8scFbpWenZgxQBvT3nEd3sf+j0Fv0YQrRaLfSAq4O1pwK6ELOTNBxRuIYRmAVHS7a6v5
z3xZ9wNHFSGsaAZLEYpY2DMYv8pZVvKl7XjW9nL9FOSTbLl+8yooWBk0IkCaILPHAJYbjqurfEeu
DwPXr/9LsSPU9dTNN0HPcCVIHVUNvqldW8hWMOdEsKFKlfiw+iofMLUA09PirNB6Th5X+X3dQmtd
LKR6tSftcAGijPPWfvbB0AzsHOZOBs2NuWIdEUsi/gc8umN9IWA06PX3oDXE9g/YURLoFrOlPgGd
G0pCGiMyEtY5MWIu7DxkEBcWJ5sHSvxrDKUqew+jJ7U0P4JPSw7AuJRJYbPcmbTzvh7ltFTFO4Y/
0lHV8wVUe2udzXPBppaPolwufV9rp/ZkV4ENsJKphd6fErjvX7d5M1CEfIyqBe8zmBVOCVAURhde
5xjpUkC7YAIeqQj2Puds8kiwkXMXIMW7Zj9GmlvEgCCqQaPxbmKW+z9EfNzEqEN5Kn8k8b8uCNdd
kHw16zIKlP+605MNL5Bfdtvmms+XYcC7w3PBWfI+y23CkYUWEHFyfwYPp0QYujWiTwO6yTncoo7b
nVe1d77ztHGyVwMSLTJ1OKJGdDQIKWr6DoMS0D/scPhUn4nCxti7OtZPNhvmh3b2Emg1UKFjhqc8
TcmYUjN5strrVsjfbKsK7qZQ9i9FS1KIaT5grkDFGNZBJcZR3XcsmZyZPZ0XD/ZkJ9bxAOwqzYbP
CuEgzeVkA88a5GVP2oCONDRB270EmrtPT4AnJH8lGekCXZ6yVnDcJ9vtDvuDdHT0l6d8jlhFJxze
01Esdmv2TmlwZdJuZ5Zb7BNYgX2CAQk0FwnHgyR5XioaLkRVpXtcWI0AgLRoK0xbVrO0VfcvlnUH
lGsyPQu1bf3d0ACWkLKnEFAhmmaq8qIDYhhPqXwfEmicrVDSVN0FGrQFqHZCIPUjs0zYzrbL1hWt
7zWRrWE1KPLmxgQ4HZQa/CjRABiMJN9fu+OLLlkujr0v7Iqg94QCbXjFAgRlKaz+UXkxF6ihXULG
qoxNEZV1PhFQ5q9rDPwxpurxLgMR8kOkOjilWHQwCwpWAh7N/LkvBAbpZzdBFyOEdd/6c2iOXNJe
b4+OUtzlOcvV4r8dlUDARkhb+4pINox9YgijrEu2mYLLTxoGgx+Wj4p1Vn8VnWE6b5XrxU16j/HW
lfbfJL85e+wbovBgGDTBw8V7D9WZwTfkgiyYb65mHqEzb4DoOfkzePgDyLqffjSWpAaVzKpvCuFc
WJgtEqZLGFXF76xRmgZnuEWopOUwaNjz7mM7DEBVj6gUYyGPNdZmpIC9dPQ8SFlSMs+tNIVhmMGa
u+7IJ/i8lqusRzrWZCUmjFMkldhVKiK9FgQlqb9S5Du6I1t1LMUkwP33EFCUQio=
`protect end_protected
