`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38544)
`protect data_block
hTX64IeLyHzfa3tJyS5DfmeG1nOY/rEI1k/lSakDFsrpemGpSDq61HGkY9wsZ/6hyq44+dT7O44O
uSXE3NA7Wxzrb+5sAox6ueky7qnzyJxc9vs2cyEdT2aBuAQUN1TGiXVPqv0kGylk606Gz6ANAnMR
5hge6SzOhmcTtRkgDpDqdSSBQwwEDuaidDyd96Vaukhjr/enKmqm15i1kMQVnzVzrewZwq1uTmun
IR2Oxy28bFQmx8cyYTQEs0KGq0/3eZnHkt0B8OpAAaoVZ4EGhlAuZBnh73MQTg8koynZB214fIY8
gD+nkT8vBNT6/chVGij1bua7L5yGNIt6e51woNV7gtgtJzsLjXC3LF7tktnPuWNqb1RZ1o4QgqOc
m4WtXAbEHd4csLNAEFYjbN6UEdoYDGnTDCV/BNGPguBPc04NqDQ6qeHJsmUFC1ULpgB46sY/D0E4
Us24mqrSlmdpec+jF81ppB2OAx79+CF2OTHJhAV7yjmuCG85OgG15p+5GAJ9DHBOJ3mkZUwlAmgC
Fn3SfmW5UlHYqAY71V2igzqdDqPgX4iyh4T4YdfFkEvOGmDqVWWq6E9PrIAxqGoro2D/tNTK4cM3
2RSH/E4KeCaHW7+93F4hVOr1IHBwMYG/BfL9rGZu7kZPtS1L3zYONGtWrCXKJ+EkheGhjXBDcspQ
UXeuWJ9NKi5oM2ar8b2afrRbhrlCT0vLKgWUeCb446zbX0kIFECeimcglT1oiihS13YUMQgxD+ob
cbSN307ZGwIDVhDjOoDeGA5ojh4SUIuVhdEh56US+s24H9EATs8FzN9ISJ8bnQWeWq0bnp0eXl31
qPYYCuKKuO/bw7iJWHmWDKfkpM5VI8gKZQ6G5Rlh+cFVvAsjvrWlc94UEmJwxYTlPW8cP93Cq8GV
nI3jIgDc5SH39bnJAHwEZCnbcFSeA13IBeC2DNEO967atoCxmf5sucQGBM560m/0Uh6Za1q7bmkT
iRzhv6RbzFv+T2mP9VCaBZA+9Zp0x1ipwZfs2mtn9w2dIqYsU2osOZONUj7ZPBzJFdrWsS8DcJ0x
kiATwMymokl1Y5sPlUhnVuJ9Oq3NuScBI1WAQd9yr3UHR3QOLVfKPGHAtLWqkRHjRXFxFgdasVFp
Lj/nubEYL6EXQ3dlBvXniWp6eBOZ0jYg8jwe1VplS95l5C+5U68e2eleGnLvfMeNOue9wcxcivdm
iVn4PteWh9mFQgvy3Falt9wxRqP0rXv2ys+OUV2U2MDZ8Fb/adzRMjNG88IYY3xXYaye2zem/UuW
IfJvisBPssuv6ByLbs55dOV8WtVKb8FyJNtbvlDmXjMAlHfdAXvvcdqTSXByf+DlgDJ7qyaSTuTS
qcPM2du1KeHItoFmDw4aRoIBjKZQVYOfAfiFamI05uv1wbmKAL7dqOhVEA54D8F2WtyLx5I9CJC7
dOb+sxZhEQMkpfcA3+54Sln3rMX/jR97hpIvUuc8v8qLTjNz9gxXAezQzwhQtdKx+b6AdAgIjMMP
PuPCEdk7cpUh7GAUr5UEoGk/IkbBy19mFm2AHIcj4Hz8222/Jez48Cc3nm6uf0OI4ESjBxHRnrXt
YqQBVLjTcHh6InOJ5vb3h/Y27xfMhEb4TZQ7qowpwLK9XdcojFDm6C6HNZkCYR5TlQ9bsi9pFRAa
hcn6+i/kyIUsBKReXVVjnwahJCrblexuysQLRwz7NjsoBjyUPueHUhJPBgTCB7opEhPnhJO6r7Sz
zkfoqup3dXwFGpRzb+Ho1VA+9+ND7KppI2koISKTBlMPuPqfAQ3nINZfMsUkIIJwXzWrl9++jyce
ioqW9lGJSRHoHh4LLT9oa68XsXGctW9qLLCwQFZD+hnumbDZOUScm9jyWiSX0xUksHdt2m1yknTJ
Zk+6ZrjaOFbyoiwMxKB0v7A5Dae3Y5k8G7DGBHSuW1wE8yBPBjLWRTRse7JgWFBPT2roQ2Gr0Y9Z
e0YakqQnmgHaP4jv2CJTioqDHJHptybLnNDB5YQ8zEAosrixlb60lEeL6/yWnI/ydAze8eEace1e
wmEOFnJ5h/XCLDAmfOmMLVCHr1Jrq8JjS+EIsGfnvrLVLOKZR3FSCgiyHAr9pDqipJxdfnAlMdtU
YUL0sRJOi4PuBGo2oOwR2i6Ndj8Jl7ARJ6Z+ylOSQfoa0NDAIX37b7SwOd7EMB4CGY5VXhYTVevB
z3VBzedDcbmLsefVQodoCy3lDV/G9uVA8XU4GLMVkPPLr4wg2wDPUEV8C+Kb9sO1sod64wJ2ZI7x
fQbcmRwig0GKP9eRvE9qhHhVdmDIsI/Cwao29jMZGDnwDPznLoMH2WLDXeebiXY2vOybgK426KoJ
TIe1JhVUuHu3x8yuog9Lp6n5ksck3FErwOlrCuf8f2xOHis030Kzvo3iqFHdsLnUhWGS/pijHQwF
Xq3VDOlDsf7eC6HQVm0alsYwk2ryBs8RvP+ALycurbQ0OXTBecez/V+v81uTBeWzNM1mPIEcNCCf
j+YAbtzz4Ty6036gGMh1dooDscczbXpMdjv0fdF6+bffT8T10COJZlKesDjFac/AcJz/QEZm996z
p/d7WduquVg3TvkevYwrjbnbsE9zqK1m60C9w318d/9S3VaIBjlgkApeEimMgSy9A7n0j9Qb2q1v
z6WLLXBlWeLhe1PBobd6lU1kbtcx64PLWgUDCHsF0CzeY2CJCkQ9Lky/H8haNf9U0kJm1N7oY96j
Uc+vcXjOszn+A46tgXkiibPI21NkfSabnmUXRUhr8Q7k5FSv54L6+YIEGiQP3FpBca4HfKgBP1nL
lyaLZtEVlf7VebyYj8fcj+t7IojRNKUa9Pr0JrSJuURBQFkfKLT+6LNAnF515646UI3muL13MFQ/
kqlS6PBqE44xOM0GTbUBGth73gvL3VFHMUalj2q33tJSlgZoFI97Zqtb+pX1/HzfiWs71Zt6t5eR
rUg1PaJBXs5XMIDvKpv9coT6W8jnUOQVMG5HFYl8/gRo+eWt/vqZfxvmIVyPlYCXaRGSCNTyGE3d
ZPqGz6K75cIMGdelOqelbKr1ktjjAVDXD86wo/+r2/f+iOtyfj2zG+x9WeH9UVQRJTzsCgqvVySD
i8Au4wQmNm1NnBAdVkhzNl+C2ccjSskHBwgJnKdblW90JTK9VrjajWeSV6pirlcAYPQ00OOUGkm0
9GMhuMIc6emmUckdUjmfruT7eOsVQdh5wUpv+eyWYyuENz9p6Yv27FR1UaCaw44T56tUh0AgZBAM
IDHwXpeyVOVZJO0Zrh5unpTIoogSWr2EL4dwdcYTn1Nxugch+LlBnTxRx0GLz+ouSlXS4mT7G0v0
hYxIJOe52aROE/8jzr1Nb3SbTELtH9wHgoMV4A+16ZuxcDdKrlSAm/L62QdgQ9ao7f1ZeB65lTuf
Jy6VE9y/U4aOcW2ReGWGLUyeyQfiEkTtSI6d4wOBJ+3UQjWg4RdElRQHF7aI9j6BrKw3LQ/RgTiF
6xVnhP2YuvfnUoMsidfhWKm0NvxdlTWZxKrULXuaBNlH4UHhd/4NZLXFGh9PUYrxnDpLq27FnXg/
iYlp3uPGXeKlqFqVI4XrLDJOF8tDJtS0AptcJnoue6peivGcNNXtT/BzCQVOv0+x+nlNvN3aY2+q
cVIwhPo6WX1EH1yYyeejN062gm+IGO5nL+X8+GOoNp81+dBOwIfJdaCzAUV2g5UbsNk8U4ZSWLoA
8Mu1E9agcXLPNtZtVtHx8zXOC1GHZLf6xgJcMQjz8qneoNa21e0sx2FSl7k6eOaw5zT1d7R3bgWM
qDjXmvxQvSr+Qv8x39FoPDB6GAJ5/HsSwhRWfhZrWfX6PYv4YxA73Vc5jtf5sCqNys3QV7M3W7ea
MJZXV6foRsw7PakDQtIuB0U0cidMkBrNujDfBp4sawmjk3+hMRZIongVraiozVzTNcLkUYHRxwrY
HHsR05iHNJ9doOaGm+wo5YRhZ9hHPHNUr112F9Axhs6zhMU9LF0Pz86BB9rfTMN2Md+Cg9KZ/zQf
BlW8/FyuO5OSamkIeP7DJQm1SYRnfiaD9NhQT4DHkI45Gsc2uAyr1IDS9rwObKDH9kfSHEnmZRUG
3/RRIWZc32YqVpeFUxlY7iFbH2rEvDBNkNWZuD1volBCrw1qzl4780Xe+z8Km3IFXqsmv8J/2c8Z
mSNt4sM/zEY1rUW6ieAFn0Ds0vZ1mQlEF3m2svzriLtkTy6l4Wxmc+a62OWSjOfk54P8CuMpeSa8
4m4W4tcH/1Gy/KJXCGM8vsGs+JMi8xuUFYizWA0j6bE19UvpW4yrSeKC6JjwLMRQsoH09kTP+XYu
+fErJ7Y+hpb5DDJylhQ+YkTnOU24ezJM9hdGnuRFQkGXsMG1nYninUN9CHzZRrB6FIcvh/AJdxR1
vao5cSCRnNCFEmsH9H+vN9x7EPQbJo/g+blDL9Vpla86jJa7/kh/7KZF8HmwnSiDNBjx4LAPttXz
aR9A+ZeaVhEuRMWm4X666Ya7zhgGnZPum7BXDm46WasQknDr79Ls1YOadHgbbu5ZV+g1QFh360xM
SXvtR4grp9ibm93LHaPsrXoSd4bpJwlkxJNFYRRwZpSzfVeCs3QeBbhOXiUIFRG3Hp0m+2rRSHoy
Ae8KA3Dbf2gz8Nqg/Ct0F1AOuoy6rBd6j+lB4JO/pdmfAwTMW3lfRR6mapnG4Pz8coqBWGdDog9l
45Xx6IZ7sX9wOEwbZaeAe3yaV3iTNoxjB2pxDNzlTLJRO2vckm+fa6AwMJ3qOyuit52X7jT8y1P+
DcILO3wo57BXGcr0yMLYN21AdesAa0JhZku337KbGRucK+hCk8MlctUDdJGB2oxVaHcGSVLQxdVx
KZU8o0aQXyI077eq11lhY/HHr+Mq8LnBB73gwwiFHS7YkiC64gDBW2NuDSGjCPk5Y7SyQ9sEII94
bAhVKy4cWLQgwWtmQIoRzpQagqJP+wtZOO0HzrHjNSuCO6Tzra4Ol/z94JXNHmvLWQ+jfZQV4DKn
MEkAxAkxECqXfmAklSOLUiTROS6YRuCJ76eDR3S459+gPcYq6+T6JgiYtg3N8OeBWKKg2UpFsidV
1olEt2+EoLP9G1viAHXyqdghGxfUwQFDHQhLfBa45pY2+xqaXwI7PMElgoriKOsQn2WmDCRroOmC
htIJAjYjvFLyMlOiV9HEn/0HYWEl8j1di69kBQen7oMEIQaX5OZ3IMf7/3mDpvdk1Rdafit8xVES
8pHGKqHHF/OZxI+j43mmCff4fbJWARMggkB6JfCey0gUOMy3JuwGDXBwYQ0aI+1Lqa7txDK54oLj
qB1MeFU9o1CrdbHxu8oLjzmJ3fWwti/aODR/hERMD0QH/XgSlesims7602WsnqIC7/cR6u9sZLS4
2i1A8nl3T4A49xQqfVXe9+fRVx0MdF0RZkvwCsuFzWlwGU3vtJHVFJSWm+wZtrWWja+mm37++Vg3
NabdHDINo0e8cb/9mkov35PAhyKhMcn1XP+8gQXzCpFsxri6g0ykVlxNCO5CnEjzY9lEWkz9Zisk
4DNHe5mDYDjNzMswwtOo9zrotEAYSh3lSw6tY+WMUB8V+Qf6hCen0PEB4kj7BVvxYw0Mt31TIRXR
9qLYrdA1XiSfl8lxUy7vhVsEz5h2jBapGFunVPrHfnihLhI6BIBygLs2YjV4htVgijS5OReW2j+E
S52rf3cZRsciJpWhdCAGju/ug1eBAvvbyhMCyNHW/cbOy/fHYnFyZQ0RsbiS3NpT9lFxHcUKcqat
3SJtczOVa987lm6TuVA1UjAMeWomM6v2+PC8Y8vHlo7VDkanofUw0OLtwm511L0EkfnmPvMt3ANK
8gv5rYgY1ajX/Ws3zOIl30eM17Nmtm1Sz/gfpoP4dL3+Rf3rCZDnDaekXjoRjdz6+mZYYp9brL5h
WznXuUY3+QQ0KTcXBzdAjyyMrLOksvhulSskrDN7RWHmLfk8m8mZQOF92QikukRVJTMJ1HUga5M7
0r6xBVldLB/Z1r6s1UljV9RlEsYTW1DwMG3nf8C++35gUo15mLc0wcu7D7hYKXnXabXwJjFFjo+t
FdCGiudBcRHdRe/LA0Cq1O/WTCbPsVZRgZHhJCh1xxYto38cdrgAFOPBxlOmGZeBabUIejF3aOZB
P6zzhGVXg+8mYLRi/vDPm4mWbCmR56CLicro8hoC1XZa98gK2RFhufPlbXyTIirpoiQHE+RXNgs0
ovCJH9sW1QAszZTFIvZNw+9qKYaWR2lv1Y7Yn4e8iMfr0q71wPRDDwXEsmzZOjzftPebtyYl2zDG
3fx+4vQg06Y9NWIsQm/VmbM1nr10u2JiH5i09quDaXQfD4x6GG+0I5Kz4sA3PTxCE1trLBEoRFIL
miPKd1XvFsyikprS2WhHVX74XmL84n9ru2j8KV/L+E6CYWPfieuRSkNkmFSyNhnTlzINeNfIOcUJ
ILZJiR0Mt7Jj/w9yCzhnhyMkqx9oilWZZ6WfJ9DWbnfCLA9Topfld39NDnGVb7fMP5dNDuSzRTy0
xK5GmOYvblkKN75tfr6z9oKBY69OuEd0FpiRizVd+p3PI7fbXK40zrneXwjDd0pxR9NIUjVUQ9gr
VseBatNuUvGKrcheNNL/kirZSk9UqWMgFQgbnx2QT/J0O/Ah/byZtrwDphgWucgd6StkHqZOPi9M
Ya45vizv5sTxbyg2KgNG4lCRDWnKB/sP6GVPM3FTiJUohI1I1pB+ktBvhQmozU31IKBzA1MIO8tX
nE93s5hEOhDs0O2utTqQ09jLYLZQqRmxTKPKR7PYbjnHVW7oOik9U5ecZr+8oTNTOU42BpItAy7v
NQZ6lELDgaevgkBrPHs0lvzdfUGZMInC0onPSBZJA1bkcW2G7cZNp7ofKKuSOQXEa1sk0Yxnr0L4
Ue56B1GVB2KC4h8jOqOxyT74/+hU8IShaYq6z7F8K11kAaQEkFqZSHByrQ32W38yHTouR65L204M
8LUvxAHg2WrTMT9iSvL6ZMyVkZjGrlj0acuYE9z3lQR4BPCWF5w5mlgtbf7LcI4vU2XfATPqjdOi
gvRbFfFxeBf+1zWC27TRXyrxKepWVa3oedVVU9Q/hanAWwEcM35W87eaxLktderAz7bn3NSE25U5
19PwETy4yhw/5SfoP4GX8TsBUoiy4OoS3kFNWj7/KzvPzrevUFuhzSKPV7UU2QACmFhTjXUn0x+e
PbfGW015vtiBNJdrJiyzx3uaRX++EtMFiyiDWW/7GudHcS4VHmPL8Q06WOM/8wEY1kgjeZfnRzSp
qb7HN9B92XJNxr3ngZUoKwyMv9WFdewiIMoI99X7wU2IYB2XHFrCov3Umus8ECGogB8Qa8ikc8M2
MQH3tu3HBkv2Fo+lyMlKu14U/RfkJGpIJ+eyHQQTdgz5ZxHafOSQcjVu/A3Bwv9Z2xrHRwdW6iyR
ldcw97a8MfqHoj+i5Y0NoG1mLV8G/x8u98PgV/+M+nWnctHDKU6ro27ygo7KkwLbVnH6EEVhSvr+
z3TAG4biCipMsbYSHV+d7q34nE20uUwXAe6wIwyRTGIGVZRMg9fHpMxOapbkF9fjoMmrT7ugjmlX
I+5CZHyccRBxnSATRZNLkXZBSoXpROf6/HUyE11AhltW/d00HFLIAdxFI3GaJeEpRr2steA8aThC
STADqoPLwjGUBmAOUE3m5fgDYXgGreEDzEThNS/oNAFfYAz2eBdZsffn5KyqvIvn+oa8eJ0pjY79
7Wm0VUe4dt3of9wYMdL1VGCo+HXwC92XUX+zd8eYKz0GVm8nqPHAvjM5yLhL7X5qTIGXHGAwas3h
HU7xd2V4x69P7Tk8np065C7nowAbZfRY9VxcOdpsKQ/VPJC/YrO7PiqcCSon5bin06WwqIGxZ/5S
Xq5jEkFYmCjKTzC5Jhqj9BWNsgYwzZG09oezefC0znOXbOtfgYqeof8yFFDisUp6BJ+X+Z8k0Upq
TQK7qY3LjBsq+vRGMq9mj7jRJleUFU6BxFEKNkE90CjWqyFDRgw2G4U/ZdMdMC1HxnzB6cHS7jG5
h3IXJhGMgCzrGqni14Q7ulr2hkhMWVGo9VrHOCnxJmU5MoIhsH3jlXPkRTrPz/CRO3EA6xYGgEQV
0lwRC0V3sqYtZMJ8P4bKugREKUrdFa7LN4fUSnUynlKKQH7PKWnPpy3Qizbsz/7Mi6q1zdaV3B0f
x7djT7LRKArxaDAxAmXKIfbc2fjOMcgNw3x6MepvA7cSych2CWSGv2XU6fQ6ZgfikSkNQxKJFbUl
oW92uIdroHWJrCGDrl9NjRHK7Kg+NWOyiiZY4lBCYXAe/nhm5f1LZq+V6tH0u/jI5jO7C0Pb0B4W
vXUJLAI0lEgnW1KT+LYJrUQzvZ74AlIoGNkrBlbqpc6wxRi9i3fiBGL6mFf65L3aVkYOg2NxkQLm
nynCNxivvcyHT6HSKkAjmMrh4B6L8ezy7LKmbIjFBpuo1WvIcPdomVQd7BISp3JMQMdku5g6mq+g
hLNue38xZTDqYL2cl0ixS/3TNrbWNeGJ5DsKqyPJRILCOdRXoGmcGbLS73qeGpX8/jaCvGEN0zHG
YaenEFDeDhm8nrgA9mnonT9Lsvq6yNdXuHsd2LG5Q3EiF+iaBPsItgSXXHLFljEaoncZdy1ZqDZL
wxZ/jpMO5a0wLVG9gixMpz8T92tnHApnJN35Z7ybWmM1VEfz1gF/0BKwSy7oBk0zlbQqiEL4+FPl
fjSb69K1HDx+FP42CyD3oPMKLvMdTJn5bhIJ6c0bLvgRb+t/hcqzBju04Jp2cStTf8rVPIubVUKW
3wLO+NxDEGCCtDyDtARmRWxixYBFLuLT68NduOVEhpqz03CgiHlG6OdaxRCn1mfqas4WHdJrgKj+
rSiJ5CU/7x1tNphgsIUViEVQpJek7iIails8D4QYa/5AS8NjPHxHb2k+5/nnVOozFiLXidhemDxG
tT1MVZDLGKgf9kNLbxOuXBJ8hh9RF+SsHKuil7KNGGOseouuB0PUlOZOTuf/ujNMYWsh2JhVwIqz
ojUhiRSKA4IPBbFIV6nD0cXfi/xiogzWqHQX9orSK4/mPgtzsHA7RuCfNFrTBLNs1l8Sye3Bcs1L
6oNyYAkK+uMy0c1gGlqNUXUcIhFdX9Wya+aYJ2hlheIwele9IPw822xY3sAM48x//HbkND2Kpu1H
CEd3D8VznjsJAJfDp3F5C1tf2uAHAM5eReWM1Bl9hChHA7QdyWHE9oHKPGW+PPIaP1SjiHGmHxD7
6OneyvrbLzO32TQ2MwmWQfhZoXGFvW0b5LPCDD1N4NuNHrWWQ4tILTCkFmTCGgOE6f4VGTH8xUQy
HMsPYnIv9szQxc3FXA8OJWJMHzkilE0rL3C6b5gWsAQmlb/auBd2fwWVVEmWt/YqMvOVCi+PMuz4
3M4Ir9Qu8AYYShoOcS6DzxjREBDZekhlG/934TsDrJl6CC76FPxL+G63R5TyfjEsW/2ssGZhybqJ
SUqDjoVhr0httcOj2K2hl5NYxI9VhbAvYEO4LzqMFQyH3P7fsXc347kfM9SM+OmKzJi2btjh88jJ
PcZ1FBYTWhBP09m6vtFjgj/LaEBgpCWOF3LPwwN8Av84TAcs1nr2ev+znqFplBXaAzQaj8Nbjdks
6ZazWtK/sLeXRWWZ3Am/7AtOM7ibPWK0PXnfNDS/aJhLLNyeoKKSnS3GUqmFg0XKgv42ZWG05zeM
y2BtGR28B2aA9KQnXHBOj9g+5YgEsj37psn8pQGxLHM+M9KATwwONd+6OOUgA52b5IlfK+TZDyXT
vCDkLQTAJuX3ZIv3NjD2nAdJW5hbQmzMV+BXwZS6TXgUPiF0mTM9IaH+FkDbf3ndU+oNGOhmoDoj
oKhUWooIGUJ2QAlFg8lzX3+0M0EYJgIqfJVyr88cQOya/F7MLmQDdoKiJix6+gbDWSKFZd4Agnc4
ffcga/YnMGNGO+hCgJvDCBEiRl7ZYPNVwr9jPitimWrV2M2F9Vp6ito27pU78SR1v/aGBj2oC1fG
p8dsPYoSbUphB6r1FCca7bwVCkgQnfMRulMXx7fdhjocsSMwjQ+3izusNsbKfbE9tb8FRbyOvBm7
1FjEXf44cvoQyXZ0svsA4yH8LVzCurroVH6iAqMFanvbS/BHDIPhBbsKUdSt4b6Ik16ECIwHLBTF
ehjrqsMgP5Fg1rkD8W9FDGhu6v/ZeoHobzKLx665tAMj2AM+AaOYe0Ey7ib9r3wfNToZvrZm9l9M
Dio04oDiUj0R33gHC+2FucCyKemgxYMXhIHh91x0VvS5W5SF5ZOOOOFNl6rQZFSFQQfqsoQK79mu
13ffDaQAno00Fd9Go+j1cWB4LSHly5rmFhIRmRcS78gdLudGLM8utIrhRaZYPO9HlbQm4CazxKlG
CvDH1QkJla+aRlcUSQFB+6pGBSaU/gEW3HNSisM7rQRlzaBBE91Z3tZQ/2B27lr3i4HKdWTgoD6G
MNB5X8ORgYOYockwcYbsLGIoPTki5mQHm8deiAtcsqSiYH2YOgPBKnTEPuOiyaLNJrDFcGETYAkL
BU7QJn9P7i5MoQw5WMebpDv81Ptz0EUdwyrGiXq9dxIQfiAks0eMfs//8I1EjhlR8jdGnPI8Stpv
vUd8af4nBr1ZtsntovWmQsnZAD8ckhsIOQSij3aWMyrlYOwuI/kNPzZHQ7gtjVNdDPvmvcn12HEu
1fJQ4EmiXpUoNknBE+/JqRjP3WZIUNJ4xo977PfbuUxe5+8nfo/JFf6n2kIm14rkP6M5NO3JTh3o
ptrTTNykw71fajqNOPexdqYRVcZqRrK5bcG/1sqAfV+L0GI/XuNoTfPYdGH1nYub7ne5zQWveKdh
7AvsWHFx/tttpcAWjapJWGkAkXlkaYrfunti+NP/pgLD+15th0t9lKTC2Xxk+37cIxHjKEr4zTs4
jDFPoPta8Q6IOW0SjbfbpcUsiknUJuMsltRApZSflY/kLiKpLtKn0sUhwRe7aoe51DpFiAnqXCWS
e3xbu7pzRQd84e+Pg9p4UlvN+UBn3fUPQL0JtmD7Y8bu0NWhbH12EDIfzKTXpqSnWagRY0ZMgS2D
/Hu70jURcsYQGCXu/RU8ctZcd96fsERb+0Dv0GxXG4cKLjmoXAPnWkkp6lRY+uwbNlq6OqujrYFP
W1P9HETMTrv/Gdq6nNFeIrofvBDhaiXUwiCplcDoK+UMPYHRfDq4QbCNp4OzW0BrHno9eCAF0qjb
s7nCBD8DN+gsprARsrBA130oG8q7odOtE9kwky/xuZ1jDgw9lmMzzQ97jcnow5hiNqS2qzERiOiP
ZnydIf0zR+4RSaDxGBPjODxoLE5aDDmuWGnltHxCRBIG6O0HT6gX1M/awLNcFR/RZ4D37vHvsqm4
+6/MRuUFQRpfn/4RSNoORocz31dymwKlUlPyIrFtuAry4f7kHjk2jP/Iw4lren25wWgTdOaruBrU
d9EIJsc2tdJPyOw6nQ0lvj8MKugbmYlq0S/7n3W8PE9TSdH7R3IlyW1aF5uMPG7Psy3+ZdY/q79N
Iq/8ceBGRGfzptR3wDv7BvfIkvrMYV2mE4XGgkGSuhTiLw5vZs1pdRjx0MRmjw2BVAGOW29fr/00
j1o06mQjiPCewfyHf6Q9TXo93n0A36cQKMCXTFz87/FV+6uMLz467GL3vJlIyBU2+0dlwy+MhIMd
eYwaA4cbGuT+uiV0hwdv8l77C6mI+7PTRikUNPNdRcisohNWQkAEjLK+khdGySTqoDN9fwsWLIcX
n48x5YumGhHwOkXRmJh9cS+rOYHtrlxL5mwqnIDr2F8aFdNKXElzSe33azspK6gUDSYsmiSNaR9n
sm+E4X/gM950V3RX7ceCS5gaElGmikxqJFUpaawLkno49+pEj9Z8u4NnhsyCys2dw8b4wk6x8fES
CYkw6otQPvoacQr8J5dBP5NDS2bMt4O14ACMB+97j99TIZKhjebVWQvZYGmy/YDCr90fVBjuZZFz
wLX0la9gvLX5y9sOGKfr8r3U1PPzxSwkJhRnyc4fDYgM4z4OE+R4qr2iLHWhQJXJ8Qvcd154LNe4
VOGiKpnhRsDCMvxKj42mwp9hTmhuGp93/Q/eL064m7eMtddJLGqYp4QGCvoq3uXTHrGR7my0Jdf9
IyrHRAQzSVegiByJVQqZhURQHKw6BQ0zsfUm6d9JUOGvfOJbi1u/tSmqI65ZsiVhNljC3eaTf11m
Q9EyZ2SjBKHSo5U4C7Oc989uoQzMkCKkDNzgjO2dTs1iDG2buF6WhECqSOcpMnDXz/jpxhlmYk7j
uy3sB9+8JL6EK8YuW4xYOFcaHaCBWcnvC15NF2hA4YTXwC4z4iO85uF+d7owZfYDU9bng8uQR3Nt
lMzmlXRUV7JM99gVGi3VcMBW+KAWull8Cygg5whAz9p5eDdjXk20KubtMq3RROlXUGVdn6IJN7JK
Ypk7bAjn3xZrWzye8k6XheOFOfQXuVDOJY/zVhkUUu4y666kDGpXF3Ky6GbjRu9sRxYsEBZlpUhn
+J/w8LIX/aGEPNhp2Mv6bX+zVFbP2xijH363iaA0bqIkkPIop5hrCpsoQMaOJpk+1hVP7wokOtye
tZBDIWUREJYv+PBDqXfuKb6eeS3Bowi/67p+AUwLDkitS7rhG3NA9GFHf1waAx7kKgqMJiBqsSAT
KfD/62JKB7T+jJBFVnAkY40EMxSxpT8gJau2vrjCXmf4iYQNDZgMHPpPGOZ53aNiN3/qX8GHy9Ql
Ti/I65XVbHnVBVw2a1HbCrlvFJoPRC7Cv5/ScPVdtitFckKUGXD8CNRaciijYOOoGHGVaoeTcypd
g21/0KNw2jfQThkPd/+VANFSvdKok8gNMwS8ed6/CYdV/8kjlHM2rRpy5EKhf7ofSl6LDI7bmoWj
C/gWC/qC/1regt2gnzQB6JJQrhrDxoujzhGLhdrO6mrzsYKvZymLoo9i8Z7kRJzJyLlGY/HtzLgu
dFoYkipHogosaDwczcZFrUxjBD4ejomURSsKiB3fS4mf1ZSZaVTL/t0k90WpFg30J2sVPtxkFqgC
ThWjNAzyTJ4F/Ze29TgymeTNqRogkdmwH9DPbwi83X6AuE7IP1mc2jcXj5AmBXoO55ajA6Kbdd7W
gXFNZZ6rTei+8JpjGZSgdvuYg77Ao9ZNHiapbUxm0vq5WptXmtOtPTmsrJ+aJjZP6ZomDaaZGnT+
0NhoxM8QgzCBY7easNNc+OSpo9gezYaN3CCltfWLurc+IiAud/wBhRiaZjfHCjj1MzdT0vR8X/nL
FRMSmp6sKIkwf4OF0HBXCjKqNmZnAUOgSCvxjpQ/X1UvhFXyq/OBMys8Ookyc1rFHn60u5nYCCai
6vUUuNqMAIPOUreXv1Ott+z9YETUnRmXZYmBZ5fPSeHhywqRIGEIIcaEGUl/Vs8QuMKSr+YO+kUw
LZdm6rUfz99oexsZe5a5S4bkw9Fltk8/Vy5Y0q8jhVjt5gT4IS2DhRO89Gk7IkSxhCgTYVAgxv1r
dJcSr4X9fUzIP0/EYExFKMp/Bqlrymh5dZpG1lkwY1Xb25GhJmIaxVeEBCJgCXtdn5Q+oRwe7Dbn
WKfcoswIy+tl3wdbqfFW5MZKj20zp9lvEW+Jzc8h4h/PLTG8UZ1gEeaCGM/XOEY1jYmxfhJpPGgC
h6E+RUO+PAxzhMFQXEVEQh562n4SkUrfJX3gm3CvjPe/b4BWYDa05oTkmjKiaX+4f/Y2wx7kTQSP
Is2o9W1Yfs6Ilc+iUxxp+HLxdYzuahSM0dJ3Pcl/vfou7fj2kV9MQCm5Wn1C6vIVALh152/OxmI/
GtL93IVbMo8YPYzcB8zL2hWZlgFnJJ5t2GEtYYLhwR95a/FL45tuxvQ9Wyr8gugvMceeBJAZFoy+
nY06PapiodU7zKBCCrpjzQGQODLeXe5GJS2MSuVZNoF59ebQBBvDHe3pyLk2kBBGwAMZEy4xbos+
AvlTzBm2/QO8BGnTKQEB+Yk1YJRXaOe56pLk0o8Cf8mXGVt5HnXbuibVMJr5MhrOTj9Rxvp8r8+w
uz2kxn0Dys3vAIqupZxfHOkP6KiEnHRzV/5l16WM6qj3KFlNp0IaBzEriv4zU34j24671dhSQWVb
ekif1z3nDLj3acJ8j7Iu/7SXH58kAloGahS0ZVO7ooXYd1e+j/36Ytw2otbIS6/V/ZgpPjU7y1xs
lkCPp5/zHs+H9TfJ2Zeb6+3TKJTlB4NCOse0Cg40PUoY5/W1yHv+JNngwhAGu8XhVvzA9G78GQNH
X3EOZ0Czp/Wxd/KBlzGRHscPOSZcbKzjhVLcNwjZEhteNhy0CtTBEaEGkGSTcVTa1t4qIg7bEX1J
a6Y6I1bJ5Q4SslvDOYVcbUXpa+hLCh5ADygHr/7GYbii3k4Qj6uZtdGzVGjMu5T9CV+/phJigDl2
Gy2sEunObGI65rLajjlWVOBBSZ7mFu2LEje1jYb1J8giSLs40k+OQY92JxOOm0UJcHGw5AAh/mWl
lDspQ4KFkH/ovENpMWMViu0cyrDMhXyHXooiIR1y0ZTt/qceO1AK+AP8P4hFPHPq4aGuPKbHbYqZ
uMmToiht2PneuBckWcoyk0AXFdlZ28vuV/achjmAXO1yIbU99XEV5ECw0vF+piBdoDNwA+l6luM1
H3y5BfoqQ5pW1cZBsdz0aYFwA3GFis0SK/Hvs/YlmTn6SWP0ReKWSmhuEtQ43DW3F+OU4SC+7YX7
2Vz1JBVjKUin8h03ywCltrcCa6SDGl8GDlFepgdF9sFgt2YtM+Z+vJUNYL8vDqsDW+JbQFi2Z3mv
I0QB5SsZwYhgGfVE9e+4rXR8NBMW5diG5EJlLcBUgMKcdgj5zB110awkiDS8yXGfT2FU+bty8lyr
+KKTK6kglEAsDfY6SnSVpBEY8jcqgKk0Uvsdlbuk8qFYXs7Mr2etcC8Rld1wGuegZsESaVCS56t4
TD1bAvIRBvFrybTXmxstY4bvJjO6XC3Xfcij0JgpGHdagWBPKyJaKlDQZpFbZWeCOm7YmanBmZwo
FbQDBaDK9gQuJeD0AyoGgP86TVZEfNYYMgs75eGdMvKIs4Uk1CttDCUAN5bI346+t4nc8nM6N02D
RaxLvXy4IF8bchTAurq/CrEL3l6hsySBnJGZRKHm92ntoeD/5qyeTgurMSVFlwzGMB3QROiVHy5v
blmCaGLkmBnig9AEUQbmoSGbTgI8UVrYLLLOwWTwM/F9GPV7JjT3VfLyqXCMUgzDOnWXMHyib8lP
vjb0iGDkR6yG5nMs5yKKEOcY3yppVXSyAb91P90TH6BTwOLOOg50yX9oHyAbk84KA8wta5lkBPLh
jJqmfMYSHCqkui7q3Kx2rs7+JeOzYpAxJDJuEY83hEQrfhqge/1+ScbXba7Rj72g5Vts5/0Isq7s
WTqrQmNWI3qKZ0394HjhxcG6RSz4FrgHHfZhWurwFFg9njuesRJGWsl8cT77n71bBeG+7FspeZkA
zKB9xiuOYrgCpBR1AlVorDCRAks2wLhna+i132qtOoIauz4XZ86tZqGxrs1JodGf3kEQWEq/tzzI
ooU0NW0QxER3UvPwBZw2klWi9/yiJ0Np6rQQG4GibBufxqJOgTXChoCcN0FuJ31R9AFUN46qU8QP
Yy+ffkC/wnN0xPrCbe+SuWvPb83YlDfNAm5TfDgd7mHn4OASRgfhvNxufe/NA0trphJw2dF7Rf7f
A3BrICFEsLzyek0yoLnegzzF0M5xW9h1i3gtxmeqTRDXvuG2Q7k9PO8GlQfKe+/Zb8XFbHBi3V5w
9ZJ3jl7qwG2KUDeHFyXaYEsDSVAz3DwgkHyy4A9L0weWfyZFzIs2o1pnvUGoY+29i89AcCMUYGTw
F5Wg2dMXe7KZLZQp2dcGwTa2AMu9mCP4OpEpzMWWwbgDcy7ZqBiNlZmEtOmC2FDrN4x876tfa5QQ
qv0PiyS7kAFi+Kj+XtwwsFnWrcyERNzyMpRsw/UM2JOuQCwEyQImypSHRebq1qcVueR9Zqb3vZa1
bARMqzOi11bYpP3xJL2u175BztHSKzuA7U+ioQZ6xVqzRzpKtdaxvxhec3O+ZPDyxhp/4BUn35+C
SVErBDaHkQOoANk7BcZdZtvCvqmNscrcidmxP6oKZktsC38CnySPb+q255+Nj8UfbnDYKwuG/TU3
qahXwI3nxaZ5FyP+9/XKpL1y0J1GhIUVhwiev3loNqehyEmLptmlkAAQ+lRgS/49qSX/s/upnZRM
zt9h9jxeY27hAVnEoy7+Th2d+IjvRWwpRNASZ12j+M6XahyaJ7oufYdIW/1Kz7i06x/NcltbPEbS
pB3rM/w/F9p66YUZCDW/aLCEhc+3u+A195GP3ftq1M6nPc+GzpdD85MzAPc/4Ln+Bo3MpfeLJYft
BOM1nmeE/hZlnnvLEFyxGkCiqiLkhVirZeywyNqzEKJ1vwgYuXF9bIpSyUfPgZWkZaRTxYaU0ut7
0u+9093bMSKs8yticaO1Pc1FICuOAYgiglfw+ec3eMaWZWhTkY69zsTgWEJtDTdOELcLRYhLXIoN
6o6JIIgD7PwRM5RKGWVcyqRTgDWBtCQYpMU1wIAL+NN4F/6iAnEicv05z+aEBBrqFo+g9imvdKuv
FQAelQpEGfLpHyKMpCXZXCXn5hRLFlazlImuCvsDJvM2gNxFrgGq3GWHpjeZaZn2FsRovbDP8k4W
BXH5cQ0jUjpQNq8z/9nJBSlwSBzGaFSkAftWOj+by97RYaynpH0tUnMzTGgEf/Yu3SGrxS9rV025
7nyXIgObdL9ih3ufwvv6/RUourLe1aAAhqlRHpBDAUAXVik606+dL5EhJHM4nCJ7VDr6MihOBN0S
X19H/IiW+lqsUf9QW9X6UqsnStnmZIqRfQ52BLQyyG2CbM57rRwKHACiMNYdPtsmiGmim7TSLMzy
0p3cVbgkJO6LEswPxiFyjt10Ntd+JL6Tkn5rIBXHtUYEsxKbtDuDmsrXxDAA+1to8/Ze2OeRy3qV
/tDY+MURBAdNGigvS0+Wt9ksLdYviqSB04LclebrhZCT7hoMLGwjveCQBHVXmXGEt02lpgTVxzaV
3/ckVFB0QvcO9OzwSIO/+2klDuAHTTSEdfD/VrQ1E7fh1Nz32Xj8As39l/g4DlZ58NIY9b+ZrPj3
9O5hPLd/aqSNBsdcNu6CFziRInre02Jt2ueRVD9/RBosSZqtVN5ZHu5EdZriDuQvP32uzP+RjHlC
sDQFkv8R0rak/gINTIWElexwUYSMg9ZUscWlCq8L6LBuxw8L+NzWsKIz5DOdYZXCIBLp5Yc7hike
xtCx+bUmIBI44L9Fgpq7J8ZoLw4ZDEY4YQp/C7D8q6jM6vLpIUWkuRkgl4aZw5EbFQUB30oJvQqR
lEy0KudVGccrGYVYnDQ5cjez6LokvH+rWuyZSoSrJ5pbGmhR2rUKLLI1m2ymK5bDzkIaHTK8iy2J
qJbG3ClBOSs4WzolDp15a8S4bIzCTXeE9XcQB4jcTgz87Ag6i1eKko91tihb0mjlmH0CboGnY1p3
yERaPyCvlJVQJMmL1GaL0z6HahkV98m8CotfGCp+aLGlNfhc4vn+tKEvlQKaxEQ4aWiF+pHmUtib
Jb7VuaI8f2goNCaT7a4V36KIUvBzVsvn4BE54dgrC92UsrxEIx2WZrc8b57tZIrD/Y9egA9vTuT3
yUAolHKwY5lSjgHZMWn+r+yA54bpC3mr3JQDyljIJE1OzFoU2xdrDvxCJqT1CQod/1HPe2y9zXJy
aBRPO9FC+Mw3NrVOqMdx3UvB4nNbMqmpbT0dNnF2LMpxzN9vW5AEupndIAzKghp97YZCiQvPXaUd
wfcO4pcqhOCPIeXI+ArJ/UJpKJQGO5+IU2RLYXWjjaMTuaL6CNvYTmRAERxpFxED02wBh15xjp/l
br03vuT35z9/1eL2PXLMeB1mE1OFSZvCXxQFXzq3o4YMr0/S9Vwa0Yajy3BYf0Z1MzFA+gUKZQQv
JfHTcM81DBjaWMSZThHlEmgnril46ExHdgqIEIZ2jTOiEv+WtSXcxfg4Ac7hdBxWjw2ugJ5nJp9g
NNXu129vlHD5XwuWkPNpe4b2iJI474jKijDaHLmi2lhOWNuE4rnVbxHnAeNt6JvXmDQ5ucuJ3Smu
bstvdTEAIdC+GoRYnEf5fCGwsZ6HvA1pB5p3U7PNFwsNBOgqwxvSb96MlMh3UEXoVGhN2QtT8rz1
tRQQ3CYE9hAp8+Aeorb+4rKOXRgEMGSFY5UhStP9/41b/oPKPghC6wYVjOPOSWZBNWw+RmQkqbWn
7WSengbFimzv6KFZt5p65icA6rSbN+dqEKqvQnkcgzeb4K0TxwTNBE3P4C2VqUrpYiMXFUKn/2dT
ijRFTzh8TuR4ZBmDofk/+VTSFA/FjE9lKu7Q210Bt9J5NuNhZMdjbm57Ft3zQPO2Zi9cewfLHWI0
0DCEO2q9CZ3cxCoBF28+2TfvikdC3eyw8CeYtOB8RTIIKKrTDF89IVvIZd7ukMy1+y+YSXKaisHG
4wU1AooIKAI+vKd25UTwhaBt8rGt9SkkSovLkPcL3KrI62sNQ5LQEmMjPIAVstRjsTouhsgd6DOn
gffpG2O/ldkV1o589ffWyHmbM5N7wHuAFGI5XPVM7+IdeLnyavLEj01EmIeV59Tf5aWaJQCmojGu
sPPfBTCIsNbzB7XQguuicFekNxKWnGu9pe/O2DF+PFy+LP4fKapz36pHaCWUcFvheqbnD3KkrhZ+
medF+X+6vV4Pmt/SG6PFmk+iltzPuhz/yLMSFoD4zMKMUH6MK7yUm98ySiMJEdEcCGVll58FgZ4q
2tLL5KArRT8H3DpNbFY4/JU4JATOQ9MUvZ5xuG0mTqCkryr8mCV2oV/kA1JX1XTpU+esAhlNPyut
XxMctL4RCA9pr5sOabHTpkk35kB6QLkXX8p0CFdZxMy6Fr0iFwSX2zrytgTZjJ4kfTsoRQQ5giqV
5k62Cbdii7GMaEziUOPSd9c3Te+H0lkMpDI/3wuKS7EiN/8CZM6JoK1Iv9wY3LaC1BPnmklTfTQa
cf5j8c2zFjStD3xpJ8ndMTuXcL8tYKk8C4CC+xptMMfMqbLjcuIbgTF5LHLRwiS7CT40VCHMmCfx
oQ85Ng6cMPOvahcVuK5XmXVgCdXdTFl7020Dp7zD779h4naPV2UjFq4csHtuxtdK6BXoKFtujH8a
esKPhKhZn2j6gLSYwrSXWywDs5udOso9khffQKTVcRD79nazkIu3648V7ncSxUX3+SJYPVhu/1gW
9IPzywrCQ1vNnzq+s2ZAvIBr8z+zvU383BNwvLS0uztVMV3CzLZF74rpTOEwWyZ1zlUCDzeNJxUZ
gQjW2RSI6V1Be2lqsh4NTQliuoR/OQA/LBrkgIIMtLpjfj3Cnp2tdJpMWi1N4RzlrBWo+Jgqr+Jf
93uYlq3taWYwW1CBWMJ7ZY4R2xv7wRrHn7B/+UCnozC7gKWZoBpbCQmca05bk5LlPjSKOq2045Lo
GXpGTVt2DdkXR1wxudcf5a7f7g85aYPmzzE7OgO8K71377jwjct0eIE4Kojy7A2yXVv74q8XSz00
ePYBEQumAP0RPD6efRrR5TqNU6dimkD3T3e6YSy07OLiuHBlvjv01w9KBl4FnWgd80frU8KktoJf
6+7IjrMGZlMgGrhesvVCy+O4n41J1d6/6OQ/7V6kcWTY3H7ghPSBECYUMYaCJsi/mJ/o9ov6mNkC
uaEDDyFt+VoGrUsLL2XfYx2FP5CK+rqcNi7bdQW6W05dJVkq253UgNhVyLYdahLdpjH7LwzXPsvD
9MTr713VcWlqxn/OMCnP1JU/+ADbU7Xfb8wQjJ761E9FaQEAiuHyk5vchzU5Nc7RCTFD7Q+C+ofc
psPSiVMudyar4zeuL8dHUdMT4lJ3Bg0c+UwvTMZ9A0eF/cRTN6L3l1yJZIF0IcTMqdcGSV/UmQHh
064sDwdQXeeUpZwjTX/0nRlkXaYYyOM3bmCv3L+o1HcRZiigUIg9bdRxfRYHaIqG7VOZxCHdkpmn
q7XsctshcFCJI8apGd8LQdoN50CoIwskEPueJ4fnAbeOnP+mlG0O/GlPYuGbPHiBb3J9GtUUmEyl
Ms3jp/zQbqQcSzvUtQmcgpl+h9wLCrhLMY3nO+iAWrahTWLZEHVjzEDDNuVVTEjOH8VJP9hOyO/X
YO3n6fX3p0rSMkQQGT7XgSx/K0oSMXVjfoDExP3sJm+WCwihsEZuzOYxqh/op7litzKh/YqmIEcD
295ZSHbV/dNBzGs+EoltYM7Z3phKVG+GgOlDb8qVgeaSX5uY+H2jwgCiXN3BHliJXVr9LcEeYtrr
w3V6UmfknMBq+6jM5peBMXwAKP2KishS1vbZLgHXzqvYB1Vla0UFxSOHoFk3XTNgKAy2rsCvEvW4
R9jwXwnuJB6UBUtJJZzC31lFeNABaqq5qUDfaqErowaSQcWSbBSzRCpv81WAJPvcduX4S8JP+AY0
r2hqQ6xfZkxu2Q8MAi1iSBgmbey19V8HuhHhKcCLlJMCAusVESfASrl/KC/2desPpSod0G/FTHA+
Qd/2BQw/C2IWkPZOyq+u9Ls/nE1smSQr9t35Fs5sQPwX9VeC95ZkspMzU2A4BP+vYvrD6vixZw/Z
bUPVyAHbpjmYvl9ivTSTPyKTmPKxZb6Wp05RrrxU9hqV/GNds8Hplz2cknFghHTZyzjG18eYjApc
cA8ObOumS0+v6vloHNZI+cTcEmUqGm4MRr8T4RX2ZRkHfnUT7cmlUtoGtDX2g90G0odli6kpI+c+
/ryrjvpdTuzWn99jMAtClOJ8xBdgzkC+fvqUAagTQkz0ezM+WX85Mgx1WPjSYzpZL6G1fgEfSwpq
9Xh64lrCUd7NffupOx+fGahXOE0HwID+oPdWnxJXWYOXZwViCU0PYZij15mz4bVAP/w5cPzl51mP
ByGcX11Du2p4f9NO/sf4yVHiMDDiBZ1r5ZfXZOdUbthIepj/JnfYeGMiVsGbJe/aGKuVKQWFYkq5
rhsBBOAk9yM4M+rRiwI3S8kCJU7bfGJW+diR9JhMjJnLneo7Ra6339SGf4ahAEqJ+THfZRUiRFpC
PJyIBsAgIa2mEnxZNzhL8yJoo0+pdM1Qe+LJHzUoRWBExS1miYqEWsrIDqTN9RFyD0PzJw3t3oZv
Dt8wheWflGWeq9iYLmR4uxH4G8fC0NrJ4tUEMbH1/wWOw8w39d/ujZ11hnteLWvZ7CoTSyjm8YwV
HtIb9aS4B3Y05oSvRHQVGpMb7zttdAjJCK6znLneNok/oN3oPSz8/AW9+siJrBHYRT7RkJ2oJdwH
C3TbhYKsRUtGzBM5KEQeXybrVm1Dep6JqO4J9A9pfYAGndijhXT3rSQ0lgBciglZM9OxO+SYJXT9
K3JYEi3BSu1ys2EJ58GI6MYbN7npkkOje4ZTcmSCZPCS6e9z3mMl5UC3q5rMc6OJhYsuzceXV9Bo
s5ftxAAnYKeWC4tKYvXOjr1P9Tu7K+WDLAESdZhVgVzzbW36Qt3v/bUo/ysm9R0lVNgEdjHlcBHi
Fjal4VZTCMqGF7UdNutXu44QHpb3AQsSkeP4D5YEyRyngIvF9Nkkq8V4xg0Gv9NDzZq+/LeXLxjD
q95ak2FWKH7BYA7XrZ/18zMeo+7XwnLcvL+iDFN6xnLKDUmCZKxj33j+IQLY7UdfCj0V3WWQ6JlP
wCi0IfKOCunGqhhS6c/F6w5hCNhMb9/HcH+YOtjGCBu2UdKdwuNN81QknN/wflmxdSmaqrHJdbuM
4/xUSBJ0s3Y4FfbNm1pOoCyWhJYYGnQcf88t+N7KoTfrs/VgsIteCcz9WlbUeHuBTInJkfzth5kP
xr4d7l2ex1kagCVnjag//nrVUnTOtWIjWhP+Q53x5sXafKb3pHpLsjdKer05PoAUjfOnFNNUWyOk
33ZmMN6eux6dgZ2WbUAxIQTufFw6LRT+p+gj3xfR5EoLhFwoKiyZP/7GOZYiZbfGlLUPd6TmGqx5
T26MmJl4xGER7/L717q/ZM20fSB5cvsstbtqYDNL1lnaqVKrJXvVhGOtgpT9zf/jQsLQt6Y/IFZz
0BWiJKW7WJeho0HP5CbvXYMIThU6SYnM/MznhHd648I9TFWf+YQ0mCXWlCyXyaLdoyeDYeC3LTDo
FmMBCceE78jtdLyyOl0oj26+c97pBixg6TY2IZQp9qbDDplwvqJVEf3tlkF5zv0eMFvIBkwO2+6C
nujWXs2BRFi7zuqPBaIfaMXY+acYLVkdmYFN9ahOQJXAcjSJjNfT8tk+cf5TTw/S4HENoAc1Q/RI
6b6sL4RJa3HiaclxavZokZZ50OQ6+UpxRSC4pcg0bTOG6wPFGJ4QViLTagjyYa01I4ghs2VHXy3x
JqP/2mg32U2HdykbIeo/ctWLNO0+n7q/+2ilPv737NMszo7Q4ThLR49LEHFqLIyBG7DC4y2agKF1
gsdfgFvh/hPxZbFPvMDnPG4EosqeAIeUwCRySkvrEkXJKp1xo7tYWHyd141ibH6OReY4u/SmSvHB
s7RdjsSRQN/KVLnqPSbVVV5flRUI6Txl1lBJlJq6xlAsiopQDpsJ/lkei7HBFzdV76BYJrwpsLdk
mkEQhKQX3HjwiRLpzGb8vFyhz5AaOPxHcAAJqbx+LdJK7ZYMk9kBoSXSeg4Pa+ALY3N8vb0useAv
oOt4xzWqNjJf4MjjKOwWptvACd5HCDciH5DTMgQhv5YdtAz1Mk2SNnVu+f2XksIpBukFQPL9vtLY
5GRezdQlujowUHdEk+3H0lwAssOQMAJpWbPgB2oe3qyHFITcHn1zduJGTIKe8x5LEUfr4mLN14R+
uvnUOUiUXBYzaF/TPlP6vmqzFEDYvDsEvg4BeugAyHBdzQjlk2kta1XNUkaJehaHjsy0xptppgRU
uZrNsS1QDrydkPpYBXwR8wH4pSsrXirPN3fqMVAgI2kELy03yLjjem6zLelMATzL9E9QIf8u6o0y
UJHRlAo5F6ImlRcZAfIkw1rkNfuA4OVqepPdn2IA57ulrgn+d3ikbDK447rjKO2gBz4EU6MrHoiF
+5TNgOcbyNDVTyTC5gzCtFmxGbAS49MSt031YIH7d2yp12SHXUJUpP5OjrZ0nM+UUC/dui8UBUSI
4ZVVPkoKX10b4jMUX+2Mk0Rof8vh6eXHPT2WX8y65ZJt+JkLOC8Kdn+94Vd9py+texTN0+6voy/f
ScDRmO/dMkKt5iMNxcVvQycGoop6mvsotsmtq4yKSEXdSjbqtb8F5adMx8ZtScz7JLq37PvLg6ki
1ydGtbGL9F4Ks7JfEn//fibdjIQsUCm8osUOuU+8S2uAn/b8+6jphWZ7lv5vIrjL+6qjsbYtinNY
65ZLPNeK5vp0v5eLHm0pCZr6JFQq6Ho8CftSH7+zETOfXgA02fhLCXOCXmSC6rqHXYpcAwz75a51
wEtVPy9sodcV9aID0hz/5TL9OMxvWhqk0tjvNqS+4EoXOz7rv87hGODcLZP8YRzR96fuav93yrOM
P/Gy2CkFuGowxX4W4CzEqQiQ4/rl6m6So8pFiDw2fFmFXXkD9L/ItMKSTaQ8VKfaMWcaAbg/hr2I
jknZ1nGqFjcTQm7WzyoX3vm955Dc4iXM/wjBHDtBmUYp0fonNxJc4L4MWz6ca7VnBEWq1bHGXz59
eQfp9S2me4r+pPyGE39gQHNF2KTKcIUJnwWbxr3KjV0sL0c5znqcBQo9EhqrQWZ/R1BaWMWvxdnA
drD1Qm4lv8aYAgXXnXQlVuKLZhbJYsv4Igz+RkyoMt93fRQTAhm9QaHJKvlBirIrsUloUNggbhfV
cTWpRnnm7ztEzUGeOitfZOkCnyWQPzoB0a36W2uHRKdVlfM4TGG3SqfIJnoeVCHYCt31cOifZkBC
3TqM52zZY1/kde2OxlwNoTJKtkWsx2JCEwhRKNCrMNOv38bAX4licb4aSvyOLpQinjudXI9FKj54
utWoqkFpFIaZgxgX0af/KvBHswdYVQRRtris3duF2uBlIDktqFHrxbedgQdROqkiWWZ1+ACNepyz
Rt7aQX4LqKNi8phqyjWAuR4xZJLRe7cMRmHy1oetWm8AfO7PovRdkAy8pdOwfszvbVQZ7Sky8Xue
91TqTam+PCUBj4rvEcn6PyTURLgabbQhBIZLZ8HpLQbwo3PmCRl5ZEH6TQqAGdwqgE6aVFR1o8y2
dKZOOzMc9ZFGZ5aOcEJgaw/55uNE5LUouX4wGQuFPaZsyCWFCs9V+tqMi13NQZ1J3B9VRHM1nUvi
WRqV8JgEzpS0ahKYlgs/tAd3s2otYd7uijuWbu9Lknj1/XaI9Ttx7b4KAH1IMGBwrPLK6UCf3lk8
QlSUWf4zoupbV2byKaObMTkRM6qA0RbFdW/jJBA2WBKmxQ1KKhso9JBN8WUXWlXNoGYoGxegf+p6
s4NPj38VSud24HTlkwgOCqm4onty/FVb3MqnU7FHjbfg490e4MAsCVLAbMfMHrZnnL9ehlE2XG14
BCVex1gNYsKq8UH8lEr7yNYgWTbj1CViJFbDmhTE4faPtFSFzY5nwJwaBnqDnBtfu10Bdmj08/G7
Btozma44SDZy8E94gSIg+jpD53bBWPZjvTCuoaReOw3LUs8fthES6L4BLUJGkZU5XqnKX8p4NmTy
Vm333fOJ3igDgPmwtxW6qAdxTEVKHRspAXn4Y1us4HXWgjGiWQFCZvkEX5acY8OFHa9rTRNxoESz
11A4gQjswv2BjCGFrROZbtmyW66Sr60GJVBRzkyXSWXmcWeP4QEkwpHpYVMEwS1Jny9aBbrcnrad
m2LLAyCQpixgmUQ9gL0juYjxgnZxtMt3kpQTB6R1rF+W7MoxRaaSkIRZaBE8B/Vo8mb/gwZOhf9R
tGSa8lIb6xZuQ6jSFb40DMosYnD8r4IPwk3WRGBlzStiYEj1Xiq2j62XlsKHBOOeCu3H2cq44Fer
CEQtUxLbBLKGuOCjdWy+YirjuZU+RDg4AHP9njhmxA54m3CI1ZINd35T7MYhlZWAyJYjwBUmu+Y5
erjDZEtg6Z+yyehRjlHsb4cvAEu7BPyYTCXKS7WzaHq+cWPuP0btsWwRkS/po+xHNinlxUVOgaWs
qHlz5TxiiELZw9lVAKfUO9bWzr6ow37MKb591CuqECJfKzM8aSkoqEL5NV8sk2Klv8ZBTnHPw8zl
/BxJfasmhgQuV5CLTjfj3gdLbxBew7ZooBbMGsMamuZDNaVcLn/OpRA5Kyps7VS5eBthxWwYxoHp
pYkkED+Yo++Ycnq7pRm+fkzpbaxj+4khlScrSrEW8qitehuecsXZrkGNQT8aL2eP+/FxiXO3ju0S
FEijvlgXvqKVinoppfLD3/H6PN6zc6XN4YE3/rksa5ioGh7KzyUR+dezCwPMcu8K+Ox+XooSrHZg
j6DfpByoznvyWJHg+KbSQvAJQXZT2y9G/t7iu65HuZNsIFDs3pVsApYr6hLohvz0kzU1vLwCWc1Q
mSq8WK+AkObETZGFiBNyJrkw1ea9I330J6klrKl8AXfl7RU148uR0RoZBwqq6Ncx3SMGacg8vPVV
JlXF2b/8Xj4iKaDyhosLc+xRJt8+WzHTpKFKpQY7F4iKd2vPslDrgV+w5jnwmcIZLx/tas8+rG+q
u6O4zS7u1ROiFO7jtU+C+0baGzPWdRDxj6uq5SDdZNEzdfCKwwo+b+Wu6jGMEdBEFbaV5Z1FBVYQ
6bn0MipKNZK4Q39ZZkD+VZu4CWsQr4dIttczdNEobxWE7ZoKKoXgs8dcZWUFWjuqHGqiPQuPVxQS
xEjrVmt78zFD5Wn7S+AqgTIWCkRQs2GO2a4o8woCg7yYvtp0Moc/cNWabqN8VJPOkkQsNE0Wx3Hg
o8GDcL253ud2y6C5/i/6Ub6HOleYIhuX2zHssqDgWwuHW+ueMDhVwlUzemcpEUwNyZZUkB0u3HWZ
taCZRc+r0R79ZAw8p9sKBhPhqARdv8H89k5A4yDxpxjRJbWvb2U6ohsv3JWVZbBts1ixmLOXjM3k
kFmXsZQI4Uye4MQfYcCsnL/yhRqh6nzFSNp8vH4Nk634RekGFB9d0n131WkcLIrVjR6yQZAZysdG
LRH+siYHJ3NIywicWiGOoA6oR+860jcq/naUUXS1o9gDvRDzg6Z++ZqQRhc26jQIj1SXFSbCQ9+N
Sxok7YiQ246GW44Fef5kMdH23B+tt6e9gZith9YwH5cKBqe4ZX/zA4nRXZPCTf5SOJAAX8dmZ285
JUsUvqaK4o0ga522+TsqNnfjRO0rCmqOOjAXqEAZpwV1dzOOvV227cimT+AiSHttmQA8KdMG8XkM
Ep8Z2v0m/EZ99FR1qaftHY1rNwsqp8Lo34uTd13l926/gA/OV3DTAktr7M8oU2zmJCr5ZDGttI2o
lLGd4mPIAyujqytbbs90WoqZR3NfMGnDjzRNBCLATQVDH3giB9L/ojj2TTx1qQ9sv7uVMwGbBvXF
yV5CLy/vnrCw+6pYqVuW0SkIxS9sCXnf+4WTzEjYdNT4jlhaFRZhZpAplJH5tEm0SO6FsWoUwRKr
tSALAltDu4K3t2ypIq1XcDh6x7RuUucjoUZoiH8ijl85LK0DTiNShWhe6xRmOINhIRubT7jtTjXg
JIYmYSYqpRm8aowIhI7bl4+1/nQYCpUW+ZwtkLfYLStv6WVNuWbD6bUDc+wpnfN2/SlyN1dIYylt
m7a+TgG3icU8IzGLCoP8qlS477+MDxKqGfwobbaYvsQD3SqRkP9swS41ZEWCR/AjtK3LsOeKRt2E
FXBKLHzCFg0dpGAETuv21GKoC77NYTUlGqggSfb32Gq7zaleB+9VoS3vlNP60Rd4fvIsflPKDmbW
X6eyVszmrS07cszM+O9qnT5O6p1ZN89pPW75LZLdQnriqWeGK7lwYa14fbfBSIZmC57tJjciFw8z
BGeLKsRWfqnwBXEHgTz0zn1CtA6XH6MgHWFRbcAjSbXseMcqNc2E1BuFcO+pB2PU8K+42Xvdufc+
Z/CFV74MmqBce1d6RZDxnGTNRl6PVZ6v82+cAoJrDxf5SezpvM1dU1vfIfYvA9W0FDwDK+lUCzxb
Mn0I41XFixcEonF/XWe7pWXqNVoQtqDPGUd0AAR6eTBKZvULGKUUq9whVT5SdrOc2yEfJUsI6rj4
timyWeopGFmiSKWINSO4kY7fWWDd1Ro95vMZ2Gq0Q+lZikw+uZyRYbgPFmb3ERuvuQBE5Kpz/QLz
opq6qc01p/KpjuIVBCQOLvsJV0rA/E9uS1jIB37WY1gDuvukNzh9IIS3w+dPJGUkCuR5Z/jiMxPG
DJPKCq9DrvYQ7cH6Nqrgjvz+oYbYZ6VB2wkU7aW7PmKM+m+gCPr7AS1tRCQ1jdEjlLGkd4GWUXJi
Lw2EQ+U06K80Jg0hGVq380c+4o88769h5W/LoDJei9g51XTOnWJ88TgK7980xuuPVBff1Cxr3sQ8
SQWwaOXxMOGI942WnwkjTNmq+Nh44LeRzGlKY67svn6UFKeErBJYXCnJMLPwrAv/8x8pdZqxrAh1
g+fBZoOEavxJxoXfWIXTqR6tUiCk8ioTf0uQM/WqHBJnZRsdoaiL8GHDlrF0Qk1Gi7538pJvvY7f
kom+9d7lBcSNZ7DJBFe4dclM6u5WxNXWnWKYXOU1J5u06rgdogEyYw0K79D+vYl9kuiuyrR7h3jq
L+PvbaA21taE4G+v9P3S0yX6eV0Vr4KcnpFvKFmlSWyTqg3a1eUFFg1Ytp9A4WL7TNFErhEpJzD5
Uh5HLnb9g/dJjCyCqMi7IxjlCbO6LFnOeL4SKGA/Yn4bxaUVLJXg8gJvlHgm47rgQSu7l5sDqDmu
9Tf56i/7FKy/5a+L/HLHH4ICJ7usde7ch2C7pOE41EGKseTR26g/pKQlLMW6PsT6VHsK0FqAm9hz
Zb7y/lB9g4OQokhM9aU8ud6kkVtvjqZqEyew0PahUdrzJheWBKfwf1poxGuaDuRtJ/lS4nlyP9Mh
sZcxvnxpjMNMqcCMrb4EnmMFW7yPGf26BSPHzgmGt+H3Jpk/gYEGYxFryXDgJj+TLpjBn5ZDMLK5
X83Kj70HwtuNXxmo3K6URYRLnQG8TbaXgG0k8bWeATnMIaggsdtrj0THT+rpM31KhiHrRbcP449W
i7zmNik48NETNrRQjwegT7fWNjS1knmv2VGCWkq0kFi8rAhoL9uibTis5XJ9p9ae2lQycUMgZT+9
uG+xT7xtrGhcevdRqSmbbRnZHg3++8L35l6ZJ2L5obXU79yXJKf4i+567oe9HEII0YYO74rqLNWI
Me0gMp/gErnl9c9dnIHLVggKMizCsOLKiBkcBeL2rjMqOZXqyUgqhaIWZB4duINx1AQnA7lxmzZr
/weiKqGZud2KM9udnRFCGfwkbrRpMO9fcdUzO3TVIv1SZ3HAOYXRd9Dkf7rBhHbckhcoSBRvSSbZ
5Rpnf9dAU3JCAnWfrsSFYCq+1+Yoto2M1G70rCRQIbkwQeVJg94Xtw5ELyM3KycNfvFsTs9+d+4v
nY5IgGCcafG1DNqLvVFvXAl3IDp0KjLfL4j6aK/oH6fwLtxCcbsaSRrrxbeEJaVWr5w54O3IVfHe
F9utYLo8VQZf8g16ltHDTweufSAVT14JQ5xWXonTzjcTha8VmlUhTr3iIzpUxYpsCAbjumPFvZPA
MazgQIrn+vWCmA/QRHiPUpdOZBSune+rTlX3vDLiiQ94oA4n/pjZzEASu/2+FVAN/rZpGE4garQX
XeeQPPrlHJFI5VGL4eHz7fJlovmjOppfTP5XoGj4Ys1Xt6Xhu60i8hW784IisyvA7rYSZaA9J9pp
es0/6lFrh32+VdClDYrJrgHmmYEJ16LHFhDusAV6bcQ/+vFz4rliDJo3dbzuMkvA8xaf4sk9HLZl
NkCJF3SWb9mmFch+2VRMyUYzSlTX+W9dBos1doNZIJDoOk5REh67At/ZLQGxLZyBO+oRCyZfLoAC
7eyk8rm+327FL24d8WUTe6dZ8WnXEKJOhwrpq7mbbWWYSEZzFzYzH0J0Qf2rFvhd4l4CddJBWMQL
4GJ0vT7V4EER8MeloFdu08TqtnWii18InarIaE92nwLn/wn73i4Mk9HOqc4fBmQu10NVQQOiU1s7
/RW8aK5tK++Tb6CnBjAqeCwGI+RH7slylPCZVf3BhMh/6UEllNzwu6Jd5tZR+HH5wgkko2UYRoTG
29QvHxSPb9Ss7R/kpbIaJXD7uBtLwXGYbYab9XZ14rLBMWUQyblR8uXRTDh8cF69sWLG2/14OWAv
5gub48epXqoZIrC5lunBtb9rlYnZhijMfyykAM67b8DLyHBd9MWtm6CF8ia2V8jlpk/GdxImqa+j
aRjJd3au3yVRItDCIhV8zm5dWsuc/ZQXL0inkDu6/6UJgXhNTRLUjbdh2fzUH7wFzT6iJsIlHyvx
cZD/nIQ87u2xzArZ0D9j+F5JbodCkwtdNOvpjshynq7jFs3vkcl0I3BBxJTAksGvBRJ+/txijksp
br3YfAypx5ob+zcp4ypUGN13AyvgiKgV3/uCRgzlwfRLO7gcE5w35lzS2k/PqUSwharVhNNnH877
xj4ZQJFFcUHf3KBOhsNszpmRsUJ3mutWxJQMvLd8nvMd7TLba96ENwSNLeyp3GdI1wCMwE5uzNdA
psKLrJzR143PXAvf+cDXwFlUEE3m/Km3qcKJlYHcKc/9/bcLJ0h6UboLyUbSxO+hzge6flzlFVHZ
Z72EZPAd8vacB1OtfT1M82j7WSwdBag1oI9CZQq5hJrUTjAs/poTHfwpKnyRIzCT5QGwI9geLAnn
A/s5KCpvDE0KZ+S8LjtkMVHclGYWJI9ifkpzye0Yc+/a2s6RMFP29NzyTUOBL+09WzPUKlw6eNx/
mEFeKv3pcJbh3ncCwBnusGyuYduvjHIFHphGvT0hWQ0c5nD/ckp1f+D4sR5SIDRFbpVkqbq03xlC
e5dSRWq+DHQkI+AgC4G1TPwxVi9OX6DCfxZECM5UE4nogpGwWBLHhGuVLdE5miveM2Rnm7vCkXdU
cJcSbvMEC+zRw/YL6TR3vNMhIoDURBYAjLY+IKLGjGXpb4wCrU8wR+aBWfn4Ver9yoBJ9WwlHzrD
8iI+LLkuMOWjWhpNh9AlMJRVy6IHzK1nTXD/1Ruw4YFLVhz1UsnBAf9iM9UR2o+aQ0AlVAbvd9Co
njd5o0xisKhDRqW9kqingU76PVq7B4JqZAIsrKTYrjYGSMRn5jrZu6nnF7rgUe/LvGrwIiq2sp5Q
ylrtvtktdYQ7U5iNHsgsUqCNt7XQ/5ruHe6eO2E7tp+XFDHzaglXSpBWDBqoGWh6G8TY8lSdsQtP
ZcQYHGrkmbghs2rEnth6jK1KTBUCVrEsdgE5kdGfXeBboIjnukXFbhAavTlPoi7jUyHwFa5hOgv+
okLKbIjRsuhecS11jJG1hPAz3C7FjF8ulON7Ipq5AYLiPMxOGlvtLcKkQ5nf2FkbCIW6mnpBSQAM
G2p1qqbf63tfe3CH9gjWKaB22Zw0G/TFJGnqYSX/YdTPGH7ZNdbTYIUSF4n6h6dGa+BCX+Yd5NGp
TITbV6zeTSqjRHRjngHQNOzQcPs2Kwzyr5h894iANm0vRktDWTKQe1UqcUcAMNmsZY9VGROQUlYB
9Gt7CS88hNG+gl+qYyCVWr1mFrgrLm+39TlcaJOfrSkGAat6tFHarJgF7GO4B+uIgu1mQZZYThpx
UwLa+deIl2oebozQNpNGZEB3wX9hzrRz+frmYxwp4GMeBkcwINPNOQtPkptC0blt7CEAkiwtU/L8
02vLN185IAVp0uUESQluOFgwsMWWE+7TZDhy55qohy1/UreuF72GuHPpDBb59chaMuhP+k8uAF0F
GGiumJV3sXQBYsQRjgGj+EQ9oeN0v1A8VVZIS3yBNeLOOAejjkD0gRkRPc7w5RhdTtzEMu10T9+o
3RL9AKbXkQbMG1uDqCLBIhQJGcfgCJmPpcRopCr6VuA/T3LaeY10p5cxMLWJQ0wniKlJkdN9jr5G
xJSSh86wmQ6eXXDdMndTMEb4S+efyNzfTn82Nu4ZkJ+yKbeYsJqmerPzICZDklR1kIPyuyRsU+3y
CTgkYfl5zS86W3wguaDJEb2qdpAwtB3nHDsOxybtuRKrBNhhXbdOM1BS/yQmY0/A48kNyFAcMapp
t83EYq2qa6BF7XgmCt5mTtwx33TkRwaDkKVyvXThFhJkhpG9OMw06/JWmVf6+LH+5PiKVKEiJcca
uhC2OX/47ZRITko4Zmk2LW6DXQnoBfrmUVbITVLu2948T+/xNaFpOWhfHp2p4yJWKEevSREf7vKb
Nrkrtx1pAkXXs88hq7tSOu28gad1DDyF/yLbCt2XB+RlFvvLKhRmU+GFy0CIf2fapF5TRWnKqeSR
3A7XIeuEaYnenzJStOZrdvnpVNttJ6FvwvYx2puvaHcWu1OWOt1beEYHvuWT8PU+ZHA3IwqGZ42W
JlnGQGsq9Rt39PxMfp8y/pXv3TdP4B1JQtg8iUCmUmsArckydM1xcbluZPeIB3A/pKYeCX10TMqt
tGt+zlc8PjWUpbHJFW5qwVEpjsHt9Ry+J71ev9IjtoeCDMkWbjaX3ZlqDQY2SGd+vVvO8uHf6Vzi
faZMC0tYVmQ8hr4E7OM4O/jH9cQ7rjEIRh2k4lunivTa9sgqxUNzVSd9bEuH9MppGlReDQZ0Ua19
MW+9FQNAVx6xCqJROqHxDyBODUC05R1r8jXPB9D2qWaUNMApcPf3OdsNU90WcS5+cO3LkqvViea2
5epM5022XSSI9mf5rO1UjFgwz4DOn+m6y4l7JoD6JaJWG0Zss25wJ7rfkAjVZ97G+fATS4XDTnvW
P+TFU7mMDxS0SH6ZmQJ9A2jgHFe5Q+CrqJ5azX1AlbVPeGW/dodAQZxFhRmNKHnhBT82M/Brq1O2
b1KZYlYL1476xpuDtuUCgB3JTagPdMle3Va/Kw5TpIZGLkCCjfaSVYe9WGWb7raRI3ol3+ZYJpzT
J4+7eh0/ChSz3BwpWbYWcPUON7eTb1sxNgXpkPJaRC6DkwLxtoWBy+G0rVmybRlM/IK1vc+mtQfX
MV4DFog//pn5yiG7RVOyBnwxlhzKxrv12+4ZLjHG0saAWbNN3cTzmicwqxB9taG2uZB79dJqTuYT
KBt3tndDwQkGoNZx26X7znT5M899/3IAzgM29aWB33uWgdJ7uBd02v+Um0tBssCbEqaQSPuH21UF
WdKoEPqrpdAA2wz/WwsltlDr3P+LPmLhrt/FHiVk+wu9neyb7jUBbmbu/ptj135Rh5PcTqvstywL
K59Yh1qXIb8RJfV2QC/PkbQEYdyhp0RqaYaX9G9FfkRWY2YaupjelXbwgjbN727kz+pkrIrYvQ3r
V0vByMfd7Z1mw95anx6JdJ/W4HfH6/kC1hHryAgHO1gcDbNPz7jr+6nQhjx6Zq6zrHJg+VcsZypJ
bc5QBWYi33r80eVCKS1j3zscmFONpfNA8AvjMeaDDRSKIzSxMNoifY8vcNDEroBOM2lutZ1ywp8R
9pzwKgpn191uZXLkHF2bgHtmKLwfUXQCxvvlFbbXoxMZuaHjSscRS6207+LpdeZQ7ETag7/ncnQi
6+/yCEIMGH/M6klD2E4d3idLdLRUJfoIZJsgPyBPvTcFs2SLfUkG1/bFHoOAV0fApfa9qfxRl3Vc
32sZXViuTT/d/MAJnhZHnpqIvdKouBLJGT3dPr06tvZQVs3IzRgAigOm4Nx939Fq00e/KrIqUAhY
6A/mvfpmGb3R0aMP3QZ/53trlcBZWg9SXLcWbg6rBLt49sgkBpo1WDrbG3gLYbm7yuvSJLKg87lb
pcpjLrj8hiWSW9nYwWLvFvG3ILOJ6e5I5wu6Yf5ZDZukI5jOGMDpDsbyr5EWESxJnooDXgA4sk3j
S/CvxW3tfMeUKZp0YFb+7C9Yrk+sRqaKu+jrsLauqr7P9kG9C/ek62oG8SxLe8pTZftEwhfJ731l
cxQk2w2G6eLGWIuhrq563FbWDyCev2LJWutcXCrtHyC4DOQ2ZLtlW6CFrDnViu85fEHYjKD3L4Zc
eK75QQiRskRPXAf7d6D6uHdkUorBu53iimpSjlR6Lx7r3d1s/f5yZthtqM/Vx44vkX4d0OpdwBmS
Aevhki4T9oMoWHL2jeC/9++OL2BIOZ8XOP5hYo/XN7/AZXCHIP0+Q5cXIFLiAwNTBvb0+mrVYtcR
/W8pYlOhQ1z5YiSd866Yh/T92vDCrRMEjVcAZENWOqlqvlN/UtycOmeHJsOvtjeX6SVASbA/g15e
KHAfuxMZiFt3qfN54qREcxO+r4mfrnck2MKeZOePdYe3GpsR+54hLBEsLDkH6+0x85kd61vVo4oS
UhhYRM3msXoDJAOs7zDm9ZbmDBJEbk5FDM+eqGsouiBPtuHHpxGM1qUHdFVtfZVwbpk/fnRBevQq
/8a7RewLHbFf2FtMtGpuSuBotS5ei2HIZKNsAPHdopZEzAVZ1W1+Hr5klGjl6x8AAb5sEuugGVIF
5ULIaikNz1NumkKoSKAIbBGRV+A+FRdVXxnZU16CGcvmYOxUwqK1vptsHrTER3poxbdslhXlJQYA
rhA03zoOENN2QacSV5jzJkzqYrRwUZDNApMTDKgwYMXX12kqgHx2Gww/f1g/mhygFmInkjzKDUSh
4WlqkB+hFUtPV5UJJ0WRo3nSLBzCJTim9E2Aaq48yUbNcOsgP70f8SjWYaqiwxxktzQh7Uawanzg
rFMmbB2HzdyZuyJiyx/nl19m/T46FMA0EL+ToMjGTFgmvHAPucRYQPrSfRiSUPiTvVcIswof6ehF
T8uyR3tf8OXKNrJxLK+FuIxTIkOyil+OivV1af/Lb2hUVhAFRPN0Kl3h0+AXoDGC4CZnYe+72aEg
K4qlf2Ztsi0oet9s1Er21eIRflG1M3zO7gbNhHP/9myxc780Ay4uIMidBQ1fEMCyXq3J6+lOyYjV
+vjJtpaPdTBSP50zNBgzy8WoGuWdHenJxMRJnE+6GZpgytWV5lTf94hFI9BOvLfM0utqIGv+h0ET
BA+P67Y/k1FbaEXPCAUry1DYv5TEtxl6Dq4BZbQEUNnTzXm+j+EiLFJlPCexaeueUPxThuFEVpQJ
UIPUWay6rvy6w41oMuMXe8M2nQ+7Oln+7AXsLd6vT2IFlXlhNPGsS2JKDafLHI9r6ZtAfg9gcb6D
c1fM6TSN8jaZBpdQVRW0W2g3Nyo+ZvssIt9OUCZpr1CE3UkjXpz9/Ha19M2CmyIJ0+ReW/fp3aoQ
jDRc2koJfWAAIaxIJCAewmMX2AQzOdP0aYTOUPF94f4nAn7CecSUunlkK1IaP2nCRjhjzNY3WD9s
9Hl1txaURBy3abuHpVyB81DYVGRqIRkZwb70y8M2NfMeFyvHKt9e3N9TqxDGWE48Z+VisXbGt4Sq
F5bI+HWZATlDyBq7YkYmgyzug8MgOtQvCi3KigKLX8XdoXVVagWUQmDi2uqaLJEruv9emxttxivu
cJuI7KNpcSXoZpY/gU6dzNQ9I9y05XqWLG6cVyPa16zihc4uJJaH5XFqhbepD5frflkQ5o7f4caF
R1sxa6hj5hoGXK+fi1XAihhaEUMdezUUUcVtb9ocP8e6aKDo4MZhCz63ASyocAVmxATUIp8Hjai6
BN8UPBOcRHAeAhGqW8LXNusUHuvRzpiS6Bhm5GNXENf+PytB/n3rhaG1mkSecs4p0M6PQUTTBBhY
YSggjw16V7J+sm0em6/algULadUYch82gPIjTtxR4ZEzuGKOuWRdPO/ue2OJScbaKQ2HfJ2J0OAW
vgHVZqRSuyEjxj8NYRD12RC9WUoXFYHU8ra8sFBDGRg4gyTakfFg36LMgbJ+zgTF5jHcpZDvxZNk
zAmmxDpPF2mrlzc3aZ3ubrZD+KQXrrL24jj75C8rSkd278D4JijdagTNduKy5tYpzYZn9hzSi74y
5DDx4nJ3dgCkOb5l7nsFQ3KXzHMV29Ts9PEkE3ne+toZGgGrpe9T/49qsiK4qSIMOIUL0oZvBfpN
FkiWxWHU9NzjFiU0mUepavRWRvKO1mpqcbXlai0wzb10ZCC6KSkgqbidEnp0jL1TLrF63dO88wQi
bDcvkbsUDdqMWQYxQwMSStZf9Lo14lOIqQcBpBr6l0TMOguvS/q4crN2mz6dJdH1smUhy9DY/Vdp
EQJMw10wF+nbfS5dMT7T1XwlwPy1q+YPXX9lLSu5Yx9h0EAJYMMM7KS9YJl827wfQ+zfDU2dluKq
JrwyCBUOQRhKqV2HWMO4pLWivqKLomFW+ejX8z7QA/m0AoW3JWqJZ/+BLWweS8qkK5ei/E0UY/0u
FEji5SsYcpgdF7O2S4fWKtY6zZChb7LWG1wuWE5dmKbplJLowC27RJlkkLJ5X8I7/vYK82Vq8h3y
rHZ2JPmJh8BhNqMLXPcSp/d3/jolJE6afajZ2ZgSOSyqLiAEAQrJWGci4TERdYSxXRMLcJlznpgN
n5aj/JM0gRmvEgxsh3fae/Kd7ttPIE8lwSe01x+kSJRvn7h6GewoSh3jKhDTxF1ysJuG/obcjb5z
OBxpFpnX2S69xVkeL1QfwBfCRkYevV+zWhW2cyxKbO+m1E+56a4X/xyZbMNcp6n0MX2pf+HfKsZY
DQqNiJtKWSOQPIy73Wm+ZTbxPIiq+ViLa1b27BDk4+Q5KfuUEbSGkjvhJ/qMqX1T3wX1o3cDv9q4
C6tmMpWj6c9C7bY4foWFFF29+2YcCM8MqeX4rofu0UB1udB/yI+nFp71sxuhhQ8G4u7RpWuEYt6p
TfPH7T2Po7rVNulqYndjxhvPvXMEbgoIWeSbFHshZICF12b9AUwaA149beqc5+HNFD22Uaoy2JZ8
yXLZoqYlXZWXbviwLhVoyhFOc3Yv4OXy+fFplM8hwGA2yZOEdHnMnh3iI38P58x6kw3Sij51czs6
JlNCqucfsnCDLxktw+sezBO7cXbamFpKUT7RXwEAO9dDnHMYqz5NvamgHKExBLKXrGCstPGkNs7L
0X969q5QYkR/eTRRa8hEECJxMBpedX13sxpSodmyOThiTxeYhQAzHYZHn1SdsO2rfnRbzA6L/zIF
j6eAZVovwktwnDeJK3wHmmCU8tRA8/Zyz8mA6hRF8BNfOtdF3MWHbIEyoIAeZso3mdTlZYcljtnk
xfKidG+yPbhKjcas5YLTlW5wQXGYpOw+UiaG3xGbIwRD9+KLGZLrGMk9d93Nho7KBeGHVna1kIPy
t9F0EFRqqt8lL9F+IyBzKoLJyWnaSGzw9LvRJ7mdMSkyRouurAAa9VAM+mm4w9tbKBNzhi6bgoxg
mr/AV4mFSVP+t7tOpNzx2gUhD5IAvpXqOjf++Hdt0fExiC6NircR0FWUNWf1cEI4qIWdDACiHLjJ
Nc9YaVO0eL4G4EGbWeRQgdjNs0hch4DvHE1Pv9A9j452FzpxcpHcceTyugZQENiw1U0P2Ri5JnuC
UK3LWMRNo+I5h6V15Kp6Cssve1ZS715Lr6iJqJyZE0Olde/0FrRCmyFYbWeWtqe/sjOyPxNfQhgj
1HbnF/XfizY7mTP/BiVouyeFaTO0ZfCysYLav2vCzwDlfeSSM5RdWgTpNv5S9KWHlv+C7WZv7wEJ
Evmz0QGvUD7JQGV54uoXZ/SWNZtfThyYfyZv0w2iKcdgHSb8CmLbCuMp4MLQ1TWV7hlQCarxhkY8
6o2s/TC1U+tS90fCuPCc9hEYWreqNJrKZzpYsCQnkz0/YjS+CWfM8wrPW9KgxAm0JNg9BMNZ/qB9
GBpwpMh1Ntec1d06ysvs7VodGJOHNvQTp0kFRahvu4sDnkotFf8uReI97+6bSYOKlWAHe+euVlOU
5pPUGRl+Jf64Wacjcw6ozJtm+YHrmm+Gtq+OvGwNO54dcww5VgV6y219zW+FIVRb8FH9N64SZ+N9
RTHq+6QRDJi5iOLSmFAkF8SaEZyMbCAUn9G3OOhB4eNK0dXMiiuFrcUW2SLcFlLz7Xri73KxUquY
GsJHFPhNHaHDcjsYtibE0ioOoCxP+pDwLpTCXUUfJZ9fR+M8c85dDyr+giZeSvjpVq51/wWfAI8K
POXne8es/DSkvfyd/gaxoasfEtie6ygFAEis5bkk7BC+lSB7i6GgmS1+aWvdjff16UZ/gU+RBpt6
Edc53fHkTrKNwFWbb/GzHwVjlZR/EIW3T2g7brMF3fTG/eaBMJ75LFl+CU9l12VtKSwHcNV1TVoT
JcsP5BEnJGPrl6FKsEDMGEnIa5ULjCoTdIweqKu/uulXJnEVFGNJp6LIl/3ml3ZcbWjVLvK8OctW
E18LQDHbvi3EuxeKCIDDxQgL7Gms+gZBsCDsvzNT1pbtymsRCVJgiDmxKdYWiwOmkU1pezbXid8d
kBu/AASEbaDysZq9MNq8P5biM8gjDbQRqgDEZF4FP7lGQD5ZcSenNXr5kH3MKgUVWPRuIpl3xrgg
poEk6TGJH6/qImO2/c6wBgmNpZwGjDEnBfYiYOWkA/8vjyXQNdj1647rhsvGXRXP2AlVVHTk5/kA
5Np7VLjehoW7R8tJLUEfd0Zrju++I32OKRdVm37m44poXGKK1+2ELZXKcg2Y0fgxAIQSCbo83WZ/
uNdnqOb72OzBM4EBob0IRQM//ElX56Jgfj1iTdtlRP6suUJ7NOmOFe1TPI8p3NxkyFH4l1CQgA2f
P/OjXRF+zU7zxqhuLI5Yb9a3GBEdMW3IKafm9Bpsa5QKHNnKtfj29ucbclylozsC1vuImRHmgryX
HIzC4FktLiu/DNQ730QPo0JTyHz5VdHv0p13M944T2nYaT7rys1ZffEwZMo0HUW63vuB5b45Vzfm
w4z0a8GB7rgsPJ0/SG09g+hvZfOJj+ay0uf5cAI0+wOOp4Nxy2ozgdf+QbvM53U3QhvKs8ie+rb8
gwq691pMRjoirNZLxbGEn6WwB7csdbh97jIO5rEBqF0sly/dmynFVy0qPO/m75jd99aiJCUHiOPX
DLp9MNSZDSs8liSpj/5wSUx0lDUDWcToFphKhnchAvkGnVvtM8S3qGgI+MNZwKXw5+E6NSE+gNlt
GjTsWowr3hLMq9bsVqrEfg56GhRJM6GTSt1LZ5KoVV7WiMwYLhKS2/5jiGmj6Zq9qHudSz/z3ev/
OByZzx00oogASkutv9Nt/bfRpqDqxWApJc+pZ7lSay3r7Fr03cMAcIqAdzD7O4Ge3erQzTbmOA9v
WjenqNgRWls5dw+EuSe13nxZjAsjIng7BpaLQjRgFJWj5htesH84JTfFu3sTzOeRSObW6tspoM4q
tC4Czfe85QWnSUkHrg73qoSkMnznTjXFz54sxEmFP1Iy9QgPAILA/N9iFsOiip04F/hc0Gkt0YQy
dwY3+X+sEwturGqFyqvBccv4KhSHsJ5U8wQGnhKXvhjxfsx3AnrpQYKvOsVCAX2Rsa1QIKVKTX/e
wgJ8bdK2PGbw76v1ZeoRMvL/8qfnRb92Qn3BM2zhLfYf4433zbg/Nbkj95e7UzYSic4IUNHr0SGD
WdDz/c5Foe45MDJH8YDS1GqZWt/JXbvXPiJ7y+2gWQYowoO5KStlk3aRC+7pgAVduYWczLEIscHV
/iNKpaSIEnbtGNVnpwSiAsV/F6qpfvgJqsIDxmHLBv622bA4O9NWSHrAkSMeLAi6zeruNvJPiRa2
fcvvAd0vsl45jvnTxCcDPrHDVJIR4oGde+vPTHeUc8LaOg4MOAnD7f144jONAa3vUgHNPraWFAf9
zgoK6VlengV3rHRwGshrWdECv1V1J4a+P2QV0gFy7ZfaECERseHsFME69le29kQ+WnmxRsCww/oR
kMemHgB2iYz65Xkawqt6aVXSsGTI+b7kQG2HphB7gu/SlX/cyUDyS0U8MjXi1VDKIqXRd9Ot4utJ
DYSExO8wTKZPB80clwEgcOZnJ7JU1zarUQnCFXYZfbjBiBoVs29ju5D/MWSt0yu8Wa2uoaYwqwY7
QfvoswOpAMuc1ZVxIk5iJaosBEJSnlaqsQ8GQqAypnFHe2f6OCFLlsf0wpC5hxDyOgCwIyyFgX4/
pcDw7VNB3MhjsIIJ4S0ybafYM90UVOYshfY96Fc1qapRJPBonSGe55cPwgEuWzk9D6PdJOFFSS/w
zJYmrzqbyfKpFTCK+UIC2J4dt4ZQLkaFAZz+UyYIaG+qlU/s4DugD5GwwlFpOherw741mnwJIDUw
FJ2j8IFtaAwQw6IhWMHI4x2LwJPbL+TbrwmP3Jhuir0mgkYhUcKXHTf79G1Kdj0P7TvC0pZxeios
/lXes461PnliA4jdQWrrOFZRxiZIUiMEnJrJxRcYmFXa/s8rDt96un/1EnVBit9CmJPgkFQBJIpj
l2vPkbcFCLG9dhXkrvCEqZBZUHWqORHRNtNpU+fnW/ZnvTSCmvMUbKfntWtEou7Ww9/V2qyVDPFI
o351bt0XeKHSO62hryOE05H+Wpgfcx0FmMrk13Oh2f2uHxyZFtGBpKwh8WwyTXpSawuUHm2Ng6ld
vBhonn/MOrxgTU6DBQPEuEeOol5MTdoefpxTQy8x/HNxHQ54lK2U5Tphmn2jytEjg7NMUzYTxlgV
fll1VssLpv2kf5JidzfHWfXLF6XYRgguILXuh105nCsBJARVLcRSIwnBt4pgC/BsEuEASnBc9IrS
eZCW5clPO8JaM7lDFBstNWrGMMCTRPMUw3Wx+pJ6WcBt9/gfXYdYJU85MRyMacysazgVRmpqULX3
0ODwJ8DtGpKKz03LZqCnMOhDjsppBirAZtO1NOlaakbEmeslNs9Pq62IKelZRh0vSm0KiJNMpAMx
UPjZ4SHjA1ggE8mnmBcKGpOf3Kl99f1F9XiRC+OY61cFPyN9qPXFVX7JKXZpOfsde9CNwzmYpNG5
YsCwHxyVPhjna0Z2zBkgnMn6YKc++S+269nBRRbOHVZgWuHGmLgMmWhG2gDNtu+gaGznNTgc8VbU
c6lWnMXfXpTZ3cFmmRii6mvtz7iMX6a1Nkp2kJ7bh06gsRudn+5w4aW2QfRv3phu8clSEoDQiGxE
2yCLM130IgGvRv2hr2+f06OrgtwPxTc1rI7L1ankFQnzyGKQEfLlthfnIHeFG0pJDTrYGwJiXKNt
GOhzN8oPpld/XkO+6cU8dnqWrTQcvRppV2yvhvdBXwm/rn4K8Yn5YXdJDtB67T1Z+7KmDLW16T/M
F0whWAR4vpLMDI5zzEghhsrEuUBl6jaOh3t9y48oPJ3WqcuNhB9eEq6hrxMxj//vUxKLS1Ap0Ans
4Cnrig6Q5NNZMuTeMRcX4YQlhSRooauiKvHvSwFV4kcJaGPVnc6Ww1pEfJgEHXZnKNRETiH/ian4
V+xoeZaPk43yG5uScWQkI3+2M2u0mLCiVrBXXkt205KSVCEt+vUDptKqgcjUXYqCApH+5sk2kvdX
z3h7kXB3JG+ooU5iKS7w1ka52N3rDiMkOTugy89l2fYpEDOt3OL/lyycolrm0R42QKWgPOMirZj+
gbvzDkEaDB0xm5TgblM+ZZgzwDhTRxDskrYcLRQG8edIh+QJws08T9rV1TLePb9hXFci2H9VrIo3
dkNU7kunOvXktKeZNC67XEdFQowKD5gxurW4KHqV3eLkKGNVmFMWcvJbVzn2XkiIsbd7wb6yLA6K
IVKvDrrJ5w0fjWLE+3gMQmtyGl1HYZLYgcN1CoY6KCpkres6AOfICiv4o4MIU36ef9qsg0BHe6v2
IcDwZQ/9b+qI86rT2xdG8dg93JxsOuBrNVlJAvJdRpf+R66MZCJ7DqeCfM77W1SU3Ozw7BfwmdPp
gEiwYVD0eHysyQThzSMU6QiYlNW8dPxnYDJo/2Y9mXnQFxheYD3W9dCVNJRrghfXRUba3Uh6zNMi
h1UWWkLOUVOTJr0fUQn4WrSiRLFMC/k1clHolP4fgZtFzBgZ0f30OgzL8exOSF26m9rO2IUQD+Ga
yTcgssWD6evdyzNFwnbIYMPGlFX7tu4YdiTqH2NAMdHMoTxg8hSBlvsJH4KZ8Yog4+38+7IQxXGK
hCrQPI0KUaXFttx5TuDnnSqS4ZLKLpF7EDdlcLzAAlYdfBHSbGqOqtv74+WRL3r5ofJBnrJDrUXj
FsBI1mFLS3NoCsxy7zv6dk9LKibGqKEQN5oNRNmixyjgHXqSpzn+kxU86b4uvIDtWp8kVJP7JFhS
mZn2SL2dT5mPXlegTPmBjCkGII+2s+AQDY/CFdfoN1TMwfkjlWhMr/bmRj4wI+R8cexk0poLhJ3v
VbGverc/OEPSCougw8G3Sd3pP/tRQg3QbI2XgUEnLuxj1AU6zGAEuI4RlTVZrnE8l6J9eUqyc9wS
HKre/zwupOgnI5n4RG/pJexdiqjaDtXRH3xR9Cu6DZbTwJCJdeKKuVY5ud50FB9RnSZ7Gc8OQ30b
1QMyD3R+ySBbmJV7UGUK4Hul68j2L2ndvLQzjzUzCPCaPKh6by05xLkfDJuSVj3zUOGHvII89uec
jOao88Agqk/cgFnrPhf1QfC71OgNQCs/bHUqK9q8Ver29mBRnCPOv0qix6XtJqpgR268fL1i2bSy
9s46XtoCRmdW7YzuSzrUVQBrBo6MMoY/oyB6y2lyjAFCzG2R2WOhZ8RgAgfIlHqkAXkTZalF00ZN
qqzOxi2R+c1Wm/dKKyahraAZESbSC8QGCvb0ULT/pR5DYSSSZV6kbvz7lDNGnXUlsSryVDnC4lHt
UeEd/6w4CqpUmquKVrv3QcbAuP7+92QRTLyZCLkqey1CMPP2v2lX/nYC9x+cOjID1VchYMK32ErY
8Ws5pL1Pb4GcbLQ9glNAk70VIc1mZpZfhcgihfJzJ2gC3EoZ9EXcfujufRABic4AQA92R1KWAq6W
VnIGGQCtUJWvLGez8kEyszMPPkVDR03XDz9g+f+Fc9++GfEmzGLa60UsT36NlrtYeLKqiCVbX2Bh
KPptRUxxNEtqUDUK5uhiDL1jSaSgEYASbIstdLc78wqSGrKovomkk29BvLzFcyQ99aTDaS4JkOlv
QNPEyd8JEAZuZSsR2HpLdBPAmMKo5LvuMQM+wpfRvoeeCy0vqSoA5NkpVqxiDW1p3s9OeBk6ZlZx
pwTC3pTgyqwz5HnttRbVcNJHUVirfi4b2xS4MrOLyMzLhL5+R7akXLqSVzvtUQRXZ2XSC6TnNYk7
Sc5nwgYAcUCyVbClajwJ0g/fFfyP2cwxzX3W4b8xLI7Y1Vyfg0RDiykYSFimtcqiSlD5P7H+pCrl
/FmchtD2ZiW3OBwp2r1RTMLCdq0/6IpdsjGtRkDyufYF6+cAvVgF2XHaS+TBnL4jQqG8TVpcHNLl
Mq/vw39TbYCtnor5q56c1THw/0ZYbLg11glajlFJmAMWQYNuQr8R8BACD5BBaQQ8KUWW3klu8NXb
J/ccLLObXZfDDj956NJikhWHU4iGvXRRog0QXW0dX0DEjvmqVhso0pSNZnTu9eNjIdz4MAKubRK2
fRzk49U8PdMYYCNPS/r/Wqx92pJhfIv1/s/L8B1yySiOirDYxrsCp8ep2vmjat7DP2EMwO8yxh0x
rohHCk9i1zEr/nF67szNWfFFW2Vccv/9kzONCxOvr7T832jCuGbjNB4L7pLeiuJPnynODLNH8Pri
GMyMrB483PcisXL6jesXDUZXy9UZ6eymwFRfS1+JFjJ3g2jWKSEcetRx5cYB4+lJ9qO8bY0hKKAg
v20CSvXelkXdD8IJIK/HlcZJUVXEyF0Wz1eZEcoU2c8SbAdE8XQWzNNp/RV2Y6ZI8fPVyDt3DtEU
QVAdmPJN3FPpSK4mSYf/+xVVo6OtnxQEdFsYUxPWim8Wti1S5vX9oynNOSDzuJ4FVXabSZ+AF+dM
GLab3DCzikzqi27lR60JGm7SlSC3NXz3ZOQrWWBCkqZMOO8C60Isi4CAZcT5MEgpDx0DEeRrkHJF
v9YQsyrmD2wuLKMvgjO71j1wWOKN3gBzlHPmlwU5cYHTvhxebHDV7GvD/T1J6/0En6UNprExyPie
6f/KVyVGdVHbyveICpQsbIRNkjCZlqVBmAxjExm+k5hiM+Tn19LnuZwi6QbxSZQTJBfmDFl8kqVK
TJa8lygYg7Ti/Y3+miH40zAiDnD3xWwSMRRjSrrqwxC7p+fgPmOFMwIBUKbKX1YCXfgCJmIWLiZQ
joPHqjlOQN0LbNc5TKvZ5nxTtgXHqmsUtaI30MI5E2Su8DEY69pyDEOTpEphcTeMH8VVs5ZMeP8P
XICkjFxl9kpAx8By/taiyONdOMin1hRq0QMwLP8u8eb758synvjhs2h4jk8rnlzttcF1FsHWM6ug
JavC5eArp7hHzZ63H0iLHlcFUJq2FMB2dV+q0UzU6qwBwFPqgBVBnDguWhDird/9LLStS6hd+ZA1
qiOI3HzHoRo0dUYDp+2Qk7FvdIcsQ1WwMdBjVNaadmgSqAPPVlCjl/WkDxwi7mUGi/MvhnenuhTd
EoVbMh5fX2aUjTAPC+x1E+bZCtVn13kEVzlietMSM550HimrQ1ZV2VWxjiP2CsCfVxSU96UPmw1C
278MX8XqjP/jI/+330EOUe06wsLICtfcm/e0BtHm+Rc3U58G1rDNhKwJAwW1QfxpgvaUwL8awRvz
xT7Si4X3RH4CGa5v7LF0A+TssSrFO4Kj3umQxTRd57a3vkeAqPK7NkaW95uPbmz0LzWG1dR9OJGR
es9DKp2o1fIzT4pQQOn8zFrT2OFsuX9vU4FnhwukGm/AwkpsRW1RnWuMywgqKADdrm1AQjq4/J6P
wDSRBeXS7YI+niwqfNCsASzXW4kFDiyKfdpZc7rrcIpfI50gcMcSEorWCb+G9SxvQOx5x6D4wo7S
DQXYdwTsjqqlBIaREJodQG+eV3MmDxVx1lAcnko0+PRqyh2h+cB6fYXQYeFdRWV9DIe2XkRA0U5m
9bnxbgIK0RojdYoeTjtpU14t5D1DuqKxIZWqiIxeREmicA20zong6wPWuIPPvxKjmcx4J8H/snYy
oQixEnhKTMwFAMBfXuX+w3Z5L91R7FijIAAGCcpfCsohlzmzPR2qP8xOuRXqqgpyzFhWemPuxNtC
p75PiNDTIiZXn171ymBvk5keV4f1jrXFZUJohH+/9Ci7PD14m2j7tnyNc23AkBfjdrpSsa6ZX/1X
J/cmwlo7e3ATi35r+HxiOwwp5U/DeZniYjBIM/GzqxkGYSfQ2GXiD64NgHLWqK3eG69V2CKl6Rdk
GcPS9v68GEIhP3cPbgS5be9EN0IeFwDhjlDij9OQUA6lukjnveDX3dV/kLNvqBfC/LbhdL4y4eoe
MMsOScgVljwvaL0ixpV4oowLcHHWXWJBAl29mmJrg5SOcJCb4zYDflW45Kyg3AJ0MMzO2qRsWbug
BItu4300Ga5XJI1GAq0qPUUjmWCJOvyN0qNDBtaP3++kwVBlFz89jgISZZf/2u+l0OxHBGsiEjCn
/jKd2cxN7n3o72AIjx/LVUB3Os3XSX+ONmHQdqvPEStASSpMt2giKRKkqD+UVGQUerw687rXEomr
nTgL+/z1gxAif0OAjbg6U5nz98bnpjGfyzMXZwR728XkvarOxJy8hEZ5OsrRSh2FmdhhofGCUUYV
RK69TlS61kRdCpH3kIPDWM2kLkYlLQdt4BtdUE9YlauwE8PtBNy+ry4j60h0f6B/UUFbf4IxXibU
lZ1y6Z05Jt64M431jBItZcYqZYO6DgbMDRqT7KehlwADly+2aPAZrqG1l5Lbtmiomb/i+jy/ZqF9
tjTy34jZoyAaCoUYnrLN9zKhyC2tlsFbNErJ27vGtKKkrKubDrc3lFzLcZTsuUxSSyYBhHnpKowb
zbV49MXUFsmv8uAGypgSqLsa7LxL2aEXTFioAKkz9g4EdmWs1tLPyS/oy+C2bYEc6yUeijGn8inv
erNjZSiyDlyITOoEaNCQW+TBlNGrU76TSZPQQ2fmyJxJ92kdcJRL3zOjaAaNE6yLw+5Ru40m0lqw
QwaMO5aTT9vm+Dr3SLLRhm3kaBbk815teyRW9OuYNxpi2+zpAulpdlzZTbx5rt27CAlNR7MWI/zq
n1pBTEAYH8ZncnpT5iMIN6q9863aXD9JO8wvnh1ap20GNAx0YYAq+i/A7LwGsjdaXz/7rX27vQ3F
kxyFjTClNbHBqeMEjb3azkHG6RpktnwWwNVb31psRKu7cCHrUzzOnb9QuezmF/jbKqOjzH4Vmmih
1IY6qXgTIfDBxWlA3AW4HBWpMAVfO2kpPHJUdAkrgbinLIXw7ExcezMPyRZ0bpMSfZEHCSQTGThb
clPAA3hMXw1EhIAI9cklmzFMrmfF7ojF8WbXVwCNYilig4FGdrcxTHvFBIcDzw/CcxNGdlqs1Dk6
mox42qw1dHFFqoSGZp+SnpvMW0COwqmgPFxTK8n/y9UnK6ics3u4HLmzjGnIh2T5h0bBKb0oF1w3
HxX9su3CkRlnBX0Xoka6fMFrHrjDY8DwPlgOKVtGtOiFcmZzlR71I0lChrEUuyLLqTkGVRzAPUGV
0vmBo3qiBwxzv/rCl9ldfs36wzu7lSyVPNQM+J8qeZ4lm9koCiqualGtaOGXQr5utwn5MHGrUitw
/Gm1bD1hzucIvwoBmhPxVzkG21ybMgMrXQhYo8cbjOb0zhaU0PmONXkYHW3cF2iK34/nK/eGKrry
bYTT0b4PKDBMIjfSSYusjyQOuXfr2kLj0nbpzungrPiRTV6PwU/dZM5+eH6q/xyU9vnXjRZQf9jH
9L8VSub/tbrW98mHw+swA3AP6aKvydlJPAQYhmkwaXjBL0DJmfdhWuWqiR45T5KjjvRz9t29/Hqj
JWgN2bd1sDjk3GzXhjWB6LlG7C5VGJGahpygnTSxDv99wEFTzuKv8EyOTKWtnbA3wIhnDF0hJgrz
N/N8iClPOlRAWX7Bl9xm+OYzLcJuhJKuoZWz2Ho0pxPGlfsKMAFZEjiaD/OfJNoqeYcXmr6oCtZy
hRzG11BP8ZVqIH4BB1RjUgPQpdSwCeG6qvyhOn4mRJttBGE6MOVKa8Fptkdoyts1V8FHsniDB6ck
W6VwVbhTK53NY6hnRMBJm3im90EGFXPHlxEpiRT68rE9ixycu3KBJdaXSFBhsqnX2dgMzWAK1uT+
uNHJGr6eFz7zs6+i32MHWKTlPTi+m0WlJV1c1uNvq9A8Owo9pFCtO1WSc3a9GlIJ7dd+ZF7k+HBn
pIVcr84cGCMd7g7SQjxIpgwP1vhGndxoD2n3J6kNiiDzJVzZgz88XFtyxKTB7uLCvtcXAQ+z5NIP
EFhYIU/wkpVHv+o45kSpV+Bhgk1ea+hCM+tWtjJvn9lpwxzgSiOO46Qqqw/hYPSoko1zZLFmrdo1
g7W1bXvCLctedY1mXWnpOs+oC238uXHxusRiKh7ypLk9OjK7tUq0/M36bZNwICEtCwOZPcf3+aYB
F74YUjqybFFG1HeKRdlSLQ3ATD+SWwB5ClbZNuUpvXHCgHRAKL95ZC+qMyt9Aoz1BzGNszVyk5PO
AuAp/pj2eqnDuZoc1OhIc7FV0Yjf6ad618DmXbVIT5GxfelbQL61hm8mZ3DspQwroZ3dsrYlmvtx
vJ2ae6391REAFhdDGdfhmy8edFSeHO6Go2ARA6c3XzrC5W3fkt3PQsCoJAW64i22IIJepm9m1ENC
yyBFlxTaP0gAg62wxNKBaNu3/ODH0Vkt10RZZP+N2p6ykReXc5mICiuXVcDvyrLAkSfN9dVbb0WP
Q5kIg5iRGMtJMKDnjNZe9E0o56OBhTC9eG+oVc/0znwnwa+ZGNmU9/qPMGjxPvmqwXqp82C6gnfR
SPj79T09DsM92Fjmw80NiRTEucuFsefFq0Ii4mftFozktFIiLZLzXFzDCOvAufx++4kiC00NhUyG
TWGQ45t3v8or1ZP3XmfTkBVa6p9S9YrLSpqHSqk9OHLLN2CLMo7e4VsvqBCSG3TtUIWlFcELS31F
gUwyaoU4hppzFkLVI9ZbpeLLbg/UXMz8Tjo/G8rSCD8466ayojguEwX2Z6vk0KVnSl9HaLDQuFGt
cR85hv7j2t42KjWwRPq8+B8MbW3obiS4Y4qr1Onjf665LHQmqPNInTUyrtkkD3t0IwtwfoKao6/8
6Bw21NAT01CwQuOLWblH6Knl4tZ5GR9P2qw1qf/h9BV6zPDG7KVnJoJBOaWRecZ8yKrQeL7mQJFy
4HQp34DBPPOgBdm+KJjpxPLahvmYNqyB4Pf7KfXJY8CxdTNFSIUjfhOHmo8rLle/x3kdtLWK9H8o
mtmbQLpxLFmmKGNEdejyy7536I2VxLO0APXYBQdOWRlDsfROS1GcXuW2934jtmKgJrnmwYJsT4no
eJQ5etSod/WtbkenhFpvJgyfHgeYN0/O5NU5mfvJEmvNNKRXx1RkmWSAIAxzHxQZexzTWt3gROYO
Xzbi1ujEDXnw0Ayx0+fT2u3zDPQuQ2NVs8wO1zRjB5dnfeHN25F7hsI7kegDjNwncD3czrSvaTE+
Zx7cFw8+u9JbYoz/XaVgBNGNkw6sUKwY5DzgQLKccw65cl28OhPD1zUYOhxFlBwaoZxIgwikDi6r
h7h1ko6gR7b5PRSCDR6ZwwO9fczx7pmfZ55AN9g2AMRUTdduh+jSbGTuZoSyYvtJFZZqWNwCE/KC
VFNf6M818IiRf9pRFoJrQVtTV7yF+e08CZI63SZrJWcAcx3Jtn44OScDZpFMHAt84p3Aw0wfO2Is
5YecDxZpW0L0NsDMZJIq+hFjYgjG9cgA9ILNvxSY2C/jfuq/8OqjN3B+MrDEmYO8l10ASXjrbq19
oZ+5iTHhLu8x0ZM8XAp4WDLkLG8yD2r5u23kUzC2QmwtwIDc7UY2YVjgXd89t+6aAMC5fQV7JJjc
ZfoP4nf0PdkWS7fWK+T0+T6r6j+2tVJVidz10kie2fRTgTpworBPUlpK/yhqZ2NqvjKL/9f23AVr
sEg6kn5MVKCFotIHju7U1SmW26dBjcAqug7ZL3IhPbqO0hVIy/1CwT6dVPftT8MtonUp54RBrfNC
SnvHqqqGTDfNvwma6ZyIQePP0kK8GC5wSb/IHtBmO7VTbIjbEeaZ1gFIdR6XAjQcfWEcKhxC1lh8
hkcg2289+M9AM5bFLnNJfCaTKe1GVknG9u33NvCUj2JMtxDtF230FCBQMuPbRMN5Cbpigki/FBFO
DVy3y3WQE7lZ9truArk87LIPl8NBRELdm7byspXGgsK+xWwgxcq+nrjSY+1XB67VSa7Vs7eh1con
uZJlJPLm0atyORBlTdZNKn50ljN8/pJmKsjK1ibLuMP0LdPgmZjCAylM4W+yqBaswMg8BqLRXlo0
wiasrLcLR/SX75EJvi5HvSrdxz0h06gZ1JSm6QaIWKSOILqdouVpXrbYw4ep0h+BAQmAXgBPN1s/
LT7M+J/zWhRLGM/G/CoAnN/jukPKJIcbO8xItizD1COlpHH0y/6y1Gs/WNYgbwYwTMu642beZ63O
IjaGf1ohjGIFIT7/a5tzTWVw4C2oW5xxpcgW1HSh/XSZ59HH1/bmqBQcrhzUKZUAgewXKxxsIMDs
FJNwFTv5sVRYOpd1Ts0tdPNhNKUAYhrlRMZgYUgb3gCAjZsbVmpQVjOEMPJX/An2r9R44ki6QERi
Qhl1ZWzx2V3R/fA+rIgwh2khbDT0RSSmq/WoD7GKdO+MHQrcRjldJufc/mMszViRhDfUs7yKUs2v
fhdmlHZIckDw5Zi8MoyLp3zBJkQLxa5Jl0+mLmp/jgG2Nz0X3zN2LzlNFgooCxoHci9hc9RVx7g3
pAOFsltlCAno9yyPJalzFYU0VpDr6iDYVFyw12oOYMRRyQ8yGJdEXI9pRn3Jr9mEV36lYZ6ffpsT
yGiyizhWUv//oFXZK0RlRihhBH1NtT81wN73TKqCXW5zWxemjrdXPU34xQgF79W+NvBNs2ujj+kl
M/gNDSgyftAs5AvtOhVQmLxZgVP1GAwQfFPSUgS7KeAkwtqc98t7e6HVaQllErFMA9RUkUAGhg4/
yT9BM19s66dMuWhXg38slATEg4AL9jVj4+ME1mEq+OKTBxpY+SYJP7TWub6KVVoSqyLQvNnMk10C
rTLA21Hnf4mEzkchNTxuJGuG85TevHjyvNDpP2lh0kXTN+Q3skBFIX7NpTcNOqG841iLtA02hQha
IBupMjBnt2sklMRzYvSxQLOKGLgRT21kKn1I3g6ALWe93OhR/xNDwcLogxpa9VizzuS4hIGEvytL
R0T6k0/guVQDN7OOnKlaEHwVtXIfSgOWgJ1pQgr5NOJrHB9rA+COzl52VyozA3i42yhaCV630e/R
PL47M41NqTfIZzaXdzCqfnvMsdKV5o+kzLQkS7MGG4WUQ/WtS6YMOGb0LDHg1tCbEj5buTiXSQOz
t664A+W1HK8wmHT0IFEswSyNw7lb8sB5S5kMoeCVWvs2RoeYBZ7pjPj6wZC3FHe2mtj8u9uFkasD
ec1aYMI8xZypVFdibGzu6JtGEMnpZA72g/grNkCmks2nSeWWTiUT4D+z4VN9psEUDh46ohDNbJLb
JFGvNGHiT6ok+QTFLxK2ljcJdQ6yOebrr7HbB+Rl8dMnfrLOwZm2nIAo0UT7Ou1uBN49dOtVAX//
zXF4rdh/IFW+IwT1dT9aXIG9JjgTZAxjBhv25Vg+NfAyYoUdEbF4Fbb/ejg74XB/90D8CaZbcJSN
NiRhPpexreX4ggxUjabRK9XbmAR7cbTZErmyxEkgLSBw+vWkW9PBRMTJVWVM9zojEd33Yid+6UVt
IGn5foRCNM50ZHRguHNikNA5gKWTi0+yydyqBhldW7Sh225o0U0j6CvJK7qd5O+woAVjh/V6hJzw
StQ+8UA2c4c9vDSs3oMTqnr9VgREmz4kyKvy/S4YlWvQzYUo8TlemyYbZx+k5aeYwa1+TsrWceNg
Y0BP+7/Okhu6UugiFh0dv70I7M0U/1M3lDg3hnP5l01/iGevJeBQi6XJdsD/YYab50Kmv42sM/GI
p0XKQbhEtjj0/VLRWQCbX79A2eNYSnUqmO0yAFYn/XMQEyRUxp7QUVakVTbcCZaOp189UCtZ2l1r
FE/yVmjc/Ds0VcsCXcklEpLvohMB18i76bTUrxHvThsfE3GRZv1CyRg0hDCrWLbNYiwALiiMFahB
qLeTu9ZLcv3SvAsyQm/8r2UhSJ+es1q0GWS1u2bnkFSq/V+7UAV2eU8hjmxoHguvhdf7PX1ffPR8
JuomWoinADGy0ayoT1T7+kOZBoIva83mTUFFnROo6CXOoCIaKeFN5v2HMyVSYgLGzmevH3JJ5wwS
GVXGszavbGkXHdP+7NWFZPtIHSQt0QFffyL8wsYXk1eFSnv52etTjtzdz6vPHloApN6qVpmirFAw
t/52G0LcZ2jkA8yZhAzzGcPBX09f08WCkGjPoKof+6XkxszKxpsl2cfSDQnzRTFMkZx7Ts+EUTOt
hFLjbwxd3rA7R6OPWQyDf1RdukbRYjbZrr7kOzZa5A/ohr1mGIjhNKYedvLBpeYsVmLC8FjLxdly
BcNmpIaf8bogfAhIIEzZORbqwaK26e2+QDI0Aa4vsy4p3YSZkNq/nwEZA8s49LNnhrB5j2/06JS/
fTs8BkrdyPQ+MPt+g+YOYbbRNpMyr2c1a6Y7h4ld4Q9BLuiE8Ms3fJ6Wbpw1yU0WXJ6eM9q1S20A
WSQ1qNITLlL8rw+v0nuX7jTLY2+nxKYiyyGB050+wvDBNb4Lje9uZmv+3maAS88Y7cttarIomCsr
+xamtzeE23EjtYIMLHVSbbADi9GkpTxHVya/h9SpSTwyhQQ1CJbM8UlcE05vdXIz53ZUom3aKcbu
0gPoWY4TNEhIPGgb+q8+1hslDYho63Cx855WIm4lbe1ONxd0XtNZH9yGFNGuqYvu9hVbYmbINA54
4V2XdohztdvEKd43TnpCSaYyiNB6vDCXaz+k9nDiJn35F1RJ+aP8D2QOm9rRKCJrM0+c2eC9YVMT
52hKjpwn3w22NbKz2fpeLLq03fmzy1N/T8IyZ4lx2OgYU/a48tS0au3+2mByv26ewJgZsDlZ9jq2
cPEOmPr5OLYyyw7D5BPcCnCKykHh2Wq6xhEatsrHinet1xrsj69ITa0AvIBQ1YaLDszzPXCba6yN
PTbMsTIy34Wc+geJIfNdL6WoqdftK1Rc7Rusuh9xbFVg0a5fqJiH1KiuAEsOaxr5UskjYm8zs9W3
b+o11NGvQhLuDX4iTYzYLMxgl+XWfXH7j2AXCbaE93WVgwKaN1frCFQciLauXdoVzf46ivSsSIl+
VR7c+Yj3nCmKEbLQ
`protect end_protected
