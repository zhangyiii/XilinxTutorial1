`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31872)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMK/PgSU3QY91fBkoay9fSdIXCM
AO2YSxjwjCCa4kjZ6EGpHLsWaRutaBcN9VFBZUxk88GZUKXyxFnz/FEntp9Y4JdD1OfzH626OAHc
i1zmQa3eDNw15stEMGYeYb2JzeHGuJitsFtt3F4PaUb8tqxTAVH7Cq0vCshswcZHqxNzvxEiO2qc
82TmDBZ+jGB7lpzN/MA1Y1cBIAVSTQQ78k/vwFobS36Sl0SJ+9LLlVbL7vOgplkHRfbygk5Uq01S
ikffXlJlbZJml3na2Ji+XmYB8lPyqeQFUUvcVDDpqGM91YSESZt1OV+l7c+UTeK9hTbu7nrhBIyi
w9+1BopnR7Qdl2vksCH4GnxhNdDpjTxc4KQpxjdMr+pvqSarqHc5vkXX98qJKTmPg9MK1y/tGjmE
gbKUxPCRbbZ+UzUHdqETyqT/oxVtuEyo080upJkuLoaZ0mVyG6lxOBcDe3a+MF3g6XAb6GZhZ0yN
gJ1ljnPr3adn6R9Q5dwW2GXG68B5RaQd4DBd9ud19e7tLRsaoplU9YtDRU+xShdodwa7HXLSS/w0
R9anhChZhmJtT2FLAc//7HSq7DI/C2cp0x23/QFeziaYD8bRiSO+m5Nwjn1VjMHGK4G8QHqAFSvK
wiF/tURipRxg1kPTbTeWxQXIbmW5iZJq9ug3NdNP4qtswJQbe/x6sl2CWZSDsMpmBYZJd54KBWxZ
Bl1iyKuiT1vBiN5ZXQvABZQiVUYye/dnKjluwAgt9FSYATex0L6AWD0v3RPa0j6t+Gn94pzuFw2W
H+szpPu5UtB3tD2NtcJmYLFYdteIZF4rZP26VsvX5Q9L5rNDSzl5kdmkppEsrf2qSiJg0YLxMBdW
6V1fhuOdJ0j+GRjGI7cJ7iCTwGy9InsQDc3RuIhCGg6PUIb+aJAUILERbwxrhJcBelgoaWkuiGC6
rfNMwezuKA+Ii+uEXsHyavypPGp48K/kCTuP9SY8cEWb4XIjbew0g6yYcy9rjvzJnS/q6FydVBhJ
YpQP4XkkZsP6xG0+AKoh9q3DXK3UlL4XW49eIB/pnAL5jO8jnO08Le2FbSNupd7DgqWUK7o2/3CR
GnUaya9rPkZIv+J2yDKC6Rresk940Aje1pWQo9pcFK5xPi0ebnC1oRA43gLq6oRkc5wgVArxtR6j
cTYhE6i+2E5xat6gVVl/BgbJwHNC6KJ01u/pJyCt6hhKxfADu3ELlXVUwZZmuYRTBUoIuIwXYkhi
NArJtrvVvTVGP3XECVnyQe++5bXOKrziBj7kuOd5MOjJNWBW9zxiRpXwSYFoz6v7g3KkT0synb5s
uWlQbd8D+0PRPZ4LdRE9hqyAYKxnXi1SIDhbt5J1ERsDZUeTLhrLnP07Wbbhl0hk0OziElZRUMHP
2m8ZY/9MDzkFO5s71G8PR/o6TvL/8TFJAdRlmg+QnS3EyVx+MbtM3T651k5hvmToQOdCUClHJ6K7
QMO8tyCEIWclHK2OP1UASbulMWVnIh7P5posVMTJwaboLdU8aeu2CmraYlBap90B+FOeFt5jr4lJ
ANCHFGYJB5AZOGd08vqHadGnSxFSzWT/mSqie2TzeIt2ZM6Xw58rYDsY4WBgnipIh4Bgu6SRlK7k
/p+XL5/m+0s1IuC6pizkURkwaO63EFz6YzhO7HSD/Hg0JpXLksQ9MKZ4SteDIQg2X1XT+WPbIyMc
erqJiA0/a9+WLwbg/OQvVyATx2oCKm+3tqiz9+50nEFqrHRYWFCdbIP8wdRmUavYyDaR7zkSD/QZ
fAGEn+kvLFlyQ1Fcw5g6yyaQTksjsn3Reg8nYROyPrdmT8cYEIV6s/iMRLI3aNYaSlV26g9ZXtXn
Ioo7TeO/w5Mf4Ld/Yq9Gc/dzOJV9IejcGxhuyMzvIkLV3ke8dTP40ovOgV1u6XS6v+BiE3y6M+A7
QS2mQywqrpbQZAI9KNl4BSdM7z1RBuElJaK7FQfs0Tllayfuiq0hLLSmIS4vtShkL75Y9gasNCo5
kFczN6yOrwAr2i5g0x3Z7xxwYuUTck4x1ZNZ2lng1AocAtdekDWOocltZWhkjVSxGu5eBEDAfLEc
Zbw4NS8sMDNih/MfJYc7F5/j7rnYBJSCkFNeji9QMXLwEaD3HA9WIyWznJE3LA2364GgnR6r8itS
815YXS3kNoVg0v8Xx81fmX2znOmJTZrwFLO47pa+JcVgAmukdPqPuumVPuwcjYY35EfqXvUPvw2u
Mdgh9tUiIqy+UMQZMYxNL+dISh4XE8ESALDc/dpvbLw0mxccMOCM3roBwnuc0y8G8jkMlI95Sf0I
Mln/h4usCeJxzq9QrLjrkCB2Z+ty3qzveGHqr936E/IXlciJcdTOOzMqKKshE0Ku6xLs7oTpC+HV
mYspOYpxdmzvGiyXX4/uVpXP7mU//DncB27Ryjur6HBHOKBlEGNP1k8Zl3tMlhtrBevdFC5qk9Fa
qN7XdbzE6NtSv1AQVif3EtBX+aCwTYO+IvvcIVFuDa9tc8KDrEp/ldLVQGUwdh1rSH4ilJI6mfGd
xWEhIw8kApUXAQ7eYaSK6/v0hW1zh9CXrrpGfDdc1PubkzvC119aNec5YysWIdmGQcroliNOtk30
g901IbPUC+GFhOopM6A4vs78KoRaUyiiITOXr2IMBReivG/EEUREeZ6F9tnS1jkMffhB37j4/X7W
cpV1llYIdtx9pPoR4yX3wwvxNSTHW4I6GxWKEeYpsOOwz9ZYzqMBmrlcgP1cm8ALPioHJBha7HvT
C7BaalzOiRc7UQGJWKhVVr/DCYz3JtubuHw87RHyNTbZeaDx5cw1ekDmlIwDk/Fxvu9I863MNkt/
HyxVfiALz0IGw8RBGe4m68pi/6c6LVgItVC95Xd9RkdXlCE9PcfaHzp7Bift+aLWCeN60rEB4EHG
/h/wSR3MaEy3+Lff7lelhEOg3v5YFAoPwQTlY25s06L4n6yFsB5TRp5chIAMxg/mJXiQVwfig0Ws
FRmvOk6pXRcK39kSLVwT3edkDk7A4aJdYHj0gtb/jG8u37wmZ/crnOQKFS1IS5UFrSKtpIpfBykh
bJ9rW2gdhNdFQi9fQtmF+QNS9JhTfmYHF7qGi4bJ3gC+edQqHNIxTzuqGpZDOpcdAeXWTwRXVGYa
vFKVBUC/+xq/awfbnm3K1GjSKzfyk6qD1ztSbHds9KM9ln7eosZYTJrYdiCOtNCP8t2HMlx3Z56K
imsppZDcRW87Yw1zOficlqCSe+oJdqHP3uZGw0YNJYjWaCgfh3YoF+h1F2lBN3WqvV5w4ucU6G3R
31duiVvJ9VKfN8QaKrNgZZWWXa026P0H0HWin+7pFRfQ5u/lcrH1LD7ftX66f+mRtD9C5QowXAs3
qmY9pNlb1x7DrG5KVK3OyxRML2OqefHUJsCTI/LE02bVR2hjuAt6+JBRera35uIjKgr+ipM3yosZ
kNuidSCnlUkadDBiqBLctO9qWgGFvYFAmWVIdYb8c7322HnHOc84SnR8SFaw+7PtaKUUHaH+1j9R
jyCYuY5cyrTPzP+iAenOyylqrNC/Hd7dq7+nW9Hof9HQlpuyXTz13WGD8BVf3xuEtY29qjnflPK4
H8xzEUtlvuU8BI6PrgNi1Mz9lWtkHDhOl5XVir1j34EZez6DfeTNE5YQ/YPtUIEF4c/eFU2MAOPb
7zoE5KJ7Vqfzf6EIUnaIPPQdPrBp/hdCxxUhgQ+r7wBc30Z/tCjJgPPQN81/v5JJBa6OmaqlzlvN
b1SHoLmFqc2e1BHPvWJbzPjJLthhfSt1lJv/1qlDwrm1R1rBgAS3gvL5XCvnxDm2yL2xoTl6TS4n
HKC/XUS10SZHhiHd8814gh21+VEgt9zSSz5CisNi5+9u0YLo+/+MODULaWYH1wrdACMvG1naZKi+
SLwmD+lfMsQ74d+jyJ6mQK/t2saedF+C54zJ33d+X6zBfpgbfE8yWM5T/jAG2V/mUrZN7TU+JRja
PCK+DGSLF0qEvQWwdlEMiBga/JiPdAWatkIbjivgDgtq8Ep7fTVZxSc92ewU+/Vw5zI9mSD+0a9u
A8iBVvhwRIOVu2dESOlmE6ebWaQkIm1WF4RpBmICoGhn4Kjj67Q7ETwiOeyKirppE4zbWBIWtz/a
uAwIY1Hvf6R8GXZPV0++PN+ScG17yWyClJbHJGQXwsXqEgmLRswJzDecDtFFOQNre6xTriVAkGpj
MlbpI9U0DqSOAD3U4XyuhSG9ZhMxmA2p641Xdbj4q4c4fHZJG8dGlw07Q/1q9Eq/i6Qa89yLmqbu
8H1bUfH8McX3X+SD0lSCnkTVdQrN7em9x0mJc4aX8r6iGGcLreUYCfj0s2MsAfq89d4EJ6Ff8+SF
gllseXhcwNKjtmgHExVogse6omcclkfo2TE4IAGYftaGtLYq+YNLBToDnsfG1BNA3cpWn+lrj/9l
5gNmd20JLXeV+jlG+aRMdIggkEsK9ObQITWJQMpNGRDsoJCVIe1AASqaLK0suI42SkrvbLruB1X6
PmrCq6gEigGx89PfWkWoqaGQa+XFUFwJDUnLptH3uptc3o0PCDuGCToSGhUl6ECYvtfRqo5SYsau
IoE7CfpHTCIyZsJ5I9tiDKbQOgjddzjB+Sgpdwi5slCAvW8DUItvvR9f2OQwejMo2Jpi8f7oR/hZ
XgKhcz7js5WX201yQ5hWNUbR/nFsJUd5wX0uQujXa5PVqfmS0z36LwJ6Jn1SIogu0dqsuvJdVvC4
gUgrpYDEVtC2zPp4BMmGah/c9s3ZShWHJXfLlvbSjjqeU91r4kMew5BM8RH0eciOE8Lxdo7BQsJQ
MEB0XIMyPaCn/BOpTRauBphIWUBn/cLX1/jLaR4zOUuM+bodOGBv0ARNp4YYxh1xMwkputSECYTD
INZTn36XzSwU1goSbInIXTYgVEhgG+tHMq/HEm+skGSyGwmvpefnomro2cnF7Yu6tjVJOkC0S7C4
0HKnkNXXnHzIlU21cLtUctuDxY/PEGjISNWuRbTCfkZ+Ljdzqajyd8xKCXLtb8fOHHZxK5/VGZXh
ehtcqMVNx7ttPDXjUsh2u/plWp1PlCgJETEfV2tANFOhWvOcyS2CzOQE3dov2oLKAZhZoIQYWZZl
NyZmQ2+FBqyXKgt5oyqzN+2mv9q57wIzrWKA1ur1Xl6gqJlxLvtEJhrgd+t/S7UL8R4H08z8R0uP
b4GB442nGjvDET9okW/v2XZqMApv/6UBSsWe29ZaJutZhMZZ3yc7GqiKkmlPu76d6dy+K4sp31rJ
3dpI6lSfD1/pLVD9qAkOd16S9+L52ReBKR6N1ItOp4ij0iWrAjLUyuolokl/QdxDRqEX1UHSN9p6
K0UtdnSdhgYCpZVeOAHVgJ/4gpflSpA5YMj65AmWXshRNOJojv3Hpk6Efm2AchRiU9mHxzxmT1ES
oxkGO0YuDTW/Nz2F0dFwO3DC3OhcAv3CKYiXrpSoeOCuN8EkEm5aS1YUVOrKlnN87KabaYSK5j6z
7i34FBRNyLIwerKeRtM6rM7KtSGN7DEo6uA9TkvUTsHe14Pj5vbi85vbXXAURJLSneAEDVV9SPxC
OR04A9pU/dUCOmezvqb6x7KZ3JR5WhCGRmNAJKMAMRqToP0aOKgDe0J6vB5FRZPluaqfbH3PFzzI
HDO9urBm6wEwWiQ7lu+jAwNMhgSQGIPcc4vu7tqiq02ZEfC5UskkgvGSHFjQYMjc18xwY85GCn1i
iT+T0FkT6w5xdIVV3Gtn8mO9pP2Jps7rlDpE5z/GtjSwccYHBkghFx33mboHfCOJhEqrlYPd6hih
TzAQGCRCy19+h+/K3TyuNmZ2THVXFFxH7bgX/WJ2gjIpx58mJqPeFHlVD0puxxM7TDuG+ZkltPJj
BuAdUFqWOzRK7Wm8t6xaqgFKsqTxjR36MGXSkeJ6AqCeLaJPdLAQSbq2Wcjqok8reqUGnX2hlTan
/hBXsWjmdgP5Es7wFEq2WjNU5pj2aBix+aSDyBwU8ieq+ynKVpa9fW3KTzMrFcV2LLCA4L2MrRQy
lbGCZ4LrZxSTRVuNi2FwPGhsvOaQLVuY+pp7ly/kCnT6iG4zMXC2ZLdZpBG5Vyt5JrZ9z6MQfF2W
XWqGGYsY+NdPeD5f3sIoZIsL0y6Dy/wYbHJ8KNtp/PGNdhJbI7IC9HUyINEL6r2KsVOUe8Muh26f
MpWo/ZtUk21RkY+heEdXM8dAFfBDFUy18dJZe9kM2CoPk2RLNnuOrhLvjR8o6nZY+7UgFaBwgq8g
M+1lLNZRXDHac4fe6OhX9/Ap8WIzG+kbtxmRjTC7iTb/PgkUYOqG6tWJYJqtccS7Nmkl4MI1821+
YUPgXbG48jfMMo05ckTMcSVdYa4MYEMr+QKYah+0P43xzqyZJyQHUlwP/laFLyNgBwm8QWXzqIF2
HpGjDmwElaLLjiLRRDrR6QtiIhcZkGeJQgvQTUJFywA8lz795DtFQ+WlUCLojTVbYsIIAb6OL1xr
JS9jH13EWvHkqCHnDTiAedfAIBQ9/8wa2DpIzityPNnxIGRcV0lph3MeSDz9V25X4WY5ouAhKAJ1
ifZ36xBbv8ZzzrJDO2Db7IQRtdrMc5jNljEG7pGyNX7bdTqfpKYrXIVX3T6NJT8mDxMh/UsXJM1h
r6UB0MwTi24tDE58KyzqycVqT/UB8JhER6wgbkMkrHMk1gI4dKOBUi0tUixv1JxRmliolh3lTZf9
NCkiomC9BxSJ5B6/mnf5EtmbJc8VLJaa55Xe0Xis1IADFUGkYjUX1C8tjMwqCWT209Xncw8GjPhN
t3xfs2pye2GcPm7KaJBelqZnPlz+NBR8h9aKdkikld1QZXuvsI8u5wDBPOjfcislx2KiS+ypyE1Y
x7knGLxKhwfn4i/CVK0Jg5L0HM1dxawiJ2mt4QYf7K0K+HG5qVaHestGo/owLsW15APxnFDFkT34
6gSyyVVZp89Kq0Lkxmz+PEtpjb5Nrd/P31pmzf1E0kYSedS2XqF8zUQU3lASTtNFWLXuuKMrt9Ff
coWJExp8kJlNG8Di+0j+uV2LXlXMUn4sOKgJitAGy22Ix+4z0fU4s/7bD9hLlzXVBTrcuNgKcfc/
yY4DPx/i6oiRHhO07ZsjyF1j49xhMjjpcNFTPNypsoCRujYbsS83q9TewlMZpC/0TQNw7hmnXfCw
h0tI5i8m8WtJTn3Qzx3ARfz0Kl7qbOJghDxjWZK1NlYdnZJeXmrL/AdyIE7oyzN7kUZ9fJReo1os
VriitXlT4jUKowVJFNQdYZeGbJh0AYNvYRYCK9nxU0dOtsJ0L1MSLQ7B9Kn0N6oUf+6hh/ST519l
QrWBOXQW5vmBV2bEcpwnZpE5AUcUXBCEVcDDzMWhZJ+zNPyaH8G2qlapTuOKO7Ja5fbZYASW87k5
i/Gjh7JGxv5zr3GEv8CPbUfTa+c6bL0VyGPKGPy86L/pRWWfcgE/xtHwWyNUQ2+UGuxSy0wM9lpi
y13g5lNnqNEH/CJXKNMyJEbpqqNaVro2fK1vRs1mngtLb88s7iyBFA/dg69Cp3Q5bahwl1QRmiSe
YkRoxRsh5L0Pk0EpD7bOtJt1fgkmNPxKYVretYDlGBGukU1+pTon+AdjBVRiINhV71SbX/8w9uMf
h2oa1/k0Er/d+mPATI2L1dP2b8yrVQw9P52noG00Uz6kddyptj9ewnEJ+ciYzE01ljzt9pPOvi1h
3EB3O1AnxUqMYP+iP5zKtyZyp+RQ7APURFEt4tIOriMQJgE0kRuzoU6RSsM32KnLjVV036tL5msx
gWfdH6NU81bUVAxzakLvIkalyt1vqVX3gOwOmr4BTuxZZVnS9BAv8M8UjVQPB0n3Q4IJKEXX1LPl
RP1HZPsxC/WvQlIM5vqs5Cp9ntn3iPYPptN2Dt/EG1YyBqLHMoXxBYEI4ynlgLgTkjFNDuS/TxNv
TjFQXyuj/SNkgleOTC+8vBRTwjQUp8pCSHJbImIe0bPY2gnlrPowGNTciI6/42pt/O4hlREWo0DT
IBKNQ+H4STczVLWZEprnuOk4Dc+V+lV+rEq6uhfhMwwMAA+x5Q/buafY0J7Hk4hTVnQjG1forkns
YS82twXDtmdSStlW8gVE7GmLVZDWo/cNOdiRMnLKvNWcS2pi93xPECuHrxGm6L1QXOKl9zs10SeM
SZmptjyM/xbAITOBOa/7CmufI+i/cOkNSeCx93VtnnGAncBgDQwPcSzYXrwzIaICZtbI295ImeVe
fYTLIm7Ey+gnv7bascnsiCq7HHm8blPEMpQumHYLIc7fhqQS44cAfmh0ZakS65R9qFjGrIRtdOjP
vBQcvCpMZyJb/KMdDnIHkcBD/TgVPMX6+Ny1X+9I+tHDOI6lo5saCixkNALQ3yuZ8hGZwckuxEEN
fueGMmKBs/qCfOZEKaGAyrUS5i3F41wwA9wcm8THnNN/N5djmGR5db/M7ClqKbkiMBXsLjGw12K6
BTgdV2oRUPG3FCNtqX7cQ8e1TecoUP66+va4Or5SEVUvaY45PlA8YqfWCbrRD1zx7C4ut54YY3Pm
7PBj/z7QqYOGht+EBaroWxLk6yT8aa4Ke4egnQ3G+chXzNSBIWGdOO+BRHIBAp2RvC9SFj7tKNJS
qv7tAvPk3ZGUHAtJzvkUqBi2zwNQ3T/SlqMGaZgv/ztt3maoPfvXbSHXWfovsmqweQ4CvgJJMOO1
qGs0aqtaazQbj1nyDxyLSsIGiXgUkw8Cktu0dEK77A55410V6P7GW2lJ0FN1WoLPHzo8oBxEPog6
/+XwGOWi4vbNARh7RO9HmR/x53vghPh0RN+qCJ2WQ8d3nl39ThYBfvhL4clC8kHUDAYpLIbusC0Z
HonZEDckedhxXpEUAxjZKnQCPahgUEICqIrVv+WGy+tDnSy4+j/o42gYVZlpE719yvPcjTCefDp3
bsAqXB/zHXAMOF0rw99jKk2pKqtOoFAMPvFXJAYNNRZePsgs5BF43EeJZ7TECbWPJO4/85w+zCYZ
ooX81BiCWv8OebK5UtprCyUQDxvJBrEe2qlX7TCOc6SADfOkJoz9YHaGTiqGe22PW9SYZ0hzpchR
KYJz8s6azYvSovCoPY3gJ4iKUZeXCs8Z4TC6ZZkwtiiNvNnpN5iPSWMNgpjyOnviYT35qKuIRUj9
6ZPwK9h3Rzu9C3TT/j1TO2/uPU0JQZQhlhDF9FsHEWTlnLCRgWuTDZwfM0rdVL6SHg/yUE9VvG63
9xL7j75jhkGfyUQUQ38K+HNhwIW5LCFerIg4plqesmXlRZIv5WQCr5U/nmIqjs6qnbKz5uzrpCu8
j1kWQ1mI3qQkWhXF4DKXVTee58rL2AJUEZ/h+fM7+DtRdWhFI54IfRGMaKvLKMtA2AdiKkFSoH5r
Lf75UXrfY+jD5ztUrt31lgR/+8c8B3GhMSfDfpHI9uSzOENhyNUCzx+Udm4ps4CL5W1Ce2kGNvF5
gWUpLO8X1lrwIFYnuhRAFhECmKMFxalECCgsqSzN+TQuyqNjh6oWZeKStFS+fhuJIhtAQHoz0zm6
TaoBVk1t1MBZ8tTZvtporXP3zWZmo8S1+alduouzR1yoaD+8rGnXBa9Zei5YffeV3r1SCgc5K6PD
AYkjH86d3KnoNeOI4WTbNGF/mCUabLtQzub/epka9AdUifnluvMqmcv+YziSpKDUfhTk4pDOjHls
svrkxCt7gmaLJzk1cF39LjiEvlKsv1DnvQSB7mZDgyzutC1W6V6Ad50tx8lmgaOxOLxcihuSkKMR
3WqdHS79YTfbdX1WD9zN9f/DDGMdQMD5fngFyHZcHfjjOPYVE5DhpF3JrOIxkRpoVyMmHAUoZPl9
ek/dj7S3pO+/b+Hu6OeSyt8XUQ4Jnnx9ImMYtI5dLbAsUcikVMJw1JoStGRkbj5KIjNXIon2ZEZ5
R8+2j0WMSXoTVyTKeX4c4lPpJryKxx5r3Ogn1IcCt8ItQbOUYdq4tWQbxGnTvrM8nhDnhMR+b15Q
VNjj85aX3kNGDi4TYmoz0Mwd+z++a6Py++rGsmYnXj6pqwvaCoBT2I7CR2JAG6gW1FvNcTwyY7sx
VBbgdzCSts9Dt141Y1mK//amGM6tfCuqB5DsaREhA2W/pqHlAfaUZ84oD5KOhFGwjkeFoh6BYgDT
9+h30kfRwi8LxOmooYUbBNfNM0i47ueGiv/GpxfnoT+OKN2qJKyZzSoJSbUtgHLqcAT1BrmL5wlu
vEcEbv9pWpRHCQPel0WOJkQs/Vo0gn7IRKKZ00WiFaFzrMlspKAbmBk2zBGelkNerQoC0zKzABzn
QzcwvMZAsbztXY2hq/c8/adm3tLO+Dv8uRFIzN2HwysM5hbrxIU8Tbnqr4nmlGrfwu3yP/TKyZLX
kUoKWeyCQDXn1IBT4rjhz2g2QR1OPoFsVy2NG/3pmMiJ43Kr2c/iJFA3ieMPZY0pUfGG7NpwK+nt
2mO/dg7k5Htkm4OdMMyG9+l0g/zUh2E9q9LXaERX2hmHKUrUGVP5c7UzN7yNFScbYqzGAmqqFwlo
jXX7lgOzH6TnIVfUrzNLShmXRjqpNsD8pKRYNfQChRYVek172Kqyrismp29acEcY3hD1r5A50BhH
Uw1/vyP+RO2umMfCVn9n/TwBJrDjw0ejKRzB1MScLPof1NAtW2bVRZxP9pRrxrdiH0s7VDsmT9C+
fa8V/nF45nC6aypGq1IKWeORv98iurCAQY2u2mrcQVG8xZ/WZA1qrYesEZ8R9p+td6kW6T+wch4n
fPaDbK69Atcja7jIKaLEBMqJP7W1/7PaynSWozq0STfS+SZhJlw6ZML0vxeY2gP47bYP5ki6c9tc
MHF9YrDGu0K72mcsw/RZZ1F8hQCLywRzFQs3ARK5Ll9XyOXXGWZm1iBoqw1JZFESWBbf9yTVu2Hi
bIGLqvcQIwgW6yFH9G33uRbKKOomTD8wtVVUC0hZyD3J3fp08T63wq/S2strgVpQnIsPd/ukI0oE
fBNXGSLGoGvAi5/IUnuy7s0B2XMisa49C6p4Uv67atDxE8aS2iuKlMTv05xXbMOFJn3Jb4ZLGVkk
zecn/9x5KzEBJmN0WnWUt6y1ENqOIJmI5g/cBuGQ9C5suowvRCwnocMIzY8HxrdcS/U9fzCJqfL+
JI2xWPHBBKZApj7IioN7H9UEMWnGN6FVLkrzpp5o+FnWquFt0uG642N/U7woOYVkOXViavQyc0kD
w9hvZPzi13kwWGYJ6uxmhdYIMLF3j2aa6lbvs7nhGF+n6uSJl7fQFMtgcDm+SJJ+m1uX8ScWViN8
qBPshX5DOnRCGgyyf/DFgwu6uk4ygCd7zWv7PMwRrXGkrymqGJypleiq8rEdouIxvZzv0X3PmODr
6dfQHGWjELm9qsT7va8dhJkIxmMzaHAy3loaLom+7WTg+utOcgB/v4qaN7FZ1Dt+wK5B0+ygwUCs
0622L8dSCbK0jEqd+iGENeFm40ofXrCOb4gFsSxnWS843QGyh86FDbOwrmOOdRI0wq0S4Nt/Jm1P
zIa3ztq6EJTtxykaoMIKpd3uhDepARFSHp9JWJOsDFnvESGeo6rUv7qL6qcxgzkfmgcTKIbTFIne
KkW097vQTiTUUa7162I95lcFl66nRY8+T+t+DWeImxzwZlqwiLXvYvCujQWIj4Mv8tbwTT9UY2/h
7TnVvwU+D7osfAJ3J3Q25UqWj3mL2pH8QKAyF9ddlk6ycOSs1JEQ+Jc/eRznIqY+UqRl1RJdnYso
p1443S/o9RYrt4u61r8N99Km67ppfdsCXvT7OP/QbCYuNDtB9R3WvfA+oELxj3ILZNn2/f3vNpY1
CtBRPi4+iOnAjzLiic+LIsAIKoooEO0Qtg/D5XI8/rFihQR0Ji3F6TT68OdnumwODLOkZBlk3csL
5lcVBYYtH0ibgNeZ+z8uTcMh4ljBYi6NVnjzigshFZnqSNRAnsAkPTzTRIEwPg4p5Oy9I6M9jEZE
zzvo7Fbp29pfVJNMzr8DWX2YJSWG+h3A5/ujkuCzrnyytMNldRTYLWbh/NCzq9y4UhNMkqZEGzj9
tvdttnk9Dc0xYcbtl9uXqbrhtCYW56hc/w9G9AgKjzJuwv+PvI0KXpViBY0mD2gA0d1cgswtSdHO
/SbS73MP5Uftqn20wWU7HQN+FNwcZCRPmK9bULn457SXsjNex4ddyKLZqhvSLLCTxYKSgPPXUXiH
Q3p2QHaBfpgov9eDQhG/kqrrmGvBY83dS4ezdshZGTtWHM6/ReC8IOvfWCOJdTlkDz7hvZ0/7Z4v
YaljSxG06hrFSpCwpPT9bK1R63Twab/ZCPxi8VFjSree2HRjrIOOSGsNJcJY4talsfgE2yMNrFPX
EmGNvDY9pkfPiAPOdaCPO5qB+QVMvwxN8P+5fV/PcFnqIeN00Q6UuQ/xJHNm52eYG11ZtF5sdNtF
iNEhFoieNqkt3NqhvJ50L1v6JiUc4OZsSy+xNwdLkPPOsyDX24G5phkZs0Ez2NT+eyQ7N+v0y+uM
oZjpRUEUiZcfuxJA8pqbdK6WsULXtiXg5E2r9eW27g7amHJukHjrmgR3FbjSSf1NXq1a5wf+Ol05
6lmRTj/rm1sc2MOaZGMrelBsKmCV4f2VbUIWp3teauZwQwfPnb59vkorC+0Zj9EVDzgMSnZ8Mkm+
fquuBKfvT0xQG4SniveUhm7xJ7hPLSCyN0hJYgE5KWW+0/unA0thDeb8ntmxdjY5vkRnG2hPcsol
kycIfvF1zfH6zB87nD/KO/BrdrXXxZUQjJrH+DH7Isywsx2nYn6DZzKacCZIzy7JeEw841R97m0z
EjOS36kP2qPEsGXpqGOan71QKBeTiUo2ZUcTaNKQpPAswe/7+PsX76uWUc6aOmxapqSFuADeJVP9
9ycb7c6GGq1GDL+JK6vz4CKYXIeuJDNgn4w4LaX4UGBsqNrjTEynAn05hvmFW9aMeqXcvIxVD58s
/6LQ+lJoTmDo1qesx/NcDVCOtfIrAjTKr22DUB8Kjccbnv82f6OFPwoQyiSacCobDS17cREueSLh
C/rj2L4Ano9Qf2PIy7kAZlMbLvIARIz3jXqCTroNe1Dkzn5KQwkAVT3RZ+eqgZeX7DFqe4kXJEQ9
XzdoMwJacAcDbuu3b1gSD4ekymHBBDCFHZ1Bx2W+bafiXnTy0QV1qOhI5EASJWmKygQrA6NeZfae
eD49dKQkHLGUO9dawCFm1yMcNT2thLDJc1q14zLZWJuGgT7qYFU4CATJiC373AV0OU1vfoTqaFCN
s5Z8vYeGNvE9vS1B+d9EkXEQH3emP9Vzl4GJY8Nj3vBkXfhmfxU+7MBILTJSIFWL/+qKXn+qhyNX
eqEFEWZCVr5prdQ59UQv+g/YQejZ97DskQ9U0VebZgQkFEu6D7nmMh22z2NtKF3pubdYca4j0cAW
P58TlEGQSEemvep9nHf+L9RKUEXjxN7SFHjc2n51PgEGhFE+EqapD5mtaz9pM6VWXe7ifQZ66G21
Bm8A+vX6DpKVcttRSWjPLBQ7TyVdDNu3d0KA30rnvPAVrguLBauy7GkRKBOAwKk+Z234OhgFPVFL
cZ5rLRaWYxnFpyj93ctjaWf6aNlUsRCtN3O97LkgfMXmlc40Zyeardq6UWO7QtmHuldpCqZWxuto
KKZ/srh0JhBeavUGFXjiWiXZQ+K+r+N1mhdVhpWKjtdfoqr5eIvYLjZTISU7sxqo28aec5z8Qf7i
ZNQAxn+NgpdF2bqwLLnNnvlleTqhG25LxkzEtQjGXxZnmvut1DexpyZb1919HfqFDqHfE7hFRq+k
mdW7pU9vL5yYvyAnTRdXOnm2JEyIDzej2fj4UMhj05kcXpdgdj0wxL1QvrIDA2jTvJhAxFf9Y4cS
T6Ykccwy6gkMxMg6mBTzuvFm2+yZQfHCV0POwpmlbdnVHrlkP3YzzvYKMb1dKQlpiEI/bdA8aZrf
05jvnIzMZDHHSCg1OTIOrI1Y/cI9T2ohWZvTqSHaG4w7Q/3uIy2fPUFrn6yl6bmNM99/0xGjbxFG
YNg+Y2CRl00m/rtVDhuoIL1RFR6CvaBZgFAVgTMttB65dSytdAAZYIcFqck0Wsln8yOgscHthYsB
pgvMZ9Dn4lWWArUpFZeBc8zgv5IsC+g7oiJpPoCdM5GdmTSRw8Ik6/h/eVdBZFmZWkjtaJOkNIho
9k2i+oJndQ3pWvX8CsHIpGmsTwxMtO8g/vFcUnGq6d2PEDBFQ/47iZQBCKIrZnK/kZTe0t3S9e49
xsaN6Ibptk0dF3M2C0HDNqOnW1YvFK106pxOWqMebHncd1AN4Jdm7qTuC4NgP6oUdQ6l92e1df/N
jAQcJ1RgWMy6jEtPwxpY4oezsbDpl8iLmFyT4/M3MUq+bykRELWgg+9hcbIcGJ91oB90fQImCtSE
mkENjEPXP5VPIInj/n9Bn1/YWR4sb+psRDN6JROafd3TGV2JWndj35IZbIDAfbhESDRkj220L3CZ
7KquxKMjXKg4Ly2sdC3D2Gs4Bg4iBBoPuqpr+itoiM2nbYwmfXvRcl3vTFeD7COUSUSjYuLaEZmE
exN0+NOanecfOyY+QyyFE/6fho9tGt048ApcBTrvtiboL8beFKIIcQL698Zp6weF93tYpY0QQp9c
NxXMnE2q88yalwjQEKBunE8/it8naykVItw0GSc4tPTtX7gur+n+TiwvGVbUY3slbh6b7m6LsuzJ
wt3vrEK5JpCoVbkNRk6sKhGqZN3gVAh0SKQ28ZrdiSG2j/vGPvGmRboy/enbxdmiXcBIrSQFQFnX
gMMVtghV5fz7989TguIYK+mVGawmR2if4hXUrlUq5Swg1kXe5NbQZkkI4bhN908KSChWNk0eUxet
TIw7/HAwQhI5Ql+ahBPsZQ3VWkBg3j/CfHu16+B0h7JFIYl6dQ6N17OkRbJotFYzD6No+dy7yWDP
ZbBme4B7Sy51/PoNQHXbGeOFFKpga4w8pVTpT/5POEPaVuAUYPUOvjBbjsl/xhi0Ru1morLajhPx
nsZYQLl7XdyXdlWWrOypi4jtweonpCXHcaH1kvqjQPYePKT/7L2NoKuWM6eR/wsiAsN5J9us+5Gq
nhvetAvlplHRvauaAgTsdOkBeVIJcX4bQXgViQWjOknydNbJmUc61DTb+XOTjSQ38tav1dkZAr8Y
mQC/OFS+dw9DpOTlUkggzauU6QIQRuTwhKdHw+j+HYKxljVE614+43KoAWdERoASDdgaDCykiXSy
IKqOOPAy8Uolol67qpYR8qEOeIAm01WqEviQakQodzHSE/ZiGpqusnTkYUqzGOiL6wdM3bK50x4m
kQ7oXT9SiIX9E4SzGg7FFoCcftDwWl5zjFBD4qIfBAuIN3Of6SBQ5XPVZ9eToJDQ+gcUSZt/ymav
2NSuxa3mREPVk/fSOA/upfSMEo9MGaoIXFZ2t/4P9PwikRbmjgnJ9E8hSsjgJT/4mu38sl9q5ze7
vuD2Nx7swO3jb6rNvASo1dyT/L01UjMz3VDcp/SkK1wn6zY6AsR42TPAXJmBlRJYoFTzGYm92pYd
RTBgZ3boaZ6unt7urnYySj7KjZ4FpZJMqhMBaerDaXn/d5axxjpHA/cgROTG2ncREEeWWySxUvGt
QpFjVt/DkuklvKFAJ7ZK2gTHsSgai6DxjxGpF1t4UB5e9YfFpExmPpYZ+JE1kebwCjATgP9FegqW
jbAZbyEaILjpKqp87b81K5NnxPuQVC5JN1d33sy8UigR80eWUI9PDhYwzA8YlNJJMVrWV200ToH+
nVK5lMqCgG3xDp+SZZlh0I/g9lLq/2cD0+MBmMp5jhAhiKNeSJtowAmGS1k5ZlRc05O4ZFfJla5K
2t3TwEbU6S2VcjMdnDZaPGNF/KRY+77LIO34YiUAX4YsMF3LXXK6w3Lb5wIwN79/Y/CzUe61YjN0
BqP00LtKmXamBCHcRL+m6O0hkj1v0PplIk9uWfsi1kF6/cTS4CYhlbk08/YX0TAeuhRnkkk8I3iS
wcrhCZ9TJO5l2MYEjkI1qyCCsE7CKON7vbzTbU3HgmwL3u69w5s0gzWpnrAy7+fhK38UMnWMUBJt
NnN6QrviPyAT3MbrnRqbmKM4v1i5JEmPeEnMx0haty7iNGzPIFDGDdx7aymXBbe3nO9LXJSID8ww
RnrMpRLwqbr8KC4vhDPl21Ma4f6evnhFUjyIFa5/EqhQFclebBNr61x3Zw604+XjN1eEAR/zj9Zf
hy1f9PfG9UNx4X4WdvbVLbXgLrsyzxn5wLLC7ZBVcn6PE8BZlX6EyMF8uo6prruxsqY1KPbc2V/h
KJBkM/bN6Dr8T5ge+0Zo4m3DGpn1sTXj+pJxn2lAvjLTUnhr6cylYTWhGLfvgeYqD8+IpEU93YVr
nzWTERKNtOCgg/pup2vlEaefrLp5b7PbcNQMQfFgZywEgc415JKLvCX6nYMLL/CB94rVCKT1IrVn
iUb+Qhvv8NcBATfSH1Fv4IKj5iASbMQdBMmx9T38mfAr2EckPDNR7IBqtVLN9G1xtDnhS5ljf9yq
Tn+vWmGRRCIdwLoSDOWIqDGFnUHXmtIEJsbdLIXRw0mlILbfBuO3By2Ca7b1hqHftgbaKG7sA6Ri
hVcFGevrWGBDWwKlNXx59NgHagAWt4CnKu4Riq/mn71KF5R5BdSi6yvZH7AWVX5daLCXX8521TBm
ZmWSItuKLiovpwzjJbduBm+VmXIJvkg8alOQS+p/MhWBniOcd7CXOOzevklBJqy4bHFiO4di8j9i
DoYzsShNKisltUhf6tReWcXSZUGls27H9rrNoLbmU6A7Hg5ijStKMsS4iqnbPSGzKsfK0Fvygrk+
Q3F6SAkJ0pkyqkqE1jv5gnpq1taOILfb+bUNKj1FbpMfxGg2q3UzNQUgOklgPcFyAkr6E/j9Cbl5
9DfOl2Qocibwj91b3HeInJUbHpv6chp1SN3VLIw8sNe7l0pfKeRCGEn1QvPsi84sl6pfEb8OYqoG
vUfZB0sDHphYgf2O0K+oDAbbbvwesWdpD44kCR9jA+YyK3wUm4mWJQe/yRNFCq2RaHp7n0JlseNw
lF6otmC9r1W09d/7w7OSpMFJqEE9jiYorzZ5LSV9RKD8D2UBJrcRcVWMm9OUHD4/TDZYaYKqKts5
mnBp3xJu8rF6wtTV3yIKlSjeFIKKrIeUmCQetxyBiM7nOtBxfYTlr37nGT1+YcRJpNGla+B4pYs7
nP/BVw7ebKqm6kDin94nFGjdYeykVPyuSGPWUm8aNMDm7j4oHu/GJDtpZejyQ9+a9yvURRDskWwi
EgSgmFqGJsmEk/VQKoJkvVQnYlpqoUbxt9RiT0Hr2r53i9nIGsaDmnRLVCHgwrfLO9qlNO8761Rw
TyRkK4O5bBE3ZobqDz7DNR1VAHB7rQsBFMGbVs3fo0m/71wBUD1jRQ5KkejfrN8P2ZRXFye3bUvG
Jitur5eOlJh9XgSbCiFI7SzWAWcnMlbJNXYpx2B/M5SGOPb8vpX9reYV5VynWG/djNwipwXCL4t8
T8iLhc8e6Zl92m+CHL3mgAlfVWVRr2sl1H7s9aeYtE1Wm3zVhIQ0LAgCAkWHK2oVsAI6/BPKJicE
BrAtw9aaO5jiKt5X5sSFmcWQ2KRmQuRAG9mvfFDXTxNXWfvgC3iKsNGJFLB9dHQGZJeQ2wkTbLzC
2JtD20dDH6tIPFWgyvAUhZS9J0DgRoPU20yFi1gT3Gxe4KWp1iiGGaq2bliV+em0nR56nvdc6qvm
KG8gjJ1iE7Do0n3clhvSKJM+VVavBcN+4wUyhzis05TJJ5oKtDifvIzisPsR5TLh055RYCqKxR4h
JRdMZzY0TUf3pKhr0gTBwDRCvUobOAUEXG6IDigRWgVzTFznNpR9p1oaGnilW1PbJ3mKY6/WCdZA
gcTkINzgUy+32Z59nOsTP/NInu4pBa9UUDUmeX6G1osfQhbQjid9579bem5zCqzvIbtUVKxIKTNZ
Ng1Itbr+oondWJCryI0uAgAwF03cdh0Y2PIo2Js7e6LPY91z4qegaYPukbrJALKQpwAih7mIADUY
hx4kVCNk7itzrawMXNIGvEhAE2TZGo/eYfR7ebVim6xNBkAisUz9Tac3uDbpDLhAD5w5QbVno7R4
xwd5kmbEkfwIfcYseW9h4A4fqoOkQKrGC8jpCpQh7eoDqPZxRJrH+i7pxSLA5r4ARCsrpDJXkx7G
9seLIsbkzQKgXH6ft0/+ReqX5asaWPFV9noTJ0M0r3bEShRwXd561gunvVA/GHBkI+j/bNX1NWGh
JABlqIk9i0o7Fjj9aL5xdAkKIo2W/C8sV1nu/Dgx2mQZuXoQOFoFawegHeQat0eRynS+k2stcGVW
ntqVLRZGrl/TPoStiDaK8MrdBXlv9tvU04fZ8AxaOr3AKGVY1dHbBlJ9R/3QTVcBQBNL3hkmWZ/c
cG/aGvVlJCN3pDg/NMCTRlpZ68t1dAUQDNU3AX1srJfUmuvS2/DGjgZJkPc60yGqNi3V9niO0U0w
8uFgFy0nxDsr+PHNa75G12p8sIKncuilxAQR+vQxzo2KLO1/7I1o2leKt3T5rpxcA1i+4VZOSJTA
UdgLoQdrwWDrLZYMSYL1Rxqp2eT5JXt4JtT+m3OEuePX6CIM93dwC/AdMgh4KGZH5T29OgojCDDd
0jkVa/l5LvHZ0ySlj8M8cDin83y0J23sQwe0kkZyhuxcWEBGQwR2h6gkoVa40i8+KTScJ/n64N3r
kVRrrA8VbKZSDRGNbTQ3X/Hs2Tj58XmDl7IVuYwueX6uOpzUypKluLf9+FkjJncUGHM/z2rlTHul
tyHUIuZ+OMLxz3zJItcl+t1E4Rwy/8KYz3xNZSdJ5pkWVcpBmxV0GIHNZuIVLF64tvv0jsoQXOqJ
soc1PbEIVxw2QoM+6b6A7JxoREbbdaewLWdToRqjm2gx3I3+FwJYOMsC+wlu2EHe955yEmoddWg/
F6beTItChDw7RtC9goShaRImy1gpcO/gAtoSaPJzx/FM5PpjTNnZtu11CUla82APXfBwaxc9e1A3
gMv641Zy3IN5xSZkNtJ+2g4NFJOJpyHhV8RmkDjZMcuHIj1THp4b5kGt1R+POu/fajk05W6S0NUd
B1/gvK0dlLzMuxMjGT8uJu7eX9zVinyp2IWG3f1ua4A6tOcbvAWeMoWubIqZjllaEgflvZoKF/H1
li+zdTMmRhvqcezxmyhWqQ7l6YuRfGeo8h+X3lvtOyRK+qN8rhrMgimA0la4GTvJ4MVFjuK2a1GV
rWf2No1MaxYftYKV8nhZb6I9qQaSQ5/lAoRdCj7UXgg/5XxHm9IvlEwZPXB7KBP4VpeTsO9v0bN2
zdMhkMa4+CmBwhaxtz5YN/mqs629Udt97zWDD1G0gKUsXEYuq4e/jBf/i3m3JwgiHZEumStEQksa
vB4QYvOdfoJe6K7gwd47eAs9heAbNG4B15UZuEjAoHXruNYMdFWP0sfv1E152+MG1gLGJJ2gSOaB
fHF+3XFGar8zk8W/5UHDw0z6w6SlvhB4hMwjMCrHw/fYJYnbee9lF7eeZDmHiJkYtruliwe+0PyI
8rtAD7UmzBI8Px1PZ3/8+OKbbvBszqwX5CDgpl2ehWMrG21VKiSRbSQ4Ycw7jwwcWGoD5GFJ1jU2
Rtb09Vm0Uqm2aT8sAcmCk/yRmpJv7o5w4DDPv2YRXXOC2i0OQO6i5jM7/UO+eUYRzzh5MyZ3YVDQ
XEIN9pKlsITPNGYajaSse7hszBw3OVsvRPkyou3uYpaF5aFUv7T4axrZeAAyteU8ZY7etyak76FP
JVmnOP2zwMP8qwT7QLgaumjLV8RzhHLi+jKUjEAj36zkmQP/IpvnKbazeaceHcMmTNHrcfBp4wh/
KndRMH4rozRKyZAuLL4VuUxy0NmGGxxWJSKPcJH4VMob8Am/tR0y4DpYDOWXC7OAvBc1TxW18HQB
g9DKO8htmJ7/3C2dk7tdi1ZAPPe2BBDC1CUDmvmLdluQJl+OIviNWSxTfWJSM/ubJXp0oVpeVNEm
M2XmelmaGPNHFDrhYI3w7Rie1ptju+YliEpq6fK4/BzITy53+jq8i9v0wKMCyNu3wWcjMdICLGtt
kxSV4zAgQDIBRG7g7QwJNQRqEnvDk7fH+Fvy+OY3kCNv8hqaBggCuQ5qItETb6QjbgiCNFMITu+1
ZryJz+jUgTZsQEbBViVBdqch5AwpoK5Vu7yvV5kk9F1nCVSHBS/R4ssArHLJIDc6OO1fj/0za9sT
NgzeEzeGJ72gXiFOilRqT9GuaYJIZ6CixbWIws2yPdSVTGfY2L+La9tJjrwdEKcKWLmv3TNPJtov
SuNmfbHeZTSHX6LYE1pAZ9iJGF4CFXOVjSXMoEGwYRoHyrhcfpyjWPtM90PyPsLGfegXFGUB0Z2M
bQphVQCK6p0SZmRNDsUn9ZX6G8dR/2tL5Kn+PEtl5L6FamZpHt9Dc4PvHrbokdsuN/5eOvV0QNig
rtjSB5qDz5ZSQPybPsOLSEL8EPNL7KBb7PJfvF0Nwu/mtie0XBA2+xZ+vYQV4Z9up34bKJzREPPg
Ex+P8qeqdkDDZ/01gBvwQtsG9VGvxHCvt+zU0GP9edEg7gfEHf+dKw4ikh+RQZ1SbuPlhi9EQPTW
co/Gn2flr8GO19Kt2vFYnfETE9CMWKvE9LyfRYns8UY1D+I0sbAHATVzsG8m8wDoyzRkac+Zayr1
PsftFp7XUPtf3EXBJvAeXQSlP0I0iiAw9Cfra3z0o6JNRk8xw6AmeRUpVlLeA71loc0JReyqllzB
nNaSakrs8YWXize97LHEUUDz+VmqaV3oaUNZkSbC+Od0IGBMhNkLsRwOivjisy7cpC/QkzWyeLmy
obGkizsEStDuwB0LSkrb0mVbO5yoA1blMK7+sziRrTcE3AJi+4czQeK428LiHSZKwd4Ao50tzFY1
J/CaeZMY44MA0jNjDtslgNH2BkTum2B+b4EUWJ0An3aNy3B6q1zbyjzKwV3nyV4MLpv8X8a76MrF
w/sTenf+ZyL3Hk5F/SB3GiHIdIJ8IiKs4zm+kF7G0bmLCX5DJAAZzqs0xXzaNRkrgzyyJsyquTyO
q0+2O0NDAHKTC0XYDlUNrmmNQJY9dWq3y++I1eK6w/+9ccQseSvJdgr83satmMbe5fx/bSVkhOcL
eo46bA4OhcICWe6y2PhX9jFcPQFnpdIrbqtgtzkyDaj14pXy1NIUYZE3SFNjCooIxqWg3orz7srg
3KapjOrW5iWWaX0I23Wu5w9vEiBs49/ex3Nv4MVSrcel2bYjbibjxo3cVWD+PVTQjtfjG7hlswgG
U7SFqecNhmMg8eCvGKBlgYmvetndWWIRHbfKiexbLgxQtI+9tEiQt7QgjcpwM/cPGGKIS3k8fb7L
Utn5KnZ3ccCAf1TRAV65LiKtJqfQrw8XHtUnqBN4R0fATXSlFPRzXUE95Tesvli3GDI1tIsji5Nn
i7tqTWtch6uixHqeqqCRQpmvgJzYJEGdK6fnLwCGJ+E+msO1jt1WTKU13Uyt72IE+2VdqtV3jYLJ
Bz2zKsz6YtNQjW3xrgJQo8FVTFP30PJTX+R7LbffErDwyhMQe+jPyXvhkF0c3RwiMnpfSzz/eo1G
rEFdmbzSz7FexQnWuU1jIR7wmIBdjaZdDjoJffQTOwhc89iiwW34Zq+dDgv3jaiaFgivxRSUKADs
FOkmNsIUXvx7/mXcBdTCRgwHUfC6jZFAjKsw0jn0wr2DJjXpiBXVaAm0BsxljlFoP8HNNorFa2w4
2XCUi8u502HYoBuh9hd449DI9wqZ4F8tvg1AAuYa9H8Bxf9YkLz7CVLZueRF9rCK0ti7gJjZFMkc
3MGQI81OjTVxgVxD1Mcq1bp3KlglsjMqmjP+CZe3H4mLotGMy7GdAh0kh/HJuQWom5dJmqxCgftG
xbY8YluX0hTLqKuLa/NRVP51jcNTXQrrH/voP+enP13J2WvdJdeO8nw7aBwTBum3Kl6NWcsvSKdS
odGK20TLuI3Hbs2fT5KTecDZr01QYT7DN2LRCwuxumNb97dCTA9xr+05CoTho6dHRPRpxluu5EQg
doh5+43q4hQGYaPO4xs8yk5KTxDAUqYkdArLpf7jIbQzEvTJKDNaTslgCAb1Yeyo1UzR7E2FsnZE
UbBxNJS0qH686A+dd/evlZgwNu1EXOsSWXAd11XA2R6OPq/Wg9JZCAZk1w7//iK5e1wbTp0pnDOP
nIrwz9oDU0uzob2stsOCYF64nYyj/7Pruno+RUGcqjd/DVSsAJqn6Do2OeN6ZtcvoCAcb389hp+F
zn00hkDQKMAapwfBSOHb5xjdPyFUfZy5kf0KLLcta4QS89/uENaDy+gj3N+eZ6B+kMcKy7lDzAB8
bUGRUWBaEzM8O08tGp1h1WtEhBhB9ELOD1nLl/g53n66SBGG5aYvrf2ogQw8jc0fLGM5txa0KxZ7
mC6FnrAlpo4B6t6y0kgm//9HzZc4vgxnug0vj/05cR6j7OB5HXS2cb5W+mKSzf0mgd9pnUZNK8cH
I90ob0ReBpePlnY97hrzQdWFk+Sus2hDgU3DIkXajLypEtBZILx4hWhV908CcDFt+JC05PGho1Sa
gD9UV9uO9Y1ea4+XborQ159Y9tuamdv1V1JuLVi9FbtwAGBvF2cJPYTXh4ovXxEkUSPWTqYWnD+R
gCmaWfE5EOZyCmTHfz5NtluHzZuL3HdVKalafa4I7ZeYgHUs9Sz/OdjXmTMeomtJeiprZ9uRH/4d
pQkrHMR4LsdEMik3ftsK8Qa0JJWCadd4SSRIqY1ybO9KIfWP5zA6Lz/JmNX+ahqoKyJriU/vpap/
NTZiif4UoDrduMX6FThWzR51CLwkZy6opLvOFIRnwbtEbIFxYRk0iBM65bJ7a1dPvi7wZqrhYBGe
UbTn8wUGWlraykSBrPLrwE1IMqfWDqktq8B2jXhzhiurZwKKR/h0GkJecSSAOYVagk/3+7iPIvVm
KpZmai9a+reJYQjyjWUVODQJJpQCUv56laXojPgXEfQ0G2YVflo+YFAldzPFkSZui4s9k7kXY+zA
LGnZ38weoL68Plyr/xRVTaswqd5ksR+Q/F8CfmHvdD6GzcVLj6ReYZ8LytGZdNiHPPrQ8XxmvfbU
nkm1K7vnRkgJdwmA4nglUlvMmBZaRzl7fNNcqbxklofaBUF9QHFarMXszJIp1mZmbV8+iaSRQxuz
+aLfmO6OpdmNkuT3AxDfCc68wGGN0kgrCHBfJGSpSpl1MpPl5LVwKyooJnG+yreklqO0AlK/y9g9
Ms0SQh7dYEQS2D6SgG3baToEKZPrIM1zsJT+TCZEhO8WH3AdWOdDEDsuIxMh87m8vJN/bB7VJS9L
XASkIhdMpX7Y8NIXbW341yetVANKMtCgIcfwDwfUxfjIkB8S9+/KE8j1Rpf/8Eu+tr+x8IYV5Pea
sk7rCHcE+e/C+jlKFLO7aRtlgzBCpWANFgQzP0zEM/fkPcnIxrkzc7uKZIFFyaqhzE8qpZX5rQPq
cKp3hgGHZDNrZ3yzPbkQqIJo6122S2gRN5LKr+NRrbHQXUwRw+L+4olY4CANQxx+a4QmW1895lTQ
uZ1OJx4BhfpBYtYbT7qKv56uXsFSw2OHgynOgxVVVpoeLDLx07OpkLqn/EhSlSJ52Ccbk0KhooiT
0PIZhkgyDYRt95AZc+ZIL+qNodys4Xcq/EyVWfWlkCa53NhbEIIRkXrg3EHj/LcdI5FIiP8mgJW5
YD3lAvBeirwm6pUrpdZ+wR1hdcck6a337uAiKRLZBFuGwxnk4n6VfxbAKlnjNiWUCwV4sk7CWDCt
rS6NbsQnaO99y1OQqwOlUE3odsknBdwJgo03Nbtj/sIWt5D25pJAxlQRbtt7yWkKcGxxoIQv0Mhz
vvJZbG3knHwSQ421YXAC64GhenKmJ80lpJ3Vzn+JoIKC/qWfXbmRY1fb7K+GraRgYbjxut8+q1Sk
MP6f1AIasgjqTVlP1qaqe1a2AX0z0GfYOMudWOVr9m4ip3tjGlUpJLG+ICpvxweRP7dZYrlIbn/R
FNNAExIXFOTwRxulPyqQY8OpRjde/9cVJhMmmD22BoLU8Yj+4KS2pS1kh43+++VKLQvGnWYlPkGR
YjsKxdxN4WBsvksZZ9nK/SsU/vJ8ubFZrniC71d6qth1CL6VLPp4AKoSDtycnIe7v4LLqurzeBSi
KsXs03nCi6jHKYFExrDDB0TqBd2ALureVcwlArR/P4SwndRrSwZ8Zy56lrChi7GioVLYsWyLVrqu
QzWXBTFzDy2XOmnmCluUT2T+NtY0AuypwoCZalvDPNofBco4FNm7m5dAIzSchGeYSiYJgf+WVvqT
PAY8rfov3m1FN+CTN/hgAiKSILoJ1SiUgcUt9DvMz5DJ/9mN6NBP439e0nQQDswHKdIl8IeIHRjh
R/0okAbs/Z5xcpNL5rZgnBfUmOBzENAXdEDqKlfz4dCkL9QJrmgusWOmv5+FlfbbHeYq1MCSajJ8
JCeFykvGU55kCkRDQjJkRWLkFA2BBZye0DbOM9BrBbxquvcz3xx2CAr/LXPyMADame7N4gvU88lx
2XPyh/a6GXo/QYJHX9tOj3Ma9p+moxOJwqP7VOR1zGVwipyHpb0mDm1KvJi4DrkaCu1AKsxqMkGe
I3FkAXRuyAjk4flGFd96AF01dJ/zkkKC5F5Hi5a0djTbunfK/4oB2xeVY7L90QF3Ry7go8wujB4I
lnWy/AQ+oQAKnN9YUa1BbuM4Wt3DR86H7wSUsgPpIpeyoxNnp8bJFmn9tP/gW8sdAgA6bE8Gjq8z
e5ge3vuE3Q2lsWN+xsh9/zlQyFOrjuZvfFBZ7CCA0jMtvlMsv12cmc0oUVbiVTzHrY8LuBEHP+a/
KwzD4eskJdwtC7Ozg+ykMGUh0C6ifx3k6+l37RiWqelJ7vGOOsqZps9FVz76thadneAUUGy7rfdj
Di/My0TQf/y86mp80jdazDGbmLQA2uNqLwd8TUkaMKnr42a0lVdFMoChO7aKfv1bHQ8kVXa3V/9X
/oRfi7xWzmmrcii41k7buxLLBmnRqjfp0x6s9wTmtQ4knvGaZeXfEoGpbo+X4JCHUgnO7joGrlr0
1pdsLnJtRlUHTGrkFMttXcProl6Zj+hXX1UYUaKHSNz9KQwe8htuDlzu+YY676hFDdOl8hN1BZWU
5HsIlIYsC1BwT7hzLpH/u8Frucdr8vfGylSWCZT3UfOmPvXX32Hg7ZidgAG7ZSnhdR7ybQDrfKh9
xI0AalO2yhgFUfcbxp6I0ZP08srUzJvoT3VYvtpt0pZ9agfQ8+MOqAWja2Xfx08Wel60FdZOVrwP
KkwDz0b1b9jnHX9mON3nCXV1VUBh9da7qUb29xi1G+JanuL8NesvGxSNELzolH7B0COSeGxE1LV+
CTg3hphfS8H8F6YXTnqPi/sbch2dRXzb/XM50IBoQhFV2aI49N3OqS8/XX+d5r8HvNBSTk9a11vH
YB6yFyCZNimDX67a6alklGXOzzC51PY+DSEQxSLh3G7kXxiW5BBqpPUKrdCgvNzh7wX1l4D2rq3e
6lSOArOpUyKNrmL4n3A8eFoQV3NzaNqN9P8xfhw2FVwtaXaWRbFAx64XspDBYU3vY4DTYbDjJYaf
PqWvbDMBpAqWzY5+pOSiIjc9O2qOYj8snnvw7ZsKpCNGfWltOQrXIup3P5Hrr2x1HhOxj6bPGjEY
FASejJSyGF4TnAhEoxlwk9RZNVuY9csmhABYPrHBGc2iR0Jcu9c+3xdeMqGLiHHWQVifBXJ8MQuA
ElJl2AO02+xQMPdi0gfKVTE0KUmlYVyDbqkJBN+WpgoOEoscQ7ISZNFhIBGeC+lTvLpoe/qBboI/
XRAhdc+nz+izPWSdOdEERtU/h3qr6PMxnLw++bujWplqTAnFLj+ptyIlX/PYjIn+iIIE9fCv0t/q
F+Wx0ZBcznHh5XkcCUkaGFB9bJJaLWZJQUxqOURn3oCMt29nsUT8Kjdw1bP0C5FSG7KMrgdcbYfh
jf6XDAJ/comvPcf3F/47j8XlP9iwL3ZMwFTpPKXFl7MFvbbrHv+3FfqB9bW2+8xOpcH5NSOEfUY/
I4Hc8bDAQ40blUlj5ahyJ9lCqGDOfPWIwIGh9MVK7W3fT2PnTj5eMMGvmNUCdHf31C6+8NFEhti8
Etkb5RWKywLonlgKPgHHmkeGVNUVSGUjCiQFYRamMq27o5WiQp/32hz3xmyOpby5BDflQgUz0M2t
J+Xa2nYT4l99Z4rnAFoUoVl/XvE2G6sxfgkmig/Yz5S3vhE8Eg9h6gf6ArF2OZSPxOnGTpTWXCBK
I4MWvC4etkuMsScEiqs36+3uAREKLNbE+XeON5QW7x3Z90+sgVPEXIKDyBj0HmQaSN0jftRx0yf9
rQWDb8yQkPIwLz2X+kbsrhjYFnTirkttZJmRYTGCXj25a9SKe+MFV6yBA2DvRRPyabcXIotuoAhA
Z5g4kErYVrcKTKHl2sZOVgu8VyMZ1tqhfrPMkAK7pG5oJjHx1f8DyrlO+NGGhwgBZ+dUCuCCm7I/
aNE1DnHw+zsrPXtfm/aJY1ic1hZeFfMsCyiaCgCsTW+nM7n+JpT4IvVXPor4A3EjjkWyBScjMJyb
bOJo1ur87/inWgjEeB1BxUQuomQlinhpEvTVVz8YRasqHklNU8iAoL8ch6xe3XHMP6T3duFSsGg2
4TbTSt21nxTOPgH22+q1G/5H6+cjpdG2HzDeRQi6FZGHlzH8Lec1ukhzI1dNW2zyMm7MyXvdNlS9
4RFtFxkagXtMaVZy3rMpg3VYuoaSoJPXyVVBmANbGmiRGWRc5ng0irtQPT+P4vx7ezJBaGrAlHi4
/t6BXfCSEV8ywkyXdx/ZZaAiogw+4jaWICuXJSRsvIkGx2VG5WibMc/r/zbGgry66FvOs1A6bwvq
Tx/WuDXSbgAd5RVxQZomcJlGgpOrL+m3nNksMpfRHWHdQ1q0Sq2qNfq6HB4Ejvm5Z6LAuMiNGfTU
CsKo9LmxEJu0/gYPP7naxwJ4I728Bvj3SChHZ1C047QMPG1gcLcUo4Vx0aVW3NXvHr7tRln+oSTp
3vxSLZ6kxLxWZeoWt5vNi9Fe1OCnAIQJLq1OXKadBcZQ+nnUg66091+RdfCIr8r8AnBD1m/Ox8G5
shQGUM2byspTr4VprsySTihJxYvMgvSEmckfpWllJ3kqJoAYYYuxlQGhNu6NNuuRC/jZdtA/JJT6
vnlQbiPpe7Ut0rg8CEyPePLofeqpGZF5iFlPUzc6VMDymieCwaK7bwsF9nrSvhOrWt1Qr2pepA5H
qB+lRqESCeHs8U3zwjweheYMcXZldcD9nC0J8HkxIf4ioS6ORTcml0LwuHrha3yMym+YtiJHx+PS
paH91MNndiVqJ+nTNhR292c/SjBtbdwzmwZl9eXfRXd657o2zLsCygAQuM6Ve+LLJMOcr0+6foWk
Pa4cMCLod1DR1DLif96zrUB/CiImugHhNSwBddrfjo3AGhMw0RjkRTw47lvWhBTbzFQ2Xa3w/HdM
8fibODtuSzsyh+AI/8/PIYbQULo6GjW44LiZrd/d7RRbhgu7JOSWrzD7s3oRxDUB3fjMZlWeETP4
FkUmE+VbQyArIPJVorzhhfVGg2AAHY6uQt0aGKeQrsvrBKYnD/QtaMZ5JqNV/treL87mp8zVOOxC
6+ABMfi2A1pcRC989lWsAwl5iAypCeq0LhRdZMFAiv3Skli6xn/mc4M7zgJmJi1bjkwIv1KA6tzr
Wld+FqxMxQPZnVvo5WihpgCFLvEnZ1eMFzu9TZZMU1YKpFiSeL9CWnLck70OlA2M/GjgoUL1t71Y
d7M5xKI2/3ml+51eESgeGY+ViudaBBwROQqNcPcMnVPpBMYIo22h925YpC8jiJQvYzMla+amH4X6
sDWRwO8DEVBizdMXeKg/zGvLETWyl/OVUuWamrOqTcqKR9vStS1eERoDb+uhSTZc21r2nUXk/JHp
A0t0c3t1dImEyXWcQKoBXxafhP982nRcan/XQNfa/jJxCRtqlBsJnAvLUqcf8oY11ni25NV5d21E
saLY9QcYvRNV/Ln2FwuZa5MO+EyvjfTdBDEgDEEltvQehRQ4nbnp6fg0PAXEjkMZWOWZnua5c+WB
YhLivMIBMTFQxbbqu9XLlh4TGtQCZl4vrGdnTK6rmBIyNUS0ZyA1ZuR5catU1VLs0iz7gydWTdqS
mhTXfjE046H/bNWLVjcgmXwf/QqhMCrxWpQaiMZK9qTvb0mKhaGLBsU6DaIYbWcsJlt2ET2YaM+N
aB/MFOBiPVLUSOeUpUEmtw//7CgxJvfdIFInyBubqZahGkfVFW5XhKtju1yiSB8WPfRFalM8+ZY/
M2GcrMNUIuKN9CvSUqo5YN8cDm/a3+22mPhc6lD0PZOhgDciW7XgAsqAWgblgm4yCYHm9RdNxDS/
nDGsTEkdgjGMcSrygJ13Y8iODNzvWsWS2MT69jKxqW/kqlF+bUveXYCaq5pfeRQya/W0+boEBeuq
K8CjOyhTP1/VZPhGeUNI85L/QN2rfzhZB0rk62ln2W3liudQvZGNQ4CIGz9j6u8gNqClktdym50m
QN/cqrtX21N0teHxLTsW0cs4W0JynaKtOZr/XrzGLxbEgDJw0hU9yvfHjyxaRZ6zKk7bBK01p6Bg
1YhuoC4EXMYKwQ7O/yZyiFaThgRO7zWMDj3sjAZ9tbaeipkEZyweJCtOTQ5MXuDKFW8cNdm8RsPC
Jr4eOqz2F3cGd8p0knU3ERTO+SxTj4d7tmc11pZJ6RiMbsFPdH7fbUEMI6eMNA8KyyI7+8npH1UK
JsSmIgdtyXYJWDBHrywcrtbw+MkzXusdK/D7A40kpYSACnUeIox6mAI/+YNjqwV3YGNdL9he3qlc
Jh1ICeiOkqMo5g+ySS2ruGsQJez0Jw44Da7WGX1NTXvWntIpdVBWrc+RHxVuFT0ZIFz06IyOqXvD
DHw5ZU8OtgsxnAeWXfNfTCB3avt5gL0NF68ufnZy9QaoJEnQWTgScBFy9GZd+XyRVcRbfo4KlAPK
mPvoHudIZFsxup82XmTqxElxazs0SsQdb9wN8XFpyQlUjzEsPl5rUjB2y+HzirKDWiHVz6EYkV5k
kaL68TDaelOYORGVEZoGenkwJspNxVfUjnbMpdQpVOtcDYwLxmUIXY4mufMqk9WpYSy4s/LRlJ/e
0EHmNiebhWOe+506fd5fiAc29eN6IVSCx1mzifoh8QZwNLg3+VZr+Om2AOyCuBg4D8GXVS8+caht
JAdEmPq79lQQ3spcGrEE1EE7U7Lh7P27Efozxb+rpRyoANEW+pfcPtwZcj7e8yw+FJToijYnYhuw
ewY3OSR36D9mOKo1dwX+cFpLdrQp9+tIG8xctBuVE03OpEudffBop3wOS3S8uUC5N9pUADlbCElh
9sdKzNAJ+uXi+aff0geKdtQiOzSn8hGh3zpRzfOhVYoDiHEJeXiaohxGxof1z8X4O29tFKK/L37b
C7sJZfD30t2PXLfr5bVC2Olf/74/ul1Dc8UwO3J341EX320Hxg/ZuWLEDatwiEKhnPa/afZLTuMI
EvTr/gF3do53cWbHuJlP85aUoTgWb3GdpNVWc17QWVJdGyx1QJWq9WX1XOPapMXx2k2t+N/Sujcv
m76ueDwQJ78KKB+y3QyIdzOBxI35o+1PNPByycjh7imHU0h0o9M8w9LO5IdpBkTz7XmRkjqT5GIR
LThiqJG7zorWg3gGoRf+p8bQF/RSj3EVOambuxmkiXi6Shpl1DgLZYoIvWskaY57t2O7QuBDVNnF
7TzTIlyMRO3Ve0+vWS5NGB5l6VxtdTokJgxy1ydvqJ5xxrS5qner7CraJ5qOPNmBDTon9b0OdbfE
3DANEU0CnncTSoJQF913uqDVfY+cDqYytRGKJsf0YMJGKP67WW6+qAHg8GHTPftbcVRE2k+S6tdo
CQDIEAzDKofLLa2Otin+rB4fLKi0ZgZVpu/NMiof27x6FoTNzLuFRmkecZDuqyvuGFtPn85aTJpL
GEG+i3cC4ISiM6f7iAXi/gDDE5N2F6U51Tw+oyf0rPKEkIVAGyTz4+XmzOA/FVGnU0j1e95e2+yF
P6sKSUGOsQPkr5p0uJ4VezBPJ42/yMt31OoHqI4zySeE042ttEXpoxqEvTlhWfcOmO0Gf8bTP4Yh
iqqKzDWcbvKErJ0DziRB18mQfNT/bTm+ewNbSFjU7RBYPDc9ITCm5MjY0O4RRbKNXbGeozN9oPsn
vIySePYLS3oGD1ki86fi+TKuEe5b738HmoTYUbtmoG/yvye6L0Y3mehjWryrjSBlsg+Pwzr03tGt
H5zj4/n/mvNNmy9vfrOtjsENiwwckCtu6eDDt1WtqqRLyjSFSasLioKYb8Fv8nFo2fMls1UKdohn
B+miAkIDtLVsdO9R/Gz3IWiSHQW9HZi7Uv5Lu75HkM69UhMdI0Yb577wvy4lZBXVD/VIMbfZsjq7
9te8LdkXaKDfper0LK5UylbmB7mtqcYrEQHSV+LV+TK0j1fsbFw/Kz0c7oX+hqMZiFK6CEsVZ+Ms
j91ko5uFLi6XEKYv1zc8QIUx9zdOsFICF5n8mg/NdkPTnOjfYIWZj6h8vHainSkEdKsQ7ZwNBMzG
4TqUi4f+lg+2qVt6C2yTwgINRMwwLR6ewUY97CPhBB1g2IKt9aLsLzqfrSfOKRBnDYTSoSkecs1w
6nk5w1VHUAQwaFZfE9N0Rvtur/wsDXi4LOg97zkmw2MJLV0g+sdxB9bihXVuLAHf5ZSg78utoJ2a
GiK/hBK1Su5Wy5YxHG5iAYxCM8EwMwPJ7dO2iT5xBR2EiAnbaWd10pVnPdjxYwK2Xw1suT1ssNIi
LHAGTY3fikh8htGXqmh3NJ0z4JPPGnAjRvKNTO+TnsjBsYyjye+Gt48fKxl/MIi9DdFJYNXWmCbK
2DtXCkOkQOWsgJCte0xXTIiVwoDUT5yk82Nx0N5u8w97a0vy1kHE0EmgjwdHOrBesc9E+4GivcEY
ZSSfkVs5w/V8veSsUxAsqmLcdoR3Q/nsh/RRtpRq0Tm3Tf5xDLWKEhHON2CgpLG6L9ACzHanDZ0e
O4dRXJOfR1EjSrIzWP04dOoBHLBFMxCCVLoX81EjWWgdYOEQL6173CEe/tIlhzgTNK8+Pnq1vx4h
Xjv6AGR9792IJ2tw3Z3ZD1yHyORsE5foEYSKTai8PwzgPGemXCneQEqh6heHJe+qjGBUaH7d1uiP
7U7v3KzAh6TfjfC+vAVNAOOpASvRdaIBYjbYBOCyCG7G9wa6Wjzxh7Oo/vMRmNuqDtq06Q6W8e+C
4D9RhE9IDM5EBNybQu3KdSMY9i3Ep/Q3al2NHYrrDAf1k8OrsacORSaqpZ8W9I6nlxPmau0XuibI
hS8BqakfgqT3/v1+QRKBjMCrXzBaXXtjG5y7DDMCTHRdpIhv2yEEfZKhA100tb1CYxFo/PzzcbYw
aC2oMuOmJnFeQ4BNX/ESPljx9g+hn7QTcWdH4YXXBT/CBnPxwB6aGRVK101MNUwO4tw32RNVVXKR
QU6WGN8QXeAscqjcZ/r2+g2NSDqJiKzL9M/fLXJunwTFhPrAVV/uidFj97cRktJy1n1IRZDYo6Ty
eWmTQ9Pn0Qp/Qsi5/uGGqn9uoshq3B47lZE8BW9GJiyhZA6aww+dUbDWQ1r6tMVfFDLx/iyzuXOU
yPNIZ74ehj3DOM3Jyx3pF6bt55/Ax+EwvcLV4+mukt04pcU7XCH3uLMMMrCeCNpS62a/gyiTCFFT
upCXS0oAAw8Bq9LSJW0U0WSf5Hrasj6oydvd+uXDJIy3oV/l43KusPreLp72FhlQoDZeQteXdyTv
9f4HmNIQsQx7s3LH+cI7+ijpdF4sA7yrSq2JnBmYhNBtehHrMtVctjS3sLRRzRitCCuqJYXvVHh4
i6zeKBhvVQ9Fg8oi+9QUvCLYPmjOH/jNBfyCa9E+LfUbMrERVkB8F3bXyTo3EtxwI3R7/f953LFI
FPY7BRDk252mccitmVIHz14SwrdxikIwaGWAwdP7syrGOii5R2LROZSOoVCIELm2v/OWvIzRQrQk
BRBfRuvkUk4KpUhK/ljxu5j0rM76EvH41OxIbUwpyGCvg0dPzz2H77lhPw02ChXj88zP6F4xySOr
Mq5orFxpXe2mshuJvmKp8/BQWArNqD836h6nN8OYszfKbzKvEhHLgOkitw2wWY/+XLiQ2CkkUQw7
LicVBMuRNmWOMaTjuesrH8f7NiEeVgmmHxl3G1+jkUkKkyWTVbiWFrR4SYKpkaRn1M970KeOlVsB
i+7GUWorqNiTkmNvBRRWyu6Jx44nH7cxyJhtijqR/xmpKM2O/m6BMHMdxzdKeLn/LhcsUtWETOir
P9gZctDpHaKd5PbOMXqGqLErv82Tte1KaFFY7VEz5V1V3AOmOpPV7DgKQ2OPE8Y3fSUXDzCDg3XA
yT8iHOquNF3ewgI6q9GrJ1Akc6DtpLYpgVLsh/PT3hiqUadUwlr0TviNiw5fB2orULbEf5emuQM7
XnB9h6QbAxrSfbaKJvcpu20nuXf+mRt5dxLbtFr9e894pS/6oCjJGc3eTcqqpVBnbo4DvGjG9YmY
QJvJNm+7itC0huPKlXOVPRXptKcVg5UzerS/OwbZHHbnIWaF8pS6r5OUKrCL4hs/Z06GubHxAAdb
u9u3vjwzlNVfro5p8LKYtZaKaDeaFwuTBKyybVSypHvk4yASsS+zbsJaXE6RKAXwDl8WQ57de6uq
ZskU9+Z1RaXkHmFodjawZSJcLHOmho2zbEGOBSciw8K8QuliDkMaM4lQADlIex2tj2WBibQRnDZe
foxTqmgdCivZ8V43eTOsCMsWRa3rvrcHFM4UOz3Sw9jO1uCgW7Xj6xp5JoYIkH9HCRU9cc/qYXRJ
6aNkyUAnxeoe7s+5JCr6HVEXmQjO61/l67945QooZIxpCp617rjvgJE90nHPdX/3rEtBgdOuWEia
hEgWBLxQ1ai8E38RNnZrZZOKizBAkcwoctdm10aWvrNmHXYIDHKqSslnZeADsz78yv6zdQN1Y5q6
5L0Yg2FEgHHHqG+3XF0ma1OI/mLiWTMw37GuJuWVMKUvwxWhL55siYbcLqrdkx1MfB25ZFo3W2U7
AKXC14ZLMRCImUwPw/N9cy9jwlqVDL8OXUwTHeB/6kTbTqerX+Z6eiw+yN2aPcxoIlxVichfd6Tx
ahjXLoqQglSpmFwOBm9x0CA7giyQwyA89FGAwaaOXCvE4jtGsUmMdTkkTuae+xJGAnfRr+3X9za/
oeS7jORXh0afoWRder/w/CQEOIUQsgEFkOKz/e2DvT3qRhjCJg7LJL6sy1lc1CQdiC8xu2VJd4To
LkCJ4c9MyBA5HnW5NIsYq4OPNronSs/AehjbRtqta5K/JpguQo/Q0cfljmrhHINYm1Ww30W38+OO
+LUQGZEIOHd7QGixjuZyAMx9VL2nto+HHcEAt31FXIDk01nem1K2Y3TuCJakBn3BOnMwHgLK7cqr
ZW4Trvre31+aJqr53jeLtSg/gwQUuMaldZ4HazULJxUlBxNISNbyGr0PkUY0BOrZ/IJqCqX5UMIo
zYuqNIIAjrHWVCJ0Wvef6GML7ASk4G4et0bnDsVlvcTxF4lVifTt4t+SZiJ4Zub+vGf9Boh0wHtB
rFENmHzrarwFosOvA4qUalB19BnqeWGLwKtA577TRHtpmEv1zH4MRrEIiNbp64tCf6F3yktfZh50
cuBuVY28cSDpAJ6TzY0bNtUtCS3M/fltGPMjZ5Lqy8BDo0QCPe0GRZHdVdMvgFocqtF2HJmM0QxZ
b1Re+d1+eSkfHzYCJoNl91FaB04nvifjtP/tC0IS5Mip4EzIVrPH0P0cx77b1gGmWQ8WXjhORX6W
+DskFR2Loartpg2qhoHeCab6o30mGhibmSzmdQDiGWOfl/W+gYwJZ6qrWs9u/BF2JwVSuOhNmtnt
EiAh2QVGhri25QwFret34u0GK28uTo4nPuupBOaGelBrvtuB7IvhnP+KSNvzio0Yd5aQjDb5hAck
pEN1oMDc2cX2CmFeQ09P3jHpWi3LXN9rm6gn1KcRXMEc4E3ez7RHGJ9jQvz8jseMo4nHCkPFzFd3
Kxq8KBirSEi1pCyKZ2DP/dz8bPywlNZSG7xYHKejIOc99VaxGbjJTt82fqMjnZStlTA0beGS4bzA
TNPLjnRRfWE3qcxJVzlvO60ZCM33WoMiwhC0vxhy6LKJZYJLNHubmfKi+1e6moFZP2oIO6aqUEo5
mRfs9CXia223UKM0QX6D9BD7WWi7q3FdNGWPIuFMdDWkYIIRwxF+SD1bNvIJIk/pmDQJWmAbI4bf
gXDaMB0iVcJ28N5zXoGzpOjQNJHeldA/2/eTsG1y3o620JniQAMKEeWFJfa4yBSsQDbI3+3QeCC/
GI0x9066EYBIVCwb6Wt52Y/Fhi5Zdh83GqHW2fo2BVNXh/A4M5unX+EPmDBDCzO5YSzGI/kmrDBe
OEQ2TYxQC4NK9q/TtDxzty1ceBORXoP85/ZWoUp6t4CmWzhYW2r6QYRm9WIVlmRdjnj4aAVvWVs1
7x+1jiGmnw66CaKna2G7xOSzr5y7qcCBAbUh1kUp3L8PL1esAjUBZrwnrgGRyOUy7r7SSCEt/pnj
0HCKzNbzsS49vZ/l+NfrVnAIs2EdlrNWjxVklXwhxRKyDkFlpl8dp0pCcVq0UaRbs5ZFI3LTJnhC
jfDq6UB4JXyW48EjioZbC1KPQufvSySxLfyu2OmI+2Sngu1VA/e5dj2PTn3atK5dahTOkVNp4gGi
nrxSc7cu0go6HqxpkRueZg2dzWPnrhjGbXQdZtBuHZK5guSPQdTTZPxPaNKf56jpLsw+s+HTxPIO
zUcWHOo35i2Ajn4zS+R2utjsH8FUnh+usIWW11S6nrIJDkItIgSwUUQjv0vIw+MhWRlqnCx1xsSU
nUt9W9sWpVhwG/NstMrt3szb22qCTRRW0LcLTbn8Sto7iOgrIp9xjoQnIX2R3jZbro9WXsz+zVV5
dEZB/Q7Dtx6Lh8wjWgvLNhkXQG98GtNwJb/jQL2Xsauc9g5BWjiaixbzkQur87ZWPrKxoWXzyrAw
1PzqXF2fGfAQYwvJ2w3xFBX2NsdyBPlQfn5JxTQ8gjnTO0fw3NISBjMe/FeepINJEFXEgXsyc60d
ZiwgOEaIBKP0zaa3vk7F6TXMeeGbWe6wa9h3WfM//4V6e9uD7SqHl2PcJ1pwmK62qKBYBZArHt/t
8JU8fq2F4DIw2b+0qNYtvEOk6m9fQRNxjrsrRzj9BPRCR+8fjR3iV66CdmS9tckIN+6AfMuNUZN5
hy5yCYoLAUXAwqFkwt2D0KdzAmglVzbnVmF/M4YlmVRxv24coexWOZdMIRq0kl92O63B+5ijVJlJ
3zyAYhSKM6Cpj7wKJnQGdkJT7hIYrAa77KFCIW2DgkGXzQ2monddZ5Hf5vJLHp5B1zBdT616a5Eu
ZI5Dr3PnpkIyt1qDXZdIo0CuK55sC4WGK86BRAooOobLx9qaTMv0NbcoFMSs5HG7HsK34McveGHP
GIuWYI2q6//FOQPbRX+7dU05MfrdVop4QttD62hR5B6kg9S8zQ4lKT7BKrkqqikvn4+WxDlE8WX6
ppfARFuu6BFnCrBp/uzoqTHET5bYMPsMlynf5dw/py74Dhi0r1HXUjyHxH7hN4FvxuJgWw4A0qNr
QXiPRfLWHjGgWOuvE/IYbpv3r5VA5wUbRe5W/ZcYC77Ip4ZoXT6Ai6OVDGyK+NvZZrKm1TjfKQ1m
FhBVtwDb3I+8DJmUkISrundo1pmsCkwlz8wpal+UF0GGwzDVxQFpzlvnXlaqjmWksbvescxv5oV6
XFt7bO4YwedU1G99cbhD1hluBJOiU7kWevAsVDxHT40rrqclM1e2a2ATdot1vRDOoP+LkTFV9qcE
MlkG8YDfrr53E06VD2HTGL0KrVXAgCvjennW/cqi3AHHHArGqLOAoV/AwQyCR41tcE4xZ8Zi+eXv
SDJ8EQm6oy4PledHDFo+84FDXXyLcPVCABmsIIcYtOjdcgPEQdufzkyurz6p0+Dv9Y0KACxUVVEs
yIuJTlUSerDYJCIhTpl9Co+bldrurVn9aVXFfJzdLkpfCxSr6o36HRNR8SyZRqdw16OeANDk4z+3
3aULWz/46Fg61WcZbbJnfaqP5w/ml9VFfpcr97WamSo35fW1wOhY4T8Lo05G7U4g5LKK5qq+6kI5
lEGo8j+IvincObP0QMvyo52VMK4p/j7LEEQ/6dOGvOu+nfQpAptWTpbKxIFqNVPPnnEbn3LOY46C
Tu/1RR9SiMxGi7v3sNzaFIj/vydJOYGFxS35A+VVwAbWOReK4rbuVWuo3u8nlkCzWQojjt1wqqwj
877iQwgmS98DrgYfzClaKoczO4aQiTgzK9g8MuNKakylb41DGnoLpn1p2zK6h43TCDz77f3ov5sA
8pmqjwJZh2kNamzijqHPWpJNY9Dc1cxMaVf0gHg6yeeWcHrqdIQ8DeSnt2Xlw7lVBHbD/HpO+11o
fbG4abo04ytWE4Ro6uE42wEUmzDOPB6tPG+XJoS0r5a//1/56obU/Lh0Rujt8qApGbZpziiuYmSP
UKTfsHxDhWtSKzhkhBePpJh84HSAAQ6R2i5O50kfSpUGlXIR0dJTPxq+d7gSYuQLiOnYYDsqpZ9S
HOelARQScJbt4tJqEoTvFfjbjeG4YRD4KOwPSVBxCUzGvLFds+oYcNHu13mHGebQ5dkWXtADgFm4
MNIUXwK+MlEUAtFRF/9Ea33/X+hHnLAAgUaDhsD4J96xlwjm07QfsRsSLMwKYB9lKczxpwMo5oRN
qpGknG1PNii8pt2ei2/6tBBV9IMEuNA5mUjqREB1ksY1GQ+NBrbF9AURC+0V7fHvD90q/InoFMw0
iPEp/ejAezOgL2BkCjyNlQCe7tYmM2dkjZNLbKKOXZ3RvIrJi1J76sq2VfuRfO97Qhdgn2mMlBtv
4wJObcz3eXVv+WvhJbBlWiH0LhQbdwUY1HoXkYCkpzLfG+esYl6uXWNKbbnETcU0L/0RhKx7IB4Q
SaAv6Z3bS+d5UIcqicYKH8JWpFi6I6k8IM0Sk2EJibzWMegvtmL8mNCfZWevihM97UCt+LMEEIOA
RfA6od+ZQ7/epjik9hON+TGA9KVj3mVYsBddEG5Mo+yxZcUEMMnctgZtWm5wmhJ9hJX//6qPCpuw
0rOt+YseWq3isV/6Abx+u/2KTQ4aa2oVnGztNALw1CHnBe7Y11k9F9emNafGE9p7CRAJJxZnatwM
IwGHgRqdnBckANcRvN0tZJ2Pj44yjLSZZcf5wzQk0kHr4RFuqy2e0kFzBEPu2HY5SyrGOzCZD/P8
LmcNrbGTvfvTXTYSLOELswmip6xc5f5P7Y7c9QBV/hXehBUxqDPx/Lcbv7wTWILBDLT2d+PQYfZI
PytndczbGaLywTvei4o5uxCRwWveBvn40INAs5Em0wtx2ppzb6E8iNg5OmTOyZvrlPETa/vyqjuY
Gd/7VeYH1He6VuUqUE05K1TNendwqc9nVpC6qqXjpe/mKrxZ9eccTtfcHVNmKpDitnhFnBJ90hqF
jzjG2B4RDtNOXskDKq6O7Vh3pzgds2XSvbYktMUeyZIETgFsd1OYttpjK7OVzZRJtwY6TNZI1fHD
SnLmUDWf1/DL1p98y3Zrjg98UVbo+SOUX1M5ztj/d+RgUqz/qp3FdJ/74AksSnxJqayz3TbhQAmM
gj8Nt/IbO8ky2Pdc0a3DgrKnXCC0AXUvEjh0bcHsVhPVbMsu9Zw2+E3VmEsxWifrZauU85S8gFjS
csSRq6PgEXdem+YEaMLg7bwFN90iCplcJDsRPIYdt9N2nlCZ0eNNG74VmJbDFdAitxXUXCqymJbV
ld91yoa6gBSuaWHut4msp58DlQe7nmd0uNze80XQbG/ZCQe5573/a4UTxPlNASAxbzYN072q0OUZ
GfKI/Y5m5hWeg6WuVcD9DS7/jXPQ1v7RAvwjY1F6Dct2qwEPX4UACccXd+CA+T2aJzThnHt4h2Lw
NDCqMqVSl6GwQAqidIdOIc2/lFqwNf79JI1cD8J+Etac/YtLAUMSeFUxt6Pmzml4r2s6Oz++wd47
fRYSFAOJQxJlM/aOc7SWIxb68FojybOyUYoA04/IU/yq6U90TOIIqTwuA5xKvlkzazmWslN4Vtgh
pagmOBvssaBkgQ2X/W41/y2wvyxdcNuKnpuY5Bzo/pJMvdORsAPcq2DbAA9hYqXJ04OyFUj/OQCy
cT3gOwrITp+BNy8LkR7saKYRbycz8yGERZr/RBfCIaklQSUQ0xwY+F4tnFjHuAlnDHnRz3K51614
66U0aHwga0g6jbcUyhGRoO+mLUofOQsqQ/1v/ebskf7OgkuhXE4PnQSdjqkRxpeQ+R2Db8FuSru3
cfIaCHVM85kbpxgQZsWncJ/5ukeGxwEIe8W8ftQXhgkrM3HWDmwhT+tV++dj35PkFS366gB70O7M
T3YMPGV5hXlBZJFNQW72zNRgDkArzRnNJHB4/s02Cue13gOECwTINWuoKimeGtJlSSI7//7QwQYW
mOANuAZTnsqGhWYQcaXx+hDcuzG631akZPmLZZFKrd5XX/1DismjZ6kygkRaadD2PFtnaJzQ7BRR
uKR5KltIieqScSy21HWe2zdPV2ZRC/j84i2mr/tp9uP+/AukhG1veAz7IPmPwQs2azhlUUx0oV0G
JhSL18VM0WRtB6cOLgFBQ9y9quCu20WaN4YAmJqhUZRWQc3wsinMqFMlUspYuuOkFfGxWvfDt8nl
j+1VkcBRo8uGnEScN2DiGlCsxsOW1bXrJGcNHq5rakitDlsJ0qzn9zT5tzMfMOvHV5WEQs1bKxet
shz7boFFpT3s6N7dttIm/AvBMmGodb2PJAsOxsFwWflg133MSCtjOZ00tVO8LyahtK1P7XZfnb6x
5xYZGXcVFzaHkvfPK6zV5fU6qCdm9Ajdj6znaBGg8iWvHtl5sTFxCAU/u4cn1v5CgIHz/KZedprz
YwTmzwFOBgromx9mWHnajDQOd7FCdh3dmXQTfTT8TovL+MaWhC5fVIZ09sXW8Osmmy5iINzI9Pya
zj7vSoB+zGkkz6WopXry7UTtCR7q5juXt1Q9d2+VMuHWFSKBaeGUL/7RfX0Qka1X7O/Moaq2CAhC
DWj/6MA6YBguWlktK+VC6CNbpj00GEL9mTgTVkQeP7bDzYNcN75C8u8MsCvi8uUP3qDDwcg0emN7
jnI0PK3rh4W0wkDO96P0DUzXuMruKu1baBtBRmckqo+TDRH82EggLv7OJdygy2HRnNBJT33yt/17
j1KdE36wSaz/GtjnIOYxcbn2y6imSA9ZdbQW2ynuTOxI5rpLq66smYfdYfz7tQHaze93Scf894zI
hP72/zD1eJDnUBgs/P27WracPt+V8NP54YmNEBZdDUQ7piH/2mBz8uQGU/yfz5C5RvOO/KNqn0vE
1LitOEkhRshfMcvo/xZF1dE9P/cBohBLE52/etALO79u2RZ9FYgn27nLCmTqemR6JFSS3KioxDlL
BH82XE8T9iqGd6OEXGMW2I6cG3Axdl6V/fZqrSAn/14DAt2hPwLfMK5DQDYWd/xVSjvDEP+PLR4H
e2+ZYxExcz/ieMSJyxmtXao6Z5Y4xhGVDIk3wa4KKhR0DnYVFMYH13F538y+PDNem0uxxaDIWM+J
KMAAufFYCVyv6UQZUKYVES4KG/wKi9s8h6cB6kc/qlSWLjMkF/ra4/HCjgXY7qe0IKN89yRzDv7z
JbJYHRTHg15CR/1YBki/mzq/lMN+9MSr8sUq6PdyDHgABNABXutIbrf8CIx/6EoYd3y1kST86Q3f
L3XqcUwXtgMMuo4yDSCdQ2kh6rQdU1lOJp7oIgA5RuICNSdOf4r2F03sAhloJEJXotltdaO54yRh
RZY/7/NlQ/FUeeu8BjfW2h0ZanGcyXMoLN9CN9BG/sEOKUeJ8s9FBk9C6AEbHnKY4P9h1ZgLB5um
/DKTfPcY0IQu6MplJ0m0jBa2U6BbSytw+W5C37u+TDdhBUXoP2V04OGQdVXl/geX1sfNeTaQCfbN
KMb4bDY/CRL/RLOCpclj/juxsECIiV6BcFrjT1yOpo93rnMuN2IHs0v0M2Lk0jVH76EZU1bxLDK8
wTFQSr+lMNnmWi7xzismAFDVzhlTtxfx0KCGYNodauw2EnaFQG0VjC9K2dOf0tm3/raiASl60fPP
FqfvmWtpaxB+asH3Bwg8llwQ3UXtt/5f4iCYxJGTMCopw32K/qScgBOaJz3l4jSVxrsFH5geHFzI
9TOCjbh5sBM+/epMRClB25BWvSWJz1UL6/12ZFJGmQDdqWkHUF0PuFdA/XEg42fQJlk/5v5Dwyix
2aoqmG9j9ImxGMouWl7HOU5gVCt5O9YNUCuQWRIF+9KJSPmvrjV20tGSPPsLCSQgBrKaqenfJZmd
yj6akBN2LbgwWxkrySpC2xQnz8raLuYuGxJeolhNYLOVlY2BtjvvGin7yBgXpgkBr9FR78VOT9PC
05T1k8njqf4I3vmKH/CrpDW8YevYx7QGQTv5Bh8Qcx34pf1DfL3Dg5qouv0IC+Smo1MpqwL5KYQc
zYCHPWsPd/bWteBlmm0bgDNBbfFuRuqfs+aWYNH8t9Y2Qb3sSBmM9hrsmqiKgIEWMYHkY0ji6bDB
QuPqOiTP5Z+Mgm3Rc3tA07M0g/k6RVx1lBOOSajj0jQ3RlxMft580WFYlWowyCLLm/Kd/Oje3zgO
b83dgXXi3VUBOHTZEVOsJ1s4cUUmAHdbWz4JU3KY4KeTdv1qV3JUqODJd1E2F7Qm/JwmDDIDEaC4
W3us1jITfzq/ClWWtxzJ12XVtJLFEjWQmtiOk4PYVUoNMivA+ni4CxCFxVUt5JbKOgHsq7SmjzPo
0tk18t2OGU6Ko9S+yg4ckpy2sP7qgsFwXAwDJ/aIIpraxxnMcTmqmWX9N535imfOpSXImKV3eYsJ
Fpmbsmnbj/PQkggzChNh2rMx4YoCnSJlmHkTfTGE/V+//165aOBacwDgqznVueFlvheOdPjuC4/a
DRqORrtBjmsooovaP3FvWH6Qi8Ocj9WYblzCIdS0eEqcmQ3GoeAgN2ulp+YNHVCxQIRwsbFG2UXg
H1q505Tjl1zGiVSlfNuIJfjObE72yiRut+gyD9UkkahodqAKc4a0vhucrg0QDz6irRjWpl2/RX9J
v2xiquPn7Zrb2oxzf3XQNRuOgNA4trqGCr9WfJhVgjPlupR+Ux0kRyKTYvWWuY+NZan4f1FL9ixX
pLaDbdJTINYwD7FkdWKlem+VySBSOkhFI/ZybZ5sWjO+Pr96ND77n1KdA5qqxOFkaLi81zy4WYdh
P6Dn9E+DxxQVS4mRv5eqADUNtofQhfatd1ciookwVRKjogqOfapIHqXjs7sM1QtP/8ceH8NFpw45
FwhKmpLtjjwNoF8KYPomIWhVf21kr0lO2zdvWK8xLhhEI6/IplKB7KCMCSKE2c+6v9/0oyeB6ult
1YkEng54NOal3KhvNZUWlwnNJXW7z6NthaWi1vc8pyq9TYfz1o0o7EUq+1gkAmno9IWHV7uHbc0S
NIfmtGKsviuSjnWZe+AjUeFJ6U+yr1mtDwTwqUL+Hu4kwY2j1gW6BrNK49Va4Y6/hwitr+pqy52G
igyMFYdx0vgwRntppiHfR+I+MZE1sMQ+Sd0WImrv+dPk4vD+OyFOlJpf+OEwLCQN0ZMS2W0NHNi/
hZ+f5MG0RVknh2JFxQD6yKGMimYCQGacRAlyYf4B8jqLNiofL1BESRH8N7VBz8TbuY0Wrmec5Ut8
MhyrX2LiGdFENcAjvheezINGZk9HHRhLvKPOv74+46fiOmbrCncBofZ5qvcT045w7gE2ZDwAlKUy
V5fX+KkMbCQHwaiG6iKnkTGHgE8+aKTkcKmE0COtWnqp8TG5aviTS1QAoJdMGGVyxqyx0zyeH/oo
Tph8PaQMMOmlaZAYML6pj7h6VgLrtwTpWwvOV63fOYimjVk/qfSncA7i0EpIKuQ6pPVNwTBfcyTj
MwMYrGHryi6kgAvqTKBjNztqOCKCWXlLH9qK5CATTUy138k74YDRkQ1A45Lp/FylV+0OzAdi6XT9
G0SntyfZ7RBBxf3QBQy5fHu3reGhL9v7HJ62WLdHjcVGBy3naTM0urLdEzFFFaqYFJdwK8r1qBko
jwNAbZbWqHbWMSxOUWlfuTqcwije7BVYzVK3Qb1PM+4If4hEq4Ccv/sLKxHEI6A8oA/1fny6SJKQ
opglUlju9RAu
`protect end_protected
