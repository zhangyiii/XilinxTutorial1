`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99584)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aPkk/LZprZljgyNzZTGF6gcxBz
LkEl/7f+3dcASD/i/Kjmzo5UztG//wPk24MByriex+1sPqTxcXlWV8LDfVfdewNsQK18ri0zF8H6
IAIuaAhwldJX9KWmFuUS5oBGXGuPxMTq1OrP0homhRyx12SrAkGr9UXRE76SnFbvQFNNwXh7AZRr
hC0XmEcK97R1z61C09Is8ldI+YBTmSydRU5VSSucQVGGsZ2LmnN9ZI88dPHwHZ30mLeTMKO8WJIR
dd4ix72h5w1X00yS+Xyu3zw3LyGgeqyncIW5d5c6T+UbuE781rN6t9QDUcfPMuvjeYCR4ZD0XD9z
hQvD2URjF/u4UQsWz5bvOxG3UTh8Q1UXXDsm3Z7v7T0amkML93mof0FPV3Npk3Jgf60vYuMHMlAp
ogZ4hITwoS76W8NgxmA72vA3g2pIQyNHhPAb9PMx1026NWGFqnmDcgnFxfdvFd0SBIljyth9qa+O
BlZeR48qsqp8NJm0kBxaTfqCU14hA2xKy3Zj4LyW+ioHWkjA8FVFM5VJniZsgsIfIQKfpOa8dLBk
P6BuwKFJ0KWgpzTe8MDDetozgYuNtycpgSecZzdCTE9BWLa0jAoX+NLWhasTPW78wntvI+WsbEE7
3NG+5wB3gCDPtVuT2A0pGHYQkCTNNVn7atrBG03PWFtYlUgkJZXy52CyI1M1ze6UB78pEJOqjlvK
+j5GvBVa+MMQEisvzeYv2xvOzDWbaSnEBrFSqXGpz9esBkF1lAjD8PslXPetsbwtbgvftSLbvil9
S4NHinkUl4U76mQvLaUlbAhrwGcOJPwhy7KmGNsAjqRIqLWmb69eIZ6H4XL7SvffLFBAWT0nM2la
DFX996CNjqqvOua0LBoei0YE9M2h7Wi5a+wlj3uVGh3C4TUPASx9C3xaVT963xIzJJTpKXpsqoiU
HgeBaWs/Wo3VaiIviYPfXJrC6rNKamKpKwD2rL6WvHVWsX3zIQ5GzdZmClFa4+rGt8MAwLBftHsq
aN6szKciJPJHuQOWxnEGZo6NR/f8Pn0hHyCOFTETP6wXCp083PS1Cytj+uqTWgEJiJNvq/q3K0Mv
ha17CT7wcoekDHrJPOgDFnyuI6j5EuAAv0itSQTmh1IG75ZJPoYQjeJvvIlHBx0tcSOFmZtVWsKW
OOIF5Lpef9BUgw3qbmwUhDKNz89/RzMGcuiG0S0JpZvCakGoyHOqfXhhxji0ojmG9vIxyFg/Xh3+
7oXhnHxPbJqZpKdzEw3b7G6gz63nHdeVCG4vEYqUoB8BrhckObSK0uku65ealbhwIJIk2UFLtuda
0zmkR/3Xn6JX0Yj4elFrmYC49DA5q8PFf90pA7QsxeO5rgGSpdtIFP/1wPq6d/mkmnIqn0pu5W1k
+VLSh7gjC9yroB/GPmmfCLvzqqpdPQzj9bxjC86zRq66UiXrQrFRvXzFPshqz4id7Hiv9zIODerG
lHKnpvAKrBxW5HwXDNkKmj9dHZMK6uoVCxayFqZZyr3Tfw/maTgi5oHQK0znEMrVE7DmaFgluwMl
P5m14tvDmJ4AIYLuzgFLQs25kGd1YZ/ZvWXGpovuriUP7hI/jqTQEmpCzSME9iNfElmqz734sErV
QZZeFI+GU74JvCsPrQN/nEvzX7WBzf7KT5eEi0FXXkgL1bU+Ki6U5uI+GWllpJIz7K+VRJ/eZgx8
W0ZKh9GV7E2+FOLReLBrR0reW0w1lC1Z+GJiParHJCc8FHG8U1kG+eMcp1Qoej/oeHUIA+7SvcsP
pBVbOt7WYJrj03H/0cxeMQG7uvCSGnZtdEk77FQqy5g9WFQYlxCGokyN8ptNcqUC9QudyTUinzXy
J85TV/oTKaLQHvDIKfh0esxFzZTP5w97El8MwAsNpENjDa6yV5xwtgQIiXKp7zD//zNA7X6IFDwQ
/EfKjcHqqUMCdhWdhTfAjV+E+LoJuTxCr2+TcxTChcfn0sS3KMUP5kohLUev/3S0VI6PYHgbltsn
P2uB6zkNgWTwxAdMVvcjEZI9/8j0AxOnITICXqhpOYFBqA1OJou4AShVOXyPVFpCmRz3mx7bJ+LG
L4zVXbfmwH+Jop/y4AgsVEQbgEu8iDIRtT3Po6MDmtlEE8gB8IytXxPIGjAldStUru9im3lCOLuQ
2IpMTkhDoVWLvj7WfrAS+QslGYPfNZD8p3lFidmq+SX9+8j+GupzE7iUUk3qb7vGYYLqz6nCPSNq
epffRtBvd/zoJBauyMJNFDWQ7oeS9rgKxKIcfHD115JLWq98bhTfPr1UETvRQYwlR60C2aw3k6iJ
PKSr5PY6fVtc7jhb6e5zjzBpcLzZawJDYifsv4hVIye+VbA4rDD5D4YsLvOJRuTlRw+IRK+S1DOl
WhfO8inIvGBth3Deul01wKMkvs76sGZGKGSdICE4Kzdi2JjICk1snUhkmwdjoAgk4M10D/zU8b10
RP0jLJxdJAHXgdwaY02Ap9i7xJHvHTifYy544wOSstobrFzu1stMYv7G7IX83vTcd0pxAehcMycF
CNs1prrtfPJODrL1q8jnMuQ47jgghjc09crwEi2alurqJZE169+g8xvLJa7jJt1GcG6seFbstoUJ
q7a2oblKJrkmEGxw3ihR2Cbj+1izBulLliPe3/C8q7kk08olQGWcTt8eyGB2Vj9OYQ/9KUnuAiyQ
fevsYDEd93F/g2yF3Wwth+kieIH66sBEw5TB0QXtRtSGO1n7rvsC5vzPqB4SwO8jL0dsn0rgzRKx
g2eV6I86jwWcPuAsv2H/SYqUem1gKOJ5m92GYfglP4Y/Murl0syDOQaC1RwE0t6CpPEXDLLh2nkJ
vzSfdEPEBnyFvByHiMywCHdJ8+4eVXFyiECa374lVCDT3YMpzBwd7ywtK4OITS3+jBQew35cPGjU
OHftczgzrq5O00Y6DO8UDuXmWWmFs+wD/V/sizHwMSRKFuxOOBq1Zedo4XSJfUjMoD2y/p7/V2DT
KLw543nS9arbgNAFkKdbgwuIKQCNyotcMCz/7FTGs5/3OXqNbXKWa1QZnB4rQPyAVAUc3UKNsIkj
ofUWD/UL19/62x619GHdOdk/4IBZQWClszGJUy0Hs3H6MOxSjd0f7SeohsV8h+/opTwwDZjTioxJ
LRLnf7PW3M9m22iNVYFkpx3WkyJYtHt8LSYIvvkP75gYTbFNXeoZD9LfpXds/02EoGAa3eDd21DD
doM06GvCpoT8NkbXqMaO+CIa9BBufHNYpoU3KKpa7vAqxQ4K76EdCvRaQcjzCHGafZGOpMNk7uiJ
MHccL1gfLEwKGWxLLZpnJ1MDtbmYrovKL39dKKfTQKBDq2USc+55xVb3GYWapb0buGvmiD2Ll2z/
BO/y2/MiZzNaXv1jCdIlCRcLlNDrBuXsjvAz6SDnkUN7+U3lPO4HpETjIvU1SBWYtrQwgGbBiQmU
oCk0tFGum+ZX6FWPQ3Qy1fR/LAdV30U6nNCzdtREc5y77rmbw90PhITzKGUgFf9pAkVrGd/97DRS
/BN9/YE3LGBRZTlVRoD806wKBowl6oGA2SqAJQUB6MPOAOL3D/yP/cYoCCMG2P4GOoDETOEE71UB
eRXUXVolk/KYhohXruO2nIKhf1gEcEnhpfbeN5+SO5acZaXqBb2GqyOvUq9EaqlwCLiI/yjKOKIb
tLG1/PbXQuM9EoPqPxpy/W/WFj5gpARPo9uMOp2nPQ1eoBywaapvmeO+anMT2bamchZUDlLde1cv
CgUp4aN5BktaXda1KiYzrVuN/fH0sb0tRnZF1egBMdrjHIojKrnXjcEgxxiv4fPrGM9qYEvl7DEg
o4kCoG4a3Aieqhl9n9fipUR4Tknd2NFmqOTsHwhPFdK7QPq7Xi5U6a+aGlu1ffxfBb7oZXnbNGKZ
pYXqAaMUjzcG8ldNFqN/r9AtMs+/eL8YFag/dcuK5POec4BZg0CAF1Sv207ywAFZC+t4tDrOK3Me
oC/Qc/YYJpw5cj1jJuj1KH6Qz73ZXpza9w8DDR+Wx6U4f79Ysx0fZlJ7EpjHEtnrwSzVMlKO/dyn
wUUGp3LYwHcElFkI7r5riNDkTKYDpBQ/qSZrUwvAUcl4iNXiEORYTyOvXP3VoWVm0Nd6acc/UPgZ
Al23ZOzbOq+a83OymuxKj3468u8FjR0gei2QmSAOeuz2egkukENrUCAlGybzYk0Y6IBC93GFaq2C
rQ+poMPNN+PJTCjLyGA1zEo7GAdQViUXJOlG0NkVqDA0bHKyujhWWz879yy5pplHBjtP4Oh38Bvu
YQlbtusSydqft1cJg9oSduuRDByvJcqtZKcoIk3KiC6UqlI+U1FA2i0th/lO9nLHdbHQhwjM5PHc
pU9KebGf06V9SXHPYmyLTR6OOLzgpGOdYdmIqlHP29OMS0axVmBFprNWjDtq2v84fM23dMssG00O
chyyMFx3zODv+QTHXtXH1sVyD7LuVCfg5PPWVQE78fkfJlb33LSVCK6AA9t987ABL1g8kVFzYajS
6IE6qEzATQOZ3ngLhv50ivOwJhOvWUMxLu33vu7Bw5/SHslYi6lS5PVcRWiwUiq+PCVQbdR5DZfx
0A490ixAZ2qRSD/XAgk8j/ESbjr9etjVASlhC5rqsLR7NcbOOy2GJhxXdC5uBFb8YBn7RgiYC5kz
Nc0zwYTkIb/jPLboE/OtxUp4Pp02ai/KM9FIw1ffHA25NqVqIVbG94ZBcdhhRCrVJxKGakGZ5iGA
eRWM9MqlJsiVX0n02WAjH2AodzrIDXtw3YAh2LpQlope4vOLgEpcMmk5afOnInYJT5yx7u3el22X
p01/WkjGkCerWcBqutaWsPGfjYXwsYe49UDrkEi1sReIp/fzUSul0haKfet8lJywWqTQOUJYg307
xocJCBNwKyW4BZMvML4Fvb9aCFbMkE2b74JisDvdzH305tU61kfr6JawnAVysqh5p/zlR+hanxSM
VGWRD+bZhK0MH5VPeENBviMspru1ZcfMqNZg4331mmEsG8sVjk0g47neLOth6sP6NneisfXejaaR
bE9L7zfpcaXOSiFZA7afkPGF7BwwODKEhG2cxbVgv0YjgKUD0eUaEfTlo9m35BPfzW7DLBkiIYGl
OueXS9Z0AJemUH8iXD3ZXqkKrm+p0P9JtWa6xA5Vzoy9F35gJZ5DBdFHJuSvGT3gug2+u9nqPXdk
OKvr6msi92wDvYwqMOBicY+xgwFQud13G3Qj/G9RPvr5HGXDKcaVNfxcljAPEaIvf9JlRNxPs4TB
OAcRiy10vJN9BpbNnbKJOAhSiK6rTUvZ90MEE1tCvDZKWUG97J1x5CPKZCfcf0Re41fWF8U0VMJk
lbvEpwouWMqYvQ6SyQP1IcssMOfw9zwz9KhOWbaotXknbtGmWScsoOnQRd2UqkP7x66D/2jbfIwD
5++GYPdQTxGLrsMs2d8sIsWtrjWgE/+4PtUaM6U0JWiNlY70YudU1CUHWFCWPeZ+x0zlJWTYekYt
RKBVcyWh9VXOyoI8ao3RlYdoWKbOl/gcQVvF+tmEbHhN0bGQSvaEicAN/UVv4dZ/swVcIYrM27Db
sdsCZPLPboRlZNJFcVdx3IKIaDCo+Cy5xTEIPx3XuN9NazNDvD/uTSYqvlx6TlOauAv5Em1wcdci
l1pyTTFsGqYbmURXFub1D2D+bZeRIVTB/Aeo7E8g5j4aqKtKdMNR4YlfX0edJmcXRDcjqXVx3Vf7
Ud4L+hngiNe9byMk7eyznvwfF7OQaFcnQn+ICK6SMdYfC+Tf1RVrhjF3bmz/IZwZ6mnYW+KjbG+u
+hEueKn5L2KZdgDDLYFTZbNsneUS53q5938XM9xorFI/cfUBrntSRIK2JO3NQlo3q/eO+ph6dJBo
exDaAPQmMthaY6MHKvhE/H9CdnW2OqyT/sHfrCEby24UD1tF3+O/xnrucpOxI8UST4Xe6uJ4Ggod
ov1iaNzDIDMPFSKPM6ipSLmAYNKH58jgejp52LMBbF3p6ceRcr7HI29cdQClv91Cb+Y4KTA1tsPD
j3bTIMepkjneJvp8jxQKzFINhHmUYoXvdoRGi1/b1IPnrBJNuqYv920WFNeZl2EAxhTq4F/VrO9s
TYd7776MHz/FOqXA8OSUtBsUgJDxvIVGQAsmCN5ye3GxjCV6slJeoDqVlqchlhz5Bgd+i+7egm3u
rkzjN00vPObey7MDCBZH0J4SKO7kV2ohRXFBiDk1wbEOtaaTIrAQxefqR9XfhP9kJdwds2GhvMCx
d0LWn9VHAEG1vMvTsHrPH3BylvXBLAiTTS84qiMJrCzczGhGSMZiY/SV49iV2wGJN5JA3ZTs4L1T
RX1sMrJw3hPXP7h4mSOMy+7Ky2o6P0EuxzLqIGYBpCSuampms76SyVT16jv+rLcnTI1BtgWnVLiK
5zPUL0SObNGXFWDBkRcry8KhYcw6QwZQQXWK/9GdLy7sWU/E+hMPjH0hQ//MzoygMCaqg6JeBJ4P
vE7gIp8u5WZG1CjtUqwlPItH53VS/AA5jcRylxxgtyuOaS6MNsD8odg0EY+SGVEzBJgiFOb/MtNU
epQhxAAwSykq77fFhI8oOOYWhfOi72WsxtIwoemh3aoXiESpRUrtk9hrlG607Uk2E2nOtbG2OuPc
lF5T39nGOhjBmE7YzoZezimktPgkTxwXrOvIgSof1J59bKS7WVq4Ra0QGAqR8G6xnjy+HVCTkB1T
s08JCJz6ZioquKY4YAVnVNd4qLNQUMipanuD6AEXcbn+diA7e3oK/SKKhsXCqed8Qq+DkcwZwqPc
SwgDk8QLzoWrSXYLlMS5rvJggtEreumTT3ap9EIpH2jb2s56vWW2sL8UyR67nyBkLV+dmKnoyT/p
7upaROy0AflpMYJq/CtyobZSHJn28RG+bms7oXao8cLj5sVKJwxsj9AHUXriZBUlAYMXjuZyaCjc
MGzNrT0cVBZcR7Ww3x+p07im+VEhf6a0qBMoYy6rBiFFlmApIhm6Ls/qaaOGOx0WLemWTjtCLK8W
Ll/ONDF+FXadZ6fnnCXY00TpDWewCsTxim+MGckoft+xGw5n2vhFdQTyuBcQfn7PdSTmgbkpBVWH
vPwsu/YsqEp/nC/uCF7WqxfPZaJzbxsUazHSk6amCAB/k0yIe2UkuDNYjf5+xlxnW56kjWwQoPE+
cIMikJd+Y5GWkvJ6lM7JqXFmSP7QAFZODipuY9D11stZQrz1GgP/7oTU/UPm/1ztcYUD2vfHCsog
oGh9K8cD0ewftyY5b5TAXqD9CUpcZ1DTTz/IvKL/XTOSVtCU8ucLe1hBc42iEFuCUPu84hSdTpkg
ZEgBD4X47aPnYe/GqXJ/KIKvVCJaNueo3HcpZMinewYayoeaO4ZGaPWcoUgs8t61k62KDF14wNDS
BTQelTIKd0gCHOcN/dTSkQmrdFScRdyl/2bNKJC5Aq4lvb7VwIjzQgSZGF2samaOANOSSo1TGV52
komBx/7/1UGlfNwTUJIk76AD5sjACfMPvBPMdKXBYwUqpx+YP0QwAP442XOYNPRUlr2WXHDwaJ1Z
k5uZCzfFaXK4AgLdKmjtsXzvmtSYDeFiBEXh/yG3GOpCxW+2TekqvzUNX7dR23mYqG6CO3HclHJ1
a4sXmEcEtQRPoD2t94Grhe0VLwnCjEwL9N7+tqn8RpledzvtUnU2PZBQTmYjmFt2FrrO8BK90VeM
6oXeuHPM5Jcu1XLm6r+pdNRgXbealo7pduNlINqPAYdgGLLsn1KsUUHP5JLDORZhhBgqX1n+Ibjt
Jf+8APfCBLhxUms7cpl2iRC6Y+RAIaJmphAWQLijZ0NJcfT/2DGH4kIOe/3jAx8cgz+sxwzkN+Gx
6HZcADOCPPXkobiN2+aXgajmQQgqNUkhyb1V+VNb32PjOk/N5rbqdzsv52GmkzGJUtVthHUH9q1X
fh08rCZ4CjoJg/d5uDM38eU964IpuzCrmp7uCM68pY+eFn1DiebOsdez7z1GZT+w2LnfNkPoUyno
MkMYc7FT7oGWrlqxMEmH8kar+KmkYswLWlb4vdYrWoNu6CFQmpG4VdFpH5K4wF+MvS8tWqRCOts8
lz0Bk+U+UpDHsdL10n0cA/zfPwTOeXMPp2ORacIKB7JQ/vl0Ork4AQJCxuRnQwbzpivx1/NhMwnd
s7w1RFxOelApnOW/JPJekuT1tC5d64pPfKkZjN4TKhhP3/js0VgmmEPQL11/U7UTVQnO0LxrpRiD
VW8hnKSZspidi7zQoiJLIOOzpx4TuE/SxtLzVd/0qMrtWkW0O4PqzqBoBNdO+6oL7hxRZS1byRdl
i7BN1sPg3Khrc/K9OltRbGW5a40xWIAw9pbgfe7VEdIEP9hQSi3PM4LLh/aF4RPcCTJ2dtdhG41g
Al0hbuCJ2EYoxfWuVpuQO08Sirhc1nGnFdoeP+BSl5y9flHUMfChbXuu+PCTb6FrWsHH9hpLu/8t
gud06/f+kniZDN4YQPan8KQi331XUXxXtHSVC/XCito0+qCwU924F689khKfBokXE6y30NTxyOaL
89pHMXJIDDmR9nhDPPzlhuenm29i/Em4RbMrKAeZUvHt1aWT3pw0Dy8KaqI6fZD7d+BxGrHSa0ra
WjeVSHJT0VZbdDT3rXPnWWpxV2rH1zdBU/BUGbKjknbUi0dOvJ2tG1dUl2D8SIHrGY3FIQrB30tb
reSAmVyPLMXoINwzqwYEvzkgU9uKLH/2AuQZOY9cdMXw2TQXEC1UVyFQN++l6izgnyzbw9vv1DgX
jiaIL1EbO0YJvypwXRP+xYO4Ty4L/jnXdAwgJXjSRdXz3/uyqZ3nwpvWMcX9Ig//N/oLgVyhWJ76
9KPzEYEcVxljTnb6ns1Ckjx77ASl28xLqpV14EL2Hzf/25CTXRYq/leNtrTEZrwQjxYuJuAnrbob
1cUFWT2ZPKiVSOqTCH8JXHMj2Spc6+SkgINI3kTLr7YhTMyKUQmyRRF2vaBl/p5wn5KGbEJyZcOx
qdHXrrGPGEwEMz+kLgMtczJ0HthtKk4AWjHBvhcMEQsiaI8HYOmG0RFIumWpx4vOXHCK17V023P8
+GQpe7EE/a+1iOPMlOrIoLugZPkmjZTd/Oggzl8ywzWW9FAEhzf78NcCka/4xxA+MKP22bmKcq6C
mFPPzR3TlE/H//0HBFsjV+PoOVXudHQyS9tJbonbQaxunUAE6MRimiLyMBsOllMtY4Dpe2Y81K67
eW1s2KGbmYzgMdQA4slS1CyJzOj9zB/UlK2kUFvBc9x/GPxoZ/490sFrLcPvSas9dfo68LHi/yzG
VzipvlgEHvj6SzkpzzBggIYsAQ+0i4U+Zn5gvMjOsvd6fXK+zP+Q4faUxXrDlckIAnQMuUi1VFYh
QWsxv2brf/ARM6THK1NX3F86u9VirUkiWhhohEef1lzYXcZlCgOQWYrqfuUr0uBkee+/YpHgyWRD
NmZLv2YXZ8Hz8v9RVDu29aLvb8zE0aTg0vi9oovjvnHDfhmgiY5KFgfieu5YgsyO/ZJgGwwBs4LA
aNMgXZL7zwgF1CzsJGJ7Wv1g8mnWRY6u3yDwFQTBPOMEXfYuStdF6xd3cIggdEuHHh5uFUJOLYRF
9Jl/DrDQyMHZxlcGoZUGqw8SvfyzKZ7vJtarfgXLM6TAt8wIQxkw0Nbq1x1X6ZVuMntcm/Rkm+yJ
olAH+ohgmnWhsTem1NGSyFu5Du1Id8qdlSCspt0qQzV0qZqye1s+znbMj9X+PeEMWFFi+gAV6j0x
E10ckfXJiG7viB6gZUc/nkXDUj5dzXsOpwtxiXV+hO6zxJA2rbVCyptmva0Gq8MfV9vmu/zOw7mZ
uC7H0ATplzgSypTKfJV+GZQTBnGIIvpF6xWq9gDz7/Mo//JHpzBcsMstrUQ2fN81s22RmJRDNMjE
Yn1qJYpb45MSszJVN7rnNRpqtw0OkVWnxZhVUEvppmphK+JT2e3AxmG3eNO7EYsLckU9auSA9E9W
bi+p7dnnGLTGdczjpEdz6/e8Ye6p2MdrKVglU1TQ7G66D0/ka2Q1U0BtK94GtQ/oC/qD9njBzi41
jgiMUegqMYnPYFx60Y0wlK6+ajsu7asbwhGZqfPbx62s+urx/CowFvCp4khdtjYApAyiIobl4bSV
WOIi2HoaVEZjyLdDQH5Who3sHMorP+zV7BurkQFQqMFdb6dhYx3wGzRFcSE/uaF9zN8Dmfb5yQKW
jFIaP+eTz/h4UG7aGfpXjgyioQlDnZMU9kAM7SrPQm6cQ+Aou2Qudo7gkg0eBpiu3jQYzD0CH/l0
MXGckn+IezCzU+6v4suUeJEd05GvoEbhtYKDWDhgBwfQhwu1Hyk3h8ToQscUmFL2PbEc9MqzPAky
hxr8Vp4+VLhuBDiB8kJoQHdJyhMUSpVa3OR0WjI8EIBeVuqxrTcGkQTxu3ALTPdV2XBbhXZ3xOD/
0V0dhQ6vz5fZrXiQDKnSnC/6UnoLXPbZOrCZJqri623DysxFyKQZggY7OO+ZeKXzN3evYQwRRTRJ
Kik+Ae15mhTo8lgu3KAF7yJq3puWPTrOR3IYLryM91gXsyX+/ji5jUkzZB6PddFkEWJTGab2J4eL
UwIkdkjHm201e8Anexh2+ln7UOD3WyxyyWgilNn8lpXhxgTE02YywnLBzd2UDDC4jlYJsKbV4Zx+
Qmou3FO4VuMnV5h6qAZxDZf0RR4X2jQ2sc82kpfTvOR8tE7/8ZD2Ru5C83GkUww6xG7aUVt5A71r
0HuFCRFzkuD8z+Hmn8WIWC5MYF0l+q90lBc5o5FKrq7unP8PEPLv2dsKvnZSkCuLG9GzyaTahugC
xZxOvo58eo4fHFtI6gK6Tn6pXIakv5bFcZJTKEeGzqWa/Jmge4Q/R7xTnWBFs50HdaulqdP7jlhp
4Ber25hwsodbnpLtHHHPgsTBzTeAKnFVIgqd3VLmNL4pZpR2FvJc0p+DuWYWcBM9csaqXlfCvYLa
vcdBYaYtAAYsMiB3WqyAw93wyvT5GM+uI5zyxt2vzUxitGeb/xGl4jxfaQwIXp2IhBB+UyOC7JTT
3RUUWemQe/HMzAskVqVwjNTaGvMnbcObER1ZbT2dwlbD54/MLmrELguy2fTXyNYH55cZ0NM9JLbj
iaF3b7Pm5udcgaAxjGYdQquwjKzGPiXXmRNel6XS1sFUxRK1yF7cEwzTaoyxZI2jkOaj7bEMbyLE
h7yGU2GmytJrmO+ijMaI0hD2MWNfFJpZoVboeHegS4rYKaj4Pm44G0fb9YpkTpOWAK2uThzLVhMA
/yAqAjMAb2imwoEseU7ycNNvaalG3bhKxgb5nr28sDB/qtOJKsYFyDS+Rh0QmeN6DhGPdTcOPOx+
WFsS6qoxJR1T3ijz9Ytg0iboC5G5LCZOgPIW5uCiuGu4/gU4lx64o3hLWhQq9f3x09Lr0odwBNBS
bJ7kRLgTe8E0tcWcRL+6JP4371IcEEDcLo2ujUBMP/Qz8aGqqTIPogaMypbn1RzqARdx2gpPJkZb
7/d9DfR5yXdSVoiTNJUdZRcCjKlsDYkXB/i/J7sq68w0FjnUghp7WPqugZV4k0E8gyHK6mdBOWal
DDLVAvMVs7BrKAH5fyeBc9xXAIcLpW+KV6Bp1MZUQyIwnm12nsqEZoibrSET2C8/MUMAxfsAtmP1
GgDtcK48bfPdVTLOzEXCXMKxEk9Jpv4vmvYvPIcQ7r/OCc4MIZmzAsn2XVgHcodimenvuroH4GFo
6rTxuJ98qzBlqqOrmYYGSSX1MSg4cEnhL7O6+J9KVgNb44qKZRVTsoPnOhmCICVk0A6j/twqTXOu
6oAHKJn/41ceLDBGMZjgoFtXjis1Dsvs939lL4/Av7ioQ/H8sMSyRbcfkiAxAj2JPcyji6okhnzW
Fc1nhJCDZYsCCS2Z+Uf54tKSxRh4vmLCMWHIBEFxd64qO93UdMSmWFnut7qFBZGnJB/zyxJoyKzD
WC84XgeIyR8LKCPM46Acb1DhHL214cIyb0GD+IbYya5nkShKOcESR20vVMERmpAEPxmGPRmweTYU
S711e43G2uAcz+u9gNM3WsDBJnxar4RTj1JGegB1qcJbr6hYzWxpzr2sLdcrYY7UemW8hBVxeqtT
ajMZRKvXhozPqBSpI89QODHmnvGzHwd8QfN2jyfulv6zvhV4ISfe0hRoqkyhmgcxCA1tIOy6DTxN
jz2sYRymLa+vnFGBZhSPKcXHQEqbBFsNyOeZewj43Hac29A8EryG6F+qki6GgsvjdDYUZ4zqC5ZQ
J38TXXAhUdPvgBddXQsl2T34ayCbZ+x3C8GeprXNw2k0V8UbGkkrzqsQln1SEfd22rCANtY+D22n
Ri6yGPh3sX8BH+FvoLj7hVTiAOtZCvzkJi2FWJ27Crt58o1W6JuuSslIKBpR4KEaqjrQ7nBcRALn
aqYzRsMLsMLSzDCo89p8dbEXkALrmWVncwfd9LISUMS1VQmDb7XYEz9U7DMwWfqQIZPrAmDzTsNb
HgM/gsl31BZTZbFQvsDckVW2+tyx+zaE4nIwOFSZ8U54OAyvyJlz7Dde7gnGA0s3lHNAWfZKfjSH
A4iCtFFzvxujQwtyQnAOPE/4VIa02LNTln9oBpLGl4ECrO7+EsuJkvuhW3D+fEgZ28A4gG3ku9/2
RZRdpwkTGSprsJL8mDjniRML82Fk573Q8uYR9QCMdoP0zJEVSTh0pnXgTkGbydYSr3ODbs0LALe3
aBcgwWnyt+cj3NFFxxchmneGB66YpA8orHcs46NKnwoYPF1EXhchakpHPIgswX4uVDHX5Otowi8Q
rNEsbpfUd377QAM+nx3eouTiSGHQ7xC67ETgwgwY95/ulQ4vJgw9YOVJyAGxDmgsM62yrmqOecqI
DpPxnBems1OEpB6ueNplMHsGgXFFEEL7Innnje/qA5X77Cl21Z0DszAZcyAYKnNgM9ApIsc12QYg
7GTtm4pxn+08K6vUHUoN+s81P7aKOxbundhjQOS/JCEfSEl2sP2VfYaQY5zB9k4Xw2O4SJPvc7mp
E1mZRZj54crpnWjxdc2viFP1E36tqPwtGI9fLrpVoZmOwq2VeJ5JHQ3Iz+vQMPz5j157hGSzixho
GU3oe9XZEZiqBgquLc1apwDn0Kd3X7vH6e1d2IGCqNJAgxhPkiNgz1H8SMecjmfPDhNJgo+L/r8U
Hu2JKH7Enke861t3UnprB2rDJuswzo+ly/uf4zEX+nH7mq/UiRwGOqxtmdSPb9wJFKS4EnqPaRty
Ue37si9ViAyw5HQye4F+ZwAdb/9Rn6solxh5jdyXuRLeSo/wxbj/OJcAIfKj3Sjc+upJZEFzFt6g
gB8TN6PPuDUfDRMR4GAqkQ+y+EMLoHPE5AvUTG+alyeYYBvDjK+LtFfh/O6Joo4CM7nqodio4A1H
6SOxltCa4QaT4x4ecorRNfwi+BUC9GXOGhafUI+13HbkaQdQ/+OjjUwkATUqZaMEHmgxyy5fwNfH
3M5HpU6ufyPwkR3QCw9c/Gl+Ytu36hQ3i6RiamBwRWJFO91LUFCzHIBzLRb4uVYsE35HDovbaxQT
57mocVwHlJByFXArph2OdHIDpASo4mZ5pOOPMiKVzqOcISLxYGv1/ryyYgo6oMgEM2bb3aS9CAf1
0+2vfJqeU4G12RUcSdp/PiisBER/5O0z9gb7X1fzJHZ+v1JqIdvBheo1VB1kmbQ1gCJhhDy86a3S
Vr2P+4tC8/qLRAhYNGgySVD69+n4KX3WobnK/RTlgtbOEQzzUkvj6ZsgxnJ7poVJUuBY/E01ga7e
hlq/M4PQBvEq+MkgrNZt/0vo9PYBPQGRMe2TMlLDgVoJcYHLPPoeyRLQjmmSg5DFmdMOhe59Rv4E
zL75FNDW7Xbwn+oIdQMRu6/CL2vcQTVApiuqK6saSsp3SA+7OhUmbyDkesoCe9bLmK8yimIYnvLW
SozRAGWjn/wsNeWcT4Z+Z3zQI3ArT6RIYdI5XJ+Oi2KOp1UTepPYXFciVBRbJNbeQ85SlCkr7LWV
OSWsgS9xBYHRWEs6OQL4Pl997N8MJzYr0t/m5D7tEf0onZLmuf8PpeFtOll5hJQfm/pKfFY/tl/Q
g3+gXYpMPIt3uNxgsq3onwgly1NTVbHIBTWhSfit44g9GpFYqKI8B+VobV0eiK+/ltxjb+ll8Ori
QOpunEdy4dnPX2Z/qofd5wrGAGRHVmn5gIlDJ6OkqsVi6Z0lXiQXuCIk5rSi9Z6u0c7+EB0kgeQ1
Be9d7B7I/cN3LmNSC04Gv+/RpMcQQlaCIjOqThcL0GASK8yDUY4a0S2khyBITB64LLa/dYKc3tDU
DiYokR76CHsxkjsajGZ9OvuBbiiJ+RLq8D5irUURx2VOHqbEIa2Vt2VK2UzO4VSnEZY7JXzaJvbG
etv2+/RWGzppc31bJy2k8RXIJx6nm6M+S/Xps0oN1Zt0EGx8l+ItCT7AHw84OxgA752/1dp2lDh4
OaDFlwrPxUIDltSq+VXA6VEcZ5LdFyqgDfeyQsqVP5HPkio1t3gf1sHwsObZmtGiKgn6qmxOKSMh
CDFslk815f5r/s1PzKhv9NDciVx+KbujY8A6EdoBVCw0pfEoWNHq/kSTARkVfra9Pjh3YhPzOUQw
kK+KHeIFWPHR7CT4JGaJTcRogJtR5eD+DDIaMRqh+k8nUnqD/J3OOQbU8T0t2r0fZsjCv+sXA6O/
XVOnqVqJdteWpcXyq2Ddjz5xz3HDBw+tirNvforSINLYPhxtIggklAM64C4a5wHRC8yo01FVOt3l
AeLj4zkUBb0n2ZyRGne53Ks3xTEaQogfzto05glTmRfe1iMXHr+0PmMUC+CHD1I90JR6++yaLl48
q6zF7mpp5hn9lWH2fFVITX6PfYmHDzVWLtJeexgCH6f0cE9XwHI1WoCBb/1m0XXiK3YaVDzD2Osy
pe+ILxyJXWViS7BwCjU8WTGWoQWzmYOM8xwiwo+Wue5HLRrMR0+0ovyvx/USVhFnUSCnNFxl61Wx
KTpxLqmh6F+3+0UFvx4aQrttB/WuNm58RECaPh1ZNEHOfuyJw2eJqBGEAAbTaUwGncVuoM6TnrHL
htVpOlF2qmZVpTkImBgkufn/WLZQpGbn+rjwaZa/dpxXQYwpjeYgWyejSrcrFG101hNssU//Q7xe
NGUPFcO68jMy83oHAiqCI+N2qtNJo+kQergenfbjq3FsJd0K447xPrVyzI6VzRRV4yQAj9uJ12f5
jKK6p9b4zxFwLPHXpgpztYryH+6R4vuFVFCYihkCEaNBdK9XNSgH0H6KWQ0hwyzRO+10vFNJZX/l
+k8HvJdviCygB900/iXpl1liKpYg7rVkPtii5M8Oc8jWmEIDG9nMxPiRG3uT+Ad8p5yk9gEL8AbT
XTdBuVp7D98DR+Xufscr1PA5/f4lcwcg94dDSKFj/myAVgElJYLrPL0OMcwUy3Lnhg0kRr5fH5L3
e0AQrcRji0uj1nmecwWEyhOB4SnZYunxCXCizSEIjdKAka+cjOAXA3hNi8pQZ9vT8sdDPboLRUF7
WtBQNEDz2abacV6rfXmydln9NwuQR8xfz9brd6nfl+WxgPki8FQQpIPptMaS/PTVdwQo+39SBaGC
tQlp/YiC+MboTT8mf6PSpDWO2IJ3VMHZgyDmAyOiUI9vfWItaDaaIF6aSCldffJfvjh7Xk+YMiom
3FlcAsBPXDJ8QicHk3z+/bqnddlnLO7UcF4dFrqdGHPHh5iv0kcgwcVzfGaX3MMoTnQk65RV9LZ4
YB6f/gRxCwPv78Q5Gmt0V0aBH0oWITnuDSj4YAOu745wYTsJJe2yI6Ss+70W2jXGza29j/in7IvJ
3wqJi2qZt3TJ3n9q8s/tWVWXGbrypvr7OZAzxkGKfAcCRD82L+qtwyqpezL7FPQOL7bZbBe2MC55
TI5EuyKESM9ZV63Noq42Tg2rg/wgSGQpKf8bnIglA85KiyfUTO0WEgAyfe2aEK6rPf0GUyPJ7mrE
KGD9MaQyx8NUxgD1V/9z5s9clbsJNuQ4jqgdnxuXlD0bEeLzzr4nr2HB4PfF8TtZK8NMTNcDzqg+
HPOJ2/pUOz8+Ua41Ep7k3gcVpJO9d4WCe7oAzWNsDeYrGSNsgvwoBmV6/nB24shnlMQZzhKTvos/
1wNwsH967CxLMI6+vRHfb7p2CiesBvKE8Zqrm76YrK7C0Tz9h7EMw4+X0LqNK6IFNthaAMhvPsaF
kiGvz19ISICMR2Z4SVOhc1hrbRf3soc8qEh1JAN/EInyeEnlIGWquokgMs87UROpQRHfgkyYeHN8
AsyX+sVWphbARP5IW5v1x5x0FjdPE1QoWUdNa42SqWPMqivEpH53Mqy5NuD9JqQrQ+emJmyNGm4V
NGMunVTFQzxWsACPwblKAGDLBnZE1IC+QIm4H1qcNuFk7FJVMX9k3+d3KHhFeAmfg+TL/NvJBgWH
0XVkNkFxchqeXG/hRNrwG1OTINGH+M3CqS315j3T5UU0jhV1HifPIQnyWLSi+5kEKP0Y08hUKfQt
GBqDMwijAmwjuJRA8UPrNPpHzhvYRI+Z6GvQYp4uYx4zEhnHfqnaE+js+u2l5PBrr/kv2LS+PSbi
z68LfUybthgEjKnBuXx46OQg2X9GBfszW2L6ujAv3Lhtg4e0rtRDEcgnwD1ImZuFxb5c8NEjSSBi
QHVumSwk3N2Axern/uh5gcXfyq6CblkK7sov1HgZT/zaGdqhLNn7C2VwKWGDMfMmgiINIScdyT76
Wtr8gBETvE3aCGmENsJsdFqF/dLO6ANumqwjPVfCjiYHpu33yWwHRFuOpMkIW0RFfdKZo07pbtNa
1tzKdbYjdW/BKyiJqH9fq27gtmcQZQ0K7ZeON/C4QI+jw9+aezAdR/ZbmoZvXgQ10xWwxT4t7j06
peTw52vJ07jOT8xVnNl1dIysPc1E+t8rNYEA045sazDGouFa25to/gwM/xcp4TiIcwso3KeKzqXC
uOo2226/iQNQ3c4xI2B0P83pUGVCMPtrNO/88WHdaGhrPXGBlQmXLuMtY9Y+dh41tyHpKFt+cOqN
YFTrE2/WgFxQ3hpPRsRd0TTJamJwqChnm8u/Qtn5mYcSl0ODJdZk97kanahSJptQB12PAl2J82gH
xoy0BGKjsJ8/lglePk5c5gfR259MzrQd4dY5ZFn/YHjTE/LDtABim4oxG7v1QB9rB+L9yvZor/Vh
kAKVc8LGr0f6Pp+FLq884iPLHmAamfWdaF+FBq0pBFt70+4juXCIyPF1ABOQ+YyHjmBIoxVoTAr2
JJywdom3mJY98e0TL5c0P+eOn3YxhiaSM0kakrlkb/EybkNU/1RbckHgCSQjGCzS3pfcERNlZN/0
eKpi0Nk7cgQE/7KyxUPUqDdDnffwjp0ombmiknyNnzIoq4q8u07gofigTp5RUL04FVKO9faKoXRs
aEZpxz3FW28JcvTVFX9q1+d75au016GtE6YpOx2FmjTxpH2s9cGcHiMm85iMUTFDXOWWrYTTUpz3
Vq2eJZEm8imUMSD4DZKa0zgH7M6L/7/TMuqFxP5b2xmSGllfbWBHRnIxkMMsdornwsQOPUImuUS1
P+TeCUp5L3B8r6cEiwOo/a6G6UFzGNCsQQnJVGxZHzemJyowlDU75jhtYNiAyaVVMs9SFXyijlC6
Sj7KZy8QfvzMAjdY4Eob4wbuzyXehOrtup1HBKbeIqCW606D6wQ/T/1SwuNJV7ev7clpzFWmMgdu
cQce4VOd+qYH8ELPTmsI4KjUCHOWNgEw6ICrDFRX+Fkn+lbLKlrEGmABZ1zpwG2AS+qGDPb1k+SI
psMzU9hizAFu7d9dTxL+MsV9RrQmLaLmp8xZxFRsLNN6EFtv+xGRbbd17WPZoaUC5ZmgOgdx+DA2
Q0ugW4IPFBrY++ZnjMOaLNa5N2xO07UMg71qZlUGV/sJ4UYsOyhfNwiISihH8n8zRYb+ExikDKP5
vFwCnTiXyTMATYnzwsK1nMbA1SrJdQJhSSwO+vP/gBfJ4XuEbxRO37SaKrHYgwXEKJlzQK8kwhNM
IZ80L7cLwdGNwgkYepwLGxcmPlsD2R/NtxDk2+YF27cH+b3oIcBWGHiScanjg1s+ZVjKHfmouAFI
6F9c6nemx6NSApdc8RX3QXWIY19DfoktBtxNCRIOev7yhefpKmbWK+afn9MdsGW/j89La0w1Vtxg
DPxuDX1Nu+Ty3QnWXqwV6VCCakNFuE/l1VxHm3wTnM4moOmirdzFUoxsGnPGNS1Sb48etOdRg+mi
iaahjZhged4swFV8/9WCs3qh8yanE11NCNzd18bPvpwWCkRPGMS6JBruesilLdI9oJruj1yFAeHf
sO5Kk0FYcgio/JJEHRQvkGLWtbL/kYgFLr1BdTL+sLFTXluyOCD4/40C4VjA7fblVlxiDCyKEUS+
edhMcQtwghD7nxyMV9PIgsxuJaMLWpbf18eLSMD3w1KrJyXbtgvFgsmPMDmyAFMZcKq2bRIDnEjL
BtehwC06b9BNOjxgkGhRQwVmdjGnh97tBFZIkeTy6wChsVx84snnGGRfCcGKxQiqYrpMEyc+CHPw
p0j7CESM5x9eSgVuY7bdSwz8gcujI/cVsSbvqx3XJUehWf+DU/EICd6a8ZiRbElBdMtGZfWbrTB/
RAPVg1A9N/6Z3THwXIG7UdG4nHiiH0yJ0qrOjEOQa9oeQsu5tAErcSTQmr1MEKkvVjcN9CY3YdjB
9xqn/U+sCF0Nr1DiJXs/WIl3vDs2nibHfVIdNOy6u9C0Nu5EYmDLRlochd1QErOOVmnSyGpsWwmj
f4B4FdK6qnaSx2H2U0hU+iR5PYz4rEOe770cBSTHE4R7qt6jAeqpBU2lYc7z306I9iaMWsk1CY4a
Bwmwrq3TyPypcAGWdIiQpk4NnDA/a9U4cb2qDF6szIkO3aXfWLbxE+wkr1VeASaDEn1cPYI69ja3
JOWyVXM77JQdmi1oQFvBXcqIW3Ln9CB34sM5YzOEJnCaP+fqk3rMhiGjojiUEpf7GIDpV6SRIfvW
/qqnjlb8czrvWHnIHW9RKm+xd2w7Y5jtvrAO7jrlCXvtwsonTIAhqyHFgWuTLcUs44ERodjSZ5vw
BYIbz+d/c0qhr6orWSfsNwnfWakTveeUkEaINfUz3OCX2jEX1bK3Uu7S8utBtZ78LAo8DIhGr4Cr
whRS8ov+dP9df17oo/5uEZL+ffL64osm+8WTtBwp2mPd6Sr/DVpknCHrJQZNOYvzmKiBLmTQCLfj
32NJvtf9g30QDty2Yk5J5/38S+xgf/LvCDXTNiP/YDUuuesZDxLvF15Ep1nQ28yUMUB6k3uLfT+V
aWCE3dNnV2EEQ+TYk/fd5Bo24QmYFKmho+TFERN6JsJM5Zk5miOgA9eslrvddKTgE5pnF5Ne7uiF
W8byb2K4jq2olHbzwL5zJhJLxrIA07X98dZKLUrPqzeliPhLlCWrY90QxncSNoBOTrNjihvCLXJ8
/Ffru/Gez0oUgdVpNQXputjZDartNBq09M7lJxOTDjZlQahkl5mE+9vMyx1h7dEfH8hkBNeFnQ0z
WxEWUZXLbSNutu2pzehUSPX8Aa7Z21ZNJ90pgxbGODrAsgcaayx9kjtdBQmEz5y5vaSTW2LpgX1Z
UnLRzBS28i/KAZ/hOwJr6CAqTbBozMjAp2RFGCF2QzT6Mh6ySlkh65c+IjMDAIxVLFigey2zOSDW
WnCfXmWJyUukya5VZoXr/A9OtPG0nNQNtUNCFUeIihiUB5YHZ53xmuBgK3Pb3sQ61b39PdkcLMkV
TeVoBL5kUpbTVY200I2P0SnvdUAAe1j+Ped756gfNj9U7Wv2tjsnlF7cK7Slu9G3PAjaELlPIWqm
5NAJ9Hn/mCrY3AGLLd6zkBNAM2Cv+BtlT++1QELbKJZ/0fFB6GYnbO+dD0wvQfB3j2JfD07I4byx
UQTMZL1FdeCOHmywKpd352BgPAHfYZesLJ/y7Z0zywF8lCNYqx5zoIIi0rlCytY3b+kP/1tVSXnr
fBu7LT/ryvuW0HNBsTOg56oKq8CBly3tKYkT2+vhfpMWnQ5iSL3XBNo326hslZzK/s+yke388ATv
mFNik1aAiOeHys/B1wcTkaTZnqKDuzLrATRT1w1Bu83ol70wL7rtI2EXszOtK658mZ1pf4Wfb7Gj
Bb/ZU6CrlgXv87Bb2Uk3K1mBoLfkdqwdSHbMrFWrr1SJ7I0vk3jKyUywbBwyuVu/gMVA8uuWBjUy
JXCGAqevxYVV1Cu/P2EKNzztjFHHYt9x2pybJ3JTM1GX0xNfRYLXcf1F+3SDAU+skWNDnZSAputn
2m/5KMv7S91+a5QQKycz4X5Z7sHwDIyTSrSc9EZ/93RIXhuN0PCKDPnu4kds/FtbuhguLWrg80L8
DaXR2kbJPYGxfv0A2o2T/LznJloazTaHzU0Wc6Qs4OXRMrohuhTYqr9zK876npl42ILhmf/fUc9T
EOKdkzO/HWISWu9to0ZvAO87eFR38v4nDoydMcap9sWhvPfLml1e2DvZRxX7ZSbNbi4JDK5d9VRU
KOs+s2C3zAMR3DSb+K+DutMNAI8y6bqSBzZCkDAbeKQvOg6QKB5tLXAOYpqpPguHn15wUaR1s55R
DZ8o2UvOR40+mrv+Zp3fLUlcCmYRtbdBWS7+SkUrImE7/dnwXzFiOT0RhfKA1AfnVCNmk8xqpJLu
Wu+yGK8h7U2R9dONgxLyTThDFAaTzBY2l2aAoWtUzK0kDDEy3GYJfGg8c2kTUygyXGH7mfMeHmv0
uwRkyoOYYO+92tcm6gBgVFD7aFsO1lBa1WFGDaX5SCUJvQ0Gem8viIK0O0mmXWoIhU5gK81Jlqvv
LVDNMW7wwgeFNeAJ5c2b/SG319/zyJa+8JInMZoGxNcxiYS1iBEr4Mk2BtssA6JJgfSxHRrRTIGO
9GScsPrtBT7N06tByevRBN20Zwuo+M5eOA3m80s2/smjh4MXROCd7+nqgaPTkVxOTO1gDGDsI8Tf
KKWOH5sWCwORxSob7/Jw3NiNypD2KQTLhh/jroDszh9z1/wehQW31IR2fZ61WEYwGC1nRleHPgyp
UHwbDMx9sk/0AqwvPxo+ndkx235ji5n/gbw56YHUX2pDOX2cCPnqQuFdv4Gn7igrE69u+8XKH38k
kpqz/2YqvoRkAPeTrWo50TuPTduNIPuW2TQLSki1iWPU16mH3IsjQlcPzrTf9PL3QdFhQtP0WINu
VCO66KJmWA0dvJ4BR9ci2LOWFUIndMwBpDrBDaSI7pXGgpLMeWl5wzloKJuD7RqMGKftk3lW+J22
r7WRTtYvo9oiVoyu/9EsnnPECM84Ol57TGiVD2DA1QuM/kiZGsWxVi/MWBroDQtg/W/ZESy/LIG7
EYK9sNEyQdnsLtENrpV+SQ1gKfRJqxWcH0xasBvMPwUEI09ut37CBxBD+xo+YIk3Bqiqy4G7Qw0w
f4MCXnfpLYbW85A4choUfIPQs9nPIKP1kXbIX+mcs3Ia1suzP8tW9q43WieuEwf+J9uI6gMkmkhG
Rkbt+5EpWNJwZEy9HvkECBxofAeiYW6GPRN1veaBExxINC5/rUHY10G9k4FF7SQdkbe8VcLAxWiq
Bk8BXNK2Ld19uXpMY890neCqLa2GBLdV5bTObN3HZlYEbiX/cWEswEffbFa4r1AGXBBEmZmRM7qa
8YKoc47Hre19pfQwy8Oef7Q1Ag1z+zWnuYhlh84MRPhgYgh/j6KaFYJHDULw5NfikSQmIMfJ0rrn
o3mS6lVp8LbhO05LOUafgfZwJcKsF0eF+greWJO7VYJmOnGPhS984EHH5cC/IYQMj2PwlUtKkqAa
AMERFv19dxm8pl0yz8acu66i+Z2oNGQQSF59moo+jkddEOCemZ2UfKHOOIS3oLcNGCZIsFvP/sVt
xibXZuw5ozjqGA2UiI35hUDG6hA80d4oYTOPFInyr7l7+kUZ5/DGBJCPe6Ke70e9ZevGfebBBWLf
uq21CGb1kb8YzEJNwoIslcmYt9+6Glc7SvBuqBpXPTUnpCX51CAlNpEXLbcdHdnOdCZlBIWUsuFV
dMzadJzHkMNkCl0jQvIVpfnT0AT+i7TiuIeAYdkt2o6IRWyIqpMVJn0cYuzBN6KweAr8SmAFg2Vv
IMeFrFfsCvUPgafQ9ZTNH+Tj38gN2MotFoBMoLp+PQHhSg+THAatlDzDb9QSSoNPpGwYIwjskcVd
suQTNQUR46mRuaaHIuGi9yXfzDIjc+wht1/7N3gxau3ScCAa2EwYlk8Nh6bzvEddejGrwJo8IlMW
Gu1kDQCoDy/NuVJzQNyV/I7bKJN+7b7qr+1aktzfBNRJX7mhc6z2Qvw2gpruojppXgBls2cJKfLD
0X7ITo5i07lXjWLd+oGprpP0m8yRxsufQuJZvj6BS+UcNvH+rNnIv+WyTWPqmI4s0n4c7MJhehGK
z1ETBLCp24oqDwSolvNMAX7yf4J00ZMIigV7cn5NZRRPdEuHzRFN2+q6MR4XQ4GfEte9zDtT/Gkc
sQw7/iVHZIJhExEVzWDRR2Wg6BNJr7Ukx4k8VnJMKyItoxxPBPjDuFTfF0k+6YOf2Y+PWXG/oJ4E
CRHXF68HsU8qyaxoOGzWNHfCG+2zMQaWngMCTLCOOOtI0DKMJu+qLNHcQw/7mJQH8mkkZRH94y8w
tjM8DXOCKmoF/heDKZ8YQ/FbIUkosso2W5mCcG27YEgvTtRwtgDX44rqxZX87MnQ8mGYQA9pU92z
mzKUuweVohzoUsnQ3FGSwwBRSCcT8SM2LIMxOoBOvR56EYA0c/duDja141CmjqQMopD75bQIbxW7
NgewJd4ZYoRbxoW7CF+ETsi2JPT2sY0KamcHD7sFS4dLhVQPwMwmxTbuYy46FjHM/Ww/gF11/sES
1Th9G9iNMce8rzYHwTJJ8VTkYWZDF2QMuqxmYoUOLqWJR0F/tt2wA+qq4uquCqvKB86OoSLToYlU
1flzpq7T1zxxuO5o2WzyZgbDxJB7kT/f0z9mRmjUukB045tmOpD9rGNl/a7dh4vN4ZaR6yuS8rg5
TYHwasZcQV7tOBKS4eBm2QNVOd18qMOVMh6OIX6UJgMZlPM8FdE+D7MqDVoOYB6qtN7ajygQPiZ1
VA4TLyiMei17H29NWzi8bzm/n6Pz1aAyTJOeKKD0Klac5tRS3Zgf+aRrRkYHp6LncF2LUbp/gUYt
8F3/UyGGm9WH/h3gHjsZiaQnTntkLxwzWPqZZsUN/WiVTd6LEAstoJP/Kvm+3h0ERNz4kj9u6y1U
7aSIdP4lW4tetC92UIVRWHSCB8fto6o6NnudK5sLT8DrKcsSODfSsmDIjFa19LIMwJfN956Qhwuf
NhC2PAEDySZJa8IiWtoP3+VE10vnEtixO/U+LUlVd7Bzit4oe/RXHke6wOStlUDETjOb84Q48CR3
T6UXoI4VmKvf4Jf/ONElV9yptjKoBbHPLS/T/9xcSJW34e43AIvR1YFiKI0i9YM1SUb9Uv44uoTP
beq1mSbwLUJzLJ0UQ2WmZk0EaEWJfXHp1EsS8mNJGfKLJscCKiTekNu/alR5NbmWIdfNxrovbkKR
9lA/X8UefILpBQApEoUNXk4CCnDP1P+f7qOZJldF7vND5z2MFMpjWQadHszxveC3gNeXvZYE8AEn
VEwBDya/x1jr8oyIJ8SDh6duzigohwSl8W/bJN9Nx0ibKyR/IEG/L8fp4x2nTudU5htNFQK74p0H
/ol/4HttggyxeIcECHvwEN0VD7aHWMA1RhG4fRe8J7XhQvhMzx1EWQV5VoeaGN1SY3OZKw+bxjf9
Tri/B3PHaJYiSNSvTYvokM2w+SQfkXFbWedeOjf/v2UmF6H7blSF6qRaku9A3d1GpF1CeCXxX/Ma
MddDk0Wi4K4/eUw5ojg2dEY6fqak4W3Eo/+6z0k+7Mug/p3yg/zJs5U0R4mcjzZ+VEtJQocTLWdG
L5o1sfoRe175rjv8yQ88B2tthb/K8MmP+L/QhSTkek1sxHvMZ3Tg6FcQfx8/GmK7n8HAKs7OHI+m
5BUvUhGmQfGcy/SBpEWqA1erqqcbvD7N4iEtuPPbDaMj7KKqhtPPvaBBVM/qH9VX6Zy6uD7ya2kN
2rjavyiMXLIz3Nq5rupdfuxrcCBxq7LFhWjc1C69/oDdh3exnXTcr3d6Rc+MsWmEMMNDq8uRgrP3
6xKCG7T+v9mmkw+9/s9BQz09kFH2/B2HWJNGXcDJnH4QHgQU04cbJZx7vFhFR8bh48YEQu6d6hQe
LkvLzow8F3J9JXD1yUgpjqLPE5+ADxUsznRW1Wow7WjQHEvP8kC6WIZaSUPERPC51GpY3P6vNIfH
zgUrU/7dJ9rX6XgsDhLsEOwfRbBJrVeoNyRHrU4SJl+Ag0eyIGdSlFnGoc7utRK+XiQNnMOKgZCx
CUjZLPutGA1/6lhsCMaqdBCWiXvUWMTUEUVPx8ijKLXTF/iyMtPeoTJDQDEBEJyIa6fi7zBu6/ii
RB2TGFCZb+ZnUgAOnsuCG9h5UNSvYD4N7M7UzHgPClcEuFaj+m1lJdYIUmAbbIrKpjpwYx5NZpYe
ffwwtvo1gZuLmCmdG8WT9X2tVyIpDdf93TAIDZQqHxb4O8h5j0RR5J15kYbqODYueOPhmKthx6GB
IFP+gl6IkAamjKXgPVVTFY4hPPFlF/wtGeFAMQyAsnVGs2/Ea2sYKn4E+Gt0fpHkGFnzoTYjyGo1
6jrzNL0gGcfZOOfRmFyIOQDI3zDpTNLYAFE/xHTtT6ni8JSfJdte496mAfBX+OWeSrJS2XrTu+Zi
pvxa+HyEumTxWZZOAM4Qpz/sFD7vf4Kl5It0u449bRuJJ1xC+ulIqJKjSWK4nPjBpgldVnY8LuvF
SBdTHDVlNU+RcTjnVF004vstOqeBluq9bYIf2+86QGLxvB+pk4Lbd46BMHRbV98CsG6nHNB0bILX
31Jhsd/0HhZt+NSRE4YNcyrDwdSz6Qb8FYVbjiobQPXnI6alT2Y9KPNh2zwoFjiLtJvB9/4lcR0V
SlJzlea1C7cdkMvBmedvXlbfF1HAbnoPZX0u2DXhbuMHYp2f5uC9e6SuXxe9GfyvPpufVYQwb2DC
xdpc9J80KY1Ta8PUIIQobVCcG6PyKHvhLMDDDID3d37jD+o8IGXLuNqTHsYvQm4XVrB3FnhvTLWG
eGEUUTAXpDLTIjfBNkkRHFEe64WO3xCSzEPfmmBlwCm/+d7raUDT8/I8Ue3+63nDblazNGCtBgMT
doZnW3w7j1Y74+BfXnqr6WPZCZPBBa4s7D+/q0YW+9zDiNBhhLWYYCNW2D+xkY2q0mpUe6vf4Ffl
tnHp65+UHIjbg9GxgF2DtoMoMLoI5JzU+oEDfek48An/jFFmWCIvs2Jz1Zd98P6V90KaGpb6yr6C
ExzD8yp6M1sbsL6sM9Vv6J+LW379Sx4U6KPTqZf4vvkj4yTBkL1rBQ/STOZHptklm7XD9x68gvL6
2VGUosHq4tzhMl3/o0UK/bsxwJv4myli15LKBNbGIkggAe6FLuiu135tGO1T/z0UEDTam0KWZyv/
7NRHKVH4sOTEmD6sS9JOZAiob1IXi/RQIozagJ2RUFwHrVGslMqJnJnqlsTPZq+Up98HSy7muYlM
XZvIZ6YJ3zjyPsXM0VkFS1fBZLir9oSNhDlSrNnNiL6CKf6CB88QSzbArw4vGuDOl3zS2PpXAjzW
/L4Vg01H8IoPO5t1yyG5v+E1FmAiotJJQn4RRNG3++JEdY8VahXjZaFXiZznCAzud0rKWKlRQ7W8
YVczs35ZNkDzOhHhiDMaBR6IoLX+ZF3HDQLVC5yRJSoT9ofISVp5DD3G45id397egDye+kTxyKNS
0cmimZAwoa+gmCAFl2qSv1utofVtddvxWV+tnREEkZ7f3qEBLQxBIG44KtmTqwPDiMgFOTF7N6Ho
knLJUHZ/lhis+dm2ZwAAGNr0xFSMTTVxqbPFCA/e4TUHFACAlL+jAkQ1dKQpUTdQCXEBgea4V1hr
LbRRmx4X+9PHgY7gEq81xoKFURuP/gS4CSoazGZr5eSWmbC0qPKlj7xOjmzJttk3ZI1tV5X2K2ko
DWi4gVtuP3Jxh0BcsaA012zK1AMoXfmxuH6UyGAWHgJ2wy5QCE+lhYNPI8Xe7wJMs2Pf3/EOLHMX
70zYYXhKJmoLmbesVp+oTIzFpRB9oq9TP3ak9b5jrUMcbAOPdvx4lLdskKIZj88rO1tNRY3b25Y1
1agxRpC9FPfW5GWfWfbEQ2TEfLBkVnbCcGZwALdG3A5Amrd0JE5J+z2dBYdETg/gewBkiImiHrt6
9Yq2jjsHB5F4R3FEUDOJeg8ZjHN0hicUlF5AVzcIVYCNwogP7T3hmZOHiZbrezNo7J/oHCCXwuzm
Q84ooH4BwUmCZdO0hExwuxf7SIa9OTitIEcxUXanN8GS5sqV3lMUXFfdnBMB6BxoZdihYX8fhvg+
NHEjVisSh/bYjVY3aKrRG6jcnes/4y8yvoszaBD8EL8ibPbBhoq2niXrpWQLCpM+nEl0q/7zO66s
YnUyuRpsiWBBUjjZ/iBMMw47V7mCpTv5Ia/eCzcp8irwMb4/HxtN+sEXRLQ3j6EaCrtwvbGzQC4d
VJV8jBtFgrPfhJYNBUTIXHTHRaCEgMaqZW38xXOyPomLCyBhNexlQeOUof75yuABFjjSqC6yKw6u
C9RtV/cHWI6jxOh4/o5iwxDccAkRKY7fea2Er/48Clj1iOls5d3/Vb7cVccWGyl1wbyK2Gw8iCPs
TOKRGiDk2GL0zwRA0N3zGRUeljfe3xPqRKwVglESLIFM+unHoq2Ksh1Ilghus7xtOtDETA1Q126g
V3973Q5+mKoDqqAJwkmwWncl8YLnxeblr6L7v9bZjuVFoerA7eYkUjsTVdHZRbVmDX/UBPSco9UD
hsyF3ySU0xQ8PZuWEZ+2h98gdAoGyxbHcIpC7XJeb+J24Jo0DeGCiw5H1U3aGIYUuaBU9lbxxuYT
049tlSSv2bn1K03VfFy4Y4k+MgpDwlKZQYIlOeM3DzCGfkDuwQIN2M+ntF0yJiGkkQx1gW3xlVyS
Tp3hOJlSAntDU1EvB4y37tj8oxhcY6kUUWBLjOUrKcCESUqGf2i40i9iHlP327jaKqo3rPB3urnH
sZtMUbx7ccjCLrqFoE/l64L1chgNTzQKXCbLfaIa/UmBvYCvFh8aU/Ml5wfD3TRppnFfQOfJU6p8
yqQCO0tuTxJhxNd4zeHCjSdI6pXF3nNbFw+PRsnueSAUNBSW0st2/MgKimwh2OgzwD07ZVaDjz2Y
5xCKzMizXCw0PdW0a51d8d4NWIXoYcc55GwhJAd2dKE8wYdmShtklio/DHevsZEAbiqNESW5yOAB
NeukYs7VSry30KZR4tG9tpuXlC+uhNwZdDV0628BlzVyIzTguraSAdGJeVfs3U41394ClsLIPtkY
lcfs5pzGnlySS/qm/LvRpRlX1WuQxKT5iXZgyekN6BixGRtazvjHGM3pqgDb4k9G6rYCNa56f0fV
La4XC9dRgk4NU1bWo2vs7bVGN2l63JIV/egNWfSrDqlvaHufuOVHJ2xJwwzHDCvPNZIJWa5Zxgd+
Pk9NUaW/59sDgnTrmQhL4VzfmEEzHU+X/g5r1eDtTFgqgj2bMTcisiHaTqt28J/SJm+vIgvo3LJq
ukvsHjy/AQlF9uVFEMoxlSfecG5lx8MaefYSjhRiqMm/0aGd3WlqH07Xj3qiT2rGOHqdu+aYqrmI
Djw2UAtnNlN5JmRl+Ttx/Q+VqWi952SCYPJsoNhSh9hSsYYAAdQ45lhnr5VvbQZ7ZvQ2FJO9Hyno
r8KQ7sBPncdIX2Mo5LZRGs683/GlevdtsGwWu1EtGvQfbnjBtYN+uB1ctQtwe41o9hwYMEC3xz6I
tHEMyPh8XxZZr/+okWlWrteo2E1VufLeKlwG0GLfdzOIJC+cIpGnHzh0e/6nX/IYp3GZWOjjRpYw
4UWflKq/JF25VuwXtXkJpQmv9twFby8VKT0O4K+aXxQv31ihsrZdshcAOJR7t+NP0wWCNA3+UhSb
1nRVMtIKPCByTkNk92YTl9JOMuqaeNZRI+bCbhpzuwqUhCEXZK9NTUKRv4ttD3fiEOoA51g3Qf2a
qS+dILycNpI76wiBoMg8m+W8B2Dy0c4uYJ7kTmDrJ9httbuhpgKqYAz+7yBCzw7kb2KpbW2fVZRC
15rAx575pSgaoBdcSfN11Qxv8q8c+UZWWOkgM84dtztwqwx+uP2/APDPuGS0EU8cOy3mPllnEjkz
lG7sQg1iMnmhmElwLOmAtq8u3oH5EqIhumtpgjVQkd4sy0RbrFIh9y9sExJ3cp8wDO3VH+onyczg
2M6HqkWfVJEmDRK+Do83pgozH5+edIJ9nbsjBnpAqwtQ+EhFqSAFJEeISDbE1LOnIPfdl+OQtgkR
rkVzY+L71cOn1s8t2J13MF7SfYHt9SNxTMVfvp0legGidvR1Hfaug6fol3daXyhF30SKXwjSYugn
uAXS7bNnLf09RoYwAdRHcu6StPmh/giuYaAVDiHx87VRtp8Pgn+B/pmAg+NIM7aqUaX65RQ/aoDX
5fd9cMwnzFljUg9QBEY1anmucpt913a5ugxY0Ldt38Wvpe4HojB5xdHVbhUhggBMOZrQbb2LCWsT
ROv/zWnp5gs6vVe/fM6TH5c6lgzv2q2KsJziiwxoKIAatoHAOPSBFuqe8orRZHC27+N5Fhw30+UW
F3R1JPcH1RRwspaXvMt4FNDJJsbFLbKVxXE7/BTSvV3nQ2zEbFc4PC8G0d4o/X8HITk63dBhY0uE
NLsDLkerHk/cf4ymP5LCwfkJj6snz95sFXL4ant+Lh9U70voDtb73f70yqmu+n7SozHcq6TZ4BcK
hsHaVWp/2qqXxxzhEqwcGfBqQz3NEJpUucRCiRP4XmmVnWlmxJTBsIU9i2/ifIccZxuvSJ33MkYZ
sqducmFzG7iTO0iXaQHxZAO4aNYQxDltwm4Jm91i3mYZd1H5ZXzFWGHG1urjP/eyVGahrWsaqDnn
COjW+xy9xHfeJTRzfmxpUmJfVernGfOsUOK1R2euWHklF6w9QstF0rSk/ChKroiwDaxDwzSUpV+h
uEq5ko/adfeOr43IL/2v+hoggVfubR3kq/8FMSFr/FBZVRggtyfeySjBrH1xLakZlD1265u0QDQf
Bi6sJH7ckrSuatMw8nxYUXdtmSQypi3wF0XS9Sq+BIuXVH1NxrxT83KTg71TMQiyTlXM+LmZwBP4
3bpw4hc7Td7NI1RMywAVX6EJZxZzMEHz+bYcp87IW7SRo9FU0mtDvIXWZ7aBeCATAPCqZFPuEgV4
J+o04ep6A6G9Do9l05jFX5qz4jpCwQ2qhmBuRSjYbFMScwNwtSU+6EHvNKb1uoO8l2QfSlsK/Jet
+w0sYJOLkgLpkG3In+zrCk2esCsFrInYulprmQcOKPhXo2WptHSabZ+NcXYx9vXq4UbYg3Fiyzal
EoRaDYp6dHs/fIkf+KkhGZZu3i3U5eFlSbQuyVG2PF+y72XI1JkpZ05lqNB9Beu8lL6YlqUg8XCT
JFhqcFtShS3CNZgmiI8Sj+kBcAEGZW9/HTxYDme4GJMdkgW63s+80zU4Bn1K87AjwFMyZOR+dvLA
y5t5Jw3OHgmKY2FdHQTJXGg2j/vXXX4enAdgNvUI8yz8RvwXTzbGJGTZBLWl79DUuHHbVBQ7ijYj
E5CUSYQ+EwqFFn7cf+Lfew3eKbF1Y91PTK/nqtLqLdSN1wmShAux6Dir8q82u6eQ6FGLqpXB4jjN
CQRGZKn0F6vqJE79awJpukJKvf2AxEI6F6u5ygDteh5rN2nvVjZ/kmUpWvTq2Qq1MR4yNvBJnZWk
gg7k9OPxjHFmZhhRdb/i7SeolNBuTzSaRWJjbYFl7mA+CN6/98xcK2He9IVC8UGRFsA6CYT3ZWXu
6+5DJMjJdyTww9FigAry0OxH9qcEDZHx6T5kGvr6wU26f4HT2J0WY0qbYChW/r0fzw/8tWaN9RjX
EQar5DGGkuWu1uAJQ3j4PceJqBmziVm6pZTd04scbn6sHpB9J06zqRJf/FuHGXEs0F1GkZzS3OBG
BYNm4eCkmj5ULkPtbd30YeBwssQQmmD4a4KlH0NXTIYF6x1Gw3P75KG+YQbP7AFU3Rsl+II0Oici
3f9uDP6nFLEq01RglgJ8tANxxDjkSOOwhdWjWfahxBsKawQRF3YViLDGLvKs79VETIZNwTw7o6Ju
DHDi2RjX+7b8lNUMwnJaqI+TfPUrcCXjQI+dwQd175jddM+iH9Twr1J6AqGnpBH4AKo/d0U9vKlC
qdqRJ3CBa0F8RH14vabpeG22P/9VVKcq2sGarFKuYVX9OOtm3GALaPVgCXjTCN4A3QcMOK+yX/Fq
7avXAipX2AjiG8uYgtYWsrBb59/RsakhO6brGPgVGX7cUUCnV5C5PnBakUVqSX4Y8rFsCSXywNe3
cBhiomdg9kADgK42s38kmFGPDcUlN/rD/rI+FXOBYwWVgSMXB0BjBD3kBDBqzSdL9aN/Rjr+pivO
JL43bg72EtH3w3I35l49R8pmyw2Uz1yUSUfIg+at7/qNlF5ThwYUMCrLRXRjrmG+GRE4gbF7kI0r
GF1BxqJTAhhMUoqTQJxolVJyi5/4ncMAs0UBSXkF2fppSt6i5yFvSFUS59M4fiFuJZZz+e9O8hkI
poWf+Te0lr3zLE8HYvryALffJeDKxWXCwoxkZp0gmHME1DbVe9ypZ+jfqZQcJYnY0Np+b63Y2/A6
WzqOHD/ECchtLTfdd29J5hH4nEqTPApFyH7AyzOCE9a7gPN9ewD+rYAUmLG0T8KhycOuS56xMZnW
zMwLTcMloF2fVn89B1N4Wc5k6ffU1VVkuL5HpZxMSWIgvq2DC+8jkvi+M9Py41IWJJYhG608CtkQ
Ihf52UFs/OdCU8fdSFdRWqbBW+HcjjBGXIto6OFjZgxElfMEMajDIz1o6N3Iqh0fCBpID3F7RZTX
GV0DPqfDj8ZNyCsUWbFur9Eyy0u1Rk9YW2CGD3m8TJEdBmYkr2VBgV5neA5j+hbG7SThIYU+jgN9
T7ys6ORyxEVtAtSKBfd5SkRwVkAANn7SA//NXiXtdoDhWRM4LiFCGQrxVU4Rpe0WiJgSmMkMMDnI
c5ZN3oaiz7I0pSeRHK9ixxGTgXjpeTA03ecPrJwXkIVH4AV6YB0Gbv6HX4b+b+YD0c6Nv5SL42os
NPoyY7KdWG1gh323PQTp8bc+kQlmJLZMFpH4bmSx0LJ5IsjEUU5Ll+QRsB48WVWeyYG2s9Gh/L+W
N63U59q/4NH4zemp1bIoxTxdbkwvLM7cp67oKK3hw37j/R4bCLNfh6VLpVf10VzV4vY8c+XYTF9X
t6+6FO5dJbO+dsX1+QjFM+rFBFDpoWNPQgPg37+BAMb37mKYHSPQ96eIHNFV5AkfiYj73s4zGgpm
65naMgO9Soh4ee5GzQMCYApOBHEPvEidrYyCHEjYkSGUlq9KBcA+x+Uihq9oQY5TgRNlQ78uTEs4
bjgrJmcH4dKIr3+HlhIitLmd+3lWwjdDOUl+fz76KhsTQJxSVnEyhXaKpr3UzeA2LlRUUImq5lgH
G8In0buMryMnNRYTkka6aNyGgiJqvgXc6f739vPBXX7W1vIQBn6slZYFnSYHfCxIglXrFdMsaka2
F3F9t5vYJolAV1cMVNLu/3HQZL40/seoRK9HzU48S41F/1d9yZT1jE2+SnWQKbWDSk5ELXvx3akF
CELq8viTLgc5ci27Qb9iv0kkmShaPyFhqT4Id5T8mKh3LpPZ9Szwk08AeiYyySotqAoTxdTMeHgz
+n6f6mNk8nKMKYm7EmVMMB9YJM/xKa++9gpKQAn2mVEKocYZCUtLO8GRY12rqeABsh0GQsUd1/up
iKO3Nkt4+XWpknkr+5Wwd4skLeNqsYKZXnHiSnJkqXIrIMzwC+1Lgm1fG9aabi6jkeblMcISr6wj
9qaEMs5MfAAqh5EXkAjVTG+xqacvfYG7qPSr+nWFQAuBMDamRPVGtrjRqtRqK0Mepj+N6g080d5H
kjFluWR4F26vdJ0AiOKEhFCCElDlbmRCdvs/mZRFiqjHNAnJ2gWswnN27YMeAp0t+T6Yd6VjltDt
5GY/mBOZlnB4eyx3BMHondBT0ZU91xUltxSH9a25338ZJsw5W1WkD4LufZuqY8hcCi7nLFm3q9Yu
5Xfda9+KZLhT/bk5pAv/t1OhchHPxK4iVqYYaOgEOruTE/FvellZnutbA7c7EYscmvYuRNmEw12p
bLHD/5tTXQ0cYnxqaulVK83zJ9B5YX50HplybYJj8MtzBiCCEq7JipYDFLvHuxWOcbXAnJNNpQk5
ZqDUQMxqPt1T5D/Q68dOvZZ2MWrSVQ4P3p6sOb5pAHbzwJr81acISaelOsPj7WrLfI/bmrMUNFG+
vZGqVsWMwt4b5WUaCo77oQaroklkfe1LuasaJMF/hhT/I7pwBlwNyTCmPoC3zq0KAB69rC7Hbk2I
G8FwXQbfIdlE7YLeG3Hu1PUybQxJQXMZsnbdMoq1OjBxYEheeSAoxmBLX4JiQhKkviUzyNQ+whBy
mB8RX4qemdkQyYnv381TCRdCWO9QWaoVQjbC5khOYH2QSpUY/rc4MyrRN+0A0RII6UXltvJCciCI
2jO0pbxvzbArrGFVKm5UPK29mjXPHrKfKFu9mC1P2hbmkYJ+tfSfWLaKWy6XzUksJFutLDJ8/Ack
BtajLpYToLDn1JJpnJjoZKiQ/azEgqK06nIqQ7ZRq9XdtQhfu/pH9zvNWPX3Od0fm+KCx+S+fvHF
osmJIpHooC9Co95NCnlnhb46hc1T2fhKq2X7NP3vBBjDox7ErKZJ9IrA2o9iu7MVv7vt3uwjS3bL
vTHepLstyf6eZP7SzW4EA4A7PtkOzVVSwiGwLjB/efXEircqm18aL0iiQwWg77ZLAhnZHGRU0mpc
2iX5hpysmiDxAoHC7GUS2zOy8Crhl673sxU7baTLk1SkFkzKC1U2XT8DpsMVH9UC0CcN2DFAcxfB
MzeKNM0SiUoA2jGlBVizVOZrzqRFvRNYzPHfiR2UzhCtqAqvXCt+RNxwDBekEnY1d69CWibhbNVF
V/nurU4IBJ5w3qDR8P9D1UP2CEj4KGlmahef/shxVB5Lx4KiJZ3qkI9No0ucQ/B4IGihWZZg5/pO
yMSwoFqGc/qG50gV3Up2AVKydduwWJCWiohd+z7fb/MTZw4dc9hYc6+IwyLepR0Mm83TxyRxtJlK
vmv41ppn7YCJ0MrCMQm33/ysfM+chaFWpozQB7AjHdEq0Qht+/V8qe8SOgWOJDQat2QJsbK7uZ82
8Sea7ifpcumDRQDs86aq4DIO3OAKNYZ1W+1gDFLD/6duZn3Y5fwYwG2KzTDVUgmGqamXgqZB2CcA
zXPksvy+z502hFrY4vG/g7s/W2IN1R/USlVOgT/n+W+SEzXhuJP8fpiVIrsHwQSQsdWNiD2gW2B1
MCilm5MXLawavSED3D+fU1JZe7zSz+WIjIHiyCvTZoGsMTrF3o67oAwSlIdtHaXxW+U/W+ro/zIe
1+RsU9y7MsC8NvbZIgGncvhdqkzWZ/UjnAAUfBpLcTa8c9zY5IibUIdVMkBdVJZx92fcR2uyc1DS
gf0j786hNRzatDYw7PGQhA3d/uTZYrKHXcNjfDyBK/GYhkuv1lnGNgPk9PRemj00yJROAiaAXaL3
F4u8oMU/kgT+/zxLW6DhVZW8dVWD9px9bpX5NvaWJycSYg2v/NVGc1HnBlQ1KA8r8VlnkD8b4Fo7
jGWMM1edooe4e/LgGawC88+QWUGAyCrYWY7ezTvm/l3tcuySXGqYUv0bC0DWwZLqDZabzL/wI/DF
IHzD1eaAuNvfaF2QARd5Hmt97NdNOALgkk9vPNvOmBkK8CPJ6LpPq65afiQhOaYnYE/p3Fy/Enac
qbyN7F7iu4pc4brtoJzWQzIjCyzZyDC5UpV7HD5vT6VNJBHdNvnlhaSGGJkxCNUivVT0qRMSFWtA
uwad9biBXV+pznp1ddDww/zSXt9loEK6dMR4VZlojqnY1l24pogqiNbytDeRk6F3Lu9Creb34+vu
V46iueiQzkyEMbVKKIaRBNzs/52qNi1EnK/ari8IMUY/20JZXyPwBLzSsYMZpznyC8psoMPBq7Pc
T1a2N8x+i2KwO8JTmZoPxYY/ANk+FZharDjRAdjRYh7GGawIGTiRlBWnkE2gin54IZfo8LWBpwpo
w+GhHsLFAdhKncfLpZlDAKslsqvkobOx3EmQxYrRUgyW3fZ0hU7HPs2jLWi7+U4LfPFGojo4HQbi
W0QwNDyV15CmhPKwxNlxjbt2ODuJzmb3ndnxVP7/AHoqToY/1QAxzZaKnemcCYfrpASNR2N+Caog
2Zy52ZGtCKi5l7P1luvkVmhDWXDrY8w+CCdqsYKp/+C+PbVdKVQf0d0KZtKfCtZl/LBooHAa3wxi
948jrizFvq9ty9QkfbrAhT5VHPe0l0Jakq425KCBOSzfGdB7uFC2keHf/sxfTwOm6cyHMvPYqBuO
buAsIeoGd90+Umgn2+qQeQtSvnooDIWAt5e1V0NSFK/UFjoMv94MKUvhCOdv4aRa/nhITY5P6Au7
wdyCMH9Wx4e88qtgku+DEOvatFIw2cC3oqwXS3l+UNDKkHG6iyMIbF+fPCcc5Wx2PXrzm70CO2EK
u5kPqYifMwO3q4KcTsyXPVzm/vMEHZeW5WY9fgaqEJGXnV8aZ/N4Fyd0NuKE78XGXu5v5MTbEyQY
xLuD0CeudqipxOLX0Drdf3is2HGRYUc0QYZSOOPXIyoGJ83NUKEbJvBFScpcVKtXsL76oOwbtfGk
NK784wX6+T+VQ8jtSuh+J5WlfZF/otNY5QPXq/kOcslm8qbbFMMGwi2M0BBeFrqvn1Zr3ZRqn3Ww
ExuEFXT7jbuRrNCYTQmtwNNx0qUV/ooCUzAFQJr0GhKj4y4BZNHhE2dhE0nveX6ehKiLfMudgTUx
alr0H45jRrG557XQODvXd7Js/2E3wuBBK8zAEi4m9egGLZSTCcsfac3CSP6Ne102D2nB/yZ9W+6c
Y+p7gLjwjibfRrnzgsZ8laABsGNcQgnQ/OFhvlLeHVwnvYnclVbmh3zM/6bhAfnrU8NhQBQ+ZRhQ
eaM5GBbuo/iV5ErzkZQCJtIBbbbn+HuqACbwO2vP6whTLaUwBKJa+GUuSGeVEy9lSEDFrIkGgRoK
6dtgr/fW7UQr4mOTocVtw8/V9aHEIWOC1wpOgeUMCeD8jLVGrTRdOF8R9GUK0XDmm7h3lOxIMMtJ
2VLTxrtRlv4q3bGj9uAL0rthvsmvgNJTxC7A1wPaloCZ5x3M2TQgZdsgk6TPlEkswwxfE011M+bl
MMLoTC6pEPytVCdFv8FPGUQXNpAz+yC+v3Lklj2x0G+sn8RU0+HUMHT6jKdcho0wPnZy6l1uis0O
NRnDyxuVz0RgzKJH9dJpP1KkAPyewVTYJ4F2qvgbS1qu50tDzx6XOj0ISGVmNtp/MRTkvZitvQOs
TYqJDTqZ2B0ESm7tfiGWbImwaWgU5DAVk7jkF8sisvn1vx9XmErp5yXw2Kr6dmMjnO0/a1L+h3mk
jHHujtbo2fMrdCTlFZZ+NdWlXcGw0PYmeYCUvPdP8CJzODSKj0PEggRMQel9fs2GE9qS/Mv53Khj
8yq3sWJ5CZ5PKclZnZ3vhlK9tzV4fW95WaqA68lyK1yp/lomB6abWfw38l5p5nz+Cw31rCay0eBK
+7lNQUiz95qxGb2zIitH58TzzWd/7PD6Wd9ieCkqSZfYnaM5rl9K5f7Bw/+0yA9q3LDa7RQE49+s
th4GcU+Us6cmKNpNgxwyR0F7oenAPHgD21L0iJ3ZkH4H6uulaE3ds/QwCdERTFLYcBZL5v11EPd5
rTUoNgk0y+FkuTus02C0M0WFhrSe+w5aJl75QyQRatC2QXiiqlu8jXc2BBVQGlnR3mLZJCRHGnFF
qhHsxzX7pk95eA9zarGspN+8PJqT0eVY/RF4ymQEJ1jqYdNVkCIPVmWd/rZsVW4B7P91PUysP41s
ufGbr3YqofX4jjmDAjZKmPiDYBCuFYlk7pDfE0jFXxNZHG7O1CcvSiGU/jtE+NkNHJOZevAmVoWH
5SpreuqH55YGEiBkdHL718p+1ELu8GPOIesjDcc3Hm0vzcYXYhyDgmVEfVnjTILRjfSKBBHFKRKI
vtDzxtGuF+KHIn4GSmytNrxSKt1egc54aF+CvF4TTqfbjH7oZh0WXPB1S5+cgrvb6zrrve6UnqCo
ZhlhTYxn9JDhSyN57JRfSpekbsg0Ttd5mQseBWxttSCIlVXCLrWd6wRmC5B/lHdzdAmhgYHFW/AE
vjoh2biiRUEewAubdfjLlppn35lVPaNO+vSSutkYV2crHPLPwzqOKDxIyk7loTYtynhj6hjViKwA
pmeZhzK10jnVyDHVRUNLNEkawNF67A59F9s8cIb9vCB/IBxNuynQ0rMeaV/G8b5LqU3N1URzC6TO
EXTEYqYnSOQFWmqC2kxmti90m1/tBNsEkEYnbaUErQJDt0ChSnkMMHQkJHT3r3/o2mLBIbXnL+oy
t6jIZvd7NlzuiI7e4HyNe5PYkobJ6G42crRuoG4JiQGoJaOlKCa8Up+2xdHNon3EJ7JMYlECiGej
cjd8z5UJXokpfW9vLz3OpKWM2/IbbAkvwtkDcT9BKaF3ak282mN6fFc0kCtlrwhBBMFDfFbji+Dj
p5v5BEy5kfeFR/Rnbr+dvT31yF8cvL2Izaq7D1il4UL6mtY6Js6TKXmMD7lYZc1uTyKY0B6TSiZc
ZuFXD21snYlcP6djLGDW73iss6KQJ0x4WtPpw6ZuA+Adu/Xg4xeOddPyzzMHjSLu12vTIobJwLor
aWDKA5GXY82E2KuBG1oKg4nnhWbxEpZPj0bmmTzl9/wcdvByqSdyHc/TTF6ZSCSWDoGpoA3K4tuw
CLdqre0rcC/JoZKy6tRwHnkgq3O0Ragk4OrwlY+/WAta1qykWTgkL+iPao8CTIqDg/1G5pqpxeOL
UOa4bhEFW2kL6BkjgnLKjQ8yMugV05SrL4LxG6IfSaArlJKDUJuAOt+M/h/nxCN+qBdp40rRpzwn
/oXZZVELzaYp8JqFxXnyBR/xaI0jChLAQu0yLy5cMZq9RXq/RwVpWlXkIEmtk8MeZ1h7/I5X4dtH
vWkX+s1sYg3dmQk01XdLUKkLl9QUhXCBGZpBYUS60mmKov6Wn41FxHstafpHPrWVitiPwtjBM2Hm
TfVKdjgX5v+kmlZwIvYMD/WI3jKG20u8rMTFVywi8fhQg74DfUSD6YX4AEsmkBrd3Un7dByPkEK0
KBwMqymax+D4pbVx/oca0DsHRacI3+hHN1GmY/SzkT+j5sv5h0rhoIuav6AvYlAJzEos+6B7cZrC
N3pfZbDfr2G91C6RBp3W4ZkZRhnEfSIfh2Oic2DNfyESHc0PRLENZVSTXBpcIMl7Pu3MsNhJfxQH
blNAkOgONRVAtnq32f+7JeJMXwuTbHq8ftzyO3VWLZD0oa6BWWEhgzXd2wd2pAu6bXPLQwD5Uaot
ckVZsf+anu6Uj1qME1N9ZYnkNB2c323alByVaRtsq/Whqo80AJ9sEmPlPZrMHZEcY4/i1blxp6EP
qeWynbflqq7FPXjdJgX297QLJ8UCfEJ1obL/FKs6juHsf+R0pQOQJeG25MdMKhWUz1kKizgQp9H+
I+7e/t6fKZBWa5e2rdLIQLpqHxYq7+9SCVEfg0wfbnhp7leErRn3qGRMYKDpAWntTUwnYfLlVTTe
tLtENeHQo9MmS5oPKXCe/lQ3XRIRzMd4bnbG1K1TNYmuY1iNUSlAAXsEZ9WBzD+9whDTZE59S3fB
ocVKMMUlCPmDV7yM1LtitB8eqiIJVhjvpWyBdDpVOcmKmAuqhh90uctKK4uzRJQmLnL9vzjTOe3P
QmYBkRWzoZixFb11igck6CY3H9nKGzZL49qk2CPcA/KL1M2eAxzr95HjMbYOEHm5Yxf7/qe8i1rJ
258aRZw835GFxZ8WR9g1WXIBAq+527kWF2LWgDnkjyz9QHIUWJEj/nnOeJk+DVYjFqEFO0gn2WJs
n7tHrDLa9rctPFSu/Fs+fSxU4KAf9JNM48rwvdSG8GLAJnKwujsV/As77M6YWbyjjx3qDm7vxbWH
RgtsNjEl08yqlPOQBlbj+SMKu9BoBZm8MRqyNh5JKpqSlBh6r+m7PMHdW1pcvuhYfOlzQtgJo3jq
Qr/K4GPOJfOxA5emgew/SeouaJZXu0GkkHvcjErasPVLUCh2V7+Ku84fa6PfOm0vgNfDYPECCe/v
bAB2u6bFoxJJcBWhQVa70RgJcaUwwTS4ILZLZUDoSbp0BJMj2tv/6RyW+J+oJFzpAcNZBU87IBSS
cpaKEYz7OY4OiJKW0fTwKtEPH54C28HrW9619+RvwcuaeTCzcr/r2lP/qIoi8lDNevi6qFa8ECi9
TRXOB7eqhBm+VB0+u6S3s/3nYcuFTnp012seZBVGjhQalZIxpqNlmcmvTPJ+SW2OLzPeQPoSixAC
baRnhEY+P0frh3BPyWu/OJhXIFmVLyp1VqAYYoqEeuoi+4yig6IDbIehqAZuj8mtDPpWTPM6k7FA
e1xu3BEu6VZtZSScatfVqIG4qh+arCP++bY98drHnaCzONnoV0TmPhnC4YlEu9YjYEf/pX9VAbA9
sL/4XmY4byX8Iq3m5HUJEwEJmH8bNTKNZjyK3cQk7mxTpoLWS7jvA3M7yuqm6l621nRW21aUgLwB
Tx8eb320elLEQ/iyOp+yZ29mt6uGVujjCG9jvRfXfkQXtoalA4urAZJ6C5GD9+3i5VUi2Ys+baPc
ys06XB0vIuQdOdmdQuLXn7TlGrPUT35fU6wvCOXmmYe+BFP8CvI+v32Q34cbcVKgNqGHK/5qLtgn
4zMm+OrkjfnGhpDC/wCUpNPN13ZWX985YEhjbAW487rieqNwyC5/y71Hbv3wUcCe/FgYy8r9OcLO
AwSmaumC9GViI6CiPOB9U3x6w2FRKY4Fpx3gn2FF0C2oWXzWt3DHPdwzxY+TCck2cB7Y9pujTYDg
+E4HR2FbYPCbYFGs2+3je5VnpxjngxW2pLcslWiqkQ2WG9w0OPrVPGD3vF9+zQncjCdcvZpkbwsG
tIKJQwmn2NLTwT3iYCd3J1V7Eg7C7HhzWShfn8jVymwWTTeztSq9usuvK9XZJetfvSAprPSmh1M+
bLx4pTRJY+PslZaCjF+IGo1+A0CfEQGaL/uobV1wY4prpCKikpD53HCe/YednSZwZunMmw0DhFvO
qCH+c6JIVqfbI8M8VHdoytI9v7WrS3VLNL+5FYHDdQJDNWPsCknl+b5JVhnOtAYVMkxivsl5Esi/
CpjZA9RimlfUuGrVUFVAOpELitp+kNbD/63d87fEqAiq0kuuGL1UiTF6k25EgYPcbWrM4us0Z4KG
0bpQaM80eLwYwEKyl+HCQvy4dirKSwyU72r/Im3HRyvSKXEVrACz1ANMIDJQLZcBLiGGs5roASfm
XX8gHLX01nxjWCeJl2Qfb2yn/dN6GLB1ksz4vCyf149dGSieK9V2eBJAEQbMYLHS1++DFVk3P1RF
Q2Z6frELobQ7koy5YTJQUeQA22k9h5HGkuBbjMcqjsaojWVuNkU90nEU34kkixpcMttEa18D/Id4
YgFJdcfoQs1HMCzpbqFxAYMZzEG41M+pT48r7tFC5W+99MU+qLaHb9ZKMDc3RggSlECfaOmFs27l
zSTe8VCS8hKmzTga4dCM4GoJ7N7Cpy+ReFmYAic+ts7gIJKgvFJV9+AKv4oQhBGifyXLmw7S6ewH
f2KI0kcHjBC9W+T+C0etO3zvV6wh+KrlftWMJ9GwL3Ddl+PHBwNvIisRMengpPhHt+nygdV4X9Rn
ZHYtcRDNof6XGUvZCsZZERZAflGq5IHU15FSWJkoCHFG32Lzanbh7NOhLbATT0oC33dm7DYRqG3P
wOz1OqK97LZAOhNAkratFKhFQClH8znT+6ynQeq4hQ/72XeBy9SMhTKd86bq1hDp9SZ6nAI2nqKK
30LAQEj6OT3g5gv3RdD+2TFDUtdkJJl/Uj3vM/cANebaCEY49mFr9w3LSWQGYJ2o9H8ZtyAKA/hL
KlZY8LGyWa/SfjM/UFNg4uH+tImQzNwqwb/Y950k46QlxKfJv7EosN2l9uIXw7HwMLg15kLH7KEL
6RnsKcL+HgHF3DNosjDwrulZ4K/jUnbF7eVULs9KmwJh3iLxIKA4+DZAVgIv8IqxUK5hFDxtX2rf
KX5T55Im3PXR7GYoGgeyZwvL2jwrJ9jTg6T3zUFae3ji5Y1Kz5RI0c6cVlJZ//TE6JpJ2hiXgPdX
bu3Er7hZ1pVBCMRgQZwp5/PjcmG+5RhmxX1KXng6p0k79sBdMcpWwKaEz3F2iBLZvcza1z373S7l
l+ap8u1sglG8KlcICTctno3yTRYNwlxnkiMpc7sI7miyy9XwgZwuSCUZ6bTlc8cg0n4dYdhAb/K8
ea6v7Yw2wctg9eIl3B3kmkIo3EAyUUGzcHxevrk5tJqM04BIkPIbOVaTxJVH3bMzrwnTVZVRfa6n
X9gN3Ah55a2R0Oo9dD3pbHr8SlBNXCFlm01JcmcQThCVhkNK9LleIo+xcIwBgJ82YjoveSzeZZTY
B5Fmx7B7ASGfYOTTngdDi4cbqySY332trLa7KAYdmzPHkjYDGWFxe01+n+SJ5Lgaw3z+eW5Ba8r+
fKVhr+d1BsiBZ5bNF/1FWKcyrhM/a/hbHoFc9OWdUZsCRJBHSlln5JyLuSAgpX6/6ZWP3p+h2AWc
faH1daFXdI8vmdBHU+5iva6o6lPO0DGPPTkdDCNf+Lw/8jnK3tXhrye4QZPKUhB4RAGECy1zuMtk
E8WxrdRSXKx1qzWU5ZwzOZ9Ma+jKFx8JXexbeBBNjkP6Leruv1SllorCBwgWlv7JmdaZjHcghD/Q
ewnn8w74mXgyMShBIG7aA7uNdCL2q0DO8Q68wJYGNVvBw8/BhuGDrVrS5UxprTEsZs53WbFBZZ5E
4LLLEUsflqmFd3NKeFCDQXQs+VRFnFPfSiUY6RAm96AeD/GWXGw0vYKJYst0QWdLoWNMs0pPzCnZ
/rUVGEr3hTslmGcMpQX6UdmWWcuaWyVlP/Hx7h2mDIrjkmHn+tqJt+XCYKgJWR7P/P7QobpZHzmT
ARSYjJgKZe2w1147QJsBp3yKSJu2cV47BcKAle3BmVnqFuNtaBVW8utJ/Kn4GhZvP/B77mh64X69
OQvkAAmncMMZ/4LD3zzYiicUJGrsB2Zfh7t3qXrS0RxdQbqiBL/SZLmg+b2Zs7Cjr6KNT5Xueser
dsPKhV+Y6CCA+vXnDkWSd5w/a5IIL4sC8KUaxOwCPCQUO9UiPzwM/W0CMTQ/Ay7/IVp5ISRJ8ydN
5GWbhqG+ypln0VTd7H3oictE/iaEAcOK54NQxAZ2YB0B+rWEcrYvyZNbHwRyrYob7LwpdwE1ppGf
XQMEH33P3+hVcbkxU+xwP4A/86GTUiIBn/jSa2kB93nkYwftx2Of9XFcIpfds/zKNBsIZuE/EpZg
ugUUP69HxrHlzWAA82cTb+p6hFmijTHQoTy24N5OP7vyaFJhoRkfPABGzbBK4p067iHPDtwT5hGq
AJT/ds3RFpVKsqxFOp5oAMOJi0LicEA13LCPFb9mGAP7oozFBv//F3qcd+FtYmjdl2G0TEutljKY
/OPnOOdoEpCwvqJh7ZrhfcyF1wnKC7os8HbluuUepgzEFWdD/eafNhr1wObBlOcx86B5XQzjTVLC
/aFS+cLquWjkuCR0IR6Xsrrebi3yZ1RvMhO3THWOpPLIcfd36YguJtB8IhjSDRhcSis350F3b9kB
8WAoiz5Y3M0YXlQQ9eUJy61UNgj03UEEgc2+vw1OpGI5JpRgblI1GezciG2kBJPRWBZinoiTlb4D
AxvVTEEbk9CPcvm0k4J4EcP5Lx77kU5TWe1rMUBw0mmnaqfX7nfUrArWEvWzTM37aPNdW5R3UGrB
QPtr1e3fISjKuRhq0aeWpyER/Pwu27IIcM/d6921z5s+gjyP4pUAiUXTXnYXFORKtANmxv612TJh
WEd20v8cmn2l6br7znyCYV1P0D2nBCKegue2trcOF4L7RSbZFiV2EKCSLMoWZkas8U4OypziB8bW
q5MJ0Ihs+Iigxiepf2fry2eq710fGkc4ekDuqQKLyQdNRZGfCwHKu3g0T67LtfTK2HXJsT+72ja9
2xfNcRt5PnQUyQsJyER/hkC/BxkzHaTuowLWO3Yu3DZWElgSXYlYaunoJVvEMWxdBctyiFQnvzg8
ZNYz43foNfXE8dJw8m3UJa7VgYUS8hJbO2IXdBsuzA3qcTp8tFpZbE4jfuW8Rn+UPSlQDz73agyq
/6iM/W3spJOSVShkE4+9tiDRyxbTmE3jbSPrRqH5RTYsGezAawk1+ZMdkdumj2BHD/nheQfKHtBa
Fffdg+tBZA5+0o2D+a9HwZv/zcl0BbHdsPShUVTDCzzdfh1wrA4raODYbkjClmSdumjUJ1vzbYXI
+BLvHC2WmEkjtuYiXkP6L7Ktm9khVxYuy4I86bJmzHhXVm8NeRm5L/qQVqZFzB5fszcuMz39uu0u
6RN8G5JsgXzdy273P4UYh15Hzrx00KtDXJnJOeZKoZeZQoKPBfCvKaWo/8u1SVfy5VdE/ts3DS6u
IDwkWQ5CeyIVlWG0RpbDrH/QVOWAzFrUpbf8gyPO7t4nH9yvANPGwGOdyuH4JHpWJxKaJ2mI+Jgm
0XMBZAUlpoBJBIXH2iQlxZnhOLawQ7sz5Jv/0+nK/WddTls+V+ss5cKkei58d/sjAkYHYY7FoTsl
RfQIs1sqy5f/4X5YWtaSQnXGIXEluzc5Cl5pUClvSMeHAEyBvbc411DiA3htSIuwFlqQWEexd2Uq
A59dVkcEdI7tWGXsvMJyVE5XGzsTDjKcLZU4uW8SWCafofAKErFJmopaJtv8/znJ0/BCKhL70L2O
Y+JwLqc4MLRG8aqP2l/5VGwh/SIuSXFy/eYyY5g+536GCdSET5VJdnyPriTV9Z/3hnDzIOC+KvLT
cS+vuM5j9Ro7Ndw2UPLhqbeWIwtnqY83o0NRKhjT5otsflQDOpwuZyq5iSAjPQ3JjHjMm511l9DT
68TfCP0NmCgbWUPmaKjFS/RAfoSWbYfeYDW5FaEHeZhzstqFRMRmsu8W9eIhL1TaKMeh9lLjO4EF
K73exT5ttw7n2PkV22TNEujHPQjUFI6ka6uJrxHVzv0vQapIZV2VCMi7ITr1fbPHf6z0RMSzKABx
ssR/d8FnIbGOwz6idTqWv11plBetUptI1R75jQ7OOVT9MivosevshudSK7OR8azkM7kso8uoQdJA
Onx+HIh70GogKr8SotR6KTEWeE534m9O06Z4eEaNHIM5U0wFeI1J1Sn0Yl6Ib8ijhsIn7vS9KiP2
wPVEcn2HfM1VZqUuLDhHNBXJQC1wq/slJStHz8AV0ReeTGEmvuKNYXi65uCeeOT7mDiABctlc70W
WYEboVPV/MiAjOo+afVtC8BwoLR9/Mb7JAht7/p35YIHZgopvQ5YiiohjuS1eMdQNa6FYULzWw/j
79ftFQvnFaEBU2b5BvDgIfw1O1M+SW+OpN5/pijkvKOQQ4Nq6IMvs/QY44mAA6KDDfbTY7pzsEXg
fw77GwSnRdYEUV1jIn1wL5G88Yyz8RknxwmmAhMM2ijg/d/VtpQaNlKcHvgXU9kG+6yOUVtFzx0S
ajrEQH+u0Qojvo9DGR6UX6c7uxwplnle63BB5IHKx4e5VVS4n+ETGGroMdlmgg8UKxUN+XoDCsYt
CMZcM5x8mn5Iz6k96FvZU66mG1psM88Y1BUqtPIAj9vrlAss92dI5OYnK8FR5zYVkAaKSkB7LpKJ
tgmghX7hnYp2st6SqRjaT/o/WSirNsViPtnALG4AKVpY2nRxmM12lOTfBtJmpqXuXDOlRrw1naeK
xwazDdz9Cf4n+fXsAJICGLYv7wO4wnudrX3uGtJWQgZqDIrWYDKVnPeflAD0+JX1A8ZDo+ec5i39
TQCbHQPzT4paNsUb50bQg4C5fZZaAQJA3wWBnVp8cFLaeaqdeq3koRs7/7bVy2CGVkBLNO7PyV8m
IxN2lQAoSMZNotSQKIMBkA0xCr59eFgLlnU/+IZT0AQhPOqZZ6KgLHQXPs0fJ6qMJHXdhwRdsSZb
vAdt1RiR8fVe5BM7LHiv1kOvx3icpRu/SDMd8yBHfMgkBe/aTuPjIw9zD+M+NmRYm6MYWy1U3qKL
DddqmIvETEYfeQkqz38IyCTdfbIOJ5d5QQOEpgpb976lX+Y38/LfLHocefsaUq1b6gV3XtDZs194
rDYerrxFMDfyIWZJ3wdIitv0cpYV8h7LvJzjVa45/Yo6dZ0DTsd6chF9G+iaMZTCCPDR1P0SQpwg
dbWkCTGsofoUbTcHZCVn5d/TjKh0l2CH6bc/WHz0VxCpO28K2YZkakbEafe5EMxheX/sr/9cRWgO
rArieVbjf1w0gHBy3jT76ZFrj0XuJGTU5U/uAyX7+HJmQ48xshniaeFG10P3Aufs/cnz6j2oiAC4
MvtjLhWHmcb/BPjeALGH3c5l2vusOZEX6HB1TiPoScR90EDu7MN4m+Fhc9UCemm+LV2PVoH1lnIQ
UTKtapWctRNinlcABArk+BLwJRKZVJZdXNHHDEETKXPq8TINpm+qx3MDdkgSdipryhmJtutWFXuK
Aj9q94A4ykVc1LRo6mYVxyvMD5RJ8dbjTt0UaekIZA+xKdrO3nBChY8NjSvtvOBulY6RLTD/YrL9
hjTLOUnNRWNt577JXpkEU46ZsYlXAEX9RNy/RPNrv48nOJMC3mr5lMRJWWYigLMSQ+3TsoaA0TcE
2IrMQ27nUdvesVBU2Abnw1IzonTDeZhebp590WqeEfepqvoCloOKG88Cqe9rcUmp2DcTDRJ3ONBB
ixeHwsQAwJRuhMX7JGTQ9pH9DZvNq/IUnd2SFit+f9Ow7xu8ACQW8vmisaWEeAPgR0Hg0u4Uu1WS
GTUGu8yuxYYIsGVUeY7fNmDqA53j5FFnw8CzbmgozUoTuXA5/xhoq4IIDePS1hoPvaoElwTREqcI
LopJ9HxOzHTQNE7MZKDw2W0a677scbjd9rYfPPpCx115snBLgtmKUFexp5tYjF+ALAaOrH7LhHb5
uBFG5nZmrkFR5Usn7sx0L75cbP52QYzZmCCmS6xKMAC8NXMNYW+KuZH1Ahcnk7sRuOnqPexcMfCE
6MmJxEiEQ7YfX5mXoAFypBp+qFWDFrvymZ5lN6fsqidpMbWIlSNyg6Efuk0j+25zmh3dgZUYvQpD
gF7+GLhgDTzyZUOcKFGCaI9UEJuHGpZBfRBQ9nuwR66CaDk/P79SF4hP/6DpIyCF3rmnKyAptVa/
qNTkliPX6EnJIvKbxsroytRz15Bil/DopIwvUtE26nJEmXf0Yam3xuFzy2N6l9VryuVe2KylpWfN
mQfllP2SUT7KCNIWTbRCai9Gz14kQq7iCrqE4vOgfU1U1zvCM6tGyo/59oMvJbTRtAUgBc4VRgJh
vp/m40l8vN7luR04K2CXbd+RstFzD5wmBsPq9urHwrqaQqa3QU9RHqxO3rmKvWo6/VcdItDC218k
ZI/NXjutS1ss4T3+1r+ocIUbvLIpvNu7R43+AHwbCjobSWHq9HvHN5Of6RAveKnDCSkFqxaezPso
u2OyMmVUxl34a33QJCe/srufZ/i+zA06S4QcJXW1rR+K+2w0shNVCG6T38RJiUXWYYiOGl5byGBV
/BTFbsJtnSJj9BFqNNpTSn2ou2dXcdVBWF9qjAuAJ0rm+brGPF6HslVutsxucdWHyUTJ1iL+9B54
HHiXCTzYEq6HJ++80ehdBjjftz2JThjLdEWEZzJdb4cM0ChizpM4lYrkfK8z4IiAf/bq2mj8tJUO
qLBwNEw2PIm8xyDvS/o7OXCZHTfASjYyZ1cyQxQ0HmyEgNLkXeZBQuf9mMt0VL9XhgRxV/qQG+4X
tvq0THCuHJHYDzgkoqVarsIhrpsbZbxlTmRBcCV/4yNTVpWO3CQd9feqsvVeno9DO4TQSi/RkCmw
I6kpi05TWbaqU2tguVmsB6m4USoYb4uIDlYKhF7OactMvT4Qc9HUhpM8DHbXG5v6ksPS/GMcRDNd
US0rJzs4YpVdvzmWhK8ZQoDfazakgXs0nRLSP9BdFvEcCrec9HiGgRDNRPZSPJlvpCfC8RT8QwCv
W479cxmRs5Xkt6jMswwTQdUn17bsk06oKQdxJNiXNSIKP4ur51BoS40umGXKhDZW4SjXs6FsXDZv
mCvkWNvScmy+SqeVzepFgid4IwE7wb0N/2BqeFHwSOYVDi8HBY9PYKP7C9+DyGJzswTksjyZq1iJ
fRbeET31TnGLhmNcMdvqyzmxg0fh99OxlD2nPpkZYRvw4BuTAg/kMfo/1TIZ+/CIQ/e0oNMbwMXM
QMoe1d6QiKtV1ZPmqHwzNHMQLnSVW4udKOwmmjsHJ6nSbA9u891Z+3dyntvkr0qOhtbCafYcjSLR
o3iIq9LcVYsE/glqsjoMxOWHGxgzLUCtJ9QynZ+Wp0OJUxDx2XYL+nqBLDmmiE5+J84ueYE1QPGR
RPRNJZn26v2vSiJrcYUownmKxA+r9FpwXjlu+USfyDipsgsqgCsN0M/G4Ufq38b4enBbD7Pbx4M8
fgkC2gbUu/rB5eZ2GgNaQYxj2eqmoHK9D30KZUmqednsyi/Rx0VTL5t7PzYwoMlDm/lEEYuiMvrj
32b3VQOP5ifxrOFfxJnXXSjHv7HFnYgI9qoqkjINvqg/NI89hFH7ELg1w4Sh60dBd1OH2q5/zaeP
HNGXWSjveEX4lqWhAbpre50lI8q8jSjirpe/Dq+C8TQWNIVdmhWQ6wM7Sn1PUvpiM773+egGzDz5
NNcmCX8aWSyJ/yjQPuAitrQl9dS3kdx2dnvJ4do2GPhIEbIyknaQPXNoQtgpBJcUevbpVSey46WO
SRi24pPNfMWItdTKj0sC2mawFDkljbXJxHOvIJgJIFMftZaazxo0lAEyd9+2lelv7ksHn8j+XcMF
IM5oJ3nPKTDgpuRfRXqtur66W2uO0vI3rqpF6Ukqkc3Dh5AM2G4VzNSD7OAMaw6W7+nQaepEBl83
SvzO7ieMOVxJG0t8zcLWoHNoSzqgpDFPUoDD93+eyym2+cZqv1uiIgy/xn9d2GSPQfw2FG9O5xtQ
MknEJu2RQX7IoE62uP1SwDbij3q2nfOUd50+wFG/GSFkVk2l6aL69pwtGuE9/9nqN4u2GMo2gKEC
fUGL5gH+rx/S+cXk46HyQxabl2woHkXjsBIwhHZtoXm6pm7pV+FNsQVjkYFRniVct9jg6fe7DBaV
kezJTj2/KHKjKTuxssdRiJ412eGzpskVv5CywdCZI4IoedRpknzV1k8R1cFZdNAg1zIJ/kjFEOzy
bGT7Asl0Pd2jqO1CaigYtkxezZ/uXCo0qho4lJuES/YO2esr+q508x+45sMz6CSEAj3FkbWNxTrt
Qey7SVCwIKV54VPs3/+0nRTw2mOrLZl79A3uqfxiqiRFwCSCZ+Mrz1vxgbnMj7nYg5arXXfrnTD8
wQS2d4XYZZAxADNpLP3I8JELlfSU/1UlvCHGmPanYniyBU2easfhj7jWYJz8am04ZvB5CeM+UcMg
cu0Y+8J+F5YC7iuA6DaXbl3T+p5+/fzjId74YUwouPmSDhySUz0eOXuWHS1KivOxZ/jqN5IS+3yA
nSOX8iOw8+7+LqfHVhsy7121j7C9HvpgvfP/sSQvtHj6okxOM4ohjtLrC5xheXGN84X+ybN6Dynr
HWqtxc1N9823893pnU0ZdbkcSyOl2YZS4Eq29ruPpjvBEqJ8cATq0YFIuUpOmMm5m8umuDR0IJ7g
mMjOosiTf/pRwm0SpDDVpZcSAXiNXL2VlURcodmsYA/KeAjYm5o419c/Giqqn5kf28/B64cHtKBk
4MWaPMqLMcuYkfd9Uc63xX/NPDIZ2BG+qdaBGVEfSxliHOJIITRejQ7KUHhQCK7GFltoJn+1u1Oo
5H7hvwV39GObv4rUJAWpLne9XXasNgA+pwE1tgHgEdn9H20t22LxiOX8EYW736vqM/XlKevh6TTB
Pyx0RCLmUMjpA4dAvsEoo/E3t8/xgFh1bLyKB1pq7BKoa/R5MNczZ4uEYqbRBodav2pDrZcQBZQQ
bjPJpjqEWQlbzu0CaoXG1PV7L7Ye1Xjw8/ilV1Fz6Vm1tqTw7+d6jJ1XXbG8vYokz+k48Agv0JmM
URvL0c2SAIl6jJXsFpAc74x6b5Z4XVRJM4BRDmcVDoNbEBvPDwyeboHkuq2WPwhqc0Y7aKGCTZVv
XqPRVaaH4q5yi7NxiOacY5yF24Z8kliw83vAokdZH6W0GBVpdHHqCMl3zQrKv8pyq9ZE/ajOLhfU
tPz9qYmzJT5fN26pV8NqbE2mgPXAuUg7ksf32SoUmHBtLKO1UG3rZfNBxKNfPYMIb2DIcNnZ+LZm
L+np+9ZnXQfgiH7G3pcwAB39OH5uDiEuj0UNHybdahz8x6TEq5QSqeW5pv+mfODxyiSFCenWZsGs
X5LdevSluTDLEh40UqoLe+clVPC46wmUr0I0G3n5tnllOxiK8TtL+J1pS9LfM4MYZmJ+QIRQqmI6
MV3Q6KQoneHAG8cl9HsfSzZazGJ6ypX/fi4omWazR8J0MU892MLk9lum0P7f76G2+pXxb1rghPu3
nA+04+SOioDLlg8JRLmnr+uZf5cUx24vdL6rvRoAWtBbwDxly1zoq8FJhZE8+wHGntHMXhnJSYnm
4DQxGD8KZot9NIvdVoWmvSV1SCNhN3pbEkzjmhmqL59lw+kPmzMvmL+lZVR70YAmQjjWdteBrcRl
WLJJOwmrPL68C/yrWPvXzqQfN1eFz2K7lf0ZmRVcNhgQeyv+mC65ORVv7lNHt0EEIOssN8xfAuUU
QqZ1CIgv+nYwtMSOr4Oglfh+adyyiXbF+s5u1tPcJT+rTl5esehWTl9C5Ezxxhz+lV0iLgffmPQx
txz4B7gjyJd/Ao6N4zOP/pgGsi+nVmNwKBIaMmTSrPKTJOL91eZWJwNwxHxEd2L7ia74gZIqNBwF
LCimSUct7O9HfKjH3YuOnjQ2JxIx1QSoXsNWLNctaLXE1Sl7Iqz8XABPSPeVX/Pcs6Cy8MhZ+78G
7XsTw4ffpwOMr9D2Od6oHxFkRfM8mCG3yp2aPsRbpqwrGzz2TKUwNsHi36F/lrAbFtMrCrtDSxcw
d4ejTQ6fz71a4Lse+ME6fM8N8BWP4bmj6tfVgUsKmcQ5VagwFg17Tz6lN/jlaNx55l7uctfITNcG
3EgcFqZySBc30jwItev+7+Qd3/u/0OZHZETTtO7tYF9zZr9amR36mT5kmrRKmUt4c48rOmWONOV2
AOrRByzSJbGF6OkAjUCnbhb3EgVBKwp+k3wB9DTDpZlr+z5krFw8uH3HNNTHFR9Qp/TnDtd7ldxY
PaQ1YXrNaIlhLmbep0DgTaJ1Vy5Mw79+Crh9ZvR9fjxueutDu1DwLVSpM2Z3R/prWgcOSkIhGYSA
m7XzQydvassG/MX/edP1uN88jv6acAZq/j2+54IFKC+0d85rGgJalGTl1oKA/gZQ9qHaAZ7dFpDF
Pl0ujFABdlmC7I51pMR9sXFpKhyo5JqdYA1cXW6ljM1XNfWtWsTX9j8pJdAzfCvNmoEZe48X0zf7
c3kHAUCORL9zvRBe82N6VwKQEXESgr1npIeOkpGXYEQ9HzkoVbm3Q7R9MvB0ij8gTjLcu3ts8uYn
oqyTaQK909LN8SOgyq/Bz4XuEdM8ZlcehvrJ1S8PoP3rnxO3vvYODFMySOQ6FzA1LPkwmFsm+nY1
lR9+OLyam/b3hvPpsh786uvk9dxXPmheWwOdMGTo3wU/8KeWmw8Xi1Ck/e6tzNKDCztlvEz9rCsz
5ulNW3KjCoHQps3+tpH6ypnAh+9QBH4tZWpAkI6KZganXmujHtQ6HnP7XtleYmvOTuai2/Tc29BY
MX/1HSVwM4Sf/nMLLRBCP5Pl/IX11w9tTdcxhf6XpC7MtsRwerRjTu1gpHKrNYurF+4LwhkTPRk7
tb99EXg33WZ12fkWiUXjJ+lMOUfs98Qno6k3TaO1IeFYWM8h6HaQyeNAaWq6MdsW/6T25mSZi1ll
5DJAvmbJRwKeyMdwZM8B3D+ISCNseWKRul3hP90chpehkiTbpZ4Nr49akXzywjG2Tv/s/7w/XGXv
1YFyV8AhKDpbgxu0RamkyGRLTdggvB0ak3FMJpJwjBD5RKaZf0tZ/ju/ToC6eCetCwh7zEA8T0FE
e+nUORa6q701wq3lhhAkc91tWjq59aYXIklPlQ6b10hE89CVS1ZiK+8/3eLL7mlaIZ35pWRgXF8G
wOifBjSSVTSqLuALKfz14RpfqMFuCuWKm+hUcm94OcRBsV9zcvcTav89iJVfoMgMHht8JowwqSlK
kIMCt+MFGHXDMUDVeqVIz7yJfbgsPl0ACdEF3T9vnbNEie1wWrjnD0afGSBQxvqM1mgQ2P2aikgt
MDhX4yGcGMxfRsPp2OSp1wfNPsGVOUaJfg0Iw2PI687hjt+dujJf3EUP2hdhGojDp0jUsCun1lEn
Jl3P0TN9JgRCaJTsBIq29pytPuEc9yIARlnnpRG9XYygkDGzNOAi+IEHP+htjI0fVpF2qDNinlsl
tNMH74lkEAp+6G9XRAhugaO4qqiWZ/Q3BF1KmK4bWeN6A+KaC0xCCfEB//3v69cVDTHJTdrcIQz+
04aeUTeKevSYoVE/lmp9BQbTaNKQqu42AX/yfsVqvfNQQgXd5QjpWfcm4jcJomXpMFhnICy3vwMc
KbePuoqX6GQ/D4XqDdtdd5FxLfQ4FO891XkJorc9mji08jq4vyb0dkWzTj9vSOzafX5JeVPYkz8c
yDuH3gAVnZykQ7cdaTMqzTwexPgFixRMEhdD+XPxbcmKqu+yYJDS/xE/JFblf05KctARwytA8RWm
bPI5rfUbYXuJN+HYQOsGQmmQDW3Ik4Kh61CCczTnNKAFAHrkqx89Nvn6qKHoZ4C/BygppTO7d9LQ
Jb9+y793ao31afwGuH9Odmknbbh7hh/kW90VQV723DLf6W+vcb69DLkCkgl3rYLuC+65EoX8rXU9
p9QFa1F7e7VWhtnpRyHjRywmXbH/xVwCtD954GN/AFSvE4DLUINmJxyTiXOK6WbXO2iLRJrLX3lA
pL4M/EqY66i3mzJJLhst9ZOuCQYfnQfdcGLQzXdf/YhZHUuxjwi6Jq2gl+KUds/f+w61AJ8Il2vB
lvHh1Ow+LaV3H8aOAX01EbnlFa+HbSyj9/mLled4vIN5opD7t8oR5SjO5nHCtT4UaKglbmZry4ec
UCuxwYyLSWXVW8+tRGSNVtb7jcSTl1be7c0DBxsJgQ3Q8xR5yrG5LSGwq4gFPqQvE5brCNI+qHXq
McmRceqzdJpCmr61VygonmvIE3Mz+1Ync0XHSslYlc6viXn50BC34wtiLQpPIbC3TZIdKtu/ARWe
vlZP4Xeob1XgbkS2x3yViTh6vPFE6iIk88dKW14IyEbVxX5OaF3x7uI0zFS6cOZCkXX1UragDNjB
QmqYpRZSh6LUAO9aX7aUGy5SH3AZ1ySe6VNb0F+eXAgkcKLbxs0JnK56AAaKrwddw8RYZf7C09pR
xrRVt0zjnvWCtPi/ECoaXcks9fLvlY5cX1wvvNrzKxYxkyIR6A0IdI93W9MFaWBiyHPPk0SczWHG
DhYKqDrBO/MsRVQrZSHdTuaTvG2XOCf2YphTLP3vFyLYtMzfpsA3SJq+4VDOUhBkHSH3r/hXHynt
yDHBYzx/dVpiJv/kvmwbzx9b9o1jQH2HLuJ/+hw/sfVS9cJIoji4YD7FHJM1unPQmensL4PiJVtk
9PWpcmSHyrlJYYr/g5diy9pTfP1U248leYJ2DovBwuHhsNyjMG1h6jFi2ThGNief5fJfmVrybbUl
QcVUPzkhKa2NdIFcOs/MVmBluTCNUS3Ma6WbygvAxdZOOqGUmBX94b8ocQjvj9D/KnDJJLxj6hBc
00n/c3pmrasbvmN4biJ6100teUalCIvfi8wlOtULGsyCNL/Ec43p32MysPWNFB9xf9w5rLRAxJ2T
2S4WQ9aatA2pcnOj3uPzpDjzesxzdT/1naTc3XmxLnHz1OMJnUzFalVUO/dS7lBE6fC07gJa0CsK
vY8sENK7KGD/k9GOQgBlQhYmslx8+nvnPBl3zO6B9lVZ5eSdsQpV/gvqEQufUrfvAZv+bSccaO7n
aPi72tXSMIWXf77vVHvnpkbTaQUK5ekRU53GXr4y2axdRy1c4uoSpdGl7mCedeMWOFdKtzJtK+B5
ceNnrVCHQcVLP8x9pppV6Et9qcnoH8nIi3O62ePX80bIpuwRTX5kfyaq9SNjRil7zOTaX7Q4Ps/E
WC5HPPzRlWXHtODrOc0o3boelgqqx4K+JoRQavJ3NN0aohZNu2HZPYfUKL7hddfX5rQSqaILklHJ
DtorFq5ZBaZSCXOKjDuVLGxyVXB+FnnVzH17gfqWQSXmfVd/setcEMn0yJqkhx7mrlBJrXdiV2sb
7WD0AlaruAFVVlzOwKi7MxUdt70JhwCUF695ikv5ERbDt2cqg/pr5XOe1eudUVlC5JCQXMwg0MYR
cuBp5o+tVHO/zUuKCmTm5zv1r0E7/usX3k+BaKemj0lrp+WfO9VD0kXAroC9OkFMuWkiz4hfbDuX
XgCu3RxG+6VbWX/Nug2dgbuQMDfrgMrZNTi+pGn49GpXKXNcGsDFWIgsOxi9xUq/za4/x+d5o/XL
roT8beRmA4WIASHnQoEO6RVtTnrqpa41UVtBs/nFBSN5wt7fQtuLiV7S56tT6dXuySg2v8Dk33pM
GWjtXmnetZhi2piFUcepmMUmBR9VPMpgnUxs1jUV6K0JFYURGc9XVZWN9sh1DSVlzvo+QDPFif7c
1fVh0OSsgHwT+pESG87iqMpaAOHSy9evsFhYevMWbFd862fiaYzGoBCdmLM3iXhc+n3RaDM3uoaL
hZUnv/ekIviFX+h/NTJx/XHt6NrZZp6BjgXY1v14nwAytWIbBsY6ptEv6DSPsz6VT8EWvdNip8kq
vy5fpZslkJubJbKASoHfAKCM4Bz9MQA2mG0NiilFIT9/oL+wRgLTQWlAhCqWROiVbLUJFtiSaHj4
osUIHRTrhouZZbW69xUenmJgYl9Izuo4a4WkMrqPHWimDCOH9IHWHnNZPYaVFdHVJtY97jFV1Ujf
SchnOajmNce8YR7yjHqBBsdPUEiUTc71yTv7vGKxC0qvIqgLgKQzBKXrGYt1zQJbkhsLKhFRyjKT
MyCMsAUUUCHuiNm+XpO6ebnnd8l/EkF3BHc4KUhkD4pvfYn+hf9Vq1Ef2Egm8FE+MBuoPiu0zJ9e
3nArGAS6QKP2MfKwqcrVwjB+P3ckL4iEvRMxRzEngUTPj7xD4RC2wht96UWDV98zkSuLyWwL9bna
4nB4zeH5oSeooyW0ngXkXK+EF6eYC5vhagrOhQaMudsi+/rA+sPwaDqVcwU8ykpnv93s8h7BKhrN
FTeb+dpAzUYRYmRoM3mpTUwPvvOCBICPuy4NTAZacwnK05/mz6tVNMXgbRa1MOtfxm63K0otLceT
EIC4xA0eR2MP0KuLNw744vXmVEqc9YIJtUjMsiNk+EVBRseGRhB/sP3ltU3WSdrmqGk68tIo2NMo
+LIA6RxGCt45kmHcyQaOgZYtjUH4zWLYqJ++IT5osk4+y3HKUo+CipOIUHjQvnnX+qcwREcebB8E
LX3Dzs/zXtcA4FguajtmJaBt4GGM8zdgXccL8aLUkf70Ny5LB1B48xUjpujiNf5wKyLiTZ97NqzK
bYIpzLC4SniYEShkA3B8N9SHkP25InPQp43cAfyWZxD7nuK6ggR8gzvJltfiBNbGgBxWwa2mclo3
eF+1RIV7svJDbQITYL6MJKnJRgYe93qFi9jdD0JxlyGczvECtWnqvoDEG1WitCbOJOqapxDJkwwV
3ijwZukx240kaIXqRvBNKoBvyUxT3iB3OugD8q9ygWPWqE1aXCwg/zvFP3+5Ww47pUe05MD7LwrN
jzsuvkOzIjAkk5ytb+lO+HUxSmopgMUpkqcwCd3RxNaRF5y0XK1LbO2uos9rCyDDzemhCdQDHdkT
6OfUSL7mIzIC5zP+dsw5YA16Qm31GVV73sU9RYdmcEVoa2h6++SyPAKkLfB7d7QNmoKlNxuz9RPp
tVvztJZxdIK6P/EY3eCtmnEh/LyFSStqVSE0lDqdpo/TVuHOZDPXkTnt8hPwAwq0+5UfK7L7Y9A+
NPwo1Yf/H6E7EXPGx06Sotqbve4o7rp0EpdVW85gntTTphE4iSKafteTZNuYneQxNPg9Us3V3/3s
8iZc4+1Acqm9LzVRTakQTj9Kdl8hT0cR0YuL57jjlsO4zhpfQgwYQEoWwOzUzVqhfIUtLlSTmaDk
v2tP7NRSUJ8UoJwJhOZAT/J4EBMHsMDBsnY7E3TWnUjEacQZm/q0LTCgfBZ3xD7qUL+uuC3ElMSM
9TU+BuWANErbtPZ8ZPeM5+fmuDizWxCL6FfKt885l6uDVGcumLAxNURvcxJPxo7wrg+HmsE8nsvi
mV6WLkY+0KrQ8g0FZ8/m/U41OCXMqmP6s1enDVq/WUfks9NCdlBbUdA7QUBXMiDOX5I4+5x1nskz
IHsb8JipUmjDrFKT6nkmCeFyBKiSpuouPHcN17uvSMLwdBCNr7SkbsKtQR783jfxWAl+3m+WiTLw
/qPvnKX0vBbqQa7XMpSgFR0QOmSdPnOYM0H+AcEB+PusF+Q/jH/GpVHsDBkrYXGuB/lEP9FPGOs0
cYDEpigygU3Cf40ddj6eMNJu5XCdKUXIUJsx8wXMXsnonbzG/wJWRCtyg5qDP5Oa7f9z0DribssF
ddG74IB4Qm/bsdagwMvH9LpQTUJ7Du4eD4TIDTc9BgWjH2p74QAboalp5CaHY9NyQqhitXB71t0W
VvIdYbWnx4t1wMA5HkpuZ+0kXMK3Tq6nZzeA/0BogcnySFIZ66sTB6l2c4GTUnWEatdqRnbO4h7f
J71s2FCdQAbe93M/iHMWQPXDOTfHpZJMY4hO4DeWXMsBADAR8PflXGa11dYIdvPWXcvYgA3dVwKJ
OSYUF0+PSmV6IpBSlHVT+agSDyB+d5CyykGlbQXcXhowIUwPft+xAA6NuB/t00Gp2oyclNvkRJJ2
nPKylI00J+eWsGPsXiizAxqT2xLZwiqyQtw8h8ULthohf/tePXAkFgpkb+YsvWHs/p/1XUuyApH8
mxgXA4XbZROoZUEX4ZPj7sc0xSrDC/L9UY1pBCSuZfW6u2LfEVUKAL9bq0U5ZHZmGcm4mAwFKoDz
VpZNOaM6fYzYYXSKEcCtMJ0fVXQQg/7ZLZznsTDcvNOcf7JKNkEagZ9PRNszZoWm7mam5/VtGx9J
6p+l/wyOSmuvkyLIkOh6DsT3nNULhuMENpEJAjHolMBK6E3b8Us3ZacdbsTjyQUvmNqUmwO/BANt
OZbFsvw01RlOWbdhgqbq4yLzjlm6NHjRm9RY8pL0WQdPeKWgI+bCAtVBAq0tdZXe2sDIsNme25i4
xv3On9shZuTKIfw/ve5tbSQLEb5rDvocehI1roc85dFxe4uPUxnBsFXsdjJoI80da4+Et42m1hjW
sj+pCHmhJF8rnZwPhrOH2VfpRUboFcFfMESzRXHgiZ36rvVnCQsIfMN14y87LyFxuWiZkN0CuZ1g
ieMiUldniYaE8jg/m+TtmRjIweDbZBpRKy+8yFBIAHcM2IMw1EDr58C6Td+i5nD38/wp4al9FLJb
3AoBsTzCNKGQVZbDp/quwPuC3/Cia7uc9hFJdikJFGoT2FEpbEKUwQ5U6TAgvpaTTw+MwC7nYOn7
La5gAQdWVe1Z91Vx+mOmMFWivP755sM9NKYDmGD7Zhbo6gOxxfKHdhKKsQEpWEyOvIRlFVy2K6Mh
q4IJ3DEIBPiVpxKb5WdxYsBQfAw8ULEan7xKq1mtO2sutG7nLi9GJ+Jd7bP9GAkl+r1tba/LPsWa
Ro+1+YOXXLBjvneCuXCHv6bYSOYTNHtGDuAszKYe/Yf0KbgxRSPkxqZH8RRQfAiLpV6jNR6+w0v/
EAtjXtyz63G1SHCbc4fQ/a33VOX8QfYVhL1OcHAv5yJlEkTttaGE+Xemayu8NfN+JO32nZ64YTXf
tuW3YlDyL3rk/u1zLiixriikc7tACtzvWLzrnUxxF+vGl5u7xd6W81xBM007VGsLYq8sOzfXUhxz
4UebAO0vple4s+hiaN+QDP6s77tvUpr2ReKeaduUj0416nvdWto+pVXo1WExzIkzWUxLxAgq2Q5/
qv/Y40P7G52nQXfF0ByB61oA9cqz+wPL86KN9Xh+iw+qCG8wkVuxl7K8iPePToAIYnVxN3ihT+9K
3trK4GmMN8JlW62tgo4tpVjDfpLNh5++2xTjTZguCr1RwDC5FEv3n+AijPRgklUfvkX1FTxo0lKi
2pOYd3YH4qqK5ljn/nuSpz/oIpp7uAu/UnrMOmJaCQ9JbAXP29npgDm3L4hyK1xAFhQN59b0iZ/J
oXPQ6+NUe1QBcUjHlBBfhdmygp/XYzR8bRravS2eJEiS4WmLh40OSFSr7+iG6JMwgKcDuDaRA5cf
LREsLsIrsnV8l8YbH9RStOnx/NmpDxpA6NWlw8grY+CnIA4YP16GpLKZjmG+agxydzkkodFREEiV
ZgBK7dqP/kQ9kgJ5EGIN0tODeGRbs0GlQVvh3yvY2DdotdcUXaAVqrnNzEIe+VQCUK1un4PMia45
G9uloz8JhS2ZWwA7JYhSfQfQL3cLnre8Kc0PnLSZksZCr0VsVI76l9SvnebG8YYKej25KOx6EkvO
b9x0SCSqf1WLGuqHd4pZkcTup5+9KOlBqgKZ1ui4jmgJw1xMoxifw8j2JLYaRD0rfinn0kpvwTME
bV+1O800uXnyuAweBiipoRPpZtxWnmHzAVx+QJ7OOfed1tRsunGZY51KtM3KkRAzd9CG3Q4PweuT
QmlCt1Ru7yijxZcBaC7MvLRQtJLaZYkeP0ornaDGYRh6ZY4pT0wsvpmWeqAJMnQQU4v2W4JdJ4N/
uWb/CuRg15Qn5QAyzzL3eGF64kgpaHV5HQQsvz2B1GlAZyvtlmNjyEa2V1fQGZTAW9XnsST7xY9I
E1vUml1KqEk/1Bz5IYfZaQp817Cl0f4xuCYTEg7PAcyc10HsSybm3EcDjIlGyx2GmmY9OZ+Cv3u+
RpMPt3p1qwhNeBfK/MVwfERYI8ioCe1cCh5as1aYI5f4GOk9WtPsmC1ck5KYxziXs3vdgCpybN3I
RkMZVgoCSZ0fotQT106h9KDd9AXS+CJoWy28vGWEjy6TKbO7GrWgHSyDiWGBHkxXZQDAy/A+ovt3
C96mGMUUezJeT1ipv7C4nSZOv+GArRVkXv2jmF1W2S1wE32/lUwzt2q4+mFI518mzra3NglCDDhG
SFh5PnuMAUabPQX59SjU+x5WLUF2tZmpFhyk+bZJlSbJlNwGTeoGqFnDPBWOgWw9m9yeS69nwSGJ
vZ3bHhqrHXLWUJ+0F5CWqNFALfW5Cq4GodGc2j2pQ+WFEWEXTCXMSF0FxPSXL3orwco0BIYGFZTC
CleApxun9OmoAULm4c27+rYdT1g0bR5uZvx99UdvyIWoPg3Ne9iNy6ben1z8Pi27ELJ/cfYcdfw2
lYQzQRtjLm8ogUKVq+HFDB3kqSO6chLkWc5hb/NprXauryJUnlXr+Y+t7ZZyrIv6+hBZQPrYAh3v
3GAfHl9sPoPGfvAsWMHGDJKhGD4zB5CMsb0Na0WMjB+czCaGxyRwelG7J47JyoCxbnlAOldp5yTy
bY99CiSfiMLRu1xF3jXgspuC0Ai0G/D7z9PiqQeQMDLaWLT1F3Psy1wKaG2mdhToOmBdycJM0RhN
ttnSXgsHRrKh0+YHXE17WM3Rjht1VHVlZY0fLAmrzvjJo+lmWA/qX64w6FPI5FUaOqatLJOtvtQu
IXwgVKWZ47CzNCwEyVu7C1jg/PuTIw1pXzRjdQmQpuVbfRkTaVGOHOYuH7p+HC+LZKG9cmFnnQkZ
9ImzBizggBx2gc7xAYs1apr1ljBAmUvOUfIbHAf9CL405rNXmi74bh2XmQ/GzREl487hZmc5vD5J
PbWMfLuqSbpveMiRhyQN8wVRf79wi7jTUBaNyn80peC2/uPqQC11kaP8BrwL3lPHnspN9r9lmTcn
Qm3KlIzQfqCQWK/d5tNxk9cqiTKcBoOEOY1DY7W+XyLW+ZLoI2thJlyU8rnWPRWJlQae/t712mas
viwiJ2TIdsZCeGFSx319yoEexesiMbStfDys/TgozlQnxwW9RyvzBp/ZI2/MsP0pp/buE9MJ5Gnw
LNlod3+k1dAn9YKzU0DxRwuL/9TvOUJR8oLqW9ivaOh2FFIUdNxmRL+s1VZ9viw/k0ZRjf+O0NDh
iyAmgn2uVpChO8J7xRsjMoUxZmp4AQI9i8l+RPLMjgoFTUPJKtJKVpRY9mZ+r1jslyXOPKmviGza
zuSi5KQiJhf66ZU9W+YDtPVDWBGGS43B9jE8AlVuwGcHjykYtRpDz4nqXq3FI2VIQO3dC01lxT0j
tEzJPTsQRfM/hYs1lC7E8qcWJmYJSP+IwH2SZJXbRG6z0qQLL0fKRRlv4XtiL51/pST2uAs9TaT1
cPVpYbl1l+PGjNlGxCuDbkZUsPPu15yCb7p2NBJD2lboO0hd7KMNJSk5hFequdD+G5rDUUcAI0MJ
xtOIP18n7Ggk959ixQJ2xv6XUDujpNYYdltqZJr7X8CzkHI8VK7v4kXoa65InLTmeZnJxIvl1RRd
j8IvTaQ3j1jq8XYoe+KHJ/A4am/d7PuezdAWOrkQamaYxa9i/a+oWTWRCtqE0DOPL4J13jq/y1bA
VNdVX+x3v1EG5nf3zWJW6W0jorVKaDIWTq3nSsFJ3W2/MuRCakK2mQHtKw3Lk57b3WuT0JfsJN90
yU/MxKsgWb6Q/rN7Dn3IRRKFAqz1YFgdUAOrHgOvRWBRul7URuPzYpTtcudMU9QgRjv+/O7Qp9Ri
s84dtBNBgaatcTbGm9dvZIuCRz40GOELTyjtIeK9XbfQLdXdywanluU1RIwyc5KIWcaMoy+7oeYR
knxsBTyEbid/UkURxgC8qwDM9H2oSm806F61qW7qUGvms6Ntd3BOZ8ALfLzhYPBUreq8Nvk1LswI
h9Yutz1bpjDERGb3G9mOwDoEdIXYCJ+Ak3lMw59b8CGaDrShneB5oRF3X52VWDAtLzC7+sw5lBkf
KndnKFwgKDz2DXGibtoQoF6/MbMs4XNsmbrmGNyW2Pq0UTkibnMM+3FjYExu+Al99Uc7jXd75Fwy
M0lmk5fkLBxULqXrel0mxSxJbc2g27iLYCuqNrARqebJkI70OC4g/cKq42MLqh1OiPaFMn/JamlW
fmFD8/FgDtdvT1ag9tlLTJoP5P2mCJjPYoSclUyrAPqAHJM+ZGFFdqS9/A2p+NVi9fPBrzBmXqM8
tR6IB7SZdAMTCB3WJOX8dXFtm7+pOQZDt75pqpQ5b5ks2CJxGRPe301O4SRnZcAWGLqNxvE3TZ2k
dTSA24IxqwNNmACBKZWD3URlPqIDAlHTgG5WubVtHiyFLNM87IAvY3uswy9l4dSjqDaf7vaNBagD
qKcQH4OKLXG5UOeiJNRNRx/6tp0+FWxT5AnXKkU1NGfFC4pBrC6ODFq/mk0TTmm9jCoTVEHjjLt0
cdsKpIVaVSdJeIyhKxwyO5/NX9PFIsWbB7Y+3EEiM5zNdYlCqK+2O3KD9RygaCcFR7o4Ap9vgOoq
gmwFBGEjMPEbIG0t8GTniOQwtHPxdGS5qawlurCHc/nlNbP8fihReR0vnl9ha05PEL8Bwtru5V4/
bFdUaklYrHdUpnrnVZw3ThXuRqGlLt7iJ7jQLR18WkEsobS7/2Mq+Ej5Zdp3fD9XKtZyxhRBKzgV
7xP0P62kYR2fFoFLeuORTSFGRIgW4F6KbQ8tTkIzdO3LyNCyd5ZlFvLE37DKvAajcVILRACK6ASf
7das5Eo2bPYlJueDmBbG0Hs/xj2wNAEqeE/3R+vwxAl0TKNzS357lkkQ4XutiopMsyGIJywheXZf
OyrFgwtMVMc1bCq9ydDh/ySK/N2EtNTrltBm445GhitiXslVd7pTFZVmQ8CozFhB58NW3wV1HVDs
XIKRt4NXPTgek5qLA5WCarXKpnPDpdpLn6cAryorJiqYLijVbTyddwKqf+u3qK7dYgd5xyBH4Bkd
zFr6Rfbj9Imw/E2ORG15pM8qNhaf0ET4Can7Oe/PgepJIBLJY/fpaqHjn96hPkCsO4GXXE3yCCCn
lRMWBzDNuXE3T3wJgxlViCffirPz3ncRrDZRh2SzwXYhOyorvq6DwhhQxxk2DNo+wYr47EalpaQc
UkfZspsEdPziRtimB7fwv6MtZvPn9H3DzFcS9F2x/lDtCVyJcyEWlTyAaRnxV2DvQko45shf8uZu
TCQQllJQF0Rw0VC+9WUi5fyybA+BFJeYib/z/sCTAe5KF5FngcheSIY4OrFiAfPmhm3Y52+uQ8UL
2tvR6WR4D+Piq0nBM6rO+1x7QiZdxT/djADnnMhXEmm93ZzVPpVLlAJC7bq0bY5J5EnXA0NoRwno
H7zIGXGVI9zKBgpVU4DvT/o0vRFUfk+4mxEHbXlhgxFfGCTw7LJmMq8ajXkWK8SiZAL7af8bC6Re
1SpmYw+5U4I2ZvXG1pcBOd6qC8qRhjkKeFXKsEkvoLTJfh0SYWiJsreX3GT6fFz3S8H04asv/HT3
gNyaM1vq63xGChnCi55qVGNbFPAadgyYV9oUrOHTg09ZXzR6x5Ic7qr3x/NDxG7sDDOEfS7+pKTA
z31F03gLaYFCqqy2uy8xHUWQEjoaG1o/4fkDbTa1iXweZ08G8ecR0W/o6uYYDowAvDn9OWZcFdnK
+VBqnMMLE3nrxVQlRZtFbT5Vj9CIXk9XOdRfzjd/w+tiRH3HFwIMN/JvwA/IQoV7HJtSN+v8yPVt
WcUWcofwdz8R89jUCHv5Iauv1QeK9NACV5Qwuu9lDGxvs+b8CHDWBAzc9BgAFGjobJyDrqNq22I+
tgdkaP5By/js3IvRDmeS2Gcank5TpSIQ3nQSGa8tsXKM/5v3WYv+Y+4+N6iRRsjl4puH5j0vNe07
zQ9WH6dJzmQh2NdbMbjUYG4DETu2N4FoU34kLyaYYeozIrBNgW70E1o4LV69M1ERlhKVl+7+mpj4
9fK3lhcd2sZfvpzM0BuLRYwlCJxvYJF5zrcpe//y+lQpdxIhtSBebx/vd/2Vp1Vujz4Rb46mkgfs
LQWO/ONilay2Ix+m3JKa2ILa9Vx41+i6Ub+fEkFrmFZ37rMIJ8HIbZOccwa38aD5dThjoyGMI0n0
v8WtYN08Uzhaelutef9EghQP5qIRpEd0uqyJazyG6Nwm0w1+QC/pieYeGPe0VXGbRvGIlbVKrdIS
TN1NW+GvfWu2Z9F2+VyS026mGhH7/L1WGWHn+2roaPm1bTcF/7MgWOfATLLSJUMiscPon0v64aUv
uYZFDrFlGtHgRNYAp3ycHoghhvPmvzceCgd9Py7sEJhkV4fsOD0rVjXOdxqRnHDkLRNFahJ7YaVL
ICk69OTNKdPi20lQhWsvbRteHtDINDHGLY5Db1ZFfOhx3g2xbWfULP/BKX31eE/M1DQbgzUn40He
Rp8MfE3OQxJG5fhbZUFVLFdiYsOwT/tgbUkEEAKNAoYlM9fNkU2a1u7RueYuZU3OdqtHnDyIXMPm
zgJKTRNEfbM55n6f2D1Z42nearegjyUR05SXOccHUytr1bJn9lufDGw3VKCRM8Nr/jMrz9gOkdMv
9vngNTDY2y+BdBPsIXr48gdL2OSzG07qREdpOX5LTpdzO8Olfg7ipHvVy7LD0C/WwfzSZ4hNjc/T
CMrnzzB1wyGlyuo3xYgD/PW/WZ5ZBSrsJ3d3tIlGc56Op70XFsCRbdbvjzuwsoJd/pYRVilRPLKE
4ay3kdjro88c15d6I7RU0RFI8F/tSJMxe0gB3zLUpFqpaC8re39y5hNtiBPGOPkGt6Ya2ADUU5hF
UQxmbZSj5obDuP/p4ZbIiH/Y4aUQJIEO1W1YdjmrSWlRTxYdcmHuPJpJxLHFE95uce+8JT4hiJll
BLxuDO/0MfracH5P8byNaT4OIJIO6d6r0D7c7Mb/J0LV0wDQd70pXG6+dJ2UNgk4/YxOOIZLaF7P
M+oGoAAZJIW6UzBhrl7chBcuvkaHFWUJsjM71M3yc/kcXWR0ZSs7OHSLzGMo4+kJT6ubqzmxO8Nb
A8QSsQm04sLXyktuM1ubgVf9QpnrqZ7EkJrRwPI9orjvdEAWMsZOamNaQa100UzuQDUMwLR4lmjB
KXMlMrQ4A+Nk/nT7xw7S23Zy8yXh+Ym1oBtQvlyoseRzMt3F5bVmtrda2fLjb0Iq5FvHy0Q7En0F
oo/IJSlOI2pDjg1CTAVHY3jGZPp+U7lc2LGSohfSyW+fHNBGmb9/4ReqUiSfHSb0Kw/i5L+CU3dj
iir4pM5/73P5Pxzmh9jT/vFkzl9HbgwwY5ggI6u90i5mu3acSc3+LB0jcZAy3Yp1yU4jqgtCpzXJ
NLxWZ71NM8MHEPefB5JxPy0W9d5tXRY6fK6TBip34fK0PqLNI2ld75oG8MxW3Ju9RlWkdcGre+zL
Xi1RePNrlqRUdayFb7zqO+06G6ZToRmYxHEFHJdYYwQ47puQnog6G4QAPf23P4E0GyETy2GgKxi4
3kpfzRFfh3qRSuMFarRzUQ4d9PCBswRQDol3ceot7jl1nmXxZRdtrYw4yiSKH/ur+umQ2DHy9mf5
TebJWsViyN+NZ3ItweIScQcUQbxd89FXQ6wJe2h1ueMt/PoLnOXukjfcH/DhK+mXC/k6jbpgB+Hn
TnFm1OE4PtHQLszZIm5Db6xqORpZYINSGTPC5rSj//YxqidFUoFYQJFpvEngOVUqgNo3dBYvtXix
sE6u744G0ibt0c3XiuDnQYoyGgQZ8H0dooFmtAUcu9sbLFaxwksr73MfnVjOn2LbatbEwO7fIGj9
/FCW7U8zHA6el+FVf8AjpwNTfZZBZgnbvZdOyrQsN8PsG2ysLhkUQBDKrwp8tpzyT+YF0FkPF/Y1
1ZEQQBTqFIzJpIizJEZtbQPFr91/w/SKoFFHEjgE60xzo02WOBxC7uYb7xkKX0iow4Rg8ia+Izoi
mZTmg+JgBpjJp6fUyKb8FXHQta2sPnVnUJr0qOGo6TBYetwj7bUN+hEV74Q9J8ws+dYuQjn0iJq/
OzwlTz5AH0BpxQmZcT2zp4pmXE8wPLmRRvAv8MugKeU/MUD/5rLXGqVZwkBuioXW5KGkIuCGlw+X
kJcC6lvqY050OSH3kzaEA1jMXLPzYV3HQ9xs8isD/A7PXfVmGuC+bUShsZOAjZXoSG2NN6+5M2zd
CTV4GZdDRbIvkW++sBb3MM8M3XNluS65GSpAh4pXpgu1JHERKtQmsAEr8Rt4KhrbsYWgb5zA6GBO
RCtGt8xlr2/I6PPspXHOpf6Ay7VWQ02Z1WIa80/hu9TnME1iCe4Evw6SQjzN0mDqGtH0/dA9kMtU
jMI68bbVnkEQctFUFJnZusiP6cdhS/jCn00Gy4/QLjBmS44HEtkw9DBFwUR/1gWE0s01tA11hli6
2uylr53IUGDyZ28xm1oC+qI7ML08sN2Sdjj4xkjVYbSX9alstpjtr1tj7Cj1i1OxfXKylauI1mDu
ylpYbHtIMl+gZStlV5LvdlKfo3pDL0RzM+lEEDoKTc34K0k4WqtJN5uIg5B3dgIcTIVMxitOzdAP
q/5m9Ikd5UzCI0Ufqjqm+TsOSwzN4A4oMmMboONjx52RFABd9xppmF8hpu/trImZyhIhVB4vTr9/
HM3/9+uM7NwEJXGt2Z63+uB+hB2Du7gvOBDKPUvFraXvdNVbFSdWEkx5GaZsrlPzab8UIYp5iulk
iv30RCs5sxLmFvwb4BMD4UfPqWRtRwf4VTotFQfAB6d9nfjuOiM/VjBSmv1w/aRPPzl6ntKBb/os
YqE8GFPcYjBXmI0N9Obb63SJ2uNeHZQxvdT1do2/x0jQj3CujI26A8ITgq0A90a2dsuF8AN2o9G5
nVjVeKjPf149lOo1JVxEpCla8mrtG2wUo3oWbycsDGQhAaoKG6WGXcuizHVb17Z6u2JR4QDuvJDH
kxKR61pt8re57+eaGzJ+pwzYEzpaoe7VCtmoDFEGHPpgiLlbJlR6GqSlOqxVVvHYUSzLrNCoxfbc
Lo9rVNUwRmmvXXNi0MVlpW5Tq/pkVsKVWYOy2C1A/yeOBAA2exUs4tNrWizGrZPtTuq+y00s8Yw4
8jVHda/xcUEy3w6NV4poV2DTjZLqhaFoWFTzd0yuCO84UX55Bmq3Ba7XMoWmN37/hlLbrIH83B4M
5f2TB1EqQSUP/pvhRCxH7t9qbqH2VJWeGSMtqPFhtZrIxkEs6you5ppYUzPj8gfrFyqvWD6GayMD
P+aCYrW8nVu2wjUofQfmb2eKpNhQFiNTj1EK8N967Ka6suchF+EKycKDZy3jsceGuSNOO3q3Aevl
bIMegnz+LKA06mb36Omsz08dkYOr8s53AV+gxDJCEJn3zIdpMFf5xBkdMbx+EfWOzJHY9KaKtRKp
6/CYva0PHw2JYJeVwQZp7+F783KSI2UMCa1VkxbCdhAG6yrTIJciCi288/BKO5HrZgcucHqdY7MK
hQAg6l5/cq2yLoUkvOj+B+tR0ocJI77Ve7ifLy4kHRpRwTG47TYoMsPnOkGEurThGS0Ol4R5zVXk
FF+spiODtBakxD6Y2yZpCpWHspDtTNAvbrl0hkAdcZ1BUuCUaGD0+OoH18Uq92tv+RmhaLVj4g0F
2u+YNlbWm1+f/3hr1nrAt11M8lZi2Gj9kEdQiPhwrK5jq5+C4wkraUm+hEIDskGkxGR8esK9l40h
LSsxZKWN8HHkAigbjhbn2XHHzcihoscRZoTfACFHFM/SPxeo4conhBvTYRZw5ICNoVutuXzZfTrP
4I14cQOgAPxSLzjH3Om0kFLDsLUDSg0YCBLT90iWG0s7xCmrn0cZBl4H8/m+IV331NR2CuQwE/sa
WJBGGIGNnnN1Q0CwnWiIpSYjKvwJunS8zXAE9CWmwUJDF9powHrkOf8/LC/o2mAd0/nu5VxRX24b
vhUQyfAStK71a+GyZXWQg2NDzksWh+F1CIXTK6DxoLGTpAsyQEuyE4G3+G/SWovEFwY9EN8ctRyi
knKt4MBSn0D83bO48VOLRWGGtqMASallGk5K5NH+b681Bkd3kLdleNFqPMgVKgtIJYI9qkXXXpFM
Gx/x2P5A3bIH5CMWajqpjZg2PGYPSnx680MzccvYUrYOlDe5iNftvOs+W3lJYGgMhVO9LDUcvXKG
bwv7FmCFZHn5rt4T5akL1LsxV7L09SAGFJXmiayRc0J0sZ3owDvXvjE06n8uIwLi9BsygCurb8oM
me+n01CTWaXIhU2Cdh8kzeAqYPDj4JF0jYc539x7RsIQhdT1GyljAEdZpZ0Qd3Qg4+gofQOoyCsY
GEeejpqSvwO/+xJauz1/33KYnIMSXs936veLbrMX7rivv1C4M0wec4Ye9ssCO0I6WBXJEjHy+OoG
uqUblqNCko6Mk6EK4Obes2mPwm4Qg9ZEQ7LC8Lj9H/OUqlQuWaaHS8/brGeDrHj5594YlADket9p
8p4MghDq9eHz+FZYc9evzBYPXyk6Wwv8aJZixLee6wuR6tzPyIEOSo2o5yapCOX8nYQ7ohpI5wb5
Q7a4ISUIN67VcFG7wIaxFgcbndvZ0B52YbkjR8WS+vnm3aKtGmB7SD+kWhYFlzhmixZSVziAbUGg
jAZ2IgniZx8MQamWWf70Q7jC1ytb9pf0L/JfVjyaPzkVdd4lPIxJEbPKm7mK0WQB2qt3aX4whetE
g6AzjDFzfPx66It1FdmSiVPHQHWKhGKIbonlb+nLqipnykpF5NoXIcEXzqnHIaq3fChVgTCJDa5g
Qc+Mml3tOVjQ5ePb7EWP7sosfJUWR7O49ujmsIR9c1LvC1IH+3+JwsigGWjn33ROfbwFyuQNHZYN
oVsv9MTAs7y9kLQys9vzCY1rDuGoc/zUEv2OlTmdjemfmurpDWeWX0LhoT5X0KLEhBx/57PSvHRX
5Pp1zQu3PgS/LayOLcIQ7ay/F7ud237OMmBYERE7VjtZTylcltz2MdtOQkZbVqpX2MfSzx6sFqFs
h3PQBYerOJqwkPaCVK9kDeV+Tp+hZub0JqJDHzWvjtNVmsrjlFAck665v2R//5/JGbuvWEGwDY9G
JPCtVhO21rQOm129QNHAfSVL4XKgP4sSrX0qTTiqMppuV+kWdYisbBnYZh69+yTCeGNG3UoGbfjs
5ddkLgDlYJsVQdJUId3qNBLFttuPfWe/k4OI/ROhOJhVXATaia0v3e/FbkXYFo6EYHgjHtSrNZWC
6b5jt3asl6zHrz2EShDBqw1gi0LkrZ3g1cx5zAZjFrRFkkKCr887cNEMPYKUeT/rWKxinIQAy9sF
uFbkvlehU+No0t9/95d/vvrucvMjpVSXyzcGVYzZEaZCj0tMBzhZCqeWhVZba40/+Bo95PJ2HlFG
kuywqMZXsFvqcBbRup7w8Gs3/42u5vmfXLLQ0IspJ7EfaQiz5XlynHlKoM1Qfe7LGQTvvmIqv0Rp
Hvk/6SYVyo63G4blDov8YxZDFECV1rikk4WxffsKCnM9VP2zjltG2HLMzu4DLw6yIxjPOeNdPdyK
S9KRIZLNU1Xct/0oCXGV/5/SW96X876Ckx3QQoHgVVriGV7LLPzYWRSoNfd+QyzCE9qI5JwYq6cl
Uw1HOZOCJLw8cXIdabAyD2tsZHkrHVYjjCv+GNLAGbFweSjpPxo3N83bknmYFtW+p2roNK8ig03S
0wOzJJHQY/7vZgQeoNqtQxLMD3ftHE7bninLTyJXdche1ikL4vMVwh1G5gM+XpPoXqZe8/NCyTEJ
D+c7/pr+hgsFIoR/gvtNBU1Apor9IEmPOQewEjFtVs2Tglub3o68ot0BTHGVgi0IADBXfyJepPE3
gPGoq1KqYDJgWu+6dEHaKGSCfZCPDRuXClUQn7IOgRnZgp4RqjU4kxJRuNc0i+0FR9TpKcvXXl4i
EuxEZAdzxWkRmRRPqeTz4FhxCr6PG0FFwMNcKPayKkgHRDctnRhvQgi7ey6MqVXnjsqp1dcLdV2H
TSn+zP9AdvE5xU0iXNcbped6SvkOLUm+8u2G0pw9M09tbckouWqS5zlHvuA7+M5+Ef5RgUVrQtrJ
MRZQv5tJ7giP0LeRxXe3dJt9e1PmuzM1dzMArpNwrJ1FXB9wEdvo7TuBklqIFg5Df9gG7sAb9mxd
tvqtBA03ZrNcFCpmpXqo5f//d0P0wLjQ7neoxHT0dNhnMwToRLyVmlhRL2NeP29FzHey4BSgoY1I
dfNBlkRWk0b9Kng21cYZD+fl7zsuEXiQNzSk5ra93z0TalIjMy6vJ6NJSe+NGJbOEhh/k8SpuuaF
jvVqcQ3nCwokRCDmXtaznsk5szP/ndBJL0doVVdgAXrig9retD2YXae2eltD5GwEd7bM2nNfmkxY
yf8pG0mSkc9dd/GrEKOlmgIM/GDJgYtFIynfWglunvDKdijgyzpvCVNIzpoBdqY0q1WJH7F4rweZ
ohEq/DOot2biuTJSqLyc8KUVaCrTXD2ynTQyHWQIBCpK0z78BAP3WFOghzoXK+La4l9is+dSdDrv
ihvRPwH8i8bA57Zn2fxALmUjq74VUsrxeu06fwx3eVgKgAquHTdgaVSzKqJXCdllYLMKcxyiGUmk
syALHBNtdoQ0SvuGOXJ02wVezdTjm/95zgw8lkSz1EaNsuVuhCyCia2AA7IhFppbdM5mJtQUtdPi
SaklvP4zX8JvxX6Ym3z9/s+lS4h1tBYwXxsFMTOMzPz/5UdUP+U20/0WNNegKGYtb6VhRbRaa7qG
hWvFhPX+0DSAc6hS3JZq5s5lLdJeLA+67CUvCcAJnvC/DjjFppeudKDHbaYwNpTwrfSaFzZv4wcA
xGGxGIhEEe2S77Y34Ey1v32lcrUdbp40q1a5UdLx81jBaiQHk6pTl4/8mh7l4ieoLyLQoxPF+7+L
TrF0ZzfGsEZOm7d5AGqb00PaDTMuFUM2gwnI3J1fZgPOid1A6uMAQsmYL0dtp6IgqRQr4W+j+ft+
upscTKDcPfd004Yo5if70Pb2e4Q4koogoP+8eGZVN9hyapQwcQ14uXlk7WSl+pokXAkOTfqNiJ2K
Qdj5ALd4wAcgboysYNs/XZWlah/21iVL70hYUW0AOsLHPHsgzWP56g18KD956s50+Im7lG8vbMrh
8+dcP+CpETCWVkDN0XmLo9BwmhoyKH+KzCC4ZkBR34FYfrQxryR2mrsfJ00qhqx2kg/oSDiK8jI8
cRSpi2rMB6zqBw0nz0rdWzCmpXC5c2sdyMurdkIm1TyJK/h+25sTkIUVQHuXCwQnLpP9TZJaDnkz
kbYlwamDG3BSU3D3/Zcn3x28WRfg6445uF1IPqxQ2Q6Jz7Qu6MSTUmZh+FsJzhm4yN+GZc4cRT72
3iZp0bBQabkp0IF3G1e2zR5kOgEx6mnzrqBxWR2ZXB9Wo9y/wVQDjGsq2+cQWAaUAH0BQGYy8wgF
MoCIJTOvWGBx4d6jzLRw3LIkQrPfT4TT3chgoSeG1Gm/lrIUgA9Mirxh0uEwMMFPZXYgvd6rpkJj
cZQ6Ivl/rVKC5zFA59tHRDXXHYNOg9AVbs0x4JB5zuNnadj6sNn2MAqn8z6cXhisKadrCQHTagWJ
z4gEP7PwQiLs9SOeYb6ZamHYqoJ+dR5Zj6IOdg4cl2PN5VMOyt9V9OFJr52KYXHpCRq+vDFvKFGW
Ay2YH8RFKurZ6ISWubPOAYLCgrfDi6yzLF97dKZ5BW5ve5Lyu7iEAlaQjk9nB6+s0BBJi3hOyfFg
1YGwmxm0GLDsuVhgYXPBL6glRyHJPgcAIImqkLNfsxd8mx8RrsfD7V45blqyNnbwWaWJTyDNx4OH
AgvcKXy+tzPdhBl6LPpH8XSfxFLH60CIaoqruZxHGE7nR5humStg5lalieyTypLrB3zoSbmzlZcf
DtuDTcgwj2LHklOio+x4+6bHQ/NDOVdoUoG70Nk/3fFUJxBw+Wq56Vs+Jto5ycqSh1UsqKb/+YUW
QyiilxLDrwypFAO90fdIYJHumaEuSfPcmaujLUaxnm3fyOj3DNqE1MrFgVXvXm+K09Jrh1q5S1wp
IPv7x5oICZyGIJ42MP5r6jzakayQXrAQGXD1NN1idXkQujrazjhsxK/MVlDIctODvCT13Da8myuH
t/4rI1TDwgXDPvZvyZIEzBj+uCc3wdwrBdvGQn/je5ICN/OxOvE0Wdzj7aRYtL0+o+Fxice4e/zG
gIyAfyjp92gybq5jxXHvs1fRjzxTaHyauoMBMUt4zHYMXEWyukSh6QdHyg3MQNO3TkHBQCoqtLHL
d0OPCnrAfTxoT2ZkQrfJMl8xKPWrhrLlcOsqdWuXxkkCzjsCk0T7LcZDL6U6wVwNaVL4cUzi0+nU
2l0Yw0Ao26QtiF8KSQUQGIB+FWXSMcR3mVVwufNZHz0cL/U0hhy428bUU2XJ0EEe+Gdii2zFHfja
SgqyS5xjsUpaOhJ9NfWzuT7/xakMmO5YSHnB9NlQjeq8y5g1FR0znHgbgyfifN6+v7tbI3awCFOp
7t6aolMWkqYNw+aP5VJE4LD6/l6oFGUtHg/k9QvDtZNoYANc++pOqCzsp0ZrzbBISxIHHPvscYdp
g4tHNbFQosj8yAnLIL+M33uRyMQZB7Oxl/nJWp+roppYsGGvptjE6bNr8e98NDIdMIH0joxEfN/b
dOd5rS40i720hRqPalLcentyyJ1yStS9ksUkIOOgrBRaJ+rLNnAtG6ALzIwpTiudTURM3EyN/1ae
wgVXZ+ZCX5WSmIbL4lhfIiPSEFMs79UTLTVnXk1rYbKsdYyQwimHhwp4tDofm6t09CaaODOHANjK
3jzmAS9BZJYmctkcpCihZaK4eu3lr2EY5ohtCPSw7NHxGLVrwNjBlq5HOEU+4IDkFMfltDug55Ea
1AYsLP0pJChNrn/AsBlyWsUvzM/4FJcs3MT9efPdpkZPyuvPV8a+Ny3mTvUf/7Uc1ALRZO5fw5fh
lkEPNIVP0nuVX4np5qg8/nPTV9yEPOg3NNr5zzT+dJ5zNHjw4kkg86HeyuUuqj/GUy/GwuLP5SnS
AdX7GuDfcwx+oEP6P98kAWoHwk3hzIg3NThgQ+kDrdQuIBK7vc5Gzhp2CpXxKnWmuHfzBSW6Zf9h
4sdg4+J1acBMWAkAShHBwfMg65j+EvX2Byc1CjFcU38dHPr7or5mhoAq2nwueItf1Nzh262vXWHe
HyywwlVRR/kJYvmV5FhgAObHOAHAOlS46NZkBaw4GOKxQKwN1EyVhpGLY+p9FGH6BOxuLSnR4K/n
knezUyABbMvZvvS/5to+OxdUIPDqu+DAxjipVZs9I4L31pDb6D4WmgghO3VsLe7gES8QDaQGszoI
EEc/lo6E8Wf5IVlohrN5K95KuqBMw4dlxweeJLu+Xvkb0jTBzJq5vVWLwjy+AP9Xy0iU5eavvoJ0
eVlD4kJOWN/RLdBXi+lcSn1E9Z9RHYesBZq35Le6JBLjDNPF45yP4jJvp5jiHWQWk+3cZotMc0H6
latbhI+/YVXF0LXs7HJhvQ8I7+gwZ7uPtf6kaMGKHNtyU1KUlr8sufqS98d3uo8612CUsWrshLpA
SIASdDsztT8H1XCLy6dCxt+cnYnI/dhLevNLq0HvAAHErYXC+YV1UP9tzV6URbLW3qYQ4VxsjkdQ
sn/AU33CPcpajOpM6fxUKZ7M3pR1uU7HxeDCzA9h/hQc5i9hGrsDTVy2wlGBX50FKQGex+1guC5w
Nwm4pTXWwewqUqSnoRsgLCKJxnJ/ueQO+/RctXAwoFhKxblrhPkXXmuf/gy4LhArbNFoS/vLDwpJ
FQBZ32/TunxfSFc6bSquw49PxqZ8bSCGyXB2WYzHZC+Jv49Q+xA0jkU5AFYGroLMOJmsDUCOkZvX
alyOAkcM4RoI80L+NtbGSrY1qOM+qOxGdF6GfaLlokxIZezWDrRYp4/+6uAl8wEBQQb+RPfyZPkx
yU7fybdF6GfqGStbdYWPKwcuMsqVdta12del61+S0DFcvVWPqIDf6o2amt61IA92eBEYXp2rHIiA
2+yzIl2xdRPp1Q3RRaL71W6AAUai1i1DQCcyLbHPKvdWz3SsTC2/1/wwuNLxoMPK4gkj1eDjVwUa
p8mGpFAEplpbWz8HjGFaXLGNS9bC1f65nGElMfyxx2YWsi5sUXF4KMZnYGL5VqMoccoxnmBL+pE5
00dCqyLEkda6bCeIH7xK2zhiS5Nq0y0w93pXG2APi/CHElrdHlHDl1g+wjZy9LGDM3BJg/na0aP/
6VFyUIoQkTUBfbyo8IuqvwxqX20jbGuagiXvHsmV2Xz6pCjxhve2N8SFYIYcx3YNz5s8gLe04yI2
KdMOWZ1kkhSuSKyRy14DxLQkFDgcdV6s5NqStaPVct7iGCDgrRbMBCKg8sIXZcNbcV1/ZKyUsS1Q
SphENAl40j/k7ORt3HjrfMsl5RwxET7MgxriO2OndEF3xJIqh8V0qLNwqcMi8wJiB8/582i9EVgR
j2E8o5daAnOGEslo986QoD1wOOicLlSicxUQCVt7ME5zOUMhi42P8QTMXwfsbSgW81bsSqEEhCPK
LsmGNfBNON635dVhWx3kVHGhe7ksKnJXVNzCJKqaHapmwCrLcc8K+EAihpHHIb6LupZEGzx6VCCV
MuDqmXTyS5LgMeQq4M2nJR49ctO9TYR8llGtHh2t4aueu6WZUuce2FDwLfpuM0TM/5+ttIfxlnKq
lFCyAgPl9HeUTtq9mqYazCvwDaQJWJpuTDCdn9RdOgOwT/bh2vLAZ9Mw6FXaT5wFudnOYSuL7rMo
fMuO13rZeLUb5DytmAk0aE6ORNozF4CloS/VW28gs4r7/ozWw1o65DuBy5EVkaMza9FqKLCEnZv3
2eI9CBAEErhtyUoke1Djc/yGIg7K7aUdS3tGPpabIjgGLxwPF1EDhZxmygoUJAnPvq1urY6iW5g7
PKFIhLIb4vgl/nGTfm8z2QP721gSXK6g40d+O10qNFZi9xa5BAE9JGNrUNlgIDNe1Bi/pfoOsobn
W+04M4M9gBBI74ZE2Mf6+A4KKQTIG3A72WscEqOVr+lSU/Dd7O/K9LqIgZX0JV4ftuEEZkeh73sP
TBC4wH7OsAi4+TUMAs9escAcClD9WOFojFbr4uzhQf7NY2WZM/xqSdg4mnXK7wfNs3lyEEbmulYC
CwTgD3ZOkztfnuqCDzrSzvBQ3wh9SuONnNWz0JL+WFl0pBN1r4B3i2r3DS/gB63r6cYkRe7Q2meb
0WXUCv7LpYo8DGpxVj76aHQPSBVQ7zeR7GZasii3Sx7plu8q0Q9sdXamnoTTi3A7z4wBbdZPBBsP
DyjCnAC5OAnoMUkLZlIMEUuX/Y422oQZJ5bERy7W/GLjLjSFpoclPc49skFy+chr63JvfxM0gh4L
CJy9q3A40JnzMOokeAwii1xK09o98wssLmORi5jGHkaC68K6Wi6GPrAnyNlLSOEXyom76j23Tdg6
ToQG4BRdfVXG5XXs5VqzZo/83gKBwLfwHZ3FoaKW32+bVy/vqj8kT2KFzTny/hkAHKJvDYE40eU8
xrYyAGI+7JocP8WUb76H13F+RvnQhEnLeJwF8erTGct73ul3tn2sMHqaJhiEMrznkRvj5Vg9zykm
QyvtolYBd28EgRypIndGMponJl3bThW9rFCbcmIaEq9Y8cv09AgN0EMZ5gfDJ5RxJWS5DFwUfgfZ
zFcpeFosOA/oitAcPGS8pOj7CKNPGoVV3d0olZRdPT7ITxYbDE9oNbyDNAAwlxUnKHdSnZF59DVM
h1lasmy32HW1+GbQ4dr1yQncgMC3DSPO1wjpnYLUh3bkC2axyqwpCrsy0CymsBiFFTYx80CH4ibF
iW/HXVxorn+JtUHA0bYqycl5gNMnfyxip78fQVGpt2B/4uOF8WjVWucybiBNQajzjTlfTB1FcxGq
hKw7F8f/6tboXnWjm0k/oPBCasgaulCdbXe89EwDePNcybxRLJUIhFpkE9/9QlqgylJbhHnvethG
D9yIhcst7QFasIM78OhzlfmO6uhas1dvY0oPX0ddykGTQkiQVqAZigOeKNpI5JsFrYMY8VygHE/n
DDTaT7ctqyXXVohNrOHDA0l8TTr9LBhfXaEGcoe0Fupx94CeV3VnuWjUkDNE0ik8w4yxMo78S9R7
tDTJEXzo96+JYM3Tl4GqW2G7zMnGDpw1b+cYqB/+aut2iwVQmvUTCyGfnxmd8BFJS+RiZ2Bt6uU5
NHpuQ5KNPoukGL5P3zJm1wZqO/Y5g4zLevG3jPdyfUulsrsElZzZ3Cx3a22J9ygjU/BOpW5zOvKk
HlnfGHl00JKIz0MOLThWk7862l/4l5yMc0B5Cqfsj6wUN3Nhvu1nJD+YCp309OwHoeLh6JSbiNEu
NpY4X6ZrnLGPU1+mpzFng+VbjqtMgGXVZbGkV7mokiWLXqyqP1xAOhmvqF2OfHHe0lZvb4jqk+2t
Y5lcptujv3rVI4LvdrE4VgFDsF+d26ppP9MO882GtBZO8h2OEI/S9iCoZPCt8mq/vIVgFYkjWAaL
55MK7Z/lDGpM8Vh04cZ8NduvoUKGjp5vsAjrw2T4az7KL1PIVN4BCtmnou/9/1SfrDi/HYZGITaT
nsPN4+iCNZeL9bfc7Q0nNxppcARBQhxq8CQEigZCYCohnHPXrWDF/jtLuJH5DcYK0vVJPFoS1JPF
Qse1d6P5ZkGZ4zG9xmJVTGZww6nddtQTMQOYz52HHWyMUOLGwt8u5aBzstDCV3rnwKJ13JHpTESx
+dacIC9j29qett7sRGoQ7i9yWKgUFFc9OMTDMPvrmec7x7gdMgvQAfofPXKOIUit4O04ef4DDpoz
pVBLJ0l43WiAKLFfLievVyKVKdUIK4Jli9xIEapWMlUZgQDXqdT3xQd0VYCL+mtBpSzBth1p2vqU
oFio/aoIYIA2p0lq4q35pyBJJhLGwtZgSB56JPxZ23z8pmI53HvVGRU36fTmkXwPqgEp6klcGb4/
p9tt7kcaf6Ssfm9vLf4MED4JGeiHACUGbYnnghvRNIrC+cE6TTphqPlKD6Qa+NKeYue+jLzB4kUg
7K/DxiWKJLHFdK+SSzf9ccr9TmxIOxCm+i1rCA8tB5joA58pdc40x18RdBPzuLFuiBSxl3o3ywJ3
Zl5ilStLA71I5olfoBffT/VaTzigomRReu7JlJI+NT8EVFUqskjRey5apUiZ0tIeiPPbQlXX9tJO
bt4KYX9NP2hNjMiY9DGnmXorvBjvW3+G/YnoYYOncbiA6Nknc92VaI6SER7Q1ed1+wqGEpj1bSQo
SNwPEzpWMzXmTyiXceAAv2Tkpu4dHf6+iOUcYS5fCpp5/soTjSbITaOEvI316Uw6kKaBKbM5uaoy
8cgZaioXpVl1FuutnDufkKm8Vyfm7IBBlLsBcgeAXGUVt97KNfMQtLNIFXO5+4ebYr+mWQkhYUnJ
yGbib0KAwtKTiTURuESkkUQu0RGihMwICIfgcfXmDe/3itfsO5Wa9SL8VrxXk/ugMKOQG2O8jyar
jHuRZvhcgu/Q5U+PipyuN54H08U8x4LOEkP8b6xMey08yXVQrTzZlOChyuUB2Sq/VYCnVASWwBOL
BNijrdUrVfqLKmWhhQJYxrijJwt0KASiFyCFkTYzwqqPNRZiVHeKoFHIMJozHa5rjZQrMYOewV2K
xZ1VBHn7COMhs/vk8wvTpkApwTHvjtJj3cxvQDBMilDGyuNe/6o+HTQlrIswK2cJg93me0MK4OmG
LeKtsHkAmkhRYjRSQILmEnF3L93OYuNt+njhBx7RcHRipQjnKz78JzcYdpPH1H+hIQXok1HGYXxS
KoZX4UeaxxH2KNeW3OtQnaBLFIxW6KWmI39wJchJDII6tW1GSWMavmI5y1Zr9hvgq349Owf1oDhL
LfzhjpxJPOrIiHvDV2MULAE5InlBjP2WEixBUlbvEpEdWIszXXG71f+gT3To/CHe8IxX4v8aZTJr
O+9QyZJPQ+qmTQx/BKXd/zHeYJYBQ3qUWPqPiSM04LYB66N8Qi+wL0vl4axgnkkaO/kns1ytWMIq
0aHDpBxB+/ZZ1qorrsbQHAu+MiwKwbD9vqMnJ8DHm38mpioMyaDxWS4peeLDwhhX+5KgyzDuivic
UrcNbSnKcZpx8mvURxH/MtadPRgbIB1VUGHcZLVtkPrW+Gp2FOJDXfzx86ebQKDqpCjiloXFuYMR
V95353GrBUv+tXJTJ3FK4DaU1VHL0tpdJoyBrQFelNCubjlbvdhcCFMYV44dz0yifrE/ncpL2gTL
T5qoC7P1JTybcbccW+R7vJnsYhq1yaGptw2+l/J0elonT/e9EvhUISZc9brIxXsyvlrtmKfaDhmy
1FwNbFNvmHr86Ec48GtBEmu7KANSMCTCWLzL88/SqScTAJkAaXoR/acxJl5OR6gyxmHO4YvrbsEs
0ZT0005zKgOlIjEuqnPC1TnqjIiEnLSUr9rCesSghlu5mJ+DVfT3z/5dPOtS0KJKKOjQXZYYmnV6
ADn+17gRknUg35Do30fcwRpdmP9023PpyaHdbM/WjS91JHA+Lwt+p8nFKkvL9IljOKPM9q/4wiMn
I20qZdtbNc1NxtLn43ZAWRn6ljZyT3h+sAZIXgTVfivkarMHy7S5nJa/V9Ug3wjzvg+31/LoJ5KB
E/hHhVUh5e+1N3CKqLl+rvNXTMzK1X80hVXysFyEqIW9WQhbbqL9xUZEzNfK1YuB66zUZo1WG4ZJ
Y70e9MG60wWQ52pmZS0aWcoXTQpEe+QYUF2i2xL+gJBohiP5GopVCzjqu0ZSerBccqCdws1RtWKB
bvqHqs9ypq0UwY2vRGLiO2RnBR5jeAl8otKUG3flBH9nyOHY+MejSOrwdpiQbfXN2MkPy59INGEJ
FKpBEWxIBj8kXe1QrnpAL6k9T08SHYOYyjQKHlHHOrmr8Sz4jwdTEdHxKRm86g69IZ2zxZp+Vebh
P9Xp+3nePKI8lmugLHOfwUSb+6eQSqh2p6mu/FwFBZiRamdbOrHTrmB7AUiUxEL+LPFqmrESbpnp
StvdXGbbdA2lz+pKZMAuPU1vJGrLIDYmgtCLv7RST3Wxn1qEWhCwlwookHbRQdBKRmEPy6JIlGNV
PrNoM3MizXa9H6G7Xvga6Yk7C/HQ9ZM1/XonI+hOdjNJIbW7HIpX5M20e5adlA42HIkF2fFV1ITE
+6Sq3V2yZ+pnsV5gVyCKie1fMqEwxYXVIcpGfNd1JYH2VSq/pYCZ5wqGeHjIBOyJ8geQjLBUpbfm
SJLKehol5wXnLmiEcE6I0IaOr7heCbV6AYsNOysgSdz67oTP1iuLEanhV3tkVGMYQvn/Vba6rRWs
T7OtNfmqXistk0N/Br0bjfGech4egJpmVpdO3z01hV/paYTMU2GDW7E1RLxFcKAOfJZ4Aw1YnOq/
shyFfvrsUMiL6UD/tz2DUu6UBoaJSQrJVJ0jBGr7O8O63ChL4bRvUeYbXG4eNmLboUKePbyxsCi/
+wf6LwaLIOqTEKzK01XT2/LdaJh/+9wqe88WJAod9xvgmh13NJHzJo8mcfhqHj3oWCJmiSeoZp6o
fQHnkJce879pbUz8NQpKUMa6ZSVc9znnRMf3etMCkqE6Z2GSnew2f/JmKj3k5jnhSqPQN7R63uYO
bDFdm0E6a0rV7RjqgTPerGSxM/z9/g5qlhBDEz+7H/GIdwtXA5s411zV5KNAD0qmXUatgUIAdEnc
XH/eetT/iVKu6LO+ri39xFjaK+kQMCFpg9EZsjjsn7jWD/KK3xleXLGe7AoIxn6KtnXp64N/fNta
nghguhfnhH53kTLyWSjFMfi93U4viBfuVa2kG/gF+vBepyp4fMiuD5wZpF37JTdIETYLBHVK0u58
KhvCgVq1cjaU7UyfzlkojHbCBTdb5q0H6m8yYNGZniZu4j4Na1fwEMAOXTteSqjxa4LbNvi4NLcp
+V/ceKXbGT08U9RZ0wvIFLt3EVRB/mAut+UZDoFIR8W/uX45UQwzhf6opU7lScRhOJ2YIfwRycTV
l19Z7SqUsDlAVkOthC8kV3xEJzRx+elTPg4MGimN9Pq1BJtBJ5xYSdd4q5/N//W9T/t/kW2TUP7T
YdzJIj4i8EwPWdbgw3JCxI59ZSWAhGS04JgPZK1xpTPI547IWgxqklpovna0BBpm4NQtxa1Icak7
oAa5nm5NzZquzF+LEF7m/ryI8gWliHLszMgJmrURgiy8uCWEku//9Z5PbutwPbBzjGzGYNmfEMhh
znT2SfdttOFAUsCTWBsHbmbY0sMpUdyg/fkKcOLRxejuEEHYULP89I8rvf/uk6LX2CoTjgZKDodf
caQeLryG7MlOGFa5PIiE01qKfoKsosngSPDws8d/ku/264vdw0Ae40tp+Je07Dj+4Q9+b43yHlUQ
Tz6jY5ik4wxpqPwB+i8TICWMFOcd3SXDZ6TnQaM5OYpJMFmOhgeoYtcbFBH+s/ADabZS4h3XD50r
r3cOoGvTFyU0rQN2TA7mT8tFvp94D5R1CEd2YLSbg5Oq6i8MfbwlUWdtQXHrUv+Mesa98Q32EY9Z
9eZTFUmo3m/EIl2ZUtmEoWBxb+4bzoo/jB9x52mGc4RMNpWpDhqNsRDIRUjb2E3Q+TzCuSsGXU9q
kHg7/oP8Ir1cshHlJm7fKApXFhcF1nu0rkANBrylxzOP0ibsBvQJwH6GF07wFALzLzw7TFNHtnOJ
NlJNtVKRVTeJ3jmEnNmZV84XIL+itbGz19rK0o1+1eTUxSUWnerjPxM4k/WwuyeXfuJJuLfPfe18
mDkn95RXnL/fM/+PJRM3HrqoRJ+eZO8MJ/vTD60yHKfOH//1X1rdxCmq+EvL6D9WAxr95PCDEIRf
uNpBAdhIEfICRj4xumltfMpVCOzID1JjLeXUH+pF1CzTjgE3+5I6YnyXhv6mccNEw6jT89VN6Ajx
Hl7i4j6e1ynZoMizyTitkvRrTHSD3XXURI4Ral19z/B5OoEfEHmqg4muAvnr+Fk+SVxSAuntA/Do
5Bb15CYOKoy5zq+UFHtNwelA9KXcXPRqCyFmwIeurGFX4c2FPQYyo84dTliKX0ps1IvnsiYNacM3
HqGrXE0KqGsaEoGNVIRqFEXWciH9mbTqi8XQQeiqDbEmQR4tvzrdq4EbwEgFyYbPaUoiwYYoMzm5
OAFL2Yl3VE7IZPmpBOAyVsgtbct0vUCEw7X/rRXP2g+A1WCutmBmvVxrfCIa49dArS00oXSnkk05
oxq4BlSP8jkT6Qp8m3T4u634DhmdE3vO/cSq8s9qGpFRsDjMn2Z++nJ1WoxCK283QZjrz0Yqa5Qd
6MJiVjmBfxV6Mt8PeLcbkY2oQQmtQY1mOOTdkgWbWdaqRABNLMm+/YkvmeBkB//f8CZzjB5MEC7/
GIJ9cdKj/L4nuvDr2el+LB/IU07hgKz9ZMa4ptVB3z1rpHTPw04dzwe+A8bjHtQ/N2g1PYvbt2ue
IR2K2HZWfcjc7UGCkDSMtAb/g9l7EQRS8uJZi1r8HcTVSp5Be5iVBpbQuSq17RCDDw4CMN6P5U/g
c5mRQxRghO6mQuLbJc4hrSkuU+WPZiz9ZqSy3U1g70SJfEKEYjz1WLBeg8phLTXybzH2XBcTSXFC
gbJdj5tlX/j4FiviKf9Et4C4JPMj59T0TCIQw52Eyw2zADpEgKPWrc3QCf6sczMxhWK6y15/yNUS
sRq1PTlfaKINvPhOUp73Lh/VGqgquToGkRp9rEh0M5xA0Vj5syqioGZLk6zXaF90oGhMSvWTz4jB
11a9EXTLPNBF3ECRskpRF9wHlKHtWFXphHhJQd57rgt2o9bMl8ePTIOytO3CBT/1kqm0dGOkLCIY
XF+uW0wyuxlN8k0v9zJBSrZLQAnafVeYqX3mndAhJ706qN6KIENh/XJHcf3zMd54vvMAsU9IW5BD
LEypOBIkZHXIzpKoX9y+XW1K9T6e3JPTmjHwr7Xrshdp1MejRAEPL7Jh6y225cJCq9r9I67SrOtO
0FUc9Dzbfz0kUQYbwbWxU2gzxbHYxELqhJ6m6cbuUrYC8C9vsmt3qEZkalSzOkDIr2vOMCQyHCvL
hNufqiqdioSxKAn/1ozgz7LnJ4Ip/w7SOelqo45HbVBQyV170jCy5ZqDuyFibf+4wFNPLtHIFq9l
WA/WBp7OvrksiPlInzQ3iiDBqj73WQlQic4kr7tgdIcllxkFlsRj03N4+v8r+VYQd4bJeY53oMlE
0N7o5hXDn39W7ZLdDwZPyUjoVIoDPNNsmh8AtgVibDc6TZV46HoHkcmu1d7j75cptRRQWxkeTFR4
KJPhJTjczuz3P0YevqeuNnL/4Mtt4wam1bkoDTy8D0s9oqJhLs5fggjKSty0f5NfEkeTHiIfKXkf
QaV90Y8LL4s18GeZB8D3/VNnnrAxX/y+dGSrqECRdeWIjpNaReWYqicY2N1pZhq+OeW25L/d9JQd
1PsMWO2+QmwTk1U0gx0odc/AafgVfn93FdbKx1zLXwxJ03O19itLZS1zi24uZHerhcWE0iEs2u7D
V38ymQYYsoSEHbfvu7l8z0QwbSsyQGQ5uZfUc7DzM6wDGTTcr3vbmO4xC6GP5B7e0hpfgFyzo6C3
ThXzyxhgpgo5pAkV4QupURaoWt7lWCfNX4XDHBYLPVyDPVNF1Vs/3Wft4Gpz0W+X+VKlLSU3IyS5
voQ/9omyUM3/9SLb/4vO/NMupFUEzncQEM9xXYWHgvYVOLC7mqyt2MdhrrUPQH6vxL4oGqt2Hm8j
+1bFCx0eB1lnFMgF9pUUb8tgRUJQUfi8Uc+e157Gc3D2i/81qC6MkKusM9MyhKNmqbwl4UlYULKd
RawmcHR4IUb+MoSobdK+rJhut4iSblXxmoKAE4XxwtSm0GOSwsfZ/p9UpnxypOBM6XPgbHExN5Ub
51cKXGO1CEzI3Dah1zsAhJ5cytQ5v5mzOTwp1TqiwGiMixmiifcHwDT8+cBkh/IIktJR9i4HRrbV
TFEgtENStwjOyHPEAKi0+WXA5BfWRyzgHybNA+21rbTup5LR1GhV1UNqwAsLMruJE9/S+7ckI9b9
pA2itnlg0Yxk/CXI+BQuOM4oLshCfBaMNkNRLX8ifntd8j0qn4GzbYa0Kbx+TOeypeGozRLmfv1b
9cGqrAA2nRKZIvp+aLusBBlU1qRUR8TCwAfvDrUjG0JllWWOK1CqdcH5M1PfEjUE/yazQG/A0otB
XQ1nrcjQARTZs4PfmJdy2I8uLH2lxb8nbaJMbcsL9/RG8ToSPjrThm5a7CaJqxwjudTu7Y0uKXT4
3dyYbiXZfJN/ONe1DWtY9NNOThQHQ45x6xXvyOtP4qlZ/9cp5UoQDG5ZbcPY6dzFE97H3JkbvMOq
FANGUy9XerCRButIyS8M2oESqgbP0UKO9Ow4xRVRiTM2bhkAMODANkvRVZ3uMVPa3pvWrhfwdgIg
3tkiiaOePNukrYoocwk+5MmatfPoBPb2hbNCc77SNNdzhr82bA4Ma9N4r/4OxZlZtFhXihQ+ATCj
6OtDde7rSwMdHBg9YTIhFDtyDzWGXScyzkGN9NdG26ZY1juQklKkVpqs/SUrS1qM+10T+htSFpVv
i8dDb95lWY5BOclZ3X8YINvo0ZuZmWwPeO3ODfHcbNTXDXitCVFPMuVikFZSwO6dJNH1m4jJSN8t
Y9iEGOuN6BtG8gRZBJd3UwnvjbBbLWV1qYMHkGxjhMTESD77cG2q8IzTylDD5+u4W1fvdyne769l
CHR17ZKeXOVpuQcYbVdkE0s5Giyiym3dFFK24me1iXPZSJmV13Y3DWisjn0p8Pzz4cpsjLVtAOKI
v0RP4VgYrcOhP5GOzXRSdgG+BmOXxnEK21tHXJpk+048Lyb+kwXgUrEQo9SD2bdeuPmOvOtqTHfA
prCkjE2BUk6p//8VPnogKWRglhXPP2C5+xU08ET01S23vJha5DkhsCLSoMSmzbpD5GgTBDL3mFOD
ggtOZdFa3APd9d/Klpl6QpEPxmfY5gs9tgw3XyfSMmIr1DHuKEkznoAWUG06+xC/R0+BpCgEeUXh
6YgLhBYE/6xNtnldvTcrkRIO46PzhKi0EQCCo0ohtJemznFntvYTnTun2Lh0QYfYSYgBzA9oxcHD
ig1ev/NSK5NCLRAM+bEMRCl0FPe56VOW/fNxtGw219MesaM8HRMGAQmwX2xP+FGlP+v9DX9N50YZ
eeBNWD6+0JstoKafPY8U51+uL+Q4Og5nIwLy6+sr/K/UgFCAlipmg6/OX37S+5Y0b1QJWisuQqdQ
sdry3sJnJRE/n+OYlpSnmR9c9u0M1Rwogrec6zkw5LSuYkX5jwK4Sb27rLADTmrIQ1ZWJuxZwX8V
7FW3M7qurINAV+pYY8M5PhukAA8Ke3PYSy1AD6Tg7gPXDak8C2N0uTa7ZMdok1Wxkd3R+SNk/tEU
JLhPvXUWI2tafeDzHxuu9CFwXtmszPOJNacYdgbg//b3kLimhz5YCJ+jcds4ochL1VOL1+QUajuL
Ivtn2wUscKIUS8bac8rAuMLNDXa1WjvGE2X8xPFKPM7k3H6mTB2B2UhSLEmW7mUtrm7u+p1FT4jf
bm5z+u7RXAHCyuKYOis8M12McgGV0p9Sp7VgA3S4QsfQQhKYxaB1tG2zmU1ecawelrdu/L/+4a1t
JefxZdec3AKtZOU85EMvjf/FgseMsZ1E+s8AgqUkJi2YAsxiqJiVpWvbfZeYtidc1KQv0bmfeY+A
P0LXARUyPbvZ6wk9xeYUvk51h/tLvFhtkTnfrs0qxXHnH1WX/S5YrDbGU9nOxZdGZxZwGaMOvJwZ
9G572bRNUOYhTVgvK4X6s8ffx8yloLjHT9euSDcZ99eH+5Hy+z4+rxl7+k5iCs932EY29Im46Uso
O/w1mpx5q3Srx4rKAlaNIl1dO7K+vqr0odEd4JNlP3UAvtVW/PGgNbbMmnSlkYnk3ZU83LtmkjQ7
9ViX/kz6IzzyBdWgZlKeNGmuU5nxRVnugVTFDZ4icvOPqu6oCRHfLtd/UDj3DVQz9QyQ4nN3O7zw
+EnoK9crtEwTNb97M+3yUU+XlJuagpttYBda5DUvYS/7eNMZu6garlYjy4ZP8KjvgbfEfo9GqxlU
lsxWkKynjJNO8XiApaaV2EkrFss2S/VDeX4UQQT9UkX3w3HxqX1v9gus9BijoSYypbzPyAxllX/Z
r2skqowghQ9/9O2pRLbswBGsaENnjiDTQzQIpNgG0iAejrH9YK1VatRCUe1hWVpvSNCUKlVpIO8F
/uZ1wV1y7TX5uKxRSPdzaw4Iip18pTzbi/oHDg/8YSRRdLDy269ZZUKS5XnPDXKz0QzTCvjzXcEi
0gay8P2opZ/0DPH3I23RncWzb82vhTWLYH7JTjaMtcOwSCKgw6QdOEAPea7FG90zxMbmMX7p1wm9
BEZF5uAkp9C40PRmVeUrODK2RFHdQupXrZOsG34Rybcr9jdVVEWGJDKbqTSqTm2nFUpHHGbtH4AH
xBES4fIxDIMzjNqjPKB4GiTTzmKWphLkSCxYLplaeerlp6yrP6aeeV9DlWKrzQi/8WPvwOK8Gr/M
aN2EEdYSiL87jQW8va7OFftWiBdg3W++gWPrfKNl2NMUxD9JWqw/lkfD9DzuI+/r9JiGIVh5Qb4T
SvFZKCc4fz0h8tBSupsvVhXUaXvQnSrA+30OAywernz5IYHIVzY8teLSOOMdxY94OHMT4XjEkG06
qAkwSz79DBn/7BQcUOkyMaPmTt1xgv+n+d/zaIYZfP3QyQyxYiwxFrQQq+4PGQ8gzX6FOX4yVA2J
c7VlT6hKRNWEANfbq30byYywIspIBHYxYL8gU60eFVvkYlQ3Ik6liXFXj/fnqblQB06zYkatLATu
FxT2qtHYHzkIbMfsl/4rZLr9b1+MiJxl0fz3qYUSpAan+hERk5gFsxF9zTdIgOTctUR/0FonPYhe
WPxwC6/uzGH4tn5MXm4H7AWTl/xbmJS70Ii09cd8XEhMVEU4fH2BTj1xWa6RwQVaMmJg3dpwa1AF
A0xd+2uXxKZJuDDxzU5LWjM7nhnNI4kgOy2RANVzwNsbVC5dWUsmcQJEMfKsNpS8v0H8Un5h5vU5
oA+aj7+ck5oygs0i5eHtMACqReuluVfuwxUIoGwZR9xhNOWcUN+9p+8sNH3teN5A4Vgy8KYFgdyZ
5PP5KDLJ6G6TWBW8Io7f1Ydt4u0z7Wz7f4xDdUJ/9Mln/iaTs2u35OOmNkc+WVCmu3Z3tastA585
FdXLKlxTJ+gJ+F9AwDdBr9lyAN4GS+VOXf5+a+Pw/JuLs+QIymjk0XfDXk686zR/Vbs0qtZVaNFZ
dvRI+hNDDmpThPLYYRLIkSjYDe64XgdfBe3qVfLuVm3G6BMXCvDn6NZw+v1MwyjyiesxdtgUT3v0
515VsRsEW6PLp8QTyZoIe/1JmRAKbE0EtzUOGyx76A0nNsHcMJY2WMpA0JJmhhpIgjGVpUmik68F
1nyTbyn/M6E8TWNHVagCBCYt4fanmhrNaTpcpwGm+emmgzzpylQ+Faziy8L0ZQLoXPcDlE7VzWt9
9K041z7CezD6UujBOnwyRanUMii5cNYBbt1TR1DoBvaV0hdtT81+EZsdPpbYPDHb2DwQN0bbxcs8
FOUsAMUQCjayV5qIjrtIwQc92cLNOlSVrtVY1Jbr4PgBlB/HlMs4+BLkTw5/ZGOpZNLG19nuwcQG
JT7lRQyKg8jX3y04ZG3/ZRLLe36XpslLKAgQ0Wrn/2iBTNFtmYi6n7v6XLhQMsnG8dqz+hNRPh5H
OKK1jmd/zK6jVGBS0m7ivT2ivSN6yL3cxLA0rEE+DqSNAyqibYjYxBtfaPgWeUvzpKP24bcQlK4m
FNSkTvJRqNi1jFHZrOcmiaqKciAyF5BWRjPNnpBlHPfz5k57/feYT5hGXJDFYOYFyZRhJZQ9Tjcb
eGkiVlC5s0/b4/YumCvZCaa76N73al9sjZpWYor+7P2qCQIJ3MI7ElfCsIalE/AYZ3Y4Flsse4mm
J+fHsZxFtSvUONxHTxZTSgoYozJMgYUdThpIIDsouzOQG6SIxVgEwt8KNOXV3SREZ8eoQ9Zbi44h
utsZMReVluuzMqBWffuZ7dJcLH+VTPrZjgkoWfZz4HJhw7CbYfgyNOAxRvMHDgQfyGVph2LnBaPS
tj8dYhRKKfNOUXnqN2t6z5SU46xNJxxF+rQ/3NNiSwuyYMn460gtZRhEFS5b9Jz2o2wdVhR+TTma
Xe24vGh9MzC0crHcYKw9M1ZlSBbZWS/vgfrd5ZR8CZD5KztJXTAqWtej5eqfXFd8IeS6s9UOSdF1
ze/al7goBsVT2uKlMkhtnHL6Mg94CKKGaXSq29y4tPKCoth9sSa1bpD1GPmtqxyIoNuZhU86n2yd
kHstidzA6AW0pOe35hVSJFhY0WA7dmvlrDdATZNbDNl5mqct+nF/UaJa2o5kJIQhmWqCw9KcNhz7
Gx3J2Coeqjw6f+Cf+PDicGQF8iY6oLch4UQD2BwIlyhQ+gjwoZK287BEnKYYWq4LLceBLntQMJVH
xgogZly34CDOV+2D4xObuUnSn+D4sZJ+0y+0rVKuJPVtmD3b0fP/WIQ1ozgy8RKicxYfxAuuojbE
zZMNc/pKkcUhzrIf9F8YOxnrmENf+bd3F8mxG2npv6Lsd1korjPL5il/NbuVdhEKq1z9rBZ/82jE
RRRb+VIqYnBhKgXFcYZUCmQux3nNzR0Dak5OiF/YsUznVj1moAx04y01dfnRvDwq+fZv0eckm0Dx
mBY7/MFsYbBqyMVQoG3uDCn+X3C3TUUiC6naBLLcCxLyVOP+qaw2mQVBVsKWLwkl35zYNWKSuM4L
yZzajzQ/W4cHv3H28u2dGXR6eNtOi3Da1wSM87VAfS09gpF47gjtH12kkciTJxVVMzT7wbNMS9E4
re24P6BAda767e/yKHtjWkTtkJcS+nPlKEVuK++CwvmblpxMizDpzXgp5zMsuq9H/iCavjHx11yz
NBOU9TiaC7ywuwJqa66arqZrYpgCijRoQGafK2dPjTSp6H9l9t6rx3xxAADDO/w9eDsazrr/6ZTG
zki+wPN93s7cj3929/ot+vSFEVFO7FLPKYc75dK9qlbn3kf2GOoY8HCL9DxdDk0z9UJQkZ+FsGIA
ljsW4I60ksae3rKBdeHYX5g8C3osc3VvnmMNnCKKbxN5JRKuF0WieVeEJeS29rf+5wFSg0rZ9IQ7
TJrJhbvBcOzf/59b4wCBcX7piQa6c7qKfs36+p2gmK71Bqw5+jKqVcHryvY6kwg6vLyADR0aeYPZ
d/WvjJcq1hsM8iyBA6vIKMNugwpdq8maYxovsioTZlFxHl5N88l9RGkABONgemuzIl9U6WtJPvFn
JmczDpfnwjJZj0Rh7lnTZ6sFoDomwORNzVe7SUQ2fU+56AfLhX/hkVLP4xC4GzLrBsuyFQnB6+62
7L7F0uFLW1R/ejoIhAzVZ9Xt10Z8B/IMEkGKzVBXInJR9ZAVnYmA0cX4xT1HNod27HaJXN+dk5NF
EQs3SFow1Iav2qr/ZcvR9EPGS5d4ZGpnsZXapej5UE+mGMCapYaTL1eJWO7GdSawvJYxfnFPdPzs
IYnrRVaPGEyEYFGNufD4s6ysGj4dUPJ1YA0T4n5uOD0ITIz6cY1Hdw6wRjcCxEgh0gHB1TkOpuqE
ordmQ5ntAB38FxDURy0KYB4ajlYjaSR0IbFWt4p/IJaADY21swQWNG41AaAbwMesSfR3G3pw2FSM
RARvxeZ8aCu04B9Bt5nKlgiNuKyVOr9m15P8R6Rnz5jj1+W+UpneHKaOR0+ZW44YAcO8YqJvbX1M
eRkZbkfiyVQOLP1AidodfySj62P/SWVFDWeFabWYvmLMWRNFAbGY343nv/n1xNViJ+A1NiYESdaK
AmESOChXtu44wWLJl5f2vfrx14bKLLaozU50lR3DFiN3OT7v7Ia3cEY9bp6IFmPwpoRetFDK9g3B
hdruCHv+6tvcbrLIzEGL687vsnR/usNZrT1aZ7EMqp4Z3YIZWbgrX7hmoLTa0faBSn3gJoE8CQVm
M/1XeBQvs48svQ8EajnQGJDI1QnbGT0bQ7Q2xnr1UVapdD6IjfxtTzTYn2gg+WGHY1Rm6mR6M3qV
vK4Slqc/ZP/fGErGx8P6lnuiN5PdTLG9QuKRJe8u+KbFK/0TOHOdjiYy0HQcwXXJtDZJ1P/fbynn
RX1zr4ZcAxo1olcXz6PUI07m5FX9fYnqKaqqRG4x9wWkhzBYLHi/34W9t/Gh/CcMRjxfbKBKNQH/
YXKp1H0I8eg4+4txuqBd2dCQMQLuLthWAw3jxqX2PmJF9Yv3OTc3ppDNFfTC3k+CXNaPE5SviRZr
QYW0HI8xcMHYfxSduNoBH7HX1HNMsP5DwtJyCEmbXNSkvR7Dg7b0/7lK8Mj+o49xfn0sYa3Iait7
6LdAWMvz3jXrScf7WiwWj4QFACsKXIYKSzCFRCWTmZmIkJSPduzW8I5bY1LbAmfbbCsZ8zNHDArW
ca20QEnq+O+H5/7f1OptIJs3RogslPlO5zEh3fLUDqFHWZcNcnHTIaFpA7QGc2uuz4sDzlSl7rUF
VZ+g4emWannU33eGfdz2mhOoTOw/tpBBDXG4OtFGg1+RvmF+VgAtdAV7hLsPpxzYgpnZixE8wQ2l
x4gmtYk54gaCA6S6c9m1H4bby5Peib/JCSZ3jPMkyaqaofOQVtnOBtk+Y3aL7qQhwoz0bcrOugcK
G+vAp5e9jYtkXXdYAsaLFkunqFWjLSi4b3yWVhWIdWVw9fbFeu1h2A04DvAcwgLFnjtp9q1VApqQ
m95iKImqvP0Hm7cSUg9BcCL17dOqzvN2PiFxlHgu37sxEOwq1KacT2uH+BOYBwzbAg6ZyXWEkuZZ
IHUgX7tvHFXFpkkwJ9KfvUTWJhCKlfX0MmfpfNTfQYzvqadJ2qJh35z3Vr38XAEYAdpwEkOIFYqv
rt48H435fdgf1vNlbd5U75BOcjpuQsuGI8g84exBneSkpHYD0IpUGPnXXGUJGh7zka/MAafty0aP
2wG0APcrbglyBY2plJz25PDKt6Th4XEFkkIXL/vyYR6OIoffaLcVPBcv7Qgo6Ior8Yej76d+rbNd
BvGZgxHqcIgVWsIWQDdSWH2y4swoV+qEkyRxmGcho+hQIbrbau8J+8lkmwlrA6Wy/pLYZYYRnzaA
6djoovXYjLuDV9bM4Sz+FRMyAGLmmwyS1ubsyjvL1j0xZfAHDaGHbo+ermdvjILQATuGONLuzTzK
72VxDj+kCNacUL3AF7FB7oZsaN4WpjdfkX6GYz3AwcF8Z9eIJnZMPM8OVV58Xk3ypllqAiQ+Sgzy
hZMmsCW+qOVKJSA8mgiwUD+Phbb/GmjqSsLvEPOT3Oh5zl3nVjoxKERCoPCCqIcd+iVCNvHhM19f
OswBJFlEJi0FSi3jauIKXcXsZ52WGUaVYs0GV9r3z54umZDKIWcSVEPNeDbn8o2nuHRgK96Rb++8
oRbUhxhK231f9duqQlv9IdzDgRNeV5isYuZBAhKPztTp8dXcGySatnnM1EVwZdPVBIQKrr4rmwaZ
aGtsKQi1RzhCK0gOxp8J6JidNgGVK0Y/CNfOvMTcORvBtSC5aqmvNZ9teagBCQRIoALmFSG3OS/i
NicEH2+gXBGzR+ODb1alYRm0jml13RfQn+2aGd773Rlp/bcVqFU6fXB9Pu8KaG0NG2EoNkkjEMsG
sumqzVjEd5zoGJhKMUsePQgkSeVdF4z83/krTH0e7bkmopTeCsvD7eGT76yFOguTMsrfBV6+MJT4
v+FJykobpySD8fWokwYrxPhXCyMmC6sNobyExvHKUU+cadBGAu8jzFHlmgiy+eJt2pl0U8LsQdMm
rrxtVMEOZpG5hXfDa/YbP+l0jMh5rcBkWPT0UurPndcIwCODl4cgtKr68rFZ7VGkA0BblDaj/rN1
22z3mb/gHFjN2DCJACq5arzIwNyDOITfWGUJWZDejWP774JyHVzWMJPnsi8aiiFdWnQxjjbObomf
22GLqWb98UbHZxp183kGO62ihjzCeIjcoK0SUIAbX8hxpxr7qSSOHLi5QjTHSc8RY8t/rNFx/X61
kbmDEoo+Ti8TELjp2E51JJCBMXu7DDlNrxVbXB6uK+VaWVOJc1EMJDCxsjWbU4DPnMQD/1q/nYvY
T2rM7vGG7hfpGACK8NdJ1mbJUG3nQpeODd0ol1j+SlwdkceTTqZOBuqKMJ3wddZZtZsTZ6R+gVZh
u1TZYNLmFl+jQWyBZNk78ViT/lLcI4uvf0eRQIn4xRPWQb39GxvlDk2dbPqrexLxZy6rVNEwt4jM
+NOxtoWkCK7Fi/srdKA2IgDQsb0cMNk8Q3Dk8eg0zur7tt0CjE3xg5yLIC+Sg51KLgfFL1kwm8V4
LTkMWKGeVgPoGclmDBJdVnYztxU/uRALAzpBvnhMygOAzpxxcus+uPWKqG9sVpq+1hpYL/V391pA
MDq/tlWGbDq8tRnIndXLLSjkvZAdQVbB0+LbXqjKvBWFbelSCuJ/13VuJIp0JvoubTYoSlAhYvvD
Y++mspL0+08BT8xjv1NEWuTUYzTpDxmpdgczwD82nMRHEwS6pRPLb5CNqzwfViMlEpyE7TgIav68
bL09plJw7CYDga3b/z3Wo4T/oCvFlivxlhuSS5yntPLujvcxOxUIl+PwH2VheQYa9LOCf1aRiee3
n2x76kpQJzxdtDC9Ut2a/6vUGIh+j2/7tRH9e/zEmhO61G22MNgmGDuUZW14eCYNVfSglkop84PD
DKxNJAnspfTLuPBFuZ5fAz+AmPxG1lnjZ6miB7JXMIa0ywF6PxAf+3n+1n6L1tJaR7h54l+K9+1n
pz6JgmXRk2Wqb15nkrpvgGuhFkk/3WmeHT3Khb5JD/eQi62e0eoI1h6pTBDonC+3myWcNt2Df4Dc
5Q9YuGgKd+x6nJ4dpr0qArd/TgIuefbuNKHGasvITaoAURJOyFOftvo4jk7Obw7Wzy213Ri+rDSu
i/h3XyIOWofmYnOy/s8lmbnVDmDnXPlrywSpHzjk8dZWA5dOLd0DAHjmrqnes7bdznq3RyiIBTI3
JbBOPbf6jm8q0JnCSPvemQ07q9rUkEXSx0G6L5ea/3atCyyIkSMPO+tPYp9a3gnoOSZuyM846TPr
s3HxJc5O7SMJbDJ3t9hc1qb+6WoiWtjwGWLMyAK71IdIHUrtnJdyBL/fW0p2/G2hjw7oLQ4i7PkQ
gsP/6M7QTvoHqowkEjYrOXWvdd9WVol4PVifET4fdBKfbiMQ8tK3P3eSBJ/gW56ZVi8QTKoMtC2V
Q8EhpuitKNyh8J5aVfpi6R63ikH5/waVA/8D9nLe94KJdysxxDfeGNPoJWZ5rsNEu6aEiaY9y3YH
qKY5WVHx7YICXxQM7VQ83HRhkz0d8Yvzdjvwcxf4/hI2C5rHlzyX7wBhdYqOzxaei6liAtEf6OFn
E0uLd0SEzp9kKOSVHAXvsbDcKyM9RbJ19zojjaXRaHvlfn1GjCv0im0KmQ8mKasz+8DmA/imqZLV
iw6YNQPsKGI94KHMgvTHWiAgS0eFb6Gk6jm1E6AaA8W+Ffl4InLlIsafMWZqEoMhm5w1b+qvFk8F
V/efjshwWXKAL3TOegMf1bceF2UC5ApTVxluhpCvGrWfjRnIAWJDZuLACOJHcBQl5LvE2BB7HUp/
lbjug6s40o9GRR/EfmlvdvcywfaoYVNbFrklUbaho1XkMTWPM+hgsd4QWJDD5gIQ0mlAJmuTUiry
KN13IJ8gRbwc9yiEgYAyDHT8YqwMwFMYnl4uctdgZMQc+aL7tYyffiYWPztW3Kx1InJDQzvh2sMK
GhjvLVCnDdE2f8pIpTVqoeAPVIpLaIcoLntrrYOsHkCsVmk7qNhXk17Bx7GS3/F5gZPwHoVxalOW
178RWE/8OZQDAHRprLCyZXpeA3Hl+Fia8EQ+VNZM5gEr8s09MxUj027NZErS0rSbEmUzmwREczgS
35Io3xFLT8p+UKykt3M6F1A/nAyaGa6UoCC7WL0L3ly0fRL4mNtAgoJ9d//sJC+skAXudvc47HOS
6fzFZR6k1ehZ/dDvwwwOM8pahnfQ1Ap34Ja3O6a7zKI3VqAHkGG67eghdTLAEthnZ5djQYo6BIvS
4QMz7PEGz5K/cJkcNdENLi7UvbG+esmKBpPslNRa6xPxEBSuyFWHJGcacgbZO0WEB5IWPkNVDiwl
Nt0/u2qY6OJTbQ1S7zimK+CktDp6potQizqg8uKZHuieXpTd7Oj1p5OhXRSbkK01p3V00T1+VNle
DW6GZqKzbVR+9f1y1gUsJYFxXCtD124j8U9eeBz2RxHHS4Q5JtfqK42u4PPNvlvUcKzAQfFW7fno
L3EpaYNd85HN3NJCekVoFpOuvOuwalRvg4hYZWRziMUMX6MLAf2re769r2cBJ29M16Mr+Yo62gkE
UA82aVZd6Pc/V2gGPR14KEMZfzrkUXV6vrppaFv0FQNyELc5/k3FdEGbCMzockc+4WnPMOOZC9WB
lhUt4m27KNtCgFTwVnQfKqv4vWLp3RqqQCQaem/G2/otQXO3974saHfcFHnhTQa3ddN51YYHmr4o
hITSiEGCBwtpGZeVhoqG6ZPcIoPd6e7+dxto1ccd3aAcJwPNf5w8PO2D0Ut7wEg4BJId3EyKLJB0
SdiBRbhDlaYYUdiqRVGCTUFblclyn/JMGcDM1SyQV+SdKNSnV1hqZlyHCOZ5xdGeVx/Un9zc4eFA
vscruaSI3rtJK+uwb9z2L1E5lK/65XLtmX+nH9H9MEK8zqP3LU7dJY4l52usyji3P75Ry/X6p/d3
0neOmhXH19ySpo10KOtTh35ywmS2ooVXoA6iwyKnyxIoZvK8eVbjulvnEf6GimwffK69fhI08OM1
1bsiVN1Sm3No9zmrd565guwW2J7DSG1XIysE9Z8kXDdSmjeRk2z+2rZMFqm64mzdNfdJtHRCPsCp
7ozaE/8bJNhI9qobKqGKVY8LUWwQD29lRBDVaQcufDxBK85mvOL/L7KG9VleeLK8uyFgZ6NVeKPP
jMcru5maGeRN83fGOq/9nMjnRVIR29g0T+a7dqteMOzvdxZLvhVlUZ5df83gUsjtqb9NwLc/ntIf
iPnSHKObjtEhe3Ug9ei0xfSlkEhzZPmaLrSU6q0frdr1NzduSZzS7jPV3+WJ5nGSvr8Pgfiaz6aZ
BwUMN427xnqkdwdn6PbGCMkdJi5q/K8kETISNPzkwfb0ZwR3ZD+DkUwbw0GEjNxhQZsIJaRRbA/4
Q7ENtwnMj088fOYkusu9Z1hweAbmCbE2im4GfSn1hXbVakhV5rMvF+YjOiYbs/9FXp+9RXyhVwRI
KF3kxz44TUXBIfQjNGtB5lIVE6uCaWkkcQnk4ErLn8mSN2EjWTWFF2iaIr22918BSbESwc/7Jh0X
g3Fuzhj5PaXe+IiNvmMfaBb3KzfYpnjg6yg6Cp4Lqg4h92sbGQCjsPJWcblashvjiumj7btwkhKw
/bXXnGR+U3DkN+6pJN6oxyrBMTLWl/sym2F/VJSILBOkpSsQpQ1LF8Ps7rOkvFO9IoKHQhM6ES04
QrzZj3Q/Y0V0vPK3xn1eKc4lK0mxYQBVQk3al9TyjQjO2U2rc87YxjBuSUM/FPpF96xmYteG1paR
Dpmyz/fl5vo0KvkFH6gRXhuVjXsRUyJToBEYo6WQA11i6FKooS9LzzvvAJU2IXyunQUg7MfEL7pW
LDC6jur0tLaDnJVqQHGUf0Ljt35rbdETVjy+BOojvyPze8aPU6XY2G6S1x297/3l2rlokczh9D9c
hiR5EXUFW2wlmj/CwUXheRLDIZL4Ebqw2Qy83NU4os6yAx2SW27PFWdGXlIHjntAvlBKbOZOM/4R
G0sMVmY9iub/K5/OZ8M6ur7aBRTkudUDOKO9CHxASXWQ0QH/m8la1C4zli2sxsaMUMDKjuG6pnSa
zEsKgUeA+SJFKWemYdajLB+p7Ew1fXlUdUVLtU7iFxN6C6Ee9GCcVk6PNkLekyFBiQTfsNEfM2JN
sKVdO+F9i3gA/R/Sc1TESFer9aTiE50YOGF2QRtVVUOHvZssrikb5tW4BHJag3p59WQMBvu3cg4b
5LGtbfpKORM7bZkFzi6YslejNr5RVBpBuiEEPUm3345ZyEf7ldaCCjJ7kdcoaqLiUbsZZHEb90wy
gPBZMog8iayun7Hlak00fNIOYzUh11aa8u/mo5QdRVdOJDl3WiTX0m0gUvsdeVYeuyVtbzZorrGs
99Wrl9hDZIrekasl+2zCsCZu+xKESUIxUZxS2CVKfWzg2oaHnI0pXlX7kcTIlvYRE4vvR2a1f9Or
/XsMqYYIDIL5VGCssgydUoGxzYivBRkPBi7zlWEXmrE4t9dNqnJ6trQ2buYkytMDyF6lU7U0lGWq
8ulbtmEM9D1z8EAe9w9BCpMHufxC4S5TVJJJuLIEzmV0TTw6F5Zabt0Smt8414bayUNfNGe3teMu
x4hl0MTEGtDMMDcDhmaYXcismt/rekQ8aY/iyNd/2724hMy9s8jY6nqQ5V8Cm0S23fptcBigSRgi
tbWkElMurngmUBIahNj4nVwQ8h+6ejVtXZeEKqWEmn66PNy+BmaUbQwwMBYnEgEHoK6uFttrUr6q
yKEn/akqtU+0+leueUJA3Nwbg4qgFTdjpxzeAyksbbX4xz6AeaRZprP3FTCvihncH3kmFWYCdAWH
kBDI51oE4XtbnZ2XHiqcNFR0EL/K9+WRsISis/Xa/cIoNEyHKL3aBZWiul5V0DS6vYW7p4m3K2As
VSfro0C+y8DGzdp+NVfJxtBA7Az+x6v9QP69v1DrEpxTOKIqzuFQLEN8n8AuJUxDPpuOREZdbgOM
StRFI/2LyXzQTGtn+ePRzPozRwg1cFBbddbwSW0MTSwBi/NrzitKMHMNeH9PkYrkhHVVy8ZAN/KF
0TeG0PNpmYaXLYQoHQx6d9hZyhlbUU5zmFd+19vmPeutzzMoCc8CgOVJ3kmQcx8nBPJIYQ2IyXuU
RjB+EbBpKWF1jxYxFic9lgjEiroFqPFlegyFAKRuwTYPxlA1MGVyuVwIwrehrV33MyXl9fCH0KBP
hktzQp9gceQcSeHkQSJZH0C+ml8gcmho3RJN0qzth72YN/LS7agIRPkCKy4fJ1jaOORxUSyYHDs8
zKn4bQ7tfzmw/PN+LyYwHX8545wNUhgulNTah+OY/jTdBVXEJCBQ0GciaY06rw125QVBdsNzvmwM
w5ObAUazKldzd1YKr+uF7ICM8L+BFaeUPuULcNLD/jP/rc3niASpGScmUb1jORWQ0L1ovv9+eYGR
WUzclUGYk95KLQcsy5mMMECueOX0ChyGuf53CrudJTPwAUdpvM8i0pvmlxfB8VXU0UkVALOW+cNG
pFqmGWND9JY2LDDsLGum2wa2AhTXGq6DK8lKw643NQvwmwO7EdKz0T3MDy9oDg21Rf8kHItBu9iJ
iDOv7PhZ97inIDEvxq4tC06vyuj/m4bgmQaSw9nLzmsiKqtNfv55iuXILR85Kb2wcrGwU8jZ7HQ4
fxyad1VmRuSEFPQWXMMqf9bTpS7Aja/7DGkKMgG2vcNqwiuWDUEg9vY3V8IiR4xNrB10JK1GjzdD
ZKm01jcefEcChDoAokXNNrLP1Obe7G1otT9oQh28AjS5HmrOAYElU9TSCHC+cTMPqUh/thAgxLno
C/zs8g1Pk71+0QfYmxvG3JIWjGbHnXMVmmc8gig0U2e3pGS1Gqu4stDndhJh7CbCijZ4ZlTuOtVq
3mCJ8eLbFGzuvVFFnCUg70drvNrHXHicef7CFrK/zpB1ty/J4POrxdc40QZ/aT9nMw+CpN262awJ
zJ1PogN8WgP/kz5JS1VvOKwuNE3uhCTekMxDDXL3XUs/6W9KH7+4DUjbnE96eqiV8/K7XriujPdi
gel1Tk0LRRI6CqD14bg1sSdLoydwklMIyJu3s1LaC2OyXY4FDMSxQoGYvXU3bUAG0ehtKbI9zLJB
jDPmEGWU2f3MYGVGsZT9iqPU04jKwm+gCoM+crda2UpcSQwQtEzgLa21JrGqaU4BRD9fNl1cM7S/
QX1ogCXImPeSzMdihOMiTOMO/jGM1IvRXJdaBBWLGSMJNKzxFQEKzrSBl9dZN13kirA0E/F1mFQJ
ITKjmB9e1GjI87ozLit71ADHgEn0on00++TN77t/BgbMB+Xd6+4MBegPaT139vovJchMmugZ5oD9
Z9UZS76/UvQUxxZhLAjxTh7du2W8Rl3GwB0zRcmIMsw7Bq+zv/R9xa4nqB3WsCEuyJKANtuH2T+u
id05NZcAjofJLulkrAZcnZrRJVeu1vRUd50DIM8pdYi7NcPiA4wCL3T9B7/tnQHuxwU+h0QjTejo
MrYVLclAv2uijoIseMKiA0RsWg6UKxvO7RVFSV2AZinY5EQS7OIMOsaJg8BKA6v2G6o+J6qJkFE1
SD0UXpWRIp0IBHO5UgR4XVYx7SGTd5ogmtMp6CnuaKm4XpJp2nyKpP1QaNdMSKR4ycTNW5XtBHez
gTEusWerlyIfwJbxqF4C+yN4U5olLM8KbJrdSif2K9idxTKdiCkp7S4MfvEQa6/bhhGhwF24c/f/
2tvpYf+F+qLn3f4Mv29Tt48VZFoKAb+v0jiZYFpFIsiZHtXZKK26goMKPVD2MCIAorej6koJO1LR
otdvFBIlPHZ5BGiEM43TsnlVwf53hsYU3rMVYL9VDaLD3liQaoeRosf8FIUtlqa9jA5f+1o43GRP
HrvjUcjt7s5Spnd5npjg2pDsZ8nSlCwtGm1GmyXRlAmmHPOZm2mSczejTV6ECXnJi3dIzwakryZk
AW8sygSEyGv30FiqYRc2J8y1jYEBrKJdHNYVLxJsd6kGvUl9yFFVSL0kvkgjwBq8g88UgF6PW7gG
AzjzM8HyyWTswSu2MTZ/eUuUC5LTLt2575KpZzlKWmIwxMYSNFq1eHs+EYXwnfXDba514LjBDOYb
yRpqtBWghCDLSTvYBGlpgFeWjzzyUuCzeVFpkWoeYujxHEjIiq96ueT5Wchanyk1/9jiWhgBN3mM
ZLvrASuUCHxlyznrl5XL9iU7PHE8JbjYCTH2ijxicW5M/M9oJ4WOSUGChSIm3IrVFF3zCoPK2KE/
xAC3lTrOkvk5s0Ihh1VzblMtvIPsahAFGzxo9r7pcQTI1/da6agmHsj2/P7uoe3t9FlgwJ3OeotF
PltYOG3iExDdoOe7IzLFM+Lxyyi1YW3AN+lcurTO0o+xAWamvSSrESOzw6puk8nV29RNHVAOndhg
s2cRsUuiVcg5+z+d6TS3aIrDa+LFpy72b/XYNTt9A+TFUOke6yltI0lAA0upPBfVmsuO2oKiCvsY
hiGOTkwHbY7umsxxjjJAyBV4tjoazHXZkIMl5bVGyD2L2P4ZeuGoj94Z4spJIlM08YaACXw3g9hs
e4m8Z0xQqk6lwvfdRoMidRzLHuBIAjyUzNYAcX9j7SZMnKF1BEeAUGG8fyZFhE1Y32orft9US+9F
ce6icg27wGPDxMDkoXg0C6bgJHjDVY6dsAbRcWdsZRVoAZcZzv7Pkj48k+63KSJOeZVmQyoKaV/R
tsO+loJIeUBN6y72ektjLgCeJzFu0sfprxzld3zqtvSne/81xEWJypbaEp6bvVImf4oA5RXBB3ab
rGUoV6CRGR35hp9LV/vuQLfZ8uI3m8sjfSUxgE8Mz66tpQOO7lB1Vuxz8Z2l15M1NrbVQJCLhIU3
a60jAx6AW6ECJWlca/ooO7x4KSP70dUC+cK1fL2ki5NeuIAkQT7L7edRyL37e23VZi48gzbso+Z9
PulNnrZ3UfKSwW01OmxP52POK2E4KbvvgrmSORS0UosgulUvR87vIfAkz+sYvrBwfcjebt//pwRa
QfKMM/JPFuy5fZ19S2nqWj7yRk0KvnS9P2zDEIW0q0d1V3iAvIq4JQ22tZLxwuiLHe4XYhP9PwgO
ZEg9FVTX1UmI8+dliLCiJ/HP+5Fpfl9dyy7NWWT9M8jPGmh66qcV5agUqF2mwdEKuX+1zS4qThRv
tfrPgifRvPezYneUyoy0EjMli5Mge03UBX30z+M+qkPqyYtTKETZZzTGX+rqj5wwGTL88FNU1NcC
/+PiJzGgXWw4Do6w0VDoCQi2xZ6qVCNAKHfoGjCyJnjNLsSL+hFT+F6MxEJxrboPB9gZE4+doLDb
fGB4q0ED4WLGB5Ig32q7m1Vh56i4mv/cKYthMmCBUM7OW8XyG0PX4PfoAjmAJYFiZmiU2RmwwaMc
VkXZ5oVzPcn0g2lvbLfoC6nn8vAVKlvj29pbDuAtY2txnKaWQzcUXtte9vhXBe4o4m9i3T1VGqfy
/hoLqhEJcJ+niU5NL5pEsWrSSG/W54SMWrt3EDFlQBe2lsKk48iw5Ggz3dK4FDW3e0V4IWQOPYEZ
W04sXgm4sOsnGQYiDpAYJkwxLDOUne97yQG5I9OASeIwwWfsOhnedIzMRnagkhGijc8CPOoCUr//
ZDDAw5Cmw1PJtxpJ7Z7mr+mNEToOcpKmn1cas9+YserakiqTF3Q46w0ZEcmu8WMv0qit5eRzldei
0GycBw5i74MIiolyjHUpLHCKplsqmySqaMn4k0kbsLf22eRDpFpSJpmb3KnOKYs1nHMUEW1cLcZL
cRG+zu+bus75WfTDACuwqb8xD6dLrl71Rlpfu93ssZok1IZPlK8GaC1R+yCHltS6TAXBMGps+X0b
t+/9V+ZM3nUnA+gq1FkfSXVrFbfFei7AUZMkvFBm+uGsNlT77Ec7asAwu6NJSuXUgxpRXrYk2mT6
2ef0yghuqD5taR6uWItgbydc2eF8G8mb8GcziBlMIFCDDEwAbFWr6tPvtfe3YZPA2/RqRJRIPNvW
T6jhThXfoNpeZhWUtFRqGJw76nx+sUjbmFa4i76+7uK4lnMdZkRCR4YFcxW5oYsYUhcapCTX9gij
m15qKewWMdjRnl4uPmGR1RhXN09nWOGTvAoOszXJkkybUPB/XuXvJQmsMYXUYPNeW45osvN2OjBf
AUVBnN+Zn2DypX2v/KYvfLS4EpwjpfSaNaD6/F2Cyv9kPum3KUAMhmqTRMAkKaoUSjMTTct404+z
gxxF+dSme1iFWGBbd2eSjLvnfm5i8L4YNO/cskiqutC30UetRsgkSXFDgakwM05IkL6oMBknLjV7
pzKDsz7ASImb0hCMMkrZbpV/8GY24ADE2aWt+GTngk++7U9diLHftBvebdwNLOv035NEHnii/RxU
UHX7Xyjew9/Hz2LXYV+51rOOfLSxdD0+XMROFZauk80oExlkv8nTMtRAje2z0sernuYmsnHsDHOf
UdAm2xEO6NkkpUd9QdU1XO/58XJh3Sd2ViALHRHEo6Z8nLEcXexiePcjnAEF9fnDH+b/gwyolewv
YL/Y9oi05Z9uXWl22u0yI3k161Ez2LlpzDprV1enVoHXwGQRlB8LttdlxE9ptz/Qt0SNjJgrHfiR
NPHawj5rTrqe25jSxbwuuGf6gPr4jqqHDquCQDSAH0XW2/3iIxI9NSBLh0XSGG3OP7HBREtxhWkc
pKnLEtbAPA8EOmB+i8ILAWfZNXRiPqZYe52qfzObFDap4zf1HJ4jsyE5KIiLFVxiHuTXVFpoF3mF
+yUgERAP/gh1ovDa+Nery8ISwvv9yVJv8ksum+rl+HwY7bFzpR0hm2ZMdRSzVBk1S2wIk6q3aYHN
uFSvzPIRP4uAzvLBZp1NPw47Vq5KixKYpWfri/RpRw0FGt9/QG6uTxl6FFO9D+gR0NgMGYtcTlbN
EAI5eNDTFnJBUORmkXIqudHWDU6p+qS/TBypcqC3xzOONF4HYensr45HPp5AXhyB6i9RqzUStsW8
vCcCG3kohE2E2Ai2j6pya5nefXyXON+0PI7OGZDKQqmSBdoAfBi5Tf8CUPFt1l9e6QkvjAC3c8Kz
J8eNrr/4A/ZpXzmEFMxucs+itVFMYQkJD4ASnSi2aschXzVBgWicu6gdJJS+D7mowuMl9wgRyOEQ
cBFVcVhaWiBV4sldA33Kz1esb56vN+gTPqomd250eZGGIdHrFDAjGgLQ+fv8jl4eKOy4TixNGC4m
vqGfUFasgY35lH5x+ScP+6vf+0E2sqvXbccXFzhKguTf2tm/n2w1vEjTYt9inP+mjrQWuE5mxcCm
4XjJCxlP7zRiHDolMnlUsO1oWNGPD8Wvir+fr83ENTHAgUlNSgcfJ3oHNm6mWFfo+BWrKvUak6VM
xJEafTt4epAkOIJJ5Fblu+RAU4EGcuzv8qC9NYs+rFKvcrxB1o7jM64vezYyw3p1/TI8DCfJbjdJ
UThaxD/URvEMm6uU0kg08hZhsVsa3vlj4d1MyWGN9cp7jsBJLgW0DDeES85HSWmNWOnP904DaSBE
94H9DWH2ngZ0G1tX0GJj6ylScAx543MinrSSQXfSJbp1al+NjfNj3wcavPbj0NwUYjTaIPuBg4vN
GChnK8+zb3Nka6MSS2erLq/im2S3yFo5DfKv1EZGsXe30aofY4kYKKopzxWCSyLTz8gzV0GAIZmn
cb6iKj7EV14t8QuRYFgiYqdeK2zYGZh3AiWILxcuV5OgKu2WZZtPaYLj6xfCuJgU2+qKdekGyPdx
8jT49MRSX1kfQTYJbF75yYWHqo8IG9edDvj/haWJM8Av3thrxCOVOxLop8sGhQiDgyHdUkZwjrWB
DEoYYgI9n44Brt3/nVgF5R/fHk8WKrPCeT9EL6Cp4SJ7dwrp2G6s55vRrNSKQg/rZCDSJjwVGfpJ
7DzFvDqcF/jASweOxVaf0tqrjk1iyO4+sk4Ug2lHmOZruZSLtnxMUAgCQtsmeTWXyzsE50JWbjAD
D2on6nZrWHc/0wVFBkytxojJO7VSXhgHJlSz2jYwOKz0jY6S5NTEmuZqNM0ETngyC2Y49JOyAZpm
NzWuWoP826aOmp/VVlwVvT/nBx/aecw/yK0GQ/fZuIxyd0HR/6NGsXzQgT77aov5llBG+FBxB0Rf
CxP1P/XFkh2MgN/P8XbWvmsyyw+JdGHFgxqzeXlwD2Su/BFADoAbu4sIALlfB8qL12ZR0ZrMhy0u
hGvHktUpkvaxKdob1P24rLA8Z+BsT7wUUQDSonxpcuv/EtJbHKib0VV2TmJUu8x59Wx/3Oh08Diu
o10ZaYMujMeHtDusN9ftYj72UeyQrHQDHIXyslGyL6h8EirIgnBoaDr3TfI9eJkfshhvx+vjDYLq
J5gDFchkGwGOrGUM3Sa7c+Oqf9tLBEatUjX8DpIQTlg3YPyiXUJp/XbzTRZMOrRq50AFU0nr8rDL
Pqr+Mp1H/7P0Q/OY6lbd73tEVsn4rUcdG2akezICGqXOYfz9TCRihzfUpGMijZ6oihVvXJbqAuEJ
2Ib2mOdEPG7U//4WAAl/4VfDwCPyh85ADgV94vKV2ADVjGoTby6XXn2A2srLlT3lDYg2/+P7kaHG
OGDP5bnnJbfmUgP4vUNJH2KxCdvXPsVqhO7dnz5lAl7HrmDnIwPkxYDgry6RxK0OE9CBo3pmMGxi
Djl9a5+frKIMcMTANrisme6b48fuV1mHfvqAlJMu2HmJHMtzOiSX/c6CMeIBGWLFwd+3/uxeVrvi
oPAPTVGcEpFIJOzIsDttJOYdEQqAcVW9n8P0m3q+Vbs6GSZgD5PZ6KnLU/OzigsJVRKR9I4j+Ntv
d3CY2ztUPPdiyC/EG0D2RdLcSBEDzWxoKkOrtSrlIhCfIT7NpZDHiOengjFpIQEwJUv9kT4JKKRN
GJ9x9Idd/fMQJZwGCPmSUriQutLLCqFSaz2XCw4MIIZWi+TCIRVUcwlYvPr7ACrPrYgoMZfPSfgT
mCnFRoe5h6N+IMu5ZVlBacRp3ejtZyd+oBKdeSzXBKw2fDTY4Mg5xBH/xqvISrWjV8cJCnIN11AE
mZPw/QcDTfThtzPlKN9BpBSXTxIDg2//loYohomlxgCOSMzmufClKGgpWFEOymKGJblovMmVugeg
MRxagJmTJrHvrmEDsipu4jWZsaMw/cufJhkulR36uXh8+FWGAnGJuV8JCK12PeU+01RfRnmaswvB
tBo4XoFitZnZXfm0BwGigUd9QfxxqPWRPEb9UgGeN0bLav13IC0a9Qxw9CC3XBS0iyRsbTkLxu1x
2YsahgYdk86bfdcc0ipjOyK7MiZDzwBzt/FhU2jLQ5T6pGnbaTlD0FwubQlhX+7VMrPDC16tiZYy
y4qbi3VAX/kl4RkdLhOo/Mt7oybbJsXENZ7EuoobKzKyxp0E4p5YtGenphXU+zhmSk9qwxk1Q/9l
hdxFKgtrQDR/YhTerx2+BjMWVWvB3RJBNRRWkovxE1VLRTOpbzWtQ95FJ5bUDJtu0OgjMnoy/yh2
R1blpPS0vqe6c3P1dQxg3mb4A/0qdJaxYAVoV9X8QNeQCfbc9g2TkotCC9DKkyuB/8eLFU1DDUMQ
fqIZgMVPATd3tlmfv7a//Hq5MK/5/GouNGZO/io1wZ6VaVUIDcmJhhCWplCzn+Es1yEXp9okchkj
yOiZRMDD0S3q54WvUDNOYRC8ekR0mO1gU1QN3bnXrxi7NH/9CNMYchkqgjrJpKwiVfrek0XdhXOX
oSQqT8RmddU4DVipB1AaT1Y2t2SHo70qJ89n2KJiBcpK+pAi5YpyaExmTb+fgGGGTnN1bvWQ39v0
QBgAKWi+5gWpD2wJzKgONGoLshZVCzs/UETZ8neYsTfNsg/R0pRyZ0tR94r8XLxinAkvaU62ofSU
Nl4NULUXXKHyobmU8J3hTkMgnqS6tpo3PDvkn/ponQJrrHjIfWDApVMCwrp9J8T0Jh6pqN8R8OC6
MfZroVY5MD0yydnE51H75kSoIDdSZd5BbdQold5B8EWB0r7CuPcn5+dYeKvaOvUt9RHR8YBHdsC2
72SZhCv9/L5/XHDa6LAOS3t3BY+rRByox4O8ZD6Hp7ys3S1I3KFW1Fq1hw0MJYy9weX/N/PJ1aad
KS2LJg8vAuG1eTTPLi88Dr/oa4ZCxzqSE7A0Q69VaQT3gNvu1UWaKlouQ7dXeNDCBiPsVq47ylAx
Cj8h2kyTtydT4mJIn7zpZAGTiFnJ52xpzXLBlv5GjZdkSXBqUkMcphOt3XGA36EJAAy6frvvSi60
wxHZ/7gWonSzqh1P7+BzgJVgFbMvwE0nq/5rwT1mtGc/rCxVGwrPMprZ76qCiCJnoe9To2+SoZKu
YpckNg6YpyBHrMIV+jD087m107kjndsxAOGjbE9WHJgoXdHXJnSJSu1QjFnHrVRqqA6sYUq8obZA
m618zFJBjMKCbP62QCbJONFY0EVKzdcsqDvmyYzMCtGXUI+UERGWf+yuEhuoJM5vbkPFoow1alER
3m/62rY9V8l+XohXgiSs/kRiUpTfQ4NbYNZtwpiuIJaTL8H2QZ3XCJGXD630Uf4uvyExSvD6XMPl
dlVUZSjwuhMf9N4LqSkPGMKVvStKl9Bj/MC6UsYpbpetsX5TYLHZBYwmGmmLsUf9OL2o/K2M7xdO
/CLQlFayGJqOcGGea3wozgqSsKeVkiQAr9pWiywHZRb3M52N3TpXw39qdjwKzIM/rrWdn7Vsql8b
B4MrT6AIdyhTpyMPLuOxU7XN7dqR3i7aXeusQK802xRSmcR+1czDQeSRgWQ8/T45bblIjkZ4bSPe
rBprwEOOULTRAoTJpnRSU+Wyb5ZoALSfscI3+fPGCIAx1FoMMqICRcQgrkKvKEiDu8YeADG1ZTix
1+ngVqYWh6RtZadCMtE1x/xOULA6kabty6x7pnjqrtvA/Jo9E6VGo1RnzUvHAPs3cYpE/pelrjZZ
P/iCGBeKFnwHmcgZZJfrmiV+lgE7QwJFFKaWZQI7WcqZ/aq63auPOuVY5bDufvly/DDLrxu1jXwE
5oIABVOWs3MSbyT2nbu1VYoUcaCdx/wHfAHb08jOCunGt/KkqO96CPaPgqmUUjBLpdA7L2j5w8/f
LGRb6Qke36PFx1giQcNXzGuV2m0RLx6nF/G7Srm6fHqMEqvesWLJHzk7Bn7kZxpUpo1Gba7RK6HL
MdxCn4lXO8PF9f6uIrHwkpQnRPuotlvR8FZ8G6GkQykuuffWgbhIevaLlL1iZ26+kZa4iIxRfFz3
DOUSAYJ1jExLlq8aIqaADza1d9dMm4KyNwNOJUMVT92pVWrTtdrQp5tZiq14zazZqtJK9Cm7xIYS
AvtGfObsh5A35M5YhS4mReOCw7yGZDZwb3wcxzEq0IWrh7UQJTksP/C4BqvmwHdJCmBgGXGp/nR9
V6bxFL3xLyeKTNDRPiIXwTXPVUX1CNu8IfW1cese3nO7XW1WZ0hg8raFf49iLPr2JpiRA/Bfh/EW
n+gYtoZkT2HVo9MlhkwgFRAUD3z2IKsN5jcYQyyqO97w0JALCqoJ2rtGYJHWjKcPSSPGZHEjq8rj
gKWqoEuE4mUR0RxSQkjcmlJ/Z5GcIjoEnhhqjZlMii/MLyyEfrn+h1GlCB+ZBKjOdPIjF1ckaoOO
5T9WjWoKC3LK/VPM4cnonkiHZCmqEorIEha97AG3vg2x0M46MOr2rwEso52Y/ej40+Gequ3nH0bk
MA4MDW7jQtRXMOVBJ0ehXcCjOf5nkU7USlL/UDdJy/Z8oewQ+C39n2A9W2L38LbkwrW0rpxauaR/
ywRCUEXu9Hx6HSsbxNSt8s/ozVlSy+GThkZjzgpcnMkF0q33XDY97BqdSpEiduEQrVwoeQj40k/z
mChjXmgPzs+0o+5Mf6ldpuSV6vXZ5MOSUcbL5vhIvStnC6nOkqR9zKUO4C2Gn5DXHMtDgrS21fd4
n/P6Z1Bh4L+123QoJaK8uIYzypbRRiigLhvmUrjS6YSwdHBD5tc+m/thxCmwMsxqnroCI8BoJiRF
eGZEu3oq2WFbShnej78KHoDt0xpwsY2ljljCEO18YE+V63wrbdwsMchnGFSgl5W8Y8uPUPiCJRZz
y300Py68ky7UImD2aGfIc/TztgmGoy36Rr6c1IQBwfR8/xOzON4iv5kAPjgMYNfOWq0/wEtw5Rou
noukIpyvUm2m9KGssi9YCnBYdigRcVkUnFUV0jXR8CoSiXrW4ELtCHuZW06fAglS1NEFEVckrKHu
/9vQbgVSY8KYaWCtkkW+dh4olzYO0Qe6EkQcc/N2U9jWuqV0uLa6qUzabRyRIeVt7uSx4xDCXpy4
5DBUjukJCMRb4RK0JzLgU5cH/hHBSJKysiUsjth5v81x684LAGe374ZL8GcedCOImYCILuXkwNfh
o/mY15Zf/3Q42YqIaoI2Yt1o1EM9GG0ONwe6A4yfCysqvT9L+F3WwoVSrUAPQ1O3umYehSal1+pj
8zz2r1AyZ6+gZB+EM+Mfnx/ipIRf3WxJkFwk47KbxvWN8KlJDmbLZcFrhiieH5D1XHHjt9Dg22PI
Bb0GQZBAx1W9B30vBn76OJ4xthpndhaZaaz8rfUABLOndBYYlarjhc83cV7PU5MdDzx2KdhOwSuE
/3CJHAHRUKUBFJcUUu/y7NumECqrpqD9cpYTBaGI7Gf31hD9oft7W6lz6G1rXUMwlG6f8v2h4nxE
rNTpWZqtwTd7RMxH8QlZlgJX9trYYdaNCLB9IpI4vfP3gHlw6RVMZc43BNpRNHSRa3rXzAX9/f3l
qU9MLC6YzOQ7WiPnZgETWfEbKdNo1fDpEGRtvuOQmxfqGEI/y+EGko6Gq4ARHtm0qB9FJp8A4d+z
HpHKWd8N7xtnyIYJAwPQt1bdkEgs0DUy7+Oc9M9J4/GGNx8kriI4gV1GCHS8k4O/MpXLxhFvCfbz
ptR+PVia2t3jI33DAE+S5ItUNMZIkuE14P3bIP+3OnZT1GPghNl/KKVi+IXZ5YQZD2f3xFtqO8OV
IbLmm0UuKvcAwR3DYybCtYKOc9aa3HP+WnDA2nh7nGFpDPFBFbgZ6q7gunl0TMA05R2wrB4fjfFF
dDjkltBoGsHArPA/mmhe8x5v+iSihh70BS3rpRWirLoiaPYo8ZNB68eJ6+jtX5/vjaSrVH1umOMD
vdKBWsO90TdVOMPgWSP86R/AroPdEnAGTN8Q3328bjqP3Nk0SfGdxkuRg+K0TNtDJUjRHoccokT+
ZsMouD+91IQCUp4ClDCgi6abeDJEUl81gdigL10XmUvFqvBihVi8bcN4LpCFHrvjkKkKl2but/C7
YhK5NYYW+JO+pQdWqmDVqvfBZYTmO6YHCysBkj5ROP7H0ZLziAtn3wzXrqHcX+YNRFgw3uMVsCXx
zzz/WYjjvYdaDejeeEYclek3AnwA+AlkzCaq383kkP/B/tU74//MUmLeBSl33WsvOQf622MXOxFB
MEbGc/UZMNoXdoj2cn9AnSmtAFHaivXesRxy4gbs2X4KY5BYa6B//Ecyv7aEgMwSjyXsjioEyYos
6G1T07+wKRDB+e+o6ZkWvJ9w6wf31YD/6T4lhWrG9VxnBEaZiYSBHm1bqEIo/Dw4oMbffqivCL9X
zONoZxmzjtdWTRtFA2ynTEtupEKs4pgefwHnWpTUALh8lGdZXPZnTGrG1AOjRNkG60mN7cmpz4dr
Fnuuc82DWAyW3ZwxFgv41Cecx2SVTlbCeO/S5ZXv25BzShhPVxVrcIX/xVrj43ewrXnZhrhJk9sA
3U57t7l0pW2C8q8QIHETETqDVYEaBFvUNK6RhuoCceaLWTGw1rQ3kImIOcJ0GhZMzrpxmjslvVAE
ssgIdvG/ThxYN1raUbLmr+thvkKTQRhGXXY9I4LMSgPbGheztPZxPOHoU7MzagZdl82i3Ex6VGan
dHBg2IEcbUP2ujrA2vYu0zQr8rqFXEz4i6T/wowS9jPtCy/W0ip539UrWp/EOm0ZpQ2WtC+R0uMA
Oju7MQd/oCfyHVZoeCP3KDXdH1JTIRjoM4s0B1sSBmeQRgA0C90/AemjrmoD9ZrLXv6tEV+xcO4V
WbMmF2qaBnX7DQXIDnmsf7QFWfkhzYZk106SycH19bb32zU9W6wXxFb/yLFklEXSOuJZ1OpyTgUW
Q5zuh/JNXmK7UFbqysa5cq4zBN/7e9M88FBJxCSTSNTzkURLJbv0L8zyb/c3zerMAWvLBOR9wxBz
D8jqTLdW9j67/60X4GQxgYSME+MT1P9Ola5BFRSavvwlncJCLj4tn67Glhv8lzvftNGLTv6jcXXu
+W8fIwm/oHcLmAM/gAwBQEujEwNxAbBRZxDpmU5lWgCi6QwZBTCLM6gpQvPYo68trHhkitJ0oJHY
fgzD32YL8XE/TN8JESFeMnmHxQAmCCMPyE8dcraSR3nRT018Q6XAsd9rCvEPMTy+4hyL24o+L9Qq
74yIdWSiWvIXSH9wIcMW0xxsGf9uR8bZCe4yYqbdBo19FEiVeLB7F57jv5O5VjrEPvLmbY4GwcLk
cr/Q9GdUW20Df5x3BsvkKs9tJIX9hwWni+1Z5ENaDEysScY8/pfezPgJ2f1LtOOp6A27N3iqAEAt
D+e89BqWGlOZZbseXGH9yvTrnJrRP+qyZ7aWrzgCw3xA8235iwjvC2UBl+ZyigXZwxfzMjUwvhi+
SbemXUSM7S8GKntuPyUV8RLZwyYYXMxG9AKzGsLtprsbr/2mghcr7kmcT36ku+QE6kp9+LFiQX0d
reIypahaHykxkHWOruWMQXIkYFr5G2OA5i+H9Dp8YmccVqQ7L7MJibIF7/SmwusI+sV9HF3ghWXx
mw6SLa8ZFlfVxyrWqdwAhUwfeSN+dFHs7DvO/kaHYLRHF90pjq7mb2kr1Ofjrq8tBp2C8VE5OfzV
B5I+iFAtEBkQ5y0hbSW6ehZ/mnWiUKXDsoahuQ6g6aGvbsl7JTHPUIUtqXkDdJdga1aglfk1INMH
I6T+COyoW2DgIzHKNqcRzhLOis0c+AogILcfEoyTgeJrCRFmDqT8YFx9Cfkrx/MW8lSuv/FsigsZ
XQ9l8/IPWWHnrPUgVZ35rqhZ4QPI09JZkztWv/wMiEf8tdTA3ECX0aBhFRAbtsgsOPJvnkJYpNtw
YuSltnOjvnXRA9X9rHGaUIoLWvrJi1X13DGgipoPRLC5EBMZJJNDwqIWxCRBRmvOBNOuea6dBQqD
acGVeNUXL4oh3jHLxtZ6i1rlR0c0DSDt1tIVzZ+xMcRdE4Q8M5zR4aNifX+2hCBJSCNBEnJoNN57
f6+qqvXoJtuonJx3tDI/EG2M1yAyX0GhzuAgMabiNtOYXsq9T3zUyfhONpRqH1Lg/XFC/pafRz2+
Odr9YiGpGiYvDb+2BWaNfKSvidZEJGSDbWlEFrHAwwAkRxxcMLJLozhsIRJU/V6MpDlhIHwpnLMa
TQ0HDC1cpHt4C5niCJ9utRaMXaF5A7JMNM5mBeuXDe3zlHe1W3BWU+nQvb0ZITGsUH+224padb4M
OApRMIRCEpMiWP5QE9gWWiM7yiOUJCt5CkvttjVtyaeBhu1O2FVafDEDDr4ctDoQrar6kf12rQu9
Ax8AIR6QNBRggE79H6Bs3OZbY4vUgUcnmV8L+hEFXHSw5WknD9YrcGMJLTsWkh8O9hK3wSdkQNaL
qivwBLM+Uua+m1SESsd4kSn8jGvVmedECiQRqjpYhRVI2oP26qU13WBRXIZK/D9C4hTZQYO3ziIM
iRt6iPOfdDq8Y+mEZP1raBlZEcqGySOMvyianmOlCHi3HIs0BCK5X864ZbykQsocGbU1Dt4kgxQ/
m2+WZjPXYB+TELYBn78fMxDg/4tcIMlQPEkWI7BCk2Bfz+ZE5OFX+a4Bu1OtuhJFr/wQgBY1QP70
X2Qk2pLcz+vcoVm7Ju/UtNycndXter9uJoW9z7TmlsC7VaVowIXupqrCdX0RrpxlIZFqc8RgZX6u
kiE4u6J6tIRgV0ehK093jMkUkkI3NmirAEsK9BZhJIL0TpoRZ0ZKmruoK9sC06B9fya31nMWcnxG
DO1lY4eNK/OZcil16qDeuD3A0d2lqLaF80JcGUHTIMZpGWnYjoC9FdNrwDJRTOJZB8yOakxV/0mC
zUFQGFpPTUKaVIhZJVXF++AzUVlh7LWr4TGgssjEIgXYj1BCaQ7XjToxVL1S3APpZhaMSIDYBEfo
MS79oBvcDNXa0+rCThUR53fhhX4rLtML9FtHjUnbDk0V6mpNf06so+XiuyF5QSc5KfW/LsQw1XGv
9usTNvhyJxB0H+qBgLEaN0uIaDb74Xbrn7K4F1WJlp1jOrmM69IzAYwpNrgKNbFGKau/llRhAV5x
fcAae/48JbbYppecVAmMugg2fhEJIWzO7/ba72KHScEvRS4RhookLmw5rMtLjEUYXwW+xv7f18ul
xVtKH2yuCFAZzzeROKCsxT8yKFt8wZxpXnZu+cMPauYGYlyG1tYaDbpLp3YuDWUFqR8WMyZF7rYl
DuNB/c4oUC+3pfyzkV6fbj8UpdC/GlFvIaP9PGn1DwlFYyHtYmpwFJVzS/cbmkqwa+lYCxNy1Kz3
wq9QrveLci5ChtOcQ6IAKShXA6wb6f4s1soOFn9QGc1FMQprGfSZhbNFqExMts47eWGWfj1PENQ4
lzlIkyrza+Imn+ukPrkagL3N0sopnDLcD4YahSmeqrLIEqLx0Y0T67/VoyC4x+PzlnRKn1oRGtby
EbBV3fL/JWN6Li/og4GqloN0YTQs1a7Rb83pQzk5PIF1035QfefWk8BmmuHrisEgS+WeaXJPIEkX
QlAzNkkGQ8YQB6FOLsS5elMVU4pPme+yWnT83qoE1L/Bvm4ZiPZQ7xqFDRBjoX+T70qZGP9cco/2
FlGOfYAf8KCim9VjBnQe5TUjJ5EdPQtP83tGRNbgcnw5+ZzOvV8AXVSW9y2TRGg7FNGKhm1Md/Ua
puKzIJBuXm/gR7gKSpC+lQCynltyr48dE+InlXobFZMX3mR30HGJec0D0Jy5nJYp75mJ410R5bHc
3Q0mBqjwd+tGqHoWnRQO76bNg6sGjpDkJbn1gG7i5sYi/MmvraLWqxPkt4LhYkpi7aohT2goNvxE
88C925IIR44xMFJJomT8BcsmD2Jx7X8mqzYrmFxKmJeTzQ6iVTBh9SVs1UsEC9s9Bua6Yh+oXvL2
rK4CZBIoh/fp+09f7wO7otz8kpzw1RNB+7U8qeGgWTyeLwRt80isS5rfkfJAL0lCF3oLOeE5+5u2
VF/1wN9+J7ka0FTLM7SLL7oPaZuWg4WoMaHSulfO9s0a46JzKmx1yxPxo3zm0wFtkCI+lE5XM4jC
7L0npkfI+IdtyDb40VzLPlH7msr5Q/jYhXizFmqE8jUYKExU73AJOoVTKdV1yJ11is5/kiG1ps/D
SsWoq0J47JOqE6GNLqwkJqhDUVeHg2SaWLjdVuEPkwnA4gZh+aUfeliUzPC9eKFEtOAuEkRp2H9x
h2UULKnacHqlOxljgHEaDssxcbHBpDG2hJQGEhILVT9GEN9oln2HmBwg2Y4dXeeq/2Nq8FH8l/2q
JQ/3QPKWKzD+FQSOcb266Qxf4pTIYyNlmUSUUKZBwHUTAAPM/FyIglpU+wHON1CB84xQh45btQbG
GjdbiZF2tqnh2ISV3fV5OBhcvkiDlo5Ey4O2IAcntW5wxz+JoBwCavxEO87ZPGApvcPdc+SOgD2w
3YRQg3g9lbcXS60sQhG3THV+dsECScmehY/bDsNMJ3DoAtQwrcuI0hAMtmwYD6e5PAnEobRSA+OA
pdv5JIch1rtTlNPFfzHmFUqepHxwSIB3zam4Il3EmkG+FUsiZso16LQw+NawQSPYevq5ZbgSf8m1
hngEK5chaqqQmihX1Zc9+Z1vJfo4vGpH1+xAzW75Lp5HhoN07zm0OTf9VvWqTTQGsq3pVrswYNuF
vxbil2qqOdVKnEW9UFjtkSHzHp3qN+74u/RcFu5Wimp464R89s8HVvwcWIZcuIQGEnE7+eBLLg9r
dZYAIZyuPuxPSiDDK1LB1hY2fEARSfidhePLLLG4m93bY+cDSF5GrsVUDHs7Z1j21B+5xFhmjuXd
aA/cjQXfMzz5FL7NIi1nCF4DNyblbnz6IzJFbir7Y9f5bRY80vz8lcaJqbS7WiNBbNodYhYipgpV
cUkqHI6UBuuNYE+DpZvMs3PBIWcL3saE28AKSH2xSSc6e8ckg+RSP40Vhu/S7/7Etu3YjXxMNsb3
wAOjfWqWySsg4804e0KaOhhdgf++1IcgtED64DrPs+NJHC7y/Ouuvde0OwydHGMesazvzw9Yhxsn
iXVbhsyuGGnT0XLwcgHFmx1+6KeeRNuZ9YswZlgTmtArig1G9eDB18/jWoTFrp47bkcTumXw18IB
X1bpCR5C1VViNYSNJPgY+e0PkumII7pCYV3zyCRME9SzIpKurjBmOkvK39hOmZJpYYJvYNIeqkjC
Pvg2KDgMHbL62usZd2AUSIjhjIlcOWQq83nZ+nOv9xVJczsULugc1OcjKppuJE9X/lGhTW7n6IHp
H446k2nMdYhm1Y42gE0o3bWcPqvF2evwR+utirFe9JbxBOwPG9Rcj89MOTrRlXxNomWPLoiqwj20
k9RuXtM3JLZpkgQOZEjnIAl2sCXlGIAy4DTD4CYPKi9DqexF1iNiTjf+FLPcqU0JjwL9lpFXeod1
rIGY1Xar+nNCrv9UDWNnAJq6+B1oMMiR8HSPFOQPuGgdzSgfjEgC6l30voiONqgk6TZAu+BVesqf
XsI6mPNPMxx6U7epNIYwnxB1zTAng7DZF0xrvJYyecbi9SJEeuSz9stB5aCHx16o05/sKstZdyMy
mN6uc0qqFTIbkOZnG0GR6AL3N9UmuirTgtLA8SBUv7fRFuPs+aW3/rIOzQdscyEnPcm0EZ++pXuj
r0ewhBGXuyjvImZ9m0euB9D68PvteNeV7YkjLwo8k6m2+HYHspSDiTBLg6aJkQjLfvScKYjqGQbt
uMsbNvmbzPu8+11iiC/JWuyaG9s72zvUDvQe6uoW/eF6mx70Ocx6Cnw9lIM1GAK5TS2keheAzuUX
ZedM+Epa6iq3bEl99GMYTLKMvimEudinha+Pwlt98zqpscnDpl2+Jy8krBkqJrcAf4jgraTF9ce+
kyM0Y8Qfg2zBjnDE4Va8W1NyS5whKGDtKaZ2AXCPOqZxVs2FFH4O4MliL9KLJsiis1k+6KqlGO9R
PqDk78OucgktKhXl/x8Oi4/+mR1/eLZaKirsgEtrOsk7c2JELd4tkhAUUAAJ+IHnGF6x2dCjEgyF
XOAJW7bO1tV0hqavBlaSB1Rv4WW20/q3ZPj/8zRpUboeEkRrfsuT8NdUKh+n4nqNtGgnLhpR7ZEl
46d1hGPdwl/H/ey0Tsf7vEWreDZb5SkR2PaIT1gloRe/TmV1Ap5qTQ7jR7WtcnoOAgUwABivQWBv
M0ECtSxSm6cJmioiGt9TnoiOL+F3oemqXQydUlBZ4RNGG1UxQ1RAlaLXurApBW79HPYSynj4iq7d
cmy6q6UwHO1E2651tar0MXcfkafrLGbW6dzErZzlEtus/twKFPyScaKeRU9iombI0SNoezciM/LW
xsD9VdEr8JfhesNtojPwEJvMl+Amrumos3oRGLkCQ3W4z9C2zXHxA2/oNpNfTwdYdHfj7T4lvU7h
RntPn18AK2gf7FeGf9yz5dmpeiLCUY0B+YJaF82GSni01/XDlz6TYNbdJBbjIORbmiZTsFbhInii
UMw8CeL1qovZhDRBIsd8bbWuUTtGIUx8FhMikojNAtKpjWCAITl3aLRCEfsAXAvxSW45egLHVBY1
VfZNkYhs+hhF+/vXzbzQTNTgFcTaehSeaPYmJlA1VRa1dwhqpRhtQxEXi9dKWQ0obw5HJKj4I9zM
EyvmJ4hC26+HpPWjPFv4+al2FxhWNwoaBgsHV8u6r8kc4WKTYZIyNaqCpmTwauJMIcNsuqgN8I83
Y0YSnjyMkAIhTMxMXZj+6TxqeYSuxuTUO/pV1WPXz8eWJttZHFQ0JtJTo5nWpgglITQtyOGGenfg
71fSSRK0PZRkIZblaF9SGer+sL+haKnOuFG75jJcbpJG8bhHzsihB88/Fbz+cyp17YTv8Lj3atXk
KoCbsy9WQvglSjH4xkWuNbmQ2V2VuL20dp8mwc9J6Stwc9bPW9bgxRndqvfUYLyK67SywB10Y100
6iLgRjEc8/7PIOfh4DLCY+Jbr739W2wd7FItgXnwkxTC+ReUeaTclnqCNapczUhN/mzT2Dm+i5jj
uI3xO4HUtKc1SuCAi2iJTf5k70/gGtUy1d1edmkCyJh50RUKc0T1zhwSF2jONVk6oUS8bQ3rGk54
utCSzpYOSGCpsnbkMo776zNAOvxPhXc+EpD2B/8u+OeHh/gY3OaikurfK8Lu9lmsTWFwC+s0mG9G
mPzDQ5bUJmrkEAzCLcd5eHqRX7bUKMDBqxRYJaHEMzRhfkdNYqvsO+uIAcRmATfQIi7d1RzwjKqz
efqnyi3q8cqSqE1qnms3u5qTWAlJ+IfHt5s7D/K18ZpRB/qjWRbqj8ELAepcdg3UlKIpN6NPI5kK
Qy9mD+TpBSvQMF07sqg26yXNiYeH2/dpoPNUFIECovoUkU2X03gdK39PSwgnviGmQEGrudHEcXnV
QdONdImTkcUWcCYtUVVEmzvc95OH9JUyOruYChnko3mbYF8XqDv8mhN6R2F2VcPgNqeEQBDnif8u
BY0jUJc2g/Jd8lE0xd19z/Y8juSSTG7G7uLdumS0eLekNl4qRUpScFgGhiS/8CTWTeIGJL2okHcE
An68WA8jCbNPi207um6m8NctSu3u2rI+Sm5VX5nB5+php8dZ8QjHaC1EoYug9SQXx2Dkn10QhAB3
Y7vUYhxfEMLCX3feXzzW0sARlmCOdCAIQY/I2lqtNMevJD7QplvHkHwAfFHDfqkijVq+iJhr36Mh
lZMhib43ChIyEeELwVkHfbiWUCVHrhNf1YuyttG8Bkxe9bnNWTv4fHrAunD107OVOitkDiVek18z
2slT4KN5xMYCEQEUh6Di0E8fXdk1sUTwQ91RNhvtkavvOC0jZoyYzgCNXtEWuriU4QU7ah5g2XR7
i/UHh/khZyJQtwtPkgRX/dZ09U4PBFzgBLyFDTCRuOVLkJYneEaBTjtoogD9fHh/xgVsnWH/lAFN
rRkgDC674KVA5QSKynEWtth3DU6tuAWmO0CVDp30gcEgrinbh5iURfsB8gzy65Umocs00ofwOgx/
4Id9qlUexIIxcyuWD17FLBRlLUIZ3DbPZscG2YHkYayPse2xifjvaemN13CrDGHlD1hkA5NZ+wL4
KzBBGvzOwqX0DlKX8G8q1lK1fdkt/FutfdBegNtGhdERgcCyxoKLhT/5Es+9BgFo+aEtmPEBDW+o
0PCaOiTeEZDpWEDEysSf0+y3mgzIR8q7CORGj8uEZOKMO0nQCh71HLmfykrvCURYHQZVqvRcl7zX
iw+n4LMAt1/jr+buu1LXryfTYLyXC+Arj6UcPzJ+1FcQY3XRNGJkCRHvXb36pgFvCQ9LjwwY0PUa
OKf69F3JzTPy2lfpP0siym+Q8sO+35MZlQJjhEO5R44ljLQRRCl+5dI/sQ2tiZoqKOMF+yKL8uhy
knLCRupiCvDCwk34A8NAoDBUFrt4NUeNUauTbVc0K87KvJtO1mnFdJ3zbHG34C/FFezIvO7yz5tb
VdwX3tHy4zmyvNExKKSKuwsEmJV49OifWq/PeOkKje+nbxkW6fs//mrvXKAOd0xOzlsbAP7TU5Ap
sLu83H+YWzCQnhPn6p5FygR+aF3mFAmocTufigq9CR6iknCrHJNCSrNYbl6YiMT9hPL/XW7VBAlp
WxcB1+4cwXY5K0OK9zLxBvOGiGhhgbDao+4j3s+lMXLne2zFkX7WEaanJEfEtiNCNt9u/nslGkSy
ifSmKxVK6pM6mFMsIGoFPR0bN6CO03iELoKBFhUKoDhUPAnKRArgMR0x1dgoAIly0wbUzaUQtYU5
1VKZjX8Nanf/8gt46GOeBZ9M35pgihzyrzUbaIWraS6ohXmU1w9BUmLbyn/g7lMhYyoggMCevEFp
XrcZAT9KtSVLPI5NW5RzBYOTekA7Rp5JU4P3EQ4HFyiRfknLVHvF7j+yypLDeuKR2Ce8HbvRf0PU
ul5peIhBAq6XvDY7L33COwj86Z+Wvq6gXgLiYWstg5hahFLxv2gVoCXPDh3nryKXTXzMFrbYYeF2
nkt1cvZPgI3kYCBkwZewa2oQuSHVM5KVZim+sGIj1yXDbFf/rDQDEqK9kTizlsdM4do6PJrcQypd
aKmB5bk26x2bju6RKo/pUuhOe6PUiuhuDlmtgHz23e9UhgbzqTm8uQvqj+POLZjua1ESNGGDFc6B
fQXIfEgH+0aLFB6mubdyX7oB5w2+ZLBtiYahMHI9JKcdTxYkM+rlwVTVJZmwqIh37n/zN1KK+S4m
L7CtmsjqZgPyVGZDH2whjfUdaWCZW+nvXB/2VuwJAnEo1EyUKux10rkZSkAb0e/wCH3/zXQdvMWj
AIOq6okpV4uSBn425iLRraCClBoG7iq/d8X1RL4k6HJeqDnoRI4MN47sJDNgiib4WabVQMW7qt95
mOJLg9jrS2m+QXUoORm+1OR7vuBaGf30Qptk6VpCh/eCkUlO9jg7p8ueyFwX3uvEljINs/7AN3LH
0Rpo90iXT3xFA9D2qKkci3ZzGJmRJZzXnfaYEjCoUqsI3BfFyU6w1f61qClhvTn0S5fHv5XYfeNa
kqBvcrDLTWVTD1sJvO8HG6RJyurM9UQ4GI1ZRBxLIp7vCuC1elvi7iazUQyyvUHlNJJNKSS6d/9N
SMMfGmTCyYx65QLCYpCyOFyRFYXQO9SoK7QQvw1OJrAUKpPkyOzwX0aiiQBHMBkIQPv5BzfPMdcp
Ob85lryM4OXGiU2MInG1ejkogYimH5n9UU9JkdUAZR5wPEh6IZsamUxkJSIQI95sbHoiVGM8EbnW
nfpTP2Kwe+ZOzNyHwj5QNFM9iIizJXLPPijwZMicGQH5Fd1rRKM89uVjZI2An/UOTRVE7QyywVWo
S7pK2r46LPdycsE36yz6+3a7yUI9DKLRr5EJlokjikPI6g5Yfc89SXb/XTJuNTBHenCEheyB9Z0I
c79OytKp5w0iSG4Qx95Rw2BkzAUPA76bWiGx22MVyD6ydn32yVM6xPkiHO9t+0Sd/EirB1uMYFsH
+Sp9erme9xief7L2XiQPZJAm3+2ywVemtEmp87SyKyRoQbM2OCxbZ/ND1NP/55/jTpxxFohedz6Y
iK8a3QxCwmazMfonxTPWqdPMZ07cSjV90a1zuswws7wn0Q3EEgu6ThxBwnqkPrEHXVfpgHThiKkK
mzmbhxvAWLVqX5+SY3lnJm/7XkRIaC/UDS6UcuB+iLD/ef1lBr3Bo/R9BnHnLBziTHCLPWYcVUfU
KPVuppSyvGc3LMD1nm++UA/uyuCXlrVMdxz15/8G8YPM3SFpLVsBlv3F682BqsbfZLY2iKtFWBP1
gzbVvRM7IovVvyk9Iyvc+eqSKePgDySakSBwJ297K/y09oatrUh4iMMxwgRemCOZ+Rf0B/k5Ztdl
5eTpv/VbndBpwubsUdqMVlReN3G5hpFgGTDgU2h/mZ0VH0GdQpskh50jcUYKskpSkjpg1uWITIDm
1FDsxUw1i+08VQkCnpI4tbY4Px1z1CM5OLvCRbF/4mkaU7oPcbIRr3D+HskssEfsI00Rs0qbs7sq
OXrZxbIfe6WVrudDmjMsBr2Ho30WimHft7GlOYabiR1OZqHmmtTH46oLyiL3aUoE6Y3z1VhZF1Hk
NDQKBBM9tdfG7Lpz0ZLDguabIRamksmqORCJSrFdiZiKWD6Ewr24t/ApNywiM9amwH2ifPEzK/YZ
yz5GQ13r2oDUKM+A0hRREpnIksltVVfVD7HDZ6c85UJgFRmLUIkK8gLhqPgrijl1oHihqSBHUT8D
lrpNKEimRQYh2r0dToGWX+Ivqv6DyuHzFCvhf7LfR2RTYWIbVYS6GAF+isGA52tLc7HAZCPQU/kP
Z7BXwyVQFmlTUyiKjTJeDQJYFILqMYwSEbaTJE4CykEkBj3pl0aa2uSa2CoIbiTYiyMwzTxm0thJ
BhFJvkcYbVzQavA6+pzg/JmikElSbuyRlFg9ABdBymwmerv9cSo0YWfIqKF5Qpzlrao6ku+2ok6k
SYFgP15ApWEYOR5auTMrr3WkDv3vtCNEqNaVv4EM0Jaj7l7NdWG6M1FDy3IJKshjmfXh6tBcc8JH
3EOUbYTXR23itGRCJuYVk3Z9qiULBdh5IDWi+El1AO04uFdY1UbPIyAlP9Q5lajkMxuHuSpLRRxU
WICjoLv6KnREid1rbxF0xCOH2rJmWhW+9sV0wXS28UNvfymvZgOpkYAMLdWbynixmp9lhczpc7iZ
qvHnVlPbB8p0AhTvIkYMA58+QfhsDUYp8YPpvJ2Bj2miPmZH1q151cdtM8wOj+0LzTpPLIaTeOfQ
Ec+3tfFZeLNAcJ2Sp+M1L2ndmAjYUbZZkJx3MHZ2F5+jydKewvguGSvmDcxYxWrEkGMcL5FwYXg+
zF1Sy17hKkgqfbzqI+lOpvYmvdSGf4pQhF4SzFUlXxsNkS/2t6QUsKV4hZCVmB02L5b3/UTLBR7I
LEyy69Z8m2jIgnik/ciDIaHJ5dNMsWi7d62QW9JP0Yv40ozYvqsXB1Zor2mRTNi4Mlb1uc88mqpp
Um77rFAwjVPqTLxHqb8S1f2vHqTSfjDg6aIAcZ8bR49PcJpBmnnkLOEVHC+Umm4WPz7H9z2lOQf+
EsUJt+FoajF7qj7tLQvIYEM3dqUylCA4Q5J40ZQxWARpEr9GwMfhnAZ1/lUcOxAJplkokpBan9Ck
pCj/99rpusqR7GUvgQboSIngUS3qoYWXEy4u4FZrUdR/aiftduvnD+Dm/5M7ZGMdA6ACK/arBiMu
FZFyzmmQnkEue4SgYAMebjKz8eCHkatdfvtIYS0rNay5w3P6KyWlfV+wWS+8wZRWUT2LrjmyX5pK
geTRUnd/+VbGmFnrwaOsLHOOlMreJztqwNfRWysHEbJpGqRMgaOJj8+LSVl1aTvGA+ivKU/dWw9H
7GjDCMRSnGGd+jykCTZuEQ7G7x5l+vk90b9UiCKq+6bjVqF4qbquwoC2ZeNU1z0fdiRkI5I1Adp4
8zDGjhHwwqv1ZuEpLH5vpPZUvDmt9mIiKu6BOpHU3OVECXyXRsFnygq1aW2JFWY7hG76evGDPfMd
KZ7sCOMv7Ja+H5Hn9+hpU/WNa5bcwiMyRgKHKKW3VPeZog1Eaztcq9lfyBaf+sT8oGD6F8pzH1fa
UC2UPNz5RtfDyAc12HcSJRfxyrYUVjE+01gZd5hm6jfk/LB3xI8TwrLACEwCufkBZr95VXXra4FJ
3LXUSfPkNC5u9fwWDebxTNy8RwpvQwM7DlkW9JuxUHVoOH9J5lJUl6oLXNttkAKwV9Xfqu4Brjfg
MqZKzvDwgLtwFMKlTfrNSdXqHC2DQZknuido1uxVCyEpKZ+f4GhUOJ0xNW2rSYnVbyhPaQGyST2X
2eUxnyHhTF2LPu16LFJ1QG23XFQRnjQ4uxqlJankMPfg8UNHjX3J7mzvrPEwlFgAF3ryVLWjNhsD
SfC5JPUzSZphkUQ1icHet0tkbCxa4ky3yurRao0UHtrCuvGY6VaHIQqr8XRRv/MsMgYvVQHYZ8uL
NJ5Yee3EStD8n1dgZsgDrMFS5UkquWxtF/p2Tt1ElDX7xpCp/Y0fj7D5I+lrdPQR4guUjTkBIcmk
FFvgGQGTeLSmAAxgNfF+xO0ZgEnibNzwHjZP30+aasgodYh0wsDg9j4DlH7lLHFSWPR1mbEs6+bn
2TUvDby5nAAZ8GcZCpxKMQRpLot7N0r16AqBBROzogTClzIU3aW/+CPW3mVLnSq2KDt4XhJOTrDj
3C2t7C0/84wGiRN6fz8X0yYkaoR9In/4+6fWz0Q3yLr3HeOJuG/pU2xeZoYIVLwx1C156hrouqY8
E91X/+UlYb9lIvLzqkkCa3PSeV8Rc/B/bjR+5xLdVocIAhyQXh+Plmh14xs9JpTtzhRS/YoaDsBl
H/iAN/m71zWbOHz7OSYVjq19v6ndKicN/6jAwH8RjBk67VTDnmNE4jCfdd1zlX4ykcD60G5CzLRP
p7YSho/KCK+sWEKnrIAdgvL4wWe9fnOzxX8IFH+HEKBEs9nGr/PtGy/Nu/nym+unHOmXXO/Ezn85
5yEmshQ2ye1pMoPyd1zDJ4pZde7PegnWGk6uB9f03a4rSdFrBvu04xPvniZwC8VOtpwdkylD6PEe
dTpWtGNiTWxeGXLIVOyfZ/gIBIFpnS5BnkUJCyDzQ0td881MutA+FpGS8sVwkYtjEE8jm1x78jke
NSeNiaZimrxw7kkXp064t2MVYN+6KVYexJSP2ZyIgau4aG4yD3UmLXQySdp1pmN0R+w3ti26lFH5
G6zpEu6mbM4d71RQ4eqamapKsr9N0qa3Gl2XfJT5CNFdiXqPgB/DKNY9AlJEm18bFYPo5270SwlZ
2lPKcIEM9wIn8g4aJ0FxhG75gARLpp/LNulnFGtc6u3Y79ZoUC5cyPSelvUVj1bkc+hPjgnEPrgQ
U/d8OB9aWcZgOHLAp+W0cJhMGXXnMeGIwihBdIqgxMLMZ7QlQKpCOA7NuwpYQUU/RGz8T1JGuM6C
s1Ay6vP6gipFUlNcbzrGQPFuz1yIqeDmf11+b8OKD9nN6BreGo62+8XNAvVM2hzmnn1MJ7TvaQvC
MjQ28oYj16aDPrXy00gn7iQ3BXYZZLEOMHeR04DMHm0zkE8w+tYoj2NtxvCCZ3tUExQPVilRbplj
24PM/rJ/6YEbpW1DCG2rw5gMCzuxRCkKGYB13sA1OKiV1mWxLqqUrlon2l9GlWs5s6VNIZjL8A5Z
giicfUs5Ra5kk/GM2avxJ6uU+sf1/pT0qwGJW+ojlcPtHWMj4yY55Re53J9NN5Lk+6kmT6X+zkmn
PSzAswGXvwFGq7jWuYcU61ymThdelBbfcu++fgf9fEgB3hEUVwHxK6ti+XNTOeXQeN0jVsXWi6Mc
7N9atWjFud1hugYFda0e96lyBagrYqcW3Q1WUyRp1wqqrE94CKscU6/y8GBEs/lvnKf82OhbngeD
T2sMoudLlXqp4Ud/dnXSuoDlUY8eYbKNjepurVBVyrQiwBEO+u23q92KlHUBj71eVgojWapn5TTH
G2nzWtIIblx07KdYKV3vMFeFCnDUHEgQ1uqMEpyPWoWjDEkfRGGh5uknjZPDNwU/M1pTdivyhEnq
8R6ttM0FOIzUAo71dP6bkuDSh8SLNf/W6QvwCfouMTUluhH4winF9i3Vo+1NBN89XEBPrwKhENm9
XYOTcOnsXu1jmyTfNBF0kLrnjCoYnk3gBG/qsBa8QxYcA2quLgE9WFip+QKCmixHyhOWAeQU9W07
s/dhATmiNgFQPdt0AWKK8tasw0wIVLcbfLReKod78RFkqBMZxGQQVnvTAKK2IdkkdTAVuUWLhqT0
xsA3xit8VN6TCNCjVaxt4XPvJEEWeUa4R/S60OUjIpHCmFHa8CoDAByeWJMrAh1Hb30i8uBH+PxL
Eq0YvVzoUe7nE+iIATaMLWtAaiaQaRqJ0xJ6UFbWpFVgWSk2ePy5bhOOB3uckKlmdlAMtoi/BaS3
3uW2i6uXeUsD7NMQYfj6iUJoCUGQA+HCpYiULlM0BavCw+oncuraph9n7sHyXZpa+mlM7PcNvQzO
BaKBfZ7xjaxsYgHGx9upnaC+nEY5VFDNGkGCC1FAW8xWbscArsK7j4ZMluV+nzG/N58UP7NthyXU
9v069G9b2ySLjaJ6RLuCds0f+bcB0tfCEZ1ICU9hk1AeCqRe04WMIO/lTP7ex9DAyO3zfEyZhQ16
CX7tYNQ3RrKzVxv7RYCbSEt4boFpi5pgbNgrsR1tNjLE0WHpv9fnLxulG8JzpHWYurB12DUHfE6B
nwdxXHE+GQmnmaEOAAtbzKX3Iz43lEUPw8bbpJb05YxOzglJ96y/hEzHD4j6Gv+t8Mo4kKS4SaT9
+boRCI39HsWMnmwLdI8IyRlTDjmM4DvCvqqxAIIhQOqHMJGIWa3aM1tp5t3iZxhkxRCqjExAwy9Y
ulo1YehUSZsOVoadk+1SKhGvPirCE7VSMQlc81zi4XwK8C718jDYXB/IpyeG7urtXyOQ7oCdBTn1
O317kMuxB8VnZhK4yXR7p08iw9Apuxh1c7JPRuKF71NN7s/mZDIfnXVOlJDe7O0DX3T90zoAFllb
6lzHQpvqYdZiutUEltqfPZwODHRZO9kq5OZDcKH642Z9j8KZLPVmyz7uXXeTNRT851gadufgYCBQ
Mmg9DlXtqVZcAEkmthx9p68OmEfX1sqKFhRA3I9vEPgUR2/eKOTPzOIRhk/ChRDf7MO6vMz0IP5i
7nbnyQiGrMBLrjsUiu/QrDGBEU9zwm5aSl8R4GA9EDnQcSb9trVHeaH6i5I9PaIOoCoS7HrE7MTe
kxY83Kl7EnNNg9W/r0tMHiqYMuT0T5Ydwcx8YYS3Q87axcWQJHPP/EsdacOlFrzliR5H9IuRL2wH
vO3mPnljzbHZqjaI6ZMBW30lY5+MuzhM6edFDFh5hDcV9yq280kUo1qs+5jBf587aKjE/5rhA06t
JtRkbSYPWghTlioEvzeI9s0WGzGCTmAM46070GayPIOFz1mvnOLkcQlSkomT5fmT5y/jtTujXG3O
1TfKFIPx0fIMUmTsM8cn6AWA7zFCE5rtYkMm5cxrOtrX3gjW2jVremH/hwztq4OW1gFiDesKa5AQ
ychcQd1VKcF5k3U8dIkAOma/JQ7Kxeh0c4XEEaLLWDyAJIvPadAz7Xhvr2VpNoUomBM9G/O/Hlqr
JTDZmgDACUVTjePWe7tBNcrkewIEFuPQ6v3vN7/ogNpXEWvW6ZV+bgmHv8hFd8Vopgpk9vOLz/Mh
ayFpnZCl/KD6QQfjhbo+CnleVWcv47GFK0k5jOgs54OXt9ulN/N++1zl28204sAngCgNZyUxXO0p
lqHarw2dwZoXNzhJecebsn8C3JXJBn2F1B5p8ruK/28UcZfoAA5XYnhTuneEWqA5aymnPycLyCk7
HgTS7JVFoYws568e9anKz8LInkijWxc8NmQzsmNmzc9kcjRhN8SOfKdCoU3Klyxq5luILovOwVbN
2gpiMdk7AxkvYsCo0hRroCtBElh9XUHyxwd4H9b0dXtAR8Crtcbng58gA3ahVToTcDY4MIEGqA4X
spVQGM9eVZc2Wrmx2409QUMwRvccJj2bQ0KSuG4nsvhRn5F8nLNFCKc1D6kewdseqZWmhgD22tRs
x4QM4fNbzsOIQhAIIZIuxZGlT6bCHkwwitKsLBSZS/XZq7gf9Z6Va2Z5TBWkdtXZYsnFVosAyjBG
cEysKmbpAZz/HDbFEzkfI/8t9+NIZRa77epbIyYO8Gk3dBk+JntH0Zmo+AnUJ+kLjzshuvBmLIR6
+yMnS/phK0Haz2iUdz7Ud+6xF1yrgzBFMl1e9R69SaBbHgPVl+FAZidEys49YCan4LRXWONnGeM8
x/JuQIg5FL0nH8bX5MafBS5e7v2a8lFt7QvlTNk/Y7njK1aFhlYhNjKeKUMLHcuI8aC7kXInOKg5
2NvJa4YEdQbpyaqgHxcfIHXl+/NUFQysA3GNNWyxL81c/1m9h/RU2pym8u+ub66yMMiVVbO6bchF
3MGdGdLPCZg9bIRViRkOVOt3jQvWWBuAPKwheJfqdqKwv/dHMGLKOEdIKOGAGRu5Ax5Jw/hgLhM0
wsML/5FKhjf5M00Gdn93l4A3l/JQnlhHnP9fphhIdxlmJ2ryAOVEjMar0kMsbbxuM6zglDzj5ZIG
UBtSk5Zmbm4iLqhQzsRGCRSJd9szQynQpYq4+RdkOoq2zC+FAkLDBaXmglGxUPlXciEHBOCXynYM
mD1ZzbxnmLx7FWX/yPgE9+zLIi6Zr33OIpL+mUuKhYrpc5Hp3TIAgyZiDjrr0GjAiBgLhVogkdrU
OUm7+jsskURhuiymiQHmxfRTrAwOxjQuML+Ed7Ch5J0buwnomHKNagCaRTQIOSMkpEyoKYh0W0UQ
LJkM73AJAiO9pmpCUjYydS8wu36nA/vcJDx4hoARmhLVpO1kPlbL2jSFDLNu/HKEvpz0FV7dTpMn
y7WcjnKOD1LJ+5jqO9IQRJKYnJF40nKINrNMzghVnURVhWTIwJTZwcGrwBngS59+KOXliX1Kf1nH
gF158u8PGSzRwpVE/Csu8TM0C4sbc8dPFkyoqpWySVj2fSbB0TJ5UJVIhQUlNJMVFtSPkV5XcUo3
oLVYawi+Q6QGOO9YKw9/xyW9csblKFrdBTbzL4Apk21gBCdYlwYt0LL4NKSBe928Rvw/l70N8oH+
z6Pf4umG+eSjY4xdH1Vsflj2M7Qj5PGvnDYaXzTBwra+7cv28q8i3e6s0jZY6qgg1Wwg7sgVPhJV
6ZLoJvlTbKUiT/HSFQ8rClI6AmZQIVszSAXWRcdK3RhLusetLx2Olax6wWlqUrLorXwY6lZOwQeD
brXR2mQB+M6L8f1nAk5c6ypwE6tE5Rn9y8XuVTL/yMMlwL46zxa9RZ9bFgpZ5oxFPSv9E1eWNntz
1As0/eD7RXLtNYruGEYMtd4msC0zRv9TofABqad6nWev/EGkUgqpiSivAPb8l2x8nBlt27khYl4Q
ILywnDBsdw1t3C3qDuYCOKjaZexpkZ7XjZ1vAGETjsBprusDM698ZlloVFXxVahmPwLLLVWE0bsb
cnHKEasE2f1se0O4SxYHST2TI2/IXmCelYvu+Ys3011Q0xdKxF1EPPigObkxcFrGM8X6+PMhgB2e
ixk6iqWLv/XiKZpZGsPH7yDoBCv36Q6NrpB/bi2+RVpFyVGEhfXqmmuRcaxmeGfPLa5WbMx9ZTJ7
T/n/VfcFMUMdh51c7unKTQTw8pOM8bmew4nShWtMeVpTssjTTGOs448SbaRk9vEx94HTIAgphpFA
63thEnznvRfTWH6C2Qg9NJcT5WqTDp0BFvdXT4aCEdT57LC4BoNBtWK4iJV8k065+emJnV/ZmF+G
pWkSWYh5pQxQi+8Cy14Vgrs5yuzeMdfv67S4lmWqVG9UREIsznXyzv1Xj31SOLmCYS7ac606s3ab
0k9D2DIZ4/V7PnFsReRmyGynPHb37LmgVBLIIxgqS8bAZKlUjmSc+Y5qA26u0kTMXAqn2rtZ5DI0
oxFNw72Os0Dp5hsNnzCg7NWOuBrEn3fl5Mjojetf1DHUDM1EO3ctdQkKoWt4NKNa6KLayqSNnleE
krTQV4iXM4gLmvj08Gp6cJfyrZf4nQERz3hxSARVIOmONUM0AKvU97g1gcZjIZXhyZWNYpOGHKy4
++OotLQ9l3it4yXcJpEb+zS3CvJpcZ2L13ZJlQ3AxGmvz/1WQrcxEOiTHY3ZbnA3j3E8/SeWKn/u
Az+UMqFcYGyFUJe7ofroN3daCdd1ph/rFnJyqcnjx/U2sy4mKm13itRH2wwhxBzTAEHwuBx5DpHr
H7UWpYRlo7XiVSR6s8fiWn9fupZFAASD6fVpARIUvNPMswm9+lO8cGMllv7fqAwrwfvhDR1nzBVL
ZibbJFmrcfrH6kgX2aMqiMbE+a77+2/jkTtZesCcPvXZozVuUboxVsGSiDytFhH0N8qI2fOEbvZZ
/PVA6avPihyC3ScbwZn4U8Xk7T1sh+H+U4BSyoq6cEI2sba9GnjQaT5wTWM7TM/05VypiX3yBWiI
77mzKG8AGcXrTz7kq04ER/6FV67KSoL+aYe1QbmdpyopAnXuhGF3Y0gXSuSXDOI5UsYyVfJjiGh9
fytihJH1TP4HpNexJFNng2ch3tkN9s45oRbkIrgnnK7HkI7sxUXS67L2aPwHP8V/QBoodQf611VR
hcOH19f6ynPUDLorYIjZZ7Z+CuImleM93WlUj5xzvDY5mOA4K5qbGuV9ZKeut2CkuQvNO9XEje+A
SuIk4nzPuv0hbBFy/8Dg6qrhuRL0DucWZfTQ8kD25/3I7sHzHq8WAx+x8rs9TSsk7YL1ibgmo2yZ
Y1RnGSpi5u0hJ7etjCMRkFcdGusM6CqUANRFl5NfI3bwZuQIkF4YjsqAy3asp1QZYuGopKaQ+O5W
gIccs+usTIg8YtAtOUCId/TNY1vR7P/2Ud0gaKBfIdFCVsXz8EaNkv61ShATndKBEat/L7HqidQo
3e7OS4kT7kELmnHTpq0kgn1Wf7B/PzU3hk46G+8vqB/KSPxT+Hq4+UvV4qwE3l3cAvTSq73RHOyD
hMy9287exHHLENo2f2ApE9yx3vXKbUX2qWhsDbr70avpzt54VIFa+4kVBRJ3wj4Vaegb97tdEQWs
U4jtkQI5lEMyRCt24IQYTAgmiIjs/9TChPsuuQ+am6hjDQcQzRKscNCWz7gniaZ2P8LRklcxcHvD
6LLiAUIS7uM3m8LuaJcvw8TOeD9BGHf96RtOZ5ulMBI/9upy0+rL2BcHJO8GaKtchfx5T9u9MEiq
h1I9goj4/6N9jU1tSCojaS0L1fO+8O+oScj6qfwDn0LVs2ISiRqH7gWxgHG36IpJ/vk9MevP3+V4
a7z175tfBOjyePG3vKCZfi4bDxAl/qSe/LO98mQaW86F6jzDDlutbdrQdik/HWNOEKORzoqKplif
3a3khkMQxSv1LspikvT121vDAOxkB72DGM3QPPlZAsvxCtoWwHv6PhGUzFhyoKCOGz+80oF9E3lv
nVUFSQVYkw6cFkI/WGNZKTT8XqlCgQxQOa8n4H2+SHRiZYXck2GLq9NAdGoGnuWkTdLReLRhmrGt
uICj6Koup6AwbBUXG0qQZboEjugw9d3LBJyfiie8y7a+58j2BmhGwkdQv4bzOqxXkmzWpbBAhXnq
xpxZ1oe/awI+hPuXheGKrI8wcV5KvOvAjFrPtYmHxr48bXZzX42TSE7nh0x64Y/X/AiSmmzWVjnP
vYKH4FNDeGlUaS4P/AHgg1hQQvE/l32xG9D6hAj3xgokuWxrsEnhhXdG2Sxkple5Gj6PgI2qVTV8
/Q2JPLTUuCZah8C0laqyrkjInCslp/fFJGQM5azDBA6XOg3fBuvVJKW5+gQPsz2JYr6QWvifJT+H
Id5WNFS0i1tdV/tsl3bq6X60OisFc0Up6FXg6FwyFJK6Bm0zMA+bpRqYGkMcqVa/yK6dK6lhSZFz
vfn8UQ7bofqD0IR86/tAIw+cbrD3KM4dZm+MFvn4Wl34TDFvZ6X6Blk4TRRnDrSJirObD1pgNJYa
XK3mEIlowrIvGtruvqKfYO5rZOEjQ4QHbcrdm2Jijh98YRvZ+u7MVMoWNjN/UnrsVu4T8tj6dS2d
3VeZJCB9PhM1HeQc4pfws4W8Tyq6Gxa85vzwdicfDxdW08rI3E0qis6ZFZu7YQo1LLyUjh3WinNO
CqtOe//cYh3jP3C1oDbgiHnHzLGJa1ha+QjosSxEEend8nPCWT/9A7BYyy0LlncdXeXitkhb9VcI
rhyD3+8hoC7Jva/sUUdIKP6sWUbFnEs/kamkgb/04V2paVlSNYb36t4adMmVIHJMzQxtxTYCtynn
qj2jo9LKi957cyUpb3ucG86xT6VtUBmF9PAFWwdVUmAQMxi5FsmPXU5Tx1HtHBqsKrFBOdQpIbWK
wphtEth/5kz9JPtNw+Kso1FkMUIpBL/1UnMRrWD2/VjTGt3BlobD2W1YmnTQuHyEetau97TtnSbf
AMwtnljWb+hI1Y3uNFBrakMF/EV457iE7dxdHrLD5ka8+rAmwaG7qTTqCSS+97et+6Fv0rB4rk/9
Sq5GiSEw3QkWmvfPomHT8mr7A3FyJzgkBRFXhXgY8vDYLpL835heQp8G4k/SnSJzgSwn5ZC0rM5Y
qq4hZfVmZOAnDbc/juSL0roc+mZRRQC3LRJNpFmxwX3oRJBDRBZ0cFQlkJbYSaNPfTkCSrf/3dLf
uvsFsEJkgwOZCjE0KH3gR2RgNU/pDIFEM21bki4iuP5qVn1v14jre0IuR4awcmmNA8TismahsPGq
d/9i2OD6nM2SnXPmy4yYhr+8Cm6nWpSTph7MlDDKfdcC7doD/cwF4cDcDvWIEnU/+7blgCEsjRG0
UcYNsc/vDvgSYHVvytp8Y+z3rQgS5fzYcLcXtGuSq9ajQ5v8lJ45U3BPmHXaVCjOUl6v2EM35Iho
74KkIwY1Ec3W5GFpPB0IQzXB82chenOsLb139RRER5QrkUR5z6uovnuBGHkpE/DKSLB0mjXmmQhK
SFLhSJ3eIO0lrA8EdnQ3oEu1oXiOazDpAafF/AzidojIpHy+dmNOSUnEi9EJa2U4ASDSLPDr5+uq
eo8zBs6WhLKmQ0i89Pm98rh/qWuXVy0/W1nsC3ZYGqufUt0MGWzaNlEu/vIgevCfLrEpwhztlBJZ
HGjpovTA+Y7DHn1hTE6KLk1sAGW9Crc5CNAO7fu0mroDpWNJifYXB/bXCvMMR8ddoDAVMQVYNp/K
1abz0esUUpyy1ktEOpdphKMg66hX7w+4HuR8ek/yoLXi//gWDFRXII/ywbEPM4z27+33fiFI/3iI
FWCXZUSlrF4zoTEGAtrn1Hb5KiHtzngFZhYWTcSom+fX1o20lMQKWLP5BWX04sme6p/bCfu3ekOC
G6h6xHFD7K/Boi6MI+/QDLSRce/KbErdywPVH6tNHW8H5XXfx9Mo+ytTYSV1FG4c8wCK61nU45um
fbvjbkliPGCM4EEbNGBw5sq8x/eCv77yOCANvfXn3ilE+W+C2lH258cxskKp++fP+UNvQ6ITyzW4
zraXanSP3NRRB/VMELlNot+hM8ii5VMK4zqEdsrvgEM6wZvOFP+BvsAE76kgB+breEn1hQPlvqfL
W93xd+xesJFFzTRjOGLHAmmYEEU4TOe9mMlCRgNWftRK3mrGu0rGQ5WTM3mtPYWpMZLdpQZRdGM1
Osm90b93trRbZiHKRnO0zCCBXMKAmwdm8UKNc+A6Zzad4JkS8YYv2emR+r+JDtwIOasdYyGnrWlo
jF4nH3h7Ko3lTTWYFuqdCqtj0GbjE+SFCRz/hgBnDCcGrRbOa6t1Z2KE5tzS1wsm6r7Moil0QBEb
laWgjMiPY+x44eKN/FL1Ru0vxGVD1AqdSpQpZS/9GfomneoDgS6lZG1RLBhPbC1Khg1jTjq+mjAY
DGAJw1x0fiBytqGTQrVCOdkaS5moNAJfRXff+NQokdKeTQz6pY9PziaI3obqPOBu0CTaWj6YcG4K
MaDx9Oh8gsLf0+mBCDgNIezeg81kB8rofp/CChkevDE0mt0JF6j7XHAyV/hCqWmZKV+xbtRLnp03
zUzzcU3p9b7JyYOGL695rGcY3MF/Xg79aTH9brb1t2IaiaKsCJjW8FhEvic09RlAsVtYKXwK+efK
wqaoxdiHM9r/tZkMM3YpGnZCqjmWyfdmdJNLsxWwSWC4m3RWZC+Ow3xvE/qXflyTnBFd4AW6S5mp
QtLhDrDHaCCJ8i6m5Lsa5xAqDYKWzEFwaHQTBXn7CUTqL7axhD1v7kBwSk3woZJXSCmu4fcwWVWq
VJ6Rp4CcXQB/JZi8MSMtjJzZqCSf6lBWmE1Qhw4ISYA1zdbEQVxhfclM3xrbIiKKqckuOeh5sCXO
xIlNdzIY8VRWBbSf+WtCerK+kHol0sNcu0mEz6kbWXJYCPFRm+oaq7ucoNQEId1vOjvHROroUbB4
iEIMxuW71vw2NPXyJFkyDekDrMcs/5NLuUehsNfHxJQdgLYd4kTMd06zIo4rwJj5U9I+s1htPJsR
Fdspw++/BcxDcr4QpcIaRhJoat5oJZRasvqOlTXO9bjcHDehBZapkvbA/3r7hf0/OwmyCmM2Q0CM
9PD7iAuAZHHnkARz4FjYJN3fiN0HV0rYImS0ejhlSAFuScqUZF/kGLZmpU2pmkc/9gTxzBiqqnvr
dRZ605mvWHbmKcxYP7W7MfK9Tb2czb2/EUHNWr8VchQQutEt8o5dVdu9LASCL0KsnaATzK5G3IjQ
ncSILRLC3Hib4vdZ7J3h+XUZzBpA9FiIot4YU4FpH5rlpKALM/7IW6Tj9hNI1VQ8X2QDkZOPlc1z
BsAsNLDU2b5DhlyijUVYSBaXFWCp1ySCxfAO8yt9CcAEP6EZAQlMYNgth8GkyjT2/F68C2Jph9nd
4krTXMqc+S0dg+5bIn1h4VZbtj8ZBNFwzFC1eL2A6Ze3ZJ7CHMhOz50WRf7aDd/w8Jy43Xk1tUwy
Wg+WcmncbNidmfuSDBCTX038xFmvXs4+WpOxBeOzTGmQzYaosijI2NxA6BHIteYTpX/0j9BbXSWz
vknEtfQ9uPwR5crOKX2Iaqg7IxmVBC4/x/t+sK28KvirdW8sV0z6JAPoWyyF376hx2teTXwIvS8b
rGHR7XTtIPBNrpkE1Giqq4++8m9wbL3MHgYxz5q/37mjzDw/wr2gRYtYf5IyBUCwoyG4CLV3YSvD
bxlxnCUTTW0PdsNPg0gmZMeRFK7YpSGqGZ9H7Pfnu5u2WHOEFAqf21SnMQLHPTwMNEGLtR5bPgCZ
amnEImXhld1Rnplj5wuNoHwZdG7a5coanLABjnMAXdrOoJGvDDJvbt5dGfDMHgBOzUfKrdV2CPwx
QoBWQxZt3teziJtjtox2s1M9LkIkUMO33gWC20hkftWPGRRyQQZeDsPnAjt3hq4hXSOOC4hBisOC
xTYhpeXwyxXtWkKT9WDFQ0Lugm/BIeD3Jblly7mOrLK2gAUassY5E/nvZjF7gacrN/AyYaEmodHl
SXd4oNdoD9rWlYjamxjImn1a3yWscuTXrmc1cEXnvbinHGwCVIjpYEdQIm6hUEKBJqvJXxKrB1+V
acCRWh0ujLmhIZreOzCe+sjRN/qZr42FWf2ItAwu0L+0sOTfBx+AN2yqygsp9wYkaH0FT52gZ68U
BONMFdVGsrIDvx09XLY3SJlHQcDKR3OTxAJ6LUZADuMu2W5oVL9WD3fwfiqAYwIKyu8a7EsrHGKw
hUpKSVXcPWuapxLd2NQb4+w72WbZ+F0mZJko8NCKl/Zq3sLAkFXWA8lWDhVCovlHdqDgNcP6WIU6
gcjNs8oy1X8QrfYWKr5Tfp+mQUBQenF4h9wqMDot5KHWKv6r3TzDKcCN6vae7aGfGgqPIvfEzwht
r30qh78iQfKSZSHk/IfHIskR7nJdKDJKKS6js4usyjeT/HTyohLZGpk33Desg1yc+GWqRNZLBRwg
AKgiL392h9OFhcGXVoY7iHVXqBCb/BTqyzltNi3wCKpil3eiDkXxXyTYPKruAFYU6dHsq5snteoW
AjfA7sGpujVFeroimwOIcz1+TR7nbSmKmiaJXYrTAyA9doQjxKf+SXV7ivjKyT6ggopo+EqTSSGG
CUxLs5uxbsxtQ8Umn2/AcjSOcbUO7qSeB9V00FSBpYW+ndhPsGksASnN4BGoKd5cGKKDTMP5FgcT
BhA9kOzW41bwu/99VM7hqLeL4+wc19KNVV53N5i9JzUvGt/ytG+CK/b2ikL1Xr+GTVOnEi3OHGJQ
QYxJu4EoFzuEmkoCC1Daz2qEzamleBg7E4cpNSCOJ4H02NhpAiFcjeMrLcsgVV/rnED0yc95iRp0
gBUdqVjrc7Wt0xR5CVJwtFJFFtnExqvvkgf3PLFSnx8/NHBMLo3ID5I85/4YEBM1/FqRnLk1lHDW
H0uuH8/ClvA7a3/MgBLYLOMjcMk0CQrZ39ZOJHK8n1Ds6vmqWqWGkYAzbMCqoAINQ52Giq7D4t24
rEfYK3XK+Sb1/d799JxN8czgzelYJzM+g4F8ZMhLVE4+tjwNWFDaNh95Q4n7klQhMPYXDCa04cpN
EzfJcM2a7EGGCOkm1yRR5EWFM5U9x/IFtikarQokRxO5fKea/bfMPy4kLsRG0uj6QzYwmlynnPOC
WwHPPyeJ/Dzk2ahHksNkSLYifOtn4+9fN022lNawciUnPLuTzy+gO3zf/88BrC/G+7BsCuSpy6Tr
JmppKx7oM66vAf6ctgnnTB6PXDxUXZpb8dxh1LiXwLT+yWgC5SNO1rl/1EKlh/XxQMkUP7dsWZ9R
sGFssCFiTv/3UWFMDdesFkhI3TALmdr/zwG4mQNAeB6QevkEgsm6S6ASjvlpukSn+db3bXKO6VHO
wWQKCeaDRFOtUaGWC/UNfLlOtxFUN1bB9kFaEYhEy9u4UiBnDvRvfFrcRmpHKktNkQjeT+nc9QQK
qZ/hFw1IpC3lsE4BkIT81+bUJoBXHoGLo7l3ffXAg400IoCAMz2+bajKP7oYMh36JJgJZZN/qTZO
tQBNsPrRQ7TKbxDh4Vs1utg3NEWqSjS18oZ3DWfp81Zmxu2z3ptqbxd4DK4NankrhXNtoEzKB+Ai
kbxfCCmlf1HtxOy+PKJ2zSBEnfSgfonmsy8Bwnjbo5K3PY9ulHCHB34Ugo4EoAJlDOWV2iNI5gHw
zRYvfNNYfnROWQl8faTTO1j2S6+XK1EiECO370Enpj+Wt/1xEooVepG4bN8COAzAeCsZEcWJCvjz
G5c/g5Ii98CmqyZDJgSfl5ByhsuiWUQfFSYSdYOPcw8f48MlVr3V5TJqz+Dm5IEih9SLVGP1q2tU
rrlL5d+Q/ZzVcnXBGWv1SOQHHE+h/+mO47XCC5intoQ0RXFIo/fZuSzO0ygNQ3F5b0/elNdIYI8k
UKexAxUnf+hosBy4jPbXjhAwAyq7meGVud1aUW8HGd8DjdfUnJSeEORYaQ838DCC5B3zEqU+y/kK
RfxfXf9zZ2IZofFR6z5bk/EfAmsgSVnDWC1MKHxHtkkBuzqLlDapx2Bl5z10fwD8QcFKVs+8xYyP
yrzvV//5rYkn0GDehuUyNvylAv7uKkAnV2GdOvPtfzv4ajEdOqGnqzYadaqtTShmPxl0JQIphd3u
mbeJMIHVcp8Ee5FiPGWNVQU76AzYMSFSe7n6a1xWddsbBuI+XEJKY+N8EgSXVh11qaG/ehl/vZ/Z
szPwGiPQWa08C4cG+2qD9KpSak05Q8qQ6kpHaqKH5Z355jVTQtcdNR5Tc2kSHQxPtXEOcqclh6kv
8/2h+Ymi3uGuRXMzGApliy/2l71m2TXzD29n7JxELIyXbPUTO1D3c4+Rwl2p/JEH8Oj0kVEhpAfe
J/bZibXAqgfXaVxOyNWHlynNLHW6PQn9INwp/EunirhBkCiz9ZkWDierTzf2g0vHLCcjdGtBxZ9B
fMG8e6cXuJNa70OJr4hRBO1epBsbE7vbtOtqMP3ZCZiSKHXTPWZ2i1nqB3elBffuAVmgL6okgxRc
8zK/lScVjlpwNPe/kjlzaqxyCNymBB6BTREBbI46bGk9o5kN03s7rIUT4mDLeAmRY1wba6ndTbCG
7tmhl+Hr6bKH81QXNxzsPaEL9L7DXfqMK3zFJ5Rs1t1ykWlkY2sWm8/vFFz0AMdEfkw79J8rTlzT
2gocTsGDBiHgWchpofI9w1MFaqMbbgU1udShBudTDQi4UxdGRnVbdG+3A5u+VjvuAl0Tewx1UuH4
BJ1dIjoqTX1XUd35SruqJV9e0ZBIJ3sftdc0VDFQLfNRYkV5YQlQ10TiXeuwHNq6uWWcVOop9TPF
jy40fmmX/ebhUdg5YTsNTJeSj1bEoKPDDxX5dtfyT5x0oJXl6Qlayl6QFJihb3KRwKIashzEJIAp
kVtD8PYoLCdYCvl0PKpgBnHjsegCJRqYYOZRFZhN0fwTecxqymA9bxcznP+25dc/0FglrsGfl6lC
5hi5POYm4X5QK0qHBqXaHnBzlduj4b9ZlUTSedhuZYMfr615medIW5wFS3toq0pwA8yLV7M1u4e5
2lX3ceuv4aSOQB8XU6Z4bnWqc4hG7sPuDUutQwa43Xtli041exqhrxmYB2CNOp3ALj0LFmQsiHP1
TlrYDPevpWztYxrbnwo+o+399DCwg3DXVC7VPdFh8uLUs5e/prBkn1kJKi0Z+PW8uwx/p95F9lbB
b4NVU2vYR++8jT5fa1zTDXH1nvjDz6nCS0qcCvOuVCYB5xalM/u+1Piuq2AhYH65LXc+gBtn037n
UiDh19zCeI8CTxMkdyrNV8k0nkClngMJUKFoirvtj7Kjnxwbtjhv8UXoRkYYDQoKW7ro+bRHma17
Gml2suiE7CXP2bzUNnxnj9gSPy6NNqUD6SaB9G6UBCUCk3XNNUxHkYnbP4uzanTXVPctntjrQgfz
iMrjjxgHb6Bs9y1nSXrTCsDFMMo6X1uN6vs/BttG4HbbieHs4bSCDPVQm/QpWeIkGp0Lheg335/f
jN+ggX9sOQD9pNtZLINoI6YFJivbLvIEd/+XJjfNbgar91SEs8JEZVbbEG69050QR5jKyuv4i7gF
DGHUpRD58BRb3amcyNEfUG5EUhJA15dHiX+BfVxUHaGhzHzJM89A9C3bSlwS33XOlBlAnSa2dUbI
1ojilYf7Nydq9jqEutHu6iqK7wTpIPojoyimEHl9SP7RP23erFDTMjo2IMOqxGVnfbqXIuEM1zmC
hkpsYdhBoRzrxZzmFMmnRqEOm5A5L7yMLU4j0kG3FYT9ctY5UIjPUbsFjHpArlPHIgf8C1OcJfKW
ghhMURiICYujuBUiNDD+Hn2X03dr7bzdLM0CIWrDYQ7+zXZeCSY1EFejxshJ3dVElqPzmYYjBIg2
Xrln/k2KiW+4Gxh+RphvH4p0YF/jDMJ/206Y+NdNB2tglGfkY8VzLz1lcBrYT7cNClde2rUUTTCv
OISEarvo+uqj90iCJBcFVnIaWEsz0lZ1WLkzLoA/r5WcZrhZII4MRlqjl/k+kI4CgbFpsCnA+I7C
WGezMe4u4fjOhirpBaXdBNpjAx1k3iCmIiuNSPYNw0KdfaSW2zRo7OXc9gckdc3jmaTQWulNbBqk
P4z+P9rINEhRHrAlWWuMFu6D/7cjAyjsl/YgMEKP8vj+DmhdLGwLyzgMhapTbs2yeVWyJtgJOpi4
z5haMvqzmvFqTxwOUeDWzWpHmY3MDbr1PMO2MfKaRBg44vwc4rHp7GeYYzchz4IkqXjipAU507IW
YdPEkl847GXmp04Vqf4qXGNs83CZwtNNyjonanhWjPnvFQF6AA1MlNTE6OplFxsA7TnyKT2SBvDA
iGl1YAk=
`protect end_protected
