`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13008)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aP0B0gUaWXB16YHYdYTkHrQeeT
kByzxROgmclqf0h4i+dNw17ZHgg4lSONS85uKTmrmSH+AeVrAMTnAeRVAxyAfN5NPuWFW82kE644
IywqVXyFo+6EjcTaT9MuzpUSuPIiC1uoPJBymXXqJqXLPFIf66+E0NgglyW1yofbtINgNhR1sgx9
DeAt8JD9ezW0dwIbuBVdM7WPULLxlhRiEjVxJrWWqEe7iSi5KOvb5fzvI83hsOJKOziBELmUOamM
/T8ir8zwHa8BgpammyJqhRLzlVnk0jc0ui0l2oBOLEZatZDKIkibZ103V0P30wEv3kgy6CHZSlsx
o+2FQ+rWnn+NLza2SdRplpZXZVeaSlrNxSpEgYaaVJ1hfYU4shpw1gY2+WgUCqWSpnJ07oVnlkGj
XgvkoW7LarBgf5DSufA7OrUOvhEovDc22xsKo/6q9ikE/FrAsfq/b6I1GPuHTq4tNmNgFLJLqW0b
o15QkRHGCFSFVYp01JsJfRhVklzXE3+toKZwdGB3lL7SLiSo1jny3g5F6camzx2bFmrQu5Czeo5C
/YTWlRYi0Y0z4kUwtLuCniSOj5fXjvS+rZqv0fMbSpKDz3yNPptEql6mPHK324bJZULNhyCzaxZu
6mfclZBjFvrJ40zJfG+hWRGPBj7lEQwK9mvMkOaLF3QzB85I/PtNnp79JEkmMsrgHxSoHMgJJoNG
GeQSVZp39h6ji6XfgW1Z402TkKgSqu9DZ/p/XrxV+T9xgzoHNhQQve11khlld5aZoR2Fz0dS6DWY
htxdwg3F3n0HldhSiTENVbQCnSgvpe16MCIUhBeebBdANdreKwenIpNtmV7T3c/f+GPQpaMe0uyD
CAdVU3O6rVoXt3dusGugSMUIauBbyvk9b1/gmJUdGw420PMi+IvocYBxDF0DyTxNo84nnK+qbJ94
1vTQU0XHzhNk+/bfIO9wIOTa/xR7TnIbwelmHQ2DvCac7jth9H9aFIFV77VLdx+lJOWqki9wagmw
xd6Y0RDu6Fnko3AlZAnPA8AV/fBoS/o9Mbb9XenXcb0Gxv3pWX0F5FX3/IYEv+LqJ0x1dnqXRtJd
f3XkTKRhmAv1RHZN4Ijf/26mX+vAAf+WHJboPQj6tVKWcjoiLGqDoK25y5/n695WQznpJm0jhAyt
n3ga+4uHldOnqkP3JRRSm/A4D1m6LtnYsvrEfBKMXTTJyBxZl5SwwWtzjpQQfAmwUjmxt2oRGiwx
WQNGqkz+TTiFQ5ezlAWncaJscI0KVffI14NwBnVogLcYtDZjOXRpYxrr1uPSV4WFyXUYK4w2H515
u1OVDSE7ERA09Y3+88cM1NHWW0nuzw97Ca/B2ksxC+9UGpBq92Z62ZAfYE55Aa4zCYLfmwGVRBoE
feQhSr3J5McYr/O7r8Ns83MgdkOnLTw3Yu6yAGgxoNDOPqr31lpfWEQ6EBJJ8ymfrpl6w2iI0Pou
3Yt8LzN0Xb5Dn9kcNAAqwxEZncjIHsHGjZgKYuGELLEqeJFypgffVVzo69kF06N/3OGu0IsB+NZF
oNQ9CNZnL8ZD6tsKknOLbWTeUN78pkwcJSqYtXBgkyD9UOx8BGFgrNj4k4z+thMS4m1D1R1APj1T
J88qHzUW5a/i6Y/y1jxvgWiDQZCX0O/oRG76lZxPz4TlYHjWusiXb9KDRuPVTj1KXsjEKkQnt27m
ekgt9Y85Eg+SKoLC8QlLzPn+Jcm3krZYv0Wv7jyISxNzhIMEnrX5lGwQHMrLaX5IYgiOb6LFz6IK
ITY2vvm+uKEKRxh+aN9SdKlZF1F3I/lQJIoicGjJsI0/TY/1NH23//QzdaqgGMK9f+g4fHgMnvke
VnsKr37PDikQLBnz8VK4rdoHartXGc4nB9HSQbY05Q0EXZTEG7wXnpOXD9cG0r2pKjjTEwKlW1WK
XwBxuuNvLZY7vEMV7Iv7VPRzudJFyIsVj91zKTZ0kvtHkYK9/Jhpakiy4ooYnNPj/I9D5vYH11kY
K03oqu2tM2sNKJHOzDo12gfCZxIZYp/3Mv7bMTL6UPp1Kc41QS5EkOliFb/hBIpI598iZnnxZiFo
nswi53iePFr4IhvL4XCufFkfN3Kjf1ozXowHvE9PaNfeJyKSK3TclZgUUJB7DxEcXSrXqocyxOmJ
W0rkdt8E4XvSQ9RXnGw08moTmC4Ay/Qm1Hk4VROcz2C5M/BEbD/z3r3rCD6G+I39slabSKb3EPL3
yrBJHvH+XBU/Og2/F6Y4BGtbmBqc+F5Cbezzs97Hchh3W3YUs4BFHq2a++VcEFyHwTHgMli9VaOY
w2XwIS59gPOO1G3+YudsX73xWFwLxSGEqElr5GNcKSybx/KUKP5fuA1KtcxvUurdTXSeBDqf/vsb
KDBcshsTTQzLHqcmaC8u4PSTzQ4l7S73EUXoM9h59/9naeorj1kALVcSetLAa4LyKoKpxpfrlObn
rL7OH4Hnjr6Xt3C5YcPxh2yGykFBndcoUZYxzNUeLBqBjfYju9soiqCkwcqCDBojqq/Z+t605AzQ
PlXjKhmrcz6ds7eYwO1u4KMZFAC4HXvTNL25zDJHkxcTZzcax8gptFOxcmyBZ9nafcZZ/+cu8svY
5OGfVdRDFOlq4Y2nRCAxb5++FTVg0oNkMP67MsAoGCTGfqFHS0mrScicIetb/lC+TbNO+Wx8Nuvo
jOhSu7tAZH4FwoFNudmSrlrGXOVPDeSb95Wvl1EHIVJ/Bt+g8jHN7L3EuP3iYbeXKJNzmhruepU5
/9pGEYnfaVZv1EKuQD0tsS2tShyClZNZ02zxc1YKjbJF/98+1kndtLO0JqmeBEH4rtJUuqe7mh2q
3HpCmfwguA144Kp23ARkOQKAzTh6YE6taVcJGIZlE51FSZyJS2qaXvOUgyHmpQhhl+Qxu5eRp4CR
QgzCw2U8MoWaz4w04G4jBnldDEQkY9jZIq+iS9RwoHGYNmHbhjhRvjxbtqzpMvHb/qKjvHeLin6o
DWEUotoR4Vrbzse2tpKJagIlmH0mstt5BRRPIFMWwHml2VAoln6STdwmzqHItJ6M1wiy2xuBiMOF
jUrBgmufBslF3pAgUBsF9WfKVFnAL01FY8FVdk+WqWK8dUuwLxslJ21FehhfnaDHm/mGR+l/ZIvC
5OmSQaWH27vJT9tlaf+k50s5SF5h9+2C39bKKqW3vSiy3QerLtGmSi6jOHgLfeJPXps+f10PwsjL
fu5qe3IpeezwjDGOXOD8p2CFbqt44kw+23UtDbUfSrJ6wAs7MWNTdUpltMm4hBdW6EEu4Azr8eaE
rOo76O0rP+ct2UXu2buMDccPuOXRwDdptZvw8V6N/qk6ER21uotJk6xKN7fR/Qy19SZYyc35NF92
oMxdadmKfm9fstBbj1aQUG39cPtIBhIIGxUtI112wstvH6fdPb3Gc/7kf2XsGSSawaj3yusoei/d
aYxfLFPeRcORl1oie2nUPwgrzeGcVBicSBcOTGut38nPCyDBKgPPlqUCYDAlWL6e/O/F+eo3HJ8+
Pv8/1ZmfjG24OpCOUChEp76UToTNv66MkIZ7mi/n1fRYk0B/bs7rZytYIgOZEqlLQlqcZ+uKP7pF
gp8kYzRYgBlskLTPWHXesRRfAklL7mcfyrb+kdJwBKowSRhzpbaokwK1C7zDb1obTNbfnr2IZuMC
4Jkve0+vsuZsZDLKWVrVL4gtmEcdpo9dQ9QUnMKbIjmaUtwMQgSCsRzJJwYy9GWDRS4tPB7V/uMd
WkiXyEPITTQxDOQV5famzC1g6uwZeGRNXKKl6Xf3srI8MeJDEr24ifgrZI5RhWlgne7gfOOOHcSb
cfj5uEDoV9nUeqKBPNQCGDJKzKNK3U4UWIUQDwxcby0iUIXu7mcRrPVQ+i8ZSIkNv7uQ63qD8FJ0
0PnuAovE/oecSIx6Us1avEcX7YzKkqjLUWgs2LZOJPMD6dk8MDoMo7ysX5Sl6Tl9JF14RntPqd5i
2mOS72ZPwr9U6SOt4tavm4B/XYOdmY3LdjECmA+G+O9xhvQeiUbpMmCIQGaQ+JLdC43Nu51CMH+m
bsHsVrUO8pxdQqrRm5yGNtBFQJqdg7cWayjf2D658JcIp73SPJd2nsAV1KXVI2I2++AhSCex0spz
H0+4Xjq4I6wcBpiB9ES5IPwBRuCAU+KNF7cxUJfb9AH4MtrABYZp7EUgpGF3kkDgbIMWWy5kI8iQ
gwoif6mSiXdAR43lYDI8ydMmi1P+QqvyE1uwf57rwrXcT9XTolTEyHeathKbcF9H2e/NusWFssxn
ZAsHucSrjOtuhevUZv1j+NFO/tsWJEgQUWwHFUSHl0tSZJr21Jtv04QAXDIe9uKviuEi8M1Zye2q
VIB12DuPRPB5Y5ZTt6VJEynbZczesS1k6ndss5lIqg4YxeC3iPwEQtab/YwbJyKTlDFjJ05Z3I0a
5V+JL20SaQEidsS8+tML5OVYqOF+X5YAnPAd46ujVVHrWIUqpcTvJny9iLXWMp2puwu15oYG/J87
uOBUIg52PONeRo/2ZROHRSCXUnPQQFvIxzzNph+Jqt5ZIXMTZJMFegj5FhwuthtnL7o7o/k8Lyey
YgY+A6AeZeXkPNrO3/jyNDHcx8ngg7j4n4zOIMOsYL1Eq5h2QYgfEDCRImFX+a8vMUUFhFzlUq8Q
+YnZ/g5GghVy02e84jV91RSbdXodjfxIQtHYXE6WajRfQd9Xmc3BRk+8Uk+VlXiEv+gFdtE1jMEl
Y4J6vlUOaVEh0nfexf06/T7jVeseoM1c9nznKqaRyS5cnfLG1Xc/l4idfhct0jnfD4xyo6ztKKc7
ZoWW//Ob3qeNG3mBXNZQUJMmhE2P89DViTozT+GQTzA785Y4apmPojF8ZI66ombhB0Bej2RInX0L
Wdog3njTuUmLQllhN8s0QQIfhHteB+eIH8vSm4vihPzrjwPyRL84uuW5TibDb8uA3j2aXmJ8sARQ
ijh3bM9ltfHOSh+gdfA2CwTtjpCuJPY18zeVTbwrjKjXjO5I50Svt+1f62XsFYJ7w0IzUqVuGGKi
IQIkrQLlKPh5bBbBhVsC9dBjmkkRCGBuawHh0VgUNV1IjwtHW05jlfEyrTJWjUlntujZrtGWGc9z
VRjyV83unGC9AEscKVLm7hTcgw1Uejk7JhTYsWrmnXD/2yniLpA31qEtSZdL4A+bEwKAKbWiQxsG
COwzFFI8dfZ3qGevBY8aA47DZ5uUd0z1t0IeSunBnsNh1mnMj3oOS89PX0dRhciuDE7dbg8+0tBW
9EmHn3PKRmNL1ipXvHIIfYuYc5Od3somla8JnQyl6jBAle2+RUahuA5yMVZLiJ923n8qhGYa7t/S
dKPTiknun9P6w19cPSXpI4v02Mjg5ALkLsMe+4Y4TqElQ07w7hiHGsu7EYCQzpVovud5f/db+g1b
nI9MEUV4/hYX4rVfPm8CDe4KkNvnGMro1E0JXv57X0O0escjc2QvaFP1SNc9KVhyZLJ3lYvDXd3x
YVU8eDke68BRejyCkl7EsUFiyPvyFYF6Vb4XpEWRIiW+qCj2eTK3JY3aS5ubeehk/Df3D3xYofdw
Ps9O02/Xns/UUZj/VWl3GeoM5uK1ckObVDlRwnQlSIa8X6EKAtGbeEyKDtZ/wF9Cd9+6zByRakKG
yAZ0kiS0dH8wvu9JtejXD0Yu3vjX6UgRJprZ9GYUKRN+1KYS/OlJ7wFri824lniD6LCqZb7L0BdN
l4AQ6kM4NrXLDT427YeMNGPoE6FY5QyFuqPLdFUJ1X71o6q6ATkecmV00kaGAk2x2TwwVpfHHpTj
Kab4Xhl93ic752GhbFNJw6BBquu6DFjJEenEJKGIs/Qq5lM1W9MQ+OoHd/On8K+ThjECiWzVBpbX
19ZnKrWbyfTNu+idotUkQRkHnMZfO1oe+p4eeCIPk2f4sRaxVoz4jtahxDdZzrqbgs2lXrQ+h92Z
MJ4JqtyCA2LWlrYOiTgfV6jeJnOT7p8EqA1r5gNMMf73uzJqRhTbLYdhoqY1V9brJqIelEZGwlIV
eObr7vF2SmXqVv+D2+vRjpT9sANMCBFzg5JJXtAYiHbLFJ8WXPAhwsZkuoP/a4pQreq3LHnioRRA
NlirCIpTHWBjIlScqQefBKKuvJKIAZwO+0G5Wa9FG/eQwqM92Ugne64Czm5BwKe1nXlS4MqmO1um
I0b60Gb9nWnTtKFce6YOmmSwUB/FFOT+muekdItDqFC6AtF+AvtUQ+LxE6jEogPrV975od5PONSK
1XCKPqiO75OrG0GvVL4W+lvNsSWCkx5ezq+J+I4ba63UyxL0UJ7ASgXjyUprZVizgkZujeNC59rB
YTyaZRMVtLjriqdEgpHVnA/Mp3OaA/WJJuD4XtLIIkizKKnJpII+saXW9Tzz69ET5zQhZ2lTxjF5
bAPXtnHSYBcyt7s1Junm0aBhPpsstcrQt7A4CDyX1wRNxsrG6K64S70LNtZkzN7p/toH2QOd1Ntn
vk428QrP2w/+RDHCWuPAXKJk1GKTaYFb9o2RlxWMOf782ar2knfS5VHhd59BblwWY0nW2IA61OCo
4OxPCxRPE0HUO5Iq4wg+HMth/Anm8AdPmfHbIYvwHtItB+bqDht1Hr5pQkOydqpCJvnPvYtauzq9
rTq3A3t+nYHY1Q9lwG9WfMcGaK4de8jHn9WrrkEwVnnLj21jZlnV0ZxET7ZlY98c02e1rwVnrWr+
Je5t8HKCBYOR7JCv6DaVwvNIAoqVP51AsGin6sd9h+HhA6aVypIaWjf9tyloV/NzduLhvfjhcV66
WNNxNcgfaDRoCt8Ryd99nsYqwm1v7Tq4EtN0gtX+WoGxn4zzDoF8M3R+yb9b+7YNchfY5n5bXQFn
MCE3vBHAKjWg5uk1qBr75cAu1Qca7g5K92MfGhc+jnnTTux0rvAu8+tJ6X+Edf5DHKiflbQgiG9J
7CTAsB9Q7zkjtJcl7OcPuHTk/3LAHhWdPeIm1LX4NVzF/kt1kI5Vptuu12DpHErhezSs6YWCLAr9
6A5AUIXq46nPZDI79z+GCMgY6Do/KG9RHrttH+qyncHGFhJFIJwAGmHFyM4TXAc56a/ioJI75zBa
csW6uOhgYQo1rVjjGg0JOHgoL2hiSo1cgO8FbaYeABImPoC6h+UmyWIrHPEva8RCDqBIIxYacjF3
Sablky4HqOOqTH3Po3i1W4hePeUWVfmiHqGg+rRQvXt3I5KcOa9BHeP8PLH8WbZnHhybI90AJW4B
ghGrLgpA0BouIjoGXWb28lm9b1cn52FbIvymS/YVDidtBow6phD7ORIC7RN96opz0bgfDpBsFfKk
C1g5JN/wmgOIQ0XanlsorghXFG/y5P9M6hRDR47vsyrhrmea9/a7kEhdCuFyvPL842LMx+nKI3eS
FvJtjqUdksjTtLmVF8b8u6sqwU6UFtHtD9r3ZhLPKmoXtg9KfoRBC245DQs/EvRySHvQuseOcjXx
5RkzTTZ3jjy69kCHaFf8TsIzpmT1k2o6SeItN2z/XLhHF+cOKcMNTrOPKzOndIfCrhVvXL1vUIfY
opdi/RQbj0WYsFBlZxN22CeeLsqS/sFkzosL0tk/QrsDCAW2e5lDVZfaROYbFV2DVaBtCaPsukxr
ii6dJlm6iBgbH592u+f2mI9ze3K3bpsNH3CfLCIYDDI55iw6Qwnxg8cyeNwWyMIdLanykfH7Ju8c
ZcGGHpV0gE7uf5qc3HOBJHrSdvYc359vywTxDuP9P+SJDyx+t60gzygUEutg3fdY29j2wgp2D8A/
gRAG1SnHdPc55yCIzkndYxPE3e9z/tEfzN9bpWTkjECzzAYAeBBClkKk4paB5YWIjvLEVqoh0jfA
ZVK4BErzQihjWblDamZIenulFel5DULaJy+tH7Htt7XS99+kxeShV3OxFaxZmv2wZlozcdBjCWZ+
ibrVwA2Fw4qpfd2/mR9C8rkmZHFEyhlqgOObFsCbVRVhAPifX+s1OAHQnzvqqri2oe0KqyF8nWeY
YkcYb/hkSqPmV/mUoM9CDDcgJQ+MssByY5UZxPuSg35Rlo8SrIeat1xZbZ1y4R/59kJonl4hERMX
KzK/D2HsaS6LuWMCBBAk190mDb1DELlboatAk2U+ynZWeDcMUgeu7V2MDcR+56IG1e6MK9vMw5p5
kyb4IC0NudHIppagDkhVyqyMLYHhl4fbHjw3zJQwP5DmLffEb5u1TgBzbzxhqvOlYpBCjrIXvzo5
JSFcaTA+aXCzM3WWjZeX0dSP3MZV5gcz4e6tELgJxNQhelnifyxFrqU+OJYBo8oJUKU4sCKPafmH
2Dufn9IKryoxUA59p75/NZadSANaqUvLXoqQoRVrbKBRrK9TINJPx//uJsJ6S7btepIbmQmJw7Ui
lEkn2HbtLf7cwgdXyCjgKBL9z+onHs1P8Q78w6U33GSl3kyvbK8KJhTDTcEvB3bHQCd4qeuM4ahE
gk8UNAIAZbbTnza8Y8OhN+gGthKNYe1/+TmfuVD5AB9HbsIB8bazOCqKyifB+eGZVQtn6uB7ShIW
OdpMNUZuhaxwTq469qaRr8EjNS2xE06TFRrauI9CRpMBCBZNSFyTIssidoQWA5JVHGO6eqyXwfgB
vB2BxeV7SQGitHtabgdw08LzDXd6ctJ1tKT2OCht/xesY4Od6hO3ra+xvEGINCjT8XK1s9Q4P4u7
R0GKZ7oa3h3BylbAaJq5fKMjRqLGkXFvjWMTc6rhESpWck6m0TlmfdsXflsCxYWLEibvVDaevwsT
E+uA1UOEjCr+SWq0pClD4fxV1IqCSIwD/hgVnlpu03nhBk9PDfmrDaSeHLKm/uh4y4ogBCKQtQT1
JmW0IgNIaA13zSdQN6wD6dryxMF48Cc/THO3QtA3vl5svNKVWk+mEYu2tNApzArCa+Ifl+x58cC9
9RTOIl2fc9Gy38ArM6S39s+PeEh96xUGVCbAueyKhiO75V2yVROYvgGkC6Qi/KAqaEirBS922Zru
Ye+TY6Q4phjpf/CHGsK0WpRIwokqgkhZ14OC//k+ax0V3DhAJqQ/TcPI2ooG2EpPNdNPYrcXwXRp
9ck4cTWqITnoGg4hzs6/cxrjxIE0OhNYgLKht8zL35OZrJfHJ+KEVNCyOw/JMRpAsB7J4/54DcTW
FsvTSEABYu0I5LqKvs/BLx2tmmXjJqpjTFLA3FqNOPrrfhGkaRxQtAytJKyZibGWAgx1mzNrsrIN
+C2npOErzVY4oGBuXXV9X0qmwkQ/aU7UIyKQa90gmpax3j16L7/R/v9Do0W88WlGrCKZwOiEWfce
kh2fzKBoB+AJHxikJOg6488LLmaxBrPcA4O77GNwoOgWKufHrGUc+MJpYZhzJJ1I4O0l026xoXXo
LfGceXZT/vdoovMcrGf91X099uQQsDy8jqLLziX9f+6qIZUHx47hD4ECXJXV6QyY2lQ4h+gJiOzW
hP1yGVP5PD9jRurrtxcMEuYwQsmIPutHpbt4inFagIVxVX9BbPqyLsiSsfmKkGK5Kui7tWDDHIA0
eBmaW9Xu5hOBy1+qLvCOIPX18643fQWKajUy9kWmB+s9itfVOFuKKshtG/SnRpe5Wetoztp+kuxH
OHaxb4zGcDpebbDjrU55ej4pFpJgg38H7ljkMiGkkLGAn+TwllHeojnqM2mghE1tPG8vjPHD+CMY
uj4exjB1GU1JGByWyms9F0oRdvKliwlIQ05hpPAyMEIoiHHg9hkaOoKrQ+U5vQVga9ofIcH0BZ2L
TEFBqYxtRkqi4yYYMh5zLQ+fJEGSVs0ajiLIwoH1KKmaF1eErvEW86s3d4unJxkpkb2QxBqkebLv
JJIQglskZ6GmqiO9cPpVueo8cyP0ZXXzO1gdxrpLVKx+QPyPIwzRP/x/j6EEgh/rsVZSK81enbkK
HThbYw08GTi/RjVybS7QcsMrMB9FbuzEEAyWs5XH7NlXRTzjwB+huO/s4/BtGuaYwfvD1cXk/UWd
nqYfKzMwtaat+LQjmbPXAHvLdvRbtvSLJLWZSxVURGl8Ez0ZuIyvn35lFNZqh6I1QwAjFQ8WDl7S
9ZuT3xlLkSzxUZOUfC8QdaYV+oklrWZdkKm54M9bfeNQfeRBvylbzdEuIbgkquF02UOH9XJUquuS
Sw0qNuWzAEAK4rLchd4NfuCGNl0J+TSytnoQy/XzF5H8qSc2SQuA18fc0o9Jl0A+dm/ZfdbfMPXU
XLz5bFi3TQ3Jlc25v8IJaoN744m0G+vpEdMPPYrqHz4sXSbIDKbthpOcBfqeTkf+lAq7OG2e0MUm
XWTkWs7LMG8gLWzgi/QEryCMMmbub89tfonU2WLEzS8DyNBeXNj60RV1Xc+d0YWUXJawbOTH9xSD
sg3FK1palRgTIyTAIZm92pZlZPYnu7Roff/MBsVfIbFL+lryo+IP2H6+RyijU7aNlpC5ckqeJTOa
Lah7+s9892HqcXgQ2r3auRNlgI8Sk937dlmT68UjZdWJpi/HLmrCNTVCb+vmctVvQppEusxvG0Jy
kpI1bkdgFQnYIPzTWTODGyjCnghdoRX6ZmfSmculY9PnrF5vJGCSgOpDbZIy++PoYNN/ca9pwb+h
TXSnO9khtCRrt25rryyYrr9M+bUWr6OIr3ud8EaDfMSVCzGdNDBC/iJPfnXYTvdTC7/uWz9v1woz
pGV+m8tzkZjzBHRhDO4CeGWSR3/5H4K+KIHojAT6sCVM1j1wAXZfa0bBXCAiP/TStnZ/UputQgoS
ESPZIVRO4tMkHjNqhPLr0XwO8rmlZK4ejmOWlsYJelRZ5iKeJAKOfD6aTOhrR6Gt1rmz1r5Oe+86
JZqmDk25bLMoZZXMeFrjp81q+KwjxgnVSThF6n87/Z8Br+h7sRZZcjWKBi6UhB7e/XTroPxTNudc
ypLjHedZkWxBnpyAy7HpSv+YmOi7nVDh8opsPlwmMcnyRo87+NKEbI79LVlM/l0iO6Fcfbbm28IL
nQbzcjckRBPNb6ERDo6fOPb+NfdVhDlHNy2QeNc72nI3H+pKanVLjstwurg883OZymM6m9bYDLeX
vsRwJernuWDwDXa7KqyJHa/B/eqqMJR/1CFDdfQzfPr2GRIkx8E23sCVgfEYC8UpQUMMAdpg1nAR
ykbIzOa9QJ9c1RGx/hz0fQuUduOb/a5ltvxQRTySNojTlAdncANN7ewSXNJs2Lpp9S3d4j82cMbt
1o2k9pl3ngSxgOOp0fm1HfKjaX9kRMyDbTq7WsAGxwjV/c9nCtmsWxIVGccFSpaNqMYiusvV/0es
r1/q4Fs46kQDJWoi1uyjoDOxxhok+CLmhPVDTlI0ZZr/Y6cwnMuuhks14z/R/YocI8AkGVW+HH98
VsLZNoQIFlcN/SgbPdnaB0OsGHWOsvLUjeSVTFgi7LhtyP2x4scEDCFLfnlspPF3GjbefjIiNEov
rReMj8XKZIexeb9IQeclWRSwXowB0rP1imG+jlL+D9zOv1O8cOhqhRloK62IBi/Wyv9AkmX7EBeR
Z/8wjNay/o4TW/8RsdNOT+8ok/J9vIn5ggctes7WCP/nFkP2WAM1nABVzqyPW26FTGgOCSJ979Fk
x0toxJdlkxb3v0+7lyz1sDv23dt2MlPHqAws1fLdkuovJoKkZ1dlR2NcYCZZPhXjWgvzzwJHlOsB
8gL1IRBL+zYIREP6X3E1poTEEjOq5+tVhVW+WfQBvn6K6xJfsD64LSuwqrVkS1mkzj1TvHxBgRLh
IitT/JuCh0BbwOpt8MsdRQYSA2wJfEG5LoyQsaPpqn2B+WY+1icpU894ty+gRfAAeoIMfCrYMTC1
QY2UMBEuTUb73zaWP6Q7x62Y1YNaD9XESB/ZqWcKT5vIILi9B7TVW0E85E8Hv31PLvY892k8E4LH
huoZ7k7QPkNFdr0xNSSCxH4kgJAXcKrDZ4VTmOLFbUORZFvFEOI3nIV1LRkpvMdO56DWOh4JH78y
YGL9L9QZzbHeQ6rTMNo9CVCa2A1E4zR1SamoBYYtCyzgYKWSwI14selgW7p7Psh5CPcPlQga6rx7
VW4VzokHR07Iq4NniBqqYUCd+RzWwmALqHgpl2U+DVn+4ESKLisI20E0cY5g/ZVY6kMwIQuqWbA5
m+vnwg6f/GJp9gaLfGgh2zKsfvBeHq0XmFw6IQsZst3amWm49qs4uc0dZmuBZkmKK9aGbDnJolL+
+HL1kGBLZUO0+fJin7bYrRHIFYYoZbVYSzy4yX9TgenFG6zYnHS/l16hWZqqfSRzFjgyVwVKF/9E
MwnqImGOVyQ7J+n7uU+AAdP4VR2x3Il35Dhkh6+alwEtB1s/cSs3aiHQ1RKw82qd7N1hEs9lBkW3
BxeVyN8cfAPsmg5mWb1ljOoSb7iX64/9fwuvq13w+piUMxoRXj4bYRn11EPIg3sNkwKXyMx2KJ/J
kuzsGL9ExkUGmzH1Y9CQj2N4Oyx9zjq71VmAzX00Ej6+bzJ2aklj9tv+DnxVIyeoaGvH+3XvFMRK
X/BWsc7+QJfE3eyG9N+YkeZonu+cU3qYTNL+Bw8yamX5zgP4v0k7wXJvdZzCytHB4yLj/F0rW9jJ
arbRSAbHAjCJ6BD4z4AkWvZiZR4WnQ/KOmkMoQrdHRkVRI1QJSXEc55t5uJKmu/GhhfGWPg85J1e
lJ1J3CCFS6e9fG26WV6mYdIEsdKlIKbQjD14w8Oy3KHVczWo9VvKAH12y+g0tdLD+Ag3uOOls7iv
LQy5AizOtPdU7HV1W4NNyWMET14SXbod/LE65NMlIM6jGc8ER0lIKnUfptsVKDF02RLR1yNhn/d7
fmlnhLCRMM51bqDQvlLiMocGsFJCzKw7HBLsASom6Nd/fgRF8xvbwDH7OUsncfeuJiC7AZDAdViq
rC/oB6QwI8TA6CXGAhiI8N/xzptIZ+klEWze4ENMstSH6LlbbIKf56od4VvTTkX85X/P0xDc3Fub
daDexnB067MRkmm/eupSXI9D3OLHr2rPzD9QvGe9/w9P/iiD5p7V3K5qgVcejFTdeYoPYsNJ5bwK
HoN2SRwb6s9WEHPBNlJi+Rll4Xc4vxclzF0plhYWBZVMtDEyeGRNekfz5VariivlbvA3ZpLA2Yzj
lkjD3EIraEnwqDQqT6bBMTHD5sPvIaRuokoYdEqiaL75ZEY0ZDhy4jKACuS7prqhn60SoXMKW1xe
LsJsUCgdgKkCSe3fSGkAZdo/bK7crQ+mqvsbtjgE4CNOxy2T2ZpSnJBhTcVPvhn8W1GB+EjrHIfa
RS/P+lvWENV1PWi85odvoFPP2VWxqeNQ2lLyii9zzMmYNbMhJjF087p6IDPyNq8HwAMNgs+l6JDC
tbOGYt9kMB+czH7rbWe3xWp1yavknXF41UVkrYMYKse5LVvQtHlZJdg0gtfoaR0vCSP7s/6oeFjP
6BIJ/FSAyeLSP4ObMAo1i2124f97gbP+7pMTNSLNrLv4aZD9XOmwvtdixrMAQRZscsyTgF2h11Ue
Tzih4cjJl4bqW9gJ71sWHEdHYruSGcCbrCe2KbJA+9hTSDsJtfdXAi7m3bjL+OUQ8m8Xf9Cfss3A
NWEuU8lRIeO5VCOdZKgO4R2RB45lJ7NyUL/RafKZozgN/i8t0FX+cklls4L/vu87i8A2NgY/Ok/K
3690T9KSdZxIO6OYv25l8k0HsygockP4QhDUPForiNropyUUsbYER3yeYZUf2TYlpEagET75rRI1
2PBJSao5eRsqhbhT14V8Zv4HYxv9GdxzVHZKF86QtR9bEIsQnxZ0YTsovwVzaRWMTtUTedn5PZ8U
JZbkNq3zJUCq+n+TulivCxdBkTIsorpT7+a/+2M32u3M74kvXOoDi3emCYm9IuOFHwaGQgoMdPmt
lW8iLuKKqy/MccgXLz7JfJnxYz4JwhvY2IpupqxdlsttyuXfqS07tOCP47d4edKCH9D/W49aEMRU
/SgAFUdOIYbREO421ZjOopEfuA0eR5ygDSkQf6dGw03b3TGsVvxwnhKERefF5cUeV+Sxz1KI32WH
kcYc6zgntxT8eRDjhp6d2yWx0v/ysZzNgTgMeB7mbk10kpnB0b7h637z8iX46sfMXq0JFomI76v2
l8I646CEQatWvxmakVWdrcQ/uuVvFvBl0OfhYsbgPw+tuRiGwYgzsFjSw9pMFWJoKbvHZstD+7h4
bWH63Vkm2yzLSoks+9wPdCLqKeSvHGA6C9Q5djsKn2SOlauVuRIQyqOk0YG8tIW0Eic2zMUYCCIt
6lz12rd/usiO10p7wiIvGXidb3NLI+MwWhWAYMCUG+Mgm7APMJbbHOm77fowLz5zV/Rs/6VD4uZV
nvnxRteVagtXXCkiMD5W4InZgvq12Sj8hppvYJ7oott7UM4jff2ziOSUPdiu6nhrLpBhi6dzfLec
ot4eLfgPVkW8+xV2mWAN891ji+mc8QBINhSAPLouZJ8AyAGvO83NB6GnQM56MFpjlaYJS+4TFJ93
NTLyvmPInQyoZOajtGRhGlsgdnvEdXSPAUQ2BZTgameaBRs9LsPEh1Y43+J1uyRI6fXErGCJPg6U
9efqVgRobI3Fhgu1eItNuLOseysDprIlxIz79z8ySo+1XLmsZgKp0QFaX1Fhq0wP4t481WIgy/kj
/Z+FAPOZLJbUG8sEo0Vih91S2sql0GY4yORoVZ5zx3JHiffCeCr1tLhT4sQRlwbzY/y1xSUU/ZDN
XzUoPCRrTHxApvYqOFPT+qFZ+vi/UaAftQNDVQSBzxFA/LxopC5pJEVi2mrYlZ3oueUTx3EHOp82
b2LiDk6UPnxZH0zdPQBtr13TPjTgJfFL+FVLUvzqeOJDwko5RYaLmcGYxeVa2Gzsh3rNW1KMwvfE
c6IVV/+g5jTz/iHKpFcOWclEqqn40rAzHXQ1QNuzXzKAOicqI+KX32Irf2QVTl8178biX3+3kusr
eFOsv6836hr3DjTNf7qAkGrCk8lChd3V9iYcEOQZ7KRDykBXfpGU7Qk+8tzpU+r1cj8AQ4+w0CqA
lDlfONdv6Nk/fq/RAHmVhX0pd9fckbonJAg72zazCvO4Xn3kAZdp+2Nmc5UwjN+U3egb74FuPKGM
NdTRLPvjQwMoP9mg2dNVH5iC0QWcY3Dj2sYCg/ALXxG7HV03UFvKZ/AZKssA47IofJ+Pn2oO0oJ8
w4ylFe98xloVwyv9NESeeVPGuYr+KirBJ1ty3GkCRF2HW8tBsSz60/QeBMe4ifhzlJIMcG8FKV/z
BqXUDYpO/W5hogGEpE6s2Ti3NfXxki+jXlRWo6YVfhKkLHMH7SqCFx+c7XnrYfx9YP/DSwPcT83h
+k7Ciey0cMYNVyFtdbOG1LzIJM+5/rCq6X4w8nlT/2ExfY6kYObFismDI2oTpszqR7NiPCpD45P0
z5qRNXEDcdzbECsgK06+0jf0B4a6V5Yt2YlUklRR0IsD/51ucVvAX+yUG9X3PcyOsm05iBRlIQaY
jvd7EOa/cieRbu5dBACs/2C8EQfbzPznfYNV1mvXkXzSXC9q7KXPzzHOsug0GCgxikCMHeTXHDmX
lL24pW6pViuELSQW14IeZZxhh+28/ciZ8iJukv1vsh40gw0E4hMC/XtFUx2kW+gPrwrsT4brWrW5
imvcjRWjPCOdNe61DT8u+PvRBAdA3kGSjbHEHF/tgOfmW5EFLavF0osXZkwRbVsnEmpR1Si+ISbv
Zozo4j5GHr0uC7CyOrugIVncIAJa3AJY/vX08GlV6CxqJ6j5HbQLEpRF8XR2qKA2xhZwQMo9N0mi
2hKzfoahmkD0OjSTbJxfo7jJuODAYAbfFFb/G+5ieTbpdbqPQG/iDpl4XdBuq+J74suA0IQCxoV6
UNNdNPlwdxC0jxh/0mFkfX4poLdzkjipGkvLLWcoBhAuWUSH6ocifFwdnbwkdljh5BNvq6gHYQmO
K8nfdbpy4Eonr3+G28XxsESbTV9iSSuaWQq1imTZzbO+mqmRzOJ4GPUsgXttlFI1eQiFaKRCJvCF
T5BE5DEyHarpSPLseU4oTx1A7lmQT0WLQ9SCDRfGO19O4zSfERrpSJrO0U/4OA7EUmm47WI7aB6o
yjS4BhSJSyu0YJQKBr5dHOOJ77XAFA9bYOUROkWOtnQJ1bKYoPvTtFXkRKWzb4S8DZWysF/N375s
gsAWoSsWKLzIJ1qSBoo95UJi0moAplGlxIyw3il8rHPqc6GdqMGlTc4ZzhVFiQfep5BR0KN2l25v
L83ot/fSeYjClbRaEiVGD9YcKXTq+PYuAzHNNhv9SywOmGwHsEmMASLCYdb7uuYHqqJkYVpbyirq
YuYyBDQfOni3tDG9iRFiHImfYnygq/VjpSUSBaqH3QxZAnkzHkHf4OJmn+IsR1fqL+KwNu3f0gv0
19OlDizWlWlJ3e6fsHAvY3nPBGtNaXHX7oPtxyn8ifZMWSHnIYD/WyDPBLo82U38Z+rf8q0raLPn
gha0mKz5AGniZcghzxRzl4cs9Qh8BhtD4qPmeWujP8l9/i94T9r57T/xugHTa+xnoD4N/+sJjBB0
C2u1OIZTbKsp1UEsZtfcNrNZQuZKmI7zaSfkL2/Kytds6DAO4Jgxz7uP1AxpcDwOduZrqiCXu/ai
DnVCs6FQkKNo81nmYR5/jkX3Lq/onKY4EZguAqpAGLZnyGCkUIgmu1cAE722m7L1Vn0TZLPPVMCI
N3VmF3BW2mdpG89PK4XoX/dmQIsqQN6h7NF1VNAk8DaDr/AvzmN5xxiH1YXwbd48aP/n9QW3Exxu
ohad+9GfvHaHaNarQw+JdZQOvo/h5Py/O2sZ6ljUQKyyene+AlhFSuy82HHny8mG2Bs6gKBC0Rjh
3hdGnsrdCJOetyIxCfS5W22xEm3c71sw9ayszKSa69E+Fc9PTbyWvGw3ATi0H76drtI90UGZ/lMO
fpI14KeZxrDGAhOu9uGsz17i1mkNPhEZs6ul7EZVvqWOZsMM7kagdHCyeTwye5IMZVnmTq3Q8Xwe
4W9lMEwrY043Ne/PRNKes1kU/+ZIX9DrFtWqirH9dFEeBnuy4072kf6RmVr6SO/bo2HUso3ZQNHp
WnY6TTvUrJnoDK8ryAy8UcyOxHvfab0dN2bSkzyWHJ1xeY+kDyWgoCnNNJzH9t1o4dmN6AhC337g
jVIu8YNIa45p3DwLYeN1Fv+FSzw/hzYpZMcM3URadSuYVQkAKkomh8LZxX0D78pcjJlgndp6hehi
bDjKlV21uTrJiR5N
`protect end_protected
