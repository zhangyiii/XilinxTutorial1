`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60368)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMKRcNvzOG7grs/8lZMh3KNjoyD
IXsq0a+K7fwBVl18Zhbp+vFGx+nLviNLK4nbLGzG18UzFbO5BR1qogjKi3A7o3XP3D4SlyQp4NzY
BIfg0Ckm6k40mHO/hxlTz3yzd5DsIqyAAJK1YQ3MBFoWNFUfmjcQDlQRW7c7EnF3qlIfCCCufQJV
xdrU/NYYKMWMc8Wy0sF8f/ss1rjcdmG2n2qlgVQ8cTz5g3Fh1qWB9OgCgCK97cUf8jQUFsOQ4BEj
K2bLaGYqIzFVKV0SDLZ7RNoeIWwsx972HeP9KLLzRhy3ttGr/zTwzKnt3leIbj2IEeDYIAI0Hon5
b05UiXiKZOAkfJk22bZ4bE23JbXrF8Os73Y6jfFkJbS4rYed/rIasDupsL6eJaIPKSdIsOwvn75u
gmMOgGb2iRYBdSewNwMC9H95osRuzegWfhjqIcZFb5aM6P04HN297dBGxekvVJq/sJO5WgG7Q4li
jL2qjI9uaUfUwTKoFr3oTOdJWUrFbTuG4w1KNNCyMOwVZzHr9rfDj0hOvx1Y+vkTySiNd+z8ydG4
L+66HZjYvpH7Q0KDDEUwrx9SYq9/4/OYwL2nRMTKPGJEyyrkP3FN502i3wvknCYAA79xeGCl/GfC
j0oMZUBh0A65nFgePbupGOWlkO7xsU7ZhCskWojpIF6O4N+c8AZ4WfUuaPdisvsYB/pGFGARsb5i
p6Kg5lX9YHn8zcrH6RxHzqZCoR01Rm2shko2yBVy5bEfPsimTYYanAbo2eheMavuWhljPBdOMsmU
cXK7dVSYlh2IdS0N37zOARGDBNFKZiSh70v+wPOnAZMgOnlvw6wolkjaLBW4uPpImYULgL/bRVcp
Vnr1Fp24rMfkGp5LyXBChHxZgdKNCd+09fF8B0+MjJdbs4OGgE5p0ZOBOB2OlkW+MeHmfwbi2/wk
Vo7r3aa+N5j1h9Wdp9t13PhzFRjs8lQ0cZv/dwFgWlSxwVlReFISr3bsELsWZ9OxWgqa0lqlh/En
ioATTUn2MoUtxxn1b+1rSKMRu8Byf+TWROmH6I31MsKkGjBOduSkAcrZdfwVAYszb8Us9NXmfRH6
ju7Phj/34N9iqFb//TQruWIf0iZgBtDivYAPRWYpXdzbBAW5L+T90GOs4YQLW2qoPuIL5D5UbVk1
Pxhaua6sbzfVdWG+R/Ie6+wh1AQrxFNP5kSdhjBsHIEtX1TJ6+VC+zPT8xLG7QxxvnvCpJ8F29DX
pUs6/uPpgWBmCWdf0NWl5BBaKjCinLTyaJRCIaBY/KgDFqD872hIWpbf/4+rkaJNEEY3CizZQV/v
15ReVD+PJxQdmMcCzVbhOUGI2e54NmM7wHmRMqvXpjtwjqaKTG7vBpASGWkKnvqtC8Pi/Bdx9lHb
JV5vRE4RiQFLFksPX74Kq0CilWW0Zm+bAHodFh9+x8d9NhQja0hgrJA1ZyWRr9+iWON3rKPieVZd
T+B4zBJy0XJOmqVRUZ60u+SNPo0+YZ+8PIY996Ocf770tqYJpyBCsRaSrQTaIhrv3qK9YurtyaWH
AcQoZ1fEHkG87f+UAT5TKsQeQWARq6Z9idmf0ZP2LPU//SuWCF7pzY76NoZx4CpmpOAsP+jetOJ+
65FRoogzr7M3sMLfYqAU/V6zuLwTFWUsvZ5DVKe2TSnpOn5WboULbvwoGJiJsewMWuY372b94i9k
O4dhS1urbOq3pbY26LU/ImF6QwDYAXaYsqk8Wzxyh8XRhtQbGNo/OtgyQR2EKOyob04Q8w1X+zS0
/kJi0JH8Of+cfRrSKZYhVIdZ1hXg73c3BZJh2JnomH4sMOcNo2mRTQSx6OZXRbFSTjnR2Ew6ck2/
87oEn/uTAjIxXLzje7Xj9ELQ3tqmy3KSP8+MS8lIcLXGjf23FUXf+BwUX8BGhX5rwSxPu3ZQhDSr
cuNdPAI6GzwQDN9Mvt8epFucIyIFStQsSl8tFSlbIgkxtI9e4Pz2RlsjdTD+nkb0+X08GFW/BtCm
87hk29hTlS74ky5D8eu/Io+Xvej29vZVqomLqpXR2jarsxTbDcUobYzEv7nevX3j9Y6s+oLnbofW
sKnt7r3gJy+1ixlCsu8aKVElZVELDa/inbmg7HL4glYtGV1y+roM9J6azYubPirVC/DqxzXILwZj
kZWt9dGJfCqU//VVh3L/g8OW0zCLAIwIEIiTiiv7za6RuljEusIUbElNfXOpi2QQu7FzgD3fmpXf
twmRHBIAcSVJmYG2huira/AGR9xwZMkwHeg66FGvM5Unb4gU4LIZrIB+gZZIqY9GSdCOAnRX2XMV
9hFs00wjUslDcowZDeBxYopsDoa0OzN5hQJWuUvrUyVqX7IYbFK+kHsucfTfpxvgMBd9ezlEGot8
DQEU76g6kYQEbPEmdq1tU5n1C3d/3nAmxbtH7k/M/o3u8zNtQZakZXhXao5UQPCClVMMgKcm3Z2D
GkeemlD3XivpJYXrL3kHsfEu8KPNjhASX6UeNewMoFfHRP4xcdh+xrMopKAHwm+dI240VNx/77Uz
yMd+YvQRSZNiboNMdbjvA9rMyPi3X71Sh1ALlh7r9hMoFcsAizDxgpGG1/iPK2k1NZBzKnM9h3Im
I3kckt/WRKZY5NferGGSgaeqEanLDsHH4FZTPxJ/9MAFXZtKWM5NZw3BRr7dKD5yefC8awRTFpCG
PQVsCfm9AuHMQ5J7Bd4LHzx+UqPfAbEr0uTGhfp8QffoIy0+9Ss2Bjo1/p0tRaAra2yUwQ7seU+6
Om9LXbO+0iDOVmFvxmFEVIadD4KfTmNiq+LJ+Jz8oMjU9Lrh/EyZ7QttXJ5iO2oE0HV0OgEjzoeY
VcEuJ1mx3Zx1MIr0jSIQd58cqa2lVNb74ldfrnsWD7nNXCrRXTRJ0bCimVNQZTIwWT0eRGoA9RWw
ayBJBcDobgvmzqosZVir3WAOMObwISoKgXcKfqIqPwSGsfVKrgMR8oZ/ch1hrKYrb4iFYs3lZ0sF
DvYVQlBe629ZMhwkM+ZiR0p5uQ+xX43B0M/s1kKUeR2uLFzxTJB31LTHFJ+mU8rKbu3oBPKcOvt8
8RkCSVf06IgsI+MZ8oRJzKhI85JukcQTvp1YY4K3qGCM+pVahiKUx0hdFoIu1eTaMZGAmQlQ3M0q
nsxG4k5QDFtW8ar6n0GPpBlnn8fp36xeuIkf2GLt9EmEkQ0rVqBL/oNXh0jiXgWuEzSrHYvQJcVG
jGTsWoB73ecTtj5ShML20oIHmy21c1ftvMQNYnea6DMbFkfb8KylY86lUtAY5nmi2iiDLzg0CCHc
71UfycjwrJa08FVMcZIZrQ5YVuUqD8olR3Z3vWy6zflgKcz7M47IWLNh20vbaqE8IL53xggnKWGW
2r5ADEiaCHAEUrDrWFiHoi4Rbx3KNuTZ2HYkukYIY3evAQREMaPTNl2NeEjBdGgTtW7sgsK6rVzy
apmTenivmpESN6s9xnLdWrc6Qwc+XcaMLzQcu1KU2c3xcIaRBv0pWHCVURkpIfbCZe9MWLytO8Lj
2uoyQtilo3ofUAG0D7azOz4Fsoe+YaCsxqNynoJd6juOCE3+fG/DWz3KoE1yzZdzv74tioMwqdzB
ZZR8jOjTRb5NNBjGf1a/3cq4j8xoKAew+nBtdhWPgPRPg4ABzBd3p7kROQoBwU3GArNtBYOh+e3A
on6whWa9xJs3kr6yONlviIUpzQpcIOYB1//BXSBqeOGpgAgdxatSoogD5GAAGddL3xGhlOGei3vg
DGDWe15h8P3Zo2hdJ4aOWAZ1yxk5uyNaLprQU+Qq1Ymyn21aj9tCT9cxAIv6szIPCKOYQvnBUkIp
A99Kqd+kQ7MXIZBoVw0ghyBb3fzmuMMS06YcKk9Q128NQYqJm0RcnWKyZcQZ0Iv3QWBbnxseNvK7
iYzLPJcEmKsATOLvJL9D/2FdT+FCeUT2NDJlboOkMkjc1dqbcIIwOuz5YlnuMhY+w+e6r24kLQMD
WNGg/o2B1Au9V/yc0UAWUHGOOvHRH6q6suAfx4p/HoaWj22w1IH6LNyOcWCCTUwZPyhRbOZ8GqHA
nYmTpNdjVx4sDIn7U5SoTjfFRkAw9AvHA3n6iMeZB3fYoQ/S69y5Y7mp+lMrDqmlkybtvUOuA2kr
BHtmQZKtQ2R/607tc6QI5xMmjqMxy8GDkZcu3/dE5zAnDiaZvYjjmukbCBXX84Ra+9MKemQw3wNC
dkh4W5AQF76WlUpXQZddD3Ekhqvbj5YFbsUz4Z+xIl8SvnpCZ57JpKY8C7yvJDeFi5Jaw5fbcO9L
Hma6UGUGpeHsiFlH28v+qjsQwNnACM3NqcSvsLFroJ35wnhOkOEF7H4Znw4BY0L1ajBwbpWEJJuW
tdSgzZROqmDSCBx7crnqOckA5OzHF+G+E1FmT3FkGQW82eXSSYZadn9vtyPfcDTDhfSZ7/UA2E3G
lh+iK/AO/Ylw/swfNvjfxFdGpma3YW9ZUtGSQ4EhDhvgc1ifRXqZwBj07F6ykFxeVigeub7YQvmq
bnPSljnE0FADIXOGu6zIgS2dzVQXtxyzeBGRa6jnpLj80QKQXNsrQ0xMUs63HX8jT6OWPOqLb5Pa
mmx8W4JsIgNicE6wO+iUPU1i/OwO9KQDWEwwgIaeiKi7AMhNhQvGHH4O5chaDYAkF1Id8ILLTRZ5
U+jVGviCVp23XBONZ+oazJHO9mp+z4NlogvEiuT2+PW2j9JlbCqOMyIEbPQ1NLaJhmI/AeTxm3J+
2ef+IjZDj1CYh8pXIMTLH2TyUAIHe6E06sAFV1WNms/Wa+nZ1XvsDu64FSlPy62xoRMEMRR3wX9O
VAxNomd32Z/DET6DZAKe+1571z74oNy6U2F3Ycw5o9spEiM3FB7czs2HYLtTW57uMyeE1/NfoAmV
D/6LPoGe/94iRF/RMkKQ+fHfiRjInFR+CaXRZGKyiDYOdVkGWwBI1YQL2D+QL5oeUADb+Kqfu/oQ
nAXwObxPudL67XrapvoCzgevNRrtWYyWLlyAb5pQtk6fAv2Qv6nx/yKWXeL7So4GF5zPXqz44bXe
qt/0lvbSbNxnrvlop4qP37tnhTPGB0CWjJYpKX36RjnDBiSCO+TPtX82xprrw4OJdvtvjRi5tk3I
njym+K0MKf5YF3ou4FCtK9/ImAW01g5QdDDrSSBLLnoUkZr8HydLZKVSrV1FHSjf/S/gtgkQ8Aah
4cVg5oi7frtDgl9d/e+UmYgYVEAbZfzsIbOZxhTHbn1bCD1S2UVpiRpNAmt7//fHW35BjW4Q1FbN
Xp1nGNVgIiwTjYZWLrEmS3TAx+UgzMLj20O+OkRavNssSn7oFevV6is6uQwyo4EDeIt1YiJke3R6
nuAi2zSMG2R1Ea/GnjTXnn8SNSt9TSyRjvlr7BKQlinrRiAhpQdr8rqUwfplZe4KfObNPzOFITq1
1sx/0/OvpR9WWbAXIq+tMdHoeRTqWeVKpHiV2W0SNjpZf1c/JAyVXspNDY+TULmq7m/DV+I9EDfJ
5SdB3tM0piYGQuR0pHpn9po8BguKf4zmX0XZAFc9PQiqUwPYOVN114qDhtFzGl6e9q8AsIvHvjbb
wQX3DFPGXYNSUuDwtdS7/LQ5vihOgyocnes5jsv/gTjUgBbGv3iUxL0gzCDjVA/yqg9vw1LoVnHt
gvDaia2/aNbih8ArmoDJySikPzrb1976QkrheoSa6JWKeA++bxgo9hIY6gZaBH7YVuAKdDJOc0c2
x3UmakrxLSL+O0g6sCRtlccFlPuOJSJ/3IrWMvuOgcTJ0OT1W4TazUrHft38UFcRV93vqVP8I2Nz
bVuO6kaqjoutGUAJUdUrKZfHJbm5xKVR1JwO8aLt8u+p1T/yyjUNKN6TVtdJeY9pRd/ekADVf8Qx
QBgWNdg5NLBIydgkrNfKtdX+exWp7xeNfj89gr//evy5izcYv4ZiEhu29wJ4QXmbzqA3XgKddnbz
nmfjCC5H+GHLd2oa9qCyJFT6/T/GFbtfFTW3UZm2N/TYEai6WL81mouwZnzUFAC83St1PlFfowhE
U0lydwldGSzwz6kUzpmEaqp6kQKxPYAxkkDCEfpyhAXkDMYPtwV6a8yrZ2wmYnDdmh6eIcWFUMPQ
Jw0GtXsP7gYAgE/ouXl509VphPm8p+OI2z5QvnLc8xYYi3qELSt4m7jG7afv6D883asJEyQxmQOc
LK6Bg+nisyeNLKMfrcFR7Stykg42lR0ZVsNNnyBiPhHRDaPRT7ESyTQhicUJevKVQRvw4ejbESgx
Lbsz+5AzcpH4TybIjqKAk+cdh41i141mYWj5XG4d4goMQmncV5LglYutD+G+rcPYkw+HhbrSSXIc
F+DsdZjss8jvtbSAMpJ0V7TSk7p0vajWi6YNUe6W/+dKLpVmDn0dr4MaCJwrWzXQOLvyVe+7Tp6X
/kJ+Sp8T7kLeiB/lxLjjVCfisrautbScrVnP4H9rfen6Uxz3TDNWgOWc/P7SNH2TdBOv0vYYo/Z7
qc9UmnalgnpPuulDug3H2m0mE99m2vN7FiFI5mNISD8IF9hyEiyUYlfTietE6wDUapnK/W0QGjM+
dXiB2bl0zYrm9AO3uL5PaY4vYcpJi92jWwIMDZVdOOzFVxVhv0ZBRYtR45uN3ggnZ/s6XozCVGVi
64AND8HSlLOQazDxdXYMIyX5D1qDn1MEwhmoraG/RsfWOysFXc0q/VatBXp5uN2DSIljyce4cyfb
wUtLujIx81N2LXwj8GUZLsnV7IW2F+WEc4YN/2f2zddDg3lORY/OmMNNEwx62C5NxLpZvtbkBrqu
YshfAeVdyW2EE/xRGuOdnHvSDS2pQUDgJbCLmSgiLez4+Df6r7FeTbuo9MtfkkMb+/megpImdNMS
tR6huwi8Ws51IeO6SlJ0w4KmJIwrvl6awf04G15yEZ3sjoPGi2SKc7fKsFywqkRsnEeHWcebdxH0
DysR1H6U7o+0/3dgf2j+bsZc4MQMzvj1pIrSU5eV69ZoWUz+tOvLM1C0lr1ez2WrSCIkhcrIUugn
BQo0NBVTRYpw3b8UB2WazEbqdXrg5phidhdVkr3Kd/f6npmkZKHz2K58Bs/a8TZXl3Xgf93twR+7
anLPY5VS6o3Jnd7kJmb2Mbnhcz/sqoteNS5ZSWklQfKYRfpapDF5YmymFS/Y8dWtJFfWxDAh90T5
GKKsTeVVkjGbjGJT9ba3jnTh3QT3tqUNtQA4A6soPgSgOxTq2Oix3qm4uf6937EIKaR0R4kUm1j8
Z2K5uhfgrXYMvz8/LQJnFXCuRxhEAkc3EdwAR5bElMDqe9B06LF8f9mSeJUXXhYsApBQfDWwlqQu
vYRUZLt5hJx+0yzRUl0AZIHjQpttC2obbG2vPhVjlAb2I2cy8QkPY9/TSO7gnOktSbYN0eTjq0rK
+kNXUvuUiEsst2bItsedt0uqcWxUKRTv8kj411VG2KRIPVXhsmAi6B0FsBZxSpDH7ppzdDpCkDnl
DnoHDxErR3V2xNwXg2vxjVt/5a/cpV1hAJgOe/WU0VQBKeIGXDEVyg1tSHk8GUxm1bLJmD1v6YlA
3x63+Yi5Atx47wGBq9t+ayh4PP7Llcq5UZ7AEvleXWKyhn7sovmIZcChX7nLXzpCj8EXC13wmRl3
GJRhZbCV/polsPpYZb1hZf8J0bZLk9hvzwGic75IoDRCH2YM+BFTgf8lfYyAlQMIu7P/QR72ugiY
6c6Fu/liGkKVVEQv1ypIDtb/pO9ZI26nwqBIKMULG0mD0oS1CpLaQYFLEwVPclZUoBj43Ai0ny/C
dA8UFNT5K3+QmD4zd0ehgSjJZ2q3fUusc2u84Qgywl5Q9ADetjY1bVX+LnjKuXsLvUdBJXUkxEDA
iOPbE7njtwZjDoziQYn53Bd6DriRWT/1xd6bvBQnsEBWSNE1aU8C+z2Bhqdg+ZGtoicrXHxiUZWU
lDJAKymls7VngOoOE22T8t/Vjr9IhpfpmXVx1wdicf3vJInFZha+3Sp07G/6m8fARajVf7WPoZ7z
XFVU9+YzGUZaOEal0Rqq/EDEOtp+rcnA0bCcgfRyTlDELKEyjAaA4l37RpRxP0VhOW4quyU9yoym
KSaDauVq3poTErscZUnXguuha2UnfrwsY0wyfKZzpRnb+KN7a+z29anqhepGvRmhKwV84h6/ca98
U4iJnwuq5jTk+C5ixw/Fn6Chu7tqbgr7UMZsVXL79CVGXI3xLrsm/yMrEh8Kj3yN9qAnZAieIOOe
X23BFq23F6g8Tr50AfdfrqIMs6OR7fgZiUJXlXcqlvZxpeNU2JGyXlLv+3AhfOlPSGEan9o5K3aR
Yr5UESWZromOL0QxoywOHkaQyixdHHQS12Qmx43hK7qr6BKfuXYhRitqbPKwABPgHKRg/lvqKJMX
HVs1r/KAQwy5AoL055sQBNjPx3/+mfAqrQsnXe2/PG+Zcl4uLvJeyM8e4YAVeIixTWDHEPgJNRRS
F8QzUsKynTGk0hpuzEnC/hIOtV+ex0SIvAsMm/XD8XnwZoaOj4++xw23OVt7JMZLtozUVvUcczkZ
tV8dS56cZQYBpLVhzgjsYk4bQJ0wQ6ddcyxiB1trSjlySq3OP5g5paVNCoq3J7nx7NWrpLrXsphM
6sv+SRhRW8OkQZZ5NSTOQ80Q6FK3axT6Iba8j3LUFQ0FbzPyM8AIlZLuHBDBjC7FMkKhR9yyCORp
EwK2FQCF7mcFrWMHZV2up9oFaWVof6fuEgJdYdXFqKR3E3/OJYhXDu2I9nIEKJeEkz1GGa2Nec6m
02CI4TplBWHp0PzIiBqYuB/nNEJKe2EilXVvbq1ZIp29LjCUoAqPNzTi0toOF+XPnod0kZmFB17T
Zv4Y2LXiwfcJer30udUkSiJ+v4wEPM5/jNQglttw4SccH1ejC7tNYXw2MXOfsXC1yG9z02suDLYK
VaN1S+a2AOuBsnzF4L4EmKW/7HdBinSPBcOvKKlUXCSJ27WrU/wyY9NoZKb2xi3Q0AGJ1G7EaDgS
SFA0gxwSGIvTTlrJNr4KSbNdOFzUytQjPILijR6qEO+7dgfn3PDqb2lxWIBSlJvaKYK2M3ssdlDa
c8x6CGqmOa8y0xD70nxyRSjbZeHu8ag6afbXw/wWjFKlNy2IC7eT4FcFDbIec/9i0pEbhkChiumg
iQ2WUm++UHuQFBEMe3cDCiC25dICwkbPaXq/gTX9dtLbnpl+q1SGUdQwVZz0ZvNBhc5cf8NVrdYS
R+Nq2aqN9eeBZ2DmiU6q21EPFPboqZWKpQbFXxq773AHSmTq5cV4UeLsTL+PcBdnQke4clwVJ4gs
cISeW9bAULM3TgVnbhACswDeh9ti+InBzkuNl060yxRObGE25L/hVEGcn3y1/kFGY8j6kWq/ymAQ
VrNPAEgYaLrqpbOun4D3KV5ZTulcAANG7sjeqgRXnisLq7l4/D/wjUCjLj3Z6zU5UBYrxbSpVW9I
C/lhOcZ9WiSS4eDPq25q9OlHTDsps4cnhgJdUgl89n8hMZd1fZ91Nbu8YVQwAq3DhSS3al8kzh+8
3c7TCwYvTyCeTL+ejBwSKmPZeNZV0nJWUcvnMSaYC5A4D0Ru2zutyoYwykgK4Q4rBcidwsoIPE3x
Ptmo4JIGEcAGWgTbY//GfQSskMUmY1oJy40EoWKtrV4/MuG6GtIpliIwpgXmRc77Q7bTguP+9xsc
3Eg092ZFFudO1mxbSmbyhAl17jXm5fwEtLmU9fu4ri9z79OkNzY5nT5CzVZGloY0mY1peXfWp6Ro
jI62ceIX5NbF3lEptwFNeRqoVAkoir1hHqtQBnh/Lp69nuXeFFP4s3IV5c2gA96RJKID43PTXKUl
Z9DjCIPrLHe5XOs1d7WAUoKMeFQVu2EchJ+60sw10uClby87YAeYtVtpQhOq3FBPmFxTX2YMGyER
CxQGdpMHu/GIC8FKq4aiD3NvR8ZXnrNPmfneLUECBo5pw5RYsL5N9JUqPXXldqVJuQLe4yhPkMIX
wagXuHDGDWg7dEjRYe7RBt1qXPIdVN28XeoSKZrhtG32wWWlThmNXxIjxVN9fScPbYQxSrTlUw4I
vuB+7uklZY8tCFdlJjAVX6EVr2h8g+Qivsnh4HX3hsvumXn+6SVQ+j1IPLGXKkSEAw5rzRWCFyX7
nFBE3Z1n2/m6r3UCT4xp9yZjCeffbH3rkK8NGZP3RGC4cH/CKT+nrdRbJzibYlIaua1g3xWQ8ayU
gaAWz/5vSZUzP1UaCYPl1gf2qYnNeV4CzRcnYhpDukHWojVky7mRpcdRD1YnuElmraJZdFecmrRK
i9AnXGcJ0SIcK0HXC25TUzKKllZQk3C04abKrc5LwLu56VGkV83M9nOPalFchTViji6BLSagPoIn
6pWer4k8+FE4MpjzN6wGPDdrFciLn1MB/6X6V4FZVJqU8GYl1cxbAR0xCOxOM1IOI+waQQxKbF4c
JqlhV43D50BtpswYXtFcjAbuEnKB8BTZFuHIm1EAfsjKDsxSDVLfANvfZddtUw5sHndlZ6fp9wfi
3yCZDW1iK0wP8uEQJWqG6EJhlFogNO0KTXbeyYyL9OfvCwW+iTOuWmBmBt9SlZdrOWYlfU3p8629
WUZYMvHJcISDcZ1u2GErp1lJpVG1Wg22Ey1/DAKpFFiUPx7Ct78U1AJJbsmA58wYwq1gdqIIsnMv
y+NE01QN/RDHFSi2Q0GVBy1ZJTvESj87ErYHv0LpMNoNhISTzxBKt5jZbiI/VLimZlf0JXp/dZrt
AdS1uS9X2EDQbXLFPKEh+10ZSHNfYZ8e0dQRT1FqEmS6Z0jmgHPh5yoytCHlfmHnlyIOHh02FdM4
nqtXB97hx/Ak6fq/NJ+twfG04akJt1vRtmqN4Uh44PhpP/r10djbUQGD26irs+rAuEs3DCJYdnJm
de1W2tdNkMB77yhQ62tb0c8s2rm5W1PyhX9SlgJD34ZRqu+wxP81ef2jrvsruWUTY10yWsS4ey+F
+vYr7NuEsk35PV/5jOGMaQoHVtowsUmHEEAmi0/LIrXYpWAQ7+P4alWQdBkJksM64pdqSoSfx0Et
oBmOqV+pXDWpDWMXdWSkYbnv2R/lFK94X5lghXon2YZ05IeXxux9H1dKJ3y7n0h4CEiNJS2KtueG
n5ddk1Aq3kzZad98Gfw8V7KQEXfU7ENNyEfE9ZkuEV5o6e4onMswue0p6Odbu1QB3cwxR0ND7QSt
thCV0O3fupYV2cB+dxk0evk+39BAcr4IV0HmzkEejRZZtbE93OK6HCspGuwZQ81YVqlChAxfi4VR
EBtC9tSCzR7lZ9B23yxCfWK5oCVV7g0jH0ZoOJAxxDMMnH+klJfIgkD82hcwvtjqhjZDOJ6bb43s
eJYy6GW/DhP+BQFjUAXjimJFNpqiFxFhAwi71p/ySK6W44DSoEWNbfG/e+x66PL2X1CSjs3zXZ9b
x5Evpc7PTxOGLZ/XUSA9zgf+Gr1RkSwuocMczqD47TL0+BBuAqdXhMq8YBvSg592sxTWLE8yxPUG
wtp97F7CIBMihWpXIuQADS+SvPoNHzU7wFLk8ChlWMPV5sYmr+/oh5kjTCxm7OkZBkje5Z2V9wkW
0PiubANNus8wvuDg9VB/pq6CMOHO7i7A1t7zDbZfB5WdznepZ7/PBZfXaZYXC5vfUswzsEG2n1TT
bLnr//1VPU6O0v7i4U8164vyeuU120sZ6ZZVMfUBfJHEApICsLZj9y2c0iS0Cau44VGRHYlt2nIR
LuxfPYfZ1KpIyhc/lWSc4lCaK7yP6qUGMedK6b8w/z/E6lFuWlUOC6P96uo4jOk3T7agF5HXbTTr
iWO6Qb2pOkLEB2tcpomncEN5Iw4wSoBsVd8C5KYWXMJ+EjFHOUgtXXZuZCVs6R2oH1n55HREVgP/
FEes/qfAdnX7GdIDk1YEilrfMrigQ0rd/Um4YRfLTyFxypdFgR1uXDwCSxnxpYMShXNeHc7exuxJ
gAiUF5lP+MWYMshapodR+L9Vyf94vzkEmY/j9GAowuQNEtGLkZ1bp/5bCwONEfwfAUQmyFjrYX2v
gO4Sdazi7Tucuo3RCb8Dm3ZyzSAFmoWJVjfyAtSxzq3ujQHTKjHm0cvaB8sjTvCZYXt3xI+MXUkk
ARqYCIVt8+mBCJbc9ZYkjmU1LSsUnqcOUZmCAuL6/dH6Aotu+goihhKnr3tLJYCkCGqjOsihdxcX
qLX+xVSn34EKxUf/zGl/8QDLbGnKubTIKRLr0UjRT/q/f+uquruL3WgCgGCdneZ3z9q+afO+B699
Zlu3Q0VHcE/Gnu66Q+9ytq8Wh7aEt2Wt/+aKd+iIo3mSR98EFkpNK6AizF78t9LXDeGKFP/9SE3q
uum5Ko6gkHYBIIZCZa0Jce0n/LtdhPN7xQQgvF5BZGxTai0FKDn1hrjpEOJz18OjV2GtVu3PvIki
3KOaewxcoI5V27WNXgd6DnKS8Y0mDYEKlhBh48myqWnftTalmha09cPnQCajX5FPAwPBB7/iNsmH
42MwIdbznbrX4eNWbQ+92oT8UmIbJMUVKPQpXYNVTfQ42eUK08v6AiXInvfHJyQGx9Bb9BhTWLLc
3vXwOSXR6a7c1w+Le2NslCZVPUuTMjgiY2MBsyDpNJtIPI/tTDWpaAgJchs6sD6Lq/dxhr8UjDQw
iXiZdZWnM+exW1phLcou9W11jFSNljmuYBkGjF59v+gx6s21zDs/Lqu0P5bItzrF4uqB0Q9HsW3A
HKy1qeAD9WmKG/pXZ1pb6ZtSwYj/VnW9Rt56D/0Adekx6vcZWlhWl3hwuwY/MC4Ukzr7jnGXB5mE
ZqGmUOb/Tdj6aRR5eoXvyQCu4UZeQxgL7bjGQ+45BlQBU+vZ5DO/yO8b2Unl6aDwOPuCDwXJYIS9
OaxnkQ/MbV+7doU5PRAk9kynxHaKgs7lrMQJ2p5XepHYl1zE/CJ8Q599bTFoMvq1HqP0108JQANJ
etJT3fsplKoHl2hZkGLSQfnidlYjdWwuy4sLRBRLMlK9JkCcDJjZSur7KyggCSW8Pr7p4Wot6Y6s
j77AwU95ukUQEmnZlSighpROMbQuN9G1RdGzRHIpdWYiQT5MC3fsUu6Ncz1NDXi47onyJ80JrEvP
jPWN2yFa2BSpog0eOuVPtTnDz/W8HxWkyg3rTyI8TFdvbsA2ckKYOQc1EdDMzByixvA9oPiVKT2g
6xS1xdisx3gK725VQBHtASmBYnMoKVstD4wud0wMkJGXG1MenZ6h2XE6um6U7WdSrn2S0Jr6chNO
bgLCL0PL8+HRoPs6HIqwLC6yo0IpKNJWH6sV3Aqlh9ZnhGRtNwNgur176MYD43ZMSACOHibNY/4w
d3qs89cB6xU3sjW9i8tfDflVumyXk1zTFMcfuchVZ8Hbs1itLUJo/X7Uic/WUwYNKUj34lew4nP7
lG4JRBp7AMSiVY3K7KYWtV/QFomkkdLFNWnbPODKjFtbPENckBLGssG3Isa+9/vR+BpRgZ0JP6MD
wcbgM2PspHyNqtuGAXHzHNqlYo+nQTddqz35kjZxBDkl1xifYdfiFq80G/72O27VNv1ZVLvl7PLZ
zBufT1ZI5MeyuMF5S6AFz8Kb4Jk2DIUOfpcnf1PhfRqYLXKrsk2o1EhJTIoYqIWZBhDchD4UN5+v
WlZjES611ndyDS9r75jLw01MEfeBJ/pBYJST2CVdq8wrtAD250nL/YfIJtfFT2C2CfIFQnmd9084
3yTMhXvmJ4BisKEN+6gUE349PKwtvHxnpTmvtRcuyDpdF5L7W8FYhbRAJSS1D5NOqR8PFyrXiU1T
1AQIAFHCEwq0EYcfTLpRuOkJwPoZWZb3mQ4T4HQ/Q65G3C30R58UZ5h7spjS2QHtPRhBdY6TPQ2p
ZNTeRYpfwWidUcY420uQSVD3+7BuOz1vN2rs0OyhQTNBzJIW3aVqdmm1zljT7wItJFEuTOsWy3Cn
xVlL3lCG+OxKt2aNuTol4AQfLjL6a4fGxWcy1UVA+bqlP2na6X5X8fTzSCU5Oh3K4cGO80dWDZp8
OTsph8JUEMfDpKCmZXkB9K56ZdmSHwRhFPjOIG12vZkYF/qp/NMvamtfQTqGOMignzMAXAcmgMai
m7KeJNTNFxxt/Y7jqpJwwmGW14FVqx6UPLHn2dSSJaONdSpYK4ID88hIa4OGZ7G3P2WJsUvpDWfU
DzQMT+QL78Q0kgUT03mY4Vzpv26a6BH+BNHDbLbAR6/8ML2kALMaE/BEn/HW4vsvyoBCoY1frv0T
8g3pGABW41T+yuBmN/Yj0GPu8gujc5FmZzV1yb9K/k1LXhHUZXgSZkgXT9o+tmajeFyncHcvaZcH
QFLrHsqYUzTTrDUTnmGBMAiBjgVdm7YQWaObNil8oLGORM0SndHSsryrxF96yDcME08n87Hq5ety
ALqQ3BGGeftA4GeDcBHnDt6Ckxyo4qGE7wHf7CgL3LIIp9fJe9pRzMxIhERUefzSBJ9AaQLDTbiw
uEccrDuL2eWNGRMTvmTW3s3119XveDqTlURsuOY1CBtsF/qq+7ke3W0lDEyq4JtIwur8NCQFE2B7
e9U7Y17nNSqeJK5TA921yN1DtdPGjlI+qjOANFYBMDQUwe85C7mnraUSSQI5vRfp2EtI0Op9i9tw
3PExjQubkbpK3iPncJmQVofHJn+lIhxoQgTnESRaYV0EdaiI0iQDknYoDa9yir+aIj0wjkps1phr
qVVBtAbSDR1hGwXSWo4nIJmBMzGRy1QOXDIPERu3MBu8uHZiw7aTCs67zO/ndUtD7iMhdnrKtqjo
UiFKh/z/GxNSKYWRY/RzisN6dh/meHk1M7zbjzAQg4qNuijqPSZoOYG6zaGXmrI8wWT9/cDCb7aU
YEc0zr7PBcedXq9Q1K1VPp3nqHngA06WP1f2n6Um7xR/K2PKYK9d+zcIZ+ZJJTJneTC3Q24Xxjvn
2fLyfgZLyihcKXPG+jjpkKrfUKvw5LwV0QhXq6M7ZMhChgWsmMkjhg8hz+I/Laq03AoyeWt1mkIP
dCdfN3JVTPzb0mrrkpnfeibnSKeoZjh43q1k57mt687aGdofyvzwCzQFgDbwN+BNKqBBZBQPUR8J
0b1YQDS9XbZDY7FTRZM+eKGHCYdT4TPy2oDASyOVd0xSATip6DsE+KEcZ0IEfbE/8WVvmo2nqZco
3ByWRoYg99lwpnC9N2U3SGV+/pe0EPDiuw8srd5W5VUqPLpTceTIWHNdLXU7rUnGxV53mAN4+6VP
Kr4R1KWg7C6nVCkh2A+OhKH9m7iMzqEfcejHbItesU/dazf6UxdwU9SHBEx8gm+fvhL9EewSZwNN
RwZS7sYcg9Ymm8rFMsPmshR82x404X6OUsmHA+iSn48yR6Rom5jtqNPDczPPBxNt7kLmDBD3fzb+
9IOpGx/YhxzU25dsmwjpDTMf8QQ29TG3rMP9Zi2nHHztBCKsgGaPrdfel1p08L6YQM2fqM5AycGs
1tTjiCDeuTUqlSSSgx5o2HrF/WU0MbMO4PAjQ4iHv+8KF3lmkK+PhaK95lP/3OBniBmct/gLbte+
pmCSy6LUhRKehP6a16S3HN6PtOljhbzpuqk+Rn3lUwNi7t70/TG1i2FiW3lEfOUAXjh5K0JsuOET
9EiGdkPNoI/xL4v7iAFzE7wAzjXQfUAfy2MZkFZi6jq1koyNScr88h4qL2OrGz7/hEongb6rhSzk
Snf/FjcAqYlWjxT2J/b8z5TVQkQu6SzHK4oiWoTm0bV+0aZZF46EiXmH76Wj0KEdja+/hgsk18AH
u3LhIRlVBS8u1nAuAxOnnpF8ncGwsepWbdP2ZcQmyVQ9zvFaKrDlgC1lJFlXRAx58yum6zKBKGIj
2Ue27APh1/Ddp9psDc2AHPutPTGaSiYqR5e5zdt/A+MOr89jYTtLZtZMtAj2EGjuBjOZFttu8BJL
+lenWDN0XR9C76PjjO3OPQRhpxIUFmX/mC49xjQyV+c7T3tBRxuLja6fiP88NXLJyAFQgw8Itkh5
N3+SqQ3uScQULrhEujoDduGYWsZjEzUmK4cix0r3Db0MmEOHhKlXu6+a7gT9znisspyC1qmsDQKo
AXEgYtnRytQWkDuTTQW1rv918/iLNBTPaOrZDeSvs0GMRonDq45H5PyA7xXEzBIAMPYfO0upFvKX
MlSUK30EHGzqNx6GcH4HQQB01R7DF6orc3xFRpOgLHGsXtJLxGc5LGzlo8PoBRNlHMhb7cK779WN
8aHnoPKrTQuqrw6t2oINUJOVuBXtheO4mpQ0kItvABixnhZexILMKjEBu2B+t3Y2BqTYhva+DzTg
tC+nC/NBh1DbjA5iRBvBEiA1C0LSz7WstAtX52XRjIjPK64RCekCpItTfXe6Y6KQVnqUTZ0Lx3kI
gQTLA5VPgULtxiv5Mslp2dMzYKZ2JWlVj/lfbzwFm6Ct5+QD80/TkAAGinfNuSR/NRSXWmmtph+g
HvFABgHRAikEw/eq1D0d7UAwa88IPRSjBXfrR7PRZfSZUws55aXueA/gjfPVer8WeywNP+Q0Upbm
hO5Z5kC+tm7bMY2STvocYWg5hkIgbvW5D0SUYPK6Ywfijt1nMez1QsYdyp+9VSM38mYNNhGM9Z6b
tLupijNK/dLAh1WLW8dykJfulEUD3aJ9TwZIUinNn48G/kneSS6ke7yJ9CT+DhUkW4BdSSI0eY0m
bG1LNBsxsMfMxybftp0N2eKuo/jz/dbKv/tpIU74BK9e21tPLxJj1DEOwpHxaACQQTRriSg19FVt
02OlVGDQv9DWjqR1ljwW/VXQtOY18hfj9iq92tAlW25pbH45IL7zn2fjAl58g9TyipRwk/b7PsG3
M2OftMtCSCUQB+AbQGb/qNMuuYGHg0kVevekglbbMJudqlSSMPEFb7tUJ5zfWtCizZoWQ++ldgxY
WTToPzsXUxs1reaLzJTpPK+gfJGKhaq9wtPQtv9/zu2NPJHYU2ZsXRwkdQG6m9Nfk9mpPZ0rST/Z
yl9IHsOBKHyiqu438Ytny5s+l8OMzC4GSqvUFkOclMIpKMRLhCldyyqDVNq1JXs2asNHePrtvzdy
9UTNrCmxedBSXJKz3HP/9B7r3OhkRpXWeDGzxpTZhugOPOS5owmiLKPjRX8Q2KajW97gejwOWHnA
+7F3mO7cmm7kp3VosxoYPY/7ckWkfw5ZPndvhkuI7Evl0hr7fwoJuGYLb3/ym95qEyhVNwNtTC7o
zjd+l5vwDarRiOH1D5E2cvzt8/c3xlX0JQeoxKWEtSj9No/Y7IitwzsA1Y7DZeYTV0MSqzbrl3om
dy0zeOfwgp24V7fXR645QN0ou9dNzdSFdrMbJohFPBkX5Hyns4udB2plPCyb5AJG8jX2uGbIuIKq
axEo9Pq0H5wInxuCBmj39lJMECpEZHtv+K5B+Izq5/kJ/Vb/r0Svt/M+UFDsh3GFFzGiq+n17cGO
3eZTCQw0J2h5a6ExgM99qAXofshXrR84M9fwf4PHPuH9v4iSkrxPT80ojPDMVv/R9iBVNS392OZW
wNvalHVTz7DxsM1Go08gwBQbTCNAttMYieuITLac6wxAOVZXFTu69rmWHHKIETJfeAChAFCUQW4V
urfdDzrapVGUjn2m6+y8Hjo18McVBJwbq2GB+v84oja+MDyLKjCMkNYPtpCIHDcG8Zdefchfmjdj
Fa5c2PT//+4kvi3o7LAI9wSNehDn6rvRPRwIiC06afNBYYpwh4g4bOf8+OwqrqGxz53UrMrMP3OC
zRp+V5OSKJwpnOLnrWCrHg8I9JvjjaCW4gILooEQD2eDzb0EguoxUP+C7jm5IDxKiO2J1MWqLuYW
Mbxz5usTDMRI/t9ucvR/FHoJ4jvsCTH7tEQiP02QItzQxhXhLZjkmTWUkwG/h2e49UbHNPToIqzE
E2jmREnykV+j7J6mVcxiRymVcTaTTdYPfMBk7hX3AhRCkBSUXwkadN5rO73vLqlW7dJ54WStdhgK
1yScDXACNo5MyGKd9ST3k0Kf0scq77fQ/ItVr1M6d736GFMmxre79psjvpC5oRjl4HPEyeugnCVw
iHsaK3EZsQA9lwVZO77/vnV7Uhg8aOAqI1SusiTq3fV9cQUENof0Knr378i8Phfjw09oqLimMXMv
Ss34ic+SsV7aVWvffgafADbSlPLpM6KCXUEElr6IQAct2HxWVr8RRCy/BjmjsZZWeVn2lUatI8U5
EjGgFKEyzS9AT13RVQJ38Tt75TChhbXmBIxA/NFuimQaxrwTnjZ+VZkLKay4/pSx0f5O1J+RkoD9
JR9+T0BcUmyEDPrR8BuESBjaN4s7Ald0OJFHneilKzhv+leYLMTuZwFYAxMm/SdoabPNy4rSVFHp
VTiSHb36y8e/aDxgFyXiAaBT9y5GBe/K68FtlDI3VG055/dseepBlZB1Ujz3mmITyjQ7yjRg3rTJ
ZDemAU5GnmuIAjF3erVjxCtBf1D61q7mi+IWbXWG/bSBThaCaV0ggVF7uInJgxFIFzGPAVh1pP8c
kfwF20wDcjJxtBiBDUwlRdqjDE+aGahlOqOMe1WYgj18p+phtlAPh35AEojHEDMg+pjJNlh/DmpO
Oglmw7+kp8d9KxpjCpjPgu1MglJkM54Anpg0wESeutSov+Kiyto6zY3Uj4cLT0OHpnjq9hTs+kT7
Ovhw27D9/t5E9UXAh4fwDGTYnUol51zA6kK4aOd5PgOT5zwZ2w/xCwZaKbbIm45ZPBFJ9myvvUmM
UxQ9MysYCHeGjnau02209TWhIoWhCI8b5NhfAEGKVU0gSkFRHf0pYJk2a/xVp5I4R52tkZWYc+l0
OH12786Fk/I1tEVNd2UQtqM5XsH8dKEc9ROU3QSwn/s3hIVotBiXqJqFM/c6W85iCO7AFVyID14g
2pK1gubRflj4C+vIBmKhesZMSNf6uJXwAREvqgfsEuqD8lajSfbXyx9MA7YnWoJqGMvWebPHA2ME
V+1z7FIthZIN+ZCZXPOQOJVSx/VdX+74/XfC6S/pxKog/iuHl20ECwZ8p7npFTYAV+pijkw5QlGC
yfeY272XnuSEpCF37s3QyZ6d3db9zVqfW8aVw7hwKCHiSuBIcnhHiV2xhzQtH64xAS5l8DkgEyie
SNLDU4odEz9Oga1BgW0tct8mJow8EKieH8X8jP6MrwLAjcpWnofVTn6j2ohhWJM8R9VHsa4oVF2d
8jD0hkDrYvw8Dw2hn/HMylVxmclyZ3IGPAUnOesTkPKI+ti9vwvgJQRVN1+VsOZUP9ccgpN0SWpn
zCx1TacoWChQtLA6Q2IucVpiyR0E95Njz6vBuJ70F2ed3TegnuqRuHiUGvDO42UlGEFQXg9lSsQc
rljUEfmkzMV9ZszcomQC51NDBmqn/Sn366NjjZ9UgYoUlIv6PLVFN1W/CdJOfmpL3nv7NJ2uyqsi
GuF0TXSUNGV9lhONlk/qQmLztAWdYIJ4VCgy6rOz1GgFmz/EBtbtBgRMn+o4/TbFq8DOWrotSJm/
AtvFGZ2oUd9E7uP23/ljjNTIZHVa69OKFC/deIl3NyCo7v4FZvFoEJn0+VaspVFh8avMVjuFhVN/
e02+vHMLM2nLaqckgj/JvxHGVTaLONe+j+0EbHcuASySI6O4hccZKdpZAclce4CEJ5WHyR3MRi8Y
0NsCqcMb/NmUTc2ADdvx96R78hLXu8iY3TX+P0rjqkG9e2gdrqLwv1Xrhu7nxJGjSeyOHVBr0ioN
x0QqAjvHkje04u0nCr2aVYXpXfqG29ijiYcIYhStsbSLKXbaQisBgZpw2jfThH8kLw65Cwl/FKDa
bO99Th1mkmHDvvHu1s0S95lJBAAM5/8/d/MsvkdseCphkY2ddN3U8dT+cf5nPP2ccAZgAc0nPnfa
GiVSbpC/ErORPGAef5XkWIbVCbasIumqrAqdMlj2FGIrjVAvzy26Njwyx8oTo5+QROnJ5RgKm+3Y
WGWkdu/4aBBwH47aSUzOlFeh3fOQGUlEGfDb3tnlvu/qaTEON1UIqXM52xzxrp6FAt/G/P0HZFuK
LRX0XhLHOqTAb5Id42qPwQBpGyhdIwIAG/DDN1YAPXGK4JLWSe25QewtkUSWwdjjZdlS7E3JKpgA
VGGi/1v7x8PPfHcj8wN0qKBCezONAr8t1UjzTald8u9D2imRsJJ/Lz4vHZ2qJ6qC+Ju3FpnL5+8s
hnvVB+oZVw8R9kse4ksiSl9zWr7LtaowAXI1azCAzA9Ry3QVPt2N1uiB5i7FYwr5kWHJ/iNa3o2j
k3BawuiFipO4x5hv5lKFpuahPZxfEyYcuibXJTF+HktKgzWTWQubUJEngxWyfXmdDuQJGiXKGKsN
9sOFWxKEDKWvFyh2WwwE61+wAyUqkhA0PWKdHnx5KTqweC6hqTyDTkaxai3rC2dNXfA7xnG1cLYa
gZu4vet9t4bGzQwsE0LJNoGiYCqJy7/6BPMxTzpF1nF1t4S5YvgrHeckpsriPWxDh+sMFH1SFxoM
vu9w1mL1z1iMviEK9FhHyyl1N8+F6Q5+kO/O7tpk7pUyGy9JkuSar3av3YSDfYmKbfU+9F3I5yPi
hNWsqX5Yr53uELOIyexOqIEddQjJoYYKJQLowfOMJN9EmJSikLMECmKy3/GaFyV6TOn6Z/cHWi0S
/cH25WlJeHL4LnISgjSDMEG0+kajM8r+t1J1ekhSisAx0MkhFSiLHITeKhd3B85NJfGkeFpnltQN
rxLwdu7D0GWYkVMjNXghb/XxQG8dI3oSIwHjLxEdpbNs5SAP3NX3ibJBkxSgWA2T8UZeaVG6AYPQ
zGOJkW2hl8As7GJcoXUPJlWbdgaulpZMoOV7WKmSvGtETix2u0CNm8t0tf9AD/eymLoSELkfoKgp
52vBYgo3QF6l7PP0fNaXj78q9C/sMZ/0XA6Z16Q6Z14CPS7UnUxsBcSnZt8j1jckNbnIZFEbVZg7
4jq2gcLV/D2cHNUJmE0RuLmAPZVU3gYI+GbOJMQGGPjRgG3gbxKZFZlpkd+gpfnMUdubk44hoMwB
Z96hGQsHa7peOVO2RRlz8tEH4zQm7DFL95DLSExlLgWubL8i2TL0/ibKX471xdGz4avjc7OwoyGr
eP1hj3eZ37Bt+qxDbs2SUS3bo7CiKOfjDIU6uzOLw88eOs8Cpa+l3rl2fyVD97GpDg7m0L2WcOzo
K8MWMPgs3v5YzeGkKFo+Db0F+UtCb4r8HnkgdvDY9t7SniXKnvQWzJV6gAKpZUmbsJKO0JM8F0pT
zxH6wdHlaEo3NuwnhDt5CMdLw6W2Z3RMdAI6qys+DoCu2VBB87VFz7dPqyT2a4/dpM2dFflYKvIq
Z7kZRgn0ThQaIcTm1315KBIVGesf5dRmtiCvUGMM6Eg9oC34g/p39Zm1LdJLRAjP9Gm9PRooAq9E
8WAVhBo1T39tlzLdUF8gqKDTTd2vwf8339K16DWWOMgs9WSr9T4DZM8S7uPB2OvF8lXqY9Frhcyq
Dw/ZStQeYGuR+t6AMnuy28ZksFB6NMeVEvUISBkUyVBVeXPWVrLqFRw73sgKrvZ4LyKJODfWhROe
tDnGfgpXODX10vEWGlmLS4Qa/utjl0arsUhJOvSJuRB/hZXIQfE888gAhvMCcpYMFRumnArByShn
oRbp5XY4k3ODN2D+ZLHCOS/0Jnxw2sbiZYVhS4+YVxDJXYbPQVAf3wBmeNNfv+rXvmRjo/E0CRT9
2uxQoVBhVZ59sF8qnrnpmkKoi0tlRBB23Y1LuITcaG0GOD+e7M0D/qCLkJxCEA48e8aSi/0js7qB
6qLf8rgYUY0jgs8+h6xYFBYKjL/eMw5S2BkSI6FYaNQhe0R05/agX3RCTmlgS42w4H1LtxvFOvRu
0llmqj6kusHw+58ukmqhFtKaZxyHbokXNFZylfkvNUuzTsm+6Su0+XNDNKeYCmVKq1yi6v5UWtXB
fFYyGnySc1CDR4y8l+aais0d07rGoTjQUnmpDUg8XsZme0xE9BUCUU3CwS0CwOyfQpys79Ab0EJi
vqmXSkMKb/sWhwZqU8QE34XBT/LX2/JWShQ6p+1036vLUOQmdmt9Arr4fUKqhGPp3DpCohwVH6dZ
M75kkz54WyTyAtk4HilUiRaxX+94eHNeYMafirxKQS0y4mph12myd9jK6wPPAnpfCiyvHYFoOO2t
LPl0+fUwYSy9t35SD6hWXV2QcbqhBvDJjJnvIOlBAckg4T04PAOS1qdeWEoYX05mrSIXVud2xTyR
gFaZQk1x6noPIOv5JcVpcIjDEjm1crdlqwZ4OmBsP9zRfmtQlbvPW/0ZxGpjY2pFgbR+8l1BZZ/e
u7swHJ/8qfOQZm6APYu6+vukQzbQUa56ikXkayTOw9BU4ho0uzI2pQhWAEmuP08/1SB6OCL26O7M
QysQUxUzHmnruFQbxrEQaxDaUNjDAdnQK1Y3eqFnWI0ZzFxBjqhom6HAqFZTSuu1GsgDc+5VZmk1
mNpywlcCVY9rErjPFGeXo7wdNnUZT2xtlqo7DFzj2wteMRxqRwTfozeY7w3msdvElOZDVz2bWue4
z3futOmXq1eC5n4lulGPupjC0bcmtVDkPsi9+hf+bZFUdxKTmPGjvBThzOwLx0lNskBVOwK+xn3+
FsjroAZFsgD0+rADXEPXO5dzYlcTl5D1Ry5zwEgPX/f8SARRHKfFb2dbZa/76Kle6OqPSOt3+qJf
z/3M208ZC5RLQUvzx3DXBWLkuKMczSAo31xFR2sUa+TSVISKhEGzciNSi99M1DhLBlM/b+HZDX2T
yKpK+aM/nbiMLcS9so3LJzgCrX/tE3FddH6oWxsBD1be+x8ETnUIbJxJz2NWmxWy+xAJ7hZZmTLC
lcgdpK7ZfDtsM916P05Qti0UEkhGCfa51wuKQSjbyU58hYF4b9gjAk4C6K9v50r+b3XaaS7GpYaV
eGZjxCIz8u6qsT/T32Mo2Z216upl6EgGq/WniLK163iLwNyVtN7cXcL/FrWq3hRio9dFQdPv25lb
mW2F8Lf3ZYev9iX7RTl/iSuFH3zax0j15J0vxLRg72SNfEYLZzvTF9iiXzRNhetpRRoYtFEQcem6
XJzAbeBFp/RWO2DwGzZum5+cRVFNPMNmk5encZwPz6W30Ux/U4PY7AKWouviPdfdJErnYoEz2hQM
XdpqkaP7+42XafKe+BwWRmonfabzl4JReVNRthgTG6W4Xm20CQ8olDRCarFg/MmXChk+HqMG1XvI
K+YNXjYMbyN5LGZSUsb3IT97C627r8TEgr5bcS1OcehD9P6lFYHkYJVebbyW8mCRDPjZ79HdHuu0
lmEzb7tn1yhEdyFbPklrOuQgfJSLEL/MkzhlDh+oSP3G/gpwyueVv/5YsrSEDIefGvV7rgphgT1t
FVhEP9l5Z+n/7DRy2HQFccf79mXvqT9KwPMNcAA974qKqq+0BvHLF8sHYxn4Z1gDReeRfU88vjnS
fRK05WB6i7d2iweGDxqqLE2CzZ7ByDhbdwV3BvLxi4EwLxH7BBkZ2Tg7Cgb/7cHoDNyiNkWd3+yx
kQa5UfjY5PaaLlzIW827RkJznQD1QgE4QC5Qq15vSmCH0HZFqRz8RWk5Ciqjqkn0xjlveA3JaxB1
fJ2bqCZIjtyMv1b1ysPREHYAPYn3bJ+AZH3LwefJUmzfsQ6cJIZXtL5hFztONihJTCdSz+lmpnmI
zw23bvuFvUZ29WJsXUZPPWtURdd4uOD3cwKbfmd0WlIN6pfqFZIM3kkw7trdTXt+XCpUS2vwKQ/q
mSPH2pqd59WfyNODPj1Wm/pu/9EgUe567czZqZvwOnf8olm+f/D0vQvjuJHjfecclLV3paquRndk
QMPsKbEy4ozWZw5mvjNFxHy0ENuqurpcMrRanjHpF3ttcUj9bao/TPYCXVokAjULfUhAuEi1Vn1d
BaLB5WM/1YarfOtJBNs2WQTr9nMAc6jx7/KJJk1i/BgFvkx7s3CcvcgdPtZVQ5DJ9n1AC6makSZC
n3cSkDkNKG+CPpxeB/xm1zchpO4BFgkr/vDB/SBudx3uSc/rUMOklfGuLr+RFrecSUxT7cH+pK5l
rzd0mIrSyxt5tbPWpND00nKS1g3+idheLj8VHdWVxAepwH9llBuJXGZWRynVfd35Sqc6KV0qVH8k
MoWa6bFqqDbpVzOUFMEpMieJSUFutBo3maqXhnDcOQJLHme2a2JH2tzLdKXf6ZRsmWxnhIGiOXE5
FKxtE9nFcGlmbzuH4MGunQDtVASfD0gGHXZ9rsZz3aN9em6NRwjiRRcIJdPrf/MjDF6z7rwhrvOT
zNogKQk85YKrObhdKJ0RQVPAUxrAHlDivTP+zmf2GlhskpvSYgP4I0SiaSkHG3JAWuMuy7L7DLxq
bFkQhSzED+iD2ck9XgmrwyQeagNn4GsFjLVJ7BAVGeIViIZmXPMQUZwjH6muIbagaw/2AehKxhWF
tko4I3he8uUzFzYxagyVJ2YdCHyIVIkY2qIGiL2Ewzxe9WDjYSXY9MwVu9lGX0eiCPbDb5nbTIT5
eryplcfOPQr6gd5I8vp91GVxd/EtxIgcatY6ZK/k3Fd9TBRQV8zhMsh4u8CGbWtkoE/50aenHCO7
PtEbcBr3B6a1QkfGRx8DEGJRKeTAW1Uc4P3Wactb4rNu/4+6sBjsCA+rlzscAzzzD3R1iCeK2C4D
8l+yOT4wAqPHR2dPf7+lYn7ugdpzHlZIemhL6KLjMLYzZVGkV/9Kg5izg3U5VBP7o52mNLoEbSlk
6PZVDKvMMlgmAYqLjSraI0ySI0pDvbJNVrOm0TBOh79yvPwkR0rZhjDnnSM7yk1XADIwyETN6AKy
SsKkLF+xa5QovyUWDeLwjZclrpVOK/j+oU4xZ6uI1HWxEiTfU7CvaKxx2gH8waIQyF6BsilOGmGe
F772IEk0t/q8GmBw46LXWYKHre6IeMrE20pQVAr003uROHZ0xRNQb6aALoaEU3Ra3Vt9hm181QiJ
ncL801Nr1wJrezbhc2IAUtAkYvtrz8wEGKOd4paelmThO8m12/qJKxAvKYc4Isaox+zc8on88793
Tmw2rsj9SMroC6KQC2TCgjk9noLufEO4WYcdygd2hdb1Xs/U67iEHUsev573Mt77p7uncrsAHsOQ
OfQOSx9di6YCiaFnWjTx69MJwa6gqXuQdDNgjR1LEq2HTrL6YEtWRVIGEnFd7YgPhD+Sd3y66bYs
zPR6T9Ca4NcxteJsJFxLQJWimX6YFef+uPKu1g7zaHUh7ifyjSssbU0HSSCfPuMg5sVAhMifLBuY
8C2O7XnCHTzJGOM+8faxEESA5BHIj2uED+kZi/lvUyTdwNz1X4DKH6a1IZ/CW6OPQ+Vmd8OsZxED
KCbLE3f6oRLHRquV/LR0+aEZn4wMUeQFBjanCzi/wnamg1OzgoS/H3G2VlQKHfB9Qyy0u0FC8Xj8
VpwzDiAWxAUV8NX3dBMJ1ZtdyxzF32yQ7w5tQ/NDs/jWzDh8lzotdBvcnz7K3NmmLT8mAS+RqsmN
y026RacVmHacetooHc6wAhGKqO846FtZyTQ0NlVjLYoWYX6/8eC8B6LlmQXtUf1BZU3mSc7hpaN6
g9xVvvj+HJEecRNKAthyO/oyGwqYb5c5M6qKDpxj4/4y7Q5WraQybaQ6JmqokA6OflkjD4ZaBmAi
ZFC9Jgi9Pt6h7qDvqGYaoQ+LwBdJz2+hiMKmSM8SKLh9d3cS5MQgdjPW7CnuqgZGDM7UheEGl5He
V0U4sH2GXqigbImj9V9ogq3MqZn2gRqApSr5VCKUUQwNdLPSgbJPCZqcsDtEf+eN2lfEs5tw4Ymn
71nyFrG6j0wySq1MoA2qMxDEQftaeypJZouovkMM+5ZMeCcN4XhCArTIe6wPVpmZ6Q4zViZSuMzN
GW+UBelRtkGIAhBBxFvmQCsO6eAK1Z28Ul4EY1tE43XzqE0NyJfx7S+m5vGfQdKLoVxFTQhmEK5J
ExvNMLtjb9W0PZkI+fb56ALSIFZeV/6nK+HsOWHCz0V8/u5jtRjV6+/4WhQpwoZdQQouVaIEXl+n
vhtOpoU5BC+6A6bqLm6oM9nf9Egez7rZCwWyDp2mdLPfd2c/CPKKA2fbqHceI0IM+uh4koSI7Tk/
Cd22/aqGlCu3kWp30ZrCUp54kb1zNARPbeb+qv5XWqzIxkE1I2J6MvXm3Cz0/3gHUSTuHPyoDuR2
jGKCe24Q2qSBCUmhaD+jPWf0ByKgYCQyiZxSehoqhXxkUU2UVotg61bJ7GesU+Bvti9pFnslouRB
bpq1H8GKvifx0o0Ifkw8mQlJNNC83OqZaTLVrPEnSMe2LjEgy+FV3nk4lKq5pdAuFa8dWq0CgYdF
Qs4Zsnm57acKcYX2SCI0Y2bNZk3O8uX6+eTcdQCt7piwekaYLmcOagTAQIjdDQRjhda/UhNAyUOw
zqjV+Wpxcd+U53oQzfsQVqoWmS9p2L8AwFeuuKz2ad7L6V37WNRFkAtby+gQ5YNGbZqvhJIH+/4s
JeZkl78PyonC8Jhcu+VTR6FPdggQ0RXVqakrpqWYcXrOse7AERRK9kzz2lwkYJgnMezli20dWnIF
/hFQSnL0P615D7w1QT7ecrVx/mrGAi5f/hS/KIoFF9LgAZsyXQfAT/Vit8XLLgnKEkF9ooga8E67
UOtk/pOf2bzEcBt0Mp3llYB/wEYcVC9c/R3A5bbt1n3wc4Ah1UiALEtz9LD5LjxuhlxftP6x4Spy
f0HlcB5oVo4EzM9LvbbNy/9atCRdvQRkOPceH6uxHDmlld19qIn0p73h79tqGId6hvjEeXgmmp/a
uwRdp3OUGMyr5UOD9//N1OYLz4YoBpWuMsHTLAmT0behMHEls5Z1Kqy/lfOrrs+ianypNWa3dp5j
jdavpB7VnOhlUwgAxnVvRmnDgK89sAVuEG5xMtjDH1tWbzhbaSWFWipKy9+JeM3hsLS+6bOz9MEs
j/NrQcT/YIhh5HW1ukRcsFpH5piuskEvRodoKVybjHvBvabcopQBBKb4ClbZXPDf7x/at9qF/yjb
uRz0laYKWS0bJ6GDdA1H5dUPPXtpKhdBoW/O/Ctj7WXXqizWUNMd1MBaSbDNXo6Wm0YLoIzGqUvm
24NdaD/VvZnXCXH2onfCBeaHHMJ4drf9yaw7Owv1lEMOWpyFBE/f9iBjQsH4gvvPamcqG6XjHIcV
8k8UnJdK+/JJYeYO2+1362H0xlNji0OgRE1O4esVFiGdhF8SHQEHDrhfZNmT8PQGXwtcySDCL9qG
FidopIoy22q8uZ1OeRq9yUeF6VlKRGghjyA0fMEMJPVvR4R0PNtanaJ5OJ0hUWWFM+5S/SpkjX3x
6zxQDFj3/NoMnANOIXh5KZAXBdySGnjfXAjlbJ9Tdo3wpItzzR3mHFCyxPzhqTJpieKRYNd3/xU6
RmYhWNz7oDaP9d0t81RTgsu4ERKIIhuZMCot+yJK6UQXlw3p02qb9vZZaYZ2Z1ZHThr/cfpAz0ia
XR70xziAxSzYkVlcop9sOhPMm5jwOHlhWuL0rjpOKvJGiYsG/eXZehdKSB0n3zEu1N1Z5I18LCEf
N++jCJ0HVfI0D8cO4SYe++H4E5kV8AOd2nAz9j9zmYQgJN6E90+j2lh/zF43kQ55UZuCmcDoB+aS
eXu8kaozIgj0k0j9FxFjmf6JEx3Z3TvOWKECFhTuQSfoamjQUr8Sjz+5WRAs5mNvSsKpKf8GsjI4
EBdf/lcLalH488avvAcwVC0TmqemTnZuPWVX0nKltk9yydvbA77IElQS8/p+3f3NU+kr0blN2FoB
FGfk0EHWVrt3Ycpbo0V9gZXEirbgt2TwNbVln1ERHT5CvTwZFK6zXIPvPvshw8T3sXWb2u8CANg4
MAdaqcAWegBYlCyQZUXwxKi8X2lRadE/v0lZrbv5KQyDhT8oOZumB4cvGpftRk3d3Vc58ZYrfRVt
zw0iZQNG/m+U7aNqtllDAqAeRID/jWsvYxmFoVkXeVCdQ7yEsJnyrLVjAqoyStb9i38xioGjjyb9
Yl6yWKf2Yv80mUBgXSi7qRdokWYtUZy0tliD+GmAZENtOQLMap8LQE/Ax7bRWGqA87wCL5IjESxa
j04ilG/GQ/6wzEyuI0Fgymkh3ZXiRpP7oQfR90dZZpsOc79th67wmaSJPFZMPplrW/3gAIhk8tpB
HjKVyPGGDjMs9uj3jY51oGCx0S24yGwP0NWasnTxpRvbdgwVvTUPyGNkTPxEpuRESu3/ErXLjsSi
UOHyD5JJ1Ri1eVX1gFdt3M64SjdzWddPkQ64Xv/RBd3mgKEtwi3iGJZPl/9nt9CssbcoL9/ClMR3
d5qs8Fq5JRIiElqJ9FkPpqfBvfnYUFsvgVboTfyHsTirycm1GnidDYyt31yK4jGGtiznaXK5AKG3
ORQN1NKntP9U+A/c8h/hAmAA24IGC8vEB+zxkR7yQQTkLBddzWw85CGdVEXMlQ+bCLoDhcKwa/7S
rCyPEi04/BWBPoAIygCWwlGfwTT30/OHfWO+brCDdZhAbwOLFjnjbLEXIDMUwDd5iNRA3L7fSbPw
bv+0CJJtWkSGYs+lCRSFZQDTBJ6bstClNqT5rHJCIrqEaHFUfIhvYCRYRzNwDvOcrXYynhDE5Vze
lwlKNLp32YHGzj2R30zbe3d7bk9UJzp2QQGjmvYtdNFstHg0/niaJny1oxGhhHHJc9ztzoLGBSJJ
SErDYjJp1TJlOflcMkemGM5vCghc+x6dApmzDAwmea4uzl6RftkEoYIFJgPopg+LPZ2hMrOFzfpo
r/nl75k4FOWVZexWSnjHYVOmmyv+9o5fWpWlT29+ttrSRuHwtoojHkwmKTA/CsoEKWAzuJcENNj1
yy4UGGpV8bzsT5w4yFzm1NRXmWivblQT7SkApTNFwW4eLkI4f6agS2EM+vT25D/882B/cQFRTDvm
htJSLIxvQCR2Y/tigJACIdBuMd4FZ4GnlqL8Fb7HLvkVzvLAdgGrxhP9yctE4Dt0ZZFzBTwInH21
U0uRNqRzd+saS8MkCbXx6mReiaA6F0EWDwoytjkwU02vNq2Pb17lgXs8p896wzo0BdHBuPKDa62/
uNQ6cYlzedxOhNfxVbxrw0sjSEa3djlIXNBwun9KFLnW5wC+yau43HoJT46/wijNJZ8YH69yVfs4
2Jsehi0lC2j8QwqtGgkqN0G+U2rfP8ejdUeLVR08GOlZFUkhZnp2ZhRzs05AlatzSNuGXwcqpTAb
59kmBnCDn+nORU8hvjXB3QBmgtURtkRC0WnASYaDkno0J993vxqeQG/MG0AD6ibG0iwYU1ij4gW4
dT5yk3Og39EHRVgEp08orH/BZdj5n7K+EInw7ZWvTY5657UIBoGz3hDbjzhbog1is26UdNxNTroJ
+z1cFsYQseGIMfIH94RQe611OGX/g3Jsc2/KyHrQ7yEczZKyWKQGvdB1wrqxD1rjN9tXxBNwWOKy
diSKYPikt394m0A+vumfd48cwCeRl7I3OwYRcf+M3182eEH77mHGdl3JDfGV4GtKFS0IsVhoUs2K
j2LZhpW/p4McUp3qbcxKlQealqdWYE9hNYqCaApvz5sXtTAVIJqIo6XJI3O8KW0dqkC9YfPbFilC
aIHw0vqjO8hft/Maq9NJd9JuRK+ZQqGqE2H+leEmhHVftqRb1omG/z8a7NSGrjwQA9XU5zCdyE6v
gyBj6n5U4mxOvxEQsk5wiyUOTFNh7Q33HSWU4Hb2kYiGYowNnlrWqSGiD3KFOqaCjnx1LdFjqNCA
EwEey+RbcdlpzoPIaybSdfbwV6aTNF401kVLJ7niM8pEmVZPAtzpnEbxCHx92XbC94Lp8ZzzcLbs
zWYNl896lZCKizbXtABk+RrCbWi2ffMhiqoswIbGvlWtaC1xpKv4fAJrqu3+c6znCkpTOLz8P1Tx
1BpJw8/DvJRAxeVSXCtqYjJ2WyqV02ZYfd1vS1Te5n6TawHMPjm2bx95rgkJWP8ZUETxto7eNway
Q7BiOKr+Rgcji8ilObyXwNJ4m2eQrHRxbl/3TPWSXVTacrjQs3Wc3ATt2Fd+2oq3QY3d7Rh6bRS1
xm4ZI1i7d8fLU6SbPu4D3Ej+1AU9DtwqBv89IQ/J0uw8+UD/d0ouja+YkUlHrUtaJsHlxihokqVP
pB5SvnzTphnP+YRAEfp/uxjvgBKMcIWUt4E0zpFBHIe0Vbs9SDb618SsJy0Ym/YUlSWkq3WiVgHT
Jk/vd0mNPxcljQk+hoahxaJ6j5MoolRjqU5WIXGCcZ6Wwsj4dZEkOrZwt4pIZVLqq6rzJyXSlpg2
jdlzPVHjqtOG3qsFeHnqMYDGzM/iq7rCNktGF95OqM672IY2denfo+rD9blAabCsUympOSzxjrdy
c4p4VlbAmICF1EFjWVn3+xmJ8gZo7waimU9Ee2HNi50bpE1LChCPtLIFtLx/tJzu3RRjFLk7N6D2
L5kOqXRTAz3XICbY9FjUAm1msOcF+Sl2eh8E2rZRZFM0TirSKJKfq3X+QNJGXzKc7uLAQD4b0M9X
lzBCToZmygL+RkPbOAeitIF4wu5kj9Z+viUypi4vk6DuEms0B4WUBZ4ZTq4bmbbfhHiLyHnf9lEL
PuUVsXQh9kOf0hJaCb5OJlqo/ZA9QGoeaIpbLxezwLg+Fvju7L64GvGQNKhVMh2ivJGzwUh++Xm0
OKqwDCuxbnFcissNk0omOwk7e80k7rMBEgITwUrnZLaVqYpIU3RCQMrgExa1ETcyI97QtKDw0jmC
uA5OJxC3WnJreGG5D3MiX/hN6+TE8ZH6OVu6dnNMXRlWD54aNQJi6dQ0T6t2sY+kasQ3Jz5ch1OQ
4lN6j1bkOKiR4pryQlL++SEox5z9SWB3/fdyTjlDXLxjkACW9Uzyck1P//Mc5MKt+MA91lDoqSPk
ypVV2G1DW8Jh45zBXR/SPhPh8nKuBzeJn362xhf3/brJKELJsBG+NfArRi9dtEOq/E6LGXUsJVrn
196+E9OJ4Oiq9OXp0XXqpM7Kr+uY+tUaqZj3RlB/M9E9itkYv7nnEDUtzhoaxVLWHv6lQbsUGkbU
Gw4AfCImNeCHWC3SdY7KQoZtBw0h59fFE1j3sojfVKo99K8a5uGwj/6b2uQem1jF0JM0/npp8j1x
VNGwAsGhMSvA9Hhws0xuY23gRhbZ77mzF2/MHyRW4egTnL+KlkCc91vLroM2pzk+DZKKVmZgunMM
lcHTDMTZ8fEnQfTbxWNUAXFCtPZoJ8I5orr8wRt8itTmttZuTdf2+GXFf0/+FUOjICvT8A0pyBAw
In6J761daoAs76LZCNPXpOExedQ3nTQJbl6T5RwVjeh8js167rdsXVo+pqJgfiV+cPRZUporzi0F
fX8VrehZHOJL6wR8Xh/FqLcalRg56RuOcqy4ELXehaqybPEvn7FgepFu1nOE3p3Q14F40B0Eefza
pgXzOKu+OYCjAI6DYa0bLK9Wy6698gMQU4O0OU/4Bgtmo3wtrTt+U+A582v4DoGIRxAim54szagq
LtCPIfIIwxK/VuyzuenV9YLZQUFM51S1zjs7u1PcRHdX4NoAE0kYPnwrkwu1/VshZz2HLUOsvIAg
PeEkrfaWBYE1AhHFiz9Z0sm+eURT5O43x6Jcghv+uP5iOpCdLr5l7652cyhlDFgDRzPDUcFIywmL
0iaybBctQgmdtsMa75xuKIZoBSBDhupGCW96LloTAEjOTmC3jEBoFOKXz0q73pxDnsNrP8CPGi/W
M04EB57vtcnwqd6PZRQ8epVCbCinef1mdXwvlHHU7cvPYdViyKpSV0l3FIud78GLU51yrzuaMBd3
fXEtQ1zkMo4m52GaeZodU7oVMyPDpS61lAVu1+O7qgHDuTPNgzGN3flCvldDjJ1cWZdJ6QC2D8VX
jhY8WwsINQdpZbMKUK22FrZ8qWZ55NueucJeh9uNLiRzhRzmcSgfoVZTWV1zD7fQNMNLQbr5s+Iq
kdTwgN1f/Q43NXzqh9UrQJaO21gVef4P5IadODvky8Ixm6I0zN7XtyC2G65BJTU5WjNE5IW2ff7k
P0Hf0917QvzSOb/YjhIpJUwbLWbjEZ6TkLDAWvmVpi50DSXFjMK2vm6JKBiXanEUS9u4ye62xraR
Lpj1+cngWW1L1tBgBX6y7zVtyIot+GXziqN5w7rN2a4ErSEPdJ5SzAdbHzvpeFslTtdqfev2MtWL
ql/1Pe99nDTOnJnH7KTkHCJw4jM9jbOkKdSgOm9CwICmhokjWXTC23MAelAMvzbFTZqeVIXfByNR
Z/0O7QbWOcFNCa7KCGxNDvHzfwQyRclodDutIS0soTD/FFq5QEv9nAfKAbAbygt0a2bZv/QndWwC
tpl3Ge+INh6iGONtC+gvojxDVa0eUGbLn5Zs+CrwmcKmS60uMQbRDl3uBAoAQqwWKbzcS0RaIGoc
uH7oLFqIk9eamv56x5/A465LaXJbZzs7NRpg7F3ckTySLQUVJ9CWQezY7KkEBX3uwKgOZ6E1TaG9
0rNG2doWPkKVtToM4/PgfRErta1vvBsXQixUkWTwMfB7RJ2JMa0qEOtZG6KTFPiYEYygEE4928+G
43u4e8iwbSh6BLsiGSGC7X3uUDI8dGlTd3I/EUlxqT3trrxrw7PY1LImgt4w5bJ++QT4gvBxulC6
9fpEiCak2WXnULJ8XFo9X4FJ7TMAobd1pkp2248+f//hrOitBL25oVBXaOiFQhAIwr3WZqVqQi6C
LAxthQCOGm1w2trVhnF+wM0XADZMYLFY1hT76Q1c7S0PBgqej0+lMTMtsryFHsckceGu6Afgz8Xv
tNanW7bAi9Ig8Wy6cHS3wnI47ilCbIwSm63DmdaS6mEZb32jFPf2ZKjJgqcP0IVJ2TwworN3ADgs
+1MB4I2HgMi1PoT57sNb8W8GV1SOVpbI/sMn7knpiqTpnvD6DW4nbGIGi4J1P0sINihnD10fOHPp
Q8c5uZUyw/CEdb7VAAZmsmUPRaUtpE2SGsPektmUG7nht7ciKvDk+eWrxfjmidYeRhLN0CrZVQLR
B+9OTPZHa0+ibjhKKu3DEU1+rRO0A3QYj2ouqd5jE3MpvucN1PAzyF+yMLk3z5Ir+myagx3NobpJ
BjbuupOyzQ/5i8P0tU8N/FJfasZ8Sb0UhJm1+jfcCtRddj6FFAiN5hthMzLZalxox0JccgsPTLpG
BnW5YoQY/vSo1R3N+WJmKjvo6jYjvfL4a15zhmc0D/mdle7NZAu1DOTj3ZarGyRbhpOCsDl+Uq5G
l4ldzKZjt8wu7tx5Rv7YaxUMLSHBDgMisLOpzxGgNNH8Gf08CF2k/cVgMuSodCogS7PJiy7I4GFi
oM96qGltFZbhR1JaUdQUKwqCPzQsIrmjRKozaLFlOAVyH9Wi1Je3uZZIi8L1ufKj86AAO3TCTCf3
RzY4YUUQCx1qDXKPvYwbAv7FT25uppM2lVFkvKvRewxoXepNfCt0dDfnI/Kori6od8qGfW4xV613
6eQr42WLZWDXHQd9nCr4QV3qsVPibYiJ4zXt3CdmLdj24FlPBUHEOJh+NhnyMDZhjZsTY7+x6OdN
ml/ppYP2tlXU+VBuPW/6Ak4yBsSkZy4QCg1XNu67wM1S5hA1bxJD1JkjuwFk5jbBSdCAFyDT7t4o
hGy993DRD2iynY1xmMBgQN7Qit2Q7nNK0XKTg0ezN+zmw7owGQwGLOwMmz5I2L54yb1UqZXWuVDD
5HV6uzFToD0uU3PFFNJkiNpVtj/yvc/7wH4a1hZLs9Xo6Jz9sU6ldl7E7VOsYZSQ1mbPaDISLNhs
uYiaQ+fq5v5Oq4ospvMdTINejJT2p3zPxKQhI9LdVfG10o9wGutJFpkCuaNRQx6xJNZHHB0r7zQM
rQF4ZKkypBBnrd3GJUS8Y7x2ndJJDhP2vc2EHVXt47+xEawd1bwv+eByxWk/yB8hur6U1cvVwAkT
4YR2K04Jia0yFelGgIjTnnmxSNYiLR3kZpJqqaPkpxW+B9+oxJpgYXyZIe3MwO4xi+UW9c3TyWho
fkP86/0HG/IhJWHJEgLPXnq9eZW/j9C5Htez4b0XDIsk2TRQWRLUVnC+0pLPZLAa+g7IwhzyDuIm
5GWqtrJGCtJUTZ4oVF4RRPRbpwip11oCEm/pmA2acbAibhCoBaxVPqL2HYUauhEMXYfYdqxtROv1
+hA+d8E9sjyGfTMGBbJhlkafYFbwH/SkmTRdmCTS5PwqdMKAyylM4bqm3GgtECo5g1P2f2RQKrbR
lIgJxi6dHeHRH7imae2N7c54xd5ot7LzmZDI4dbcrcKb88WGwRjgIuOn1/Gf8oTyFFL/etKhIPIH
bB5YwGQcgVHLCYz7RRfcRSPQUw3KVihxhaFDO4/nBS0MtdLL3XI/biIOxcW8qa+qLEQc8mTcqiTC
irlvDr3sKNpohCHfhlhCbcEbqF3WisKcur3wSWJgzeLl0HESDjgpoahm3KMG1FHGQPCxPobhS0YT
x4Kvu5BbmErsvfZAyKJrpXlL6cCkKnVsx6j4FRbuMMDxkqaeMEjdTN2vBOnL+tyMMkO6B31/3oqh
jNLezH9erfaiOBqOamSmhW+GFDNl4uvCHX+j90XmQx3liq9hx9z/NuqZz2UBI7GRIYCkJy+x1MA8
ifFrJOpFfXKm4neQBOs68M79Dl90bpAeXaBhrpL6uWf4D4Fk5xxO+brYTLQq3YA4HpPnPMecwz/H
+JpJzi1T29p/Un+PZ9XHlWAnFoIzQL1psE4lJzoVTO+YngssHuDNt3tys4fB1KeB9ysZoa+6Pye+
rgKz5wHcIOpJB77UjnGSGrd5O0zHxD7vOXp+JAjnQ3vNyAf3BbYyUcOjAU62O4tG2fXiXrWVaplg
JeTNpwgT9RLAfxaZLSFHOWcK7tOSxWv0Kayj297PPc+VVQmTs1nlKdFU1EKW3vTIzj/2Wq063MaP
1lDaySSb2rY2pSD3J9HujVvqkahAz1+Fx8M72DG6QKMLgABlT/DdrcE/+4OhCzHjIPNqJhG1fCQf
bjkGdGP2Yuuu/zZjWqwtENWmZQ6J15qCKlyf930/MiG8WH9VhlcemqF4Tt8ZXVbwMgLr0iZwE2EU
UvPAYajRWO7hZN2fuDvwZpLs8/P7k0zeXyadWgvvTfRn61jaLOFZn2rF7ZiykPKnW83TNe7SeBWd
76olEQ9S0QgGlJ9vxDCIESBsuQDLvK+HUp7ckvJCdIq2//t7gnDjQwhvH5A1u0t5Y1u+cj/td4Sp
Ea9Lol76i2dSxbSo7KXaVf7NmvDigzbLXdfegxMvNukJxsddKJHc0wQKA0j/PwKItGJYocN0MHH4
XjGvT2KHNIaOK+68yxy6bjSMnAfUYeZi2lLNFCpR7g/e4505WYbiYYUPudHFnroUVF4PpPO1ilnP
GyBvdzDtfsFRj0FpPLONC5bunrXDSoZXG3cgxvzoF5ijRrXM5pD6Hnk0Lp+lIhKuKneL8XXfCIrT
OpvcsXw+taLzGnS0fm/9FMHsHLRig7Z0uTWVfsMjTcF7+eZ8G6pe7S3mIkdVs7OCg1YPYZg+x6WC
jxvOIUidEI4U333ICRXioX0cVU94hegR+sOXK+v9uy0dQoaZ7s7fWL5X2gowXIQO++HObI07YuHJ
/mkWKbpZAyKK4UXug7hvHooL0UVMp/mOczG5gAllGFgCm5IHAk3tmOSqa/fUqfw16IN2XgckofFK
oNhJ3hYkf//NgphiRD1DePUXapX3SeE386gHjwOi+sv6taQFsSdB7rlAYV6z6W16rH0srGipnk+B
YNeQKb1XyC2p1OnwxLoS3G9qQUYsvoihBnWk5sBqnba2PWKkknLsJB44wKtWN+cfhN0Y5cOJnX1l
GRlhz+g8LO5+pgLrqP7ApegI1uQ778GVMusqPG4cdkAe8douYxzO42SYAZy/n/2PBgwG9HZUZFWD
l+CWhaOMAQ+JXw2OEWTe0gCF1WRoQCtUsTWS/oE6swi4KJScYZfuLVdlepIlKggCTxtsgY/vCdWi
/EQPZJsWR4jA4SEkku1grNECqt0LLr9GSb6t65bZvrBuEEQU8YyoKWye4zr4vtFS7pxGfIeIeBon
+zGLSnfRXrMtWLb7ttqI0N9IvlETEHAATT3N7mAvY73vtoF/Wn4wKzcQhw/X3WnFtYFraTv4o1D4
GaAWFGyLW2fx1jHL5WDTxHSKYyGIiCQS2KjHyRLduaAuZVzzEbe7SLNIQznE6XCvyTnVw6xA8Nex
W2Sn7zPjISzROH6BN9OjBvaF9OLa4l9RmioOtj21EGE9OuF6azzvgWbBctraZMzBBtBNuqn7Jenr
8OVfrB3IwXsd8z33XSjsIVNm8y3RKWSI2ni0SyAWFiTuTeCyyNqLZnnu9BTbLtTqP7KEKXB8al4O
l2HZD8nvtmFHbpc47vOvi88iQu2qFi6mE7it3HD+B/AzXgQD+BBYSB7c/gvp2pmbAvN9448+styL
qlyCIjFaMXEIWeUQepglOZHTTYJIq7jTTsNmWQe+t+tfvHks2r8ZVEkG+Q6NLxJsMMyrlwqc+dZ5
koq/f3POnYcb6xO3NU9x1hevU5zfZi4LzF4FYBrwg7PkIa9NOWkE8hhQhu5Kix0gI3zp95c5BM1o
7YWqCezey1/yVrR1D41IhxKhTUPf+Nyos+Z8YlVILIVmKkbnryBqVzwIpfq7TrqjCYveBSdysuiH
0iEObH28D3zZcT15cTEC/AUkYGRAjdWSe3IL7p+ekntMQ1zhCndCeAOXKxSGxDrBnED/LOpaNrj5
Ug42hstUrZpH44IEwPeciGF+hT+KuASvPpv/q3MaNwS4Xj4PilPZuETr16SQUmi0J10w4uWyLqcs
nB/30RDA3HpFhBRhLmzq6gnnA5/blL77GIbVNrFfBCiGodHL7egoUDbxgDz0PSkEb3MkHL2sBiNY
+lQPuyiSy0yR8W5VCbio7h1ynDbepM2L6sInZQMcE/ge+PdptMFzBT8QCwDkgbpQn9CldU1ZoVr5
YPyaYl2tpy+sTJGVSMy4YN5DUo0OFQK9Q9gDOXxVfUbolfRdSXNH+9a8UhhVfBM58dWteMZUL5ei
NUuciW6hy/Zji6fnVobfl2LNRLudt7+MiIpH98N6/jCiSMvDshBm4fQV38JS2Bafe1wF07VkwDxN
9FAEEc7s7r92QUKXB+LYzQfhyuyFGs8tJRq5exOW6/pfTjQzkVBEVYBXSxBwpbFmTzidfwOVSSo7
6yNomXhJsPKrncmQ3yq7aF6W6J+ntHOTJQWQJf9inuDXsbH61qHkopnYvAGcyBfVhfE23Udl3TxG
vNH8gn/9bLyUBP+Py0ePeE0oKg+8AiVEqB/vT3JmxX32Orf/ray9qzl0ijggi4kooMTMqu9tOLgD
yXi81lgQ8YyzJekGChrck3eAAMcwz1owH4lncZr8ysxxMo90Dl9SN+Pqk0BHt7EyD1/mnuCxARx6
FvZFVSBpW1skM62YgmHDwMLcutJlVXXcguSSesWtsmZeMudFxCJlD50AN05eGPInBEDo4muXKQp/
H5G4DC5BlbZVHtSIIxSdIDe/C+m9yW4yqf+3y/Q+28LxXIIlLx/i32tx04ej00rLYAced2fEGVPM
CuuMwTlg0YR6AMESAoi7Lmf2KwruKfTnGNN0+/AKgBoEzyeXzOX5fX+RIFWOFI0EtcDIL9IX2r9X
QUrQlnplF6raH+2m9WDmv0fBKSOs6d3Y7/nFRiRJlREKq8r5OlzfXcRo8aTjbaD/BHmDHE4BH1sT
9dFE2LkbQpSePuMww36oOo6iwQUFM3andaQ+VLq7qu0Ohu8RCzU5tbEGcjYCjw58Y1scbleJOdiX
r+uU9rMKi8Xq4MuhXpEhZMRL0XlWCvLh+33vcaCZubqI1iJTxOW4nuEuPijGGeMwOp7Tryc3ymY8
//5MK/WAn9YSyKdU4uvWLqKi8iTpHst9w9u8Fm7QGc7uhiTRHISzScd4lPVfCBMeN4EklejkFp6h
/tgNRA0/rmQqJTXVA3i+lqzaRyOvbV9Zx9K2RgkxxnFOD+erafaT85F5aw50h5GMFQ4tth6T33DU
yhq6kdaMzuxE+51rtmOCClye8mBPGnbv9PfRkuOwb5CJcevIEgDUc4JSogiahyZy+eKGRzVBfc00
a4QKZePBTtmjWEx8M6DBaoDuPk4CAgxDZm6OUNId8pLLTTuo8oc74+fHZ+Nz4bzjRBNco/Ji0Iuc
x6r41p0KuZovP8JOY7nVvAoBEnocopi+AZh2K8wKGN8keCgdEVbvd/80nwu39wmI5UWTWb1M8QtV
mBSHWjvpx+QpfQRXegHdYrHkzrDx9+GsUkFn9NtGmoN9whfBMJ0g/H7fCsxh27pOyTgbs8oH5zF8
WeTugfesMlYRVXCejYxCp46wNnm49BcWhMpYfK0JHwTnvxXaopFJJJTzU44YipJzTBsqnH06TAjo
1VGX3fZnIyqnQ7gCq6fro1fnoC4hLDIEg+56LbdZuEDOSKT3RCnF5MKIQEPgC19asnIHOZ6OTGU7
p+z+qYQ8xQs0NFYVN/m62cQMG3R2G6BRzRtCs91gbOlG8evZI295shpDK+TA0ejHTDi0FEDbdET9
umM/khJbetJL35pqFTicRNCy8nwepV+IfKOJhPF1/ZtW3HMp2SxYCH8oxetp+IptLXyxUrn3nJ4R
8IyVhJvgUh05njK2gcdePb7uL7vg1rJ2o9c4sh+2ycO6ymZs1i4hah5fGIKhUpyJkWls9/o350w0
frA3mXrcJgJbj6oyQ9mymhHRxOVjPgS7c/sn9DZcbuxpWZhqUsY2kIohYFn9NM+GW874hVS1MU/3
RTOVYP9wUtJLwdpqjTvVgfjDLtk9XBYiIOZCMNyodIX184mapJ0lrv1eC4kb8hcBkPK+JcII9tU5
zG2oza8Byex3fxNYWxeoxnRevSfXHu2rG/pqG/Me8UUCYKP9w92RjU+/wv0fsTDUHSTJAtLKJlIT
F1CVAhUlU++YOiR0OZX8S+Drx61+CwpWXa+oX8VgpCX4QvLTlWjso7EmJ7kV87UoK3ida1CCsLSh
RnKBmG/KSUCrjSj0XyrU/BHYSHhNRc7BmKjLVvUM95TDJoKqORSJiMAXpGyFazpiJWDdtaJdnRd0
MEZvkr7bvZGBwlQ/kjpLMltjOoG9JRzf7rntYiJDBO9UgpE7CMBcCFcqMS5+cd0bD4v2oNxMWu98
A9zT8TgwoP6JAEgdykuCGSKBLjxpRD1bS8Ib3IGrYPUj0+DljvVy1kcD43rmEnyrF5ycm3KSSuUe
rwJcFsFmTa4cmGm3Y3kuKAbD6/1IRDcXzh9DIPaVBBGRoDoXRcTTqRY7Gulm8rsEAtBFYUeGagYa
7MSzDUFu1XE0uVob5d4NbMH8V9f1S8ZtGDUJV5eKQ9LjKgyKl1d0KeRPWsKI4VBKmHY/PrSDvz4G
83jarpb8JxABqqE215RyKt9yjwmZsytNzCcipcZapsu0E3mpHdtnh+1PS+qWXv7AAJIMbBeQkolj
ENgmyyeRL/H1QmfqU8Ju4deLgtotp+axnIqe4hadvZiYE8VRn/B/Ij6Flu4bNoN5WCRJzTNvGpDF
qdRSa7hhq6MdGZKOS5M/7Q8GDn9BfEFTksJhiCSct8cBPG9xSlB79sqkXe0K5s8sxwTqYvvhyPFm
R7ktA+YnjnfgZV29TV/Dh6njVFKdC642odSLPlZcM8XMwDCKogqW7JJJJyQ30Fwigo0YlN/JIkwV
3BXr1hLdAxfmCaW/qeeTKmSJA2R72Hcixba6zJI5p8JIPZTn/ycxTegD4egTj0BgqI+R6bRtbcuk
q5W9lknZSiFfrzuJKrD5IpLtQS99dCOxD+gjWqfBt5oKGFPIxclWkzjyh+97r5nI8P/i6JRe49gE
hOyvFTVyYsX8GyHCNLFRyTyUc6Ol31lr37+alvr6mXnCADwOyN1GiQVYWTWqRNv0M5ln6BMnCW0J
DoW27lZ5r+k/yajJWxr/Tie0js8Wfqx8iqypg7y97KN7c8P051NF08u1Pr/yeqroChOqZpIDEuJb
ppLiasdewntwnpvwHHbllvPWilJXnyN2cbq7+rq4a1ybDVUYdV13RGCWh3ynLbTuy3Xzezs9vU2N
ElV4cS3oKWchaHK/y3+uh/8lm3wLfzhSgTfpvZftH/PaD6E2oaJpuVHVu95gGPk6pMwiNNm3xYJp
RRdeUc9gSiDmQc8KSD2yLi9gPF1N9Q+bAikCmzMmT/rtYGTFcTz8ckZudEvJrTQoewISB7ZwryKL
VubiKxWWF5MFVxvnaCP6acSayXBxfHhCFkd6yCKqyIWAD7O7MYSGNv9KPV5caciA+WiGqhGP1Nqt
eBWZeXKxlgVfxVxorI5fA/gM8wuS9hIjQSU/KLTmbEIoeIJF3nR1IlEAXnkNTLSVpHEp98MjgxOE
v8E+n7e3c+q+4ROc/2g6Rmq7C2p5q8UJUE4SU/v81j735YqdHOmEH8DU5grQq1YUSeP0O6y7XA62
1qalL2a2ZvoZOhOsfOE1xxAyd5om26Oak7zbMk8y9XN+b9amMerLiuA42KMtIDkDgDgL7voEFpW6
Fk/xeMF+5BYH6XfvxSnESCEZJ5p9r5JUB6KdTZ+JeUxPsaAI+vnZVapJ97JH4HE3V+ydmLeGNn8x
J++dK1Rj+0t5AVL7yuHDsB47DnyMCyHsOGbhs7LXYxz1coTur10q/MuhpDLP2q2Zu89EJpojypKH
mDL74wyx/VAeUkDWSrixKBUqyBpsr6GoL7+LSbjUOJ5oCwE/ER4thqhzIdaa4Er/K0mfJTnvpmmK
T3BP4gkq1OwRCbhWjd8g0NKYesYoWLpBc6ruzkdxhf+vyfI1mY2l0twJP6Z7syshvi2V+O7HOt+5
pn1iG3ivzxGhmAcUGmUgyzwbave6XGlOCEKgCZ0vxx/JHyAZlqE6CekezQwuw2T7Y5JsiYyQXFOi
2P2La6/UvegICoo2RicOlhZAfAJTeqrtTaOHolERRaM6L0Os3u8EkZ6KBHHH1QOnPib03ljuMqRe
lS9j9e7GLiriDoBKcDfl914eiY1l1baaW4nfSnf+n9aTUj/y9Wz+Pm+CZsiIfMJhJe/uyQSdtvrn
5lADY65T6xeAeORrSIoYWMbeDcerDayPpiiO6kdih35ui2YPV/cxFuGi/7JEPy/03Bdz1UaITgqH
bxucXgMXqn1XSNqoSodQ2yrVtAaoieAesKXiT9326xOgUBhql3PSMvRx5zYOW4uw73xhT3CxCymX
UGO156WUoDyC60cjE9RlbSjrCVIOfSlXKmO2iqH8pElHgKkOjbwS1yrEfFs+LWRPsqnS60ewAok+
GNxAfkgCjbSxKi40uJgK1c14JH8z5BN3u6XCM3WJ316FWNgJQyaFrzmcBfrn1v2TcQ4e3zkDGveR
bRnrahXdV6+98ednVbUNTho+/opVXJiOZAr0FS/e44Lpg+2oLzYq1nPPS+V1QlDNamY9eK2VQe1M
XwR5KDMg+V0YfsMArGk/93GGnTC11EOgXM01juA4Oa/F4fyBJv7ZpsO6gyv5MAuP6owFH+h1T9q4
ywzMhZ9N1ICA2/xR8aXpJrkt1GpwZAsZ1dJxwTehC0Nz+BOO0YWrtJ3ahrBJ1cIqLvUDYD3uNaFJ
O2uJJOF8d1umPQlqkHoxEFqY9mJ83S+qrCQ5pV6tHJJmi3jqPBytu/htKKEcaXOJqclfErPiN+v8
XyAJiGuSB3ZA3r+s/D+8HKTzS/NmlQwYiZaCyhxz+FsFQsYrxpNLg8YZo+kb9lFDcaalbPAAQlBH
hyCFgRDTwW8udbeWgSrcigj8lZpHtUvuDf+6D/PsoaXEzLC1AvHPOY4ARynZvl4yRoHZN6JnqRDc
WfcaXjwFq6qopUdCdeVLZYYGm0tRksw1oGBD4qDLlIQSZa5IFuCS/XfD8FmGg12dA3AICVD0Hqnu
X1Sv3B8uvwRO2QTny7/6aZLL+TzdzG1+a8DeTTKUQMZGlsFdJ9bUoguoUcNq7jB5Z5SXRekV5dcZ
x5RSyIuVlkP2myE9W6z6S408v5d60i9GAtbGP8KwPoK4B1A3APv7j+C5b50KQGm3vMv331FQmHAk
Eu6V8CpzZPUsCbG0r8sQEV/oAA7Ar5lhuwJcx/b5M31LDN6VOdrdFXf2V5iVzZPszIY/BggovNCk
N18LmTUh8ggDBhFOliAaVs6ysgRO4ssyVb06U6sElkAXDLsJRx2IKIDZc37nSD5qkBgPWBLP+c+p
t2tLGbOjr7WDu9l0svFEwsD67J2DtFVTfs/lE6I3A+Dv11lt66Gwxra8YkpkIiKwx4MI3yAx+6Q0
O+M1DbG8f+lIKXcXF7g45iJgwOMXJLD826haYi7RkJkX+jGFgheKz0lhhiviDKZkZ7G9UKtDZY/9
rR8b1jv5fEuZkKWXKWuSgQjzAau7CBPTDZrygr8o13gFq23ar0b+uZyw4QHFlLGryvee9HSPC/p2
zZ+ANS9rDS2xrII6ujht5htFrb7a9I8t/3rEWjxwOfnAtK7KiFuDpvNAMrH0sgx3XlRrKMZM7f1S
o0W+dRtulQWE7w8QUYrkbj/nYHO5GK+4cz2Qlh7Z4uCLVJq83HtNKx/gu0w65Fztd0EOcxMrp+4h
Xq5gC9c7rITSSA2z/rDiGSrXoAnJxy36GG363ASxXQVzXYGCKETRGlx/GVDm4IuqJcc+N3dPxjKi
QWvcbP45DSggPmTO620ut9iMFGenQoXIWTjda1gAalF/3/LymOVedGNRXYFWOBWWsMLAkflHNJOW
5wJibLaOvZBwA66sGRk2zJBoVq20XZ12CeZBWrFXBZdYqPvL+FAg1FG8F7yRoCHXKfiTz3nzlvQM
s5zjzHG3yuTPtMCpH4jJxQ7Du4268OSvQ8Frt4HjEQ7XiR9MWqmgnkLx9CpI4MtvhiCtFP/wfgKj
R68z4ekDjj+VezWQ5bjDdm4eBziOhzW+n/ykDQX/FgcvAh70R80EY/Sym49XU4qIQiuy41nppY/E
6yWmjGxoss3XJf2knOscDfqMcNT6MByrcHaSCdxi00s118v1UImTdXYGnw0P7l1omaRlf5N3EI2L
pV5MTgX+FDxv/AAGK+O+JoclwmwovPePTYE1FeTtJlVYtmRiSQs5BmM2CPniXqMeys75AA9Ekzqt
6p/PyV/4KZHGLqBP0mMSnwstm6GRDfWVTFnf9y3xiF5UuKfd9hdyKuQ9GuD8Nc1Jd9jAeERUoruO
UpwgK4jKxo8I2vF1Xq/u/8HOsvlNkfrK0fC5yNYaghddr5prEB0leEshdZgcoEiaLMuDauLfyQwk
6UupUXJy5QanefaKBv+V+dU1taWGU6er+DohrItLIK7bnfxCQdVYdY6Q2c3RqqVTB5Qp6YEfrVO2
6CZZA/6uMlU6isEQBz/m0dEXfgpnSm2aGMzEEqC8CYFOMeR4C9iQsVQDzPfkoCyHd02orKhAuwR1
ySJYF7siEzfMDWQNQX0fXVzGO1KT8bEn1/ciZv5IKQF+cRwCRFjUyABOUVEL9N24nvWSjj5k9C9o
JF/vhR0yOhYQQOSvDavbOMzQ5NhtALwFyF0uWmErf35825slkagKpmav6RvM4riimn0zBaz1+CNa
KzUmQ9EcvxBqWyJ0nfaj01ZiDYALbFcL2bvRnbjUXQu6shKDphjSaqz8Qel+njd3kmMcGQZwn8oe
f7HzuIs4mIWNN+tu852woHhcS+QD4v9NAeppG631HTyIxUxcaGkykswBDXGo47ml4AQuIDw7Bk+X
NnRsnOL8AOaiEsjTeGPVifq2vKb0nni8DmhrlMzFJbIgn8Ylku8OdJ81B9L+GvVBnp0Mf3cNw0WH
iYUrRMA028d+oNkVEfv/LcPxBLPOsnJ329+B++lNZv7xbuFqzCTgb6k3MGNoifzqG+3qBXyMO+Tq
572m1T4/eVz375FllU7XC6+Lw9mRlR2DZzFMswDfPcKhq4EoFaY6oBhDhQa7Q+UW6986GndJQ42X
bxPaVLPrzdTHcIXFiNYQeg+fgT8HpndN7WTr0Id+PBOyguDErjkLo/3mUEAG0BBw9QzwOh3Vts7B
S5BuRI4uiRVbAnVQzGIuZ3Tv0wlkJUXQVxJidTtoY5NQdNpHxRCfYJ+56ovtMGPK0NCXWO6YzF9b
6gHxyjukfhAPQQ3YE4ccRyYg3Tn2xSRl0rp5szh8WxJ9f41h+e+ZDiBkjJ/c3DY7Kqbc8yVhczzl
v1nu1+Yv2ioGux1TltOsKM/dxPSn17Bgwuu6hptuU3DrhnNwGuD+5mXZKm0RFNICtQdBQNjH8yln
6atnKnGITIQSp2jdcyFR0jpv9BpRJZH5ctAzCVMwPrfvTJ38kZq/g/UgkjBWeKSgYx1fFT77lfzO
zgkuorkdtcqW4O3tkWGMSgaIdXG0pQRvUn5L+BoQH8kMrsRF4dCrLdFJdwqVFHnm6d0ISsCo+pfP
3bwVUWiENXitIohcSVaTnRBvn9V6pLSOx7u5rs9MPss9rRJ/6zgvSK9oOL9Q0TkM5h56GqRW/mfB
wOzpum/9Dt3GcfFVHoYeyVuurRrVWEVNAi/qgDD0iAq5PGlq/fkbYcz5kB0xikB8iW5426TS/ZEj
dXxkr/5K33k0NHqg3+3yKcFBe+Ooi3HOQvtXCUHCk8CK+8aqeVjJHrLcQN+rlxrGZnimEo4opqFD
oXFLdcqVQ4BPTD++zih293Z9OA/e0RYjy4y+KWJjQc2rdhltC+NAugO3t3KcSDF2Px84HEHhNbUZ
XS7k1P9+5gFouu2I7h1qTVtAbSeNNZyA8oCZkb0YktKrgzOU8MZuoStJrY4ZjcfxoS8FFyi8H3KO
OQxiS3L67e+3N5R/4XtmkphrEqHv2TM+i2RbsAJrHsJX5qhZ870stEztVKbMxDNnyc448KX/rv3Y
F5JDFYRS82x+mQXO0UDWm0oFe+jmwnEWGP7u6Z6mW+ALcPhkA64nwEfWg4JRbEIvqgyzGD+3SmBm
mOMQz44mf+SelpFGHn87+m5Dd+4n7L+/qlq7OJ7j6VCI0h2A8IAPGXNbuXlrj75/Y8c8F+fhe8sn
UzQSBqavcd8effC3qIH1rJrV2vq9pMpGBdveSvqaUiKahfaXu21HXieZ4qs22Q7vzvk3gAccvjX2
6VJQAAyf7gcHyrk6FFWP6Z1/rcmIXmdgjEN4EEdvrSGLmWkcpsKYFpkBaha85ZGyD/ZpKJUdYI5d
+EJYvIWfYSOIef9OVgUmwPZ4Qq8CzsuzBLM/Fo/Fc7PvztfjH79IZQMPH6TtPQ2OeaADsMgk58Pb
ygWPAqBQB5KNWulcLVu20QJtejoOqYZ0TDKJEYYdQG3wATFc6xReJk1ahVuQK9ZFvHAyJCZAiAnF
2wHJD7jI8Bb5Pv6zLPA9dXwM9uSX2dUOIVuj6IYT/p7MU4s6EaI/w0+tuM73ESTZAcR67gEU4fDS
QOTop2+CIVW5zDgCmcQeDJuW8R+iflbXaYaxijZCUWzh51axJikJWr1E3lFN9dB5cdK7p79TcBLj
KunOcnDMTnTQfAdWdfXZg68/Epxm5O+/0g0uJrZ/DLNjp02Tv3QTxf2010twmLUb8n7YCDSSqr+Z
gZEkWeu9g80yBHhIcMgcJsvgVvwInUCYTBzJRufyxyy4gR7BoLWMOrpyq/UcqBXBWk6TwSh0BhOE
FQQRwXe8dMWuJjtbkOW8wuzgr3LyHU3A25TRq7kxnW5tVV6krWv+nYAyWnKXj6D05zqVhAbMZRBC
z0zqeObFhcUKaq/7nktnLJ8vaz0IR1cF402eTByPpXZmkxx7bE/bVoBmbM1FamFZcMK2k7unLRGh
ayFCmSXzSHS6qvGeSDT7s9JseeqTg2IVnLGZ6r6n7Xp7eKwgt1lyaquC3T0/XiR4O7MD7SOFzFfG
J6q6pmBv0hsjNXfnTPE+tIEnXoQoIZM2IfQxsnwQAGZb/9lUDZNwfX221GtiFJ7NIK4oTZhnwHka
RtUdgO/oe7KZHmENn8NExJ9Z8W+bHW/i1oZYSFFs6RoMaxC07GajbJY2fCqZXmbR6MAOObQrARfb
irT1T0QBg6XBSixLq+OspHmEXKEjUVczRwd50KYdZB3w2qVVRz2ivWFaUMG0UndxQ9ZddIvrnWqN
yZRwxxMsmdO/7gLNCQUbKKzd5PO8WSbfs2EX3SABOJkrvPQN1Den2Iostrb9+u5Io3O3TARIpHkr
CuYwVRvAy3UrsdNlfZUSxoUdcObd+Elzf+dH9OUIsR6mew2Z8Np3TPHarcOGF4Q2BraKYQl8TxWM
LWK2PFK2IC3AsFbBn8kYMqg6VlWmK6cJ8H1iUGLyvEL/usGkRPAhg7ovZ9Y+MDbEhH3SyX3H0kXP
ECeRiuIK1jhpgGqrqmPTPg0YwZKCxiexLPsIyrmsBmOJAMYLeu5khs5Zfujo4nSkznew0kb8v9I5
afb14YrjP2tD7BKLvPxLLA1x5Qu6fOW4+hDvbtyquG/2VIeXoqt6Mu2+hn78OYY1hcbu9QdNJsV+
70LF/VposunxOBuE2Mv1/sApDvLHrYo7qnuXfj2h3JWa/txoeY8plIyj1gAaL694XuSLp/NKeJ8b
dwOOacYK1nEEeqZ4UfVGSf5RTrQzpUneMGDlYTOM8H1GX0ZNHGfGGIxZIkXKRWpWa6KE00UZbGaM
5BLbAQYYt47+jYeWFljzCE5JrI18OyHVTNGbobyTFWYSDnnU6rFHawwkvYV8dMmApEpk3j6zVhZU
zfycKJsk8wJKYNifk4xpzzS3aO7faer3HI36xEKlXqdc2Lq4oX5hyuHcOQedGwNHjdSk/H4V6+VQ
lJGnw3iAmyvB/hRPstDHfADbzfnQlggR2lc8kPdhGbJ/lCXsrTAh8D917Ejhc9zDVTKVyIXQioQh
yH/QEDi52dZJwZYiP2uxmkavPcRYfZ1E7KdDEnKT8DYH8QS31r5C5PofIWkaOdlG91HYJPJ4D32y
OIrhLGczOcp2YP0dN5vIPIz3qQu9JilKZlAUTvBnb25JGbp9+lEvLBu0vksPkWkbRPDi70W/hTYD
4XMQQ32aJNbE6DaZJKN8YIrF+Y+bZA+twtes3yXTiOfATqUBFhwlW4yoK12aFCGoSsMLkQwPkSyz
aH8iWZ7RVOA8DH4fjUosmSVIuPwu4Ff5o52Z7ORO2fnWJbSQZfVcIY+ClrsEDhyCiUSoFFKV3/5N
xOP0nnlY1opu1MpFpLaYdU9mrqDIojB65ppz+TrSL6JOX8ldZB8Tidjq8x/bh8P4h/uaQcWNMGkw
s74sTyj1zjTd5ge1q/79T9MUAZmnYtPKhiw6dWDujyypNcIN1YaP5JMoBxNvHJmEOZefQaAfuxDc
7eUJgY9aGpZddbQbQ6dQcaz8UvXkJcbQsLHoMAebLeELBiR+bnOiMNMkvQsz+1dEFMpg2rFbieb5
XnHdMZNX/cB+g6yA0yR3rMaip4vpOWxb+GS3xbYYc589CjQ2WiS0puakE/SLIgQP2UiwlgYlICdY
jw/k7/ZC1KYWlQlxK7l4zMaN+zdOPkEutLASf1byRN8Vvg5iT/r7hxr7oiDXjzf4GkcGGKZmzByF
jVID6qU+E4KZha87mCOgZZddU144GrKuAPaq1+RB/xwvPRalYx94qRn288RTQqs0Trjb9qOUNzD7
idUYJNayf1+1HlITBkcRRlTLPrQoIjwa/ye1jv7UXKkF5Im1W5d9+WwFWbPEuGwn24oMK8mTHdkI
3uzWY5yoB1Y+FPaRcHwB+t0ydUHArHR9UmEqT2kDm1tgnrLCzLvx9GZkZPlObfTsCyilwikxirRz
j5bG9HhTiddXDbm9qqDqKFjQcOoFgQe07u05fj7/iumZIuVdLQwopQiD1f6k5LdslG62UFfWXjec
/S/jsSAzNNWJDjoCV8ywFOTIacrRJpv0ZzhNalYp+ylWOG0rNNFStf81K11Ng7heQ6B6+akXnmKf
QPCsglYL77hE8p85Hkieg6dSonSPr1mMYrtIjsgKutifxPxOYJmC2AvAuzN+h8/DsajmsLD9tZJl
kKpOMOu7wEwwMXP9n41w9es78QjGYlYmPHAe4NsCo4KowAo+DSXPMslT35vU4LEwjjMixTD6C7U6
D0pxe2UhcZVDI5cXerh8eBl2WYMlHfow2r/8/UNOvwUpD7vcQzKjp5y2sE5fBjwfr1cLwFCpMCrw
cuclhUuiujUQdGaBgEVid3qBWU2dwWJCqTGSqKjDqYR87IwLf9KRQZUt/mj2RczOBM/BV/eZ7yqt
5g4o5+9zmTHmNeP6pG+tB6M1hAA/Oy8cy+1y8nXcUm3TgGdQ4XmZSh1GUPFlEZ/vv2yxmXT3hQ3a
rh3KiqfOlsLLX+DU0oIcmY829fgLmBoBT2/DlKUWw8x4X4KzGaSZiVjNZdVLuAotLiimQvn9GK25
L73CxMtv1/Pvj6xfaJ17yh03rmuXA28xiLnpdtAkX+LDwUcfld3A9ylo5Z2WEqj6JMz1p2rRcf+Q
Lk6qAKa/gT2A8PIVIHgawtdkPKinwu+W2eXI62mjD53uxHkid3H+pHiOBzyz78OxYAYo08Yi6U58
NpLeQOVMv1tdz497r4qyux61RkBuIhQ0MPjHNYR9okS8AWrdog6JMgxbC4ZZME1m6x2DjkID2jh9
OXuTK05Mi3mheDBHoTPVNnJckswp12/GZVt2h7V40S3oitsy371O2Y2MggJ7lZBYM8BxzmXgsgV6
fetazwYUmtjTPSI8golbZvWI6xzoLFu0jC66dUArtk3IkP7jZgrfw2wgEbGUOfi5l1Zi7zW7mYRQ
EBxPDh7JfqZTU+XdtFmyfuz/drT1WRaS2kLK5q+WfVe/NPjpf+9G9P3eyygcdRRzdqmdKgG7WBfe
Xr1Es41c/bPtV4N+MahwpEUZbejffiauH9sztAVoXnq1hVWiR6e143QpGCiEGPFvuKU2Ocs9MIPJ
Ddj13eYy5r78IuTCQNMozhOxf8+WCge7kZZxb7y2458yKs5Z4AL0pLlMaggVJw7pRw5alDlTYK/G
OUwl/MUXBur8OTI4dnSC11MlCY506qd4kmVm7klqiTjGYu6oLtL8HbhfSjLwRMaS/zxRtVJUAXyR
SFj7oqw9/PzNNvsYCnIYV6hOVLsFERfBhMJa46bUuuzCCOKCDK2Len8qoj/75q1NfCXCMurIyL3f
6R3EzQeNPC5O5x6gUdi1YBXtQA5BfGz4a6ZvDo/J4zFd8EfrL5yjoQ8JADMVoTIM9Rikl6OdGCLz
bvLcDrWHAI6NOAoGRk1fLeJqd9Np9a91jF9e5YtUCk7kFpRTEYxSLUaN0IEYJFLhbL1iMtrrh0ri
gxHheOPecQPyCGf52Vqf6jiCGOqJUk9Ab1InFhpBa5KbAXOeR8V9RPWw5y87wQWSlUoj+143Hc6K
iZlNkNzqGR4jitdIm/SrEcdDBVbN8TaZwdEmjmGGcQW6Rh/8ADj48GLhRkwCG1jxhNXBZXbhv+AN
cPfmUdUBXpZZJ1vhSFyuRbzBHqTMv8tFjcyVG3Q/gSO7OoDK3EgsY9UP8jaTT1B885Jjb6oRgtVS
FwVUUIHgGZ6hJhP2Nb1O+5n2FEt3L9LJMILa8VU+hmv4RbuPJdSsQdLfe1/2/ivf3tr1SlpbRITN
3vbah5phG3DpnotXSHVpoAJk1Sz6/GHprKGxqxyOHk1v8Yy+gf4ZERx16AzD7yHnI3inAnOBlUuD
+ulgxIiN62RvZNxbc8S1daXwk2OkGrFcx2/TbPQ3W53HaktJn+oQRdMTl15b8NkOc0OGgVuSiPAa
9bwPXGp15LCw2ZbC1NAK+lhF4SFjKoaS6qWnwWq86AoAll6UIRWHB8MTQ+QzjOz3BNMy3XmvNKnP
f92RVdPUCSySnepK06FMZAd6fiagXU37+dIeyDD3uVOhtQS547djzLSD6vqgcbS0nVnb1QZWgLFJ
/y6/q1pduyCA6mrqcbSsznaOqImH3KdzJWPrnjIelVbzborypV9AfEZBgplvKTw/DmjDW/SIlmxB
q9szTNB2Nff5jIsbwsklHWVI2KkfZGbH+fWpA+/080vvyMnqgbWhSJtmFXqchA971Ty9gX+q/vf2
aP1fPv9FWwhnhtXdC9ebBN1BPtNt9uYpE6e27MkPbDKup0CD/ew0MYckxC8RIFji63DEPK4Q4H/1
NwfIyAvpGeUaLhhF0mTHf0FZ7HRpdm2YtFN1vvB4zJKxEvpH4kDYMznwJGVcb7I9AgfHAXU9JhcV
1hQs7eravnx3KzpBnQy4SDfeUGLvXWZFnmUBLp4WzUAHoYu7p5Ew4oxW7F+KOJ6iJnMXWsj4qfh/
16Sv+5Oxb+3nJNspub+lVho1igeL832HyTDb5v0JyWSJVknecI8Nr2tGdYvwNNDdFcId52K9hGMi
KWcB4WLQ/qbufZUD1e/IOEJibmjkbmYaFuxX9Pf9Jy/iefHRbU7eEDsiWz44OgsLqTIUZc/09TZH
B2RTP4oGj5+WC7s/a5C2wG0LwJb/NOIifhMlDgmbJ0RZP/ULzqct/2F7KaI1/W9MMimA/EWmLwdg
kWLjgu0Z5kXOAbYntDwolV+mGYPfZ1YkwxrRjIDN3i+8Q2d4qDRTexBxDAPP2riVwhdG86y2Q/eA
I5QBp51juxV9uq3YqP7qwzuVzuFItPeE6owOyW4g/jpKTijDvITHzkMMC3WWBZ3fhGo+FJ4BnL7w
j38j98zw6A1URyJ62pNYlwu3iOOPhN8uvqbJNWlT34Kwx9dnfb3d0sd63XQdRSoLTEoi2QM4NEdA
7cyNkj4jB1KPz5oRdApijdfdzEySmbv1v2HdFVDi8zvZjskN9rv22k+EI1On2PGkk+GQhIDttuWz
6GY0MBY6fdHk7/2PsY3ImTwqIlTz2XuUPCRKZG2+wl0R8SSOkvkM5QaLSJzXJGFa668HXlD6DeII
Ov78oS/JA8TrlG3JkEVex7K3B6c0+YvnTjTvX1Shvzd4L8QWLOT8kGKjqeOJFHH4gR/VmaHmF6Zq
Ks+QDRwmF4kZ1GEJP9JGNtnClExRT6AXrb5UmB+vC620dsJ34c82xGlCTsSpyAw+mvzgZqFEcerM
HL8ygb6hv2bsL0Mer7pat03MkTBc++H7WYfQJ9pqRP+WJvRReysOzSuiS9s8+bm2lxaqzFrYhHbb
WBbHclcryeI4UkUIo4UDpGSkN3Bv/pO1e2sdAYMa7kMdB6fzCu2vGN0QfzKHXO/LYXaH9tJkLyxF
NMjuKB8lwLqN+KzlHzgINHICTncntTVrDUhK30b5oXg9S7iWlii5ime14abXSFDuDqFZa5MnWP36
d1BDM1JdSq1w2xlIeXwSVAInV8ntddyEhpeYviDemw2kXUS7L0KzylwBJBVqJoPb/PcdO17iYnKS
47uQ1AdQ16G5IjEtovTctKrjQB2Vqr4i7mudeE1sJHBeFAJL5GHh4BOuYPjjqWST4Sw/byb9/Lqr
3yHDlhMJJv87rgrT+yilZMG95jJiwTBSCAsHCCUX2Pf8EGE1N/nc3On/RCjHsqel+C/2GGBli7ax
vPpDkN1s1R/Dn+EqR7onjzp+mcJuG5LGmV/2h8Z4qM0z3fM3ByQDR0lwIhCjOIyop5anw1XvVCbD
Tt8VmIUzCtHlwESomZkQTPCNoxysmzOPycvO3Gg6Gc0T/dygmWGYmCAxip5H+gObHFp5coQ6vYPa
aXymywBuysLl/oZkylOfTNrOqck0fAdnWGgLZi299ejDW0PiJ+wprO/I9axu/kF1LcJoUekZiHu4
tkl5Uqkhez2H12V1IFsTj6dXk7yslr2pOzQqGH3r/SyFMz20Tn83h3GKvTOA+nmoIGv6fGt08KcY
gL4+VcdIVNllLklne9lKBVwD9kTcKa+W18yQ3IV77o+n7xWBk2KRW7jpG5+n2U1AIjwSDom1mCPW
QhmeIVUnTjMyKyA5OOj+yhvbH0kGBaE3X9idXADyoMF5Al7kO8I+r/py8n1Zyp5kZ2HqZ23DQeYY
yii5a8OdZguQT4fb7gKy4kOSfw6aFY8QxHvcgQuC7L0VZw1kEI4S08EC/69TiNFlsyPU+V29ji8H
fX1wGvNTsfBWkshawfDi7+EZuu0BidnCo7OtIHPbLn/ZMo7HOJSavZk7N7rHulbwwKLXhSzdWE3z
78ztZqoxPaQMIZ1fwttWHBcz6/wQBGLQa0SDsWWj9z5/kuPO3ooB0Ypyt3XPv8uYbTS2zM0eJU2w
C7w6BSDTZgfODhkK8TppYlOIrxWrsdY8Na4DjOfLQmipNj32Pt3VfW+HwfsdLxSjZGC39pHZBUSM
9vXpHolUK2ZxQohgp3oLpuSwgjVixLtC87HRAw3JgTEcUlSP4rEmwNvrDmroQ8V2SS8E0ru7/i1H
IKxolc+/R5dmi1lOJoQ37nZB/+bpX9MABOcvfBt7YbMuBE2vGgqiDe9Wh7ToFNtm/MbpKko8xysa
2REWgCPXmGrH1TX/8sqWbFbNdDZ5/vayWw5rnXpWr9TsM2ti8SKEKKBW9KwYcgjGZJpDywXEIN1H
RXwB28Zm3W65V3gVl7Z4yVIgbnvdeQvgEiqxDUrO4Z31YYC6uD1ep17b4KpYuFrDz1YbXcJCaxyR
I17/MrqA8Rh+/3Gk4jq+9v1VjCnhUpi2qk08BYD3iKi9/kANTZ3d25YMr1QxuDEJF29/qqXfxyFz
lWll1NxCrWQVDwAARjWQ0BOtgR6Eo67x/5IuisteF/Hhu+cWNo812ohm9qTxcp7AwR9t8bpG8KVL
v8nQLBf26uViLeQmnJHA3M7bCOhm/Z7L3PxmiVyeVULXeIxHTe1SC/fwFzoHV37WweErFb97Aex3
G7KxllNNreT1TJ/6J7/lLY8Se/spdEpPjUSb5WFW3pv2WlsJNJGz/HBdoBZt2IR/hMngCWjaHDLq
UzUIDtoupOKiZYKCBdMjerm8X7cmowkY+quxSXW7hZoOlYNlWRPTZMs53E4vv15S5pJI//9ncmUM
CjVS+BIJpYt9dMBan00KnxwIv7LxKOLFnNlsS+4rHyW00oxUOqahm5lG1tp5xNty4cpuBdV0gfoS
7tFcd+kyKh6lYyqJca+5roakP40FaNB3jtE+XlD3VrpYD+iErGZJfLnz5QfTlB/n6JCNnmrkj4e4
DMf/BIWN3vX+Q8B8Uxj6UDyp7Mrogc/aiz1zsUOkwzfvOu8SeMh+JIXILFElBOOsy1mbdU+ryi9V
/rahjW7SzDXhAT96gREESK0F2j2zjPpqm0viEI/LShnAVaXtXvlB/73113UT1NAsBBWLQQoWd5B2
kcycz5qG5LLZEb+SHt3FzHMiCIzBCNcl3o4C6fG3hPtrruZNNiapwsIhKRBXOOtkC2Noab4hA7qt
Qdf/I2crINLNrmhTsz5vXrQHd8abcX8/SSJxmZ4aQ7PHqX/CueKY4Xuvxpc5/yMApsT/BwMxEZWd
QkEMTV4QtG/DXUq3AhoOWwxT8Xyc94oNiH1yAYUL8dFdxZeOhahCBI+h3UKTpIK6YXCG5V34h1sW
GHh3RWU7+xQ+nqIerm3oU77tJMeY7Dr++WzZqw/E1Rd2NucNxBdJFK0Dg3of3/YucqeibZAh5sT3
ev2Bd9OaVBe76C3KFzg4GAdzGddHdEfIMwyYdsEWiOmvnvxesn+nSpXNFTAArPgeHgbDP9loj2Hw
lJRY2BCTyl+OrS5u2rQHIzV1VQYgS7VPQ1xWJPBSwkVpfNggq0WKHLrKIN57j+BDm4Aknq0V99Sl
0rqqdCXLSnMVxtiUBVinwbUlqXCOkDXRuFPzEgUNYDhF/TNjr6TB0Vgvgss8m+kkSUaUpk5SekQA
wYCxXVhCD6UqILktz4JVdZWL7gvlIZ4WcUA5NsyzLPAu6fIXZPD0oRvo3LBhktZ8veHzGtsPSrsc
Ffud/eX5RmIPd5bOrLD1axKRwSW1AV26TYVbXJnLSz9DWU/R7I7piusCYTdlo+UHRBpLau3/w6Df
5oChRYH80cDAi/hmpVb4tR2W4ro2PfEIEbeLX+ZdEAgivrhb2g0TuS53gOwC15LST5y15/JJPVZh
pmEeqzzkf1lS4e9ReZUvNDMmHO1TfauX4y1HAN15IXNbZ+KhzjSGA3HCkADRBvlVEPJAY8JeJomD
tFYTPCdQnUVB61QBFHiM5R0fErjXOLmJGGxUx+wigDm/aUqeRjxc+oKwTv4+U7BjkqH/pqD3owSt
i5YXX3zrH7hNoGEcSg2fYOTs38OUgpKszQcyJOCyD/q6C+XtFa7hq8yeiB6iOWDYM+uv5ScQ1f80
QxwLm5N4plcPSpU7uuuvDp5o07VdbRVzt/2vERpV0NHkNkA/2vE3X0trcBCaB1X0+RMvq3Fsax6b
Jh9WDHw7x6wCI4VLFuTeutZ/47OlRSvRTwCWyS1oqYnqv0bz5CXc+bAaHFzcUSKwLwPPyZhGFIYJ
g/JoByzxw+9ufAcC8gdE83E9ud0e1f9suvdWq3Vgjx88WaRfixB3vVcW87RU/e0neTQ5LvUjGmlG
FwQ6+0ZwBUf3aP6WMMZojHEBGbzznO5wJg+Tj91h11cB3vt5jsoUpzZu1P2nt99nK3Q3fo/CsxgF
KxZsr4R2sKh2JoruMNsGD63y/QNKwevV++F/GoTPuDlEbE5kug4U4sY30eb6Gy3c38lxGdRL5Rcq
Iv9Fl1D1MKacJSYdAvEa98677yxCVsHqnj+b+YZ0WG4TJtRqgkg/nzvkFsACn9cTcqsBCBj6Lgoq
aG3N30L9pSSKwmP+axCS1lMPRK7eQ/hJaATaiJf/wgozQW3izYi74m8ufv+afKXai3uRtJ+jJtiT
qStekCDgmQNsQC/O64953neYtEgsV9KvpkCn4PdoKvjUE+hYpW9duWLfMh40Gb5AEAVmn6p7SRJf
Xx/mrtTLDhozZ4/ASm6sQsA/Aq4SB8DfTR0YVrd5k7kwILkyK2Ic1gigw7jZkJmusyAVw46B0VB5
dtIIVv0xA3pYLk+z/GvXaZok+uCuqdtLtGjQOARnWWoZN5h+UUvLrNAoQqoVx1hYQj4q7UGVMwfj
ap1YCP7gwcUn9LLjRBMFpgHAR1Gh8HXHFExEi9kJOlixuvadQ1eIzzADJ3k59e5Dal9Czkng6FvK
sbXA90JxGeLi2o/KflFnSTqt39NFd3ronmCIOJPXuCxDmDsqGhfsgP2eYEfGnF61/5ouJnDZM+nG
hgXg871XsFdSnY6Y2H4g9nuzDhW8ryXKNkjDhLudGlg2JYeFw14ho2nn3dVCHXU3eLA3pcm0URdz
0GBjNlwFTlypySspB+/RCNPFasoQ876qQSNqfIrOGrbpZLwkb93LnFucNvZ2hn/EQc2aEQJBtZLC
yRmRsK9d5Ls9IuQVrCwPl22ncRDpGmIcmDiYPEC8vNVap4Tv2tIidles5BwBsSR5P/SwYFe7q02I
CcdLsC8+5SAgFoyOrbNfggyD+7y+WXljc7agoH0RJ0W8FrJBpNvUIroIPg5PXAdFcZL92dfcW6eV
APEIgOYkwEYzqASbPIS1G0LRvUx4cFiWisM/Slndio59pCDl4d85J7JPj8+dRtczHI1W9PuWNM9O
U3DFLXMi71wU2sibAXXkaQQQLS/L7BBbWlNZVhS7ii+sl1NcPuPW/zAuZVkq1hsu4oWkC/8IGDiC
KLhqAhHsUvXs022dcGavZ/4MyfcIF+NQ6PHGkP5T7iItXHNms/CwADEBWdpXMqs5aITEK5T0Cl4h
qowWtPyccKyDJMc9egVv5jflSmt+4/nEZYdIhIr4f+BmSDkSbvnLZYCsdURnb4XKgAlVhFHSw6IT
bP5REbs+6WDcY7PswZulVjeVa2oY8XkG1nLS7wZApCuNaxY0Cj0ajeySSR82XE4lh8Tnco/RBHie
P5HTiiVqAlHxdxismaR6J9SIo8DjzkqfB7o+nq+A/JvAXMWmJVe7eZ+3gj6ECYDW5OfUZKeT9Xbq
bG4ysPZlebdDKFMDHR4laiOjBr+3XPjZny1IL1SPMSKCfVlZMuIqf+1zRjBFgpx0CgbL9LH+LWtG
vBlYhiKkRG3/AwwIPs7dUqIBaFR6mUNWGJ0Hye/EVcGOj7PETrSDJvmWbIXj7lsF3+UQSrXdBswx
G/b3/roHe8ZXpi2ER/xo6a59bW5xk67cs00C2VuVosa16GJrM/VUHx85GdjGc6xY/fBOSo8R2PZ+
tK4ys5uvszmJGE9XR01X1wpJZw+mtUaQzfhXiPRdhglMaSBKaC9AKB+ZcwdvjXuTPHQq5IVvLm1p
ilg5LgBcS5eXNXaU+eceICNxSk41r7K3CZPs/TiUtkkqSjEyUp2eAYMGjLOUmUITUU5oi89cQN3j
ixwRkM3UQw5LSJZyWzRqr3Z0yfINzKVYWpXk7y5lopwOVQz4Smv9cKHs1VnCsQk9wNWL/YD382bQ
6z+TlnwQCX78fV9YkDJr1fZqahNMy7HsBXedAjho4FoF/i0hVgScNUP9tazbBOnqGV4Ygm0G29oU
VYCskMLKFI4UP0Y/rFe1zVZxghcK8Qnof8wPV3/fnaf8e8o4j0p3oHw3qPA2LLpw/R447ISlCXuE
gz2pxF5KDmhhK2E0ursov4krOWvaDHfO9cHrfiqX/MGDL9+UafZQBk7qJYixNScxZRRYULs+5RqQ
sCvLy9DietJzWDGKbILtVyb7fOjcDGbiY+QnXtoGJ8kBON8DNLTTId8Dw/f7veONpxwFPyE6e9ZM
OIswT3+Ig3pcmCMMrYnSyzxa/oRQp5o5SpAYivy8op9i5kfm5MXPMB67S2qC6tGkj01a/YXBia7T
KGGpydlVbyOXTJ5PM6KQrnaKZpN3zyX3/4Ub8QLrroHSTebZXvBqtpFpuuCbcdnhRKDgkHkVVWwg
Wj0cIPKveozg5h/+j/4IeVN1oTg4CbUziifNrOG6ZfC5F9SAPTjkemXEBokjOAxhIgGX1zJzQs4U
vdGbiENUoEV/JayPhF76EkS5HhFQF1Zq2np8iJXP8EGHUcKVaN5aFbJOCXwz2uabJpfYmYo+x1CI
apLmx5VabrZBlCs8hUtlPQlyryxmlQ9waUElSgsG6aVk7paHZvGEbz+J9oAjFl59Mr2Z1DkJDyUs
CCvs4iQjSBYzsqxIstl7YgSNcKhJ1LTYwI7zjbpLhW1sOv0mtaCoN7aJYWEPOh24YK8pR0uWspRB
W+Ninr4WhnK2GpF+JSE5uPybRm6Ue3h8L79UY8vomUK34/xv5P1KcL4mxKPuUn7BMXQ6G2Gm0eE6
uJ7NyPKOSCCD93ocs+t/ZBT06y4A+X0S7QIxSpyqVFAvfUDmWNuV/cXTl2LaonndLZnMwO+4J9NP
IAN9J8BBT1aUnUJesjZX0P1Wf8CNKVZpOJFOW+UO9Eacx8XrMMvods/kPr9m6C9XEE+cDnBLBK1C
uqHIN/GPPwSl+Re4MbOdvBmcxFpAxDzLLMuL3VWnLF93R5kb2qTZpt9KAZbqcZfoRXFuekde9CIL
rHm0w0JWErerBc8e49LPA5sQAxF1E6rtvcrL417JvRlKPNY3GivOVpbyuCdwJuRqgpdaOjBxW1M6
vaSloh9Vfadjyu+QCrYDI5fcDcHnPBooYZuFDaDQM351hiRs3HbSwzv7djWWSqulhWxcAbWbtuX7
iLgYuyhw5XoWgNbbs0HorhBWC4/+FNLkNefKRA9FGg3kHe806FnmoPXe+pwH0z/hrFCXkoBN+Yi9
CJyHtrBCiepgqwixFObMXvzKGT8ntA+Prq8IVzXP8yNCf6S6JymR/BXkCyc93m0cbQmNBJu6pS9Q
fw+GhIdeZMUykgLUC8ckqmEAE8xQogaQVvc4rm5Hn4ITP/Ad7fiutqddOnEF6xxLBLMXW2uOZ1JJ
6nQxxlvA8sUWuFK7nUXFat+EHPVgEpn71CDaXO0nrvimyVCrFwGHDYeEjX5VF47j6rkb4yIJDAem
Jznynlb7YWIHI/+ABn6k1YmN1orbx1C3a1NSe6/zDdEr9Fg//Y04wAHlt2sUxCqjOA5kMBucVBgo
o+yJ9R/WIJAoU8RJ+GCAwUsSiSghtw+i+k6SsnM6lrTsdeDrnf+HKV39MjUDohK1sTwztEernzpd
SEbU9mXu9PAw7shISOd+CB7FVG0d6Er+6UJEVs4gbb0p86/YlHaNP0pTRJQM5wenTXUC+nsCngDQ
wnmr5NOWNwXuy0yh7bkob3y7UsYrrqccNljuLqhP2sA+wGDf1bRFhZU1ihZbH+GRuz8tJ53ZrNdv
IaqCwXoaOoeRUgocc3iUoItEoB0gvwwn7YB0/AOnswU7nWSa5t/1ZIw6guJ+xB3Vge4LtYkwvxkf
fxK8/A2ZZU/1XSG6UucPaA2CrpiW7KEIYGLVtu0OhqIc5inNbTyBB6zC+8UPm274UBqRHGDkDFe3
7WEGn0q74RBJl1xOQ+b/BYqBVevq9sUF6FPwQI15eN1FnumYigldvzhd+EKBY1LVetXidc7/BHQz
pLaGt30S73Jn6G0cT9nLHD6Y1YyDJpZEihRtyTGDqNN6bkr6zb1d5GYLEKzgXUAHbLb4yoEf1kp5
migLIPFt0PzmCfLQyy6HNk+z1w57+U+QahyxUKdiuB9fOvKwBXVHiRZMgqpu9YnCzIJWeJIB6WlB
iIrgI548R1bjsG30Nm6Om23qxNiCExI+W2Bn/npFcfJPUyoLWT5OoMvJ5kB7P85a57W3zIN5S5+G
mJWWHp/T8Y25Moqm4NVFXZZh0n6GiUUlWJBcWgewei60Xd0JMoqcAjSj9Zo9BcDI+3uEqjYsZGye
HH3BzlvdbSamZS4+ghdbZSI6Ull2rPvFyBiEfVfulxr63EEcQqSmeiKh43UwbHLzw5gpB7Y4BF5L
jEjbsaNsNGsERph1G2mp1KjRE/kxe1seurSRvllmOvVsle2si6DzZU+jlT9bDI2bat6/ifduOLl7
A7AiAcd6GROEbAY9MC3ZEOLjkIwmAqMcGn0uIEYm44Z/re3dNJQYp9gKDvEwJ5upUPRDNpaQXA2D
quBfV78hNDx7ZgdZ5OG9aKMVxDFf09zEFu9KcozVb0lXroPIQ4RNcy/5m09x+8EdeEUuvJq9Bwef
zQonI/ZxbEjkjU4dUMwVzEcz7WINH69yXjQA4veCaGysEuMxxu2rWw3Iygjrq8gNvBCGV5xoStLc
9SexcLYGlSWH2QaY5j0Qr6OBV8cxs478SdsUsLqQ9RfhkuiayPk1CpHyaWblC2ph8mjdSiXisOX+
FRtnG3WIbauoFRHAJuSz32ZrOhyxN1xmScRrBKMSPsqhcq05Ezil9bei6mS0Hu+PXFdCDNoJCq9h
TfPf7a441eiLFGsqnxDP55BT6cF+0HFFEC8WieYMulA8mll4EYv4HYN25huvCgNEHQ31Hx11Y+ZA
16EQ/XyUxxHa0bXmCC44rC8Oz7OKr7fhU4ysSh0sRehRWa4JLll0LpghFuAQWKPtL1ysVDfcy7o1
Gf+NcSZzj6lTZgkfhpIQD2vqXopKHYZRNrHP9gGbujrIAuDFEIhog/Xci97DYu8wVoz7fCuDvE7C
8qDsnOjxEabpkIcj9t7ituuixAOD+xy6ApgASuH0wEC2abcSCiTgu4wwd6Et148ZpDO20LqviIFQ
+6nhNXYOU4fxrj3Sif47tOMTZ5cxh2U166+tLExETSoYF+v7pd8cnLdVQpQGJYfnrsqAY7UM/NRg
nQUCCVwzdliMZoIncUfqsOVgzDyN2bB/iuoaXfg7Kj+tbv1rur2BRvqbQUfZ/uPoBOE7t6cR7vTG
0ndK8lizQvcXPbWieu5uA7+dmFktcKXmD1wX+TPlg1CeKeS33yu1m4s8ncx8aHdck5LzcmMVpy4k
I5jb7uqwDRmD6wm5UbrGm5Y6ByZTS3YYYvwDkSqF32aCeYCi7M49z6r+SHGdRa5mULgyP97y9If0
0q0/pDi+cT6BKJ1eraggKjTUgeErmNxV5Sm/O+nG8b3KDaT1mgvQKa8YE54sWKuAxU91T755VIue
9UY9JvV7jCwWEKRxvS/1HLJqK6nbDBRt/39F44zht5ZzPTSLzrHMBWxIKhls8Kb5Z9VoNRCLKy6L
SN7if33s+YciORdrxDof34tnC7Ot7Aih4zP66rA3qvvw8aCcEN7Wi0Q3Smb9SA/KJPQjvn7wO2oR
s3dO5BgjDcc/sRbbCFSiPvPgg0dNx/7h82Rs3D2UTBwUbTMB8+lG47sUWNMlOXdbJXtm3FlGSz85
pmFvBeeSN3V67T9kB9W3qfWqaZ4kGLFdLgqhTukEEe/7oDszMHXTS+JD+biP0uiI8wrQ3HEA6sQT
/rCR3jp/SvSgV2N2PRA4CG3TvGZFYL2sJlKeVaOarwL2bXZbscJ0A4jS0wAs7VBfGmOtEWPClPrM
9TMLUF/XjhqTZbPxK6Qio+1RoBbLvnAbmXiPPXsS/UMDbROLtvKfYSDD4v2w+W/mhYUXyKYoPwts
cbupwj3/QiMdRaIh0LsUWj0Os9k0/1B9FHHzevGIHnIf/t1yuS/8cJ0rp3nacdCn/MsZbFm0TZ84
f1+umvmkX6VmFWkWiPf0qRGgWj16tgeHpj+8LqEFvH60SsMWrguYFcnyT4EdUFrSEbzwc6LVrN6k
Cb4sqUUzSlpbYTXtd273GA27auuCctsxX1iuEYUYiKxUS4j/GrPUwp3dAkNssQcTaXPkb6b7CrgE
NKIGQCpE6CBb6b8hcKJfG+MuoMOZVYAx+sYxwCsK8NRR2Dm2Khw+tUw+S1f6yia7BXWb/RpRQzdX
J3MLDgzyJE3pefacB1johka7D8CcKpMvNJvMbY/A11ywTiRky5ZvoThsO/hi7ACevM/FjpIzq1Qd
ydRScqk+JUp/xnIukHJX9ZqkXliPoJiLz1JQQdrJc22VKkktJ9mqdsIZxyoy7Z+G13tZEpnEbmDn
CxPf1bXOlCgvGq0NRoiEQOGtGx8BytbZM1dN03kQQGWfKOaAyziuLny7qEWYiHkAvYM/03caJBMp
b1rCexB1ClXEdJypmCzbOieCSEJCy0+DPzpHbRa9yNefi8tEDv9/0xlh3JilIyxP6ALHRJCQ7W6o
juB9Khf1dzHsSXitDvH1wbGEONGgi6Kl39p+Z0jGTde8K6A8UVI4xc8bBr1B7VwhYQ5A6xbjHedX
IR0x1WAsB4yk3JktXhgeIo7NHvkrX8hHDtOZbbXZf/SrjCgQMtE3lz7ni51zfAemOvLvkgiQyRNc
amUzcyLhmQPJoNpEtUWe+acOkit2Ysd02U0jelzumItgt+A4R5SaibY6lwuOnG5fvJKaIt9LO4TH
9SDrSIhjHhPBpzAFZ/g8sH/Tmq8rTWpKdmgLnXWi3aZ7HmrR7NAlwgMF5gmUCNxPLx2RH+PW87zL
s+yX0HSExV5qwYQj+9koXT+ip8uvkxZzYLa/LILXDwB3jj9tAe/gOybiJx9a3x+I/J0y/d1WJ1vQ
gZs1JY+oYjfR/f9IfGZi2lKfMc/WBz2aYnCM3LGDQigc00upShH9Bpr9lOaNRXtV8hSZ2p+pC29v
DgorofNqWLpTEOJtya9wupImMGOqPVlK/N8MKHAszuc6Q39LCWvW3amks2F/0Pq0qYSCR1r56LRR
nYR5ZxLaEQJXwZ22ieaJ3qGFTgRWh1A54QV0subAkf7jWJm79v6NTdc+hAdRNzzWr6D/Bw4aoO8C
myuOEuoIuLJkek8GqK2lii3pTJKrBSzAmyB0C+qyaT3EKNpQP/9p1VzRPu9WVl/+2v/dc/idTXOj
OeG7qpIGYayliCDZvwdhe0sY+mmRfumNUBJ+qaxsC8P6dkazEdBUrrL38rCujdw0SKmjcdXkRwBg
kg60DQLugFbyIUEsrsXv+Jay/PE+mM1QzYqbI1GAy7BUXR3OLHYOoQR9tUMYR+JFL7x9HMVzYU6G
dYsQ9qZbhqBrS9FAOel1doCWly78V7LdLxySSggAEEhhEaefSLDr3+jkxWKEXkGSa4X/I6l6nyIM
5JGP1cza/Gkc777BAWG5ZnDnr18QYEdGNZFw4jMyyOjdQUBUXctAslW0UTvliAkC35hmLDAMouJd
0kccWiFfJ3IV8WfQWqfJsifapoAetU7dDGsAEoCAkpTAkljlLNokgdFojcsvW9yLPmb5iCVsZAnQ
oE2PhWJX2InRPlfdpv8jXriB52v1ECKFUKQ+htzFiDWP+rODDX1tfA50pX1VjEpqNohAtSbYn5Er
GL+qc2cR6oJ2u+dABCRDysclbuz+nRlNwctbInj2IhtXmuOJgtN3AmnTwQU/geVmr+sNWYkcW2HL
/uleFFRa+wVaqJiie5QoZxXz7zlqTXoK+G6CSLntkdQwiH5V+CwbHdsr0DkerMJwYZgi8V/3iY5e
JFxheM7ZYaz5/N5zcEqY2uWAqpQOEWq4Km6r8GLkMXdpPG42jD+iaq8Ne10i37tlm3z7mwqmTCgQ
SslBU0wfOLp0BHxNL40HxOM1QErH8/hai/+n+xjDXvo3wZoIWDJDF/tLY9sQz70nIqLTsz3yoY/l
n4Ht6wN1Djfx7ezOjHbCu8Q1oeTRLndSVsS4me4plqMZoqAP4fcNPVrTVA/L0s9jyMRFljNnOKIR
hHTopMAOe82xuaBLjYRQfptutfcwicaUCIIHbF1GxHiBjAGL4+P+NH4TMUC8IWOPNuCwh3KwT2Ko
sM0I5RRBWQ2XJqN70kv6gKTMF93VitNJgZPyBpKZ8OXpi1QBt/sSQ8CJQpiooU+3XXn7QKuWqslZ
LYA+4r9ay8V7LnrG/YjDM2jmtF8kLXFXyvL6Pbv/AAgbRZgWkotY5iECdKbrBwnacnHm/vqTjhOd
7pcqq85rVUCjfbO3MfWwg5U8Lzb8OjENXUqOUBJuB1cMAQzTu2HgmPTf1Ks2WtJ+zLpAo7bHYQzO
wYSOuqWHafB79YtOHAPH4PnqKNkUAEcmm/snfEITybnp4kmGYj9icq6pxZz1y3/mls0vV5SHCpy1
6ZJi6tHyByGXlKuG21W+0Yx2+YB8EmstVM5ICZM84EK3bYtx6VbadHfzbFKvwgTDDSKAo3A5c91E
BSYr6UtzTwU3UZ1g/GmC4si0PXRX/ZV5lGQMuY0Bz3c6uZcPmFZMxrmfXvUJFRM5Ep/EujpTBqvj
O0lIMFzzr83LYGJ7it/J6VIp3nUGegSCn3KSnOX56XCs9ETQ/WPXMgBiBEOp8ca+TZa0gs1GABG9
r709Igr4OopOrvWsqyqhYoU9+aaxt2hHOveUms03b0EkHu5C2ODrOfPBsoVxNPMIytGlJAtksK1V
8N7N1R75JgyChhi+0pdS6ZqRoWlcIr+82KM1WdmZWFzYLxu3nw+Dap9LMLU2vFSWyi8YMkIAzhIo
sNv+ZtPwIwSUrt8HQ88R/uGOJ1TY9BrFfy5uEsTA+v8I4+aiWd+BHqB3Wv9ikwOqoWTbPvtJw5gk
gcLKhkYyHsP3DOfPa4CcB10MjzaV4xjp3kCF0t6RmaTaj3VCbfIClrVIsL5sRN1hfu8yEnTi2vPT
Fus25C5OpLu6WSh3KNFpGGIvQyLr4uj44hoAYd+tXP4agdPYpD3NKrPO+PQycpZPafSNFm0dGAhR
DBE3DaqIW9zl4r4KRXgLkeTo6sOhZqoWwcJ4Dhgj1aO26ID2lNtEx7X49qeyAk9QouKTkn5d0x4D
GHB1df9zhsK+Ui4QPUA/OsnMqzWg+0j+2acdnjdpP6MIdEq+MTY4/G21VSU1K107Hu41aZt6ZrCe
Sq0XFqrVzUG69lm3FPDN4hV1yRAf/y+rFDto1Vo9XnUSMBz7dtrzAyUoDlb7YQZ8qVigU1+cnb6A
yCzDuHNWiEvYFZpeIVKABfOCKDn9jQK9OP5NF6M1FGtbqUdEZLBNPFzwr/2eltVre5AsDNGjmvkl
wx+Fcpq4XliYaH/fNOVVGHHJPK/0igR8IclRbd+PAgAa5FCWkpM78XlBV9wNIH+x0MAbFg12oUOO
ZXNmT48825JTnV5BfyvyMUc3IvPReyQVPa7kWiIbrzbCCoCspmu69QHR+01zq7xvmoVj8vopYjGa
deZQ9XQ6845RshA/dILJ8TQs5R+mkd0MWlAp//JYpFWqQFd+y1XylYm79W183eLtKOIte4456RDr
zHzftweOOERpzSTgazRmKIP0s6EzPxPcGUu3Og4MjFRY9fOXl7HTKigo8b9kHlwPp1fuGNPFkBKQ
3+SoYrn/fHkjtQQIdRp3Exn5KU2HvZTWZlNocu9Q9+5kkj2189+cnULH/7aKXD7vhHwzMK0cHuHj
vjfGNJWCUgp5k4BqnjWFxj2cZ2Q2hpf8hKtKKcVz0wx7QkUjBQGfX51eWTMjfbzX7/vQew19oQF6
7Ep7KwvLM5LO9Gywhlo47s3a+f8WOeVviprt28skzHhLdmR2ohhGUTdfPBo3LR3bAkiiXAHhSuf0
8tGzqx6ET92dIgndkMc8bP5Mqj2EhYE2LAdmSXoDyQ3HtwxinTwWV6wXmvhulVn3KSrzv9B014io
qVeSZfm96x7PNfoSc7AfWa58499lXNymcFInCGsF54DFIPyeN5Uf1CNA9QhQyvsTK8MefG6xMq13
IejwQOSQL7HvBl9JFAB82L7TGOw54OsCZJAHtozY69aCEVKrqk2P4LjROQDgaZdLkZqafEIycULx
PKBxYgDV++p5f1X0ZGpWZprsJrxldTOjV7ou/XfsWHzQwbC4NmHG3QRaM0Ex52U/k11toAvqkIq7
Z7qPm2re3yd3RNyS2AmgP00dCMN9BdFJqHNRGDcg2YJDcmBtNNpYQcE3wc/rKsVFQ36m3nRbkxTz
Gv4VcJh5PPUCwanrfLXXJxrR8XEgpKzIrktVCwndrAPdH+RNmXwA3hErt8sb1oOH4TSqR5bF1yDp
RhXXzeGroUNuLLV8jgI4DhbB7U7wmBBTJiOR1Khd4DKHHk4uUl7EeW8VH2IXo+CyB3NXufXrZLEC
9sHzguPVAFh4sKP0BKAxFWpxo47Tp7X59epRM5g093fDMuIVSOL14PHapraVRsQIbwbp2H57IEks
jlrpOzYl5kp+7XldPDcYWGGWW02Bi6bMa42mmNQKZvZACHQuVrtNJC97PdVHi6Gfm+Jf/ps8CYya
HglgB6mMbwFomi7lZcqRcPM0iNACkDLNDh+avkfJ5V3nwuJSxruLDt2D4tQ81LDRyCbJamTRQgeD
RhxCHDx4g9159QaAqUYQpNYJh1W3WbJnaM4RAD8znJdjdD+zSKsc9E06+46JHSpS3QAQKdnJum+s
h3cYu9MDO3YaA8IJ31+fsZ9tprZw4a5shXlX4Zjf1ZpeSC9sGpcY44mdZ21iL4IZf36xCF8VQEDc
e2oyVctbYyTrTGx56xCBXmGTg6A71G4HE5ipgQiD4MWrKIUlUBCxEwy5UPe3rLnSZoh1+X/7t72h
+0KjNi1WM7J0unWEEHhKZubBCPfQav7vWCac1YXuo3gMQ6ZXrt0KBP6+1g838aKgsUZe1hPXgwJN
gKLEp/HRZzGP1qTUwUN6OQW5JvVoQbhrns8HqWJknbQS9Wj1D07L/yOBjNOYJeLzEoK9PSAa60tB
hTKbDCAKBeIJ+P1z6wtwkseFgAFDBtIBP4o+ZycQ7FXjPOFlsOrmb36WkLR4eCfi0r6pfkZXJIPU
kJotX043JKxGTukgbjA9CllykylwZCeARkGahkKqvKtmLkTUR1xLWy3kH1pIU7NGfi2+Ap71Z4AU
Nan2pcrSy5qQfoHqBJ3gY/09JtjNyhvCx8ADvHQ2aAcdNMyAA+evb9UQIdndd03DmFLd/O0fhC9p
4/AWEvzEl7es6Nn8n9y6G5o8DarqzWpUx/3qbqzVMstF5R+39tzyijW1U2E9ofNpbtjV6XZqqPm1
BTxHejMth8TRy/+yGreNgVWF1IfJUHiipepn2VA4lcWyhk5uI5LVJMf3TJXFvv/iAGUEf29qWuXd
SSe/jPd8yjrlkODhvlPE1iwXDwLaWu4I9fRVROl0HtEXyxkEIgnOwDPd97WKfqqTvqDY+/Co8mZv
EfMOCJN4BBuR88MC8JLbqcKVfYM/lXguJe31ErOz9kQeC5v2Pu4drT+lkqii4Uu98pjyKQljeIXw
MRYprPuPQ1PHL76cZteqOhPQ4nlfgtBRUOwN3ABlTjeuq5aI7HBssrnpvg/yoZG5NJCDHxNCbeG7
Zm/wOS3xalfmZ3hJyzxL7O9dtbNyX7PHd0cKNUiZogoOejPnk6s38WSk7/BuFwWLA+ERUmYuzeql
x/wolfl+Ev1PaXoygPHKbhdsitd0u5fpEOBhSXppEK9FVNJ2QATtKk+JBPzgFvymAW1amZvugWpe
joWbsB3ULWWUTDKlaxFgnuIgv/2dceppka8a+6Gb3cIiD5tWy9ZykhRO3E1c3WWH4y3Lb+zaAY8J
FG7xIayn2ylyTUE2/0deBdIFS+obZghNH+iQhwnGkEvHtedYO4uPfN50GvqCVDh4ns47NeazzXIp
lgioR5mfo9ceZL0YVq/Ngl8KWi5YDXc6mMgdxjOGmcHbCnWr9V6dtVUKJJiT4t2E4WfoeuKJONcw
Sv+nEc4D0RXXQqFkQhXdIYUkbDRQYS4iyqj4AoBnt9Bj9HOCICNKbrH/dF0a9xPI2tl21o+pR0RD
I6OKkAhoge2DegVdORCtlLB6bCot4uymG6HlbURZuCqE+TH0Hxu0nFjlHI/THAdM4PxVrhOuA3W6
ciM5UUYJDE48VqBAjiEgWjM6oQRD+GrYCajsNBS4GeVay0wgrgO74TSZ9kZ6hTD1eevNokUtaKcW
dP0gRHNbV2DzFbJ3eHASrwomQv0D8KUm/T9B6JpzHgger0mQfpajKW3g5DoOi5QboWsNu3EkNwTN
d0wAFZ9bJyIbv3KkWswgjHQ0kjabMgEwLYp6Au54AAcISfmzUlWrV7vWndgaBB55sO6FaNabCs7P
YBeZ2WBgshGL7aGL2aqqEOIi2UJroRuHToGLHvk0qVX/eTjg7UdihqsdW0hX5/qn3d9U/3tfiTfb
3qRF/n+D9647++S9Xr158xkAB/l/FHZOOwFSmsO0TvWAHlqpuClD48s4yqchZARyXFHD5sBUnX/Q
4Twi+BwSD4yYo6MXM0LHxfU3C6CZkZIjxDAQ/33ppLui8Uz31H6cGJoaBG9HD8Ge6QuBJD/1cWNB
Fa2PUa8SnzO7LjyEAAKhhgBREkxpn+eMZrGQnqJKkcAyy3b9U4J/q2/L4Kd3Et5FtWrs2225wj6W
PxJsCdPGOGSs/3NER/UvfwXPbYEyGmktjXm6TmpW9MfbZWKGTBAr9iM3JfI/moJeTVe6FuNau7L3
AcnT8DDadI1RrZ3n7rnRYTv1Uc7aKSSqpbU20F4r4d9EggbF0S7D/zqb8ZcFXLcajbp37n18gyCS
9IoAqCgF5bnRwA8XDm2Z+gcQBGaE8V1LspdYQRLfDBQVjH5WTge+M/dHnU3HGKVFeHFFPG0J8WWB
RWXO+wf9RsvLGiZicBo0KFyjZGleSOEonm9kznjeUXEfm5jL4EufhebHnHwcl4WLGXhivXyAv4Z5
gR3FqNpt1/WzsEWoyp0Bcy+ccIGHWUvs/G6cKQBmlXHJSqg2Vew+2KBTrcEQQlpFHrumgYu5WRAs
JMY9Wd8Dh+8U/iLfSgB9rJrW46j59oniD8pUy4jOqfzZqrXREx8iRaBHk1R8/LMgrMmpTmmSssXC
AdftdaeP51Vxlvwa6Nvmux4Tf7evCFwlq2eJbofSYLCsBPO43C0rH18ZqLCBRTY2vNqfkzmwvQoi
zMesvv7ATVVm1qoSy7lSxtT3MwvUd/nC09ppeh0V1xTDtZh8eZ5YRNpb4mXETxbodEqYVO3aaTHP
5aueEG+bqM//9FPwLrHwXv5GAS2R7mJgxWsrACX5Hb8Inf61F39/juAlcWqHzIzEXFI47H+rrxqI
nWcAR9JiAnc9xWqATONoKOpEe6fY9wxOu7ecm/Bgl6F5fvMYWnS7Tcy+q+UjyvMdzx47pY5kiwHl
lZQJlTRYJQWSEprjmVyqTIOThiiYZemRErQq56C8h7SR6dwuB/MLhj9Jll/B02oGt7x9gJZBlHT8
dYAUKz8AJRGjXpUow6U+VM217ukHJBpjw6fbTvTeCvhUuhcxxoBTL3ZobLe2cqLdkx7hxHBabmCm
E9J+f0i/b50GvknjTNfb0TYO8uEK0AAIvkjqQ231rGQLcKt7BElERT6JV4d5hrhfDhbKglo9t/A4
GGKhE7k+TxA0FJQM9UzxhoCFCcAw+KntF0dhjmppjqM8X8C+Yz7llzO3iR+DAkW6UjI0eQxluH1Z
R3tAoTEaX2Zs3k6VVZMrghRceV+HaLKz6aqOHW/IPXvmvC/qfKUD8CGmKuAp2I7nrq6Ak/H/Nxfb
jm5iFer06s6Z2+r8eIFwacDMS6e0RLHgS42odoe6/j5w576Rq01Ws/AfHJ9+DrYkk5ZNhbFOHinL
BmoyGi/KdRsFxJ5EN33AAIsFFW2Wqy0GoDzI4nEgZKaOS/656tN/PONLpaVY5bPwd9kdviohr0qV
6GdBlZ27igxXT57LLHk7Bcj/jz7dpSrgpEn8QMnmiSMi7LpM8F9YRiyqmKNZnTho1EmWfeP/KpOd
Ke9VyzTrJ/uO3mGhqc8MybFgcJMjfjIZHttWuZP979kRWvdOezKf6OYzrmiOU+UgK6G50kUsebVi
B5Y5h1MvyrOnTDIlT9YY5wf6AGIIuCxQNDPd3reg5wH+cjO6mq8WdTdsTGJcQOK7LyePW24OPTvf
MgHyBy78SAlUy1cOhrOIcPk/ECArCQm3VfE7nnSWpCNSbungkFmnuO6oElABvN2FfV1ou4Ob0eGD
0wX/Pljs4Ai75sj3W3RwKMOuuHSu2kkdIWNbyqonvrmcTyL5Vzhd0Grq8WqK6gBu33p9vHm1NC0O
eRQqo7yuR866FOl4l/pdBC7JMDvQNqb6OlvX6KIZ7joG34heEcwNG3SRkh8MfUfi9DuhRr+hH9yg
+5ogf8CBORZ5qJTkdc+qnDey+wk8YEODr9O1R6OR9S1YP9mu7OkyFFPHEJ6Xpw5EwG0GqdR22sNL
mkkbQ8bn6n6UlviV5O6pKGO36L7roxFEgkY2QP5U2HFJHBpQceSAlzSUGVMo1YA8L/HLrFerK9j5
ua15PnqtKO/TN04ryEgvttgzz16InASCe4l283JLjKKV6qbFToxT6epH77GL/+gS1QjJdLvKmg3D
gFvuPOTLOx1cXK/woAD0PH3cb9J8dvgix4yZYG4eoNGLzDx9de8ZbjXoWBekiW/SBfiKe+4i7S68
TB0y3u3GvJZc+Pj9mcfOQzfWBnrODqGPI4fbHRXWAOgzdU6bsHEWdJ+b7QP5L/OY0KyQZHDSHdn0
gaoyFQs0AMwzGxsYR/qnDidT15uw3hY4li8GLGAknK8dmwvg4kH1XyGWcfYQytMCPzRxFOb2hAiv
y04PDIoklk7tRvVdy50BlnjUolyC60iXU3OZaH+L3fGrvswD+pKEkEuD2IKGFoXzgTsqur7hkR9i
/1ymSaE1kv5vqaZBxARD+3lmt9tEU3GNyy4KK6ezqpvMADfDE+lA/mKnDN1LS0BJ1o/RV7dPd7cz
G8RqeILn5fYfYj+YMTioXnl6hmtrhpoVQEl+eKA0665GapAxTtVG4SWqPZQSWbODqeXKekf6vm/g
0AzAhRm6VW5csURpebt8ZY4FkRwMtMECM+CZIbkaEaXnF60MNoNOo+TIIAv7ANr7v+shpbh5qINE
zyv1an9cLZQ7w9VVlZa1r4Iki1EHMYFjwAeQwq3kdN9jPfo8NmrinEty84vi05Sq3HdVYUjw7r3+
Y9Aw423ZlLIqWlz5a/gJp1ZJs8zwhEaVpsm1VTkDWJoxqWVSEV+ayG2AGYvIQujqZkt+206R0wtI
7AzKNbUt6TJmu02JxV636wc0IvIX5QZeCxndnKJp3rpbDh4fIikaf8n+IbfB8rVy/N1WIjxhJKxK
4b0quVEwmwIXuHAheNiTSY3vvJsy4dLrs7ZO5KitaPRKun01yhsaP90mVbA/E6CuPjSjV35OptyL
yGJxtkPGiUdCmEUyuUryBIIadD9qz8y3eNmGA+S1D2V0DgimFSls5TZF2tVos1i03nDX/BLss0Ho
n3NkTQYLePeQO4hoWAvxm+lVUUWzN0EYdkbzqxMt11BxEaGdzh26o8+puzxj5ujuyPLpSeeN/toQ
JSapVaE7OlDGEx1z7gbCyWJwv9HHgLkOG3XMHFRRjEYRgHjzHWwE1LtRjcakvfVvKsAwN4n8/Q3X
w5s6yT9fWZP8keawNR6v/PG0h6k4fCUxcpjCLLzMytShD+/cIjUpvloKt9KgOJiarUzVtP2jpn+5
6eLxUITohxIp94mQhdqimFgzJmP5cCpoMgRxy+tOshcu3ySdmOmjZ3NnCet+cNlH2PhbQRWXFV81
jtRz5VgChZzeybxLDa7nOqTAfAVq/K2LjC9GfeS0ZZgI/zFslGDuST5s+jk+KETuD4HgfNkxXKNm
A43XFvafwrj1L11uZcEnGkAjuzJEYZF7gsIIth3dIVtObqoUd9yw2erY1WEzfpVm6jc28OGu5+u3
+VkNo5i9DNGmD74Zg45wJLs0aAaMvH+Z3L8bExwIBryMCFVXHoCXalxKrmCj/kVDEZS5I3C0leOu
xnyTj+n7kpibmIR6D0dA+kmc0by2rozS6beUhDsur0l1xomz0kKw8YXZUp/hmu+evNkynGH0/aMY
tYcKetSAcMUrfGu29kcoNtyU8R8W1mzQIXoHc1R+a88oxXRW51mwzLIkyyEJcKAR4elxXZQveyJN
thysHSXgb9WYO+5izY+RU/nUwNCgqkY3xuTN8zF5DdlcMR7dD73JNDQ2UtFxisE1IhYzPIO5bbC0
6VPd4tTbYNy9lku/IGncS5f0dpBiPYxtWXFKwNJ2xbqyQnHQLpPpGgDREk6Zxg6M+wKp+iWU0va7
dltYKMW9PCMlyUR14HvZyJFGqaZ+SUPxsAlKd1CvOcqPHrsXY1oNDU23LD7kyrhhsdGvaLZxj23P
F0YYdedpc0VyCWt8LLhIRg2/SIzKzM1exu3IzwZPLNAGMhPSnek/iPNUWUSHud2bEyBTMcqMVKNF
apQohny555YkUc+gK41qviMb/ZFEaGSVMdrz80nbl3kUSjotgq5wS7cTpYJxrNTrtrsNudarNEv/
gE360UqJhtu3QXdqxPIQ2TA0Zu7oOj7J6KeUwlzs7aRJMih91KTywgn83NQcCw+tcWiG7IDqEAur
j9w/o13xGDCnHKGCFokd/J+2tIlye9CI62H6XvLiNtEvyZuQIrumD3QibzAc8xMqWPuTgvRU8fBA
ZvSCgnt1CyFidSfNU+As34PkE2GiFQ9wwduusBR5+/AZqPFWqlloonl4Q0TgKopbmGoH7ue2qO6A
pip7U4PmHbH0l0twqTzuY/JELtReC4VVQvtHcgVGtHvnTFhtWLc90yVMNMBIxvOltteDY7mMwmQo
08OqufuMlWDrkh57FWvVGX2QxBbTYffRM30miAgjZYTDoVoG2JZTwf3SQXzq2C/6sfjvpkuVW5J0
yIosFO9vE2FmsYJfqxXJCcfr33ctwhmH0VmVc9YfZ1zEl5ir+y2KVrbobBBL0TgXf73DBD+yS8Wx
uTQ8wgzk5XB9dk44WkOpUeQte2z2ktXBD/XCl9It2w6LZbAOZ9+9WjSFSzAO1y24t6Es0LJT8lno
8ch8RnBPPMkQvoSFRH8gWOs7hauJ3juQTBFeVhLsuTh9HAM2tt4LaUTPXiXRR/QiWoqS6l2B/aHq
GcWOdB/so1gi29zGlvuPeA4kQJzcB8jERFUn4YHEm4tFHWfLZq3jj3cx0TaxfCckaLM4kO0YS71L
gHWobnL2CjfvS11lpY2e26qBcbt3ZijcTiwTEdZ9V3yu0H5eaSxSHVa4ARWrmspPWKIF7Ycs4wV3
UM4I2LmB0DB3VFbkWsVV/WwKneUvfEMuB+LGHWlywCw1mZriSCUEf0hi9yeksUlVbpB77f7Mc+4a
55XP9DzoEHZYlMqQgSwfVs4f8wZElKs6aBYRCTJyGz8rDjTCSaptgDilOnMf+jbVuXOl+QyfJOD7
jqjkxZmgasCjGPnD+0h0b17NFc6p5mlg7XJ3t5T78tIMM2qlPC0BtU50SESe8tmtgE9So6GpTgjS
7DwNdjU2Gq8m8Y45RcWMmEOHE16Ik/b5KGUFslYR52kLclCICaZwhxQygPLrEHEZl+qTW8dcg4R9
d9aRsxmMZoG0/LAPV922PTBGKJnMCtY0J0XVEfmlqw52pftJEZ/GdDBz0Yr8lFQJhVWaiXtmVjea
k+DaEb0lV+48ayJ0JWjtZ5OY07ZYIUIIoLLLsnyJsZiKRxk8NFGZdGuk5YDRy5b3xwFJKMxPATSv
bOvFdFyAHtr3j/R5UnK3KGbnWNeqmDMVMdhE2iKcgXL+lM150e8Gei1I+2e1crMNzsoRya+CYHnx
2nRwx5Rc4d3jSZ2RN+6/ErYcN30PI5a9JI259auwadQxFgVLmvdZlHBouhPDvVqkIeeJ+WSexI3v
XsuOINATfGcVbtlJ1Qc0CBmGq+jQMlcoaSR12aOopJir1SNRIhASdhFsbM3kUAoJgsUJPh/AtebZ
OFmTjrS6Ks/p/l11ZOsLiUDxmqH+Wwm3F7CFE241BDiOSI/ZAQeMTwMKanCtHKjg3ZWOA883jpW5
9LhuFnbZVeWAHh4tOtQE6kS+H5+3OpawryblN/5OIMZvDynt61KZjESGlSEBvDItldlvPMuCI1wX
iX8/duuthXVSSJw2huWQnnWxGWw2/zyZoMgJeWkR8vntwrFsfgXT7hukrJGYnC/uRFtwbvKWMhW6
dNIN398FCjSNWXktbEQO56SsVv3lmQEwbgj+VfVZXh09T19md/M1WmblBl1Oqzkh8Obp1q1J2XJ6
1jeJ1Xmmo31dLBSfxajpgCaXhR4McDri1SyP9TTLTaPcPmY9HAnJjred9M7Go8hpqFbpR3nYAFLD
tdS9CPPKzMTc7d8EEYTH3fP1oT+Y2cAhAiWbkseOT8K6zrZ+EeTAOtRIEHazoj8N9/VaxaIK6StX
FvvazNjAlGMMTvgXblQibqSWCZr+nPb6inhL9GqQHjJzDYBzyvs8lReoKx6FBYAUZ5XZaNC7d3c1
Q1pNumgC/U2c7O8G8Qyk5j0LwTs3/8QwXH6KzXqq5on/Y2+OlJwqDyeY+ZW516N0Fl/Kr/YIMW3O
07VgMdrE41aVlawObuQmnitBsPZonn+3z++X2Zy6oReGiMesIgCi8nRi7NOv4WiXQ+3lYVdzCk3y
veJmxkeKX1ltQZ+5TT29NZEMlJTZIW62OCu6ntPgg7OvNcGp0rPz3MtD5epO5zR8F1IV6UzzXOFX
Ln7j0PmRw3eMSO8aqfBDXBe33aH3uMlHb0TQ3GUUwac6CPJ0gk7t8qpugBylK0663txrKi+t/oto
mIesVdp2iaH6JdCJPORJ/QrJdGhAdaGLjovOunHIPi61MKGHC5GGG3J3uACxf/zoE45c9desWEbO
V4IcH/dCliqQtZ7MGZxwhQsCPTPj+W4RVSI/Rn/MCxxceG+G2dOhD7pJYNZwnloiQtT6QctSFeuU
Nl31kbRnOZzWp7NCa8f9GTfdwvSOgoHWR9MR495FrGQfZ5/sNeeXvvaOilNqHH7IdshdWxAiFL78
orelVLUUfqAaeDktFmuW4SbHvQD6Q9P05UyAhQeumvUn8ieQRVhRWNakF/HuONrycGNOxEhq8cWp
VV2z2lHCMsa/qrQKz+EUGxKXb2IwHsB6q4UckgqGdI2h7Ahj35yJPMaqYLL3OUKQ/PKUsl7PIY29
UgnAY7DEt9OLRK7XsYlb1F5EgFFyiIjg6hxejXIhKU6gJpml9YJ+1LXq8DjPycIciTx0V2YO0VLF
QYugWjLIvtxhgkk8f8z8S0Pilf4u9TqrOPpWa7r+CTqkC2LMUYBEH1U8IswmyGI8LhGECUaoxa+I
3L+KiAPfNM29XgLrKOBQfR79Qj/RTBhbgmSftlAdpGWgMwit8YSKQdQKQ9QvfHfNXjSvsJho0UAD
9etjptlArOj1NsYYH2shgxfuffTsjigwk9ZNd7KGmrExQlSGhBbLrPWn568LYE7lngIkRnpCiRrO
iO+8s6JPi2F51UzlBBhMMvIrj8BLzYSfZ3IVDuOoP+eCm//ijtpf1xhvFz/u7pkPAbtZvJCIdK5y
QBunpfn3k9TK67fGHOgrQ2LqeHXRX2pbxQmEFV7M7vKP5MpT+pxQeVuYQ5LMNwHgaDkQ6VVoGR/i
f7UWQEPfAR46B84W7XWStSTZqBrbrgAsBScPUz43aKEdgaY5zpiJAzT75msStopuoLRTz/03Xi5/
qr6rAnbCwc9VP6IkVBpZdoIo31/f7XObI7d2tN3vRnD1l1r+xT3XdkxEDMONsstnfqvcpeRLG5ml
b1MpygkS+cPFHjvYSaL8q6le51sSLlTROHZGgwlZr41IZ5XmEGdaNvsuiKpmdW5KeHpIL/Y7pfFY
+UD5YClSEfP3F4/hqtNmjKJll+H3bShCysd3oLqCnJHVoAVpfaJQ1x13cGPvy7aNcK2N5N22R0DX
PwICY3mn6eeZ1y3gnznLYm6IKEtCb044BU9geeowwrlee0neW2SYhdK7qJtjrjPWwsfTUtEBUlr8
qMTTdU12Q/Y1O5nZ+Dr7QgLYGfLqmsJHb80cMSbTICmj2EUGRTL/ZwOjtvsZyOwhgggBNZnbXwL6
i3oO39DnMG5vStleJb+lbXEEFUJ3QGwMDdJgO7RbmFUauWMlx9ZAzr54/nqwOivN+wQ1TKJVmc+3
oyeBq74oHgkr79Fiy/1+Z2rkB43MqWbT9Uaf/xznswI0lxwjxzTSmZL3LaMkke58VVJUnl6S6McV
bYnwMcj2s/vAOzZuZFf7Wvp1aOwHymSoBo6+hzteIvEUG2V4Ca7zGX78ZhcBVSJTv5RO7OCPZI0y
CKuN2WDINESkHfWOqUwz4ox0J8qdtiFJQ0spabTSeKVfWBsENANtlV3QnXC/ynk4TnOir3MU66an
TE5Ho0zk1MLOpQt/z8L48y+tM/W8BezqbFcdxZy2o36YSqhjE+eIa1zhoz3nYrz8cmES30ryJ7m4
fhyTRw5znlQ0jPXlZauxFFZkSixUTzOXEWYIt1rz4eE5ZzPlzFfy+sOWBg3luqnYJu7dJ8NJFyaT
aG7z3fB38DUVXeXjB+YAQr1U0nvN7XXXfIk3adspRl5pnO/mf6w7cFWKRP49ktq9AU3qAUo3wBdP
4C79LY98D4bO3Et0oKXe9pLbFBX1pY8UQlDfq34QlfaFQ3SHmsDaPpQ5Pip06kfDidmq38HkZ4k8
SxcGO/BUoT+ekzzB5zDPAMr9BQUAUzNY64WqdWEBI1BntZC8ldSeja9lq0mQMwnPkB+M/FjyhjnH
FGMEZFSgqR1BoApPMOVU/LTKfVS/cg1mnHqvagkSNSWlmo9S+LidqymZ+KQSMM8EHT61+X//g2qW
go03E3/mklc7dy1f6WFzfmNRYOIDZ8+eZPk9l/U86LUzYwak7jgmAOzKotl1cA3/BimrRiRnKNnW
ZQ+tskMbYpVx7S53PQPXm8gUFm2uqdjkG1FlosiMvKkFX4F7CD+B4svjhH9yNXXbjpybPSFrXbHN
3I22cSoElordwna9OUSmiYKn9Fgd9jDFuP6KglhB64KAAVyu8cME6FN9f9Dz2rWXZcihO6pJ2kbO
4Gf5LDGqrpqw6kqeucyhzu5lt9W11lF7wDscsv/Q6qTee37pSL16/eEOjoXiJsTKGuQHwhMu4mh3
lT2Bo+Wq0XkKcRfnDThUb0r3ftNwZPg7yV6wrGcRushs03RuB2ia6g0aDciBHjGjo+oOnlNM5Z59
eGAok9bO225wM14sF3Kw6xdji5JrPkZhPRTuzpRCJtI18cSdWaynat9i/aaTiAiEyrcf0U3JdTSd
nmkq5gXVT/9hdKAtT6q2tr73rltQcmXIvfSNPzQRSgcj4lnwRroNBiRdavCA9k7/bjj41kK8teGw
uWOegz95TZbTP4ll39a0QTO0CbAWdktake9lt5FOF0ETUymCzl2ZBOeMFsNvhCfEZxLZgkQP10vU
ViqfLmHmmyax2e7nId6c7Vm6dUTeuDmxHbY2/8LQccRjSBL2QUa1AW2bZjUcoUamQ8Trpjl5rb9R
n44eHXyoQAe3ZLeHcZtafQAvoXpDPD2/O7R6YIN+4AEt4HT9yxxrJlCtMJRbj1EPUVdnvCv5es+U
Li4kkOXV/8B4phBTLX5fFJQ/qZmAggVr2DrIhbDkeZmguIf6xe6/PcBKb5neoof15rOId8YNrN8C
Lsnsi1iVYbqcIkWKl/59D/eJoqxklp4up+SfcjrgEJX0s6A+tizMZqBe8ow1lUaHTJvEZoKeIEcK
luT9jc+5KfqZSz32RTaeZwyiPeNs46os509R8FopYxplvM5dAf3M6i1XMROIAj16fvhLqqzhNpTj
IRjLrLmTEJym2eI1gzN+GKmShGoeVcAbxz67KzabEY4Q9EF2GVu5CmYEFkaHPyx+QgCEme/5Er0y
PE/wfJKT9B8o1hGcir8ff1iM1if6rp2NkSb/PU+rjdZiJ3O2iztOuCfeuf53lCs92SFlzbhWwM1I
YcY/IMBt//cdpIaOS4ma6sNbkrLleqF1xr/lyiYdevekeJajC0flAL25fvzf9xhAv7njVmIgIPwo
eQ+8FMjF+q59WYBTJ+3OEtaUFzk9qN7carrOGC75ob6JqQDK9YgLYHTEyogWVdmArih/wtq7GPCK
mMH3YRpbxK0xUEqpMD7E3xuFkRpk5xTR0d6K+DJYJv9n5tLN7AtwqR3e+wjaYxrY3/wQqIpkE+0W
yROj6jBVhEzmByjfKiCAfNo+/YW4fLls8ZOLbTe5tma+R5XEbcwmezE862E8LgOqz1GzL6Q9rJvr
PRR9UbDJ9YLc1XkyDEXqBjhPp3NMXhOlvuD8Lv6SfSYAmzvZJvkwd60W0dZQVovywhQFQ7KBPX9b
dLgzE0MrLD47Noh6gvyZCFjUYXuZYS+XzZCotpZ2Cm2T06LZDJafBCZ7VpGIhFYgXGZZPJqIcFct
cGYYvUFtfq+lpypc90iqdZXhTthJOwIhi005Ugtv+232CFG962rUyF69fyLtQEWvBIaGNJ/C/U3L
U0NIfw29CctfLSwraqSbZo9CsNFnePrVvxm9e2Ls5wVZKLxK6fO/AKMUALpNnEJ8uTisgA+LdltM
0iiqiTtn1GH5D9QGjPl0k59VK4FmtsFnXO+3Eyttvc9dDsD3UvXZk4x882p6P5u+YbTgzAYfTx04
1OH/rc1LQvYA1G0lOhr8cXOJCgk5y/3+/m2dyCZenxV87wv46KzAybD5nBgbHuGzuH/MKwxcHEAo
lqHx1F8XEteS44r8ACpEft6H3qFKnMnLI2Ihjoc/qRC6a+mLNAUad45lopuIfOZVlycmO1qhwzvp
1u8I3NBkDWkjjOiPFFJwBpvNQPIQykX+D+Zbt9RdHGF0J0Gi2BwmidQozNyOPEs17m5j992hEu2q
LMHeQi/MSWtevD3RYAvSI7ZwE6c/9HvetPlJfgYZx8Sn9VJVuFqTMA8/tXz+90OXzlXg8CjiX4m+
qeCaHfTp2XNgR5vV87iVWdMkPL77SxVs1x+uRZWop+Jr1LrCrnlbp7E/meirlnSH+hoV3/UILzBS
Twd1h/R670nfavu2/3zaxxN5oLkUuFg5hOjhHVKjh0yh6hWgn8hzb/Vsmp9mp1ZHQi3O8DhYw/7B
OjeRqQYve2ToXSONBaezMyEKWq9JhnPi6fnfqdbrXzm1FjbGu3R1NJa2X635JRyBvTZTp7Kvz2sr
YWx/6NoofBS4bId2slpgcvkXU0g1JW9z6MljxuRFVwO9b9xHtf4/IYxuci8A8ZAJ4o4xoeF0j8Zr
7HpkRFC8EH87FxD/6RCXV3XE/fjgc5dK929r6DoSgrXIxTIKF/ec4qlTF0XjkFCTm7eLhQ+RvClr
SuSa9FnfgpKxu2y/NaLqOF1em1dUeQH4WL7UeDXCQqirln+FbxrhUKcov3qAvifraBkThBl7RHI0
Ac67RM/S2n09/Q8DTtI6sr9IJfoA08YPAdJSRc8Q4JgZwFzFKZMBw/8yupIjdHlG8OVJCgLfzx01
7yNGRMBE2kTZS1Ge0ekbxz558n7nz9PFs46t0Zfu9G6Wp1zcPIbdQK/YnzVWXuYG/nkLHH0pjFQl
EaHmc4VGno92pJmVcxPs0YeNiGShpRvmXE9uiwJugWe34MfvOv7IL8dBT61IsqE56YAngIv2ApMV
xJEAOR8suSkN3dy3cKDpuzGsyNDOXc0uSTo8xEJauuS26c3A9ymnvNFlFNcDWTLYOOsy6zgqNsxC
gScwfXdavq1kmKMXJqQ+p7/ecuYrRxnGZws7OIMSc2C9MDiJwaHfujgxnwhCeBFtLiz0cGWhif1Y
FW/4P/TjjKBjWfyY2PUo6og3Npc37lSKBLcqlektQ3HnsXOx43MnH96FNPD4/ljKz94FOQuZWNSa
uXBfVRY0ZiSORk6UcGp/xVSQNa3YaLEQxdy6NlZpH0rET4dzrGIijcQPdoITWI6MY38VH/VMnB3d
r3hSy6gsJElMx3I86gEdqkE7dp0x6GLQ3BH3exu2+dH9X1gPZ/4RjSc1/5XhI+I69ko0sXQOdzCi
HONGgVTlVe97IOJe1mY5K57lsRRfW7ziJ5lZozce+v6Ue+j+xbOst17A1DS6gW1MaSwJYWrflstV
qzkdPk6S5oD7JwH3xRgCUWfMFc2sTElCV/vhNFob5OMOIUpK+9GzlWJ1qZTzUgp1bw7l0KrBxkNK
Kx5ayIP4H8uilFSaGuADwQhb2C3WpNpoXQNo7ACU5E19PI90UeyRjath5PL9W7XESsBjheAOqSIx
wwSquyWbduE6TEy7DMuxmxIfk44R8PHYaaDp7+nsXYQxgtECijajoh7k+oWNNUcJDv9nba1FvjVK
2JYJWWzD+f72tkGAehTp0C87QIPKwJ1TUMZ+Z9o3Ln38sdNPgqejYRc9hYRVgzuZR1IwSOPeY03B
z5K8WAbwB3EpWajkOEFBuwHk7UWzbhUjgg1OmKpeNUw7YbhIy8T/aQAWmHJhDk8PM/XIZ9hlKuDA
dHiDQabIi/sGlvCnCIzdjQKDUif5u7T1rlkxivot4X63OVIJUAntfiPQoc4VNpodq5eJXvK3afAV
/yzxeBoEgQ5ZWrnCs6ileq605mUJcmLFZcAaZCUpBcKPFWlPWfh+QwZ/M+wFKQ17jWnziFbKUgpG
PijPWIu8oA4koLQDJ/lr60Er/5DPCwCjQqreqvZS5ZDn20yv4VIM5CXppsfOJ5WloyVHXPSSQjpI
zQAdN3yib3iseJiqX4+6Dh50O+oo+TWQACn0Fp+LXh1Nrwyw/4B+a4FjpIN9B0yEgCzgfHkeJl0u
4YrUij3v7z6bJHEO/2vkm0E+20EhauVNRQ7RMnVIAWAc3K5k9VkwlBzGuMNtZgfNEQm3pngx+57e
oQOEOSpOLuWxu9MkQ1rSyq3DS45mc9WE83svGNP5HMqfa98np0AOuv6vcIFKu045oosoQoydJslq
ZBPxQHW/X/PyNxNoC3uJXgP+UhYmHFdSrLUncvnF9wiHeu7RY8CbOK1ey5AMarOcYqzgt/mYDwmx
oRiAZm7GzwAz67Fu4sZdx+U9wzC5ouFHWkGX8+r71ewOZF02V04qxMG2p3DGRUAxq0xlQnJsn85x
6R5DxNTXkvVV6kIJdPJwIoDmFYs+nJhk4afBHbxbX+ICs8oYa96lzDkk9v3ht6w8Ijbi7+bEsG/V
pVBtSknQ0f43r6KUkH/0VFMJQW+ZHp3YOUzGThshy6k/QCJiP8DcLwJ1opD6DcURrrwwhmO2z7hq
blMTL766dfuvsYbyvtABBlhdU6jbO3jtRPFqTfO3iqn8/9XdiTFbfX+lDWyIcM5OYPMBkwIHV1va
PelvodKxD70ZSo+Fy8oPsqdfriJtn5J6E6XFSmYbrjFSigAklxUFSx5+5N7DR4M0WlnQktlhO8d/
5Y6CtEfgJLWa6+9CjJsASqI6VVCV6e/94Bo3XrkePh8puazhrKwdK/5kjH6GcTFpzGuwb1LcrMWW
fsS0l14dnoFfRrE2hkrKVENbahFy9krWWgC842s+3ToGrSbFMaQQWl4ajzl8B0gpuVHeByhuUP8P
mVUhYc6KFbjjn7KADeqDrloTMXewRb8EN88+BefVVulGmnybN4KRgvUcI8wIJ43eA46IuuHIZToP
pFvr/J/tPdCUWOmHTBk5aDppN7CNSsTXESPIrcH0T55C7a4QvN1HeE37ZXIP/IFgj+CPbeGwsCQu
kYZPdv5ZPCpM0U/le+lBz7517M+B6J5bcmk/StlC2DnUjTPZB6tkUKrB0n0KRZ1vrYd1NFP0w50B
4mfE3/c=
`protect end_protected
