`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5088)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbkV3TO4Ee1mp364NJ3ApJ1FbWY3IB
02vUs3YLSDgyj9eZXMh4yaqzcKbXOgmmjbKlHV7VT/2nPr/n176PYqHpH5WOQgLDKVcRyUPmFCqo
Vp5sbvSZ4QuceQ/e7X+XUNUhZ3OzLPWnDOniYwtTagc1ZwJD8OccWAo3ob42xNhq100XFAgav2Ka
svIGe+t+WsRZO6eL54E2sqqxIySewOzEWm4PIe6ICW+nLDZcICddalIcZYbYiIdS0JehmWwv0UkN
pcwtSRq+STrfBz+r5SXKYg04zc/jFKH+OW5ygtJTcL8OId1LA0QdeAXzErkGkr9IOv6Bw5jNMoGK
JlA+ymZaWWvovxinBl/9jQgvA66eg65RGHI9LRwviz5JkSXnKONyzUrcjyIBfCLJphHKm5JQTbI4
tcMGEhbZrc47kOjgRSJQP5BgF5kqX8PKp9UsHSRK4zoyuX/ub2GWl1JvwYgM41vqPrC/jpRTNCeR
+VcjSwiGjfJNAVhMIW9M4adVOtE932xqVomPCxaUt03fKA6uy1bcq7+uebImZJqYqBXxbILB79vr
A8NTZ6My9U0S28Jxxc6oAr4p33fkYtHft7paTiF/WX2T/FbK9HfDLBwDUlP18RVl+yGJNKoxKnnk
50FTVUHi9NgJ996f91ChAGuTYYpedF57/vO5Ve18JhGO4SgKOGm8sZ58cC691M3gzRwtyLcm6LDt
cgBdkMAASA5KBlqf0/BD/Ubeu4WAvvpuumivbHKqvIk5EArwEro/MaBnqrYedl9q3rW96TSyvR37
0nWJ+RlE8YeliG6I1nXLjPnJS4D1xsyYcCwMMyKMyLBb8eb/K/7zuVrqN0ziJ6AZpL98QboSofZf
EH/S78v7qJtHsxEIHynntBcikZ8dKTgjTysIYPBXwl5ro/8QXz0MQakhvtImgMAbWP1GLOYcJr6c
RCVjBnq/ymDX5kvEhPURNYNVvD1vCIIrL4Vj1Z6OzAkeQU6Vmo2dzmwBj/yeoRTprpCRYkAY/olc
p+t2ZlltQ51vvEWljGotHOEP230S91qd/BB+myTN+W4B1z1HVIM8a7isQpcTdRuIw/jFyQbhr1sb
oM41Fw8f5rgDs6F+WcKH6lT/ggpBJNA8Qx6JV5K3QEziOKPd31Y5zHjV/IMKonwFBXgNDiJnqd65
c9wD7WH9U453RZBdMX8AbrE8tnyLXc9Srx8oO/hRoeQHQLTU7XGtX4nInbLBWXnM6peuhJWb+oXH
Ud9XhJg7nnYKnCfURgq80/gvDIJAdYFCWKjEjoWSJHZ6HdCcZesAfWsH3+IdxZlNsCOB6BbWMrHw
AKeXtvowhbLEVl3UhL5Ozq5E7HzberxAMZwaU7wTDY9I5NZUk9RiyZFNO6Ofi0rA3y9nzoRbd7OP
7Q5+31gbK5vO5yxAm4OIdtqhfS87PG+8iZ95VNQlAZA7ZtdR+JUzajpDVcjDRqnyNfr3QIX/99gE
aOvaTe2PdOHZHidzCv3NdUnhkiYHhTsO3wKLsRGxvnuDAJXB4W9f9BonCz4YahaHuTIbwHtL9Qao
5NfdO+/XFxbsXU5EsqYtNgQrEl+B1apwyzkocjOy5cg4NoV7XdMwW73N0sJ0+obLK2gV/HEkO5WP
zQoBzPkxE7RC/URVTVsgIOAZs192tm5BoFmimQ6z8BSGdMxhrvH+5DADKD6fBJRXvgDKA0GBs3Eb
ObKsjKpGRRrF9YUUJAdEjVJFR9w/2FtibwSyfRmoGkFf+w84Yy7ylRI9NrllY2Uzi+8XZs2c8AGr
Da/hDn6yk+2B2LyvUQWZydDSv4nyMZtW3sGiSaa8zwY0x6nz2wG1TIPRX9MTJAVnZksbG/UEJSVI
Mvjax78JUjrH61YZ7sWXfyxdvSTJi0wPl3dEZfw3PN2TJqppsM5YJ3PGj6uOu4K3gvPk+8RREiuW
4Q3+Tq0nYBnjv0V+b1gFYpzaf+jGJROKeMXOYsWruoE+B63wlrEQ1znjPDU6vXg0PxtsnFslsJTc
C1Xc2IF0LEguRHi1Ed7LWy9RQeip1uZfaZ1x3K+SmCew22KmJEbOcIEX4nJrMlQBHMhGN5gO/3TH
D6/dFz/pMGwjTB+tqO7mrjP+ADK+924N+gjjuE8amg44k4O+LwVyPd5SzWoUUIS0trjsw2ERN3x1
/AMkQHusQdx0bbSL8eNnDEapymwi/dsFXzfK1QWFuqcZAxfqOx7k4HIfp1foQUHHwq5g/eIEdLVv
WRNbOohpn1d0y9wFjiokDI+n/550KPdiw38cx227w20l3Ud8g5iG9PJzlgpsmI5VHaLNQf/hLQG+
kVeN3JVz73YRaEQKsXPyK+SuQNPIDkzXVhs7HcAFi0xoW7snnA19WHGWihTcYCu8zlB77PJAi1rn
o02JE5qXvByHJ69PhDJHKOkmhbbDpgxOJCXAQpIHkFnu/0mpTkV+5xYrfTbQmZHgtsM3Nm3U0EsA
Qj3NbH9m5/gLmQVZswwcc5B+816CrK05KnXozH2olnKw2y97XZ+TBGcLm2DI7SoXCz2O/wwHh0Qw
EOBf6gy/leFjRDPvGzMbaBs8sGUD4cRynNyxMv1aQA7uABCAE6ooqYt+o1iqlGdwXKKsuy6ycByX
1/0jFZQpbtCQ7PQiy9H2zGbvDRWhw4yWL1jJ60v9DuKMIaelUoN0iKwfFdNZ7dTnxNrHjcw9Ufe3
JhOOsWD7nfXhvaWZteWRlkj7mAScorH/lHdOGvEZggcO3/IfPglA4+6VoBVSvHjzUAbqCVxT8Duu
KMjJKEYyuXRkh0sRDU5bYc568DchnbaB5HyZGcGlPclB2wV5bCHS+qCENMMRkRmJWXoEIaljiX4l
cU0qC3A7tcQRsKmpTX3c4VJap8oEv5q+my+zRvpAAcYjd5uEHy/7kMO/ii0MGa851hNMoDlF6xif
4N5PvSjrbuFhhDGttnLviPkPOKQh6ghfi6J9dMP1O3Ka5ClflVy/9FDhqN+0o0CWwxnHS6fC8lLW
aLrlmlJh7PlB/wW2nNJwYTd1Zy2WXrCLAFfnJQ/YkF6hlh3lmyYym2P3KzH95IkAOZR6w19Npd4L
8km8Ug1H6XsVtM8rIGGAV+ECZ8FHWyakFeYpGb5WS7o/kTUnn3THF5ynIJaia2yvrPCWIwlc1dXF
BDL1tGaw9EIEtGqw/a+m11s2POp+Fq+pU8eF6zXmtvDrKuurrqVqjVgpzKHolq0j8RHu2GbJUjFY
NHmrVqH0DVsO7Nk0kggb49Tj2AtAKxFZELKNVte6UqmQAxMYlffFyvNP/sHUppuxE/G1P9+aZxMU
FRsiXJgE9pKdtAZQ6yeAXndeTeB230IVVNXeRPggLCBckif2HzHAoUaArzj7MAAZdnyU9Ss6bT/I
CcuwBpISZkvfQAz37Kao
`protect end_protected
