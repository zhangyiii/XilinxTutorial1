`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25312)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAGqLwGYSI6uQ7AcSmnVV1T90WbP+Rd9YkulszJCNk5h6N3Q+wasJ2wC2
1lmqeBg0TEsgeiT5YVHod3tn/tFU7Z5lcIQBZUQjUri8anpblsGL+E6bMlQrZOpN297EIj9quRki
yr7/Js+3eICJ0jK7cr5bZfxJBT2ggdWMG3TUyG655N9iw1adiND5L/2lYLAoHm/hASY9LOvSvjHf
uNkNze71ZDJ7WAXaxCLMBaJ1N0d7EdoGiPfE6q07IoNPk7ZFmLBbwHvBW2OKLNkqldtKqt4rUcMa
EQC30pGZXGDQTU44iVHPjrqkPT5t1KUEgBAA2puzf332dzLJc22E7R3pCdMdcxm8g2sJnbBn2OEK
bA4iT8UNWWfuGynrCuSIjK3VhIh+XPxrrAOzs4bitUBEemWOtvB8lh+NmDKttRlNmO8FqqFwR0/5
/LtieS7ToCcwLHWJGyJ6YVNXmd+NrUPuwWPMQc/778vQCBpXQ3QCVXkUE9A4FFd9vrlxvUz/BuIM
QZWZXPZdBvJWFkXozhNXrHWScSmn1rO0pRa8ydRH8ZPw05vhyBF8w1AqGFO1mZ3HO4cBIwdBuUHe
EGBbTQNQOWiEZXMedv50uM3g91dbRIY1jg6Sba2JpLDhEcVsQkX83GGDbiYzoQ6dPPpyeJIKxK2Q
6DIBleMyLjyRxWTdpxylcU97ycgDtpkQZIUPGPbR+aKJfSZql5YoiQ0E/MG0rbwG8YC7jYoSjYZN
NzIjSHimPxSB9as3mBnnuPZZUD14mgATWVEqRWpzmS4PecKGoSo2BxfrTlinPM/6EzBPIjqupn6J
NrrxzWElh/PCdb/XRtOZkNwyvqYa7yJ6fsyneg9ctxH3v8vVvUeA1xnCPJHzJMw9bxtKVEGb6PJY
DUp3xyN4lNAPwtZ0z9Domye8UH7S4qkROWiyR+ANBE9+Yb56HRODwpk6Fb61erYKVE1CLdM9+kO+
KVJ0zA8PJbmh3u303tgtN+YfPKpLEdVsKYE4D2MUTJRF18g1ulVmd4ok5tpSFNkheqXhXJUd535y
9dMQtLgIepS9M2wi9CxowBjr8pGRUQQ3ZBrB2v1LHhyaSui8FA+F0LRmo9CBSF8pos8RgpZGWhf0
NG+WP1kg3wuc7TJnPjL6kOQ2XJFMdicj7w5NbqUa11RCc6tj0x0HRuEX6Ihfg7nrrEYXvB4LcXXq
qg6t51edA71qqIDjwjQNakQJRPCsl8Cn6TZnS8Aob4gSJkOPCucyIhiw599Qoksf3k1m5Je49RRQ
COtb7lVE9VYBKS8yktP1F5n7N30HgjA8XXxNYXzszwQpHPmS6ur1jo8l1zjqmPItBLvzYtUFiJaX
ykN+FOOTKUF++ENRwryl7SZVHV0l54haQzmgytGBlu4SxVmf/EgspEp9aUqXVKq1JtADC0Kzw1yf
GQ2RtcmsJX5rK5VQw9nzTdi9m1x3/Y7fBXbhPqaB/ot121AFyAuKKg69xHc42m/nhxofZ2RaoK/f
i28g+Ppl/GnAceHX6zxPWwOTWI0dEznH3Uj2n32ckVLTfMf8UzfrYv0OIdYAnK5UYvl/2sJ0DQqr
ZhJyBkY6C1fFq5ODFHLjvwlgo1QZ1rjGiTddhI9ydun02JLSr2Ep6V7zD4YZeTRonRzk+WZx4ZAL
n5gRpxUpjrfLLOGNn4Z9eAs4HcmGbc9adLdyjN1Ts1uV0L39ErzdB7EOTbKcGYvR8nUtzB9HnWJu
lHlE6VGT4rckjIKEkwCy/SLgdETPc4QyUysTqw6yXuX8CiWfv9gnkXIZqa6BGAHex8oK0LggsRwl
YMHN+wU2n/vNKrK+dw7bbcRysYTrSkb2+BMWfrKk3H25LhCeIIv+5ebbEiSO7SHpzVqyzQm/c52b
lbWCtlp1TnqRc4IZK7tdMV0SinW1xEl6M5nwe8+ROwBViu8HLfeItxeCeQ72fm9Aup8KUTheqmf+
9aXqAEbKACXZHjYbBAiAlqThpYjAxNAkWKqeXb4nyMOpE6N9jMmvOOOHd08CGGLHcvHZyxqjwRp2
chiBX+FJ7qn/ifmdQk8j9OmB41L4X7daQqBNW1OIdXbSS1LGLzeOOeTN8SC8UednspRRgzEyh2u+
KLGJs9gjbxHwLd/N8w31vPMkJ3v1lWpnnHNLCOAOCEqzJ6U4LL83L1KFV2v2prn0L9xULRhYKKHN
zBJ7L1AWwgdCM9HiICcxaLsEBiWdxTVJPXkXHBcY3utD/NV5DspnRgBBj6xXsSG5WP8Ygn1SW1jO
WlePOQBd5cLZB+oN7OdTV9S1clnA1fuPWCR59pwl47PQaDrXAhHcie1SIPf8A8XJjcVOROg9gaJX
vF94MATQ/eZg9nHXUax4efn0i923F6FtXxi/RBTTItJWRg5S+SZmIaDwRcxl82uSXFE0/kqaUXhr
n7PI+3R4UKKMw1fMPT+WMmxjb6m5eg9kpm4QcJqIqn5ouSWto5grRHV/3heCsxsRLkLRuwfRpeVu
zfNcqSRoxz6OMf3M14kgok/vZ34WGo6iBAqxiHU15xrfY4URd0GEBWbC1kq+gHqEt6R2L+i4AucS
rFbAbqk7BxuvDhwl5uzw71jISws1WqbDpDIfeDnKxZWnvr4IOZ1rdmeAadyZxypGBeuEFHDGyz6O
V2S2L0GpG+qxIEMLslWvoCuX7eywNDM81m8M54V/RfR8WUUYfRPWyOzIWeik+BPRq3+4vIVF6uIK
M/JKQktDQUh/20XI8Jdtrv9CPN8VUVYGsJymnPEbmOSiML7mT88oZgiUMxVRKP9PlqyJQ7RaqXkt
/sBmd/hJzqT6bqX1qOYsmxcV7a5yufVWXk7yycSuJqI0KyqtSucOPYSPb/CMi/rIPMuURAdcxjTA
JlWs4A7D5zqkaGtWos3KvuAu8Kscf+GiehZ701AUtFnKhItHqPONWuSoFe106IoTiujEnMQTd57t
29ouWPzOX9lCeDgdsFp+Up+wV2p29laKRPiko3eevf+8HoetNivI6qPe2XdI/I7tu6v9+C3OSA9h
IWHo4HpPs3XVQwIzFShcNMLp59V+hKYIhH8W8EsK9/HltWgLRpOCP4Vu+ENj+RvHdXOyDsT4mccj
WD76L8tc/SNgGasGtmjPJQlNY96BaOutQsoGgiuZkyNak2mOlsrU77+pswUNdU1HOiUl2/iaHCUs
JT1Z2MuAc3ypisj2+2z01Q9SuokULcdRx0huU+GyVmvKYW8e7adsSKtziG8Iw72hOD4mYtViuF5C
JF9Z5wYIrGk/lMoHsu3BcPhti9VEwHWx0sbxCK8nbWepYpQr2wRulR/0pitCaXDHoN5i/eYthXIy
ga4EV0Fhwy24oSkE6d8OUoPCSjDwZm5fYpaX0xhJu6jsjpdYInpJyBrpsAGhxEe56UC2HbmxTij9
+YgXhXIPLDezMPL9nNgmvM24wO6PbdbAyqaI4k1r6KHpKqkF8dEDRFOxXrmHJpFJd0G7YAjXmYts
VjtzcMlt4iLBewysnfZYETc3mNipnjAV4bkqVITARPPXHgRWYNuI0fvmSSbz9ti/RwUT+lGCxGlC
2fz0Q7aU5e9brSKEdoDE+vyFBXlhmVKGJnkuxIiLDP+gk2c4avgtW+hI03SKo1uLOwnlFG+yqoL1
0nZ168MV/lrFxq3VMn5oFWDE8GaHNnyfE2KiAi06WloO49i9oL4CGbAzH5+WXDk1Z0hhoYjpIhXR
5QibHHlgAHUAEaWZkLXOcaTMwGaUlw5LcSxDM2Udbj/3AIuQQu9LHR42x2+mwJfKRbellqZ2xp+P
Joho2OULvd7QUSjzpHfws6oGGk7dgjsqCIL45uPtoSsEH7IxOUxzxcjPv7/aaoYU/BTsZkg27lfG
5dx/20pwQv/RleENn5GTn//HPxlKDQDIzlUOtSki5lA6mGGaFiDaUmrEFRGfTChTd2pcQ8IGYD23
DYtQXI9xiZyXejeY3vmi2d1hbU/irDx00hGKKtjj2yGfPwV75Yy9Ftuw5nr6dmZ2Z3sM3QuhOd1u
vbC7lJDhMRdeIhHcdS1ATO24dcJSykPwf1AxzxmrQeLf2HPXjl/KLmE5dKX7hyW/UZvjFKYvTuwD
76+nmwvNCTK80BKYnufkBMIsNkuwB9Hrv1ulJt1S83pzTTGd61FubmzjCROQ4dcDl8wB1TWjixR/
1JpZ7XZg9MJlJMsy/vdzxVggsLutFPaBCKlGIyYEDxJWfjGo3KN5yU6Ab3DA+f/Fw7gCAQN0WN3K
9qAJEzzaP/lLMguaWh5vqGyU9y1IWz82SnWIeVM2ZTl9aYvilgwY/wsifTBrOVO312x1mwk8Ouk/
PL6d5hwZs6Oa8rc0qsY+0mY3Yp1CbiY7pI/Dn9z8lxSAsfQiG67mrmM/LvSy49b/MqU6ah2m/K88
D6IR112WJJX5QnE+y5zv7VlTofOJoOSv0tbUJpv21Or9cGyesAHgFrc0vX1ou3WCngE/7mv3F9cK
J0kFHh+wZKXBTF4FPjkN3OalsLK95SQlNeAP/BYCnrXr0gnqUjAB80KL3tk+S/vj0B8UZ7APBUJq
ixD7CpYbbGuQEO4pVXG6xlYmJFEvQv98IPmEs6WPYlEDfFbyJ/YS6dXSoUlOABrv0Zfm6HwQICk4
5wBVDIwBezdPYnF0Ju2njQShf+jR8LmaPZVYafXYQIHzMoubfOGJDRC/I/UEKrmlKq07llR0nQAU
Id+80wgsIyIpIoyRh0Hskf7qoLu2bpDfw0Wu5xC4eE3PLica6DowESQ8yeOs0vTJowVMeyDO8dWK
lKj0a7zcbvcQhYHUXYxu0Rfmj3DHoakQRWi90v35J1qmTtRpT5DTUSEBY7aI4K+RmBZY0E6Z/VYq
VeIGSOo678ZnqlDL22Za1wryfcTLqkDK+1D2z8tDCeZ3KOB9cXLKSYUwtjnvyApOIACNkBw64SEU
jMefIiNlNyudy/wk0SGMvkmP1BKGjDfOQG7hBqULyygloSDHVPFkGBRaYZq1Z/zOvaQPfjgYg4a6
s99PBbBSMWMnDHk0QJa7UG84Y1i20aSMJNq16OFzQubRjpcGea21MUsWcNTFRh5YTrxKuPqQ6cxF
xY5NRblqTN7J9IPZyZOMXbwHnRlxP/UKZ9Yuc1+OW9w4f+h5wPob7yNnt7sdB6M27S8oGMD72Hv7
Xh96jtCw/EzNnTpmLhbFsdSLX+XLxrIryvJxQUeVjCTBWw631Wf4o+KhVUM6sR3CJS0n8sEv5OYf
r1zslHtErJ7EXrmO/7y90OCICkD0F9WY8lKkSWEd5yXDwDqvzevoUmOIZNINefTDKpmA0J4uFQIV
M2B/mlklnRMlNyIE6JIGT7R4oVZ4fCLj8en6j4QLMuQWfYM8IS1MhBXzOdykE3inowyCAr7WSjw0
86Ixl6dB21ELnjuBQJPahlbqswEjgb7OKn/bZMQL1TU/6k/UjX/x8GOnOxqKb80zKKybGajfTOGL
brfptW/NpyotyR0nKxelAs5y03XiwksZizKmuM7IJfb72nNlw/6NRdl1+6hJOS8t+b8EtyhCrzrc
cwOlJly9aZ6bgHgUGKZu/l5qE7BRapk1N2dvQGEuKsUHUwlRs7RRCed3+gEnTNp/rrqhN9Cn0c2n
zGin47mwjolYlgoUfYjc6gEaMrWRRwDHRUYEsrCBWaylXRYasUYgQ2LuNQ8xMxusIak61rT7NOzr
iqHUvW+q/xm3Ikymj42xftoesz+koX7Bi4mP4PejxxP4NVdDCtxGfN5rQUytd8jBEx7uYd4SgzwE
+9ME1WW7hfRw0XP7hw5O3eM+20Bk3J7Q+a7hIiQPBMMYNtbomckD8C/l1sfDx/eRR5e9ZtKweSE/
ECc6PRAYCHEUGSgdM+w0iVh2ADTfmuWLAQuFw3rZpqyX+2E2eYmrEEXBLmg3MXtSWyfec0huDrjy
rBP9bxGVQBSRqUBwx2rgTvcMDTTkHCP4DHvcn4/utCNxwcj1e+iEzCCxhAqRSLyvsm8iHUFfxpBy
Nm/HTOvONkupkHM8WTBVomeZOkPe6xTxU3j8y51chNcqvJ6D/uZWNBuMUz6K+aFyniBUvyP/HiYi
x89QczgjzyHLe5Ot8gg/Pk6YXuiA96vZRgISFEcL2Et8Uze+FSw6Ijdi9qh69a7tXcRy9lmS0mLd
XkLlxbWqv6pV/diMNFlbpliQxDxEm5zdRC9FFyO8bKJ79oTqCmr/JcBhYxAMPRV43x7HyaayqM9J
daZMwflRiLtoDigLgcRPZWELefVxXgCCHYS3NlyBQ0Xd4xgAP0y+P9uE3G3fLsldZ3ADA9hEL9q4
6jbJdABW8/jhXPDrXd8u6ZbPWzPHGJpvZpmFOwja/95J2scu/nt+RI3r/xtjZzQx4AaC1WcT2ZPI
/1qb6V56tDjk+SP3CzU8vzyTcyfHUn5ZifXmDO67Nc3Fvdkw2wqs0h2pV/ll6dQnt2ORZanU6pDJ
m46iaBPdlNINPSZoZ5RlPIiGQ0Fd1oVwbyGPdV0/6pSQl/w5w6vOaZH8eTEC7bguLY0zQtyewyVo
Hr8J4l7AT7mx6iAE6oWh16XXBNb01nNZMRkK1FFQo0BPr6sdrpZZfW2PLXm7K+XneFNM5bXp33mk
S+mEDELCRpBxzL5+RsKbRUD8f9rGz1g7WqSAgEtMz7elJOPHchPcbAUNdiAFGDDqgXOeTWjBsaj9
2FIPcbTDrBG+ahQO0YKIXnwGnGYkYe3lxK6prrDpg6GugCsGeNBmibzdvvX+t/Ds2bLQ0JCxTVYZ
3Jpa9AT3oOiIfAUxP3KPEWo340Hsx6d4H7sob/VoBQxTLDF62ovdMswXXrEq27s+JshXoOuvWyxw
bQGCRjDbBHGftrPDoup8NHv7ajDTWVTzGZmqHNCyEeCgsAvNQEvSKC64pYUZifSvReTYWJCKe7z+
XWsPLKBinPos3k6Qie1sIW+HPTgH7+OqyulXjUS3TEy+jSuqzAbL7J08L6rU7rf3kQg4HC9zU4yU
Sha9ZoFBOj7Vua7sHIJsKlv1MqjZ39fFY1xxDQZU9elwMxuH7PEt+CmKmFhWwPvVQHTZf2oA/XPh
yjke+g9G1t33fOiiF2ty4eXvOVfMKyf5DdB1UBEDop5mnIdTL7n9A7kuVEzsM4hZuUidZXM/kCRk
g7ATaGVL3RIDNvom/ssbaErLFvjvH4+Gpc5GdsbwqrCWQYKgJwOh7LdM+FR1sgLJ8XPFPE4Vpifx
MQoq/s/OdO5EGK82/FoiYfXty4i8FFrx/BrhQCjr5nuMsPQc+II1iL4SRrE8hYiFuPyfGx240QwS
UY/nIZTTqHqPSBp9ExT/LTGwrr0DXKXToOIXZ4UwdrzTQdCS3m4hduopdETCWu/6nSN6QFBkCB+z
XFYNsbLs0l+TnQk4ukhoPq5BuqRfbfdzAJFn2/8ExLgTZhSmy7xQdGdbjfTf/8w1u95LFjDgPWur
vh/n/YT5iiM9zktIqz6Ucz0RUCoa0D7miYzc8Zvvs7MJZuWk5YJlyhRkrgEv/DFpcfW9yN+OtG/V
TaL+nH830impFCGgPLvFSMF8nS5riUAWGvJLIR69NkdEx1sfzud9hZ9hCMpgfjjXfCaR9lOpzjO1
vaw31q2ciNMgYSqsiKchApCcY6yTUiPJjbQhU9vEStHFLxA2QdA6wEeJVw6VJtIAVOOXMWSuWQmr
ayz1us20BbL04Dv4Lg9Qa1E8JGC17eHXJtWDC1mlnZkdoBgb7lFmkxTLRN6FzjO6iwm0APv+Pjph
Yi+YicPVg+qrcz2H4yCYt9cbFRVLA/muTjw9SN/aUgCJX3Voq6UvdnCMnQiaHByXiwcSZRl8fMuj
OURV5q+auigjOg8GxQqlioxNHlnBTiXB4yp0OxU3YgvWa0VtPI22DnKxuYiA3v9t3UAmXLCmDY96
dLRApdRd9MrGDUqstyhwZD9cUG5mgwqRlyoTCE8q6WDIB0KG0yZu3cKVQF9G4nr0zVdY1PW1ryxM
aGomvpkwgsQg458IChSNmJvbme8+8uOxRa/rAxLDcfKr0xFHoRt1EsTLNDEmX32oMEWdnDJZM7sB
rjn/paKcBpSvKZIuWroT40ipbOZ9Pl5ZVh4eqdl4AgjL3wLuaG8e+WLMUmPzrQD1Ti1Sm/m1A/ME
PZ7IygU1JoLAlJddqfgf16cGwaVEW97GzrKuvxey/+8pXi7FwqL9t7DM6Xf5nvXfknhTaxK4WXVa
GyrC+ukmyxKBlzwIB0/+tR8Z1I3YMUUPEAg3siPe+xpy90rYcAxccVM4vKvrL++7oIyXYKYhPpIL
980fYl8szbvBttGJvRBt05FEyGdQp5R9NadNiwPUFlTcm33X8zxwEYMIannRyZdMkCzrEmU6/Jgu
tEAo5v1HmcZ7eOi+ad4M/u8YgJ+LZQdDaQut33bksqNZzu1lgjI7vBv2yWYDIfSWBAQDPU0mmnn2
R2LUbA+PJE3jREwWOZy8yfZ5pamBIVTpfgXNWcnDewI+RqdflDjDb5ltBSvGpZkHMs4B8SV4AqUE
MjTl3YD7BBen9TdREdK2yON2OFJSTrUO7jnAYnCwHKaM44JCrGdgVm2PVXBBc3kwZDw4NS4MZLvD
lkz3kZaqOiOyp46A7sbf7ib6ZylEFyIw2MiSXFVlTqO/lawZu1Zx86bNGc4rlr4LJdaIxIAjJAQq
2Z3AS4czIdYkG7UnGHHqHC9PBwUYX8nbxHfe/xMemyXKpjC+oDtbtDv3/d8fC+oiCe+4N7TiWPXh
qVUNpRR/EgYwCoVE6985Z7OefZaulTDiaYfeu7Hm6rpjZNATWxvng+4rXjffDQplxhOjHJOWozAq
B8NqAqIHj3scX3DLqwK6f0pZ0zc1dR5W7+731kiHM9DAtvnzbbKB9a6YeMPi5/SWHby2cPGrgl6x
+PiPNJ0DfLSuqPgbW6OxCFCmpPN+Ep5JCR3K251fOnC8qVlrgfZLVFqZc6EYV4Vfl/kAtuWp1OQ3
Syz2/oGrSpD1WJuvDwkjopW20uJeIQf5SNefVWs2BEoXDoXMCxRh8w5CAEAraO9kpX5m/KZcJX1b
pTJat9wA+h6wGGtFjQoYUl0ljTuEDkk6gz1YG4RvWfqBCehJBsS1Jvs0BOGx4+Xx1tXwvNzi3a1V
jPr8OhZ4L9dZA16zeBtmUpG25IV5RZkO2SvIIisvCnddk6qPzPdA+5uFV0MMOyFguWuqBxOVdCP9
gHLPOLTRhRQ2U/nHvIkvvUzev6HzTrU0HRFvcsjDlyAMegJIiC/K8r13LvFoXDoQw1Nclpqa7AiV
UmN19Fm3Ng22Mc2990IRPPFQXbIcloBkqUSeU3tcdpRHQEVuS1SotZDy6aPyvkSZM8F7SMhF6vVM
FODP/ly+YGBn9f6lHW7L2dnrjM5Gs5Lu6XvsgRi4StCaCGSYg951yiT8pFMwFryZ70KynOG5Wnf6
DvQ0kT0Z4jo7SNSu9U738s5nJfcvB7WooX9RnjoD80XC9SQWIn1BOeIH4D8lAU0z0RINNVZOmGmr
+sYAX/1iLnYOS0t3M18y8/MXvcKOqNiPwd3fgmJuWSzqLTHyRn5qK33G+KxPe+weKOpFFEMPzeLC
GJNn0vIsdsuAKkqQIGexhcAlLuV4UWnwHqPIOkg5wartKtjAqYHKf5ASZoeM9V+LoHkSEZFzfiAr
4v66oxkp5Fnqs9Tj9WeOote8JhJ3Otl4INMGy3oWLUY2kFAkWoskI7HuVnz0Ol6cvfg8wfEkAa7R
cTnAb8yqjTchmK+YLox1JumyfZZL77s+uE9n4A5NJpypbekcj4I5HRk4PpzQ5P2aAUXw3xBW7eRM
zLr9+jlBs/svkB6heyLSJ1/wbNVcZQctJr2R4fZSfkJFYdM6t1g1RvZEOZ7wNuVp+upAM8UWXl6q
j3opbQ85n/yBFxF1c8Ndr7yWE75kS2R0njD8k4xnNj9v+kvGUYN04S8Te+AmiUwC6xsCYRP9oIZQ
4aADOj2ZBDomezW0o99oWltmYHbOtdmEfBBEatjVrwEGrCgCW1nE90Mu+eue59VNJXBYBCYq7qto
T2tpTaa/0Q9Ma8VfaTnSZgZ/sBm+Vpxu1NJI8he54AmDEyt2cAGjIzLXOMvK71HDXVCncvPbkKI7
NquIJZcxM/UxVHEmwMOHKHH2TlDHGyLtyFnOIXZFvlZ9x2O8pcLWy2+omYGMC2IXA6pxQF7gopC4
NIiCdcL9WanqLEXXQ4IZODF8aRzhXW65gptbMVqoas+jLmz95mCrc+tNQcMGhTZQx99aKPtdw5eC
gh0CYjFn5f/NhFoKT8RD8tmhsalFmKxPyQqdpb2oVSXYoHsZcrjyWMNqMBnILEbSuXC3B3qO34ec
SUm4N+Fkm3PEFmJu3eOf5KsUwpHK1v9L/LjBMxVbBAueFbOjI9lP5NKSftUAr1UuBHxEfXhDaSxR
kaONzQ5uDYLBDe/m5HNUsh3I9RmP+uns4oMsrboO35guox4d3BUu982ZwVFp9vVw1MM32m3xP8tj
Aaeolbc193OttEQukmTzYsRcAJ3S6SAnnqdR0Tq9+f/s4US5y327mhGTDBHjdmqI/XKTLEjqpUj5
jixwhvuDpjx8+e8NaqvWrpxcA18cOlLyb7Y3gvgsRjSTdsXft2cIBNHQKZwZ3BEsxi29D524K8kn
9g3h2WVP3hVRCXushqPOz1c5IFJeFowboZcy75plyvzjiOzrJb5iNPj5OSv1HNdHTU8laKl570zJ
IHt+2hKKKFRUGv9M8WyTsiSOiDLwBDVpEttJMK6Efd92Nq02Ms+Gb3nxhx0TSTITOzV2ujjlTjly
t0jYCUam+gSZKeEaLC8gTyPCqfCwDqlaGAFIyFaR6QCorhpR72IRp61BnAqlMTLQ73NnLxdGkb8g
yxzjSl77X6At0nG3lzVCoPWBEmOEsrEugJh3hCsnQIZdYhnSRuSt1tn1HnMWlwQ26Rhbg1EGYbe+
Q375EeMLV3+3elVOeWPK+3l4rvzD4VB/SHybaG6GyLEacS6KoGQEusEs7SEVMr3odgLohLEEwesw
E/yPe0NYV8TeDJxGRaEPRNu5RUMFFMwFZVYbkYi4giyDUOsxFMDOVwgLoa8E6dCc2gYMJSqUaU8i
nyy8ajv5QK8tIraQ8mZVGsspENRI7hMFzuB1LnvXNCdlRkV0eXJSoC05cn5OWN4v/DtNNfz+nGkr
egofK82op0hoG9QTntArfjgQjPvEzpmuWkAORZXEJsll4lqqhviLO2sb3eJtW3E6oB3ZuvmX6ccX
i1rFf6rYpb9vkvHowIQv5Q5/OB8cI5JRIeZo1q+mupwWxLKqk0OYCe+5w0qf7zRkdeON2AF6Pqaf
pmGA1xmuYlm0a2FHaxoVXB26aqj8LI+2GaFTy3EghVP5J9SYf8PvsHoGVg5iZu9OSSSt4g+RgzuE
ZBj5o7KnWcUBqU4B0WgPTWGu4105w5eVki+HI5XvllvlhEIyh3m6fSod1ob+dLDqi2eEPsrJqkVO
zhrKLNK6pYc3G2ULr6YZ2TRcVsMoeF0Q8pLCYDneevx9rdAV2periGwSLrEQuVOlS2qiBWp2G32e
/mbSSu8yeNpzxA2KLOlmVEXF/j95f0RxgIU/e/OuIMbqOALfjpzxynS6gH4ZF16nlGERntZ/GOBn
KwNebbDddGI9a3FfMgABE8rZNzvSebs3urWJ01bt9Grd+D0Yldya77DMqikPTpZxegrHrKpyVcmb
pe0X8JfCew07nTNNO+InItRPpkhoA5at3jinDf80taAdgDXaEdfBMxU9c+XfM2NIkKsiYCCqH6bi
p9u8ql7UeeuNOK8O8gBsQji/V2aUxqx4nbORpGsqwyiG9YEzntkol3TkFp5HfBCzac1wKYa7tbjW
nm6UDK+UhAUW1NtUvd4+f553CCcmN2jzDRCE4L9YtAXfiIJ+eaNfJNUJGJl3i1SAr9BikRNqDF3n
+/DYcVzwYoTRJByVRaWa5zsbbIHo8P76ksXi5sreQNZ47KOChUMtnf4n2Jsb61fcoJr/UROSnOM6
A4tC4wYOHQZ7gXv1oOgG7UrkiQk5oqb7/ATRzl+3tpsLjKZJbBVYJwMp0KBoxvImpOwlggKK4oe2
zPDMuFEkucnAfIey0wMnyrs9YG0GCswFqbnihGja3zfRkL49TaVu2XOKu98juNQ21x/O0lKHLeuM
JNK97a/zN1UxxjsnlEVL4peGGHi8uhvrXqzQHh6gi38trChP5qB2+Zu7uSxhM6a00TDFhsbYGsPc
h/gRaNhzAjgR1b1DNjB0kiFb7neTZyG42qMpLOd5YLngfw93jpOcDuNPGGmi8tD7w96O2oDnSzXW
C/YFaWorAZHz76uMknOUS37ksVQqfwVHypv4rErx7V2tszJLPR3iiKSGbwDOy5H9nBQq3JkWs3Ma
lGNl/gNMrk6WFk00GFRn5UL2Uc2eB7n0CGB2Lxj0AR8TnZV9nR9rZYyyO5LBsikVqq/n1wCE2oZr
ubNu36Y/E7hJQA1rocqYnOsLDz4M3Wy+0MnnlxJn11pQfl7K38aVhvjZOkZKRStqPX4UXV+AySTd
5JtI0HmE1HlRdC33zNaitbZirSgCqZVP/rXXdVS22RyMpW+R9puvdfVx62G3D/nrd10Q58idVK90
bcX+Gdoy3tq1EB30Rhy8xTlQ5d+g7cCnZDbKANxcJ+RmJw1LaZjCSPOnFEH0LxdWMLLvgQYEf1c4
yiGrbDGdCY+WOBH0eblcwkUVg9bmpJbQD0sq4Pw1UwzGf4ujVBbLeSBiG4bEIyxo8U8WnnR34nXP
WE1GrImtrDibND0RQYtiI1dLzAXaXM64PhMRlwOkmHGxAnLZ55e5n1zp90Orj8ZZB+n/JY5jl+7a
IVXcmnJd0WKtVc9xEqLqf0yWfEtrgpEQGiaiiS2EXCH9o7vlu7+C9h+Upb3wICrKK/MdbyfisHSM
sNrt+OwBk8MQSIiMXszUZISiVX9rRziCBhquiRJXcVKlHaMzolNoIdwzz0C+ftvGc5Poeua+PLJJ
Fifbg6mo9jO/dQdXaH7NxXpa6TYXU2VLZWRybd6wz58EBg5S6rTbKxkWnzn7Vx6EWjP543kHBn4y
elOsghMcC+bhAC74WZyGFAjZi/S4/j1RAsvGYmHRHepzn2bQSutFeLkNI1o5sBBBIIvqeYT3MLut
ViqKu0WV6k2a0m60kgz/iPFgdigAEURxE5ovjy1afersw7To2JUVwUrLB6kcgwJAA0GsvZ/fN5sp
mU7l412GKfz0V/2QsSr2aiKRI3FBpUEOrNxS6F//5wUYSqMr8sXFUlBJIMPIh5fgacxl3TcgntxY
0dIx/8oQyF0nqTBf9yqSaXzKp/HgfPHp+N4GXnjAacRVntHmS0UpTTzNIDkpMwZxb/g9azB/mxqD
qODgV1BGo/pnDbC1muJjgiZUnflOJZqt0HJxWwBmbJsWLgrUVQwahI/DDpxjjwGF04ikXLFnEgr1
cPdVfvmKl7DogWBF8ImP00f8kvuuwv7d5WKdOlsRFm58P07Z0aKEMgsW37jy+6PRbSAcJZW0sSwf
Ls66aLrnCZ4pickuFt2Rj4mh/bUqvzu7Hu0vcNKjbNA62zobEzcsVW8PqjS7bUrRsYW36RMndr02
QQXYfbIDhVX1MjKXzkvy6KeIjKd1p59EtAkWEjzgk9Wza33QvinPZ9MhszsLcOw+i5qs6XA5Mx2l
Ssp+fAAQ749iLbc+d4OqXeBZFie1bGeQV6Rols0lEcK0FRHw702ao+/mFl3N5ni+UpRhm51mIHli
mknLzSgnDWOrtB8JPBTR2i4eJbPSuLPM3Xt3H+QkrPkoFnp5nHz/bB67z5zeq/8TywruarFZ4zTY
Rf/bNfkUIjWXBtkW/mSEtqOU6ooekbY66ezHIaHFhLFyfmgt75JNuotlxNo0fV6Rxrs5vOxf3Tdg
Yoko6MkwmIi5NuYY0CyqOp47yLKFY+A+d5MS9ro3v28TYkv2CjYW6q+/Z6tEM7lYVVPis/K/D8EB
KSEJ8vGKnjF8u5b0b/3vQnc6+Xv5waQA3FUct2HELZWX0+EgxBGCEOpDkAXXHgG/bEKmjT4nmCmO
MWoAcCNiCueSspsOKFHaP6UsNxDEIQiiPN26R+FAxuIQbSyUZrH0nBv7W8OzdRC1ThFhYt4kwKLu
aNZ9MofqCM4naLMed6YK6qk91PMh8upLkdBo1UEM9wH9oEcFpFH/9p+QnAbnUyw4dHkEPHoE/uNh
KZuMi/wIb0EXq1rx16oMGZ6t+of3XPC91w0sr1SHJ7Az066WfN2fLu506HLVLJSLtL+R5PIlXmF6
H9ZMG2CndlpqnnTsnwQl6sMy8lG2Dhyd8V4JkYWPEr79kre2JqmcZc57UHCCHgZFeaW7expjPnr6
7apHHhApUBG20mOE88BLVQn9dFg/OHIEU+gkHE0eJTiwPztaQy3TZPFhyLOQh/H2K6jKhubMACKD
KUwm37+lmaCZbEtk0GtIUnIp9XHQjrHFOJIHHDkBfsrMTJDQ/H8vl7JcleK2iJt4u1aKxOTJC5SP
YV+1xVIQZwCMZUZ27WoJI8FmqLg0DTuC08K/0C/g4VureoZrrEzMXwE7EAy/js8h9dsFJWM21u3Y
Yaz+SHtE1X6h+nUARss/OqLb4iyeta5ibFRNnK3UL4cDdZV+aalObaOAkxDwgARY9nMT+PsZ5Eff
z7h2mGlYK1F8ro6jVIoips4FQppIvJo3Vm74pGr7SlQ+SvOtMmhHgnmtu+IHG6N6/6AnamXCDt37
//RpEoqLUC29o9am8t8/F81Q7o+00KwCz+XZ592/rCl8YmK9WdR3aV2MR9/HKl/7kL6Wc9u4+evq
Asi0uA+DBXVXxAneJROzrVrjDGlD4pstVOdnQFow3PII05Ekq/Hhxn5GosbzVKPylqHiBbbzRwJa
4KIxgUja27mMvCP1UMb3udhO1qFyrHTHI7SsTiFZlf750d5WSJkdwLGt37HJfaIHpU4pr2gB4h4K
SXFxDcOP2dK0UIyX81tlJuc9h3HR0VhI2avyixD8CGqfEiS2//vAQDBaEPVXxKbGPfjSs92bjiYv
Xy5K18AI5HFG1l0Baj3qmr0Fnye4uibs4QHT4P752YIzk3P6N0NLMxa5350XCh1bp4/NwVNDq12U
R/KV4tbov9dKn1ORe1ATjAS6CleLx/BMyLjHG7Du4nC3F/me70zRBSk8IcB45+u3z/QDJE+rsukS
aycch6m0vKj36omrU7eFCJfrofqcdGitGHXJueUMxeX92vv9JoqBHdHw8Xe09opCbh5e1aIIDfFy
KlZuRhX9DdYgJABuoBcgNmglfdrcGnFMsZ17NidIusNSt40pLdQ5dZlaOvND+xrJB4u38JNnn1FH
u4d4mZzlZd1mjFUDyCZBvEj3sQib+3tyqehc7x8BcqA89UUxSWKSIDSXLCqOnlGPry+ixKBvuvbj
HxInloasXbmewO/oiSbEsLHJEXF+NjzHDbYIef+9k7P+ZCdBDpTN8bNo8KlIPv2xdA0p6imLuxzL
BaQCE7TWm0tDPB5G1aKZpK843fFKKif8j8uTjeQQqyaQypnfs4J5seBsKWAE9REH7VUiu7AbTBhZ
ciY9F1hCDlTzpRtjzztpEieG+RXvqfLqDji3ekPO/mSLrw/hi+29JoMHpxq1TvMFfrvK6JDrHag3
e7q03hqcV7Us4c5s7aeLdS8ayn/3BTjgto97WFIaMr01yTfTnnwM8qc91GOqW2dlsEflOfSi1TQX
ySENG6rTAQpdIbJZA9EXTgn/wswd2gmqTJ27TS15286tb/TR4q6xcP+LKGrXCsGmt8ZgqBU+2SlV
S7Wig7FCfEz51E/V45qtdm10xn594j1PTAKAXtiH6CXB6q1S26IsFtsa4gfyozNhQv4Ps6KNAEDm
joFJn3aBoz+G2t3mplP6sdzTkQQ8swozLlNaTkuxS+U2lceH/6WcUCyfIKZtZZu0YWFYvGI8+hEY
Bc39NLgEaMTf05B/Ups23c9yeZFOXTNdxROzQUs93bgd/jeM+8qhH+deC56WHGACJ3bm3KJHbXn3
nGKrunpja2NDoNqoZqguVvvfprCXwGZuopKkwHSoOR+FSZhPc3WB6DPnH3+8JHobwfLQ7eBtv39M
Yysfolcc+y5KnQsM1Pazfz1I63Wuk9tSdGVCHR9z3gJJRdfDYkOlJs5GwAvfDHAb5J91vEVmTSe2
X7a/oqa48Xx08e9B7OLSu3l6lF7Q0VwKqFG7tyaHbX9AhSNyQQHILfPtP0Qi4Qr8iF9UxTP0z9QA
uPeAaE146BwEDamC2DUHHJJjgWHMFi1wqyKSka5wKPDjMLEqHMyurYWmBInvwOTVe3rBacBfBdXq
Xgmb7JpFJErCaIcSznsfDoDdIGDiDu3aWk48EN057NTVZgi6XFFb1DBuJgEB4en6LqQxShnZxQt7
BKaLcZCNXiNpQpcXyU/5hjfdlQ0Bh5WiKxVqcmNMcLQvtOjM/DEwd80LPpM22uuTXGDf5WaHLkHC
0Jma0jputBqpcIEvjVDwo8KlNoILziimqnmX3puxf9WmqUAFEhRfQU4GVBAl/uwQv/b5PQf70qKK
Rd55F+nRy90KiYOQY5lkUD+1srpQLHcN41GRKlgW12RmJfNHXkAspzoEFFfXPL/MdkPun9IuqpcN
biHpAgwxKnBnleiNCIJ3DFDP9C1xcppcGBZqT+KeSLrqMLI1INhpsDEIgPgemK6IK8mNXO5An6tq
qf2ikpAgQKOXV4qDRSHQ8KIoVQ+Q9dGAu/zADfxIVPZXfbFy2v3ek5xkoQ9RNTzWkS3LajZ1yt9F
L6moPxJLQReTb8eJ8REAWTIT4N+6T5EqBuTfSkMRybATFWr0A0JMqCOU/sD/ocw6Vk66jcNCvMn/
AH6LZ+QezMWipPEkdWvGpXb97312m1s/wHvG+dcwLoduV3646g1mFVr0Qog9thtqj/bzWBlINyLl
EFtfXLiOd6+fuT3eaO9kAPh/zYNNmglkLE0ToXCykwlyIuSh18QG2bF+1MoIUMNt6aKdH4k4TT1j
1wH8Y6KONVvGqHDhM1C6+3cDVwNs6KHEXg1GSFvTRWjzZGo+m5Ovl4aT+gU/vX4evurkVBPQ1k/c
+PJqKFTaYMlRnSh9z6p3ik0qXbRINm4K7BrxkdOGza2lANXNnFhSEqEOrSg0Ev97WaZpE67CWT+e
Vn9d5RUMy+JLU3+kea8bJUEPIyGRwOkEAQgbuCB8YZBIYGfHKUFCbhs0IhG02T5eO+7TPtDY7Oom
GFZLROp9nZ4Bz0NrQ/5DLhYEZeSE01ZwvxwK+OJENbLdlbCXXiOHcyXvu2BP6bVu7DVxyD1efZfi
cYU2eZeZSyBayhu4e5FzcJVTS+kXyDE568Mzwg2fdJ7ZdtYV5X8jfo+NJE6gbxqbweXW+nY5SVOA
UYARWgLJVm8dLQv29KM4OPISCqCLAw2J6MkV7awAkjHX6b1Wt2SVVqqNbbi0arfpqM3Vm8EXqL0o
MteJOiSB/YQbhfh1EqAN7Qs+jfwRxxOoPVe72I4XtYzbjDCQEB8tymrgeKnOhiTRWUrIM5Zs/n8m
YheVXcQ1rwUYWomoKXwNFPcw/1kRdDyDAOZo7HAA6a7WyZvQJUnH53cF9nvEt6kiCmT/3yRcuaGy
5lPEn63Jj6Rl2Fsal5RONI0nsZYHRbwbfEbmBDNupjUjYPD6fPod7+56Jhh6oHUxg9+Hfxv1XTDX
haWNGHloTSpx7im3EIPBNL7zQG6UoQFjz+4OvYgZlIyT3xJ2KR/wE7Xs68+dTOihZ96LBO1m9wVs
r9T3qEZW6lzTYi91TLJmKn3Mro6OKkWdMLivrMEatYGEoCQ/m4/KPeZwMlBM87ht3aBV79WKP4kz
3xdYmsfDuv2NTPoP+II0BrbNUXwR7DVGG2aSOHvdJgE4pk7W+1o8ivT/YDehbw+SKWoqKDRcf2kB
/h2p21iUh0e4INKDj4NEsr1aFTXx7AARsTrSIQKadBLrHuvhLehPApaB4wiOHFryLmdui4icJfCv
nySfswIDhuA3YDsGTdOmaQ9fzq7PfC6QS9CrSPndGWZA7rMEMxzleYduij/Uk9kjCtAT7D6o5Bsb
328TD13HVSWG5LP8EyBZNyimGbqNYLMNm8lnX5uD+g9aXcIa8d9OjANIzzbea9DVYBBwCbufLiiD
HTEPVrwJO5BcDP5qMXSFlXVfAClyFRgBCG9hY+x3vNgooxPHqFUYhT5QzTc+NlnOScKp7kgOHkRf
zElUm2mRjdLjsmqcSs/XaZzOT4xKj0+Z9B4ueKl2N1NuvSytmK14Gi/kx2xt4wXhQpD1icfrM4/z
NuRNxmLZqyPYmGT8YCgBNQLRfRFgE8s1PWVRaVj2mPS5SF9EzANQDNUtuE4Kx0PJ4ZYmR5xB91X0
9laGnrbMduCkHOf1ZSvIsMWUapKP7Uds+7nX4NdtOdKlijp5opGJrDG+tzWbR7X7NSAO2VJlg8o0
CehaAkSQ3DQb0Q1NTh2ZDtZfxVLlFvXaB42Lw0yar7WjgMRidFVsvylH86fqjONzqagaNtcLAIzq
nyizRnKD8WzTVDicX9oZMBxz6PiUSnl4srt9yYYFPz65mDiY4InJ6MSE2oVK38uWSd1J1WJZjaNV
3xzTH/qYAXQUztbJKLl1zmxZK9hG2DpH/ukTkZdA60J0X+4oj6PZ5hVyhWqx03Fm6qSUDwVmk7yq
Ycy4HO1/z9XJDffGa+d87PobLRrRQE+3qQcAfzNXitYuVKXlRs9XtWD9q1yq6fbv/XIrwZbNGdjc
huz7+FgpJ7Gf+phMmhUr0P3hB3hDtgGL/5mRA9YBNBxxG8hOTzJGjPnEoM3F2BXqXn9sqrvdjv0N
0q2ficbvN7vNq7qM6DGiR5xijeFRCTVxpqm5EQ3+QH5fkg7hHpWWPGrUl0txqqVGFJh1qIDlQEu1
iIxb8bA9iIein3ZcHJGrRN2lYlzVimkUnryKQA1y2OIjHuIeK8mhDho+Oo4T7i0bTzp00KvS8YgE
hF+J+Jhp4DOaf/yhwyVAXySYyxo2NOiCYCEz7KGNnuzPIIiY4kFUGC/y3fTGrxQE0PQbRp+HL81F
6m8eZmcfnZQjeyqZrLkOA68RaxbSF+dbBog2nsowDQ6v+cad8qsL4yYL3Tw2+1ssQtw2b2DntXON
E816hzI2Use05O7Mgjs3kmdhTpgj9KVK5LE1uLr2eng/MnDN9YwPPD0GyWqIFaLCErznqb+f3aRU
zB0KA09l/6wiLZp+fRhYJLPIsl2lWA1wWcQIgBjtMLIGDPmAhuwnSOcfJWczyGy1N7Pz4ziDM3zW
/AVd+MMyC0ZiiuAIIrY/ZMpxO9wE0XlH1nPr4XTRsnyFmFDdHzPK/M6eKYsb1a6TGL5ZJe+wYcV7
fc38LmLiXvyGpML+Q2hoaB0bWsqugGy6JubXVF717YAo2VgJHMIImCbv+0iJq9XlO5Hm3kh+iSsK
o4P3Exf0j3nZBZeaSy7hcNb61YxWf9JYWOqR2eS/COXIgLzwll1o0IhkSaOFu/aul/Z3wdlIYtld
qIEeN0sCA4ZQwtiSJ0jNtbxbCmL5//PhObzf/Mw34DxqungNZXpA3t5mYrWgJFgANNaS1qm/A4cz
RZQheKHu83ADKlBcvR+amcnvD7olm0NYivKXzffI1vvHcMeGSlfwSwMzExulH7JwgAFFgHygdlXU
N20/7pJvb4QFPXWS+Er54ABQF72p1F/lr0c78wo6w5rpVNmHWFdny47ina9nRWPIojXsRrE6t7Ak
7kUZmZEHYQaM9sWp/gzzRi1ov7ItYZipal7rk0ZPuqlh2D5FPmbRNam57nbemni9fc6kEdguxqwm
oijvLUHB056eilvFqIci8rMP3dn1WcEEdFsI9EaHkS7nVGfN836uDna+D7TgKowc3J6/5TneXeP+
Jvb6J9v6kTidGqieODm41d+HWSZNXwP5YiV3wsV+HB5GADD9k6T12C6UHz3i4edjwR6KWX3jeh8f
8wHwFLZ7zQpON5AYBXOQPC/Xm+qfpVJ7uOk9Dvuvb7pypxd5QO/T4xq8m2C0bsVjDc5Dd6eBDgpu
RMnxheZBIoATfNMX5a3hyGcH9fVO2z7zYbd8ekNgTsJdEA0Eg7HPwYDL5qSaBppEL2N7zfamMOOn
Xpln0N/CZZMllvWA2lYBnk8aQlzBS84xmtBMf9OQDvd3HCRNuUSBVMNvEYvfiB+YaUxdC034nII/
UxpzIlvGIwZXad5uRM6v1pUSCgBvIDEU8HLxKgFqoKoxT+9QICNQ7EarBNC/3lxxnGVQr/70aJ/8
I6GV7E2xdA6fuCoJhGNzjhlYHcgeBkv5ecmx2flybOkvMLBY0OOFiEJJyVDC8uFScnZyuq12D+Lm
kujJJ3oYU7iC9ndwfyyLOW/qkWNKvQdsGkU9zplOZG2wfTbknDhKiQ5VR/rTbJ2lo45DgCn0l+Eb
LC/UccDGayUNcdnIKQ+agd2I+8ACsx2UDFAkdmb+a/xSQ5KOul2OHOPYPIEhTSAPZGCM01b8ANlX
Sdgdz/l5tgojYTSOvrupbNG0qWCpIyWqJ+pAfQkoqJ7W2FGEARJimKYA3gtjJ6xp0PvBH98565tB
L/ruQdj35ha7HcTu4+oE8HnuSlbIBWh7AsZlo/QCkLxVA/zO6ojLe1B6JXTnNmaOG0+HawwCsF7D
/WFYixTupinxPal2qt9QFkQ2h0u+Soq56IEYQJZchuEKqx5f5vNyk9GJNyG5HddJhh4BulY0LvUO
XZsgrYi0WoIeAJgBqkBUD6X/OqN5KPwK56URMWkiSucTTCNzsAM9GYr6cj4t7jOepItghTRTJB+X
sCUvKh7LzuabvKMKkPd9vPxEMNR7jrIEMm/EHogg4y9enN17V0xDa6tfvxYxFXoZoXkM/ZPZvKvE
tMQ6HLVHnpdKBf4UUHQ5dzF6G0RObPP39jH7/awMaucqYCyMMD9fdH4OL2JvklCeH0vd8wgecFUv
CNZ4gIPP2FxHCLLCZWX10khdQfa0yQGKgLiJ4pBgabynm0z2K5eHbXlETRwlHzr2rRHbeBig2QDc
xTLQTJabjA24Q/H35Ym83ORwCa4IFeazk5aDdaresuY52oxr6++2dHSIya695UIpN++/VygyJ+ms
oWjtAffgFrhCIHX885KbnCuyvMXqe8W8+HBwUbBUS8jF3t0R9QgqU+FEpGa44/TZWBDfosJfJTg4
6XWRcSApt9hHHPRNJJ1kwrJOAnMkCn0P0NmNomggQ3RHuQ6TRRd2jRHzzVkZCMFN0HUqPNDxEFWI
xYUXanl/vISFGdEPDclE50cj7J3j2n6fU2qOsLh2rVos/q5HkfoYeKITC6G3XpGwjbL1bcZwUX+l
Wbkd624lztlwGqIEf56m53c4X9ofCYCMu0xzsUgkzEKv+F2VpeUisxi+wIgMBICl4pGjTPo60l2y
kA5SvU96uByprzsuZ+D0fHr8lWs80QDdg/dlfMxkINP/PMaZb7bkodPwBYYgAR5qUafeBQC1mJMk
bELIFiiOhyk1wq3CwUHXQtFsIvMCIURpDWYYqM0C27b9C3EG5lj4AhJbKjWxGBjKdH+IKSvTWOMk
T8IvE0hhfpnBOfN0/vnq5WXL4NfOpBIoGysl2nFSJdGAb6xjiG1W3lWxENiQYrpE+z6aKf/5VEiV
icqLPCz1qFB2dlkmwISKGMT0PrFaLedKTF+nr5SO9hNfnLO/FToS/bMeqjF0NxxlCD2yusP3M+iy
g9xgHMkV+RiNcqY/teyeekCkC3OTio8KBPBTIZTBQxLfSfpSyoUTKgG0slzEZTBK91ovMuDLZWR2
p41Ad9ucMzzTNvc4/LG9DcHb+dmTt118fA1xmOuBzWac3eV7MqMLS2bn32bkH9CkiffcRqLxKy22
+K3CHppiXMHdB7nZ3gfhCMf7HUajAIcrKmj8+7meacdbxriduCdTOFzzQieHeSfdoKiCEYmf2ume
olCvXIdU+uBwfELycxlsRqHhcWgCnXuN6hDIYQZF/cqGP6Wc+gGOLQP9oJKmmuXtwclhk4LZesh8
R8PJTC+GfNlvE9fWW/rzBOdLK3RhMtBPNRZ8PoRJ9vh5QtrLUJZ7xIdVzxFAyZOilMJ0jdK8Ql4d
3tr2C8vMxRSSQSUkKbEr44dpYVCUkDCrRuGexvxWFnahRF1vOD7p0vI8kMzTuoCQ3s2g5utGFOxh
//ldbzkG/i2C4fXsUFs0Zudv5yhs4NflJO6j4+43FJFZhiIo1CsrFQ0UxzzkUOg+Xw/+4UpW4UI5
N+rt8gUARh7X9icXVoZS5DhjBZ+oIjR2umCZOHf/rMD+VzA47KE7vebl2e/K/MFp8uxd3gn+R14N
5b9nI40t8PK3OcY/FP5X0Z8/+ohmos3zfQXsAUXI0uOEHrHnriTbTUd3g7gvLQGBLlZ9zwLhKvvq
+rMXOhvD7a77ashaaSRQCFNqYivh7fuvPc4Mczt7X6DbREphLXKYEdHdVzZ6WVHRdRoENKHyPJHy
56K9zJNOlPwVdrtZFP1+/X/bwj+gCF1xElHOddWrFlhHJM1gwUoCFTm/zlcaBmqygVOiyVkgD+q5
d/EsZeQz09Y2sm5VkpCjemyf/XuKZ3mwa3IFi5HeVwfF4KCjkgZJAp9AogdbdYo3G82PHtKJaOVr
HPy2Jy+BpV1zXAookvHvc5MsxqgIkqfFneFXEZ8ExC6rzgnQSqVpbtyBLUuNjRJRYMtVE3TeMTjr
oq+momQPS2nMSlKYTfY+QoLuECGceMJxHM2Ts0wWp6GBHxAu8GcYhCzlwjSOEiu6uRkfqYr730vP
HK/iit1x4skMQl0gwQgu7ZjUSikNR5ylQ6MNNSjvfJlqKMEiKLTJKcmGZG1UcjyRpXa7W9bKDA1m
mgq4dmbaIy2OLbzfLxCXWd8Qch3DGXrlNe9gIpOJ5vL8Z3GVHDWyjJ9PC0nZ29S/FMe7QADp4m9p
4knPzXtXn8zbijTKh6PGaDBeVQjDnC5/iMpjhkCSWiQ4LYuZIT6IiS4GiIvKYQrHwrE3n/2+o7J+
o4ZiIk8Zpe3QwRckahvNAYOTxkqlCpYnGQk/N0bkQIXOtYart1ix+0LEaxg7hE4KqVhtNEpxI2j+
2tzSf1bC/GzozFkkWyA/syU+USc/+Q+FNidOvP/sAzODPvaF5uqL7NfVA4CECSHlWfGBSUXlVi0S
dHQE4eMSxbgx/3uXfiVbpJBLFIRmkYgFQpIdN2wcgsYHOn7vl+4EtN4nfv3bh1vTifYynk9NVuQB
e0v7RX31rjymgTfZcClPeZ2MDEi/uxuiHSR9VsunftJ3ZcHA2Xr+5hTUcEBmLNpf3tUhEmEPtKMW
oQDSbmbB+EJkh/pITbRlMEgS7HaPa21QSNJC3KuG7obeVdGQryZmBhodL2j6P4UM7c28IkFmgh5g
S6hlqlCDus+QklF1XWiJtComaRipF+sLhI+PbF0fbW+8xVjY3IzurrzwmFbQKhcG1szEkrWk8rT6
dC4w/2j+SZGA8mqCPjLFPa8ya8va9B8KdVadKzSGcCz2jrKJEkkJmO0OTKGXdEP/2Og26c6fb6n2
rf20VYNmeibp8x8zh+GkEFUx3r58IrApwOdO6Bbeacjw5DcRBjfoOxgsyiam+A/JBiCKUSWqnkK4
uEIVDbz0A4zC/6xzpEx+ZrtcJIfz+fogbKcHFvc/tdLKMp5909aFKi0VE4K/LXDIpqCAu2K7PZa7
L7pBqV4uOXoIAsYUVgNng7e5wWAUFL6RZpd6bJbl+BlFg0eVnP+ttE9ozY4zfNDiOde6psc/sV0z
YcXnZboe137TczcWhopQXwM5cBjuaRRAbOM76T9/lWZPKa/SO0CTk44LUicMZDYVDXNfiMNN+RdT
b8m7GixH87vc/raPMEb6jkcOv+0m4+XZf7R5SiuMhq3J2+xWjzWi2MTkfZmMA00qw+tyn/R5ZL1j
J57dm6fK8QVshLxcsvTdYFsLZL/gc/gYb5ETGE45WtC6H0gaPg1ZwQHK/o+z/6EWIANtQPVfL7WG
dWxa7G+brg0Cpq0i4w1Cta/EUMM1FHcRgLop2+3e42R2NHQUVBhOk+X6Z/wNGHvrGvDtsQs6VSwd
tycovS+IyHCNNKClX8Y5z0bvo1A45JsDdB7ucdWXdVXneJHji8neFWGF9IIci3w0cJKlq7MZbZt8
8rUOZPyIqzjtHADfriiKgCUISwGwtoboCHqtQ8/CnLL7LaK5yy359ILZ3y9nHehHuwUfmJC6mxzD
lCSsCo7dPZkms6m6KidqliIKRqEqzOqlOmapYEztcBkm2KQKPbGWqKl7l114zqOfFxQeneb2qQLW
XDKa8MunQz7Wzdt/+M3jz+Eylj1SN3rT79KmG5OuLeNjujGPN3l7KL6x1CULtrBTRIl67ewyuR8d
b2PsJqnf9Te+qw6lZYm9SltBeUHlqGxSmFEMxMqjR20AHt1tI8i0V602srWjIy+ZilrZg/flucRn
7/Hlftex7GmgE+58he/Pn7MgpMdJQbf1bmnH1M10/QzIhUc2aoBKcUjUJiiv0s06hoI6WyqBGr2L
x6GzEqkDPNxc3MucHBXPpnUGZTqgo8NOtUFwYBPkE6ojDqurbN6LIN3vgwDttFAjMOGARSHOribD
tmrMc4FeRssbM5tq442pzXnvhNutAb9XhOvRX9Rz+m9srslU/wu/TwdbM5llpEthoT1imPxs261x
EvkSMo/AQM2JDu+hiT1eWZJaD5sGbu2F7Iw1MGoaSskMNTBbnZVA5Bc8B0Bqc87FSU9FGk/LbW1q
1vzG6dJMZVi+7gK5Cup4JD8bZse2gpyOETVt/xVqlvBEa/2Qy9nM7iu/mZFuFIlae8MkZ++1P2iy
2BgWRt51RK9wF4U0SQlA3jRJTsPvqlWRSyYfl4Y2FhvobzcBYN7NWnlbNZz3lR1pguqYdWzCVYEQ
miV/uHaBzlrlAymyN8NhHOxLa78Z8dV8ocpQDMPqw182/Tyz05jKon/WFC4RvSzghB3oWFhvDGWe
ZOQXdTTKGRwRmv0y99/Q5X0zxiswgXE/72L8gX6yDNKQOSVlRxjuREcvuGHLcD6YkigQ3wIQfY4X
+vjeUFnH7W1pWhvz/jfpnAzC39bM6uqGCxizTjl9hUxl95Afk0IRuezpzIXGiRAVQFVCKZ5fyIoL
0ptEi0l1zbouyiJ8lzjQSu2ZagKDKUyLgybWQShfMlyeTkLHVt6Gzszg8+6e8ZGbgnEDIWAmUkX6
oJoEWqeqWM9JWzpKS/7YCWSUfJDt+t+YOzGjCxWrQRlGpIu0SD5cVgSe9g+ZcOQFKxIWu0KSY99f
xu8rliApscIGMT0Kld4XeeSQl6Eu8+rLl/UKloH05WzaRPP5nvodiz5E7dIvF/fvg7paE2qeBvWo
IUCtSQr9Sn7RMnjUwJcuAFCz2LsRqqavZLgzhSco+U8YYf3338sqaAIDDRYcIAHwMDHLdDo2OccO
LGmZX7e8Hs3MLcuebF6m4w6U9Gsi61tXhKzhb6OCg0KQg9Z+8uTvhl+GI0uDdd8wLRbQztS69BuB
bnh9a9ixln51fArEgANXjoZ5gm36fhZ0xE99X+pb74631jXuEU6U1XkeZyXjahd8tPlUoN3Aliy3
vm4y6keW8CYV/i2OQsCxqsb+x+2GFfAu/8yjEQ+GbVCS8qaszDAneh7Y82lLqpz3xc+39dAKg7BP
SqjkpuU0GZ9uqkdRzTBxvPC4oGf9tzNyUWzBn2yGVi7UPJ18h4b0S+01KuB2pvX7MRicLckTT5Rl
duBY2fNR1ix7RaljNKLaECeecjzfoEhMf2nugMlzEJvI1bHi50TUhMT4Vr+uFI/T3T96Vq6C9AJ/
ReSU4ssKBSfgmJmnTn+OKgN5s51sbfaFNYA3IEK2KKr1dYOrg+hpmLU7n1zSUM/KliruByQDXYbT
yeK2dFR13/bb9BZ0YBpdCLmy2h0SauNKqbkX7KPIY7Id9g9b/z8mS9POSbba4rzHgUtqPMnZQ1dW
ovdjhbw1IHN4s2swVi3Ds2Hr7aQo3yE8UWd9HEyCFzMH1wvcgk6NXEyj3rbn9Goo401BGyVZL+FG
IYm4kRBJ1CNw7Zykj9/kS2TSQ78XBuTMTqkQJb3vA1t4sduWSpi97yuJ0nPN5Ot5R4AkkoTyM+ym
pYVg/PKiH67gRL5ej3CfIRXc+Ndl+z29CuX3kNUuZ+2JLNUw6Czo2wYOEgbwb10uqkWdg0bTTPCz
59gzAAr9GwNtWGByYZzKbGdao05/F1Xf7Kv/gFYN2NQy/kBRWXciKDMXHAG4g+kpBwkK3OdyY0JO
dlxG74LW59ph382ntxSBOySzWUZNM9yfi55QcbAINNPqreVTsxcPclV4eY5b8PmATuGe3Oc3xb2s
roP4nX+aEijSqxoyZ+gYB6qLIxcFtAHl0x2YeT8q7gRbYspdqw8Tt5WCzewmlNjsQZq32Kq59Kic
m/4Jls/MCvvn/2Mn0GNsrrZeAZsX/oZWRYEjai8m/T6vapxwwmI2Hz2T2Tq4hgcWRCG1SrBezSAd
PmGhAxEqvzPkmISoxG6WOMi+zNNav1z20S3jdzjcQcIP/gOndn56VitA0pLbmLhfZCEYm9nDX+iB
0kLSTV8YbnjcznWiPySwLi3hvHg495nOvedsEuJScVPGw8VIv+EyNKlAANTqiiuDr3pAONmJEzrm
iNGYT1HSZwV5LZOurdstQEz8i42FhyIMorvZ1r3iSh3qHFV+clK52PzIRRDmJ0l8P/Q7OFgnKlG/
FUn1hZwaTpuCHzg6lCf+83DFQIOw1KvV4dGmkJY/AbUaVAWPjaDcMVslS1GJvDvCELV9bDwsWyhJ
pHxI5KB4ZhuVyDe19zTe07aoKc511Pmc6t44fxd9hvoEySK7Bnvqi1xUM0oh4cZTAFA11ZyrdPIK
FMxbMlfNi+wBcElTaQB6IuHqKm/MBqZ6CqEmW4v2a7QiWwMzirwi8wY858NxVe3plnfq7IEkX7Xw
rzlfjrEcmtCJnQF4STQXkjzUmIdeLstIeVdC1HiMOcyZvigvpA9mnTdDBPp6NnTPxNtPGn6FgH7s
Dr+dn5mnY8getE97C0mUoGuFoGtuD+I7PMWaJfDi54w3mW4CjSCNg4yVRmmCwrXucS+nBtHaWvW0
fYpgTsq1PuhIeRFIqR12cByqN5W3gZy6YXt6+QAEj4+jmxDnVwnOOXGWb4a0KC8JJL3vQ58+viGF
EXvux/iQIh2PtiUqov+JyUq8SL11O0Mzka9QO4CiD1a7ZZ1SzbpMyzsxXDYgOFOO8cgTDxEYVjg7
lTkLSGAImUH0DTb8ryJCCTggZ2rz3V1HyZtBd7C7TkNyBOK2AtVb+qThEMcpEtzwDL25LuunqVpE
+RhPqleYQGh2QaGlMQJjpc8yRYy6FVPm+cf3al/0XPZEeZAmp4GXlmG/0opeqDd56ONBwh767aT1
rbVkOZqMnH80Q2GC1P4YzBokOk1SBKp/VRjV2VIrCM+f5zHGJB9wRMiBYqZpqc/AOM8Bgtx7m2Wj
W7eOfR9GASQ8fz3+nU8DO9+5AgJrTLo4ojVFvuxjTRhk46Sycv5XMy8Pr1VABgB2eAY4weOkzNM6
0Vor6Oayx+gWvZ/vfPWfuUYxj3csBJu1ZimfbCf/k7WFzAMLsPQbeo7iboZZ3rrNeVQZLC+RIHbM
dXv0kc/JxxYRvZY+PDQCrAoPgvcS547nlW5WIj9ajOx5gJVCwTcF5spW9VzdczWUadgevkgMme/V
uUlh1JnAwljhe9ce8/goHHY1eiKWZ3T2dIhbD5/6f3+hNpD4ASC/tJCAbqHK6uLKIl7fV0F9K/3j
zLJkySNcLBuU0D7ahjW+cfzPU+kPN5jM5sS1C9PwqylCmhN+uFhEtEhYpJsejBR+JrNR4JjXTEBX
Oez6U/vW+RgYTVn/adKuUdBkJioT0rrohs8zPn9knmjQaziTNPsbm1DGV+BM+tlmqrK/cLzwucmy
WjF1FZ0j4lZ+nQDslA51A3LFuxChWfWLQMvcT2ZBrmL+8aE9w+VC++7GDzLS6EdCXT4yY8QaAjd8
qsdtPR5nBy9x/knScxfppCc3SdHy2SN4sSUnAbTxS0SyjTEzI2kCrTFB1e8kE8PYERx1l+ADPfl3
xIG7oR/Q8UAIViSVh1EvECunojyLjnCJXKoPA8SIFoLtb/3zrKE+h/tboEKdOMlZVUqLh9yvcyqr
rnZoqTyUVF7jkrQxyHVkUO+iSrGm4eSc8uNM/Ye2wCYq7BjPNU2VMKp4suIlpe7NxNfTPP8pBNHT
65kWynHYePpsoHMdN0l0r+oJZkEp/F0rrdqMTCVX7me6C61BlzimYGYWi13nCq67SoHOdupaCxF5
GaEZnaqIe9W5A1S1zGD/MJBiqiUEOTmdb3nu9zyK4zeUagag8LCAlpGJl2GQw0Xk0ZeiTQZVzyOj
M88hEiQj+IrIMaDByjQFFV7ZZpsWitKGX2OqxOj1zk0ZqXk6kyGTXWDvVcN1/F4UhIQHvHLjMt0X
tAD7m6HZrJA2onpWKI94JkjwABgUUI5Wz7QQcHss5bYRgyh3VvyAXw99k4K/2K3cM3ynyky0dvgH
/9zPE9u1LzuDxHBRsnuvOFXlQj5P3vDrIt/IK5DJjBRXy7qoxDCE/tefRU7KeG+s1FdFHj1KONMQ
3dlyLbXxc+Rnc3wu43I6s9+eTi20FNcRlhIEqFEs0l0+uEaUoBh+/E81EVhX6vHSkLAymP9WozAJ
i/j0hFeagtwvOIj9xUvvetBgXpYzODFmfSZEE54aDEuupLGydO5DYBDSWmCaaiEhPLjaqWpZjUZ0
uzU8178hBEJCAbOzCPmyWwfJncjIkl9D7j0GVcuXyVEmM47TRRYnn+JOWwGKFYO1mxbkVz0lvjvL
v7nqYwJmlFzo7uuO0Ieh22TNBSEYrBDsH/uiruuemlpRe0yvk6wlTHg3QC/EL5sFhK5TRfpLLBRN
/wke5EOaLED6J0bMSWb6/dTaLkfGG8N2CijwEL6MKNly8gPyrygrutqVIArboDPNRpDwrPmzCFwP
kkRTRdUtX/FZixcIWKpo9DvMiwvXAeMD8hUXIJSNTkKK31AhstlUtpLg5eJjKX3hV/pPG+v/W01I
T+Q4rnKWgu993Cz9DHn3cBgGvlSH9kdSMsSDqJOmAqeUp2anKQ6Z+wAmWQKCCoENPNml7NRbEWSz
c1jun5wrnHtfRlukn/wh8mMdka2+1bk+cU1SR4SkDBRhkY7nRnouuanhUH4rT2IOnFX31oaqRBwv
o1eZHuGS4lViXqPvGYrwu1PiIxHDlrVFugHUU/Zk/qDHFrwyr+s1pO6asDtyny05jtIvf+MLbYXp
yQKkTIVWyd5gF0YDg/A21if8hOJn8FC1YLuA8u1eOFuj2t+dNt1KcJjFZ2Vxe4rwhRKLvjRbfyFR
AXFiltV6Ky3ozn2XpAIs5OHWOxggbOeKeYae471wk45AC7x77HpMBqnFAyCK+4EoQrLTe9tUMnOi
+4Y9keFHqE27Yk5ULEjd0QPZhzYou/6Zgwejv4jZAxUqf9Ts/ifkox9LimLqTcmIpOmWL9NXhmUH
Wq5kEQbEaG0K00D4aMm3BDc7sNAPW+gt9R6LEfbPGdkZ9TUPsup/FRT6evxzoTsnHTrWRFBGdZAB
K6ra2FoCEOTKouNUoWHya62Nv3PrfFBpCQSTOmgZ8+kaOLK4Adu4JvyG3v0T/++RmWp4wPVdG0Z9
zFiEaTs6Mp7DDHR+I529OGQ5H9OULhvKsiH+bhZz6Acw8WwJf88ht95G73+EgoYbQwf/LHKpZwzs
BPli/3lyA6nb0DDx8ulG9dvT/nx69zhViSf/v+8x5Wv2Elz/mQMrQ34JpIc3x67ZFXItLYnSBskY
H2EcDsA8OZbyR6kDOlpuQOdnJLH8Z7Q/eh1FhhiwAYTLpmher+5OzdmtyvKLeRGjwm7kYTexhPZV
tfDHtbHV5B+2cKJ56UsDOpTOIWkvzY/wWcPS9kQdZxBjh6h3A0wO00+ihA+nWsiqaD3mW15DeJLZ
Jkq+DFC6EJm9BzJlhPGzacfbYPWwTlxC4YpxfrybDR39yRyUULzN0IMKT6UYI4kMqWQABP2EQMu8
Y9nrk/6Py9vxbWUTjBdec7LpSHAx7C+3J4cHRs7mlovFwBR3MQKuhTymVWaZPytM1o4vZOOXnfYi
IpDV2nHGqga9CUrAbJMzFYcOQ2y83DkPfdfuPS0pf0T/w/R2gm3oR3FTPVZZMh9Z2D8282Tw3QNl
pW3ovnpBFOBexuZSyxtfAlA+I2iAWQMQ4NwIgtNoJVDgPbj35iT+0eLNSjowwcZpn9KdFp8ORiSK
Kw/2IQoNOED86BgFpLOQk9aJLb5zAdHverElz2ZB7cn69Zym0t1MwLpPT+r+lxOwjeX6r7VmO1L5
iCby1NGwwiA4azgoagBreZmmD1jDlo9HAeqPGkBkmSCmrLqgdH8Kpq5zVowd5D+WS8BPu78dkXTa
f02vp/ZDFtoHrKJ8R/aMrDG+y102lxjFS3FzRQUdeOifI8GlFs/c8PUBzmpyayVwb4b+NFAx6jqL
WF8+l/ZwiTGIuMo/h9LW0dZxDlqqHgIX6jiNecYnw1Tc1fQbcTo/WOLjRckCmiIyM24zQHbxjJZd
Us8rmeMwQgv2RCkA5GDRhfSaBapzcEuaAbAHH+q6tb4nt134EMH/0AXbfnzDu8MYMc6qEB1tFVBn
/6SpNjBR+KFW49DAn0KYOloHH79v5hHYLmkVjIY/FXj9XemvfM6GSsGGh1dQqsC1L8SH+s1Yd3S0
i6VHQVo4WIvYSqh7rLmjgV012MMKSlfaBiNS9CY77nQahWkLQt1NUnPNMTD0K7iczopecBaGesrU
A60wYQq7UQiMQIaokdhpoyTMJRw4ZJQxPKOiZtXEMFGhu/2njViFJsENzmnQDDdF+A7vxDs7TCvb
RR8lEbSTwSo9ata/AsSTCDRCWf39q1O+SmIMjhYtzqwVeanfb+Nk3qPLaMetxIU6nw5NAhbtRSFd
xoagLoLMBAVm52RBTnRWOH4yUhZzH5nivrv/eAKpfjI/PYvwSj2ENLr21/jT8mQXmrGCaM05ofTG
Zm0iyEpmMYUpjJA8fC9l0zNEnYq7af4CrYb0dAaZRXU1GfabClzQzbE0Y+QG0CWQ+BZpYrnDksTL
B7q64SEmpHoZR1CbbxWtWskYhSFmJxV3MAdE8RKbPr8nqNogB6hDnWanAmXTAgJeV5uhWnCxO+n4
fyGXTi8ccbOYfPWsDrbhKVaL4Xzg9JuvPmCVtn+ibQwFpO81xN27KHV9byLDzquLSX+w7pr2jwvj
yus7XhAyqPr1ky7aYSznKbIxj7v6Avdw6HIhO8jHgcUVC8qYNvjQHFygHTtWJ3g1yX6py0zdpdhT
kxDHZr1poVwN4gFLtut7STGkcaxY8dJyPAlQgFcGtDG0qQ6vlBjsG7APyXOPZqQBQh4xVSdCWCHo
5/4HOhDeilaR/Pl8oh6HshIIaJE86yILaHxMzyGG19TFQXrS8abrzerjDS/qxKL6ZuVdwKupCNat
YIYuE/Mi9Ca5Impn6+VcFKHmI1QKoNuSBebWBnvFC+2b4TKjSV1BauEluwwG5/i/16OfK9AZIpEG
c6swUbka32r8zaNIK+pifb7gM1RXFp8golBgWkcL/dmi2OSpggTZLFAWGVeK0uwidvTQ+qIrjFmb
1c4cMfkUc5tG5Iu2+ZsBAt6oIr2Xc5lrO8OMtr22J769xVzmK7EOugEjnqtNTq8ukdjERRh/Q8Sj
V9qSNa8Mq7WokgG5UgnwHFOszfS6FpxFK1Kcunp7nBHUB6DPd0JDtm7MDmi+tklnyoD54gfhXYr6
TYyjuxVq9GaK4S+gGP8URjHgauZXBxSwSYfoUnEdEvFCnuD9orsgHaWl7bjHygXHuq15sQ+PyVdO
tgBxnjBSFroy5rm28jmfsca5uLcew7bgeUiMYKQjddmAV+h37lwA71j6X27amoRYW9C3d5U1qEkE
kl4NoODjsmlAdFL6QdensfZLKJZk3cHU72QDwVAWCv7kqPTpCSdiWJTwlR+o6luYUTyQTRboTxmk
Kic6TAm42DiWw4VfOdxlnU/59l7Oz6hDzbJrAhF2mN7c6w3yqRNoLNLQn+421DarZHs8uloGxfBk
SesD00HTgI6cmgjJa9mOMZWLFkT0WifKdJFD9kFAXxH7RKyBk18xyjSG8U9/RHAjaZYf8eVL0C0p
cS5syOnRgeBTBkexeeDt56sOMeqPjZi6uwrMZhTyzx6bRwMARfXGzeuYgdRXo8X7ZPgjsw2mlrcC
HzKgZdllaL6RgO2D/YmZct2D/Mn2TMSPUGuneTppvG9lVf0lNkAyjd9rkXXxBhBTquQBvD7uUXD8
FxT7GhtOd5q0IebKfPuqyg8SrJNlnLQoelQi302dIOOTaUuTnr8M9/tNMioZlOSTfOklAKdPmOEL
Ogm83VRPhDdPTA5aBQLSsig6X44alEzbQWvLNgYJZiBD6cZQYqPwYeKxliXrozCOG5HPLmtd3j3D
pP4sg1SczkVvi/UB+pynMQCjfod1p4KqNdy0Y0TkgHHNGCGleX1yeLMcmWA0wddjySI9EcJICSkC
OcVSBCQ9FIqaA5/ZROIG0igjOx1u2neH0ankM5JnhA0ZsYvHI1ZGLglYsE5grtxqWcCNFi9Va9mB
0GGqBvOvr5CHGTlY3hx7cdWKfXw/vlt6kPtiRhoKRBuM6DqfGQkLE+sRw3tLlyAOSkGX89pQL5yb
DoUDfTojef0z0pEXrUdciFEtz5XDLNML0cczirN9b7om9FWYba1icFFTQT2lufJnZ3Ry+hWqsBKs
qvmO/W5UFpC9aov8PDfRrMFSy/MqFIrLZZ+yFwVwu0Mh+Ri19kK8BHfxAewVrC6mFag2pGeTNVCo
XYW02erRmuVMw4pZ2PDLlGYAANOF1V7nrk5ejyWCeaOII6zuMakUuTyitLdJhevRs+vIzJU6w5Dk
BvnH4rWpMj7ttOP6eAkIEvZLt+M8lt/e3zTATNa7DYVIfOl6PQ6Xy042H9sZFs18//Mt19+TgGIV
2vEp2q8L6CwUrDMXEA+DRBjhE3FgT5hzer1+izc1BWtfvW4CWD6GqUnAgc9AO01oPirJiQixJ35W
YHlm6JN4yQvlcl4Kgyzme4Lm4udgpL6wooo0re/1mObeKZ+J6o9QlGa0s0xXYtsJMG+ZjrhGpX2B
mJdTURarzgZ6aSn2n86rwcZmYJxRt9M8SeItvgat9fw83Grm8/TYjyd//yiR26MMkovEMYbdAQwk
ssWOxhLW09XHRvXVzTHY7QoylAhkDHSReyoTdGjejzkwcmsCjzHAhaN9xFtwWvsNcJJtf6y3x73K
AifvHl/VJol+t9AhD1W17farYqU1tB96SwgdtpnVLFVj3Fsc3XP4TmXOtWZat5ol82eKQgP6Ao/q
eHOuFID5uiP75e0K5TDxgDPi+KJUUe8xfMExibTEWLqmzmRmM5Rcya0/cZO3wa6aeVhNgIlxR6Eo
WAerizizMYU4HelJ9jryQbXVAbDxkoXfuY5iC08ueuKd9Jk+VUD4aDiQwiZKN38f+u0iXZ1A0CK9
3EfuRCFr3qs+mGiPm9whE2WXMQYxLnUKVq9GtJMJZCaMW1oddWyoH3HFum3goZd4M4xbTHedY811
Esv7p2X85XA9PRD1JoLVsiyT8fLAIXQUYHlMZqod30/wYJwLZmLTkY+OCzLTuUVSGSyQD6PZe/z5
2S+FeQ==
`protect end_protected
