`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 126576)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAPydDXdC8S72zaOeXPH6GqTSLNxD/XmlXOLnyvM8WWttu+UcWAVyr+cw
OO9Grgn9f2aPyuyOZaQ9zQDoozXvzj6t1MafgAk932r2/jaQFOZPAw63mdU9IDWbfB5523Rh9uQd
CNr6E91SPNLmdXZMisfVYX3+p/lkRR36+3ptJ6RoushvjRtHzrlgAZLnpi8OL5gIJVT3pH+nTVXG
cXz3e4d3hs5fsvoNBssTA09GQ0op/34dSv529qJWT10yqVnp+wv+DvPTRV1DYvTaJaoc80aIVwhw
i4B22aX0FKLIGTyiXUZPpOGZBQeDigYARLmgk/uQrpJnk8S9aktSrFNaZikQ/rQR+yjyGcSlzNXr
9PoRcxuUxfhiNtAxpL7H5nxv8ueibbjyS5OYKxo0PgL6SVzhrSgcUPn5CJpJrXVBAc8i/ArssrSK
Cdxm9IqfQRr+mfW8pbw6XriR02v8sSj7ynmAzzxuuSy3EBHoamrfWxPEym9LBlVETlDfBaE4jQCG
tLKKYdHE7mkwqv4ASQj2MDXv7R4dQJggFc4ab0lsJncFv724rJM4nU5koInSMhd/lRNZr9iXhLrx
I9Z9eYP3PnI0oZiQ+JE3WvtO3hUDKPh7NFbozBb6T3LB9V3D7WJIXi7L2m8h7PurtYVrZU2IVvf+
WQYlVamH5A30DgHdD1r7jnxxR2hh+TYcJxx3YpRF9L2/MhTQnUoLC1V0R3DbHZQuaVrE8AH5w8Zs
cigXLil/6e6n9ILLRF7ZdaVlFGnZx5tghk9mSBuTSiYDtPSGRJpD2jeu2Zg8TIrQ3bjzRuj0Y3E1
b2SY7Zzgru3cdKyVfZbjEcYoCJmVoKQ47nNaWbSHvDscfSFXm/aIV0d2+41rJZ6yOooMThUOWYGi
n/1ufqGPgah94hpOeYg5sfkdxl8/9Qlx30Xc6Nej0sqs+8Bl5/KydtNRg2GPrsT2MGJasd/MBdFq
XaN5kMgEQyGk8PGa8HrqLB/CRu5uS+3MELlnqhCDnTfI2c64A+GWJfJFo+yChVNdmLVlBEYizJAu
nhrq/xLnChg+zOMICODqxUIgR7J17/BNVX9KZaKABQ2I7qXrtgbq4w7tt8aaniAummW8uz7JaDoB
wgW+p/AWgAlv2EYGOzzlRtAi2l4Z8P0IPN34X6sP/o+xUyZRUZe7NtoKru13JLvnsIIUweNJ/iZ+
Y/fznCWA06GcBTL7ZqQOSdIHdVQtRzIYl4fTGFIjIHPnzlushdy9qzKW8yjl1yfeFx8r4q9x3KWE
cqDAjPVVeEtjM+HbIoZmkidVhF43s6WQvL406CCwkThJeDL6wHr/wX1puLjj2hE6b9lSW7MWpacR
OPKjI/SqLAmL6QegiqG1CEyF6DRNwJovkWXWdEOtNOyfhjcVs7qnn7b2p9spx34GHF4wqDHwRtiX
t/QdVutXm1hKN/AJxeivEcMRvQNlEezViaP3s4LEX+63PdNk9Rcr5sgldMVEgZ1VfHFWFoOQlWxO
sVPHaPKztD+jDxGLwEoZkz+WhtX4RNy9TmU8t3XQjMEyISt4BX8fwR6PD+dgRAnQ/zUR5dgIn6u1
83FV4ZXf9RtWlvTw4c8uBrzMHaf2MGZpre76BpegbjAy3P3NzJdJSlLKD6aw4XfDDuPLFsd7vQLM
Z5VfQ7KSWnr1USLHCzV9wBRQ1xSBOy0vPBG99p3EItagvSeXGUcYoRzDi2rIExTEZYHoYpj5Kiut
4aw8vbKhVO10RF7irBVxiLUfOMjnq/+MOfY+w3fJUa2+nk4sJTyARUTuJ9+49LWrcAYTeIUcjGli
ZWkEchkQjkfJJCvg/C0pwYyCKVB5dwm7EhZqtmzgJeX79kReOsvg6lZzAWAmfon++tzX25tVt8Vn
954Nwldhq8txLWhoGD9UyH/o+mWRvaIl4qVLJ7zEv/iMcb28ORefyfDoK0HnUz6gy8vpXvfBUuXP
Z60B141ZxMD+1MQdyV+ALFB/Oc4zlcDX5pqDuWhFpRdegSpMDfP4MylIa7t4ROWkZ/I9IZ4OwCba
l26IDBn0MZsEJYUj8EU5OT+sLu/MgJ+kkOkPagWU/w98k9x0RVZ/vxe2DPHniQDEmhkakb6r39Yo
lmg49sKaLc/yryZ8tZlnxwIka4g/X56W1GQmyyzwLoe7/jUK45W4vl9VODjjjDNT1i/pHvnNYs9Q
aag4HqJ9a/xK/EyDWjiJoh1h8OSc3fnqA99rKny0Ll19ivv0Fnrr/1tnYxxydNFNgPS4PBWvdxZo
6f0cJd32W+Atai4rne6ynJvjdYUxyEvKaa5ntNP6SO1+LLnpDa4xLz3FeiS6t61nA/DCiFnfULTn
a/4ILG4owMAfXlqJoAJcDzOT2Py/t/65SpZ4Iji9QRYiadqZE0FEYLR8AfnR3gY32KdWAAF4cbKl
buDISp6v7W0KNbKnY7Yr0an5jtfjoYS+vMvgzedEQO3RbTIRqEdHN4Elw5bqxGGZI8wVHyn7adZw
8vF5Gb0Wifrt47XcAKmfI7CuQphfhGY885ytKyaZAI9TNFa2ivdrr6N9ZotfpymfZUm9/YqC7DIF
pcy3bYYsE3+NXyVvbUDNvm2C6hrd8ST2Wu1iUcXDFQbC4UCFHtoauu8kSL9snGtzHDJQUEsHDCVp
TBA6EPou0n5s0ALyQw2bmkfta1n6QGhdfSqejw8KTH4twgOxMzvm57AT6CiyEttaRSCbohkYZF4z
1hCisUxCDgZo4X7ulN8wTCKFxzlHp+ogyWNERRmhCyRtbhbMPbv77Q50Wx10GBHLwewzpUKI+Tkn
EW2gAdbbmVsAVPQwscuZqHzIT23PoBjgpF6b41A8ZGXpruk9Hrs+hJnrDmKFNuc3yxDSXG5Pn+J6
38TwbsCmKQfzk5r29IAO6UPcPkFu8uNH7Kki80uUv+EMnqV0SWH79+x3bBbqdIPBctb0yDV7nN2T
N9/yCLYR9jTV8fMfG6XY1vVCdhkLa8k8wsQlhf7PY/ocZYP+X4ydHLvgtVHQql4joXXQZjBOVyeb
ZewEG9AfGb4RqeFiYf7lGEr6FNxHpvR3fAsH+94zE+H20ipLDj9OrHPwg8f2MbB6WUC+LFhDB3uL
s5CRjzaoLzIyq5MwbEsBvsTIhd6eCEcUBN9n12IdXKz7MXUp9Vs44RswdeTTTUL2Tsk1hQQtiXJR
Z3t+6RMx2DsxShX5ABkFGy6MqbnQ1jtoDObn6y8gf4L90kVGxemUYqIFTV+Os2EPDjm7Oz7au7PE
5xhkb+kUFKaeKICY+3Ccjn0OPqxgcOxrXQCmgGfVrliimqtVebQ18tOgUzWe9RkzaZpO8rDNrHvs
p8jlC3bw+ciPiDbgbEcUM17iFBpbmn/7tRgryT3K+Y1EFNtOaKjCtOAJR9fyMLM5XflD2k3YKieF
uTHXu4RcsxG8yzzfwaT2UrYHzoEt0Z1AoBUaXYhmO93WWIaqzFCG1w0skol5BWgmpQntDEVV3GpT
R+8armGg/iHmzbNeM2GCHnTAp9RM6/0zsTnsw+CSZv229bz3kFs48XeLt9cZEawmxyYGySRiLqMT
RL+alzfKYy8FP96PJdMKsi7z67S0cwhVQi3ii8FN6kDFWjo1jFEx9npew8J+GrPNGLVrBoCzbCDe
+BCyDYAFN7mGGFi9/nYObUk2jkBuF3RPXYjBcNAVQ3Ee5m0loykQm/hLaIEIYIQta6A/rxilriNx
fGQ0ldh37UCjAfur7NnoLaVB6y4Nay5kgJJecr8e2X9rsjd/kObhs2zvzpiXd6I7bEBkQia0VKa6
0GxRX7VgF3OkjEOIH4a2KZZqC/LMYi2bRv0C1UsQ35yHmTFFzJvQO2wqNSUII4qCMVWYO3yLaGhQ
JA9dG+yZv5hJ1ttCd0oeNYcGDjpmYfiQvuwWIPbuJ97t3XapNU6ZwdlxMyPH9/92TUar2ohQuQ/a
QTMkwHy1Sr6S4Jgh+lKwy/FrJfSvYGzeJAgpgE5TET92Jzp9vtkx4oWcs2HTKFqa9R7P708iqUhy
Dtut9zdkGPHiSPTc/WjzrjYVn/fYv7ybKPt4KpnIPjNSVDyu5h8C7sFW7/dVnZcR4PZqM/3R7QGg
ifkDMTW5PQO9vMRxdXlkqhgAiox1coIFb7i9S92H36wkHjKSEgu6T25DztpXiXyfKtOW5CDDHTTb
b0DEN0KMcQjIfpKsEZi2gzOohuTao4Ks+6FwR5QJKgmiePYVAzLUPghNIaX8s4aO6CoxHm7Juifn
HwEVLZyGKgs3mJBurYgF/BPpJ3BapTf66jLcbv1awqCTyRivjzo1BcbW6erwA6xI+zoGI3alTP/O
b6wocksaUkEuEfh90Ikv4LeFMINO61vL0OHfUFnWeXhQlODYbCNIu0TWQ2xoTKknbGcIbM8pkkIM
xw1CS3QwXYwhlAc/QPZH3jwS/ON8O1MJ1AR3zqJQcJsG/7GXDAwF9mBTsvzWNdHtHAMzgnBgBuYH
Zkfup46WvRLq5ftGksSN0AzqikW2Bar5BDKEbjc/LgmROdgbH0oFXvo8P8SFqlkbSrXT5Q901wO2
y7F78a78vVf+mvwus/mGIhtOYP+3KJ3p++tMfhW9miM9pWbqfOfZsnDT6b/iicEJI/d3bO6fTds9
LdvMq0h5DGHgArffQysh5ustmVKN3iahzQdeRi0jVj2I8joORhv0RBvtFoc8xx2XeJ6i0ficec5J
+dseHVRu+8ds/qepbnT2vA3t6IXZ+6mBf8U3GDb8h878ss63A4/N19jdqk+sxBUAmmslRIil8ayS
gkfflsJLl9106jwj8+vL8B4vzs5Mrx/tDRfMzFaK8xlu6KMMACjz1arJcrJsZ5l6Ymrf0vVMLcnX
cVZlOAwFQrHpnaqnoDZHLeKxbd1zrx76xCS1/g2zS8ezNh5D8ROqpM98I97B/xeaTn38470Axl2x
q5N4GtjNAH371bSFiFBfq8oQOWzRDQ5p+FqSvy7ziJwD9kA9oXwRTtY/dDe3G/gijJDGapKwULhW
c2FT6AseXCcyMQJFj3SkdiPp6Hg+DTNWRobX24aHM0w2JTeO0VOVPAC5FCFAk9KZiRD3y2Rkhbs7
9d+pbiEzNsKkFVThwbnDTCLarn1XWxYZmDOVcykvthWQY+XgS3i2cdHATLYeuk1vtkReqXt3Tj+v
QUIL5csmb08LMmxmYYPrkFfD7U8nBlom8GxliFuM0R6n9oQ8/1T/6yw5EMqzPWwMG+T/G4uWI7k6
G5/mpZ9/0Rxr28T7xxcLki0yt2rQ+vCyjA8JYUsrFJp2xOiqnz3hmk1ZWp6BKy3mj2EO+x33QDrU
zvrUXXBw5AUWxXgoUOOBsMiNMbFGFU1lPxGI7nKoNHOi6/k1AnQQj5j6DH+NBicwtDu5nRIntILN
4ydiqFt288mVDu+G4RkxaWhhhHG0a4oHykb/PpP11nZGPYsOQ14o6McJB1gjqkO8Yn0cWhu3fnhl
BWeKY16ocsTrSkYDghUOSen0imWBj7prLCpnbcPe5P0KGBsAo+yDChKuFT/zfYxgmIZiZn+b7jNl
dKkfIwUM6z78H/flev2UNVmHGinIxj/5rx3C79iaxqVDq9CXapJUHtKnx+CmHVleqZFd3Ym274H1
0ZemOUV1geQs51Hk/ufez0MZZSnSVOoStUjEaJKm0Aj6eY7phOjGOOKXATAAtdJhGO1cnI3YHNz0
DU4iqhGtu8rYdIJUHp7RkU5BfdQaYkJSc4FSnj+XOtOetCCTZ4bUAlN22XB6Y8WSkiIYx8J/Kb+5
dXLt+g3qfKgwh4BLRpNercQF6qz0LQQxrcsrHIyKadYMtP8nJqXjwvp4MLZ0ZnNZZ9NljMV86mWR
mAT6DjtIwJzUr6NAsT16sSlZl4HNGduNSyouKgECwMASxyVOEQ4L1L0qTRbZvrbEDTnB8BY0VmNT
DZ7wkT6/4gNYBIc/sbd8W5OYAanSC4zVbz5Ol41wUPE8qPeIWjgQ8U0o9wtbhErUZY687BhM+/TL
dJq8NlOu1Bco3iFPHRTKgey55ZW/qrLozwCUY2JzMQs7GfFf5E5x9ErcL2LwNsfqF71dexCGw65T
tgFsTTFSoEylidIjEMIKdjyPsvzqYagVDOfqTIyJCMhvDqxGgBcvWwl6Dhk//Qj0j5KMEBr3eEq7
kTTNjAm5VEMJnkF6tpZkCt4ftH6Awgt/3AmlkdTORnrTqJ1yXwbtPPETzAHX6V8Okesosjoazz5E
iouMUSdkNsxV1xkuFDu46MCVa7ui1a+dsxhVYWnE+u0eHmR6Pfh8ILYO8iPsmgJTY4vMoDcSOZfN
ZGbtQjZb+JK/UU15czBVSXzXeRaLOi5S8+eUmy4Aqre7AY1o+vzaw29ZczpOiP4K8eqeS1d4/TAi
+umHZjCXrMQqXY2y3ZXHmqir3/3PU5WUyDpWF9AZ5UHh8csxpaf+uH2Nk7m2ugNiwXytxWWeGBcR
UfR+o0Po0CvvYPv+1sR0JYDEDLzj19znYJnOj/WmHT725t9CoeqGxX7Yi7P2Z9r05L0Tf+gEmiLw
exgO3HxkBxiq2OG+msvg/08+L6PoWYk2GdsC2dvpXV5HP4qYDe5uqB0XOd0rEWCh/fVa4RDyU+is
hjhAEw4l2kk/4h/H/UI77J8esDiAtQoTRTWIGhmiQDMPVJsYEI+bE6HYt4vlFRHLCOZHg/IAAAsD
l4lmDW2fF8gFAP9ACyLKexuM/jPwxKRo3T5bD2XhdMwKcGYDOHKkZCXGR116vtiwNbmDnszW/n4v
Kmuh4s8N1FoR9MCbA6tgtCOLLI00FOcIApiGHKkoiYsJApVsxp2/bRnZchYx2RAgpXotUmlIsf59
SPkG9JYdgCt98OjJ2bBPJM6iCj/AUmv6M9xNCvRNpW1nVcuC5ChY5Zoup5WM/kxP3iBQHTZWTPsK
qIJZ1OgPZgVRbPKSRtyR9RnFKexS4gxwP32EiNgGJVdHCozDAfFiA6Tzr7g7I/+G4EOrvrKXK1q3
ykydDq8u3TrQy9Yq5vpK4YBwJ+hz9ugGqJiMhJBp+bNJv560vL0Mb0LUVBsUsw6qTPPazOSqQJBv
12Xi7VDZYOpwQPA6HQyEtn5qlpD1AflUJzWpTVzEBm2s04ieFD+GuvZ7cusfpQfjni8FzwsEmI2P
moRXkDnUwyKBvxaRoK4nHdLpz97XxpmWaNztudRurb1K4mLoVxK1SNzIOgvsiksCvHvoa/Des7/b
yaIqxCQwdX3+IitfO8N85jIi+NCh6Pb4tfAFzUwQI8+MDXPz+eRO6e39sp+yiXERCZ62IB9MOltC
MZsJ/g7VklG+Y8K6jlqLN2YLv/j54zsVIf7eJCV/0sfYGV62Ol0ZZ8H/jOgqifGvpxMuzREK5bM5
FaN6jpJs9bis3gH329qFjOp/AftiyqzvQia7xaWTPIGFaQVdnLm/wsJe8dXLXkJVzXi1WeHZADxw
t0HVmXTfg+gDPQyo8D8UcP8OBcjEVGahy27arqaGsefq10Qs7hsd8TLIvHv7pA+WaQwsYQCD4bJS
zqDbM/Jw58mJ+VimRvJWiyir2hqN16/Y5LIrA3jt8q015sszulqR085jzR/uEukPWBsc34pestD6
hJ71KzP90MUqMxZIWAAtobRPZSjf4DDO9kPHgtuXi5sxbmA+taWF8KyScufsVIWP7GM9q+Z0q5zE
TtNRrwbSpWBzz6/Ieay2ZnRlixHHdNX1b5teM0tXO/fF0/Kqoa1jAzD+dxhacf4hTmghG+ypIdEB
BVpHLn5BlyS9/OxzI+nGHwHyJa4ulAZTjzOjyfAXB040sDvyGatxWgpiZyZS1COwoCWU47JjE7Kx
+bDs+4qg7aizeP9Jg1/rrMjUqfujsRwVCz5DVMWo6TexY6idxHjC8wHWVntLtvrji/ffqvTuMZHu
xCC/8yzvrV2O/2sc2K8loqV6ruWHtoMdRZZUVI+SIu42uOlZtdnkw53de90gZxdOyLzhQ+vgx7tC
36zy/LJ2sVm3laM0RJdDlUSJX+6g2nSGlrAxHQB5uDjG+agR2dsxF+Vy4qQL8e8QY26oLlG1ZDMl
bcJ9XSes//kDf7aGEOE30vxcJkUc+Ak/SEEMCgFimWSNCN+l1ExPc76probrhiAaJUWh+ZkhaLY7
9gcrSJ9NdF0h57l92DPLOI9eDkMLSSQas+ThSH+Th4okDcBFf2TIMoG5ojnTlsegefYLbC6Jj7h6
gIMSIMLgkKM5TTlOclpipUYlyWhfzqxB3D8ldHUDXILrR9193hEeUUjp1Rvzcjb3J6iX6jBMnZNs
U+A0/yyQXT6fA0fkJl/yk28ksLk2FwxmKB2lzSNc2rs8hzMfOJylJcO0k7eKmFqb2wuLS3v/p+xp
HWbgZoftxfYDmVOqOgLa9DUR3rm7u4V6kWzZOIIpe6U74YfHr27N3YQoqy8DhXMj/WNVy3J7UyNz
hg4b5Z0kG/hW8QTSHeY4FIMNx63GizQpXdX5TvMRojvHC7otuHM3Egpx7xabiqqzGjRVYRVoJt86
RGf7BV7VZtDFJxfeH0SZa4NCoe0CXnnRSCtpmAwVTaRCs4GYpi9pdN2gnNxNTCxeRtzdtX2hGVw/
tV3Jflz+Su+268rv6nHXdhTj6GrlnTE6tOcP0heGu1mGq4i0ePIqhLWxAHX1CZ8eAQiXsLE8voWB
/1NJpVnmF+6tGly9gGfvkjsYAHHXqKMIvdbCeEZ1QPIwfeJTZkrjb0Qt2yWxPk3B903LY4PF9MoP
xBeDwMl37lF3Kt+0bi4MNnb6rnOa9bcac/ZyQMq5F8/Py2BB6TAGIxxrJE/mmsPrC72hPtVmP22l
bWwKa6DqYB4TxvHdVXa+zoaPILSJ2Gv8q4sDBnnGCOlHwzSx+XbA1oxkMXsYl2WAHANPI1TlvDfy
vcBjJAZmq3yke9t2bIjTDr74L7tfK7W6yCgcmD3bGW2khpPAXqf5kc7ROQicJ+1HdErkBH/k3jGJ
Ga5R9s7RDjrNlrhQoEiFVoVWjbtfMecvIVm373eIidtLPG0gzf1yP1P2kHVjCrIfGr3ZVVjsfVyM
OjF1NVrtG0zDHH2plWyoVkQORijvzIKMtyOzR53GJDrFIl0nlRAqqgLtmAiN0SYmHuEF1q62IaSe
dVymG7RM58OXCX3d5zrGC5t5FEBlsvX8BLh2QuaAYDG0ggIXKcjtwQJte+xBl3mXJkQ7FbK3bLEr
46FrjiNbkM9lsU/O4Ek99NWnxyh/1Zi7ZnDD5VrxlZL66wf4rieXkqwZ0U5PXfw/OwFZURWlahoQ
sx6U1nEoQKdn720+19bMkY5NDv33lD/9Y+PEPITGk3k3JzoR5MWlAWd4TjhgrzQpX7F0EQpAusT9
aXW2x0HojBD+0umf3i4BiNoHi+7oZX7f+ODkFCwzjYiYsHdfGzOoVK+CTJmJBOiT8qoPAvHk6qAS
aqiwaOQT+sXgJlD8nnsO0DNPLUaVg8r+yjC0vw1zBemzh58PQan0VKHrs6/YOFtkey9Oyjq/6OJn
l9tBelfxfJJ+q4i2BuD8dEP4qeYeLRyz1MNbO1BsTLGWBikVfXVUlymNto/Pir6tGh/RtfiKTAeL
f/L917SGEzN4KgccU/Tg3On1QW9oBNXuu4dsD0IVxQSkdy7oRsphdlJ6DsJWT8VHlXRKYGLy0wYX
XMgfFhcP/d46YRzZ5emJYA9q1OuiIbcDuomvy7wIyf47fAxdmgi83z768KbWxFMHkcsIwQjPmOMr
qYvPuk1hj7B53zvHzNKhdzqCt5wlqOkl1UMWkJw/2l6nJ3Jio4HocX4qH3ZG/zuFR7ahRpdVMOqE
c1vNGP1U2lT8rsP1tn9mcth88WILDp+o2A6Xh3ncHu4w0s3vwJ1b/F9qth+HQDvT3D9mXMOiNJe2
UzVJAaaaNxzZ1kPWXdui4lkhsvW0jUiSsfcytf3KcdUUlTyk9AjQWIbB/7udSYgx6q/1FY1uwNSF
LlpnXZ+fUQ0esVoyYzRmN2h/LLfEAAmRs2dHuYRHGc8+qskhDTtCZ/5T+AodSfKFxDnyuS0GlYag
i1gaMdKA6RYghX/iqTNZgqEWMcE94yQIXkpT5jTNj3/bAQuAuKYHUYOFZk/hoKQ7i340zk6fufg/
c/v4yfXgwnv5Irc4LF9IQd4dVLv5QlqqrsmfLTm4ce6OloA3MALgFAcCKSH7QI2iyANMoe9VLQuO
sjzi3IEPVgA9JwRjRaCzRTiqAdyxF4IGYMqxKmri7RDCSVIO5lNLtEkWzPbzsOv5fyyoD1HYIppa
gBbYY1vbBiqCmsP5CKUgvW3nG1EZu5wSawKkThXfepjra+41RPNyD5459+9/xYR+7MtOmk2vFf40
PqiLSIkJLQz/77UPgeeR8XoIulZOQnXrmY9iLWpLvbgGpyCUmpO1BfQADfTlbRVbL+7Jek6CdQtx
TeT9OJMUf+xF2vT8DFNBgc0Uc209FvwyE9q+Okdvc5lFEJPDZRnF1wb9J60v6TxrD3mhGi3NB5xl
kXJfllf2ve6eEays3khvtM4mqbetRjOCTQ1b/GModhJQWx332zFD9duwJGoTvVj4mf7qcLthJWSH
qFr0GORv/v9kWWzcSEiRhed1HpIdKqy29KaM5Z9qtwvmADCQvRObc/v9bIAy2D7z+sFVNvZp9mjw
FfQChr/sIXuLhQ4S7nWh/NvBD4CXaxo7ZIUk4A6KrVFepfdwZnXECbwW9BKs45PaCRtTBVs8gGjW
L1yTmYl+DcNHz8/LLEViMUaIk9ti2Wk4YIooyGp0X5XaUBb/CugSxF/qe2eqluqGcPYR7LFX9D2z
TtMChpZ7Bx+WgQ6wGeixJJzebF2LZVWkn3k0IR+kF3Qygy0Nd0H0LRUtSU7k+vB82kYfcmo501Ck
CJf3JDLuNz0DKMK9I3zLhZ5wJYWoCvgBBVetQwjKvG/WRJe1XQypp5YLQKD2amYmdugwDJAAPS+J
vrvQpJzJ8rhtPhBW4XSHAqYZmxFreqExA/6C0rWGdLNztEJYnyGPJk5lfVfCNdqTwlnUcGity+JF
/h0IQE38TKsiZx1lfudBF9BghLfC7H8ygqaGj2m01A//7slBgEfHBrcrXTWZhVcNNzXHOisKrtM2
V8FIKGJ2X+suAFQL6CeNH67SvvyGfefdM9HWnmXwFHP9Y+gqBsOF+DFwcvQLPPEWSotYKthN2zHL
JBhPFmy454k+AUhMlXU+bx2BouF/JgEmwjiitsS8JAfVlkuWcl1qUoitR4ZEWSe29mNUD0KwYf3g
H+of+CWxD0aoYb0OkztqYUufl52PyePx+hBKaz06WDw4+X2PdTSC4GbTyimIiKadex5KPLUiHaK0
15x8WaYcc0drjvUZ+ARZ5WY/riESo20RKMfcFqt3bzf30cNc1X1ycMLu0l6JeN94WQxIqG9yDDN/
F2F1ilfQ7HYfJWps6DiXhrhoy1inMKVPSeO9qUXTbmdBm3tA2NqMRUTNLv2e6yzWORo0d3UlxUtw
MzjfLw3CHL2zAqERleSouOQppK1DplwHA9CUrO0Zuq3GRqghWBOauuAA7aKer7FOC1r7CkNufpqR
z+WJSkBQ46I30bEiBR1o6SW8nb4ThbtC9patQakChWXyN0J2RS7rSU+3Zy07f/E1XR5hz1hiUOMB
thsNqdu5uB1lw0XD9TMQRCsh9QoVaLjGCFQydU7zRF032PZtNBiyQeZj1FcIeTotJob+k+dT2DRQ
vfQmyKKCRhhE//Wbk/q2h99MSwCAB3C1lIRuNQSBkkmKqwPYfUOdEw3sszlnxauB5Hxmz+gFhFfL
M48TiIkYqeYqRrCIw/l8MWViFwPf0lpro0WsJMXjb/lZzNpuF0jNIBYhffK8Ijk7YHFyYF3hB3rB
g8FEw+tIuN0QUxb1nhAcJ4iZijGkc/oKybeZuKSu12FDn6J3fxxXMNwVQmH3PRuyKih0coYELy+G
NmDD157aQe6QGQSVD433ZsYdDK/G+278B1pZuBHyZJSbZC90qUi9v2Tjr0llcct/g5hVNV3NtrX8
bgdybjt+rhV3cNJgQZ/4E9FtesmwvTPYnUQbrTktSCSnTiPHgawgRe3ew6MiRFDjEWrbbcuu+Tw9
qOcutC7pEF5d4M4O/IcceMNP8nkWclOooPSshKsTMeMo2/iIsO66OpDG7Kh5YmS0M5BLJ/h88jTR
gCzWzp0DVEGvORlgM1PIZKaArHDR5JyPr1MBileHPopvixcMOFnc8qdGqbBK3GsrHhJIOGGuH7SS
OKaNTVf3+PtIaASktWe0SFf8E/ZRhqpBUWeo7nrCGd8l7xDUTq1LnwBnI0qPaj8HE5vLAIZddnpZ
4fJ2SJlQEshI25TpgjiyVo+7RHsYTqZqVcu+/arU8ytg8XMJxzevfooTItA624P2dT2AtIgXZZ+C
OB5I6rtjehWgot9GhTGNJ2efwYWDARfA5+zzuwNPEjdn2/+1f3I4tjQLgwe5aGacCJFAkKUOfXYf
KYs43vV+cQvCgq+8GncdUimR494BkxfYaMTL2LrBl+Qv2U7yHDPwMF/XkI+SnT5hDllreJj0fEn7
9DBH0MdA9j5lIf8OryYl+mw9Z3Ke+2QmNeo8WTOJYQTyDOvj8K81A1XxttLfz1A7cbcq3tYwIu9c
E2/9hS+tCDGZaOz3kw4IKwlvTWxDRtCO+Q2ZVxX1NHfWPpWNCqf9FAYJQwITaRGG05eptYxUm3Ha
G6DucLHAl2dxLtxAgnkNirmuTR+WeNjK9eShyH++1Ye85UvOKLE6bArVXbZd2yEDHHjNGbyIrXPu
ZU9tqYYWyf3VkySDt56JC6nfIx/8xjDYNHdlmyiluJio+YIe4NTU2Fkun4S57dS60DH6WxhQUcKd
EHZO6oxMXgBwOdV76iy5hQN5Al9a3onMFLbxcyz9DvDg+dAdukMsl737wvBdIjb2TPHwOb+vSVIH
OmpXYyJTNnOmojDFp+4WcOlZw7twX5BTMKeBeXe2r8ik8Pe+vLDlHQfD12KKuIgPk8RzkllRRp8T
H3l7+zrC5gNgEzTOSqf113UX4uCp2DjQTlumGvewIUJVF4uafwdT3weCg/h7nZm5bmAFlthU51gU
MgEPUd/K3Af1blbdVqbdZvEIxfS9kDXWeqoGW5cALZMkta4GSqlK45yvO7zoOLEAd6WO8PQSgOnb
1EfisVS+TEkPOL+x8hp2+N5PMUqMVSOo1++WmT5+blSLHS1MX7cQu1MTeNVjbKgg+pPOi132XF2H
XJfU26eF44VFmRlJS1QYjHh5hCaXW83+cAKSSHAl7Zy+vy3w5gtViw4TUD9wgU3wKvQ25YxL99FI
YybfADUHlVFb8ekradyZaAwFAz5EETZO4m1zTWo0uCxS5DJk2y+dhErxmH5YaDi3kZbuyUcMYq9b
lTKcDsDdBi8UphnUGj04UvFGfTnGeRHIb2d7s7pOIYUc/b5L9dKTer6qSgjahYN6PvVxyDenJrAq
6RPjkMVOsFDW19D1T14UlzbZiggA1r1wVJWg46I3EWxnN/dUFswJAOppxjHoMBmA3A6sHqniJ5jj
ay2sThVtyZwK4p8pTElV2FWP0A44c542QpxuOQUdDJmkjNst1JyjDsvwY+sAh3Sa5YTf+raMWnVY
5MqodCKtcy9mPHiMbYz3q1eOtPWJBrqD5+1MebOEJMNvqNJiA+ydpNUHKnqyIhXSC2s1d5zF6ySY
73h3PJay/r4Fs78F1Plb5NTCPHd/U33Gljr7vzVGbP5kQhCqLNCv3x2QUDOc08NeopVfNqPyFcfD
P8tI3Bcbs1VmGhPtzckKqGFm6ewlbumQz60EcF3jEjcZQbfuvuCw5+pvy4DstcmOfvzq5oJEfJkv
f7FBN9eh5Ws+eEVLuvYSXJ5q/IXbp+A2xW+HsFiNJHZmx+2EfEuaKu1xMqOHALhOpbaYiNQiLrgI
P1a5d1Yg/mdIWNaIeWg/MdT+7hNkDa4JDKsOjRnncF/VDZbY2vTSCTpPhOHuo+xqK5t3tPe3+7e0
5mkdq3vDRgT75epOqs3oY3Pdn44A4ZhlUYbiDlJK6YsBH7mKSoiF8NhFt2SenfYLW4Yjt0cEikIQ
0qy1Ug0W+kjuu1zxWrxBcU/D2UJ7Xr5Sc3xPdblW/etD0llR0Mh3OIYcBqzz4fhZob3PM+aqFvGl
TXMO6uuHZ3Ky4kCf9EXGGNyXCjaVkVxxjO6aQxU5uWp4wscij+QPeLPC19FyvlhMEKHSGlyxF2sR
afv0BjP8Nf+zFf2Hz9MfQFIC8CaFp2rZtI9zmAFq2ejRqVXqnStetZ3M9NoiA51GzW/ztONADKIn
oa9C58vPsepRj9TUR6D2bTf8Mr41cPEZ9kaEibsEqPjk2IuCJL06k13t69D0cHyosIPkjWKjxX8f
nnAUt1w0JLNG9PY3T68R/6U9RLUnN+dmmtE7YiCOQsBtKf6GhbuJoELLzH7Sh4JRh/ywzPMteIFH
aRtlzfStw9yAsuKVbqdWoXBd+rulfnz0NSzZW3qRdpmx+xxxvrXXHDCVxMxrE4ATMPf0O9KGNbqj
9IKp8usbZYykgXnisFd7iZwGr/lLA9HQdS7zy8hiOkH/n+wsreTVKpOnW0GTohVPRdOFHrXGTRgK
oe2kIBEDHiXpQOAsWkMbVzinbZ6LQ54MYoO96tbtljYpq29eW5vjYJ8pEPmCBJ6IrhZDR8++ZT8U
TYbMEQFQREns0ZEoRBPQXl7MQJ3/dA0gXGUk6KUHTR/FSL6accbD7lwUb/YUFQmToACuVu7sdkXY
0nOxMp/eSkgwqWTqmjti3Lw94m5EGPKgpQBuN2T3jhQlJJpqvbYomCzrpGtBjIaAiz9Zfa+YEG/u
vL3pkDGiggziHvAR6BYu/xl1tvzTNcJVBQe0Iv9TcsvAiZpBUZh5Cs4MzOTkEz2uPxxixGHKM9uD
8HDypCdyEH/dbUKd5OTg6HILgnktueQapLVa9C+3lzrI5THiOPQkTTuZbQ6AnP5oP7KGHFJg7eYS
Pk2jSr0dWtZHRfKumI3QdMDP/Lv6ECbjQkperFELFD4D9wmTzVrl116y7Q+D82ETKZ5OeoVSP7zv
ZXJiLhr2OI/171F/hMRTb30qEirIcLFfFX2BlAP8I7DuRmCQ3wcD7KBPC/+WjZzUt9vDyqwXmd0p
z5I4XJB3z2bXyEjrIsliPPweYqRVgVEQ1dnKWIjiJEFmnLTOcPzQeZlVglpQGjUFrOHHQUcRWVji
leY+g0Eqx7rpt+7I7SOvUI9zqaivAanN/Svx5PPxyrvip17UI676R5SXzkM/LojTp/mJsDggh5If
Q8zFB18gAcWvSAHJbreq1abo1FG9GYm7pWE6/x2EVTZnRQqDm/NA3C4W2/oB/uNHw4TaN+TOfoab
zq21hLu7j2YKPoEjO/GoulE08SV0YxufV1iQJsuMbAmS8VYaVsDUJtQa85V+xVjkWOsGsgUCR+ML
+t0smGAus2X79MBMs9JPwYYeuFv4kcJ+hsGDPWeAidUdBCv9JrHbmQQal7d7TGXBi5lvpNkLJbmw
gDrVmocbkA2IwYGCmFkVSg8m3G8fVrEZyphZAObqmVnww9iRQqUaBv7FlSLDHEijgjLyJM5ZsDSY
hwL0rfr3rwOB9V/zsUSu+M7WyV3JpgZQw5QEuvWy5AfDZ6rjF0K2lJhQrBJLKjPhRkGaDCTPnNZz
dMT5eOydYAUu02cTIoq+egTB1BFBbVVcY7Mg5Ci3AKI0TfoNBCeY6NqN/bIMbPgkVSNxX2IH3YgF
j6Q2m7pKKd5xMUwN8cStt8gMwu+o4fbJ5+0m8OOoMbHO3uxS0DgLEHjMX+j1dE0ADq14l3gsdAwx
csCkm3q1EeTaQB41myn/xgAiFMaila6Kz2VuZZOfBkHTmFk066rODD/UjbGJUXl4p+0W4VSG3c0q
iXLv4WslVis2sl0Us7+6qAhv1zF6BoGf/l55wha7Vt5+JUDbYdwXA2LMM/PyRZwjzP/X4DuGLZnE
jAOX1R2ydFqV6hkuevg92Jyv0NupPJhUe17hdE7zwTgsVkXzDhARz53KKe+k0AKmJfB4DIjtv2PS
pj9dCJO2dTnK0ugfn1TanOJMtjmMOOPavaFjdrUcbVbtJAjCqSSSgkpX49Y4Mb/f71Gza7CHOvJf
1R1t56gKZhcFcO/YwEwStmFLIF7ooRPAIV0wHgdAhASpfZDzgpgjPJBIchnzTTbezrWsMWggmI6Z
tKliY2o8YLMR6B/TAqT/3OO4hv/fLrELFJsd4ItYQ1/OKiyCt5hBebxx8iBASVYaAkRcq8D5Pk/5
bQqAdRrB4beVpum5TNHh/PvAOV8qzhy7jWO+efbI6Y0+kbXuVd7KMp56/GtGdASU7XfTohE48Yk9
I4sJ8ttavedRmNXd4VJCt4C5zIYrL7ct7lW3QO3VBYZcwfhDDR6m2KBZh68R9ZtaKpoXdt/4lGDa
cDxb3lGGod9fSBNdOiJgslTnMaxknVaVdvY3mBrdZXSIYRpPhoFCO+GN33F5cYumnzjXh1lzCcAu
CC2Mp9g9X/F8zbJmvDCl0qqD8I1NiKK45KfcrMQpaUrpHRHFpQ9Ha3OmhUnhDi4tVHNw0SALQmfv
/ZZQGO2s/n+mwqeg4oFa7/GtjuQV92QCCpURRq/Fe9XMe03p4WMq1n2TxDiPNO/V+XZMZkO5vsfh
dCUOuJd2pKFVfmLqIYDE5B9cBSiDxQ5w1jUCJn3HOZJf20bf1NZx6x9oYqyoNO4YzaVtaSkRi78Z
k9EDGc3QDPMMtcabnstQtXBZS10s/sP1aFrvBrL5OLmdNM/V/g2rbqIRRQZj7Uv4piUjFg6+u9kP
SPv4MaiW3/80SBVTxRUPhVt0/2sR3nza45GdZJiYjP4kWp0b6bnwc1cLEPZOoNo9+IYHetBYP0Jh
xyed5my2gbebeE3m4RiK+PoENPHFAO6/jAkV+Mxt1FSOQRgUEh+q7TJahcubi13AYkFR2NjY7IMU
jWgfxMsTOEjRggCXIEAmcUQoYDWS39aOQFTBlLYEBUR6gTx671u6jGz1IjhqE/jI+kTsVAW/+Tll
DZPS1mzONfd0jGiZX/LuixhvAmSSOhAj66x/cCQKJTsGUiT1akqSkYv3msJbJw4tWDqurzsLU1RZ
Q2h+wNbg2MVjnCzASii0eWE9s68liwdFLYVMLyNT/Wlk+RS5XlZ1Q+IxHqNPODHLm6lRO5EOogrV
WWRcQO2KgXBKrexFBIX3e9yR3LeS7A3j2Ray4vmw4gWtmcd06VugOrM3BBU8UhAq/kfhlsbqJXf/
y7FC9l9YSKKMPWDf6ONY9AdAxTV2bk0Cbxmlw/J47+hD6X2ach7i1ZXVP0Lx7ivAF69cMMR2jYmr
cRaHvHAAIRkQXdu3RjUQyg5xxBBNLu4kvVloRYtswhWf+gKEtlR09b/BRt2/0U/2c62hafRdG7Qc
82yvnSObBo+JZIvdSuco2PocuRYdhPH6WalAdbvfDoFklUnO0vFct1jPPPRvThZlGTVc8KlTg4uD
i/oojo1Ddceh7wfoeBODCxG3cquo3SFhnSHHNfhnSMO/jyj/Sxd4F7tZJhCzF6I5byDuAScjHVdo
dfAuGoU5zQ9wWCAaAdYLdvcLR2Sb3ex/S/yhDNwLXFdVa7PushmRlkeNeJ3aQPjeu9hsu7WY4g1t
JcxvP4971mcWdam7zQ2h1GJbdPyYy8NgMepcj+5zLJJzc9oReVuBY669W7CmJ41xCcrkp/v3QgF9
yRGrP5nPn7PHALfjr5CXyGDEak9F3mGOLk92c4b8n62QS0fILKFFviSBFPGyt4ArMF1kA4yeUKdV
FARWYxBN4r2f7f7IfmynKyhCDdw3W/VHWYzaND5ErrgXDrhIwGxHPHUqKbXLVCYM9hrez6+VhF9z
iIlZZErpkZfK0QLUCOb0VL9jzUiqlG1bXplX5GQPmst0fMnU/WRfQ1mk5V/9Wly4CG8pufaP7qqi
T/A7JY4GkBcY0klYD2Dj43ehQFaYOzmbFbXTKjK6ELZQBE7yrhTHYfnM/OvQdakyiNs7kNoOIAxS
eO1mSjupxiRG9B68/oznJje4A9OUW+WwcgzHTC27kL+z1FSd9agyybx4W0N341AprixwhSMvWUe0
8ZleUgdOMIacG8Sgs/XVqW0GTJ3Gb7R9CKhNcSPCznoLsPy4w43Y9BZKv7dI8tIa2Mwf4nlXUddn
Ianjd10nR61Q4sN8RZmDZgO3WWo2FCYnU6EsjOqEl9kwLwQjZ7wxxAlKeqxxFqsJArvDfy5Iiqzu
eAMxxLmtlj8k+7tmuBH+VVRoxaDFZYwXdJxhqZoPZ583qnfG38GSgSu1RH4ysUr/CLhN39pxht9I
nP3DXEUF6D3CE7SW4kE8qCsB6wn3W7i3XoWD4NCekv4gwGBdvKRyX6Y7f5lETBczlNgElD7REfte
uCGbzeNU9/xx5Z/lAKuMkbBeJgKYsV0a9xSByIIF+4TFHYcw1vfCZCRFM23sqQQZWrDgs9OTib2H
s3KGcTdHQPU16hK9CrVBEynumPuVnC5uZ8ZGV0dE1WTvU0HmuAD+O7OkTcOa+EUtPM0M/vUD3eJw
FUQsY8wR8mho/vVL+SYq+pzXOramSjaBd1hoP37caAIwjvONFooghJUObN6foODCUW/LnwbUeIk1
TVcWWy65ihLps/SSzq1/lAkRMnRwBW0nM1ejyaV2fhQ12S8rfORfMzVKVlOZeSjUBGLhyxY70akx
iEM/b1Aqny0OqfLnFeRa9KO21VffSKgk+Womt77KAQTkpBBVNrcEb+HF25Pg13zGDXwH+cjXBNEB
hYy6Nkr+vnMb0MLKvaMQIyWkBt7zsfnrIH7hXGGhNz5oZFc8Usd5IJT9/JYGWEehyrJvfB/Syz1l
a3es2nG+EAoW931pdcNslY7lmj4Zp4xsT+93IRfUr7570WwwFCO6IXR0+SVHZyUex+cDuTRVYgnU
Qi83zsy6vUCLEDdgrWMG+GgwqXRP15+wPZCq+6wcZGu5h7R5UIOaVloEwQwGFXOqaUQmd5Gn4F+I
7GzeuTjkKfLEaKVa2ZC3go2KsHzC2Id0gD8YhAQasw1c+Xfl6lx2hM+YbU8YaK+EibGAKH5V7voK
Q4lq/FFbGaIu0fNifbmc8nky6CgZrbmnUO23cX2NlU0uYte8ErJ4fBg6B1jFMcP8WcUAJvmD/93c
DplpwIGixixGC223O/Xehd/BG/u074NJcAXkzLsPKpmUlX07006dYf64UUqoDI+jEEpd5ZDoNbED
DwPMGqunvz7YX7tjSfw2uCSHXA0rjPGcE7Ppgn3Ufpif3Vm9i8pxFsq7PI//SRmKCn9akb3kC8+1
iJt5txjP9fKxzyKJxCwG+GZGWUeeFqPiSIWBJ1GDI87acqQ3+dH4XKnouJDaqIOTIl3XYaMIdJyw
QRPn9LmzPE654+Qgs5cG3FtRiR+hz4f5PiLIjQjQAv0i87kMz21Vq3j1PiKnz2QQgYnTnpj4c01R
ZQNsgdPWibJfPttG5AUlF7eBJD5MniL8rUWA5A81kWjOY2zZArafHHZ90aYyOtaDeOvx+U4nx1As
WiLGNI9VY/YrZOrCQf64HpDrmLkTZYLr8MyAMp5DF+nISOgTcpqZVSskL+BLrlbcaKuZQPb8Jqva
INJPMXEFN/hBpU7vLJMoq+guFEvYX4yskaKGtVvY3SWgEwMmE++6hEbsmnAwRV6rgchCxuDVf0QP
PZk5S0lxmeN28AdHiJF6d/doECpH4BkJqjR97XquxwuLmHxiev+OP92Pah3N6P5Wm5WQp/oewkBR
/Mz++G8TpwAIGinfJfpicg8J+9OhG2nvcppjeQfQwMk5ByCwT8GOvDg36/G2fECwMIb90lLvDWxs
AeKYwKMqWt5ywou0SaeFO1zt/ZDBs1XtcMB1RWS4vSs9GfLg8KUTBVrwYzDePerfhjx+qVj//VNP
T2b8t4wOevxbMyLOTKUu6KNnhWK7Q7vC+PjFf0T+ch6nh7A8rBZ8LtAS20SgSw/JRkjzJeIyZJIM
Uq0bq/bZ5nHRdihqbilZHdnRY8lbI3P06LqqyNQEBkkc5sJnBnbR6B3rbYoTr/OnEW4HP5OG0Non
MO4kR9QLSbTMwqI2ige4FQSgZSHomRZtgMyKyoYapv1tAzcfkaUG0RvO1yKcZBql4flIEoLi1s7G
7VHAOtDRHxJNq6WyIH2bXc0xPOitKjy3iK3GxRlh8bya72ENW/ejsWFYa6uY49UhK6ijdRwMb4O1
Fc66jTc6PO1RGkWLVLFQqh22zd+vYuQ9B+LaI1eOFByQqrKu8Ca6I3a/7qSFFlvDtr+koduBKlA6
KxyXoDHPdbYCzpKHzbvpOs6u6UUPPnBfTvKueK0aTbdJK23OiWTYhnYZAoJIO4WpERbPQxJz+hNl
BLpmgUpscRs1ST9wIg9D6c19803J62AAumL0B+pB12rdjWDuJbiV4fJBOUhvPmHv1lFD7kMZBylk
5sjL9cvyn5KKvzuqJjd08vVRf9tjoZQPenIYos2XKnewsCOzHiwnOsP+pc01vaDh6W9z3wVm5zaY
oxWp+zEqPyD0BQ1LW1n8VnQTzlVF8szZBbkokS+g4F4tkpLJJIVG9QFMcKe8lawZJek/rTr9zhPo
N49zS1okCYHKWmInbQ5+NNIWbtPTECnmDOiZDFD11igJ6KpJEO8lOu1WSBbthVE3QLDDpoq6OWcY
R0kd9y6+NUgQQNjodEzqN0bV/APG59UxIO7i2PdQTH+79clWzW+JOTZXf7oJu8+9ioEErszwC2cw
Fka+WMXB4NbQfKMRb17KP04LtCuD7e5Pr3d36HVNRHHCWP2yiu+ptU4OCJMP/YyK+oRcFtj/BXB0
Ot09A5QJBFUn+OoClCrJZcWDJdsb6KH9UgVAQahubEdpKofS9ahHwQgbCUCdvoVbwo/+W5ms/nkL
p2tCxyx1xmD0DMftMS8ZJS8Y7K5+8BrlXNmAZ7XQkSK6opQza1MGi8y8K4fatkyD9VKuocCXgbdr
fEzWkjJWBiIT1p3PfbVqnJ12FJFMYkaSr9TtpGIUmuCp37ZWUTSrKV1qOHN3pyLONtW0a46AFEVC
Ka1x2rOatvBVdiVycXGfDMPYzq+hrJCtZErisHIlUyW0ngsqO1FFMbxAI3XZ13z8Hi4C77ikE5YU
sZ4oa2Sl0TkkgxFLOsvxO2tbdOqrBFHq04sEAb/UwzKSjbfi9MX/pYxMlE/UnqqIkemMLTRPKS4A
8hqEMn0oCG9Pxu/sNYAmL8nCVVYNPWjZYqU2aV7vt0quhZspJ+HFTa5YpjPAriNpQFqVugNToOuw
mce/473nFN9MmdY3aB8b4PaUDMEOiosRXh1wfQu82DYrLFgPDk12cxy89ibqr63yp9v4KOT406OD
Uy7vnRPS5Rmk+3a279q2sv+tLSDd21ghrC6AbcE/+sb6R43UCrViUlrH5DCspCFMAHg68OF3AMO3
knUAzszPGldBJBE4eqVVWEgx1HTL2kP2HLG+Un5cYGCqJctdZZYm67Y7XtF6dSIqtTq7FhO4Em9O
EQYGX2Q39KlZeDBM843rFmhBqfOCPvmBOnmquuBsfIUoES5zI9Adm+USoaMflP+yYgqS2+GalstE
DhHglFcJnS3kisImEGYlKEQFr9+UyIFkAHNQcLPxsQeLkmCO3zFCOBirq7sxPkx3WRTIAe6qIWkE
gBumBn+oWwV0qElqIBaHl73jpBRkjMFsJ8RyuoWbyFH1oEDANBKjN7CUCqK1iXZZXLWtTgd5iO+2
QtceVH9v6uBC7WxRbcNQ4dY51pxHHDf2BO9bkwxfudrjCggELUJgyVraPcmNG+iIc+kvCW5J7OA9
x0CsEekUlpsRw4wqWvgKGFAkrJWR90smQVtyce1JCelyBC9Mgs5wIJu4gKXBufomS/7jT0dRqy9r
CTKIL49YvZUFtjlU+NMsqmsrwYaAG+xllzS3GSrYJqNRVrF+4A/Rvz9c/p5xBm/R4kfRzbjhCugv
+te3gt9ZCpe6xOhl3cL5w8Akl6R8RG6U4zsY0CNKwVgMREEN2n1D6X2J+Z4qjk5+P4NYD8q00umC
sq/ymlJkcZ2APltBugFFPEzESdpD6T8bMl4j6yROtbj9YHJRUz8YUqsCo7V2HoBcM64LbOCAUPXN
i8R6vU2HZXb8uz0Ddp3zOXz8FujbMUYuXsvQgvH8NGNepOspqYpL1hdqT1dAh93ZfecVQikrxFSw
9pvyUX0MK1idKtk5yCsHw1IY0fbjVW40LLGq4ygwIVrSqIBk6Qadj+gqmjQmXRqvsQhNV0vWr0xM
4s3U7TqqfsucYYv1EeaP23f8B2NjvPs0vg0nJY6eOY3V5OcSC0gbQiKXBxxKhqaMeUpgq2RWrmcT
n74xrP+1rkZBGU+NT8rzIdjU+EWvGoS9PF7BB5cfohbzfS2A8WQWsPzGo7/OLr7ffVGLnD4Gz5Rl
i5d2KsO6wbRYkoWx/hidSLn9+PraLBaDAwEMWAO5kuXvuU67O8rRmvN1rRsEdHN134HRzSUX98+M
eoxucotwBu+5YbsRZbP8FciQB9Z1d9GMB9dH2nFxnKRAkCnsYXnCvqpBG19BUKyIpjHfte7Pn6gD
NyaM1KY6eH7o5XzRtdowq4qpjBtnN95luWIigB2NR9PHZM61o/VtXRI3dG8FvJnh3mlZ1lB/Fmmj
xcaLlpQWS9ledJPLH1rBJVFeDq48zYLnMOPZf4XhlK8EQtstBFdBMK28pHVfN0oD/xOz9RVIyIan
jZtLBHGJTgME2m3UR0etDCUsjC+dMIUwZU+6QmRl8M/8LkoseInz1ajN4HFs5Ms46OeG3ZHQffRR
lVsLMBRfuVeInvq+fwPyQyeyCkmcgwHU/N8diN3KNAgd1pjW8QQ4dzv/XoCCHar1c6gYH4U/y05q
oNMDunIVjeICGVJZ5BG6RABbvKjfpoN1FKk5/SoVoUnNYGEEvqG9Svi9JcQ92iWQwNpBLvCLnKYb
QV81ZdMgqt7kWpiXZWm8c/DWW3iSPKGCJ42GThnx4Bx4mkxVpOaqB/sjQIN+esIYPWCchlGTDh28
DOaG6NFIgu/x3QFeaBRDUsV2PO6lAPdagdR8AKLZl18eyfEymNbCDu5LyKtvuBaSkFKFei9veJHG
YOl8g3ouDeSoI001kwJt7h4HhIR6VAVsUIEdyWZcs+j/NWSScd8cRRtfs+3nwuHA8d4HSuYGh6/J
7iTw3gRajhVeFNwaMePGXc9NkIjJnFKbL54dmE+N0oiRWsMKwNKvMbZRwcYEcBYddWlRu+IRa3+9
lmyf7/lJiY+x4U3XpZfBYbdwvwhRzk2vU1JHmxbXHBM46rAUjr7ErUpWGwefU7sXdONCb/Q8dqsd
L92/zqEVSFQgcPLE1QZB5z4o1enhCYq2Bb/h9W2mdeIbz0xdwZLDJzGkvdM+AnFLL1azVXx3F9oH
WOFYxl/E8WPye75ooB1CxWGxpfViPHb0agOe1rPqLMV8ZNqlrXm4LhM/xUO3lbvTZ+K8S75oXiCl
Nf0eh7h1WHGmYgn/zzEctskTYNgtBvUobosmbZYp5wJHWi9uzzZEV/wS7NWO7EbEXoCbpGzeIPwi
hPRo8airnVP0U7gBSEIrC561iH2HRqumCExvzXrg4qj1NrGNz30KtIj/6eRu9avpAJM4qzf0K1BJ
TXud0+7Avm9mU+l5DgH0ISiKja0pjMa/3hmWcbJOrCc8AP1xCRxIi19yd++JmlUIx+palaUQPk1n
pvG/90Npp/gxXvOnZ9w0MgsSSXWV6zMGI+0vJcKy9+LOjoKzkCPT8hZg6LZDxEzFZuJU+deTvyDX
FC9SElnetwL7SEJz2IeYtytyayUYmNSeVCT8qoaURm2xQuZm0qroBID8l1jQH895dlu0JXaxp+n1
Zbq9D/ugDNmFsqj0PQAsRhwzgT5DhbRUI1AO/TSqmtFq1jShEbNKJm7tWN5hMpKfW01d+YL4MsgM
d7449ZP8j5m4H7Wp68wem7A84BAK68DqMpIy3ltLTNqn+66xGLMSoa9MItg3uf5cRwI8L64Z3ZWj
xez6QndllSMbUW2p9ZTvkXSo8M0nKJ1PMzs0jdndiNzeRgcraluXzCkQt3uCCwsIx84ppY0PG2S1
eZUZvSkQF9n9Fdj5MfAQdNETo4NQUrCXgfQGmyQCF+U+247MO0duWwoyKSmO4sALojnPVSnCDM0J
iJpftIUUp1GFynh7z7aIpHme+slyVW0Zvi6PpLCZW5KHsOi3yJMHCqbmcjBcx3J8ksTT5a30Iq92
FfVQpK5wHSn6fEiGYkNSz0SOs0ocYRUfugaxfQNKKwzgh+YN61z34nc5D/MhYze7nCRyDZgijQXo
11jujugYGajDTDsuLvkpdZwrh1hHpsklav4hhY/zc1N4xPbb1Zi6hlyWFwxGkOvyFTdKqtkMQAG/
Ik/DTG3YsTACJeAtGamAa5b6e1yq/Cii9mrU4WxiVL4Ve5SF0wk8WKe5yucEnIUeycKNAwrK0TBD
hpA8oBwbxHAKd/owrnrp21nFDVu4/ICCoZZ88HRinGs5juTPyCYeskwnB/K3vxPzO/Unq764joLf
gcJ7wDDCp5wWi3XQOt+c7h4sC+TVoxka4bgqNpQLTePm/cNQU4Dz3Y1+iLE5vkQ9ifpJrZanh6Xj
o9eZubL6t0ya6NPpzsngIWu+T9Y/hqyKgpazvyScIvnwFG35fdQ2uCLGBGTqqnEKKkvLU5weyk44
KARLMrwyyeNU5UWq2HwdGF9nl8GNh9QNMOOuR3Gi3FEvwvsZdgNaMlrlFh/a3yHEusw53NtNBJY7
sTH7szv4iZOt6hznkbGYKv87RjggODPLRlbUrMqAfAZ7I2eY8sRTr3QLtD/Hm208P7KULS2FDdtC
reaA3ssIURtwf4wsJjqclEp0yVnGyjr7Qr7eEX3SIpFXGFaGv86SfgAiv4YoR3f8x6MXi3KJMguj
0s3LFkzc8KXQqf6rHf4rQSIZmhLSFT7ZocsJ4BxU4fKh2jYcQt8tAK1PAH9HbIBVl+r1b2hDHlFv
7Lx1U4t6FHXFK6ORym0EPKgJRsSp+eBzrNFtdu5VIezqVSzAZq4fP77T1/T1ZAsyW86KFl3er8y+
Js0T6ji9mlK/J6QcCzBjom5mIMacpcmw0mOj6aWkPemsRlWczjCnnLNY6KGp2NmKrjBrGWqpoDzq
5uoRsYl3c95YGhJ8yvtsY/HneMSEsr7pYAiDsxyXznJ5UPoZgpL2D8VaMVAu/NH3JFFVcUbeFFuw
iMw18oCX2SHZI7LL2mNiASSJttxF5uZ6xmfS8IiKIl4zsv5LssHkAUsNXaT+yWdRfKRLdjZSHCd2
snHdL2FHf8w2t58RAWQGu/koLXLJp1Lm1gpE/aDGlBnohs9GwpSvoBd2lwQbeMFhSy5DpQ6Qe/0o
ebMsjNsm5lSOqSG39wViHj2ZmR45u+hkx2K8Bc16uTCzIB5nY71fFuAxFNgQUreSlKZ6T6cnJvSy
AQM0H65Ou8hSLzzjbH2gE5ltvpuAQlzEb1vAWtR/PgcL1d1Z5FOx/V8o9SdrmqvIuVSpa0osIWxg
5tLPGmsNICBvK+qfN1Q7oqVVUHjv2yPKgxp/R9NLs2a24h997aYqDkpB0MuKhV67y3/FTXanAl8v
Vz7KV4z+O3HP4fYNyfsjmlD7SgtDoR7CG4MAkiQEG9p6R4Z0pDx8vlWTq0Q/pC7KL1JSmcMDMbrp
JMOn6nAyXA/NmdhC2Y9OnYyMkpewAQPzTno/UkrXn7Zwo13e9Xn/oSF6UMLdaYkuigASOloyoUH3
x2DG7pRAjF8fxKxoYZH/HYZVH3tWrxfcg8yS/0Yn331lqyMecXaOjE6trpITNHdaY67SWKVJxTcx
6j7vCFwY2vf/MNtBwPqyDBhailn1X6YA2pMuVi09DltBoogjd8Srk1rPiffnbMKgYXCbLw8t31VZ
KdpRC7azflbLVfa0/iICZgPV7P2U4UjptQz63GqYEZq+hUnRIviSh8xfjnObACY8Jy9VvJALSNXX
R9AXhTwT41vCdzhee+ehVqq/u6zlkFEcTNgpfZU4rkKUvlVU3wTbPBLhczKZP7hUeKaWxpbRfV3g
93FjHBYJAkD57Ei8kV4P44FHv/HGoymo2sbF9imctWGTZvfkpK+f3jHod4/mALnOBOPskq4b3u9M
Y78hZvipb0p0SlLMGlYKi6OxObN+/KmSo81Z20ys80dR5v2t2YNEHNpe8nubKuCu43zFVWgjB+ji
IfB04Oj7+ym662KEUI3YAPTEH4toA8OpCbHC28ItRP8LGuuYlXwqixqJ2jiKSYydUac3tEb2HzeN
S2lZrV2qq2AYzGszyexRJ0HLbMK3V2rJEm7ZcX2aGGlQ7pSJLiAK4hnm5ahf0eniVOe/Jg1XcCkB
91E07F0rBqYGi7WnXMnSaC37sNFwIFKKCgRgIRh3pxa14dDvKRd5PnT5qR/jpI9vKCltyEKvgu4t
r6yMEoolewIMBKFnRDDnqP/kh7hxqPimsFOYpPHw5LZb98eHBr15nboiYBSmmUApFMEp2ylCUOcU
HdgQaltvmSZVNkG6KHWspuo9JmzCzWK0s2HOBakLZOLd541YrAFyDpbqs3Fy5R0bXAn9HB0Zc0mq
JFLUQB8Q5e6LZw+aHr7bS62t475N4nqp7uUBrjh1qbN6izQlz9BcAkA+N6P7bhqu/DOBJ4paAQwo
+GJuQYfq6U0Xj/7gvKj88rsIr6wv2AdKQ1Rzud7JA7QyJ9Dv5uWLIPNOk6FW0Q6ZciufkJqTexkd
9Qoz37aJ0QzMtjmCyizRmeNDAIeNi7pIdU03FaOPOAT9U944WNmHUJ4pCdK9FGVPCcv+aVGwFCTr
yiyrX757a7nYNAarAJwam0qdLedZGgj5om2khIfNQnRSKYgH8SSfny5Jp4OvS0vJpzJFda+R4a5L
ykdwF6f8f9wLwIJ0Y6qPlsBIxFGXpI5Tn5nRY3LM/VJiRoU+6/ScGPRORn0lKtkktLyc3zwQVRU0
1bi4yN1VJLktE1Os4FL+S5WE8g6Nj1TcqIPyXDVfE38CO7D6lCgm0gdpeIjKSKNyA4fdjpjiChPS
sdz/UnJFgBn/6deKV1qvo95ad1oE53kOifcC2t9DVaa6nzAjmuRLlkmn05gJGBSHWAYo7pRY1Yu/
yq9rGoNIWDcN7CfLZUjza3t6zM1dY0WevKm0oZHwjN07br9C7HsdEr54zVJGTBshap2Wc5vDZXHv
7zV25EzS+vJPN2mwkOEKGAkC6hOeVydOWkIB+qGem65J4IjIDp3Kl1F3KKmluLknJicclupioIqU
JGsg+Rb+HrXPDvmie0v4ajfiCde/QU2aQD8uK4iJaiXgE7tTOCi1tuMqZomWeMLTP3INTlsZJFXQ
NneDP1UVHT1hqXB7MKYWLgooKe5eiSY+CM/Sb5Mwr6nShJ4ld9WKujs2UFQSgD8i8a0ol18mSnpB
VxvGsQMo6iPqi4Tbqtm+fZTXfMNvn7yz2WyDardI1IWAAcCCc+XxHLPr1/shhZyxVabo55zkZ4uY
SKmEXzQRYfttcuxrkFQi2XZCJM0wpxIiO78d0XtL3U0MLBBwdNsLSCU3RQkk4gGmsSrimZ7t8xv9
9h4lTfBxeIDibj1VUBS7DvaQdzHhJ6oxA8g/Z867P2ebagFuXnoKpuHiUQySteqmYRXG2cZRXElU
itrT9s7JCg5LQP4pfVDKZ5E3xdkEAXBjHCN/hEXwDdlJR1STjCghDlBm/DAAZ+tek+yvCgfLoPOG
qsgYz7JhFMgBOcMZIQweFgGWqutAAo84MAoVEPmgPoRwv48GfLel8gpnqPox4vshr/hIUvuGnfZk
3GyObB5XPAxMUvIkTaz6jtBjRD+7dlSJ/OAfoEri65XxMfpl9FLoBou75l5MGHWR03uiC77JWmyS
3NmGrZD4ZUrrfj9kyu8K6nNmkEWLqam5w38t2akn+Xz6E1deyepx6kq/PVz7dLumMeBwmxjXUEed
gjB/ETst+ToEKkM2qZXQHH32Q4c0UtIg4x+GXjq87owpcpleRMrYcCz6O+rFJ4bmnCfS9JATKk4s
+Y3Gk3KvLQzIpolM0IvWqSAk5QcVwi8ayxroj0llKsLncWz9vKSkZLe51GLRLkZe3uw04piAG77h
fFKUTeMg3xRJriFmVwW9Gxvf79fqui9xy9JnqjGE1xTCAPg0izZoOiCs/m03NgjFYQmegUaOFOj0
al6soRsUEr+21Z4ZctrkWNzOH7+7IdPwlaUaOL7cLDT9Lo5eFhRDD7nIv3pd20JSbHE73xNUF/LL
5HLW1tFpok4i3jUNCYmEtJKl66NDe48i+z96v0RTRa2lBdS46NX9j7T0GaR2ohUKO7MzzF5GU4BQ
BUDYZ7jHWd3VWcno9r5dvmPqwvdVSw/3BV4sq+W4Q4LG3k3duajCupnaMlKIIAyKJlITo0A6RE42
X5drM5+FHsrOkQKIDmDxTDg74KLuRKgc3cKg/gfPVaH3RfjlzfhbgEtx7qok2IsdHDoedys+9ayp
zOwBNsHbMHLlYBhexUWTE/wAGXDHxyJYghn0PIH6oJxrXsebeuFSORwTIEafSaHp0eCK7dGXVRA6
vg6vlebdG8r9HIb4xP0P4MPAeWW0cI4TPZSvcBB9Kk4NAblxZ0YUaXQaVoeGqvL2opXZ2OpU0COO
/i98og0Slo4tegJHi3wr0+FWW6gXmqqm5/4TOyTA6tQVp9ctmVgGQoWUHKphlBxaw3IF9AwnHzKx
sondNijAjFkwS+JxRrf8ctw8r23IWbQ2okYsvbjFjv2vOcaBbH2NAywAkAQbUq/c/9VdRgYWwpZK
9imkvAYJ9SkMLYalzKpBFR5G09SBvI111fJdxEKSSCMXqD8uTOnAlxElOC5FEwoO/O49ByPFZrgS
+6Zm5++67nXXy+j7vQTP/rE9ObGK4VcKJiPVXLH7xr6vhncGTV+M6GxYY7f0jTM1v7xnd/eR4F14
qcfcy3LmxIzG8ocbIsesN1UGcdqeVUBP/05kfYmKqNCJcYqi1Df+iPN/rmuhUQR31/2vqGxVsykP
xjHRyR+xHa92T2RolW8EE93Hl7XgTd8mhvDRFvd6jMy20hHPy6aDqK5EtWmArHdPUjX0MEML+PKa
wNN646mdz6/onlgsp3nGqZIIejlo5Sp3H1a0OrzRYpfk1poFOQiiHloRQ0ZdcVKz7Yw4jkxymnbN
D0GgAIykh0JB8R20vgvHFp4DbqBTetQRxqrJv77qJ5LVeRAq1KRvLMd8ewm4kVxdD7Tt2hGL+Jes
QZJ6k1GIAqT+BxO0EMmWfBKwPC0NXOJ+4Ldqj86bEZ1pZMmQDeC9Abwy1LSaEf5DbbWbpB1yID/y
xl/blqdJRFSQkdrob58gEZpnHe47Nv5aQWCjLz9pYtgaliLmxMnwu9iVkvLYv2FL98tHSWH0vVf0
MYUEU9yt9Y1+f0ww/Q7kAJs8zKa1bK+x7e6NO4Pk9et9OTp2wbTBSBVYAWXh7i4GN/e3Yc9eh9Qn
p0CKPCu6tiyR+kTKt2XWvPMWyKo9oOhNBLYbgHYJxz4wcMR4SDv9E7Ij99JJ6GZD9/oRGdzn1p/h
Xk0fpexPM0fABW7bLQBuWr76gA+kM6waD0sE7LEON/J5CUdASVRHGIMun7uHOzFkPT4Xyc0eJBGl
7U7Bt4O8TCnUa3JahS2YEsmZio/JFPJzfy1CRljDiZcX8FZltK9H47qByK7/myHhB/M4jRckGGxu
0xpPgIp8c798BS4XdklqpEPPMGTG+E9AHKad3eu7cZ3ewb9CIvKQXX1SJzYo4aXLOXQj5MiIBlAR
Ey5JsUMCTwOzmyJNLC8Mxr6ahzytJctTrv7nvnFuIU8CX+ZEPj2VGybpNDW8vmiM8D0munMx8RId
GoZUOQYY/E5myi0BjtcryHZVtvV9JYcYDM7Ccl5580Xs5RWLH4b6tLlmmtkO6H8NxL7KIcp7l7KG
gXZATcwdfWAZZKVTmegCnZJxo8XX5MxTMYcz0A07uB6X/Otc37f5y6lKJc6Swgdk9I+QBud8GuyT
F0kaMzpxmGft3BlO8kyvh5UC7RLFU2iiMu9o2nVxwOPrmmkv7s0YSesI+2H6kkZVG+5PUSEl8B8i
AFOpruR6TTkK+SgzDLuVOGnb5MdOVIrEo5okWBhuT/4qNnMuQSxJbF8Xw942AkdZYFsrM4H5+mwR
WhVJ34qb2QVxwJV4Q9NDZnMurk1+CH/zagmZCnXBnQ7uBcVOoGWPoXcvCcf9FHzZw+QAw932FvC/
tuByYWlWNTWQ8qrrRWoh4jlNF1EJs9jHuXstjM6HdlWCYNeJ5MJ57e70+bQA7D9kR/gcuHVmSM9S
mfKaCC2y8lfGIKDHwbRL61Lzn7X/S1VsMj+mFwQl5QaTZYelSRBGpZwmlBQHTEOfuLD0FY7dgBlr
dmm0YnfRPG8RY6RZbJXn+QaA/TtSdS65ZumCOEOLK8DVDDSlf2u7XA7uTWLJUfuAQWbc7C/dgoFj
Si9qtMMmOB1HrXTbXOEfmJ7zErSe+1uNaO2IxubedsO9w3ogry5NpoVgwtYw+V28HEUF6X1Uwhb8
AxmHCLZ1+zHKiO53qLKbPw+RjE8SqjlZwl4kTJPx95vWs/b4IEOu3/SpABHhz2ODog1K5lOjiMwB
WO75O6mvJPZ9VS6cxIgTRM2En4r+fD4UqGL0yg1sdXMVvqDnrF50bZKgSiBwOebo7OfFlIhQRb/w
1IyY8K9zc1PXYeMbs4AxWRb9y7gD2U6hIapymLBS5S4EccclAUBQbsyxme8FhkS6TpiW0HkwPy+v
fwaNC4az3PMRgRWNFNUTy07VrfmisKfk/FxEfCzFSNJyuQBIcFuzjYl41xBfetaomPkjnB/PKkP0
0YZdnKNob3mbE0BUBLaLG1SROm+xHnNPFNrBGgOU5fsTxqEGLbn1njMOfb/AmjACxwYG1mn1+v2B
n3l/x0YdCNX89cnUH/ehhMKskpo5QQNCkyZNRcIARoRNdMQlASyFZhjY4KFgXncnqB8us3e2Uslr
W2LZMK/v3YH/1MWo6vWDQBwsVWqh2lHTiEo3CAq1udDsA+g9tBe9PBapgs2Y7w5QyFhVpQkza4Z0
RFPivusWwiUTxg3j36ndtmIV/hiOVsUPB/sAl+kQmCb+/hKgvUdbL5Yq4IWxQtKU3P2tok7u1b1D
URNdSvHmWKhLr4oWPPLRkzqSBRUMpBLUyhc/MfkhzPWFvTy+YOdNJXdaha6Xn6F8t27F9QKrqOo2
cRnaypDPLeNGWbBSG0xGOxRFJqAOxBuMUalSDY+5PL2VknDoBP6l3Jpb801OWjwpJdOPaoSQMpyp
i5hF43ggZRlA9L3TaQM2dfTzWeONw12MsICPuHezYMi2OAD/mJoQI8FJ+Ju7KYhR4OYlVZQEkaY8
aydoQuft6slfMfMm8mfaZX/AR6r6abjbf3nE/8Y7D+yadUE6z3+4t65OCsX/VL6v7/MAmy2c0qoS
LZQ+sdMRSuiNf8HMbYgxAPFco2vcJ0xVi9/XFf7v9VYVBKE9pmk+NyEWl+FPyJ9elg3TIoeQ0zuS
5jLY5AkoS+C5/BdO7VwN945XYA7XqdGCXImFpmrslYY52Be9VTs7X7hryGiKGc/Ie3RIVVamEtbY
DYlcy7avo5hnQOHNNe/hRTU9/kANbe6LogIFE9jAgL3r94l/MDTT6rsUslC28J4TvMTu9qA+zY6a
QilAkU7L2o+3OTbqzO4uEn9Sv951rIJRhfSMyDl1S+Td79+tPALuRcI7AjngiDcpXQKPMdzvYQ8n
fnL/miHRaTwLJEeON/cPqluzDwXxAyzSZSkVh2ND5VMLUnrRKgk6SW1KzzYcVP3I5Mop5g2D8seA
VmjAqC/fqzQMnh7KPlWVyHS3moY+7Qz+HUua+uOJMqD+KWvVTD7tDANPmTmKfc07RzqCWdUQC8oP
ctp+siuaeWfYKdovyqdaBbFzRi3PzaLUiID6SN+kGPCDW9/PiQQtUvtAnCUdiP2J1YACugxz4JSF
cE4Q/tASlN4T+gPljlt/+TCtCCLgq+WpaPs24ipbMnBHsAqlUsj8XDEFAx02o1yCYjZbHiN2NLVb
uJ0ODL7zdgjL9w6QhzNGwHyBaF1lKtFB8twSu8wkXYxYswCu4qStkyBmkqm5l7SB5ukxXep845BL
arSR39G/++zTg/oJuGPnArGe0gtszpajvMlEjYR5pwYWBJRwBUZkv1lpKHSm9aiQV50OJuV7GOgF
YacscnQCt/baPWn+ZEK8sXpQxFyBDX15fhB3SjoqEEA2SYIsqEHN9a0uTnD1yndfSnAfHz5BXcPO
+7640dNwkfWbwvTwvKFpTCad/r1JQ2uK6WePvAvklWFsNPrxplqH48nQkq2Y3zfSmYulnZX7bYTz
1Rf6mI3BWSHTbzM3mWSpXnyQxjT/ZttDTfrK0YV0R2xxFbBRVZO1ZLNInDQhoPsplJ0WHB3MOIUu
1ZXqVjpppYGmhTThSEunyUpWg9qQFMKBF4N+ldfmgT4c+ysHdz+yqfqJ/wQ5zF8Aj+J4u8m1Mf9p
+i2CtvuA/BGEhLTn/jJw8VXiTxJyeOFLHGvlygUoWi3Mx0tQmEO8a28TaAEXi9CmifliD4PxAu61
hBN0B6mdVnscgXp67iJ7CgdERQGaT7oYMGnxPRmAMlCpnRIraH2vIBF6SZok258qztoibqcApCSo
BAaNbmyu7VuacVK5dEW+woiazKjq5WxNgam+s94bbiC+cl7NsNn+bg/cGALmxJ18vitt/npqFuh+
milhR8sgUjRA0luDaao6A/sZsGUbUwnTVNwWwwTdlLiXXH7eK9q6eobOXHkQZLsC1+6xqt9aEgTJ
FTKODJuuurmrF45SX8x12Uijl/jgjp3+b82wCafHTyZxmAjSsThhsvUosD1IW1rv3pj5sduZVtkp
CGKHBoCw2Auds+5m8qfFzA1zIaCP9SGBEWPTnjDpWAiC1oE48RFUWKCQVp+nljwQ/J38XC/BtC77
ctp0JDNqiTwowb4ByusiU3yRHUhsK2voA5AagvqW6fSQQP4bMGlJgfPAUCBeGLRohqz18H88FbBH
YVbkyqrEGp34lR2HENl6VdYnZ/KsEaN6T5fCD4slRDCM57cvUVkFJ8x7oE4vPQBpFI4kaeVeXgas
xHx8kYiifj3Ao2xr+MAOKNyk4S4U0ag6i27XnMyL/iFg4Fm6DdtP0wADp6XZtQBSYcsby6QoKtts
S+y3rra4OFHCiK0HtZGven50GHJF4f1nZQ95wLhfWv1ajUewjUrgj7/mZhsAfl32Az+86hUU4ZK+
+B/3rOiPdF0lrjWqNwQpSiIuDphL7fOSgs40m/ZhEOal1hA5CIDajZlKEJGycweg4cugghXrEmaH
VnjnktOXKEYf274+xFt79siRzqa/gk/PgA9luEe4egTf2mla564KR8AAaF/CZnrbXpTbttR+fVU5
BrBt8szOjUujmZqrWmSskiqE3V2MeumkgYm17cO3Tn2e/jYuRDfqurZe0ebG7w3SF1LJT4YztaCH
BSLZmaJoLe/ngzYtTsbAI4LKqb6E/TQdlzCOyVBcLlK41RGg/p9NubWKLjzbZQuUovaNfH5yNuU9
5EobAYv48B4KOgFs4vfDIuHq2vzQQb3CznMNd7LFxciK2eOaeayNr38sefxsa7HxULwi/sc7Zurn
K6Tu5xooKf8qCERqt22dzg3TUOd33EceyL9ykwiu64MQ1AMfulnHdBOSztc68QoIgASyi/jsu07t
vbHojUwtuJOHPb4KgomtCp898kYVL6M4eQBalo5hzaAzIkDXaiSJUyUt5Cjeq9Jc/IAH+272CYjj
az71pnqA5AU5D8e8WuxYBYBCGpgE+/yKtDxTWFnAtb4GgYzEa2W4+RV3b9HkNyHCl56p2tPVHPpO
dGED0CG0YhPFy4Qm54sAbiyklPZGgIba+ZrUu5OgshXIlmLEOiqhIIjd5EaG309F1A1O9breRrY7
H4RjHwitKerHmfWxVD+18SVEkGJy9Q+rNvk0L/6t3C78J07+fxk+L6uCllixz+7sCGJJAMKTSuTa
HFX2pynyooSnFbRgz3tPdHrzSQpdeWMbGxNQGADBbT9L64stPPoQfAF3d4GKHZeQmEqGygbs+D8Z
txI8QLZc3WetD4srk9RNbzf+hkVv/OSUsnMI88UUl8Cg/2gmbdqr/2iwMaodhBefL0qJW0HfhsfG
duEhZDT9dVHxFcFrxpZlwT/DmQo0Pi1AhcCzOLjAHtIVz4YTg9ZFBXjjwVcrHcDbNf32JOETIORS
DSx0+W9DLw59Kw4v8hAoK4lqbaEq67Meyl+qx55SwSztsIf57I19VygEZB5VTSotIyJQ3yBZ1Wqz
GA+6ZuQEG5vILd/bZHX9E8HwrI4bPG0m+HUIViH6Y5xkarrKZ6GWM/DhSmE5h626VuVhHw+v4A7H
nRlVsoAadn5O5ZAyrawrnNccPToCJMjCXwNs11qiud/E+4Ijoi/0SlE8jZ3X+5JM1WhI/GvgfsE+
4SNFqS0N/O8OBHAFnEOsMzbpTD5ExVPhZnNmHCquaEUHDhhogS4cs9/7ORrJyZ04Shu5xLnyMVGP
jDFKdWULOMg98ugKipv1Q/EarEO5VmibHPt1Eg9YsMJxhZp7WjcZNcGSFM6kfgmRt2DOTMoglL+W
f+4Rk4Q5ZwMPQDDAoaoeGsca8r33mzY2yZvgeveqMm/Xoz2YdXV3b/HLbAQIgPqMnaTTCm+m4kj8
2OpXo4lTnWhugsnY2Tw23dOlH2LGDUFuXEqBH2IAr/Y2kHNZyhVd2HHfFuINzsz4W/gf8f/sEKLA
37yqBVvPOYEJvwsqndPdzIvVr4ZSDcO6nQqnsPe2bdLx06bpjYJSailbu/3j0vjBHVXIJDKHdblI
iJ0EG4w7eqATrnuC+KxBSNTWv9h6tZ5t6Tfbnbkgs0tWW92JiXNl6k3egmm6JqVhW61BdqM/9Jlj
NWiwug7Ht67UU6/KzmRPjM/Q/C5pQJYN4rffoolRYRT3QCiLAAJKWxrxavAiLi63TlPSjU3WsSqd
zB1G11WX7xAaEzcdsxdfB/seFduZhpiUqC2c4xHOOiXSXJj6omWUpasGWNqFM3PQczfwWQQCkecp
Qvbq5HBgfBrfjOFrHioRcaCZm9gvqyhiQCQWjnisFahbc/MZB1O+Y3zDKOmBDK/OfbXL17acN/rj
rXEGs/VZ9hf6bb27QZUVFB/JhoU8o0hxnfqZiJgqA5y0V2pecBdKjQENL7zLldy1w1ZTHqm8DYQP
cpX9ewzuEfVmKsGXG0CdATNfvrr5gLt85D6MAS72XVrHmhfOQzNLsFcouOc4XGuuFbkchkYjAjm5
cwYBxNV/y7Kt2Jy01lOwAnUj6s0U5Xn2aFCZToqU2PcJ3mKBlW/TYcwRpeicr6JMycrbA1eBgZkW
97IC7pyXvkfKYgi3YMZwn8UGGfjfyyZIgqXOLe7LzkF6UCR/M2+khlxiRbJ5nqDsAIxjhC6n4v0j
Ek5REJ8CZXXW7f95JcMr+HYQBHfK6tH3w92/nUjqL3gkhcJKxxlhjoWn8N7shYW9xkv55gHP1HcW
+xzMnaxiyBJpL+NlBxbFn6kCgUUEK/8egeS3zF86If/UVEdwfm3dGm3bsS/9IJXHKRgRknit3kVZ
eLX2YxtY1a2FYPFIuHo3VXOXS9WYWOzQb9jZKb7by4Hgy1ijqKGl/khGTELOBaX0p0uGzBXqopox
gUHqivkpHFecUymLsAMbPet31L5R3s4IdD77DMrxjuZM7AVqf/npg+5kUgU0Czg1N717lqqtsboa
ZrO2SubKbrX2pxWGf/s9Flo3q7zKRyeaQOW35F0bA7il7R9M/Exob+aKTeY8T/Awu1CLvPrIGN0I
fhjiedYB4zA3IeLZO5d/vec8NDooeW8QinlOYrrjYwAA99XgGD1Ma6xzI4Ha3xbhCm/9X0Vm9EKg
n51J9gJW00C7L5KJ4NGwiqVDQYVHLoujQocPMT4RLg+jqmyjWkS5xmRkpmh5sLuJ8UBgS5ASzUZx
8HoVPDIP/ejslDl777GXtZXRvNpd9ve0bB4rnYbsVckhrU+XQ0u2ZFIEU5NBDZM8pmViCVgSExrD
gXA6xgcmHlFL6hUZYy7ZHGoxQCymLxwJAeTMeIRWeX5CpojbXTO84LZNzxWyeWuSiuraAhHfUB/4
n4bZ144UTRDNRiHiY6x8v88pz5VUTPl7yJJk73KKQXbZUmj0Xd2qnyufWkSYhBd6bWjS+0mFEr8k
2hddTvkT2FvHu+rwH8AZrkiUHQOtB71dSNKer4sUnjkVEse0K6cHkbnSVu58juSVhhFcsJLbJOhk
zoZU4jXciJBEpY2HLl0O9XFpNU13wWcFAlXghr0ToYTp6pD6TgDqO+szEFde566OOfcNQjPGZTGS
NBluL27thp+YP1aDLIP9YXL3ZkHlRZYoJPGJ8nmBrn4d2+1B5WYWAr/YRKGyzBmdyYU/Bm4n7qC5
73UioRiuDUnVk3vnDavNZA/Or9PIxikalWXJo2g4ZqrOZfBevgHAEYcPqCFXSYIEE0VZa2UQjMYY
D67TABPfrhaPZ+8WZQDoNQhUuU8mBBRYRJBHgk6PP2azF/rhaCRP5nNIJ0l2768Z9ipU30Q3eEmG
0m8yAy2IVk4oBiekVg1ZHZ+QQOhLWL30YKouA/x2Sydwd7o1uugMk1Y7KBQKyzPdtXpw2b1WEemB
4juD8ns8VI/mlrzULuyOd3wXZ5CMYsPrUlQ3HB6ylDP46K6kMiZbibyWccNOwzNp0MhHoBQeMDHy
+adaMGnSNsvE75bGp+dBZD97r7l5/0vMOM8q+zMVUVsWZhWQPDcGgFEJGvOjQJtIQboNMTw4hlNu
nR8Se2wLUL+oQxrwxMa5z3LERmQbswboW0i8OZBa0f8REHoaWgmFdowylMWCeeamM8L0dLt+44XT
OIyo5Y1nFyjNIk3P7sjFjWRNg18SztEE0j5G3GLY+URe538w7ENmqQMYrM7jsF+EcqXdROnmj0Ti
ANdaXfrqwBzPNL7+JjJjmC1PBvXmasMqQ1SrM2CK5gT0TCa2Tol3ULh3WVU32uVkZM4RNyJD1O5T
QpqO40U3ksAWWt21zbQ+0q8S2dn6aKP/nxlCOxLqCFp774wGDGwpFqCxOw6TjHQIt0/oHJtYMaXK
m5ODhm8ta4ttQa1y07HwjOc0+flZ5Jc1GQPgydrrw9E4gg1G285yALaJPcjbvDnnhPiZ30MvkdBW
iZAILyoDm70+GwMSoPU+MFoIfFw3CPktdKWw8mcm0OGDsvTQWubZkFt0ak02E8BYv6AI4VeG1GMb
l/94fneFpVUqbFkLS6NcBBpH7aYGGfBO8HjfFb1JVUq5pASKi0WGR3y0UDnJfm1H/VQc5tuE/d42
lGro4MSisiHM9rulUPN7hrchmC5JcNCdEQzaMJ7Us9dk6xo/BtJ5VXrx2+8gE9A3JwUNK987N1b/
3XBnRTZLIEmotqn2vks+4Jh+6uV9RFhPyQfZUdKgecRJ13hp1grrtw+LsLg9ozr8Ko71D8Hrf8GL
bvy4jEI4N1ud9U+340ZFrRPD6zM2TMH5pnlXXs6olRO1P/NxRLA+FDIJjadxaWT8uPZCu7DTozPP
UAsHL6PnvFBsvpSfZ1Ll4DIqMNtc4ityWlRr6qK7ARYGpKm6x9H0PwIUpdUjkjdioZkdg/L/0EIK
Cdcr3vLqweq1WbSx/hTMC/45KHCLSV4tQpVAPuG9tiJzkfqnvwYzFwVikWhOQ7brXbSHkVkAKrx7
VdAjItzUL6PIxzVf5Cd0RcTEcBPgMRTQ/E2gOUQsWbAh8igDB8+GvfJhwhdAvpm7KEF/40XnTPqf
vZndY6NtKdBAdfkdzLQZ/UsO5k2waGRPfgJNj2LdFGBBoqS0Bhyysq3rhlJKEhmklDuEqufrO9lX
GtvKINSBdR4hpa8DBlsSx6MQ/rp2NyB/fEBgdbVWqwEzYzw87L3rtsaZOyD/GAUYrh98ZbJZXzbO
6OxmI0+cmKo5SdqYnDhuHqYEFFqy4XRzCbC19ak+0hsez1Ew7A6QZh+Ya55jL1EGeByOlGgw+5JL
JLx6OuwUSXz4axNx7V+qHGWFtfdWgTae2UEc/CvZIZYvGaj3yMMsz8vw9AnX0F02vBuWnOh1YP6m
UwOVObtVdLFmto8IeYQ1Ts7gQvJBcyDlWkBnKt4yqgCBHoY+CQKd0+6LHT9ROMpqVhNUg/zz1af1
6oKcKyMbenM6+b0+iaG2R+Y8WPIEQJkUdpLdsIbG98Vh91sUELiH9DpXbXGhlNhiOEJIetDqf5P1
EDdV+l0k+zHYugUr8hleiPoextbfVOC+fStVFZl9e5C/kJJa4pL2eBXcZnGW3BPeNHnZhC5zLohS
9EbYB1iFlD376OGEM8owpULVFL0O8xcXJ2oLZ93EGlZ7n8npC1qG7wr10w6DT0BTQ/k3DgHvw3mK
UCSMJavh3LcDKjO/4GQAJAl55DdBx+iqdUhp8BkBZoqMrJ0IKRp7MUkLHohSr+Mc7qS+FOrJtWSk
al1wBFYvvf+CGfb5/A33RJZB+MU9zBBG2uab9WOTo5yaxeCDpo2qb4x0PRmKTy9BXBmvSNUrxOtB
jTci55FcqGqicDRS5DajHKUH0bdwVVF1tly0gJFQBRAUqvVzH+GoAMW8fqeQhn5FYB3C8HYR8oW8
jRwTGyqIXKbO9l/94GO8NY+Xz+cfirGLbPPMrlTem/Y1VaVFjWI0EPcJQ12JQhTWQFHvUmfIagHj
uw1n39tEjsfI2Q0lVeXPrlgHKNz3HiCybUFVJBzHBaw1gIt7Ng7D6rkG+WU3Sz6WPKd53UDh0Wxg
MTXnT5yvMCpnXTlm0pKNtDUusRSyw+xbgHcxQ946x2JlLJHO0u5XA8lDwhv7ir8GKOy4L4gSY/6N
PJCq83zhtZJuuuUm4FrW+zUZIFcvBPMK9P6uSPDDA1vwh6ir84erOKvWY65QF4+pznFDkiKUT01p
KGnI9CjxXJm3W1Q2Gx9+7pfURiS0ovx2Id6DR0KmG99bG+x0jn5D6duLQaRE4s5pB0gmCpxSjmeK
p3VgE4IX32tCHR4j62XCfc+jlTkOgsPhHrb74HneuuOu4Hha70/YnIHBpVGy0Xhtc/3qY+GaFn3l
FLIgN2PkkTz61K0Hv+dUhMjbSf8ZFgNfc+jPLcCifn2N5lAYYMTHmag2sMXebvuJM8ptO4JlWgnB
33X0/hhj6BmGmIWGuH4RQkWIn6NTMLFfp4s/qw5S1XOkMLxoMquovxqcBDKr8N+HD1euezlkh7hG
iTy/rOyx2Pss2v95NxhGDqj6EWqUi90Z9rdeTjnEZ0kGFkiOgMx99puyAVnkSty/9tdDedZ0tKmd
82XFZFsbyn2ufyYoUWsyiLNjzkYP8d2o/DBN0rsOAVGQsVlZwgKWzzJD8MIGV2wUt5HF/bGjQ3Rk
TvmL68D/uUc2G/0mI7Rj23v+VZSVlP1gUDw5hRT9vr1EStOtHxx5s3gSG/Wwqf5QhaJgA1RbYrx2
pW4TQn0N0maw/UaXQJhg63IZ7p/PTDIkUnBd34ZJD7P4h4hICYty6diMyYcKZf+dVH+6K43ldusG
sS/sIB5fCIoCcoBbGF+Vik/njc5Kvg/BP/rvuIP7BqUxl/xCxy3o8hZXGpc2sAjDKrGb0TwuFYtV
BRuC+dItSTpTGZk58foWzlC/EWQ/cdYut3jd6lFF385nH+6xACL8/sXrKVcilAypXyNbS6HDMtrU
IrEl0Wpwo9ReiGgYzth6mvMjX6/4GDCXJbuCmVVp81xVMLXf/VoE9/i6Lt80rUVQdroiNRxkT7hQ
VaEzssJWSe9c/Jp+bZuVmJ0RhL7+EqaAeeIgnuOJ6Ir6GObmRuRFGSDXMPrYidNM5axjFDZ+Iq+q
evND1j6mOp5um10CpsHBHdF3vTcz+rAMAO7pBQrUvCSi/qNbp+3E/vO5ad3LzkyxEDW4rqIH6ya+
tkpfim1IORrGQzAFJPibWJWn8UHkdzhZACvxIHBYPHHHceCprtZMmRzdzdgJ3JLFgr6VeeomTDxm
ByEdNW2QQ4MrDpH3QWiCBkkhg1iG4Vg6iZS9kroui2tbrSeS6lCcYNQpLMz/RY8NQ/fpEDbE7IY3
LFdQD+bp0HTTAATU2mmzGhEA/0V/iXrETiW09o1HCb0QFa2i6yVzt5NIqWouV6RJPfnF0VGa1gpn
5yIn+OM1NUGgslClnuJ2+18VfwinJJ2Apl6TVjqfHT87fhwmw5yN0y6RfXnyVCebERyLXJyTCTTU
Jsq2ErxpRFPeg6yjsbxezsW3fF1vmHX+0m75zQU53OB5Cym1Miu9ZtvaxL+Zryjgn40tAPXDblju
IHdS1T+NA6c9W8I2q0uq03BxaiF7B7hdiYg078SmWFn4+OKUKFTjzuIjKO//mQAbhQSQLuSWOsxs
1lZdHcRSoQbkS7AAEyFj5N5nKGy41klILYpXJQM9cqWcfMqTtkk8y/mCDhAjS+Rz+/8mI1kOL67Q
DaKX6AnGKwprLA7V4zxxbU+XDFDidBuhcLSYofDWCTLYu2nIk8MX15CQ3fc4NYbe5mznrOYMIbrj
77O5xJCpQKOxHwLy6P3HFByK4VUi/AwsvthveL6s/ET+XooxcnLgIWF51Mr0Gxkp3cYjipLxob0O
ws9B7RRz2rhUWCkfWWc5w5uPGtPnyDYjuebr1mRmcX3GVpFPV3YGEbHcUasddTgnArK8wrwTJ8k6
brpEMa3qYN3ctCpPDP8S3FB54UPnCi1Y2ItL/93vKhETxGWrMlDP1d4xV1/hxxeb/HEUAuFnk+1y
cJG3gmMfU2e1p71MydUxYWp8AJfIGjBawZFCUJ35u7OWaDtj6YG6FzBqojJXmU7nZIs0B5P+A9PH
38ZLbcuYJBTqFJeOfyNMHlScwqO98z4Ok3JeBYm4+4w+dPgiEeX9y4tuJFiYzkMkCeeuUJhDclRa
b2Ux/PD7tDANmOZqhnFxc224md9aKGRo8+rFT4ZdNGcyJ6m0b+y4ZfRZ8vDCaO4W5xCOvTCobiJk
srhggfVYnZrHh5UNEODSiWcDSzx1w0XTpgyGtIHhsMaCrfcNloJRJ0+BTM94ulIu3lcoHfRoZof+
gL4qfNbaUJKoVdNtLiNU/W5VAzT46spa/mTLJeQsHeZVySbAXwNowHrCxgNKmScGy2aC7HQkuNtM
yCt/hyVeSAND8Hqteq8uyj+/t1l7syz9W2KDG9up/HKbSg7vFJps9py9ptoRC38pH812CRAagOu1
W7fPZ1selic/GMxfm6zP+EPs4o8uwWTS2ysYWVa4anHPv0CkB8OcLb2FiciAIssZ1dUtbWq36oqV
MgYLSpmCvYH/FLdWeEUdNKQw6oDfLKo3zJaU3ekfmNmccGvySuRL+6Ij2W3y0BCxMNZJOAweojxp
xlxGH4hZ2DBRf/l0gsENNRjUYObMRRir6mtuEfE5AA94JCl1nEOzHfEzF9hc8fHUs2tm3l5UXQCs
zbCzaiH0WDQzzlylNx+bM8D5XK9f/Gdxg0smv24GHvPORSuLX1UiXFcNHSmM/UaAChuOvssllf3S
kLeisiWiYF5AgK9I0Pd75cyYEZlSpptr12v4ajo8GlwUYhxgpSbtAZQD5wuBk+iyWShbXaNoIMuE
1DZ/w5YQ4c/CyCEH0ZQrEgDGGWJHXAJ7EyDzxSgLxQSs9yoQq6WWB2Pe62fzS6ilVk4dxS9qjivG
wja2p9fKG6hm9epUoogv2eHoMmeLrQ7LDk/OUQ4ddP4NxX0jMJbVTKY0AWIb2F4sP0SxGVfIPlif
/p1DQq6XpBZUWep1byuG8zPhcYeSCAZEIsD/Pnx71tqfImnl1oQ0buW/FIlv2feCVjOqHvj4wby3
7p7EW5kTyWuu98HyLTiRMzJ+DY8V+97TUgDTT420xmND5fNw+cg6X47SOEIvvQ+b3Sz4r1/ezKrd
qEMCWLSk4G9ENVDcFWPnqkA3U3HMEwrbmNzOXJLKkkWvl0ann4hkUAZhgv37FMzBoMnaz4knLsSh
8gRNs4hQscXfrgmowvPV+rfATVqKaSQ0442abk9qx5MvlIiKlsHEfcXHu4qj7NnCEQja9dOjXMEi
4udxhXI7zek7M72IPHc613JLMSEJRXzig9uU7z1RGgOZk4UANMEs+wLnbjL4VJS17dyDU8Xp91zd
DWoUfoWsl7WtDYjYdOFJjQDPstYwCyUdAqe7FQJvFEcb5J0rcTp+7TYAQnNN9MBexjzHGXedf6Ei
ixCut9WBrq3rjc9dWuyVFUJB3q+GXf1S+/iAM36IfwGHqoFInOn+FjAlSc38i3xj2IY51iTjU5D0
5PwsmKYesz7RwFZKU+JTcGD1tkSeobQyqtIROBJVFElQZSio2QtULWemT8z8GuolZBCzn7UKISM4
DUJz4WimognOm4584Uua+wHkzea9ShTxs0AWLg2NOs6rCFH4QFqV7poSgiaYVJ/pt5WTAqE1lNdv
wF+9+HfKK/6AjHVhYCW7fUarr+IZJM1jR/SYZiMJOK1tf3BA5n6CtOH8nag1DqL5Aj5Tn8tjkEYQ
aEYDRap+OuRQvxzSyyMMtno46N3865/w8bNAYlb5Xo9Ys2nUHpzWpWYud+JarYS83OosepeePidD
zlv5+g8Nza6ugtmO0WbVJJ3fzkIS/i8yTSjhodfgNRfiGKhIy6hrn1Eq3rNCGms0DOgGSU83lQl5
FYuNvymW8LLkswaI/FSbcj9MLhdKqjNtv9ZG1A62ZUhafQ4L7PcgXox1ndxn/E40EN+Jk7Sxhcd1
GIMYDggTVjwa5QlQmDKZsrfUWK0BPR3T61uaMjx+Wt7sQMv74/Z3dd3TIFWYhBakYmVcoxye3Ws+
RdBMahcw1pHtRHYw1FnMvOw5CMslZDg/cikC88BOyQPgqsaQn5QVkqc5DbES4NLTf8dxMaGIBu1o
bLAnfZJw5eFVTOR+PkfenWNW8xUOZ0SKNrX5OJEnD9nHqcvC6tZvxjKsbheb0219QgmCv7elSEq3
/9325seATmDzhoNea/9i4a+ytzqJ9rJGAFwWZjl80lBe+Ne/yEzDVTo7v/yTa3RT3WVuy+e2bZ9S
OgXZ6WMMGWcdqhcOZlGGeM3hpkeb4J2eLhzmFnXf9QsniMxySRK/9EL7vgb5jJbmntWG4K/ge38I
9nQr8/BA/eiwmHavQdW45q/kq3qiF2VWNDM2NzqPm608pGZGipMvFUAiRZFI9lfOmVJc1maL+h94
makVVePPPFG5gEGQYE9uPYSQgXf+GtKDsK8PhzYqV7jFRN7dN2ZcsAV8wIEJHytAt7TT/cqEXWe6
3iwyz49sgzkcP6PLhSorrEiixBf2gP0mfbq929bQBInJItTDRHJIue1J2xMT+oQl5viNnRm0utID
I4X1NKK/WoUXQyE/gM0wRrFymz3CcpcEHzHvWFprAoGAozVstviUKcoBuawdDf2Em5pD9Mq3/qKd
ogFFqMRSlUpKrneaRoQiH7cBNSRAEK9Tgq2BuEE1a7dgGNdkImoYGCGRxI4lIdDZicaZkbj9iNMc
lkwsSwp47mW5VuqSJPFkwUV1TlOW5Ao2EwCMpvLZyijIRpawF1ddQ4+BKhcwfUfHzpTnWEmzvnJt
6iyVNAFgEY8+iOy5VOGcgAw318QT4mh/xgzJ/78LixJt5UuOsTGan12eM32f1mJ0iAW6Gvd+XhLX
UkuVHiRMgw/KnP8+x2TktDtTgu2LPNXthRgJ8EZsXQFHOEX7aOnmpdCUrkuZeKaxlcAS+tUAj0UV
z/Od2Vgbc2fnJkKbpDNGW6gLawq5OZOTthQTUAAqdA/a+kQJgxYLhSkKLX5nuCzwZiMrlaKG9p92
cpg+Om1o5RCULrmsgAk2b3BtmgJeIOHZiciByWGO3DfI6b+4s3D52I+pgRKGavpTVljl3w/Mfx51
vr55oppNldP+5CAqL3B/icm8ga/AqlUo8cNc+yfUPDQlW+1uA/iGMxYDOwJgUQJcq+MMUHsFdXA+
EIHam0wUGxGaFFJBnZJIqTSVuohv3ye4P9vDGLjdlRKHQXCk3/y3Tq/z8k8Rsn/hnQ8sjcK7XywW
a1LT0U9TrbeR3rFcDZkXCme0NOeVWMPJeZy48tCWyn1R/0wgxIALa2CY0PLzdfYOaAaMNtl0ghAF
ILGPRfpU29gVMvGvCoNr4R4I/WkhFrro3ZLlQiyuBI1JAbusz5AyG8rCEV2z+8PNTdDY0sMoGWlb
ADUNgpNWTbFUbj1lSOnk8HU4unayckBfr56pWJk1Zqm0j3hapjr7R3FOM/PaKz2uMPFzmCYVAFUy
ppGvpMCJ4yqrng5TIuCXs80mwMU2HVtpsJL/Xm+pPtDclLxTUO/dDUSYTlIhPkW+IPDH2jo0yYiP
pIPB0m8l+FZ2a+bX62+zmjd/XQd1LvVRmBO1WDpCHYm80KeLy4oKfeFi1Ja8/jWiRx04jmflnHRx
jwgOZdsoS9/j/E8t49bCy3wZOn/yRuwvkNdfVaVcgtkU3yEnnWCQ6o7vvAKdYEUVbk7C9uxwbr58
H32KcD/cjaUBB8fAqQCUT40XGbK1Y9/UnSjXHDPT0NhW6H4XeZKZpaRbefzH2weKGAxrK6oOmU5S
0RYIPfd/f/a1FtIBEPzVUPIBDDn4aFuzN1TNnucbRteZli77thhUxN/aFbL86fdBJ4W5LyzFietj
7ra2IpZH+Vks1Ef7Oaw+6uer/txHz6xHpmA4xH9FmVd8d3u/vyqzWGgIvpi3nJE1CcbdGdC+roEz
9oAgD9etsYCKscyA1VVrkWYHoSMX0C+pHPiqwVmoAet+7+tDV8IpPHt8V+9KUFQYbFXhWAmcMFku
G1gAEsRv1dgjEmR7ZuPTeaz9eCTj/JdUCWwhqs88USgEtNIBxstiIadVAELhzu9G1nUv1SEW8ESb
XjPCJ2EwiJVb2wgdvywktuF9KR/0USnQ0nXOeyGN6a5egJ72BVN5TKIAUZgkdyc9cmEFCQM31JO6
QAdW6SbNGcJMCtVmT52tsxJdH+xG9iPyRvgSUI38Kg3b50a5UOAaXZCO8QGvPXjZeG8+niFyuxoH
cQjUthpM8kouXK1ddK/Yc2v83XjKK+fldcKmBv0/jvw1XQpYJt9VvJswaUk/nuxAaddSzw02Czn3
wEb8hJcWDvam1Q0PMVtm1D6NL5bT9PD06c5+BgRs3gy1CMHO1Pie98BLO1G3QhyFCAIB7M/GA+Ld
F4bcqziHqOdK3M3AgTCb8DaKZgsk6qOkyuepD42LxilhZqKziuG5bmFCMVeluQnMbVabJJ+5PPoz
TJDyAsrxbVplUXgGtJtChVOx0XbCUYV0KqheRh5adBoU4XffE08bdG8CD8WD4NCylKjWPyx34+2z
NY/pdHDh7RbdeR562Opp7YS+tVRnslyIibjUEUexAxpeJS1dhEaIvcYDJh3nM1Or9PeAS49WEbYK
62lCx5V3gy/5OQtGC3sjgyC7RTqCu5ErpLTejFfteXktuGrY42Qih66po5Zvj5sjlj6BC9NbrNF/
qLHxRc93Ch88c1HPUOCCm0NhwWlH9Sw0XfmUJ1tfwPTfjpl10kMDo1q1/F4FqgM+AOQZi8lFDtnW
xdSz71BW6HjB0WHT+ToS6MnqRhLyw8cAj/jkVJaj2ETYQiQTOmOZumjdKZQTp/1N749lvdbZHz4N
T+TkOAryfzsJ9tOBAekBtPRoXs2s3SDXEKqxRCb+1LvmWlvWZquFdqQq34Tp85TvLmBLU37Sh/56
o3ULvmAuFOiUhfGcptW+bwwJY6HZNgfx6OUvIEbrs/X2x6BbqfXlb5L7RX7vPob3ATmhJeNBABt1
DtldRJUUBlIuyeuCzZXbbH5XG+3m/qgvfIq0aN4Z5BP/kYjfleci1TkfELcS37hJKQfwe3aoH4gg
32wPEIX4mOY3SK8O/WxYulnGyQE1TrhEd+Mv+T4EDkpdWpw2mp8PhuwoL3K8WINqfG7MB38UUg21
pZWdsM3RJfJxBekn4Zbbb/v8KikGZtQaXYEHDZc+NBf1nbp4k399CKJXNMQujXDrspHQsdYk1lyR
GUyT7xeUaQPZhalK4+VdLR+tRB0fY37GgpF/7eCC0pdZn85o3NKk8wIKUDhyWJrGwzES/WXsyYdG
lYgIWRZVDclUjFuTLbtSLHWwwytuYrGZLqEapoi0rkem0ix0ra4lnwb9ZSmETjzjRnBeWeIN1mZj
u42EHEFS7rjam2xKfaDSHrMFyr7RMhUpH8A4gqs1MqSUA4wC8cjtmrdzWVjH3hf09O5ZULYGasVY
B/1ghm/KGyhlHnTLOYZsX99n1uYto6hDNsgD6poMiIUgG58A/3cFjJALHegLvF8upR1+pJ05BKYT
iGTQxbS7VsDQEadJIV6iR67FXW4A23JS5c/3C/feblaUgi8Kk9IMCv2G8Vyz2i3vtL5VKwL9DjZS
Ni4B/iDSSjFwc2wYr0XWDOKAr8DOFVyOEJKim6G7B4tprCs6wdEAzNTLuRW92/DWkWM/BgC1//Al
TVXXtqKZI/bTrwrMuPTJZauTLzimkNKt6DYNUT1HaejtAMWCe/W5mpmRm2E42dVa9awuBT/waJ1L
R3iLycLNcpq6sTwHrAL1dASTKXZnoweaA8Hxtp7iUgXf7h9FrwTbZcGqHWZt3EAZznBOH83VZ971
Ds2VbZkCZhxb0OycMfitByI4INfb2jS7c2Y3a7mSyZouaWEY0gPz8OiPQJUgfyQNyYW6o7HRHg9N
WlzkczQ2DKOyEkVaxr30CPDe9rc5NBmHMAfQkJPNuRNsdb3LjEVOP5L6nhtR+V9QmPcZfX5rBaJp
Xg41c7TFhTlUfJ0oW6tChQVwZqwlDKYEuAjTe6jjhzz1MHnKZ7zH2gBLvNPjEt7EVTQYmCcf1GM5
Cxn+rZpR9gQtuDKs/hxLd7R5u66ra6jwmYGkKQg2kTP/HYtFdOiIAWzBVk3wix3pV0LfQt8G60lG
hd7P6Q2dcQmwJffLYy9Qo3yPFCGhRf+rbwyJ/r6fo3X0tgdblhrRkh+B+gUvj3J9uxzr68Y3kkHm
r6gg8fXih9V90Gb3bTpsZ43tPWZaLp3OZo/8Co6kw++EpABytq4+5CPVxLA0Id/PxhGWtJPLwemt
Cbgqr2MKROod0alywWM8MkO5MtEbZlald2S5stH6IJXwtl1AHN7M7fMDz85qgwSGQZ75DLPIrkSB
2GLbNJC1bE7Ymxn4PT7+gsMIO2PHyONQAhyPZfAKnksE6AXqnYQU9IKufGQ4WrKKCfQ5rB5vanV5
kGNnlVktodL1heWmNvWTISTvQ9Sf84qT3cS5SOLq4rmyhwoVL1QXTHy4hL2zYreJURyzpXYNvWs/
8qkPq17zxbejv6lv1q+tMpsNut2ycOLvBYmSLtXk/9NN0GwfgmtLHC5N7booHszzB0e4FuUobKgL
T7bloqkWrB+QZ28jYipX0A22wqCS4nGLVqThwMoDWL4Tq19jJOJ92Ekap5X5uJfe7h3gxql6Q/YA
znKwp+vHncOBmyYvUDOaAAFzi0CkU2zyaG/L/exJpncbKXpWfyKzbYktHdE2eYxJlWH2SnEBJ/CX
6goK9BciAeY4W/jVzYBSgwpeC34zFRnFvv5Uj2i+vdamJ+QMMppdbFTgnz2KASPivi3nIKGj/idw
4AKbtXT+ykJyaLtOobFemWc03uLFyD8+ntSZJPSbcKrucigaZQVHjLpx8g5t+T1Zz79dtTnqpCte
okjddb+HPK4oV3Xkajq5eJGZN1pvXDyPfHxqzhqOEwXuoTA/eKunuYFlAOoZRKTKbjulIqwtpbuo
T75g61pmAmMfBbf4gmXBbagFsDKFWCbmNxMed+mTO44kN/Biog+tQlaCbWRAZV4n/7w8JOwMyGi5
Etkfg2RJlJi5mIguf3P8ZAqNcZfXbaeuu82NvdMOlWGwqvTkWEFQicdZNdc8Czu1ksikmUw4rA2S
7YXIp4UvJJT1Sjg7Kro2AB31zY+b9h6mob5Q5cwl1YkbdS4Y/ubqphJy8xB1IuFbcB3EZwkIOhy/
3VYpom4FXbTO8rpYXKEAWXVCfNGQyGRpcqHuplFwpTr766fjam2OqeI3I54/tAmFml3i2LMHvOb8
udnuzmh5JqPdvSHz00RJV/pbXNRl5fLMLKyPpYms7ZZ4VFkUsP2jkpb+nbfcB5pS7OxpSoNsFQxH
tHSwbKFaC/OwxkQGyHYXbKF04Nste0L7T3A+4Mo/Izcpomw2cCEnBzH59F/cHCbAI3rEuVwhjcIs
My7gEAR/0O0ycfFDJf4+xw6nBy50BGV4EOJZ+jGFwpLwy+zX33mIqcZl4wAvX+my7ho1utgPikKd
JzC2qPoIVOeaPvVy3P4gjjnPjNe1jm3cbdZ0bv2zGULkz3cL/47vi6AXQqsklvMKu6EFgyrFTTJN
vv4CaIqOu+cL9YxcNYWUJy1Fny1zRvPX0bfqYLlrb9GFyjXyDCYtrpEBjrwBcIV1Nb01Lag6z+RY
QZY5vJblxRcwnK/oXLSRSjYRZXE1EWIaqd3F6i2mAQkEz1H6XK1GZGIHDNQAM56QQK6wWxLjbm6Z
clnWdVTTOhKazpmy9Xkd6axqjt0OrOl4dg789ZQo1YiZrDnzzv5C2FFFln9CSU63g//7n+nYYj87
kB6PuLtaEUbV1CNAdD/lBl3Wp6PZ9ANC2vlf/RKJ/U8no9/Pth4vQwvLuSHhJReihlk/UHJb8wI5
9lmIckt21iz6mMQ1Y7NJZ47hq1iYNKgSlg8SivLgGcDWjgLrtlcEdC8Vexd218+hLuvXrswlw0Vy
AIOHQePct6usiOga23Pv/6STfLpNiySgASxXVBaIOBoXtR9xYN1KyTD/pT9/03bWFlSklzqmqJCL
r8wk/uQ/QE76bpPbS8I4fFhHGKfHGANRcEoK6kygKV2NPM1mQH9KDfSO9LCStXeLbg7FnqHi6CfZ
Bp+8pBRffO81yTwYniRwPHXwttheJpcPuucJ2vOk/KPei6rGTnTXod40k7pwUuiaYZ7ieIjezU7C
0EfLeUbjHW2DkrEGl3Iver82qguzQEaXwfnx0C3LaN29j4VK00SkGSFTx9oCfO0/vID3BaUhrIua
HoNnlwgeoIME4bxg/X1yOfFyPI1oDz1mFLi7Z3uXa2dYay4QGVtn9EDAD1XySt0YUPFj4cVsJyaW
SRTVAsNiUkWOT0g5C18Zt3MpB68ME7tEoqXIYCISTdAU0IVoKp2KpGSrXzk6Xd6hI263YDNSCQ0K
gJACiAcmB3w+PKeovMAwI0lAw6MQqkEn+u4r3Vpvjs9fvgMxvTVSKfnoflbXDrra3KCBlbiYyyjJ
7/jzJP5Ybc8ECfx1Esb8lUTm/L0Wkfv+rUIz0OgXliyH1F5j/2coztL1Puf2WqJZxB3whKRFqo1i
TbN9/00yWqMCtxfJYFFNW4b6oreW1yA5V6H2ac+tIv9I+96UY88ts/XW0uhJvJQkgbqGoCL+ZVyF
aOTtcEsUi6S8kS0l/qJutAZEN2xoiq8ZetsfGs8KEJ3Adbo0DW099mLRaXoM8aOvmJ3smsR795bl
w6Gb69ZcQUucrUgSwl90aRbjua0EGLR1cEawVwdCK8shonMG7u1Sf47B1j0TGSRDh/vBgIPZDX7m
dDIx/3y1Fjl9S54Srx09gTKA9bCXZO1UR86zKfPTXf2sZiIWkEHX2kkp1VIa7Ji+ME7pHhLXatnr
k2CfO7RqvWSzbxhWXINrl6OV40f4SLLpvCg0bX00t0BcQw8Ye3MxSZZAoP3k/wSqjmhBUaoEST/+
RaugzNO6uNfIJnZhb2FNhejLdid90inhuW4t8+0PWVAXMLoOBb1TjayYLJ1eNyJmL+8r5D0lg4wV
HyzA2DcItKsnZKVExOVsMPRwe18hfiBcOby18cjpvio0UG1vsPkUvwmIw9UKDugKJTvs9eUBl2y7
R9Uu9mar1gN3HKJ8E70GSkZqqK+KQ3YIqeJGWvtMJHjQ39lyrl71Ge+5L/sW2kqBTNpg9LMKulPj
zYdMHWS99ot2Hse/FUkryXGCFYQPW+584hi1GT1lZJzQViRPr+7UASDhESXCatfY6z+hlen8g5Lj
M/nym41dOw98tT3LdRxzIk2Va6E3LU9JdSWQNMvC+pCXXDsMpg/S1Gzmgg1oKQZTBIPe6Km3sSPY
l0TtnxTu8S74ZTH1MKCM9uIsGxMZPyclG/tnyENqk7NkF0mTW7qbl/9co0GHL32oA3UfHvtFzkLS
GSkxU9Osvud8+2VzUPsacFYXtMFQIo1khIfS3I4MOHt1q46Vg7A+guW326YGT0u6OI/7WBfE+zcg
lt0aIBWDrsP3ZOLN/0XsTSB/fxJ5SHw/KGwRDHPR4YUieKFDB1XVHvQw4IE2FYSaGRXtCi9zPL8h
MMHse8dGHqJOjgukfkhEGAHeLbJ90Mjka0zaVkG92Emvi/oBZFxWasJV47paRhzYWjABWeboprtx
zZS7Jkh7tahyeriDHBaeEGZwEFV2vSwZjNJxCCdfodq7kcDcg5OU3GyJCORxJ1bPdlR9VnLtuDIh
LTNK9rLBy8htFO5wT+BBd5OcqUGc4iLXc+6HzqhisHNq2QET1627ObfuD4LT8hLCwYnFDjhRhRoH
Gk13fX0PFwhuj5MbZxeJyYxUYA0uOwxDZQ5d68OTrPCezxnuRHXLI6kCh454l/NfFFVIOCmz+hvM
y58T1d1pg6E4J0lUigdQsvBgR8Azip2fcKODPIVU8WBXnj8Gx8b+Iv+lPCKmTfKiUgty54Pu6Bfa
L3ArMJlcyRNkL3qN4tl/X9UtPq5ZBmMuXWZkJttqXwnSR1IJ0WfwM/tGkgMk686wVjijxdCR6cyy
Ra8reLsHY6WYoBWDuEQx09OsrA40aMOeJBr4jdQRvxvJX9SnrT7/xRtVCX5YMoepMDcGl5C7kqsj
R1PYNdAnV1wpTBpC3W6JpOIzYRE13sKAateLU5YPitXG2r2clOiHMzUlTbUMFZymSjbPs2HiTDl/
A2CWqBCiN3+mVzq1MkcVnBeiQ8usUclpoHXbinBeS0d3JEA5hMKGHId9rlOsCACLCKlBXP8DByar
oEP0ww8qTZNnNQQy6E72qtGi2GeJC26nPXS0lMGH9K4/6EPYMOOYl0+gk9fX/iPmIsWY1aL0fdp+
arLAzh+oXqFFS6k12bGXIZlsxfa3zSQBTi+XkzbGn0v34tWj9BABdK2pG0iLEIk3WCuD7RxnR5Gv
W2eDLBoZLFGJl9YP2Zp9I8aFhguSaWwhN9M1mvbvdQxy8cU0YUR/b8o8Qvl1bLPT0x+YI2hwUoqI
FgqqCvxVOVE8c/36W+HtJ6TDqcZd3oXLusHVSDHgBMNFxI05giSXrKHAHhj+2F0MYV43eWgEZbnx
MEwC+MoZOqGMJCnIpnQkZD0NnW6X+yRe4SOPLSJgrGssPZh9d54uB0GXzNSpVkws8ySIdAcFP1ro
8ES6l0VH2CP37ySSkBYBYKFVL1yb/hhFVDSuNi3UvWRLGsK/n57uuVGIeKBgNZo5Yp5cFhexNLSH
HEm05enq2mgaDVGIUybRWU1Kk6yCqoCbOj5MjgeOGvEc9YAytzIIxR1U9bW8CbavdfHQ1uPKj03f
BQZmZ1wlcgBDuEbk/IKjholHF3pJcDDRhgvjSOtWm/XbHjgfwi/RGt01/UVvf97hRSkjQztdRrUT
T0viEoPrBBb1Dy9onOSSocBWIGz7EIZM0YXxI9x/WxSbYvTcof2IO4xlMxi2ERqs7F0ObaMZEZjB
gEa+TijTxtKa6nhW1pPhbsfgIGgespYBZ/QIat315clCxA4naBcrLFIQcKWbZd8B/n6VZ94VjWmh
0KdnDkKECD1N8LR8vhJTjt0jbg9gIsyJiZ22ZhwpkIkwx05C1o8SKb6Hn+D2E7a6n7zzdrzIlmoo
6oSVD0bdzkrbFsUFeG1a17edQbjYBYN3QBqKOwYjPh/wH1CfBf80+svFIygxwBOziiaLtvI3WYKa
9j5j7pUi7MmXGeA9O+Nw3YdawbPwDKXl4nzcEthjIZ8WwJOm+n7cFLPGqYzdcHEZyFjSIUE0DUuK
1++QnOA73GrWTIhBPewanTddjaJ2ITVYl1Qs79PR5GGiVTZmYwFKtL6TOubFsNqyBedfSRGIa6xB
GAQ2eC0A7NeCAzNmuVBIgwDX42mADYm/Goiu+IrJ1htp1+vJNRKh3+AfBS0Bklf++uQ610Xl8f+2
NEM3YsjwdhVO7M7fGC6jH1ULWpAn/UcNuFi62Rh2yZPTfT8Z4/8eQT78zGvroLMMuwI4sjUZatxA
aMfBmk9blJBA2KHIjbfvUZIPv/yadpldbfhTdoITznO7DbrYaIhx+G2sY8JIHR2fYg9k4D1t4JfU
vkb6dR3OQ9prPRw3y53FLs3gB34je0DYkjd6OEH+oO3GWH7TYGw97/Bsc6FU/ir7gsEOZ53djFoG
WMT790VXXMnKZ9K7PStWpmRSvO3H2TR3fz1ke06MaYQn1Z8zbyitcPdnPUlRBOBEMv5s8XjN0oUy
jBXn6GyXwP19bYfZTJHwfGrG3sYyeFTSIS8CedAtJFUKnjyyVd5aTUQ4PkKKZUcqwNKgRTlS99OE
9JBIDhcdPrw5VnFC6gontjgtGv0ql8dk7o7LEB1bs/Fti6GRjZLR+Qvb/vFHYmtbeQ90+dz8zp/L
vC6gMqiZ9zwl6G8jKoIuGOgB8z/B4miw+v3qTxn1tMoQx50WHC5t8AUX7yy2D5f4Vpbn5+phz85Y
rxXxnod1Q2XXlPP0N9qtN0Li0PP2vTc6PpS7dk/CqpbNCvohX61d2t66imJePib7xgIskJc2tTsT
ZLhXfuU91xE1M5MictemNgFrDK4fDrAumcDB4TqB4NnTLR02BEkZCQ3otM63C23vRoMk7oKNM12x
4fEXDRqQc916bdh7TBLPujIX6w1cXoMXPIqvLeMdZwINDI10ADcbA1ZW2mm3nYZIzn2Sl4T4XxaF
1izNIxmBcbqWAwVMHmBZdqglCEsW4QEGBLNWklzDEIksi7GDzGnMrjX/F6u1RPkL/fpB5FVuK4ne
MkndqJ1U2B0WgWwwFfM3AOWbHmGfhVlJZ1u53pX64TwnE1xyukV0k4qbIWQX+5nDF0FAQDjNRsjt
qTMb6K7ZPIe612avzbbfr4G1KmpUggP6okcJzpuER6oTpBNH6/r+/stvVrFLVID1yLQbqKvdvyhR
NL55AzJ9H4XNluUtKAQRD6Ndn/Bcr2YE0bNOUUXd8kOCOOcQANKjSaam/aLF60ZmMVjB//8qZ4bc
0tfWKDb2TyDGrNTV3QkAcevDgiPN9CXzgGShraXfxP0NrV5NVB1QRKSH93vb7hxActZIOyNnWoup
m87wm6QIk880kvNmiPsJtJJKmwdVNYtQiKLSJ/1CqhzyzE0G24JJNmDT4LSyc1spsf/Hmp3N8Cnw
bEmpz0VMzuANBxlppU3XfFGscXyg2psUvIU5HDxMX/nEaC/4UVN9D2+imd0vNxbSaUxwZQuHNMuH
rYnSuYD6rYgY0ZWyw01TWScENiZ9VYPeoS+LI+49ZifpOxe75+58ZTBEvM0RfCJA52VsRvlrIypR
dp/SNLpRUJK7AwEjDBKPmXqPcFHl1vQdn6iUJ5kqVxr1ILXDWEcsRzB9MWx5ECg7ChDLcoAJiDEE
VY6pHNCpveyZ3jkneNVcGAA0Uls6BjIxfUEtSEpfDQzW9F3tjDpFVC4x/y1k6OxPDmfmGfwcsMh6
1L7No6wv4I86tW9NuygbOZ4yjetUZhrgO5yurR169MgW71tOERw2m+uHt3oA56GUP7aIjozl7ujD
CNq3BioFJcwtjuBk8EU2xXXCipywYxBrN8gRqbT34J0GerGjq5OHky0PmjXwNw6Y3P+qPoCKn876
rWAnJ/FON0ScuzrE56F4AN0tcAUTmy8lvkSget4GpWnDDAzQ/G+EX1bypVW0OXVl8PSl7iLEfJ1r
Iam0wlWzZYoOVmG9ngymtjcIYKOl1V1ekOP4rryszUCgYlwYPuyPR3cn9lWghxUudOAE6UXhFRUb
Rr+ayvAviHIktvaX0eltgfKFJQGU5flRpcoXkNZPZJc0/1VeXyZIC55KZfNrwlKH+9CN1RVZVbGF
kqkQrB8TyZaaYsdrHXyzXYZGRmvtfB5wYuj9jJs8/354nQ7DIQD09tZ8ycByPT5QYeESbk4rikyO
T+SBvEkoTpgriJuybjKdfdi5A6SCOHvkBnU85h+oTvhPRbEb1AmrLYuTVb0y5pDU3s83bqKmwMsw
WJbNfWGtZoyC1rUPtjSJEuMRzWb5bImmy52scncTs6y8OkkVBAq8hMFvhWtzrRt8L2Iqav8uLS/r
LJ5Ynh3nKHbb8HAPGv8lRbZ7tMgav1eCA3uW3HNhmOXKauQhqU9xtGzyo23hDPCNlLzw8FSt1xnR
m1wbVA3X80XA73NfPdmGh7adva8RhXQPw1twkvM/Cy3cpTotM/ceiHAGpD/3mchnx+gmaPk8mlDx
3boBUT9V4zFcUuUoV7OopSyDxgIMp5t2NZHNLtN9w5CUPkZCTskC0YqfncKLMfgON2aN3voG12ym
IUfcuXs9Ojl/pwsZEcMqx/9uU8qY4DYQf5uJ+rTe0xc1Bz5e3J7MJ8zaltuGoj4qoKuNETwfdTGt
97lwS5MpTZVAJMlefZcGGm0Q/RChA8VGO3mLIPXaQcgCHxH5Mp1+9krA7VHKXU90oZY13pdEXTAC
rHfFdsE8WahFx+wQgZrETQkxUO1jaqJfZk1nwY+9aQcKfJZht2jSX1eQ9xRp8c8Je9I+De1rb5ka
JbHRLTcaKdmZaSnzSkR7QMf8frxGeGppmeHym3+tnP27jXJCt0jxgkSoRKwbp0XIj4E8TLboZc73
oG2cEUsjbKiNpluRAxoK/L40otV/QuRot64TvU440lTzIS29VJIuyrQW75lLvox0h6ZdTTO+IyOb
XAEX2LsIJUCXO499qRsgcb+FgqzBWPQV3AeGFLE+fyzWCiKF3VZQ9VQY4hMmrpbUUjscGaknMlD+
niZMQjxaYQxDPyfUSs27t19s4qj9xnNVukwNrPpaeAiVEtZ5E+eBAzU8+tUmvMrK9276brnjhqb6
TuXWTS8yKyqi5PSNAUeCx0yjdrqnbmRvNMfgUrtzTYdMDgLz4fUjTfcfwyR1xXi2u+l34bfh/PS8
E6dBA+VSjPVgCEjf9uPmm1qG8MlFdqcrZm57P4mTmeJwO01VNYO14pfcA1l4+qRNfaSYuvxkB7Jf
bfm+Uai41jk8xI5Ljjp5rK/FcPE0gavseHMmA2g3e7qHUNKOWEi5P/uJMpcJrZNNJWBGX4UTIQjm
3vOtvk/0Q9hRHekrPN2Lb8SEyMf2jM6KuWcMd37VdpGZutncRR48TBGANYQ2TQtQ1toj5ydHfVLI
DNj6JdYghpynYHV6jKNpM1BImwCqiCcAo/vb1d+WaDyDyHHqlmhHyYwY8egjv3h+CAGom3bxaS/l
/J1X/UL18sfbf+8c70wiG3mNPsS3tJnu4dIkvX6GllsEvfa0b0ktmwTp0MxyCFtlIRULJHoH+CFj
CIFXgT3V0G+4bmY0BHNs3WT6CUkRrfrNX7mZqOFuH+3HWI3OJeHtuUgcrJ+Fi5Ldj9N2hagunTGM
MCuq8VyR+ZH6D3vNdrcjj+pwmH3W0wjiR41McKCl9JLHbeZX3KWI0CuyngzDvF7Z4lp2B7z4kFCs
Lym0LRTVOuXXvTcEdwKd3AcpmkLrpEkObEp8wgYgexydlAkSaQI6Q2I8cBHQ3HdfGfbkU9ZD9eSl
lNhuuG+CSRCPbDzylpr7sPhXhqMpTYWfnpxjZ1KlAku4dVm1wGi9I1cGEI2LVICiyfwevLqrXsaT
4RUOUqFiCrlp+JpUpephJWsl9Sg7CDGNDb8LXOIcStAShN1Wd57TT1k0BCIic4DSXc8yC7EV3WPe
OV6vIFD3A7zCF9OkQ2u+5NbCR6ylYuT4YebkkO7CTUMlSYOj6qSJHJFXsVFqVC3Px4YlsF6B/KV8
d/pNzmCJYrmnUAWTivZeScYriocEI+zsctP5pUccNIfaRekISvTxvZc90uCeJOaV0w7LCZfVFeJw
jL9GB88FQI+Laeg7YG9/WtG6nMhnMprBoB6PD7aiQQB6dSTDnoSDduQMJrMthbgZfZb3yRjbkol9
6rx52BlpcMOL30LP6WiXkBEtbBHrQY8F7RmSRmNbRrnEu3wPIJdESfBaUF8ZxWHNB39VwVhTr0RR
fl1KrZ/6sJrL7k5D06Ln51iAIXGlsTbM94jXB7apFDfmnVCdG+FXwqiv2WxW4JFYaHHPBCe8e16V
24ttBwnQk3FbPf9h8LfEcIKJkhufJz+JGCoHkIk0/cVwUn3DlMNAN3XyMq/lAI5AXd7FFTND9h2B
T4lod5+kNR2KEiKfDH7+RIcL8UPYVAzb+fOHdjpzh6h8UFHCo9rXjLvzksJLlgyeW90/TEq6Vvkg
M/e0TG7thSlhfyVg2iFA0mlI7TP0yGA45FaEjY7W+eJurZ7/6llK6xWZPwY0H1MNmBnk46S4pUSZ
Vk3xcSlZB2rKF5K27VhQVO8SZqYQQjDpZRO6zyZ8EUpOYcIWEdhPQtZzGMnZVKmPPynN+fItKD97
ERIucDUy5kcv3d1NJUULWfOEeqrBzfpplOsP1dnH0xD0OBczq5oxN4mvENOntFVgamZowgJpVdtC
/maPpjAzAgbWjWug7u3es1OcwEdq5lKP1vf4wRUHJKXOkIl4Z2RrX74HTbfKqbCYDJlqUtAWmXBl
cqvXEKT07xJLn7UTWX9DFQOtY8xWjOKTKnSUoI+O2Nn/6FBL+Kx7DjHHpl9Pbcuri7sAj7Iwvseu
+fFWKBLvHqDOqxgzIVvIkGbm1rhuFP8iDRCog1f9wL/QW6lr8vnx7cvhFbsLtNNrbXlmY4m8fWoM
4IYn7i1j0RFJcFH/fS+78udn15eFRxHixp9SqnTIpWnd6TxpVWOI9ItUMJJ18/H8lqwKLZnPIanH
1iLBI1OHs+6a52S/xMuHkA1Q2U8I63P1gLm480/XVYQN1IUyuZ3bJIT0VdjYa0fPFXFXUVYzEiij
ozTPM1igXPM/oRjioYUNmjB66L2QYbmjfsrKq5Is9+uFHAzcrfvrt3X8CXoeI7QmkMyyRiMd7YIq
DVUqMS09OgP7P5pm62GyAB/f+CBwkbdpZ+jGM1+2kOgVFaS/nNP9ACa4HeQfzh69/rxGcxalU167
d5Cs6lIhRqRtyoNSVPpmjOfsmhp2vcM0FfwzH743qEt3+x1hB3USDWHtGTNAdDqJLvz/a6BjXWtv
NkeTONJIhN6pplG1Yb3N38C2F8OsSwhfd9krOJUasKZi3nUtFYJovw8KdwbR2ocP5wKImG/zgAz/
4HCq9BVvsCxudokKlXeldstXCBSP9gZcnw07pq5GCbk6zFeXRBxgZDqWPQAhb7UzvNnBhdt4Pvf7
pX3HC2K2X3c2y6FqhN/SuBJlSh6VaOegRUx3A7tI2y3ncE02g0wPzGJK/rh3722zv5uFRFRNGbzw
k4k+fk15jgsXUpKPazyr2lDH6W+IHje8ZmHWaMmAai9Kxz4YWDmzHDC1q0AgcoFzGDI43YFShqLX
u2hnB4adHcsBTPAeYPQRDGV6F7qlUZdvlc+tOIrvE4aOpdy8eEnG+WP5jCSuLIIyJtkRo43gsrqq
kxsJGokk7JIROGlQ+cKL5aAearFPsF0Xe2dyQ+iPIz7BKxv8ERnykNINyybVhn/+qyfrgfV6BWby
9CklK7hOm/UNEziMAlUkmGJuE7m5QWxkTtDsm15Cl8XC7FbV7Ne4O3Gdvr1xS64DLkmlEl3Qf4n0
Xb17j/WDNVbPFLSz0bvrbCM5uWv05tcMk/bNS0DBpkxVIC7iPmeLD8xXXwsSd6bEXxomU+KtHkPR
Ot+zqWPqi4ICdm4Yt5ObVMaoLr9q5QD3c9Ml/kRvxvgQPTzboay/gMsiqgfm2DwL8eF1hIvbkL4D
1GOicSt1d1/WYoWP89H58P05ZWn8aXqCsTYdQdSO+wxd8EjvjRmnGHLt4UjadJojS75pQR6bZFxO
3wS5xX/yBVjXkM97lWDxGhAO4rGiJ+EB8cwhHjh3DlCgikIIv/BrCS7JWztv4CR/JtKPj+NFIILl
gNEviXiuB59XbIvUs3WGtfzm94utcrllcF0CJQ0toIyStZx/rwj53syuYOjEj3XXwiJg2Gs9mLfr
vzCOeWg5z4tD2xKH1Rv0cg+7736suNVBRZq4Eyz8rxe1+t2u/ymy4YvRYnJChmBotBp8NGzS47VE
1SnE3R+fj8NGEvcQwqLPjTEmK+7/IJYmt2/N+FBdzZ2TJz4rkI0+lEZeMUlSdAgsqDMHcfnvfUcq
FKrIlZd2P/tqGlkNXQQW4LaKwBtQtLC19fs61UDlNAjmydAbBK7jCLrsc/5cP3bvzb7sDxjMWkZ3
Frq7F0fNNyFM6bO8nHjXIl5mjCExFMurTks2H3bjxO8/f3EjUvaFOGK8tXVlAje12xUHzxJTGdpT
izLnP1zJ+vqveX7RbCyqBxJY0icZ7RNPjOEJp/yJADLjL9N7+3QNMDiYMuows22eRGIq0oO3uASZ
Nrxshv4cUks2kKAX9O8fPbBpraeFjXCFcjQzZAjHKH/tqaU1cSl6LLm3ZdBqSYk4MKt7rBDuJj1P
0WHN0vz6/ulRldEo8o2TLtToBZS1RhVbSI5jyYhLJsfDg+bOu6duy9uz6Qq84OTFfEdv5t/bmhzB
L2GhyRiI1lAj7qkqDC7JfQmszOLsv/SOdy3aG4ds+94gPgW6Mgm5CjIHkFinUAcWGXtADFoZkuXQ
AGgkScqrFcMPH1y75oo2MhMXZ7t/V7pSkaEX4gUbH/1HR5M10kEGaVzsgibT/ayeUfA2jG/TQJBC
uyIAU4pay0LfarGW25VEOCf/pykta6FALv2qd78phsaw40Nh37mCFix3BEIW1IltVJWjcWZ2GZwa
nfhGP7M+eKbGTQouEojpYcg0TUWiv5AHegiY6PttyYtt+B1lCFaD/nDYNFVxnJlj4DzLZzj0gyv6
C5s4NZBeWbI0BR/UEoW2jRlEUAehoUxTBA8hGsJ5E4qTHLsyeao7tMDDWJycGAOTYT3GNlYvrdkV
xHbt5/FM3QZTX9ipxp0Rp7d+IjjjGsG52PZgj0NIaqq8YPtUWIzKlQOczok6ynFMu77Muc1SpgIg
sSGMBgw5knZ1wTefmfwZSyjN8CIE5GXnNSdds/adZpdEqkheo0A05K8GAmCg6lUk9rAuMHvpLLh6
FRqJOiH/tDTQmyfMkhyLKJh7lodOimInQRB69RD0KlFUoQC4w3UHGPzKyKNe+B6ZvxecLTh+sUnD
nrUcTBlEfM6PR8eRQO9YCN8hxSMIOXRh6EFmnVlQOIiZI8W3KbYg8bkuWBPYa78mZMdLv9NL/kZD
M7gWadT0EVERRRxPsdx64zoddfBb+VbuDMmyOCPvY8//pSiiyktzsdkdtAAmQfrUZqRnKgEzwsA5
WZ8vBut9w7tl35sNOPCTfQc1U/fSx8t+7Dpux1wHYPEHkdyr+KZulEa86xcpkAlnsqE7avEQZ0wy
1dLPuqQpRMTxrfZFve2+b8uBRpIl4HdfPCAQHWLLeGRP2xTtQ9YP/o1+tkW854xPC52ES7hrGF0i
ozvN2UCeh4RvcyDadyWcOAn/x/ofIJixuc61HOn13UjELEHSeySPFSdi/ptOwPnFjHP9G1nF6jM3
wSfsUwLn9Qqwdfo65mAdkjkRNJkgXDARo95ArFY1Qk5WdW4OQQmI2iEJj+hIu4QQVihL/ARedUHy
5JWWNitNNutkxV+iwv+Rqyk9InVTWjnmVQtp0IXKOdaVDCoPmga0iqkSllXuAo7Oqaq1DmzY9Jxh
/UuQDq837dy9GXb3N85+OWMTfJc1WwBKgQubu68ddW1VlNpxa7O+dykY9lGvEgNOtfejxndzAADD
wU6eQnI5t24KSZJ/ftWNMVpeXyM/fC7ZvjPqm2Sva0zgZlPBOJjRL1c7KDNUCySNRAxNKt9Vp+7E
bF79gffnhTc22gBFu83PttDxEWhN3MnnyAg7teLuYsjn3DDgqjqQU6M8paD/HLtWvB812Vcp1NzH
z71+fs11P8USMSVwiyH+Q3b/G5+oElP7EjXybZ70TKhWyFAbwaksyeAJwCzp6jDSX2kv2UIAjGR3
zifGdFiVrityOqtHaVB8yVcFIopSWXwC6nZsiliOeVduhwSKiAEoBRLxaVTlWzZ35AXCEi7d8YSA
/i0xMrvtwgcFMk1ozwgGKfRtFcRBzn2gWhOW+99GVoVLIMuyC42OM8KHLQ9GU82fbOqubI3n5p+e
J4DS1hqmeLGkBuZB0LpqWaqEiFvUit2gLWdoEQN2g3ZcdK/GFJ9yvwdPlAaD1whaSvcN6g3neENT
JtZtsppr3BP8InCI+eX1G3TiZWuqk+SZjliaC42cgU4b+PgXeC4fiKaOlXZbKyDzYxONw1hhpHn5
KgvzF879C+dER+jdKfl05SrzqALJ/ah65ZEuXC79iNUrkgZlsB9TK0IWEmRg3mCyJXdRoITqLLgV
CtrPKCN3uCyjUHlonJ1btDyegxZ8gb3MqnWB+V8kw61O+EpfSznTN1L43OxSc2GR+o1H8gH+1WGQ
oJxuIs6B8KGQ6BnQ4cs7D+ymfMg13VbBm+L0kktzoIDYcgA6SktQfuZAdXKgkkY9CGx6WZVK1K80
EJXCBIN06bkiKX3IJQcosMeV2iA/b1bXqOt+vmuD+zunahslL7kUkvkcfjdK7dczM+e0Sy7fFqDz
JEknZtR1gJQp1Cj6XYL7gu63NuFxeFjChG2gdZBiHi3jqChc6MO/WiXoHcxbcSHslxyrROTCmw+s
3kao1mw/RrSwzLOGmP5Sf1RONW3bvFzcyQaCBaAslMS80auNeIsDtjwWCj4oUES0Nom6RQZxcEL3
GMLGeBrtYPyl9H0xjdG+iI5zXDrm6SPRHiM0FPGqrOpIEVr75sinqZC12HA0Z1f3K3ZOlIXzuhJ+
ApX0HGNuwr4DIURDuSVlNhZWtV1xGLkMbCrrCz72Eb6eGTKlsp3PMG3RXm18bGpQL7e+w1mMutDS
lXkWOUrVA9kMfaUKX6RnljlorHF0kIV/BlAOcxOHI8T2hn2Z07rbYNZa59YnKhXYf2GunMsVZZtq
RLFgcPEEiPR/3LF0BJr7E6UivAFrPlZ9VuFdB4JxzzbngycIIbThiBN3UcjHJHzG6JkJkgC3YgdP
M09T7xwOVwpLQN30TVIPvM/3H8TL7G0D9yESUfoPs8tk21VW08Rn2s2CRTwxULy8ucHw91ZuFMBM
MsR74NVW5nVqIhEeok1r5Lqrsqg+8XrxF+44EnWrw8idxnagLgvWm/yMb/feeisC35tUbAvX/e3q
G83j4739bbRqkZukDCyP60fPX7bK3VdazE2wcIR4dXir9khZ0mRprlpvXlGbN659KQv/4/f9aN9N
lO7P+pnwA0sE0FxPfBUv1aqt0rW1quHA+IrITEaOIhv6ACX205K+56GSU7D7EsH+clmfqn1XVeDw
HJZFcZKgd2fHvRcDu1W9KtiVQqrR9xSg9rRACk5NcOuUGwAcKpaIa3ojwDQn3YBbh8T4AJ+CYRXp
t3p9dgWqvH249/xu46dFJ4oVV8AZg0saVssOdnk72cQfSeXXu22zzt9RccBipszhZGLHoI3ZZzJk
BTJcqQRBqO+h/WQk/mSoe/Itb4FT8E6eJUT/ocJNM4Hpgm1/rYFiro0vxfsmG2tb72w3mKHNlbZq
M8ttSVKrbhgSS3V3fUUWMLdvYTjc1jICncBJuPiktE84T7Nb6O7sDLqVuMH6SLMHxdvPMqGw3X4w
+anrWG2My+Jp3PAIAAQpCOebiW7/gCEnOQdo4/AHzsislhNQa68FEWf0xptjPV3XlI9dgbr4DBcI
Ga1ZHDLD8mJSLl2jlxNQxd07HautdbBejnT+l33ryQoLlRTua6jtN8OKZloCDwKBV1fBFmvHycrU
QFo6yo04rXSz1XDaYeAyI9QufbCwG0QW4+6lRd3Kw2JpYhrHQSxIkfMbJmHLUT/LXXvC+nTugHRR
Q84dg4MslfoRa3PfwO/ZFzt+1lukAmNxhe0MNhq+ztoCc+bu3Nq83FPPUxdp5T4WHVE0WufM59h/
RJ5/0ZBkQzplTI7iUkqNJVaJLtpaPFFbpEroB27omzIFnOdMu+kB5uIm0+jP1hIAeeHCEyeecRGY
XB9fe3Hn0MtcO8UpjLsw/ghZwV8scd3evAvhc+c4FuJX/kazlnl+en5xXhUdjUW9MWOI3YbEa0UJ
/42UUUPKlcbmdXAGV7vG8l8W+75X5gSSnMusk6Dk4OdEy7hdHT4IhR1kfuozar9ng3KMSnZiuHDA
pWR+Ag2DFt2EfK1p3L+uDYhHp/Dc+0DStdHBnkxwdHMtw2LjC3b7RYgKo4ODZONiKKMu4XJx+yxY
++mhb5WqDqN0yuk9wooo1FtD0bxUr5OILOhdV7E+Hq3IloPTStsH1c0bwClfRw86Q2fzJw/DcxDU
/FfG2tgiESTtz44CLFsV6tm6pXSSlJuoXT6U8rUqbN1nW/42JV8dx+pRTyP7msdV5SM+wD6OG11h
UZSqLF8uytCkKS/fE8L2LSLg0y3JQXphoIm6p9Ot3K++n1zlI6p1xS+Annb3gF9fUpKWmONrRemX
+0ZFr+EOkyJn2OXk7qi/8ccv5S7nm3kg/y8Eduet+8JsvfniBuMln8Yquik1Yqzu+YGU1Ei4zY25
TGbIGU63Epck4uA/ICDLAEVD3LQ7k9t9byby4qbhzeIFrAzLtoDtCqDCW1Ip8+R2xV3KQRmglp2f
3KUB16sawVWyrIjHp0zzRFdBZKKWUG1uXI0/7qjXpfULp91Qsnst0vIyFEJYK7pwZ55TP5ZaBwFV
N7zKKLxGUS09FgTsS1j5YQF8kAbxuKBfFrgNyvr8XZwvgtk5Avtal+jLJ5jR2KmSx4eFFLr9Iezf
KrqM+YX7AGFn/m3kSrnoXDUSxF9D00iQYxw/eONLi2KVhJDfvbTwCIQHo5rq1CC1hHW0EtCjP9dl
BVnD6MpyLCgJZcn8uA89xC1x0tEjGnQm2C6C5yjj62hTE3NtutDLy8AcO4qRB6vEAoBLbX73Wh+V
8qkFWGnd1UftH4G9/0CiObRNRFo+TNyr/NolpSG/MBSaqoLpR9DNmJjNewR3oHamVo6IgNU4/w84
IgcqNq2TCnY0do6Mpp7dHxQxyTS7A1sWSAw5xnBc66IQXtxYtIKhemvBtKgH7hKAO3qAMvcdqB0x
JTAVznp22DWOm16xPb/M0rhCyn1jaUvnlOuL5netYCv6MaW8SHHRZJOc7MIZmoobkO3vwMeH5O7O
V+lbBR6g1mayWdOdm1c0X2DovJEr/LDkLB/rGHVPSMp2bRukS4eJlfWkbCrOxc5SvSuR+Pu7wgYp
exBRm+exbi98RG9Cq6YJ2zqoKIjKA2Klm51C1BoI6ko7YVf6PcuZTYKAwJfYEgWMKOBqSaepYB4j
4Qhz4nlt+YPYnPBTU61GCk0Mfqw69TvVgwlnIncyMBqGGEYT47T96D5gmmkTNVVyIGuYAUW65iqS
UiSiL6TDf4an8uSzk/xmGBoDkMGlk7cBMIzFuqIA59uUbK+TREQXu5mwdMOBhgry2j5STHUBQeuI
ixvnykn6mb9auYy/VI6Y9iPstRqvK2iPKCyV/GSVvcusOunPw0Nrk9adf+ow1IJB6o8mO6uBoxAZ
jVCLW7J186AafQgw2ZGYDt5Y0RfLcXxMxmalN8knjDKFuOcYvxKGXg5dTcVU17oM/4updAaHru+Q
FF3elHr2OqHRYQ6c2wyF+S5cMX+/MxG2EVR6/qJpZX6pLhpSmZTt+6UV81u3nvQYmpL0GTHzAJ6/
VVq0b0BQ9MO9dPQO4BTDRpSoAWqdmCGjm3Ifa8GG6ucV6nXCUjFsaEXH/CCWZZEuha5kUf2LylKx
Pj1uznSa5q5YcJm6P6BUYvjVlYkdNxcPrCNS3lskSXcohycPxCuVSRlw/QKCboHpTCoFFSqu/Gec
nodjFuE6l+iRJxehYE9IthNlIpoMXnpSzGh5z8OcfUI9uCCvm/chsdfRM/NfyX0uxzpIPVVTrKoY
SBUxkWx4lIkI8qt/LafQ/8RF1OCwi/+fMjWBsQXMez1MqjfPtwb+dVFPRVbeXmQ6Q5kZbumkndN+
0ASRQS3tH7miGQFhlsnidcejrhY/cM3OuCcMTky99AKijYag9Ln87bfUTsnI3j+6trTBsg6ctnGA
vx9jvutdOmcG4DElOyUW/sA0rrAuOxsbOEgDT5ZLJ6ER0O4A5MpQD+JY0LMlASt8VGhkTp94E+iy
EVDE+9nfqkUELQfZC0D8fa4Vadol240nXwVnybB0GZ/VJgc7FKGOKnkOSwzDFBDzA1PbP5xqtWNq
+W84C4cnvX50F9qNt9a4gxgCqQkx/enzEwRVR0ZHbqh/27XbMDR9XdR8yY/4w9aaF6byq8DQrvvw
biAxKaIJbYG9tV5krCszywmX+A4YpAUokHFL659MWw9RkM7y8J6AgRBw4viib0IBzKWfZNbYi6NZ
hZUlhtkakZ/vUYuKiFnNQjTPUbZJZ4n6P0/PY+IrGDS6OpAu0dGDpa6mjNd9ggrvT6V4PKNgXj8F
l8QNQg+9Kc5Mc5pYgkt728hT+iqkg3m0GJ1rHz4viQKLBEDX3720aIpAHHI0btRKIoGKj76ecFLJ
+sNR6SZVESwofF6geNWIrqj7h0O+QcnH7EmVnkeiUrDdC6DXXZvry8/fzI71ZZEiTXwtfI45hcGW
X1Vtnriho79jQtdji6UhUdHoLoA6jB8EjBFDV2+9nPmp7xgyee40yBQNzh8b3IF7h7TAj83qDTx6
YZJyVRKDG3JUYix1EEgVHsqIRW02isIti9Qj1dqYf7DarLQF8/nceBuT3mTatfquR2jgFOb9PmWC
CxIjx6PsKGqFvY3OLfqhIbplFfLLHQtlrG2mxmcJDglTOs/2fKN2mWRuxbhe47bubSBCTczrd2dN
eUO7bucIFb4fqOT3Dk1GCI+Xe/Gi1fHAZ4PLxZjSKZdhgUTx1Du1WtFQAli0ne2TudgphXids3QM
x998nY3qq77R61lcy5z09DBT3wZQJyDQzUf6mUtVAdtMWsSayWjuB0c/PFyq3kJrlim7zex59WPh
mrc5fPni54+MYWkRy5KzzR4cyYLgqr/TnT1Vtgzdwm8tjb6ii/Zi6NcyjWKd5RYLoMUDyCy9pMh0
7cNER8E/tvH029EyfjVIyJDt5XN9jpzY2GrexZxcQQ6moMqNQcRFfEoCUeI81y3NhL20laUIhl3e
uSUVhsryA3APIZPB29p579FKCSKWKO58xjOV/JoFeyWpVjToSxsyMWvAYEqi85yTqrVPvnD7JpmG
hopT/CJA31WPQI3wtZ/CCJ243y/FnQw6+n12VmGxCHZ8FaAAf79uzG96rI8UqccQsZPv8uqKA+Ea
pEZF5LZmqVnUsAgq6fsOHGOIbY4TsgtJ/9s6E3AqYFz9jn0K2V2Wb/wVCGt/dwzkKICaeUhl+7NT
Xtwpk+qHZnfkRbXBKoXIvX4A/5rIPjwNFxaEDITYITHc9P06Difk7u5QAldU6J110CRMxXa62/RU
4bR22/qCl5HJ8r3QjlgvvYY+2nzVf81cF6X4XiQj1qHARy9a/Jd6pCq4mTT54BQuNaTLjZDLlEat
1ICCyXocg4wS+lGD1n7wIicDI+GxBdhTjpLVLp7Cn9ltC3OMoS4ZQa30i0MRHtMLK0aQqZ3mvyC2
KmiGCoQe6sP2H3vB9qTLM/sGVNYPWvggdMhKJdO9nJDdRCZfTpX7ZjyousGvAkgACk0xfU1/susj
y9H/MV+4ogEwUvGjWyocHrBTpuXvErh8guYqa+ljtPt6M6xbUPLZa/LO2mviQZRMKVoDAYl6Q0bt
uzCkUv/HpfCk9Cs4TsNZlF6ofO1TNBJmqoJVCYj19ZV4xoLCvsz1512n/M2aQDZ8d6HoMUse1xr2
QhUCQLLgEAysO0VQIyHB0vuRnwMf12P+KZtfcnj9whEg0XG/gvEQDq689n6DOwC/mi5U672vFhov
B/cqOaSDa5UKnwpaWcM54ixNL7Lh7IJSWBc4GqoBTH4EiEx3kcXhK1tCBSM4GsBSoS9mYemjuuGH
le2VtYVX9B2YsrYdJsUniSbRVOtSqGD/5E4R8MjQ55Mb11x6pJYH8kdi5e9YVdH/idZSARhUfbGz
fAaS/8TT5eAFL7BN8J8h/DpaoRRBHTPnWhIiWzBzkpK68Qb1M6UZ7t82p6VoUgercxheHo50RnwE
PCNZrMsieFdf2tcMewtWUGA9O2OMRCsfl41B8FvBUFQBharY/aLKvWlxkF1RTBqqpypyHPckDWnj
8uevKHPsE6InvbU8p6CTijVON4D3FXQ3KkPWaa9/nHumk+hE2k1bYaBSVlGC6O2Ye1ajNSLNbU2T
4RtP7Khy77WbfGH7kOGAyFFnJxf08sYCN/RetiAzCs8pLF06F/+ODxHPvsxMjHE7ipo1eSJUHg6F
Akwhd3Ad5UCEPYgCpfyBM+k3Xjf/j7PIISFZWD9ii5+dd0jTnoUFMMBhMkecDvYtHiJtK5+eZXls
iUT9qQCQ0qy5KVYGwHqTp5Eox2EjjXIYU7iB3Nr6iNd74WdY0G4ObBMCRn6IjNZCKMlPCl2NMRSh
T36d2EK95iQT2nCXkl3EmessOlOnG3yoJhqtUSgjTpow3HDeR2Fucyg0GbkERNdHOFYY66vZ96a9
Qh5OhO690fX2sU16Jt3XSq5I/8UexGmWi2N3En+Mtt2WOiB/EkDGMy3N6f6+H/ij8ZqOFyWD1/Fe
3pAzcvY/pSNAo+/fMaQOkvM70EpLa9NV3MKzd0fF9bqEBcJLgkaJ+kKoxSrZLpzHSpNpGPFTcOrh
fGJ3MBvmXcBLxlZueygAmuSiY2+Q9bmbIKOUE77z/z8qabLmP5IoG97A6LI76SsuVB2STwe3Rxit
0CXcEmcQgLshlri0jTLjSmojRFo7dfc3kFann4HzUVczQRKEpsoRU7VF3cPQI6wn74zzWpYCkj4J
cNBJIzOQ8ScTYqng6htBPdCDygQ7h2LSXoeimhJTI+VEUBYeOEg7MqWelDkJrvh6PTlRa7wF0neE
6H6AqLjaHKgt7mYJAbZWAjw/f0w1PwdHoO8hY+aIcFK0+mee58yMBBhvnwDgqHVLmoEvIcmDbIkb
QLAywYjcFOvHtTXlhyPiv6SnZfMbYaUUh6I6oxJEtsctiYNP/N41WnqCBnv8SKvgws1+e0FCmLLi
AYm7GhgcyrvoEKYRQ4H03BynfMtwf42SktM9e3b9QUD48qgtCtcYmAUDRt5TeJZIKMAnBUiomB4+
Z3vjTEXvzufHvo/PUEUElL2ndX2isrAFSzF3hoDCkb/arsJoA7sGvQ9Iy9OXRmPt2/NcvbnfzyUO
KtVvRmg99MIsZa3tz964G8DCnIOGP2yTAd/71UE+UswOo8N3R2l21TgIe6nfs5+Zz+Pvc1gTMZwg
MD2+BDx0ZM3sy2he1+KxtfMsCexAUfH5+RxbxkK7fAEHVFU0/6onLoiXI+lH+UyUqTe6drdL1yvN
C1+/s4Liq/Bay/EL6t4id2zsWOCbxPYvnckY4p++fSPqK38QyU9PhXHx+JLeVfn15sUBqwfX0+Lh
vlbXsnU0fGBcHocS/N+BkQAtSs2swr4uIJ2vDDJt9bYlc9uVpqi8pjVqqm2u/hJCj5Lj1ZzxULjW
NmXBPRaavWLd/w6m/WIZxu681/GDm0Hd0cKuPtpZd6AwKpPhdhtCmMQK9m1i9mS2HmYSqWHpbpEb
dgEHNXwqYEEWDxdGkCizpUPSP/GuCWrgUReCKkxGESVDihjCvE8NseLhjKOPhQ3mLxaGpCa2TplW
MYmgHS7+4+BK/q3UFPYMQH9i7Lb1+URIv03CHhOnPLzXI5oTS0e1fWlZTxonUJ+hJxEO40HbWQlv
bSFVH3MfoagCo/6++DJzGL18eIOdbt1MjauVZNW82pt360IbgoY/9mGxjEUXDR7QdAVDKgC+nTBx
AFHRCuJwT2smcLJLQ3BtYYpa1OTASmoHDA4IP8FSlFtLsck7PzxfpjcDFPRuAe1XFP2/4TgjLjYf
RzbRWeSMvWJ6kUMaAaVHy4PCHKHStel+E/tQ+s50Nrxg82j81EHwuo/bVkB6JA7LcWIRkzlJnSID
pYGHdP0G8wbYsCmfb2z5a6/66DM/m8/67ZTj7B8T0VqqZxBRtYxCIsNEKeVM59nZN7s9TQ/ZcKgi
HhK3APo8D1B0ntSxVZ5jZp/AwFk1bAa69Wyt+xWOlz35xfnrBvik2di+uKP8HMKTOw8/d8d9oHFu
g6LibsLHej+0fZGvOV07wsOCVjEXDpsRzbV2OqhZ3zX9GxAkn283lKQlIouna67HUWBSjnMaBjrF
yWT3oM4JWRegGD1O0b2GCuuBvMI2XoJQI5rkSVJ9Mp+oBXLvps+ny4PCSN/ymOKPMnZES4qHI6Xd
qXRtokXhtGnIAl0lpjFfVuvSmsO6gsNLwjS8rvaz0Yj1u59RewONW+/rN2uRtPSkjnbzzFop2A4o
akaQte7aAF+oEdMUjZ6A1s31RmcHoILLlwNhunOr9QNknFmQZ4pCWx+Ax1em4KJXy+gYCNd1pdOy
rYvnjn7DXaOlBapOe/ZIybtcH2FiA+CUOsiRByon+m+zAjpaGjdng6U574/hG+DUVHlRiZEvfT6P
Z7NaWeNPxf8GqI740pdml1zgF+zXjNf9G8366qQwX3x9YY8j5l6n3H/jQnZoG+UAI+ZAwAhF6B1H
ilBDwCzifC8rvuq/S/eXywV/rED52geDSKiWRKjb+M8zML8zsUAQjDS+wIWfzvKJ+WbxC+VpY/rk
IV2buwBCIpLwu6+9gQZOdFY/IXWAVzRThocq0OV9xIhxFEQz4zVuC1XyqN1ZnNOUADWZTynvodX9
o1R8UNIjOeCOofnjOSeXSrswNFFdjVbnJJv4+HHt4szjJ4e+ZXxZT7UXU3YhS0gMQwhGzOncrlpE
6Zrjwd+B6OfSMcrjqlpj4sL1Gd5ihI8YKeEKxCeXQSollEYXcAEWd1x7CNhAeA8qSYcZeDrAq/RL
6yZEkvKPxi91P+OCfIyLSwitusBvTfhIjJXUdvekibT2PWSiJcQf2FH9vWzbGSg02HLExMa5UKbH
Ou5P5i2E4qTjR5h62R+wSylFC3NnKN1nO9EL6URfcAgWFJouEM71L/7qUa2njOSb9MYkI9CKKaNg
PRyILYtzD/VMtMYy/nWUxV+VmAb/k9RDHSvaCQCYXdLo3B7+tKwOSQOFLZNa25dy5NIqDPlc3Yc/
WlgQS/e5o+pkjOdHT7vBemmltwk+hWa7AX+w+AlYnZuv7eXZKiur/ujX0Pubp9cfF6d/t8E5CYs9
D1XVV+Amg2nE6INGPm3vUpJJID3O5vS69Md9GPiILJJMPNCVhX1PYgU5HB1RKNl7ExxmdJLIQmGL
vru+ueju6HVb1hWmRfgLzjh5WR32CP/f1eVu7CMwiKtpONa1nm/MDK2YQ+ABQZNOqCfl/xavd+qX
W13WWoIgAKlRNJDM4lEwk6j1Ri4guTKS3OqFiTEmGfbdi9ug1hIUYEF/aHEySoV9ofEowSZZdW8d
kFkSCViY/vNYiO/vuLvIJUz9fnRNgNrXHgrKluIQ2rjavbx/JplG/kVEL4Ph6YY0e6LIrZdmAM2e
tNGC+VGYEeSRV8kqhBVEFTtY580R019/cPinCq0a8yZbkQK3w1qzUoCZKMRbZj0q3ihrhPCzcY3P
kFvzRXDz8qkzv8b3xQ3877Rn9VIKetPFTTCSUy8ixDegzlvfGpaCWKsyVrE88UPf2S0hcDEWeI4B
Mj6/wNFQ/eDpVOdeX09btiTJeuwCMoQkFbidlx83df568QXThHdzCAETx7gGGEpoD4yASXVkVTzd
78JvJ4apOGIm2FDtOiD73YSjqYljkxHv67XlT6f6gSSBCeT4JLYBx5FwqkuQHpi4+ljTqj98Og3d
xAEsAhe5nDsk+VEGWEk//MOynUjuBtz2/nydMDA3ReQErB66vSiCp/Mq2mFBFM7kadqmJdB9M6jA
qwuHyQ6fKIYtK+IbTppQfHqPtfSIFL6AqRc6ljr+2RSFW7Yok4apxVMnJcFJoNQ+nFMj0MGZfx3B
8KrUMdjdQaTdx94lFNuvh+STErnlwPZALhRYH1yNzg+GutZ0K0UuMHIUX/4NzPP3N3cSHLvEty51
Zdv9ZH22Nw+lal0btN5mmLq/4bab4wD0Ksomv9dvZhTAA4dIu6/JNZgykU4c+g2bKBhQ0UJWJ0e8
10scjvKCxnBwGjzC9xxJzK+HwQSMUjIgum+HZ8Ad0uNAO3DLd4edjqrzvt30xcurjEqTqE7xAroo
eNwnPU41e71ie0VKYIBEIqQimHATQr4XnPH4J80R13fbpo0KhL1gNyEqE1yiHl6Cl80LtPJ23cBz
ePhHk+aPxuayi0QXkFMaeZLI3ZkbFxnhF2gImJ3KaKRVDxRMT4Erq1IDK5/mcKpfWaeeXQARj2ld
DKWoVFwpSv8Aqm+9hu02RwMyRKwI4+mPqD2Y5S26yO3MGFnIBJ8n/tPH9KOJMiyIMJBmeFRbai3a
OJoBS0W5Vv6IZgYzRX+FLiXemLMhOqyxLbxvRqJw8SG2h2vumkbuBcU+Fh8jTaSeFnwADEtVsItr
yM3BUeezfhas+uhZ8Oujd40SzI02rZgu0urfJn/VCpF4fUK7c6QkaVzXvfDtO0CaDmc8U9bbNChI
AxIuiqUysxirmYXvqz3G4PO1rJGR/6JGSX+atLcry2+B0Y5YHIFT29+mx7H5GR4g3pgvRlux+TzE
E+uaYrb+Q5OrBqg/Z13YDJugzNYxU5d8IpzRv4LkoQxKWMtzE0zhbtTRQ1c2lzkJ6DayIZaFxjfh
SeztdgDKHZ6+wOzyESCPxyqx+qhc5shjCt+miw0XBcnfeExOZOsV7yqm4K8bSKGtuM5gDqDVJLVK
+/rpttUcATr6J8CsqGcHOkTHCI0WYYUFLOwKRErfKidVxfC0SoPA9JcHwS8p+CIKrux14CQPQhpB
k2NABpXTYBVi0hlR/Ly9A4jBDlvQwRHLX5ibjwJvZShPGciNqPOei3tPzw89mr5dU3JDJGqm0p4t
oy7Blkg3v8Ytk6YvQ1tILdpO1Edue9/JxehBT6lxhsl7NbcL9noT2eyMFtQt/7ipcbceu/Pi4n4V
BrxbiOytPGgsRrut3D5u8FFxgVzw4pLpMbzKq/mlNZJM20K7TtfIPTAgdhsKbzut4IqMEKaNR6oL
WALDB1a84Jjtjc7l2exGsaCVOlLMP95hytS4XAXK2K5R0PLRapCfcMHk9ZXoBaifXnW3WElOURhF
MbQDvY8yWGoKVcLpn1Ki/yZGYyY1w6iLnpSsz68ZfFEchALRxOOat0AGPfE6M2sDXtuOgipIt1bZ
/wNUx/K65nyXgyUmV23O+Ms70xJGdxJ9PTtnIe8lvPQW32vixxobzUmWYRQevCKOnVm+Px6tCLgO
haCDrNdTX1I+UHOSVWDZz00y9VAfms7gs3pQ9cYTd0DN30O99WKpXAn6UzJEQS5fnliAdTKkR+//
lAXfNsh3UPrHVBHwuNK0nGB8z82Lek4yX6J5/wCP3cgnP8rL/+B5yEUfwAUZWs8eyCcVF9KCK0zk
3axZvHWbC5FXfZf0Vs9v34BZAmi1cv2Igxvu9EI1hAwx5NX3iDkYdV/YkFjWJ8yuUnZj/RphCocS
XY1/1ODFLm8i0JwFQuRU9qTRehmU3lvyvL68E/QbkmxHAg8JwTOGjGv06NPxpamRAccg7gabdC6m
6CIsE4pm8yPQ5JWGmUb4qXCS3ziQ1xPmEZjHCwtsGvBS4FPh54phUKSrInq8elBw/4MxQ1dJ43ry
Ni4y57woxALeekiOHHGlq2pNgsFT1UDE7o2ZvUy8LpSX9R3rBsVACvWAjP4uTlMdYL7/7k6y14cw
mQMDuACqkhkT8xLx/Ay20jXGBJwzuGFrJ6N0YwMv0EbfqowfbGghXDIzjk5XkGVB6GrIDJfnGJnL
gsaf1y8liIQsLZ8N7uHJvD/+yltA/wj9//Vx6nbZZEPuXMb9wrZzi7aZDoW/jcclFeS/qCIVtSzU
hlTtEP04hraYtHXHXpDCcktgNrjzYxgPEES8ecQiMSsxrZQgnOG8LDyntfiTt4l5q9IomyB9JM0d
0TQ7t/tSjGlN1SL8YPQbJVtL8kHqqkdVaHm/vkCU1xOnD/JXhWS8zOA7YLHA6TIoKvINRaFxOvxa
TG3wCeEoQ2Rd+IsGdOcIavl24Ra7eM5C1SfPXetBvp6Uv9L9X+z/UIs2bPub+G6F+xuX5K1tMa8A
oj4wkvjLta5aVD3CwgGqnYyccj5uf+Rf2A8bKee+hLujNDmnK/ko9X480hJC6ukLdXEQhtYzdSox
RffiFOTsYPmemwp/iIX3OTLNNZc7nw1qVI1TE+rXUJ9thKpUbTJ5Cnw4T/iY4pQeXfT37lTwNDfY
2w/ivQuYdr73IOKyILHbn5MOed7tq+lJ8LE96PoJLil0sj4cIctOsT+m5KlugJVxLPd28Yik+cR0
uNRDKIsTRrOsGyBiO5xQg7KcRubxk96jzHAKJCqQUx79IWbc7IzB+P+jnLNWAR8tfQGJVsu9ISZ2
d9NdcQRAaneFpHnF7yx+Svt+/SRlmL7thtIHVY7fVMzUBIzKCBDzP4uupeY7vdgDeJQMVrW7vZgU
NLCPqCuTt3tNhYpR14EvLjPhzhFr1eriB2nG64GhmAwA24dF2D2SSKvmRF47wqVgLQ4cw6RUErw/
JjNBFicnZFjiDMSAc4ewxTUkkmNUkaGiRQtC85URXTBku+mOHITauQZDElg0fyN1qmzILhCzzDJW
DmUoHHLoMVOFRWVWKwyJzlTnxdOVYXxkH3zNylzJ71DSt0JODanlma2Tlrnyrk1mI7i1/O1z81rS
r7anj+Jrv9Q7BN9iBt6nZi3PZr0P+l/AQjLgiFOXd2DYgT8Qq5uWMbKci3z3SORop3oTUVILeJGD
+VA02VcI6neS+yFLkGJQLb0H16SyLKpEhN17qzB6S95GO7qRUR11Ondeio4Ak5JCKRaL9KtBIs2s
6jjNVo64EOFBj2pYLH1H7lvelsVelu5TI9PYGDyTR1IfF+fmKMxXZWp1kWq7P71tOorofnSjssQs
+DsDTM2EHzYHXoilAQSGD6tmyZQ3ddOCVRvNCu/IH+F3NUCDsGh3sZ9s76R7qmUeByRAJzDoRFCu
Rea+fvg2+Bal/0R3/N7eav0xMAeDZm+GTXXHwZP3EHqIBz874+6Jxsbdp/j1xW7e++Yxu3StTiw3
c0zFwtIlG2ZCZgMD7eQRFNxsocq2Q4WaM8ydwj5Y+LPwNDOWF+KrCIEeqPwNNjA8cGfA5132lLow
VccHX6OxgF4S/KDw8YWGosENNvV6v18vqcIAvqVRFO47P4AQXbqcbSHw7DNHs2KsruZbVVucwbTg
GAarRDW1kL5HEkTrINpi+Ej+DlJq9W1HoXs7Q8fsFClEjpaLcR9u5Qh1KYyZzq+h5uTP9AC4mekP
woj7yK+WK6Xvk6V5e9urAlTPXOVtEJsvObOtNYKXcFKB96iNVIVGd0/fTUHaNnKJsGN0EpiuCuK7
Tn3vNuEREmn/i5Yo08QtZWYPEu+Pz+VVD9QdO1ZVRZfeiRSqE/dNhmhDKUukjBs1NWEaVQRSZvjH
j7NlG9QDos9JWilA5Qxnpt546K0sf5xF6aUCGEK+YNemryZ2/NPYOZtldu6d7k5765l3wy2GNeJu
akL7DR4Hhw/PuaNgwC36TemOfQQYJGN3Gq6d65VMGhf3u8iaj9IyYHBg9ZwPJctxE+6oMC956VKf
m+jfmUp7F9zoEGKFVmGF0MQgOQRa0+JIgzNIpPhs+lw982M2J4t7+Dcp3mqxyXqzWZonj4VyD1OO
6ClVUcRajdpSKbVv5rYkYRXjc0/556oNkqCA1YP2uysBgbuvYKADh2oBHaz4kjZztp7JiCW1jmVN
S4zIQV7vYWeRpqLSXJfCD4iK7pETo7FBcy/4LAu3VJ2C6E3bMyYJC4txPb+zoxtyf4N8B8hdLEHk
IKWKfIp1aFAM6k3XCSP5X5aS1ZTt5YDgVKl8KM4dSnZ00aw66Oo/qu9q41xIg9RnBv8bNwWz3Nmu
+mRr1barbLLJM3JxGKH5nh1LMrJ4NMYzgrv0Pb6zRlKz09IpFQWogosKRd3uj1Ea4+BlhPjgEkOS
YF1DoS912EUo3AIJX0gh9QqxvE2yPuF3elZAMhjZrvbQvgBOEzx+eVDtW5bGqGOcCgjps71ldZJy
vs0wEfEj+cSf38P6FNI8a6Iua3TXnY7k0ECpJzJ979vff+MhKDcUfpBpBip9VRnULm2lAiyiKQoR
Mcn6rDYJK8GidDEDrJ2qq7wfxuGkeoG3dS7HFqPNgFfPIU5Ic7ikCVyZu9ED+uum6aeH+KeiIOy2
MjiKfwDFYAom62ELR9oO2yLFO7vJYyP3N1ag4oJjW7bI7A0YN7ryJT4ZTUurzf/kbIdTsMAQ32Jz
ZVwoTZLhqOxaz2GHMfoQjSqyaNLWt5kOC3hfMO5/OD3wrKCWuasFu90if9O8y4rgxTPG009UBmwD
B4dmsFt1PghOw1uoog//2AiVvAvYniKWpdZVBZ1dMyHBWjkLh1g50/9tNFGdQzs4EJVMLePfhG7z
lt5pechTNKrzzMeMp2lokZQRG7zQVGccG/fpuG0mHyZdEmoAktgPFDKR+E4/Wm8s9DuZobUv1BDd
xvA0PJaUWfv8+MatE/6oic3yKK3NbEfXBqvUTdI4ALv4fZiyiBz438OVuYseUygd9GMF1ex5BjrK
tMPhpEkI7RXfJIosMHBGd4DGZURqekl/GU7JZAb6xFK9IuBUr7GpeWbxKetedqRHhuX5sTZPfu/v
rPqp0tGRg2TWI24zm1yUdBYyK8faFP8IXUVG6S8gSIcgHYoOlr6B36wpUYUgvnNIHH648yG3deU9
iBIRkr4+4XzVivBasIawbhVO4csGnwRZZAsoer9j1d1CJ3Ixmi9H7YEkgubTLgLL39xFfIAsPKCU
+dTFP9q+Wue2L2bLWMRO9LyhAFNvNiIydz84sdwin26PjLtLmL0j7FL2TnUiYCkw7Hy2PQ4p86l8
Y8/5yJt/DkYQileoJrTBr9GUGXJ4xXfBUoYOl/lPgJqG+zr7i+/0ZargKMUmn5ZWQrWcYe+HGjx7
v8maWYnleV5bK1CFjoXMUvdGdjIdenl/swmlWY3u7qS1GAKf3hK1m7OSY5fMvhxaObtNnHFr1iDu
Qw6/baCDoRrhKdxt9DZaTzWS4kLDdehnHn1LW2MjMNoXcx4Oc4f6ZpwwaXJTmpVgGKxLkl+xLFTP
e2ca0Aenl9nBCcynSlNI7+nJQyqmpE68aWUJKbgZ4PbEXeQs2dyXcRdZJv3xIr4CMlUOmjESMEP5
Ru1uhVGaHej6PeiTX+jR31Vt7C/qn3Lj96lLxKDofAvRP+pPMvNzevCiX7ZxWTn5wtqktZ7Q6LN8
0oIXlQXnEefY4c/i3mabrY0Idkt97ULfok8h7tIvuE+OR4jVpSrWYertFG+rqRHdJbpKUpbFbPEp
0JiPwNqp8M0/QHpgaDijJn9J35rhgOyQDCVo4gHtWAF2IypoCVZvmnqczCRjQru0AlRQ4L6pxo5H
OUIAS8CzFSkZf9WSQPi995UDanWRbF0GE50sbuz+Fcpzr2+rmw38KVfsui4/jMS+Lu+/daVplC2X
nH8kyEF5V3QoDvASPFMcLpL1z1bKXLCHV3ZobGt1MYIcQpUFeh2f2iXNMuZrrMoDVWolLjP+UZSs
NFeTw8jvckV9+cAECpf7P9XH5wliP/1zOlSHRy0hb9GBKVBpMfVQubvN8k/Ug5m/8WAw5BUOgtuG
vZoTOMGWdSbl3rDp1DPbMGsmaNeQx57vo2UQ5hd7ADclErKvBdUReEVrQTye0p/pYswYFDxMqtjQ
XCD91SnSIhut698vgmfoeLuynw6aEKYmQ7epMTswC1IqgS+Jf/e9rM80dESj/+eyVVxgx5xQ1ZWF
VMJxbhwAvn2IRPm4596Pa5pd5lMFRzpfhXkoEanGLsAcy9pj/wh836d7/3R4g9/l8cSL1JsTnypU
3GrU8rQmDQsxsqzl8LuScDbTE2ftyodvOC0f/a8nD6MkvkSfWei514XOwubDwB23LlAEtTZmmc6g
6oFFFI4cbjlm/xFFPvtzQwIVc3Fh4SZMrtHm7s8hCgtcINXqTxESWd5yIh47buylURqwmUeauY0n
eSNgUJt8fhDAZta9dq6MB5Q2YWq4N+PiCkvR8iPtV3Vd3TufkyP7M6w0hLnVoquQJXxgfxIIeS3h
AOMOxYDffSzVB8n5OXMsUxHoiCQrmwz/BdE8kTpFB4hZF+6BemNQDYhQAHs2GTbEzd5G1WHrpssh
UMbNGup1o9Z+2ME535whlVJHdLEJjtWCG3Tw4JDJ/CWTq4aQqlTBYslFHUChHr5lCSzOXI/qb47B
Tu2NVZ6boe1BAQ6Cx892TZrJtp61W871a7AjCmgk87L9vHzh2cl7pBLXEDXJWj5ObFC+tBGWfaDR
NnNblh3INJuLW6+RnE2zWwKs+ZsimUNcycnQqcOhXoHs+jP93elc71US94cqbPr0X8nFlQ05R8i3
aOReKHpL6X6xSEV+x/OOUelQDWCqLUqY7kPuz3UAyybacTL84aL9FoMM6RrkrDijg41KXbXXh5d/
x+gXq2nrKHjntcfJusUY50y1cHy6FGmCpAyiP4HaGSFiac0YFeFiiWWYgs+XnRelcQYnCOvy324V
Me6cDyawdnZtF+UfMbiCTPgK+ncCrzx23/WFrhBgciQneovZnf3cQ1ZSPj/c5ezIiHY8962RFDHB
l6Gj0nNfcEK/jFlSJMQt62vu1pkIZTK58grTEisbK0wy8dZoAOYPGNcIu2UpWxPbvFyGEri9Xdd0
1ProkK5JREoFBOKrIUFrcAX9LEuGe84sHNf6E1gpr1qsA2VZw0m5O1bJPkCYfUIg3iJvZzeW+vWZ
iMcwuj6YC4/vqzLgnXZOIpEh3Xt+ut9u5ntBV3TC5uhN0DLwBhJ2T4WC2Kquv/35PiHZsb0wUu5G
jKK+E6tsu9ZiAvNI26iCooDZIVGzkwPoyLM7oIDrGxdI3F1Ygav7Zq/pGnFJiCVyhZ0m2S4TCpID
pN0wvQ0em9aRQakw3S8FVIm/R4ocJb3uo3Qul5jYa3SrsfhoXFr5ujNvJAMbTbiYB6DvgIv3vuCJ
var4tDJIuwrljUAsaYGSxNKO5u0NdujwhgyOPa7umR0B51TxaiAMwb1CI8mc8OMSuIbIH2+qYs6J
hwdJlRQuHLwhL4vYLraAbg34nOLt4dFXyJdI9+dsPqrUiC5ln7NQQioMLYNXWZsaxvOvRdk2VAE0
8kQX5VzYY/SzJ/9MFAciuYz+oR64P/WJBv3KIHBTz2EwqcJwLLeWKWx6CVMV/krpr9Zw4t01VoXq
0W9zqn07bAOpR8fky1L29XyDUeIpMCYJ6QnnaB7y9+g1hp7vfHm05NQYy59dRqm98KOCw2Ncx9BO
+BaSwHku5ksgGf21Q4dBqT/v8CHynmbE3kpv7UqASjU54oDjL6aXY2CXS49Gvj5KztZw8znoeiDZ
0sLUDGBBx7oHiNJREcP2iTocEe5HIT2j4qW7MfG19uie6KHCAnF+Tf1zFg7N80RnrrzBQ/N4MDfT
k8FlrwRmvCWBu0XwrngsNYUTDS0ldXvNpoZ3IUhBH3sk2SQR8V9HUcCD+2OEXH6iyi7UZlBWYHsT
TNemQqtmGkbvwW0V/rRjB+ZlRqIR+rVsKs/HzF5y+Y4YOdD5Mr3PSojZkdNPHatKRZbEb1L8EkNG
eePIYsoO8HamfpGmmzhZPXqm7RshSdHatVmi5GRiDZTps/eRiT5oLKLRvTczC5aKn+5tBBTyM0VI
9Ym+YJSrR56K7Au6wMSIMsj9M8aIlGbz57MURS4ehHlqQG9kF7SK29bs5G8E0KmVu1ZMDovek/Wm
2kz8VMAElqy6opb6ZZ/k2kdBOb6MV7hwcUDH1rSqo6JdDDJNVEV6duug4jVfibg33qdGbRkhHkL9
g6Nk2QrqFUAlIcAuZpPeYsR0deZYyWKWp6s7++KUwlZbndLOKpx/rKL64uYndnQxA++fyXmOpjwf
0W4j/piNAs7mP2QC26Zaa1HyeZT20fVoXhsuHgUCg0p/xzGNBp6B03bnHIjaMmmc/p3iBtzQ8jdc
pqMb9He6U4HvbcHWo76+nfzD4m6G/yFLoa+sQyRs0FoxfpSik3xA6ZDCJqJOM08dQ7Gkk2xPWkdb
+a4UQxkZ/Nh5Qt7ujF692rWeex1+j1MoJWahLGevECK0H8rXKyTJKemYsb0zkpCWitGCYKkkLhJO
p8JxZDuybio/WgPPvs/RwRFn/2JGrDcvnqAeFyqdgXwuaQWy+vL1+eAXROebGO7hnX4jN1vVSaxi
0UDTFBxszXHbqc8n89qk9v0XJYzU9W3f7oxm0ihR/EgIhGeCRO6cQibprNURA90r8WFJlxTXWvSt
uYftsEY+EB9eGzV1ti6soZxDtbiX/6wBhXecj1xe8m3vUUiifQdtOyO/9uf/Cepvis1qcMa2R1bB
t3dNqlyyMabt/4No5uz8Vd3oeDCwNJ2NbCEe6DpmyygHXkhrzr/tSYNgh2gDSz1JF0X9WapayH0i
I1EaEEe2iJvmTxoYPXmfLI4UWxv2HL9FnPyIe9lje5fNzCbpFmiZE3E2nXs/I1xpW/GcCC+1j6Lg
rBaJCHW7EK1yEsTYG+EAMg0j78c+2qjSc26xGjPvjDsCWXQ6VzcVMzCSZfaqBDelXKA3gjxk7VfI
eMXMgg/P8kWvmVkgwEx0r27QcnjEQmbEy7qyjboSGZnbqD7sBV0v1T6P+ceT0ahTCHmcR9GsS69R
ebCksrf4OfaoSNuPhbB4Ajb57DfI88Y5HVCQc3wR3vZBBq9Gi27XICvdnlRMcHACzqjjktk5RMQ3
Rz/mmc8lQf44un0t0oTjJ5nk0mjruaL8DHsHFhNo/O+LohIYZ5fDFgicOzFbpWM0oTctB031V0qE
DRuT9w8fa/+GwUnzS5g/G+206aWUXhYNfYPL0UAMRu03aKQeuqMSa5iu4tDrVbM6BTlMantEsFpl
p0MtncSjh4wHYGHtK12eDkg8kD33OjTanHiFELYmpJs6cI3/Qq8YW482Y+ihG7hxYUog75b/HSRB
b18gB/pb61A05v+g1iIz/2BNEazeLSekERmLqqBmYwqplDoa200+JZLaW1/nfpzvAlsz77/9Vnl6
gGFwkX21I+xkrnyH0USSVgoNsrHkk/wpgCMY7uZZCEITi0zrLr4A8wKCswbqs024T+nwGZkxJbFB
ZplFTznS0HRlIGbKpJe1GOlYb4fHUNBvusooB/v0FH4t/nIHdD2lxcW6sD7BtfjTi4nJ7QBUgFV0
0KNF8auMAoh8ihZykXdOdgIBK4Twwtc6tiEcEonp81nwURwf2ex1hOjz5oWs9VMJPa77s0gLBAg9
HnOLL5HBY7TWM8FT9mVI/1e6C8GTAYgYb0wp35EPTvseUfQrVgl5OAaj5obElj738MNNrMM8TIjt
2DvENbnX4jePaVEg3l7o8DHWrepZU8C7VQrIX2dfTTHMKqVoR2Re2DSfJwgcZckQDW9A+F+U16Wh
EDd0xwpht2/VvFVS9kvZ2vI5n6IIpBx/D7ucNh2s0/Ntur0HlRVKYaxgo0vbXF5Gd5DaIdU7Xv8U
IY4v+6kzEf4OwcFbp5X5/e2o1duR3u8LS0eUVfWSA/CxM6dX7WEmyzDd+3bpFe7hLJBSILgrWuRH
E1558d9pfGTxX1qhqaMhICZJs1yo0VsvqpkJgQjQuyn/TWi8If+pCNM8CZKLIaOProWlX8ArWSWf
C+J8GFgeLOhr3RUMjy0d5parh6N/FYGOz+/ooyezPxBizy/rlsofeMIOWoTL7gWMlLIP/kpTXoub
W8Zr6Wq5WK4b4GsqNDe/xzsm9vL7bG74pGA3+VPdwxTeetkvv+4v6egknIbHB0T8f8WH5mKXoQOJ
fAd0yF5Ik9lK5bvT+MYX1ZSeGEOTZuywVy7gPNOIu44FN8J1+mzwTsgEAuoWf92cOgpjn7DHr/LQ
KmZG6DLMsD8jm9tcM1tGPeI0/+w87BT/K9ReSccxn+uWyTyv4RJAEFobSur+H/3+chqkEsEq5Y06
QK6vlj/61yJq7/UvSCGhoEaCBuoip3l0Jsmem7LDRuOtmARawFDI14g/ogmKzy2fGCkqKipuRkTk
GlS34eaiLkBPEORlydl4RgmNJ+eYDgzQoSSUuZRS3+Xp4s4HO1POrte48xKD3yHYeytLYC9OE7zX
Hkn5Vlv60VnoyGqMmqzoNbtTxqrhRzM0MB0s5muq09W2+g1agmYFfCpkF77wZLwleRO4JBGOahBV
kPkOxwvC50kZcLK0xiAmAgvO8x0uI3+UYGTOH5fAAsp4Kj2B7diGScGm+VhrMCplwqR3p6NbN/ZA
r5/Qfd6Mqix46MT9jZVfNBeGKr/yeyVhIarZ/LFdh8v4lDreHY/3LBVp0WdAV572ZnmCZtc/PFkh
82zaQxDQ9Xvs1sooeeMdJq+Ca4EiLJkZk5olDbi9rMqFhYH/OREtYel+G0I2ncGYkbMliPacn9kj
LDDCEce3cVaUyR+VoUuMr0OP5As8Dz94Qh6f2Mexf8HYfh8WA8Ka31z41OoTI89JNFLJKI0OPbi/
mB9ONOrtBZ1GJenhsz5AfEnXVdFMmpTx6SY4Vug80AilFNro0Ernj09LLH35M0TeqJAG5G90fyJ+
xfpZbIuxWyLzNDE3+rVaI4+frmGXECOooukqcTTgVffhhbozcxTy7iVQhR5hBnLxOXSCR4YY31H+
8sFL0li3ny4M3E2WEWKrSyzV33z6drlYh7uV729VARIf3NMqzgnfWbAYGWuoa9ZDo+8B9qWXKeob
Ty0DRhCxmkTiiRUQDP02WBQUS8b5pp4LOZeYQ/a4UqNIFSoF9a0hTZNmtbePvqyPvFrMQ771/oI8
Ko+P2MG/25XTYD9U59DuMou66sVemA39cA8Y5xawAWnfpjt1+v5CR9q0LdROf9L+BJUZSK/BtFfF
+z6kvASuYkfbA+Vi66WnWf9Jsmy8Fu0AyaBt6CLPgg0s8Z0D2e4cbDiA/nQdCkQ3eKfnc5QlC1ZD
V1JEMj06dfxfHThjKD8fUaUXt+VOqmW6+WNXaiOs3IH3aZ+q3UNykWEz9xDp8lajAJeAlk/hh9fN
f9MS0rbveRfyS2NqfMbFLUvpKg8BTSNCMBOrtR2kY8ldHQci8qYGHhwPXDMmmGoSbs6CDK625CjR
aSTqaWUU7EmZI8zAiogdjMJAyOia71zjarDx+MdKIFJ4GfqyAiPOb8d1c0v+Z4NZeTSdEMm7h4/F
pZ0unFFcCTnZW9VBBpyYg5/+wUn9jcVXM+BGBB4wxoJ0VANlX2F5yIEdM8/xaMS783pakka8UeBH
ebUrAifZjrF0dAx8Jhp91OT7Kvuo1FgC1559o3ZB2U2RPnzC/scfkeim7OXU+6ZfS2cDp2HAhqRE
BoyYKeAevHBkL7TYjuaPKAsBxzszZ1Z9Qt5FBb4yLetyrBNBbk+QPDlu4nxJff9z0VJb0s8Silap
4DYTUgbPUOMC//ZAlVZH05k3dgPl8xJFU9YOIpR6TIHf98pKTu6CRc9zALifSQRZH3p9tPT7aMCW
EmykZUwR0F6XsK70/53thKM5cKULMrjzSiqV6PeADNs+OnYEyzjR1Wdx/t6N/It/05nQDIK4SRxM
1zpDyI3hpE07+EqBAGxKLGRjNvxalvsnLsslgb+EGrTlxv2XwvvKd1zUzhKGAs/16JHnq7A/PcFd
esbBXrt802nDtvnSjzdDsnkcJ9WnoUNT2xn4OcB/yyFeZRjnispqqL8o1limL8+EM073bRSYvWGa
tzapMgZwozh0reubajBWu9RCVql5iGDN+A36NegmYXoUYWBbNu5xsk2yp0ZZ/8ERsKUvKLzjXwjM
URqgwzTp9ahVI8GsYH4Zi3/YKWgTm91pfuIvzKN3lNcymYBIXfSiVLUDip7JgsFVfjpBuf8bf0af
Q8ZlWgDIXpNTZN5qNjedLAknRHxyzhRq32aFQ/1WDo9F8pL2PyFSn5i/CQ56+mrojFoWokZDyZFD
eghTJhNo45tFlioz51q1UUAG4043WIIJnzBoUPbCHj67Idbx81QD8S2Ry/qXxfyA5yJqStYDUM77
Wr2iRB1tRF6wyS6kP5E/DQ/CF6abnc9A1uXY7bK2RIWwn/yymlOwzcyymlJTOjX3l3MqKvG3O2SC
fxidMlY1wKOkZUJkNeOHbBMaCCtPgAchBJaO5rBue2k7TuyZcZGLHSBx5Uo+3jLI+ZLBO+wlHw6Q
8l6J+zJW5hjtQJTjoOVZHpXHxgtvs0Eny34Glvkge+2JA8+FKUX62BS7bbU/LrObTm9+u9RmKC/f
Okst3EHFS/jHJgOBAn6Q+mC1Uixexjo931IACYet9KmGfJhpQsGpV1HKWgp56LWCi9k/8TDj1pR4
CSyIY/cSyDWmMusN4k2dRxytzbTXIP2Iow/P8FJ9DFVISZCQa4E+xV3Txp811zgZZBlyXy+LlgPG
reklHXWdSRdeMuwyirfxpCGzXho6909zVEYZ/X+z4SDxWv2acz7IAydakUVmXkXzDEgGK9xXbewQ
KMJwXr62MB2/03/kpSn+HhPqQcGrlEOAta/VV8yA/YsQLhY0V7+vxYurpzCkHLJU59R6JYxoDPfI
qA3OK4miL09vSizPsiAfYTg1VX96bJ5d2xV0GAsT+FnfAflzoHTbPfZDf5YuRCanGTLPl0df3oIK
Y5DZwDb7woN3s/zQZHabcoikX79cH9PWDLKmqpgGMHuGu28ZhSSa/1c3Yz4Oqiq1ZjvzX+l4OxSs
YGgnf8d4/Vd/fWlQE/+3nE8MAy6Utd/FVieYzH1HTSr0julrs2gspWUl3a5mV2ZDefxuc/aY5TYv
UnmW+Qs0MvlKYIRyuW1kAm962y56gpJabORTOEveWOOVpVMTqYLednyrTikYcOnTU8Wxgg2dV6VG
ix4uJ8BJhhSp9n0SIeoarR/ZCPkp1v2N7yvDANs7k/egyUNumTCsiurvThnmZWsAWr6JE3LEGVv/
Hxg4cQTQgOoTvDGcgo76V8jSDVfZrLKKl63o7et06vdKo605x+DU/hUwIEW4eP9qsxbn/fJUv3qe
Wrsiq70U1qCwUIqvWtK1QOnIKQjAwwOYhn+GKDIlnerTZlv7eYie7j5JoOC/y2OgET9SDncrXRb8
BAB+/QUsUyfT1LEIJA8u1uwWe7cVmGk7pt4JE0UPC3reOpFsAnJjz/wb0RxFGTVAiXwrWhKL/KH+
CYQ9gP3pPg2hmZU5TajC3cigQnvlnjmkb1k1TFdP5XQEgRZ2UWauKr9dlZDfGoh0KBuSl47FSbl7
tpT9hWu5tAhKgelPEpU5g50I6EiX7TK/Db0NShgJNwpmmOb/JyYY0cqeisE5R00JEdakesZhslZs
zcPnkUmFRhSjqM/EmRLrTOhHo15eQuYkEU6e+ietEsHYv2+Mozc3W9Vv11uKnx86DPKUJW6V6Ne6
CEVacG03yK/LHlRnL26uMQYTnhNsp+cGOmhu5B/M86lMdMX3HyFuXU5IznFSfb0UcI/7fUWNTpsz
lhm04J86ZOcbhax7Un2Vd14ojhc9PG/7Tws9GuRYLWp40CTHESreML8gG8J1GF3s5X8sGGyIbLvx
rq0zQWIXYCep2W1IWnXpLN1g5wRLOwFNq32TVMCQMo1uBeWKn/AFDFaRVVFo2KokzXMRt/JPFLcQ
3HcuckWwRq34emJV1o2eNtM2uCwPFGoQWD8nDZLpPvWW4/q7kparm+2R/iWQRz7Lerys3OuV93wP
aoUhWQGRQRqqozoHWpkj5PAgtT+AT0mjN8ctAxEO6zWswoBjXYuidw2lRe8JreUX8lZ16ekWT8uj
76r9W5pv7E3t0pBdHBKV8T63FGcFsAcQAMoiXjp+v0dZYUuJQZ2qrfvomNLuivJU6C60fYmEZldR
BNWr6uLYmkgdSNoWos3ZKKIkxMSqJOJKalrgCq7ANnROo1OxEqTEve3QhdTs6slCZIIM1j5yLsx6
5QpioI+HCRWXg+mpLUxf/OEFEiXtg+hawDLlB/VCmo0rs3ePW6u/3jSlFEyqrjvDAI9Y+pztvkDD
ApotqssCTwT7gwfx2lRjD0Pa7Eoy4BvE50QZoBali8HG1PhuKBZmM/YJ2bNV49LEQV5Tof527upx
jSGbxed1JBzgynMK/CvMOUX0BpybufxD18ZurvX/GnLGIOxQbeZnioQacU8oEp8GtLVwEI8bI76A
GLTShQoyWaoH8WLer5SFP0Ef+aJMkfSgYrh1NW3P6DQ/AX6cC+uwl5e+PIAxtkQHZFLSn3FMwmhg
Je+5DYKmTXRLblzvA4FQRKgCRz1HdMDuVXRvakIClUdL3XsulPlBRvhUrQpOE7V3m5D+hBTccg3e
+uVubuyMQSTzZJJlTN9jXYWIZrF27FOuEM6UO+4udK/sjF8GiNk4S53igW0UV3K1tvdItFaeXUgs
FMtcjk2IF244BAL8ZO7YUThig0Tg8znCp3VlEq1kbIzqWzJfPwCLrH/lLbgcbUHL++ERfzgHDBKb
ru55ZavJvGfFmY1I+fA+C0huNZ6x3jXnKq4xjMhIXv2ELrkC6gdV7Q6gcoXhctgpJmXDHtfky7mt
q8+undOPKZw3jW36pnAaQn8diaMPuTrYZRvM/LGsWBNS07IzDk0mLIjo7ajqrhQh2QipnVRAO5Jn
wc5oSr+Uj6SYkoXKFSSacV09EUwX6QynQoBO16Q4i47wJcs60qcJfH3XvbW6IxyLYstfdtYaCXGS
yKkJwzr0fp/RQjUoETFiwCLu2Br8kMAQVfxSEHE4guOybWt0kDvoflWyjnpizGKBwCQ22A2HTxh6
HIB6/4Xx63M+zj14Z/1QGRDXwtmTey2WmNQp/r0DRn20W5WEnOgeghdv9f8hdNGj1pFojImBC334
8sRuyQ4cgaDOun+P9KVQ+8N0rcFE44JXXNFBSaL4P0l15uRFT+VY5D8mObvGrz1CKx4wyNfNBfYH
IcXRmCxAexeAilfofSeF0fgTljRabknJ9O6Zksh9eYAWBHUQIn1lCHD+Fho+2QW9y6ueWuMqt03R
Ez1JZPKFPhI5R8i0LtWCDNZk3PtdmUeP617LB23VWzDuy18r3FQ9kQOCK49xvTIDFnI3sQgwuxG6
zEWxAa4LYRwjc3apWQd7A/CxxiI6InkBx4t1vfGDpKPcUiBF5bCOWWNs0+9erkZ2RDdwqllW/cAu
F4+ZfhYSdWzCCcrsbDWrAZwLUJ1/h1r+E5X1y3u9jr+65F0rMkSD2aYOCAu4N/VZSyszDimliwWm
mOs5fUPXOgS2A18+Qs9UkmM54dw1PTsIOUnxTfqg/XwEr/i/bDys6vBubMmFs5QNEG/JoNF3O8TJ
4NxwqQIwrOTEVvQTi/RdGDS+Lq78O6UTPr/NM96wVf40S2e29rG8IcIR4f+1GHxM6LUjCI+PtiXx
xoqEKplQQrvL1nwUEhzfZ/Bq8uU+SAoIWhDlbQvUQk+COTxCBNwwoHcjcMPKuwiC3cqqvJn4qjgY
M3UHJVS3wUa14bhAeuaLzeG6AP2025fonlFUx1vts7EmofmXS1TvSB7FWP0r34iHOAlRzH+Ql+4e
FOo6Xf+VvWQO+jQm20BJA1UZ1ayzDhib/i5GyyIvowyZV0/MmKdH11LhTtgOaO3SIcbijCqjvQlu
Zs0uFtrsIB7PfxB2cJJI5NSKI5ScRVm2mYJpFyrh8zYNQv1gd8K8xYyYxSnxe0pnP+hY2oiKZhKX
GnCn5FKthKecUNPpT9z4WB9GgulqStOxSjbAvaDrVUxyfqSaND9v+JmYofBoMcSTWEt1qMwWpc0k
Q842nmDUcU6C3WVpJZwi7AzhF5gpbhuN0hsv3lgUDLjPEUB2jM7hJ2DVKkOvdf5tPh5HjEfjHpv+
QBjdsKjcbfpXOGGfyOj6mHkPtAtlCaKTtK1ul39C0Hwa4BT1NDKqBNKKmlE8e3bOzBR2l8qE+IsB
KWZC2PYMH6Kn4yJrWw3cn9Yf3na6v9MC+OMZP4TQulDg6IWNRjXc9W4XOkQSVCPFpJLmyf4AkQVP
LzZj/7PsxeedAo/CLdkPRtb5TO0Ua+vd/f2ekhBRF1ysFIeDRAdLTf7kIWoZunQPyrF0aLSWMx9S
WiIS82jGkKIV0AjZTTUS9Fag2ZrEUeo1FUmpcQ7aSjn2LIFa39N82iaDQhBnKXwF6tsIUwF9Momm
gdKyfEEoSPibei6KCzSRixyfKC7z71DmErDwSfJxgQgzC+XrBIFecnJeM+DknEjz4phmzzJ0LXvv
hanwnsiESqkDICAreL76/t31Lg9ZjoqCgGQtVaygmUUkB3An48etGHEwiF2oyZQ2v3yggUHAbK+S
7itHQUE9fI1xVXLU9QWT2QQLHqXBRXPE26YE4sUOjp/gx8FhTe2xMEiqP2Cpj22gVyKAls7vT3CH
UxkykRv8bjinqxY4e3BvObYk0dSKfWS6HZEGB1dV28AuY8qXze9ezn9S54sSow5F+YbM6oumXymk
EhT1nTRLZ9AM33/TX9huwWH3X8rScj1NGmGl3HjONbh5QzPXi7Zkkr13ZCjRyWGnFPb5UBMeC4p0
xAteB5QUn/ZJNrI/UTponJIa6vf81xgY1Kj1Tpe2HPtDt52ng7WjVi12c7YmC7UYhPwbeTZCwcjE
0Pmb4XVWzeUyQ27dk1gkRma14o8gqkklk4uypYaADYxo/3R4a/EXO2NeF9YXEHRrY5vrwG5+LyWb
UtKWVIrJAep2Blv+6SRzel6S1TC5ZNvxcTj+7pohHQBlbEEPeIhbwhfSotMV1LsTtcvL51W2IQ6D
TNkSB6Cr8Fktdc4POWNigU2hjijcEYGsfIccRmailyf7BX5iQoWZuUpkGD5wzDM3Y+2Ud2Y2bBj6
fC19QffH5IsqawJHyfSp4eZ+5H1vXCIQMrmsiqR08i1aZCGrJdVrbLYrcn/Bd1mFToh130Iqqq4f
Mcu3fElosN9ndY8ivEJTYGy2m/8mzoNO51OMcCKH1issPW+kMT8WQJKyUJLKKKbsTfYNEdSV4tgm
Oz/PovY/yNgjMtfOrMWuqZsAVVbRr3vr2xCQEuVKBmkV3VGyJ9IPO/SFW+acWcAAOYIbAsNkL6X0
un0wOlgstdg0QZKJwj4iXz8kkB0RD6uzz/NczdeYssc+rPtir9Au1roy9De7UwB+QxDcAVE21Efq
tqvvKfmJaV8seaXPMzqmyMIfh64vdab3zswRSUh9xpV7RMqr9LWuGfws9wRNhxOXs6I9iKbsJSgm
j2KRVWwfegRp1oxduHVGzn76jKTyaGlaygjiOsp4K5dO9Z4vtlmu8K+pfCnbxABkYKMbUZoYvICT
vefX8HpyFj0KjHz+6rQ75cvMQShtpg+ZxvtnEkUuGjahpXVRuqCi4d8PpW0QquiC/8krVEA44phA
OqHvUrN8jHESOhpq0kd1jVDymhaZ3QriJNUTHDkKvncPQOxubkocRvrn6b8VKl6Y0qAnCUb51bB3
vG3/BBHx1hX0BAuXpLLFkGOj6vAF/Zfo/JR8hQ/x1s32dXStYg5JxRFHLYy39nXj10L6XjNIRnvb
TWQQzrrbywtPKNEK2cVmU8fU7blA1M8IFNQqaTpisGpwYN066+yjUDKb8KBnLI8rtpDu7OFXtB1x
gBeJI//iDTzMwGQWgs8l16UanscXetxgwVwxr5xAuYnqN6Tib3KZvAbAHN8l1lIvLQvFM6inQ4Rp
/9RXg0evqUIKP+0uJbJ8sc7YMopsVaOoUBmxT9hcq2c0yXbSUHKOT9Z+75k9d7gGUTDKb7lW1RBs
YXbjzGHfWukKEUSFfUXUzbHmtAVosH9JbRrTGkyKxXy/ftE/Nnor1DuwVQkQq1ogEcIToAGd7mqi
0kjRwcOo1wj7Yq25bEIshMll75w6ywzX8wz/WK4vvHxK1oyVMujBQhW95ljJyFBofNijmaMaXNxe
XMS3lfzWgkFiy5FSdiFM1dIc7eAr+Pnor7gX4SBKVbc9i7rUKnS1zwtxznUgo2cAEZkDZq01/sCk
U3JGVbojSL4uFvwcJ5MRj09AFyQNcMqZ+elkSEoFPrU4Ayo9HJoc/VrG7JtZgC4vsJJJnOUd1HAT
PE4+cmTPp8HpoQDz+KHya67JjzJlquH55l4W8FH4TzUDW8P+RC7OViUa17ANAJLNUP0dn1TgupvH
BF7j2fhhXuhvNcq16ZwRq1SNd0Td1Qx1PQ/Kh8B6NMqiAEY76RA4+7KGwKwDsVaZd8CxqbHiBaim
Joez4b7icfRtRu/eH1vF+ZkEY0os2peLZ66tliKYAkvTKnmk71HghKrK/jzk7ENQ8Acjx4NIGsax
QuVfaRUbrwbK04kiB1VdtO44X5yoaGxBm/ihTDvhVadKe9mlA+5loZ/jr6O5o8utIy5EBqWKuJyU
HO4MBrPZbFtt5nX1P+LahurnJO55vfh1CBb30IgjpKg+TpkzHbCFamogJN6Q/cTBPvTGgGJlWVwp
t/iZOL9Nm8hX2NjvewR5ozQ+4wDD2rkaWERIOktfVRhzTy4MMvgWMujoyewZLIqAafdNuiAU7Sxq
uJF/+e4zzfmS1IvSsNTHIkz8CHKjFwWa0xN1UjNeZi118BDv0x15eV7v5vNwK5vBmKg3S7vFfBr5
3mPO4zXjzAh20/VaXSxgj8RHTFzw0gDyU479Ewpq9YSRGhglS2xZbAcoaVWr+D287r106ibH+Emo
AX+S/EI8QfZUN1/sFSKAgy34dQic4qrNsFOOVjpnPyDQkTUj4uVFN1vkmo/5q+wyf8PjPkB5ITcu
WeoPFZjuf3dWdYnsI24VbWjzOdPXYOkQcCvkuPCLhDDbgA1c8iPyHdpF9wAb5/7gz+9joVHYnQqh
WE6KPOcgcDLwZiKUQfjjUQv7DgIiAkglLLo5w51b+r9vuvVtNJamT6yB0mPKzw0hxOsGJK1x12tO
G4nNUUGF23cbLf+gZc+KEeA4Q9rgDw1pq+SsY3aN8cCP+h3/i9dbtyGFJERlwCNBYnEeI/UbFxa8
ie+ZeUnjf+2qVVKRBSm/9WCutjrdBTb/NRlB8TXhfea/bv4OGyJmUQX55SW43EC9RAN1WcjT+BeJ
VQHjJgrBsaXDX8DExnyOPuaMa8jd6BsXXioscQPjcHZz7ggTEwDrdK/dSIIsj9rYegXIYrREtHgf
n/gcXhagNN8Z59x4m3sMCQ5XY8KCcxFay69NpQHA+f3wmgcMyAjGS1D/8hHAJwCL0Gt0TpaVrGeh
7BibOU9y/kactHH2ZOlFbFO8dFioJkeU3EPqxAjojOo6XsyxIe01wv9MKSYDfqL7CXNALRazj99R
sBVymAs1tHT1PLwM24omWPkszOwETi6JhcbdkTmM4RQ8Itg9YMfaX4AmK+iRa26/EkoftNWVy2qY
fhd5VOkDO77v4N3kfVSzwPZ0BH8VjJajzkznQxjGLkRS7ZkyItcdF1pbryg5xgWaP98Ns2dnLw2T
hRJrgYYGTb3StAhkFMMfMgbgbGZ+4hT/PO2xc+wacnB6zh34wiYDdHn4ropDrzPE+FsG/eajIPIU
Lh7hYYd+GjOYuPurmpQQvGCZR2Kafbn3QiF+LYCJM69vmOs9sUw0NtmuyZZnZNkM2b52RM872p4B
P+/DEfs9BXYTD0DVIhSTBGpQ1tAFyU3AugMercGE7HJIkTRpJJQ+m+vZlRAKybsX2U3zkzthbiiu
VVtv+mC+KkTvrTVvaeSmYRYE0/fxZfKPGqzGynAQu5WI5BTlWWAZk6x+8KMPKgKsvSl93m5aHK31
qlj0gRzk/I7ZsUnq5IbeoSJiaI8+BClNws4dff7PnlyTwl4QLJcgzrk//jNUK1I+yVBGhWAAVLR9
xM/MVuWldFbBFAcIsprdUqEO4ps0Bw0QlDydLLuGIu27XIKvrEyamXE7JPKmAgC5kgdY0lrfgmo7
0j1KC9DHy8QKY3ZsdTiqi8G9bWCi46bm/4aaNV7sVhIFMWI0vy3OQzhEzuE0giNTgz+oa1HWYqoV
oQddZHEyWyX27xgQdOaFQTQ0jheJ87k1Hjupc9Qli8mV5yi2M6tJ7WT38Gx5N1+4V/s0BHVbnNPi
vFOSVNhKGCtoIprGgswpRMqEyT+zNnPckACcMzTuOKnjGDCyCGkD4UlaElroixEuKVnXC4+JTQts
YUNpbWH1Ob8v9uQCxlI56f8vyzL18ogHQGUG0RnDbR/YWcX+orlKhBvXx9uFa2pXQ2EgxI2uKaC2
AYVgPuEh/IjxUNcPGXO2RpUxjf6c6Y46uEqNOnniGhdG5kluvq38ySwJujpwSuGiOyb/oBB+Yjyq
yFOm5ffEl642BObtGD8qtyoa803T+89Si3m6ls640+mg2qC3qKAIYaH+y0caC6RgkXuZeer5n+0L
lpCBOoLNU/SYcN/i/RWFRRIqgRCl5z2pMZBEmSgXaX8Q/iJ+P5CItCSyncO1azMyXUb0lwDn68PE
F6hctLpiesIJEgkBfvQydjIWyHmlFZHmDTcOJADArtdDMjm4jGim32vduOsErUWFaScVgZaaQ6ZS
FyiTr8YEuGzb1ANSNA4YOHj1bSIg6Ac/hJY/Htwvh7A4v6Vng00x+C57m1F2AmGtDRgR6RetEp9+
xIvtV2VXQSi0C8hlpA7TEA44Nndrw/PC2MDxcxaQAdZTh/ketv6XbHpv4wu9NMd55DMxyQt19DO5
WQLHAk25Ix3fa3hCADLsRNVwOyqpZrOtQZWhJZ5ufCXJDeIBN8h3e1V4252xBfjSHRa7sSlVbAZl
TQiNFku5C5O3NFXsOB6BhZq8xOq126Fu89uBYwDmOGAY3jdjFy9rK2B+PfdUnKeMQTLf6eb7mGHg
jv21Ao14iERMgTJifMrjs45EmhyLCItSBhxNKJlhhG8rKxac0HgWILPi8U33xpt1fjvmnoESPWAj
o9ijYDp3tv6ZG5lazW7umjlCA3zqgjdwfXnZIERnj/y9AfQrOyqot/FNfP7UoliKqBZYpv4VSjH0
muYczHbU1uP4Q5z06PxOVCezvhSfK74cnlJZoMxrsBCP5eSrHp8TBh1w4P3UpcVbMs55J62btIix
5cmA64h4sD4GO3VV27CCrfpejysJs9YSdI15Dz6V8ggBe+gaC5rLUf8ZW6nvRXusXWJGEO+dbcNw
dsmh5oxaZqSOm1kJ8ohKEAU3KflzjYfbcs9LQK8guT98DOgaZEu+5MUgti5N4TMLNHWB4QANPuwJ
Iz+g8usc58LQ/JPbVjPPi22PEjWRoPXY+dENWV+PpwGeA3tATrSLYjQwnle1BAP3y8+YlehACDP1
9EIvAfE5tW3v9DE9ohKmucOpDEY3sRY7F/mt1dL4RPLWM+bMEvx1DWES9L6yKcnFmJU7KovMyYiD
5oYg7Z/5YuvIT1WeosQ7Wh3VQjm0X99bTP+qAEOOAsnA5Xd2J251G6vIgNu6XFGYRGte6TZl1X3n
uhZHRLKhpz98xq4UVXNZOzbRzrOhXGcCBAzvGKLIFhiYTBq9F2Oz3IbnuNlJ5vzIN87tEuI1Lena
Y9cyiCWKTunGbDF7bMq0hYmh3i4U0w2bMB0qJ765PmHcHaupYDlbzJoE+uMhIrffLYRiD8vP/8DV
m58sDlrFk/pp2oE13NJzFUxAB8fZPsoOtyxLCUrwrolJ3UUgNRc+/vyakXwhgisVl/Tw3gA9slDH
yC78JWeia4MYDJLizcPytdWHNQXKVpy1pVSSFEHoiAckBSLVAT8XJzvj/GKWgmUcg1bY3Gzvwtxu
ab4Li/R+Fpju9NZRAIQ2bEfB1NqhIk6bdbNQYXMG+Annt/a8/ONXVauC0f1mEaSrzYd6dE77fP1f
A/ehS29CEe/0z68RR+66xkHZ0+zXIf93qui8Z2Y0Zv1fxP3YELWcDr0O9QNYLeJqI8jj3Qip9AP/
JJY9NjCSwFl1hA71SQ0rPKgJTbQB5C8QWwrYfG8SyM9CpAhXwWhnLPEuIbQQNAAiM2dnqw4hq1HA
F69tq92EuMF+WcN5XWNznhJfwua5VLKvnZP21DJpJTk6PrEdpTtBpTVDKJymGXt8YyD71OVVgiWN
hggY/KCFKdmftF1P8bYjNiGvDsppZTynTjoScVjKjnjt5XekUeg7fTL+X1NBEsTQD/JyXBbvVCGj
I1LJzwyHqk2tSzp3ZbUUOIeNdveLv+YIkYfVWtBJ6Ihf42ok8IB2POWkOqk3I2lCuceOeZ8WYNug
XRxe5IlmcUySatuX6yywU9QVtwLgzm0j73svJ6j6+9sbi6yTditbpEjryP9WLluyksxzMitb20ty
zKYXXps/zAw8JJZKE6s8iELx8+LdEzdhoXnrFl9qeG65JUolRXLlRJacaFF5fa3Q7+a9+IT758EN
w2MzZix4Cac7h6oiOmNHXcbJL9wsOlNsSrQh7HIR3xEM7lyjHGS8BSkcq1OVdu2Kaa5o0jksMSNK
WrH6hRT5yINf/YuOJssSUUxjXb6uJyzpA8PigqpHylE9fVT5bGayonaXx3s3Mk3K8sxh6a+6yjyN
QLNDnWjQ0at/N+ClGwBPi+SG3ffHOGH5xCpwHU7nTCJ5MutMZkCe3OR/N9Ljka7i0HAt7GVNnl4q
4I29mkBqAoF5RBsdJIDNBuOj2Q2U65BAf18B6E2zQKk5qV+hulQ0ib2k+OnEL+tkNZMUTjXiPf97
by1ICSN+gBxRGqXj3gnnFHKEwKVcTeZhjaU5WkS9Dk273q7ue6LTNeoXKKFjR4Ct2zUxD6/47xks
P+S/ytlz3hPwI5h4Fqib8NZHJSSjeFO+PRaYGJTxTFrqoYwnVr+gC9Sww/MmP+//Zbj6BN/WohoT
uUtMG3kubVomxH8+YJEzclp+LAsxf8Tll2RylsM1p1QwowDIznBpo48riol4Tm5h1De7rFZ6wP6r
sKl+xljwdU7IACEn8OUmcqHNfB3KmyNxuyP1vwVTc/f21A7WtO2hg44bSOpOREw51hpDmuZAFlMX
R+L3JnRoYqW+Ss0effw8OpVDsNQ16dutwYqQ09AyKT09EE2ChmGZkL2iJBFUWh/55Ldr43F6zDBW
55d3oJEOFF4SEUou6qYQ8fLWInekn6ywIsB4BlO011I11pmQcXTuEjlp8rmc/uHXEnOWjWWvM3rR
WwyaNM2U6A0x2H0iK3hphlx12xcu0BGVN7f0h1B5N/P13oKCZyv46sSsJkt9ZuzaCrlGunPWyQ0E
64Kb9BK7LDOtR68vL3S44bilypAyK690YCj+iY41yfTcMcx06HgVZFy+UIt/FAZHw3Hnk/CHak1S
X5Bhl6xWGOmBXNC1+yHf/21xFK5Jh6xhKe7Am1TnaA5G8kVoTg8tqSvH+hmiZcSMpZeLAxyF7ZgJ
AyxNvheBaGpsfS9gYU5A21weNHRqo2o1zdyotru1hZKsG45+8i62a/r+ZLd8p1QEPG/ab8mkHvwP
cQTwJU/Pf7gghMWkBvVBp53rDbQNsK9I7jR+ESNWzBBzns+DGO7rzcoRWlxtcfrMhNTX7kxJPE02
N3ReHVeFFr+vUN85+FLJNcbLEgGcoiXwaYx8WuYlFherNrVnVQ0mUO168fpfunh5m3jtawYo4Esy
TknDnLgFN6RnlQ+V8BpdvzpNtlQkt1i4pyPpqgDgF6WRrar+Us7VfY3UpuRb+buCPLqfy51atRQK
Fu53dldv8ijqN5oUKuZ+NbEFuKDmI0+Ys0jGEMOPLluyaZJJ/pzVMDAXdaCsrjlD5eWgr74/r5Yd
sDpJMqMvM/b2KBVUTtzeltXUG1kMzq8zpodqsFKlLSXcg3rojV/w9gYc1nIzseE7YfOVj5F9EYtD
AtrLpoymlp4NV0coqxDPODdNj5zySmN0pymstqnn5pbZzbhQ25rXtpB9YDILKb7YuuFX5ySTb80I
aV9NMgkGovXBlYUBBfDZ486xNBnCy06SBGX1OKnC2PqEG2hOufL99ttjFo7edU0iqoatHZ9PNteD
3Mt5CfJnn3N4X/supPnh5xNACpPeC11wcIKZGnQYL91NRsXdtyP8YL55QOUdYFIIbop53TyLLnsN
ryA4J/KsJrSRfYLW4MTWUM4fbtWwISVHLljfL9khrIkMsNONK3m1qgP61VuFGJ76Fmkbshq0ECcg
u5GCN5TTzZENAD+hyJJFLqhV74QYMzLtg7PfgE94bzhPZVz1JGluPubDfih/MPboHnrSOh4g4dGB
liOTBlyuth27lq1K2LNKjafazR0EPaoAzoMpMWXouQbmVQKPFp9lGUfUM/CBxu8q6r+VEoWlRCAM
alg96dl5JOQe7QHUHUNToVBtghao+dRcrMYc1HAqZYAi2W82Uk0HbKTf37uqU4OiHOzSnsSck4vq
RyOBSycmejs8YRwQRQB5f8Xk0W/9keaJU8bLslgazW4x+qTMhx4okh6xMKezCUNpws058TEtGwMx
3AKCQ2v3rN0eQ9tNqn6aOsMt9JRu0SDsx2rYdHVdWhFx31ZTMN2ejQtZEnar6uHj5yhBDW8r4Rf+
6ntdIMfnYYRPyrWP3wIDJWoX4KIIMI0EgokH/h1vbPTxJfDxRJ+2Zkn9OSrzZ3kVy0xVPSEjyGhJ
2/9/I2zZSY+05WU7gq8j3jeZNp4LGTKYQU4GmMmeL2rOZspcw5+CedjU3dq9qjO2WR+4N5QPH617
ll5XP4jaD2rWVHb+rQfOJPGry2azRKiYNMSyDrmQKFTmh0RnXaHByoP7M1Ohvih5eVGqX8EF6EpN
duRai3rEkPBqKiUYlGpENnF5SiynMec+EPaPqAWW7SzgV3Dh6g+fvzPztbWcJ3qOZBSJZ051QmIg
unxZAL7UkJCiD5c5yYwxxJj//BfIN6XibEMrl8vHMtgLlcwxfTZZUahq1s3D7p+mZ5bHpgtQVVmA
P8ItDmF/LSKkR8AER6OwFjUm16iWTQi2RhZTuROtJLg2Ut6DgUbn6N0TWC5S9RV+Ni3IBfKiJLWB
Jui0nZfbQW1d5PQK8Vsj01yJFGX9mGus4cVzw6xRVfsSWgndVHYTXoqmqGJZzohV09ewx1F66SJb
hMRRWJp05J+0yXdyUfU5wzRlYVGQba1KZC2L/WAroYxQRL7RNrfM29vOSpdtYYIwusYZ1fv545Dd
xVSsAJS56LWk9FVUqWa+FE3Dp1iu0wjhbKi/Dp8X+a3QxT2A11dEmmaBZ7TJ2Ribpcdx+2ec9L+9
9v9E8SorS00ldUBQq5Gn8X/zWvoXy2vUB44KfBkDcQKshK5a5ve4dY2Sayw2j4QU8+IANvCNXCwd
u+K1qL4iXb4PED7pi7tfyDgGi3WYxXHAtQLnF8YA2QtsKssJXXHPxqOgknR6o21QSgmrSUDSFCZM
/KcXLGm5ESiVG0y7OTfaCY/1mvZV2mCj2FcYGJtpOifL7LcnuvL9NRqr2MPCBVAPEuISCxOoQ4ZO
WJi+dAYvUmfZRAQGZgWPpJFERnkvkNc1ZdYkkeQ440KeRsRy6335JSbs1SnGgUdM5eSr/Vix2kA2
mPioMBBtIkg0ICCRwYyq4OLdGAE1HTN2BzsLi3rt0agjz5rg4gsh0+rXUsjXMyF1n1Cgz+sDUYUF
4mLYgFlbY1uHil+ps3jDITXPvrSdLXAesTruSuJ9rtd0Vz0N9ydGL17RCyTMLerC1tGmRQWG3iP8
x5DdGaorznZ6bLWxj+wT5hhENFb+DE/0AMFyAdZA5OQW2cCWWG9eWL5sgO2yEnHQWQq+PYLwcqem
SP8sWPutFxHIQy5ZuBQlS/YOXsKKFjrKsZyNJoaOXEv2IJJWCItM4VW7XibNxn7G5If3jMv2icGX
YEH07/kR1UYpxB7s1e8MJMz5X1JhzqIps9NFp3OPgeUTdxF1ed3QA2qNQSo2JWbMuGIWl5OIk4Pd
cGqdLkpQY8Aej9Ookt/3JNZLHQlHdwN32Ar4LSCsVIfikgaz1TAFZlXJG7w+jMLC2Xwy238k03Sx
Ycqoyp6+N2x3hy9TXGpzJtVsy5XLLQ4RtvcuqA6KFinx7NuaPY/4OCfLVUXv3HiCRL1Sv+dCecus
FqoV5t2YvlK+WpG27Of5VCApWV2AYGb0a5Iaj68nFdJy9Ca1qCmi7M1lBAhKwuOSbCJNnSb5/V5B
hvGLUkgCgEDJA5UYQSFnBU92s4L+/1Jh6s7jC7Csgpu1crbtcbFeBLL6ywF9z3nsgT+sL/QDbyDM
mjHYQZzlUWjMziu0Zy6YUyTDsawqHqePD9bik4mKDLI6AiG8fzpqrD42w9BoeU5jS5GiZJRIjRGi
zK5xqr67Smr/hUDp+2+0LnkPmTa6YxtDN75ioQmnKZ1BVPcGwfH+QFAS6TbUse8qRJ6CrU130U0a
+K79PxApANlXMYw2HCaYO7R/NqaVcWNAPskB1wyxMn1MyFTVHrCJ0eaX/In2ct5C6v6sa9B51iiH
dbjDBWwmWATBOmTkc7ALdRvs4D2QnpbzBt5tjkAsHNVzvEIrMHzNVbOH1/5hbw0IZJynjgDKI5Be
YnudDnBtszJOSIg87WZbf166TVASrNY3q6dPL4hS6O9IYa00Mtv7JPM8n7oXYDub9ho0cqDSr7BR
ymvJbTM39h4VDLyKwloTciZBsFHeo1hBoKXTGHt/NyRS27DY5YOIdUlILdlZouCIZ/TjpeEc2/nz
nxlAT08q/UkNIixW8z1EuWw7UbD/LNtRkFUGZGDrsEUu6H7C9/KlseLUG0lCseDr61usbtYGzRJ4
2W+bAkGV3kyEfolcCwPHJqyTj7dBJRHYfiq5/Uaf2yWKl7EZfzhV1jyaqvrAILDUwcLJ5M8YnahZ
uaMrJE0iUff63g7ixvRGgcc1EFLfTXHJ+9JpVxG01W43OoTe9jtgebIqJ+OIefUeBfqyvY+atkcW
euda6s1mhF4TwOsBLSeAkp8UtqnlqkdeN9MkPB5xgYV1Ww6JWXl7QK+0YxvaprHeQ+TYoW7RIUpO
mhjaJQUXUJFS6SwC783BI9The+ovH/fzg38DVtmC8GD1gO67+h5VlnnCK/8ZYfSV1Hqn8lVf+Ikv
loNkLMQxUaDFVglk8ZrIByZSoiskkjvC09SqfEtMHO5XN+At093jq9stv353USAZvIY6pO5Ujsz9
352VyGMCVmU20B/78LFXH2pSOIFswckS8UzY4Fii510HGChUaiJi9Y/r9PFVLiR9aSzPDN1u1zNx
Z29wER6e+IexHEcf0+MxbAm3k5aOkrbloUS/5ZV5h9PtcqWc2x59qaijMep/eUg/eVGVsSPL53RY
pMU0FDnnOW4sSKLF1POY6wxngHn/53dZWgoP+KSwVJ6EXQrx6mKUcqcBX599lKJnBxqaXUkLiQ1F
RiXK9t+ILQK2A6MwmZnrvDg7cVuE11SbjTAxRcIWVeRA/iKvQe8TtBmSxUneaehLrx/hV6ZbPNyn
FFHNSy3IZmU8AkcEp4Egqp1hOsjy+D7L12SPrkHJoxrGLcjIAUigrqRsdCVF0ln8fxQQC5vsMiBn
oRxwdhjDhoasQaj4inR9pFkw8PM3NEIRML7p0mIkfsezdSk+gqiW7JLH1O1JCljzJK/vYwvPs5L5
KeirMY4sLPGQeBwzf54Myhf7OJ6RI19KBdB0MWLsCi30H/cvjOjEAObr2dvli0D49LHZzXg251O4
9IKYTw4jpEu0tDo1xnvc47G25PAY7F80muX3G6CPN+geabtKDpJFjXzRXav3h7uK+TWZfSM3a1Yz
f1dmDUx+Tr9tLw4lGmC441EhDNF595F49Vgs0m80SqHjvJqxHZHhpm4ASNL26/0VlxdsP2S8EXSL
QSWKuKFLcqCVToQbyWlqBjLUSDKIyK7R56EnRSG1sfb7/NPmqWktTm4h6NhMQDnrxwZ5jKlCwhWn
AesKfBVze89iBOuBXHSRe6CERSMaj8603PB341VyRMzDi2PHeZCzBVpS5v1Tt5O6tq254mz9UVWi
5nFWq6JXgYJpWD7KNW53wfLeybEQEAG26D0wXewAuHYbBUGjE6ZlJZRIaTesya2YLF41ZUNvqj+9
QJqM4Ic3GCxz7znWWhaoIu+ro/PGjCTg2vfsV1VcGKnaXEZfE7/3frXxmlNCXadsAbpGOpZhpe9z
mxDAgm0kdA4gDlAO7B4OBQCtgONiI37lRZXtL4zGF/8xpMyEMKyG7iZ0Ml6VGKFG/HRHuQt9OAF8
9Hr0n5dJYZo+1Ye5iWdvxzqEzufkQBJVP80USvqE7/aQtq1g0SgL9VlJPQiRuD8wRSbju6LRi6dZ
uPzESL6s0U2mE3EswGkKmkU83DfEH8XjDycPObbWgNhjLyTY3FMBlzHf3EblD81KzSagf+KNpbin
IjWRFAxN2phImt2jnJbTMnsmJAIOFuZ8xfLKnL4QMIqxc+rVnlCxBJalpD6+i4GRMgR48mXc/OXt
6QS82sYoU/jz9AJxLA7oF+QvCa7sHCvAsUX9teBfkMavV7gfz5CyBOcKFra4UHuFn8nQDdApqgOU
OnzjX3DNw/qjD7CitHs0aUAIFP3WB9e+pv6IUenF7NKKco1g7q0MS9LcCoyH/7sfbynjtzfsa2F3
NebcYpENhxekmtwFRQJ5u8MCAEn4uVUQUWJSKCxqkEyr7xkTuF4vvznWZ7m3zlFNp1piD03+WihO
Lrxy4xk1hVtpHaorLf3EDWPu9jjCvBNwYLjIUhGyvfGl0OXqJYfyxYU3NLADmiEv2a60iygvvjAK
JAzxRzc4yy4N0nLTvVIw/ERsS8XKbjRzZ0q4wMDevji9hrrth5jkKwsDu369uZ8oSDWlZY673+CK
aiV2eek+wzjSsB09kQJR8TWRX+zHHQsDscgCDCRW9BlKZSwm4iOMFOnZBvStK+ucaLEVEGD94Ox4
/KhjyEt0/jEkctXedq4rNHQZHip9Q1k8TuQLg5Qb0AdPWOGrppGSUHYExNyLOdzwbLt4PtbiF0U+
XLtQrwsTEmDBUKap4wg/BRAiDBOvT5DrrMMRpTbqv84+ScRHJroMO7gNt3eX0BuiO50TxY4RZCx+
NJI9+lkYgt2Jvd8uLCtg6+b8L0lEaYbCVHSjko3IYcYhpdxnFa2RAD0ad4WUAgDI0dWJxgGSb5xI
giNT43GmFawBSEWU1iRNfzEmLiBWOEPxn3/4fOMBHrFkfAxBtaDFUvy2Qe8mnlQugVRtiDTbtzWq
/qCwxll6nqU/P5CLIMtPgTEwGyfQ19r2Tmg+CFsLU3CfUD5qhhhEYYsaVxr09vYxTnblaxNo9ccp
NFumggbQjf7QYHM9/2JhLf91Xl+IvbmeXGpWyD/SpMpuJGFrbIKNJ0FRqdoyHsfMKW2iXkMWm2cv
eLQPtHIWCMdlnaIg0iZVwnhKuUYfeKqgUgIF2dIajRgl6fFibVm49IDP2BHCdJj7Nd22ohgMvBAX
acby+QyLHsIPQNFtmI+KOZmUGDTDELzllm0OEPoPsK3He/waoEwRyreuJT+t4Km/Sbrcz/I17V36
67f2rpR/ZfzNQ0hvM817mj2T+Wfc8XmVFwWNs6UXlrhiHqh/Kg4dG9gPEWqvqOuKOgyJ1Jr3Uu5Y
FakgSER/eVXDJMzYrXa/2nh0j8Eo0dM/ObE698kYVopma4ie+EYaxNZplr9LDj1XRIl07BDn6YGg
Rl19YPKVS2w7PAfnMAWU/YajXryoUVkIl6gL16fkC+fh2xq/aUPqQY/IgOuGPqLKwstNCTN5Y8yz
XcTyjfBA+TYWYLuo10btFuQ69PX/PErcRl1hL0er0FtjwgCM+PtksNbrJ6zhaYzIT6psHBlyDGwU
4gqBQnGvz78w4X1IJk4jqDJGcqBn0x4SWTs2Sptz/hHRcnw6rMGXt8J/KuRQye2fVuT7JVXx7ifp
KP6kAkhDUQTkzhrJQiZ95w24llfPTE3uV+8PIrPyqE6s5+FpUdHo+emiVOL5bqcw8wtMmrgdUCda
l7WAgGfVzlVD0Wkt3Dt+mg77bpclZRERpga0lZ6RmaaFLmZeayr9AkF34nDhAakx9m7gOcu05KVc
4dQRQRWLhpmjn+Kg7ZuSWE+FQar8acJ+6cHldZCoRG9sXOAA8eGLxs53ZGAEo9p4PqrzD3bXhcvd
MGT6FXigsEpPoDL1m703ypD/wZUfsElQpaDmgtUN/2//+Vkt/HYtyWXFQXlOKJPKbWsATh3zajeQ
9Y8xoJoZhMbgP1TAmir3XMQrb64oUP9wwM/ikisQhol7px44w4UpLiPr8U8JMDpGt3/gxw49ZLx7
Gwbcpssoq1oIN1qUHqrFVhTiH8Y37JBziFZfnngWMsiIDWBrCKVh1UTcgJXPoGe3+EDAfb9JtoTF
zBFd5PPTeb/PWXEd4Pij8sEGtGWdpB5pFqdUksuOEd9oo0SNXVnXzGbue5wY2g/W9CII2UPq47Fl
JmLHyaNB/tgj0SLD0DZsGTs5qXp35IZBTUOSg83u4anALQ0/XHEgU0YDRFIAdOkX2yksDcKacP8v
7kEAoYymYQchiHggqBlY6kPbG4529F6sWF9/76A5hljO6RqHfOyAwLnXP1Rh2w5gOtnukcCk0qyi
vZt1fwqBH3Br7jLJ4dbwGQIxZoTfXadY6fFHjPMMmYJp6Lc/kiNo7vwhfnkGmqDIRsiSBs/bNOqk
K7UBWjrQ35iLv9E1aVZtJfGuUEs4c/gecShNLFduYeyGD2Dlo5H9SBOOvlS9OK19G9weeMKh87xd
UXZwFaJ0TfSIcYBBGilKMyo+UFHyO1vCsZ5Lxwi/sWwEEB2FbvTUmb6Y43+NiEd6bTGOlcYpW8LR
kgJnbyqyD7TGLTBePVVd5urqfXEqRmBmrM1MFIfIGpUzG6oWGtQNflUPSLMj7LsGqK5ljrrfaO8b
pxEp3+kVqRzx5MPeY1bxmxAU7H68KJU1W0pt5pr6WK4XtKbpiiRH7ufy2WGEOfhaIwak2/EPZH6c
D9q4TEc4YTT19IK/S6X91+3o7ywakFwHumSo/3qUQBap6XSp7Rw3z7pkgFwwPRtRRl8YpvPB1ESr
AxBviYep6hUIRHbOL2WVLfh77lZsCR2S6owQ4GN0Ia8QmGoIqkUiILo9PpDE/hDuhJQr3tg/Qrms
1X/UdJj8rwjlIHvVxej8wv5eyzMf8MYDKcuyvWkhxrHB4WXd8erXjoMBkLVmdbAFLoYKb80wQG+j
av+oGLnnvfY/sMu+jaWSFLdpErBZQQGyxVNdz60DVya+bA9wlmOY+0bkV6E1IKbWV13K477c1EEg
NHgV1kObS4C2Co1g03UIJ/0d69hWFXZlDFa3VG8H4SMCAuLVWyXC1Cp6F87ZM0uqBmNszOGg9QJL
4EObOLSxcQZwLdA3kG4V5ouNGdIkRzUYwd3LI3HNKVxjQzxWQIPg7VsrIZ7nYCzM87VGjH4DiZsn
769sDU2hHDkkEydTiiH5P/WjSSy75/VTua8n94/izoYP2xU+R9Qikjg3nNYSzblH6tGQTfEDxWjC
yJVeJiUDGWGfiMVlMMh6rr4ViPoGD6CkzH5+fr7UEOo2mNbwtAmbjV/iTYL5jpYyUnMHt+STEBmY
4uu1YyA4fDBA04tP1yrFZ0UWDgnWUu0cHsMzXXKomrU07zbzj6dfhlIkMI/K+YFTjmuitVgwVuuQ
VKr9xVlcq/yiCTj1G2g74Zi58u2LTSNNOczs1b7S8xJYMJ/GIwD2mIqLf7R5X8d/s1XD9YWCtTRB
e2sA7B0Rs0v84KfOoKP+J9FAnhAuma99eB3iJWoQhTifIiH7P7CHP6jO+dj5ZznCZ2WFlG/eKtFN
5/MJDzU7V1hopShVocuC9s2ZpUUH+KOYhi8Fa3I8Jg2n785QaaYuw3xIR9gPV/dTMD77J7ddx3O4
6id3/vX+bQabk32LN3yHTgvTp9rSYMFzM8eneOYKo1mvFtmLdd15lTLhvl8EFIoXjdD6GDH7rGoC
+BZCx3iaUnrpWJjVox9Rugbv4IhFvgMBjPw5QCIfpp4R2RsJNHgYH6O527p8SwkPD8zEBg5cNEpu
JVdsYPfuj3fuSquWviuOyHIXE4Qn/RcvABIx7qQ8kkeQVWqoisfnakYykVq4aDiTfHw/GAEO47jN
Ze9l4D3SamxII4FIkcT/RAeC+7MX1DCybvkYUjHLySTrKcgngwHJ8YXJ20lr+lfeYu76A+5TS8SE
FJuh2LhC7pbr+WOEsZvVc8R6WRQ/bj0urNJ1RPyWTuVJYrPdbmvG1sSSFUHB0WZz263yDhfKIyBQ
ZOygv2uSsvGT2/VSC3qICkUN+hJMYwdIRCoFH+mTB++iPPWl//Y4pGFwPGJ1oQBRKGuHI+u9iZKF
ARybE8DyMRDwTlyzObDL/zxSj8y9QGvhMp20pJmaQUS4IBWJQM8wywB++ssEZPvtxGwQu+exMupd
XiBmOeF0uW00RlZeHvWOZQjLoxy528WVrfbGJU8E0rVyVrUqVMJOowBpcnQ9xCFaX+bQ8hXY6PPk
a/ERK6KpevHKGkpVqHTYm79jOH9bp12vMNZQcghN+8LMt8vUFIFs057UqCNJJZfqwLHCOZTvwJ1m
g+coDHYiKm3lxR28q3zKv8Pm83X6d0NjxVqJ81Lxlu/jlgiyf2EgqFRK5shrqv5DrdcbovwAS0dL
EpUp+7aNG50viEweMG7PI4UH6euOroknupOjAU66YRBxpezGCq2E76JypULfJ0n9vNm5LkYvapT9
j3uOjpXyBEdhk1oA35m836PSIP6Cu1e/Zzwu1sHrrLedcf4V8K0Cp9UvwRkDRcqwmOPPjqJjUoun
Gzc5DoHYh8BV1hla6lAgr002wbnEfS6sgZX240nXVgz5Sp/CNHFUxt9QlNU5iM4OLZ/55HVTdwUU
ZV1aX7rQ6Q7fwUBcp8zphb9GG+mPbpUFSEELSARXy7wOSfWrBneqhRpPODufwBvPpET7ne/uB3rN
kVmXWuIXgGHEEWAO7Yok/GiUi9TL9f2cDjSeX6zRmLc708FBQKyaP1NUW+qwQo0ouPPvS4001VKf
c7IvvxS/4HvOAzPISXysQcQbnivS/+slBtrhtY6aYo92PgEqJcGrXfNnLZd2ipNxy+t7zma/9cGh
U3ORJv0ZvEhebqZhfBGzr9qQk1XX7tYa9PPu2Ab2DKksjfi6/RPPGa0sldIe22hX40KVG+BnqoK0
JHZ02pD0OnPXCKELBW0pLvyUJGlo0YVYr0GFVa3D/rbq8fOsdSrayQ9C/YTasmONd2c/5EceMyZj
2JtT6Tdp1A4XtfTf4d1X/aJztR9Q0oYAPsGLs55DUJ1iirhApxElBxZ/1PdsZTrPYZ/nASxo/bPT
DNzEwlT+NCq2bDGj1hsLESjE1nlDxn6c5xrIvZhWx6+8es/1QAdTXEGuClz2t1ssc55OURBMIvyr
0AFMj8WK2GDPikPLwOuFs1j5E8/3e4bEIJOre1DXelpYU+uiObwnrPsN82EBENZbqiIlmN98Qkxy
IGjh2ifAhZdgQhgJWfVy1rWmg1oqZyLPdbfaYLWzw6UsnxPFVb/TrUkGCZQSJNonEH7o+aOAmVKG
rQTCPyGuB4STp5HO2OrfovaJ4gDCzR5dE+q4ZKkdkeXoexffOFMOfSX5VFK4s4FWL8VhzN+eAmlq
BoYOoZBf7UXfoxNbTlCIma4Fl2Qa/ExAsSLNsljdxoroQF5foL6y9pll8oxhsjH9C6FhsvkREsQB
U/o4GZwbrPwx1orF5yos4BrWlcovhBH8h6kfPL8H15fBxsVyvIHaghHrKLdN2SvhM3XZXvE0fHaD
C68gWpSZZQYEqhSh4kmeVtP1GNoTbfRL4qKduZVlRLLBahCElYJFHMDxLF/AjgUiqstM2MTNXRAf
OH37ecQ6BoI68pUXoKQhexgekozLZJuIP22ZmxrGOtSFEvj7nEzUHRbc4SXHJ1DX/NZf+9QyceAY
UYtL/dKnEuUjD94HB/WcPUWCcLVJcugZq6fsIlZ0Fr+IGHcnajfM0o1uuzSVYZR4pOOwu4lyXPSX
0uh0xoQ/CoB0sdUR8i9WOeNiM66Mx/zmbC3/C0L09tiOD9ZnoqU7ZYxXjzfW7Sgen1hHe2XDfjEQ
I9RlResaJ8ZsuXru4E4TIAg5C2gwru5J1osenHq8aGC9kEIQ9n/6kmkehzwAsfAKY/YzWtd7acmK
tqyhnFa9uCouwthNB9r+yL4seo43gGPVe73ExJSTmvIleFdjoMt+sk4VD1l+MyE+db+8hEHYmUu5
/DE1huQQX6r56/41xgAsyVac/iNjeHEgBMDzfHq7CojLdd993W1PkrNDFPMs7QIexdmaY8X+6WZZ
JhC1Hzse7bq6Y0iq9+OpHqiHHNkRvK6LK1DH8dkMMk4ps503kFbWQxlJ8BSP3MW5c4FPCzeMU1CJ
P7Cbvakj3OKeQvXdrwOJ7IR+kpfrLM0UMg2z9nkoqjBpiRJN08ny5f2yr7QxQl9S6frLT4v/o242
mAg/YloamZBmpBDVwlYf06D1Rib7WR9r6X8fA1QeBry3Mqj7pzxNJw3SpVj5fvyyxs4OqUScFyl1
1TtvTpX/jzRHmtERvkNf/e4w7RsbwBp13MfnTIgzKfN87xZM28y6oa3/5s8DyA+TfiWq7eIojciu
lb9GG1r4dHfHh43k2LHYvnmo8+TvJsoh6IfgnRym2Xxf2VNfSvf++OHy92JkaZDB39AvevFFg/Ai
9e7BiwCJLXNs9JIYt5QSd6O/F2cct6WKmdv7iIzDuVvtSubqHxytTmjukc+FvLBzT9dWWUu9H1sP
4QEGyo2A5uXMK25AIVNy8ZbtzNrMS9ljnQZKmqjwoqyy339Z50kIo8a+UW4L0y0H1dy3HKbfZ4Bm
bB24yhieFjJtntpfyQRVsg0iwO7FUlylhrU+7HgK+zRwp81NUNn8tmBqW4A7zGgLG8uQ1pDv2lWx
tsCNm3pWoXJa7Z7kfdiq7w/u+Chn4o1DfllbZPR5/PKYzjXNm9WvZc2YxwSXCOApYp5fZqyQhVhL
NlfXS2xoANGrUPbVMkR8lmyt36hGMLCyKh6DQ6dEa/q0cGLgOavvI4DnUr12U35rRUJk8EAPeh3w
52ox05oKsVIGCDpDUwoypZ1XgP5tt+L8TX4FCPA3jvd09aZuISTdJJd6PP0gB01RKSYM46T2mwW+
Owmf7Qu24JcN7eTDEh5XdpLaDR9JcalspUeIMgtDx0voVNs0NpB+vSyPto9mV+G2ZU6h+2dX9UPX
LlSaOfIz7ndlbxlcWHTVZaGcAYMRmZD9NrTEIno4Kk7iuHq+v9QWdi5TCCRA78SmHfqrh50M4ZZr
F9sace+7Q/ZG7L3Mcrnd6o/bmFsqb4aPTFgB7/DcwhOD33jyGDeje/3VJ5OupTeZeqIT/GMToOgG
Fh3FDJ8SxKj/T+mMSvo843OAm44C+cTM4UoOR/sWGriQOtea2wgK9zr3CMLBGrTH0KscN0Necyhm
qqcLOzHHeEjoAQE5Mz4p4WUEzV6YXI8F2slsft6phb+1Nn3Rk0IWLBSdiUbsInUG4bgYAaXfzeRC
l7XgND1k4ma88KstP3/QDhb8vpRTIjBKpQaKtc2xT/4oGGkUfqtNq6Zw2yQyiQKjsrpkS8JvCDms
GA/GgiwbuhuEDpFWNOK+iadNSVHbaMUh4I6m96yj/xfwb0HoNGSqzMtaJZp8+MKDuT9zhm2h3J8a
Ywyk9ADwHTA3ESZq8n1BPdzzES41B+IWdzrUvfEaig4J1Oxiu7i0UJZ6iESqAmHiXCjwwWFusSUG
MM7iJp0hfB5MZEpgGY35XlT7dfDCzQknF5xHDOA10pNgvCzackIolfEL3RIX34gOAlGMjSQ4qRBd
PV0JkOtq9MDuifZItLtG+We2fcCmndkmqy9+p7+FmWqkBVhP5ZxduwH/OsX93I4heR1Gs2r9WuRQ
5WTAOTEHd0d9R9rqL5QFN5GRiEkLh+YMm0/9cLtfjJh5un89OjuaHaV1CesEt/+X3rzql6RsyOxl
zrY7ufERKajyKoCYLMKBBOCafxjGIguix441hiwda0hPI2w032HIEhKEjGfrhd+VlEM+QwSewo4g
/YnrIXnpN3gEnowjdajXEwkr8DxUuFqo+2QlIYQ7sQG3snPSXFhbwjaWe5sXIv9eFjjRLEjmFlqt
GUC4ZN9RtLLrX8qqvzTVryFFevDYDXFsaoOga26xpU2YOx01TD6kfdXojsbwDeuFdy0c8bM5zDyd
4Wza6NOGbAxuT6czXpyBKYHI0p0y6cp9upcgcb+TaecC7BFM368TEtpsvW5uubOyUzqFEzYa3+oS
oq4MlEAvTDoDBbrqoumu9YQjapgIEgK90mvJ+zOCJ7mvuyi9FexUtwY6AyuJLdQpsHMXbiZw00lP
4ktFhAthRrHutvZ2DHGbzxtn955tlWvHcG6gwBddSMyCDb0TqK1fVziH7/wLc8B4g9de+J+HFwtb
Cxu9JgSlZaYan+AluaWR8IJZelPjNhm7aZgMoNiCL/AThQusmagzp20KpeHN7bUsLe4UQ/GPpHWV
c1L3qyI2yUOROEWMojCx4B+AMELEDE1jf9ZB6b7FpcIbT3UCdUaEbSwwY0ABGCA6v18qm0HT5F1/
BiuRqglZN+Ke7CAlxZezSikS0vr/H5D23HNT46IQGe0xg9pYuE1dXumyxqadtJVP5S0IcNW7HBsv
Zczvvyg/VhGWONKYkbGYmAX8ztxeLMO8nKgWtuVwKIcRhqYqimIh3S/VEdsRmT/r6ve/A0RTCEn/
29mA6GhyjxdeZO9NncNcwuWHgZg6Gnss+Z9plXQ5C6wGCjxdRVFEnTqSULN6m5GrCxUi4r9xGfrt
/Jo8+8QqI2fm93BC86j+RZBwd1ZgGKlBrxcZVolBTUOYlGrf93Vt6oCtOjtif64utjUdg0x7kcek
N3Jz0ZV7eiaBSphKn+B4JS7CtuM7xcFh4b2AtwtQJOJZGn323qUWa5WdZmjo9VpzNue81oIzZeJU
ti7XtQxmpwxaT9HOClz0duFKrfTzwLqUWgfpP5Po0dX0GmWBRGQAHIZvv2nsMZRIhwq9Gm+eZ2N8
SN3SKgAAHGq4B/KhHFbO06ieIPIBVWxwXA+VgQ/fawSVVybYCtHj+cM+fRpWsaFb43+gHUhzF5Zk
2TAM6LY8tGqAqlJ/pgUvGfCsDRfpLBYXrl5i1yxBjoPP9/Tz5nFa98G5F1tjCFSR26JDOptyMWdt
pc/ePDCsH/XXZrZUTFEJELioJRo9hvQjIofmHA2A4uoN8PxqxgNE4L2wYJT5YQDw4eZM9aU64Yto
gP2tXUFR/t7EKo6bCEGltuJoE9Ei1fvJHNjbOWr5j6AbtkKE0nF16GuCAZi4M/01+OLbtISv8uWb
QkdgizLE6/HCvN/Q5nvuKbwg6FBdWP2ydUdPmMz+GzVq1YXrsX1PWeP3h5dTnTQ4apl/DOoXB6Tz
/4TThJV7TeyL8Y6qIisGTXsr9HZKlL/EDND1r+vXBXPjX/+zsJG1cX39+1yIeCuu1RPnjGnKex8M
0OHuXKHOzxYw4tybg/2HAzH7klIM1jk6GObj6UGuZNWU7MAGf9aDvtJg8a3yvFVOne6HzzuBqRkR
scCOLzt7vWGc2XxNNO/0wKphEAIyU/iOecqBYBZ3dpBK0Ff0W4CKYrXGmuDYzvOfMQuQheGdFjbC
oZNuQbTMf4x9AvSalb7W6z/YF6+Ixdt4ITw8N4nXwaTcHTM1MTZE7a8qlSFCqN1G/3ov3oeF2BlO
FAj5ni6bAwSS4vBN5k/lOephxuqyCW2GN1G+BnNVXc/iDUI9OvWmydx+g2qvAdIJatqBmxdJan68
MifwfUynq9dh+lJ1A4ieimX9puLMD+kKFoss1EVYBnHKeSf1qUHg/jbxqN9c8SZE3ouwR7Nsyk0r
5TZ8UwitXJKj50Xkl1S1LpBS1m1z5+2eoYgO7NFABxxEJQipBcD/6psZrDuljX9sPtMIoLlURx/w
ilYItw7GYUQyv0WNDCU6DWJhc0YT3RT4tjS9yOaY4GT6BUpqZVd/D2K7fIw/CWL0x4J/x2zKnpZ6
1s4/DYXrKMvbf0xIaGCyJxyWuLJl+Fp0Z4pfDF3xawGtUeWHEwThUgPT5Ed72ik/LROqJEBydjUL
8SkAJrz+w6xivTMgmmkSjX4/nuY4jAjoy79t+nk+VcMGHVz0WY7BDvICfjLWWVYfXKrI6caoWikJ
bqb8eXcGzwLe6Qf/xWgsc+STpkqA10TfPpHjmR+uUTeyKQX8Go1e5e3myvidAuASLbA7GpP/vFOv
GzMRmowMfQzLO6SYLRuECIZRoVktC6912m2+mg0qrRIBkMvENgu2EYP05wqP3EjAokgIaOtyZYeR
QSKn1H4CZfZTjyAp1oOhPs6dkj8j/pl+vzrAEkYeGH8a3YFMzLfiKXOTEiSZMdnewEdlFCDy+SI/
Jw+B/IHT+jT0GIh/9amJCOR215wA+ffKSPM4kv3hec+MyZKU8kqaIjRvmCeSOdcJ8/+/ExmGTcwD
WG7FC4zyH/8nAPZBczmI7QiDHMYcxtOW8gsvVYPvuXmEktQFFTp2cdDyIbPM60tpbM0BIyt04IoX
CZQAnLoW7vl+1VwOt2KbThWHuAETFjbtx+SODuu3VOx2DEukqaVuqtIhaosYw2TYD5hfLfjosDk7
kImXBZ3sGVRFNBpPAjDPVhpKw5oWQa+nqQrnjSUzOwNcKeTQA2OX8EFsxZuhivO+HhgIQGUWRuae
CdMSwmNoSE05R2E9Sl5bskPusqMyTp9xZ0ej6sBTyxROqZZN95Zc287QTcon8E0yyDQUZyXFUXgG
IbimJVsNY34LXMgnqixMMSrfwhnPNQl90HA+B6X8/4P2k2RtfRkkitsNYCpglbmEXL0+9aPdTFCO
WhgXQtzl/akz9y2Q7haIFkJZGPZM3LfT+zF+VmEZOhta4tZAhfmw1jDfIxHW2lyOzQ9peP8X/VOT
o1le/w0A676VMK0B7QN907xxYmz5ahVOayv71Ut2P4lu3MyIht9egTAsOGpnhGJeqDrgerpcBYth
k+X/xPJGZs7s9G681OmrgfTFpqE05v2a8TcNEWLZYYgBs7Y8f5JbErSYAHxmzdaxXTq3mxyMbDIz
vNg0vmpMQ5qF7VyZp37gdFMSINSLNaVI8JgZj4fcI+Is++ePcCvHAtp3vXd9cvF1EBWS9DIxW/JI
PT4kJrUqSGR5OeF2eSJWaoVynAFko7WWmVuBc27GHtYOkAhxafck9b4CN2iVQQ+Oix2gT0Oob8S3
CjGA1uqn3FFeL1RIfNHd7PZoLwyf2dpoo+ya74ZpLtTN95a+j7MOz3ygYak46OQ7aRt8sxlKexEA
dou7E28l4fcYkwiiHR3WHfzrRr7i448BSMyT7Za5QdeiKCbT5T0YSUF2uTCUV50aBNZvlBSCBGzK
WQTbHpKpf9PqJqXrUOftTzjRefPGV1wZMi7tt2E/ZZ5yPgTPKkfUAYEIUvb8JQS3HBseKEgECRa+
c0+WFjtlZL5agUhUO3qfxaD0eI5RyAfN+srUssY8lbcbz+9UYwWa6gGB+sib3y1WBjNdR4P3fP/p
AonvuoLFeyk3aoksGNjlDYgg69z4wDQaw4FlO0sYnTmurHhFv/AN5qFHZp0OLHia5aV7YnACR5bK
yZoN3YPnvjTRc31Bk8U97GGIINxKMzazf6YoleLIDlIGEoJ9Yrs9mR5L1/2AA8CSwnbfVbNAe113
z5lVFG9ch7bAHp3n1/vFRCZ4lxc/MFjL7vnF+vUrgxdTNKfUtVXPLSpww36rvHlHHSEJ8j7EZoGx
F1QWqFBKCJqZ+Ggnls89imWCq2hIqtMGmUpQYKnXcroi90YxT5GJy/5Cu9+QTPjmhF/FGALo/atP
lb9MngnxIf9Pbr90xfHdA0oDh3NRGcHHF2FfOxPnZI7zbshffdKFPZ1mVFd0QNC/F2MyWscuoq15
dqAEM+aEJsIJhqaICeazfmb0pGMFx2Q38a/NWl5C3pMFRVO5ud6NaxQU53SEnjlSbw/n59YO7S+P
yCWvMilEebBwwrJ2A5AUTMy9qnpc3DrsGaGS9mtUAN3SZyzHfBVWNhv67TPSKeYKC/vKPaZOM6y3
93jGnQC7V5FX5ujTVIUxQq8ZLbVMgP2168uMzknKO4bL2IUG7kVoKo5fAMY06acgb2666DP4N2rC
9NLcmc4cq81F2avwdvQjnVli23ISY/xbwebC5m9r2Vyya+FjBM3R25elaSUhyIxcTQ0xWTUk7eAQ
V0mR9JNLYNGB87Jo4mXOgi8eThK+uQatZpWr3qRNNxHkd9c9uiV3dsvo3wYjTpKVxxZuoujS9Wo4
iRf4fZ+aRF1dRrbij/E57GMgBpQiNQx308xZmL1ZhPbjzM8DjHJc7iBLWa9hk/3pAMgaoOrzmTrl
Naylz6qyw/FTDKC2ONm0sryLA5UluTlNPE2ibm2uG5TseFKc9hY/VxZOg0/HLO0yyITOAS8iS7oW
nwHpacYLKp5V7nwwdjRQ4HHI1XlrqX1m1OFinz4LgsKYAXtKGBmKypMKx8bmhDaf9z1KVwqnC0ZP
egEC0bRIRsPQFKwtge0t/PPdZr3Z0uCq61YCVhNHF0umYnu4Kj7IBzPIa8Q0XecDa3EiNwgwnLZL
fhSMtW+ZYUUnHuysRRYUOn91XvhMOGezmYFWA2Cm5legi9MvINoq925AVHXvmkP4prNUg1Q6pnaB
I+uaU1CKUhUtP/BnmxvXnPc8FFONZi44UqDK9u579IOFw0woUfMxId7J/O2+lqJIpUOGe+Eeq9tu
/Qb9dBzYwJ7rOHYi2IDuyDaEhOgizu+fzk5QER9TrT2gzFgYdrxTuIIyKCrfSg8zYfhPpFbBNZoU
SBp44JrHDRQVmuyTn0LmYiPTDGHiSq5orj1ObzaFFPUrnsFtJoT0VKv2WEJd80WZABj9/x6bvhv4
YiTQoXVG5LRKsuxYJ8sBJky31z9aK1EsWyryDMZ7I7W5jph71wjJGEYKvFMRtozQiRlelfpv+s0k
7Cb9lVp2a0JgBhdtiJ+qtTtNb7o8Du0PL1MuvF3RFlFM/dy4oZh80UKHzqgK7QxkqKHDrbaAEVzn
baX2whV6gmS8F0cipIZ/Ceir1EL5H2+2IoJ+HhfuZSNkMAbhzgtD5PeoMAcAvt6p5/TacEfb6Ut5
w2LNeAqvqMx/jPaZfaX6WoVmUar1FLxK1dMIjxeBg/ITBpMlF2/JKIpWOqoqdSr1cUm5611ANNIE
P8ll7O+JcylLw+4EX6hln0WcqsuCY6IcU+PO0V7ETQsrtpmB+PR1XMsJP7gVS4NaCGlESnHngNtZ
1pFdfCFpgOu5nd3mwPjH3aAVc18Z8tW1VzPY0mxd31luldGhUcznLQeLh9ARG9Ic0FXnrwn+xDM/
KFosPRlQoSmmPp7z8pHzf7nxwIgSpLsjvR6LwKczKIi9cxTe3bLK3wFgGWAQt5skaZxi/1BNENol
/LSPG8X6MGxgIgLUWoC6gkwrdl4pndf4dYvcVZxl5rEmQs+NQ7RsWkzUnEaSJqqRTGeL4xiYJHRc
UBKiHPA74v9DAQle9PNgRAqdhHLy649SLoAx4n8UI0ndxWwfdtp7X71WApssHpk4Q/8GwmMWUKKa
P6ClZtRS81PM2H+Wfsu8QR0n25XtKnJczhTQiZKYXat3dwOhvW+OEr+Guc0iGBNMTpk6wYfLG8OL
kA6kkj/o+W/WMRhIQEXEy7IDdBwMv6h9/CuImBVnZJzbn547Vsgll6bBpmsVJZ8zvo7+KM2imAaI
WphseSMDp7/8vIrFKl0e9Ag9r/IMflJRtQPZ8lYugyFTlekRJdITrnOWrHIutSzmnWiMGLcxs+8c
IC+ULNa9iJ0rfHrG4sd1BsfQETR9J93tWXodW8Z9G4dG8YuzjViZkUpFG9QU62cl+3sexGZceUre
7bjtKIiKpQPwQNGVpDQ3wSkiPcmXX6qiDetj+RYAWPXttTtbMu/HV0UupXCccvqTKQr8vHHcGPW/
W5MAM4C+GH53RBcEyFyJPv+6pYnGfPL5m9F/0wNXsXlrYY5kfLP3PEoTdhm1t/DCV8u0F2aEqW3L
FDu9pFA0ZpvFP3K0XRoS38AUmxx+KNzxet0ONtuUuZVZACKtw5LJAkAIFW+i3+f0r5lyafsuLTTM
knLWIKA372kmqCs3aoDfv2VKzRzfF5tY7L0KYMzsEg3822rvWkNdZaQIx0ydtfzF4mMkP13zq9aP
5ijKx0KYJ+rU9JoSQFcbC89R8K7bKYDY0KkiiC1Dyx5XrrngSl7Gcs0BpiUFCVaT3o3cZbYKvh3u
idMkzBIajWgA6G8QPaYIgKYpPH5iYN6/U4fGLIepj+Ztc6u45P6dbcz04+mLnw7DYR09H4ujvLa0
JmS3ywSPAfYkRivVMAHDQi56clyaY2spdlR/YzfsjK+PTVYrruABWGMjPLdO34xhIXHU0tmpIgrY
mJN90i170k1ya1kUiFAohzHc4IfdeJPxZpnx60oKtH1JYCSCXK5aER9qO+0mh/topIGizSpFjjfA
MHJigViD5UfaXaLeD2Yo1XqmftmssZs2BY0fZyAm+u/124HGyOtCEerw30yywLsiZB3pJ9TTn+WC
1gn8ybFbQwKiU8fM+LGksnH+WmFgtRTjkWsIDtB9HUGB6aLd+lRudTsUoDaPQUusC+VA4sTdY6N+
Ill2LcLT/JR9hde8WjIGJKMxIUFGldMb3pJKvnbjETP5xGiPV7zjI3ieSr2LBdJzxv9g48qAngiE
uACGMFm+AWcxv72LQ3RMpoTP6B3mRULcgmlOE4boIC32lUOmGfKKAgZqd7U2GtQI2g7unIvU6ZZy
zGGS7Il5yMmdxpophrxLjKuYk34XiKTFS8kxXiIzxEZo6Q+o/K6Cy55zJmkk0LOkNku0jr193a7d
7BGjiZ6gfcI594PVuc5yKlYinkQReUWT1xCJBEyyHZW1BUimCli/pb/c0AfZfNJOTxtk1QEEHb2M
+SnI5mUy4l5U60Pu3n1zzHgP437n5is2RbMpLkVjLBhtfwoUb/68DNm7FIpC4gSbwQQygIbkFqsb
F9amzNr0Ny5YGDiMfNh6SzN1CbILXQQUbH//h83sxPBHYYB9VGt6AZT3Tcb6H/7AeR+qvFJE6ZwP
g7lARfJSawlxjQCTHXYHL4k8QOImvwFqbXA2R8ixqHR8YW5fioIP4AxVDoNvYxJNzHzHxBlwBBDW
6V5cjXYmk4PaIBO23QRB2lMLE+uOKoAh/mDY1Gf1xGI3X409bpWo9ftXhcQKbArXHKXBVTyfUQD7
c9An2o+ddmbRGPc97dYLsxL0oHZN8yI2GPgRG4+TucPzK5uxO1goB1dxlcST4OeuUBX8AHUPe6/L
Xyf+Pfa3dt+Dj1QtbVbUY45pTtbQqMZoyFeIMiYiUBaIofhn8M6Er/SVN9GA+rpEUMDJ90q8+hEY
TF1t6n7lRsHqv/uusxUC+DximTjUkjrPWX5FTkxKbvEUaUi0aBtNqdkncY0eRa7FXP66CMjlN/2C
5fQVS5Rc5ga1+g6FMNgEtKtKPqC5x7Q7NiUezc986ji0RzBt/fuMGJf/qkRYXaJCpo6dJard7mT+
OjZnJC3EH7NhAwWgHf/2w5WOfEsTV1p4or7a/dcXih0z60hh7tS3skX8PLQm6hiQDeOT3cnhrMph
MHregAwmA7NBFgzjTcF+Diqzr2UToSAVAWBag4pkFjD4nAzSCdH2RLlHWx5oXCgNOFachfsA0yAp
B/2HQd1dZwAT9+xStvbGeRZTGbJDmR7Gz6JGpbvp696pcwJlpIKqTDhBR5XiqJVh5ioFDp0DF21k
WRwKhJLl94NWihYA8dEin+n34Dgsop2cGhvN1TwXXmcplzvg4fc6FYmXlRg5URTJD+eqFo0MroF6
EAmbBcB7sp3jViRVbX6XMiAtMcGhE7DfmPXcU2x8U87aYb/JnQz60iZ+6711cmtoSeDTcm+Axwa+
ZJY4BkwhEou02jm2Q7IDcVSzbOvrZuGATa8xK8wxRah0MyQ3gasAooTbSiGBb3Q22m9AuV3lD7iR
c+xhlnvHnTN4BBakXu/k/ACMB5aLCOX6cJ84TLEKqZ/MZn9SrC4u0cxy13FMSzYEfX/aOfeyPHyt
b/CHLHGLwnTEuFwuvqCcuXvJ9R11+3duP7GVsMqki1cblcokzBhpdG2Smie2OZ1Mu/SuIjhXhVsQ
qkXz4JAx1+1iCOIUOWs2itd/1quxeEH5FwiXDg7XgmICIUDXRamJ/+jt+CClUSJwU6MkPvPKXUC9
O/8meUkgV1XhBNUFfGDPWDfpfEQIDGIZdysX4g4ZQJvp7v/aHSNxGhBeH8ecd9UiuFTizCloczSY
Ui5sFL7/it4GwPy2dVFlwapDUAHfpltSq8Vpu/RQKwFSuo1JtSBg+DnDHC6c99W7PGb+AwaERxb9
UhmdFFRSuRP1aAOZfZz+fVJqkZRiYVpe7HQxzXHJmfWkUlrBXCy5Dv6msRQ+aobsqZVgx6kCVWAZ
aBNu2yIqoXXWhvPdsdzFaEClQ54mZquuE9ANk9kj5e1J/ZsGm+y7p1JjMBYsJCZfEcxG/wDRrAVo
oEPpISu5FjYCvFEJaCRD0wFXOI+QjwHIGO7p3uCiT8hFN8qXcSEY2wyqKgIu0fx4SMDm/In2dWGD
U/GPapN60fgQc4KLCQgceS2AtVeIFZg+3+Hhf4Yt6Kqzw32L56ht2lwoIuZv1zSQPOtwfQ/4IHQi
YbLegUCRdS1A/ZKqsTIC8Q5hc4eM9PCCV8I8YxKM5wY5Z3UOZ0QCHuMwHRvhMobmahPMnAHjBUF/
k7VuFpndFg/s8bM8AkgilOJx1EkAUErUPN8DrH+fCxZlbv+d0+dexBxWpf1VZbWd9w4cQZxyn1Sb
W1pYZY1gn2qC0FkTxc8jzh0fi48cRDGEJnbdnGAXfVO6GWU08L5e88BXCu2bifUU48c5V5PDdUm2
r+SOtCAG39w7atresDbH+A4AD8ZIu6+JSrNOXgrN0B65MM3KaLWQtcDPynY1SuusDBOibR5/59Gr
p3C3mhWVCgdnGIfC92lPMDQhXZ0pmBzL8M9kxepPGl/CRn5gJ31xsJuiFpPZ2hD6CWdkAZhtLFIl
x5+74gjpqe/gLrWwHYAufzz+Jgz0jrv9wRDn/PCJ/uUqzct1cqE4kDfdSbn/LzDydgugMtcTLhLL
n3TKTTbK1uHTRfk6vAqHRFXnpD2t+dcUU/HkazPKUYuCb3p3EjB0BW9LMQznfTvch3Ucb46K27j+
sAt8rDrtzDcvW3GxgjgcC50Upe52a2Lc0t6WM3UX2GsLpOJam0b8TJR/GWVxNxeiChV5WHe0tNwu
G7+910eBgNkHGpOnagGnjkRNOCu6peXkX9eVo9b3j+UTrT+q6KG9zzQst2g+uoe2AocjU3YofYob
YzzdbE9Wj7t6Um4SkiBLElYJ1aXr1/T+9MbgBNIv8XV0EoUN+AKIBLFZzdYsjIgX4FjTLOiOobJQ
wpJ7jpVBzFODvLJIt8AwJnY8ohKQrHWQsjgOOCVF5o+6XUXA0Xe3sJx62NmLf8efA3PAGJQHKXE5
rRs1aCZxW3HcnzuZtjK8guILzmNrmfouy/RVaT3RVboH7YKUvK6zZLohILQZ1q8th1G26rn6S3Dc
HLpwfsMWCpiPEMB2k63RKtNMFK/Sg8CuXMj94EDy5aTFGj+zpI6KZlrFw8sNKh12Zd2rp5X3S76N
MMLqbaU7MNHtDBc2BFnPmU7Z8B1R9OMv+HQVvmM87vADT1OfFgnGa3teiF2PRYL+sc5CAklWXj+S
EsRxbDPfXgUk2mgD6HyOQ25+QGkRL+b91thMI8A6iPElWcLJLf0P8GypLXpRw3P/kD4u9Vq2F+xo
AGNidm4MLPNyifbw/0O1HVJiOpGRt7Zo5G3fs8pu18YJCgQn9hYKs28tf1A3vliYPl+rXpwQbjg2
Iddn9ufBHFslVjreenDAFYaY/f7e0gi3WOz5toi49desfZ4aTjIiA0r2pzpOrbx0xrhSoJolKb5x
71gewU3oRjuHdYBg+ePJogMu3dFepUYmtXsVOHWYD6yhVYmucaq2YJ+qaHSYNofXIb4WwY3IGu7Y
1+KW5DV6HUIUMC3oM3N+oNavTKiH3oJnr0cUsGdIyI2FV+5d19p3lpmFL/JXpf+lT2yqTIcbwhSA
YBhgMIglX2ckpGw6WW7fDRAHyojcBB+S2SUMnqewdsjykiWCfvGuH2f5XI4IvofWwcqWlj7QjKbh
ZW9u2Hz5WDjV5q9AgakhYl2UE+YMo/HSMXMfeQP9/O/5fzQc4xWd6ls8Zoy9St425LIFEPNm0+oz
lLbgdqBeoRHVVpmQew261S/Acb7qbqfYK8lipEMBxKxqTRmjdFUk0DaBMRwOqWbxO7LBtg9kvpSM
5xDbC57iyFDnHqgaUU0devT3pM6rLIhFv1joPqOYeHrK662AlZKQA95gfuR313X5o656+zpf0J/7
17PM3wcUv9Sm4Q+mP/KwG7aQu7mNoD7he2XCmKuUCMgWWt3UUxXYi0i6fqt0kbfgBty7AWTyW75A
L34DLX1q/HqbboCxv2rtquagriONRaHu9f51xsCts77ELIgmGko5/Z6X1pGZvSTYvsfMmYfRnFS/
k6Dm4NSOFGPsHO4WZl5Tbg0kjlNjF+Y0avc6/y7X/LEUAZxPNEj8vYUQiaZgXiyZsfovLCOVXomz
7yNj19TD937Ej1UtvWhC+5+y430Dkm5Qb5H4FgOIUUjNWu+iqGKunCUc1EyWQerajbEbsifl8uf4
1KTkJ7Ux6Ftoi1JIA9WZAtgzPwTAQYsHIenZ/L3Sq1ma7AGt1nM5WkBkbnDF8OzgZvkrTTjE7rJw
oDJ2RPVkA6XulqP/U3PPp9Lo0WQYn+cyaPb735PHhzNZeFtWWbwg6Dk8DjR4611CoKsMPW0d0nmH
GGDQ3b8C2oQM5W8R+GUA8SsvaQNw66ZFfYZI5dFqGTaY6H+HvKYpDIDu9ZDdHth9BR8BELBtJ8VR
gUefzmeGwEXcOBTLzonWW1BhPPAf9RpdmNJNG6s3cvAWdXbM3ACR6L4xUW6uyTIWuEu0IJLzGsRX
UOfvfGZOZMPYaFDUG7Zf+4aArOTg73hbvcVjnI5d7XVp9pJJchCoSaI0TAZogMBpOYInOaBXl1Hh
TNtpwjtWum9fsOIRotADMT1WfAQRoq0JjYKcvWVWbEmegAUi9WOqQPQKlb11bh7Lz/Vg9rPVVU1x
2oSCgmObSufJTmfg+gyN277WeCBeNROQHijSyY5y5yH9beSvXwDEll8IHuIAh5VhIspi6sk+R2AG
cPDh/V5F4w0tIMdDy6ceO5O/P3l0oF/TPsbxLXjp/9VXNUOZoTDl+qrbWMH3gm12+eVM8cwpnDQm
TuVssV22swVmntl3yx/BZ10vefyhGdQnzdAYrx45lHyBbLa0bjOBsmlV07W4d9i8y2xCyEArSkfK
pmgGPR44KsaYOVoVMZw0PZBbYAEcUf49uLx+tznVp4ii09JsYMfoSvbFwh0iWCd3INFMQUL2WqZF
XdMEhAcogNRfDVGIW/5DRoYOtN4VOIzx4ekBmB4uCP52hTv6DwhMOwiyX0rj2B0ZqVIFxb5A5a88
at29pVgu0F3CmLyi9dV7CNu9BJUAxC/D6Rmr6/fIxsCQWDpOmBrfbjXbpU5QLRXXvuw2k/1pgksl
UiG9PwqvLGns0NH+LSIGLBvjIOUSLgskKvI8MNH6yyGOWyMO+Mnm/OFj5kHsmDjzDZhUQkx8zmsN
+KkYLMM47lqNaEkQxbw1OrILlQ/wkh1/6meyXCHaPPHO6JQ0dbQEeqZ4iPU1B3qSAXAu2ePcxI4N
SModP2M9iswXjUlrYXcr+7GsWw4UC+IbYxcy68z73SdcHeIop3HxaW4OHWXtzouY3qMYMV+XLwKf
cG6MutQ1AyblrS9+/r+if3uPgD9gZm5TJr7VpV0d/nl7yb5fYjQoh5VbiUs01ztthRlyM15JtUsg
/vcLnk69ofwo/+/KGMKqSZtUs3Ja07kzVML0LytfK4DF5wc2f+T7DaFbAdcbA6KqIPOtd+La2MVq
BS3QkDyckE0q/W3fjb2W78+jQVOdIz+b7coJciL58U1W8QnmpmqfDP7Qkz9+u1QWxlUSHwSxIX0O
Po2Ir7BUdnJDjE+u87p6jljBlTY2cKwlXyR86tDrTa9ehDsQRB4xtixKyWWbZv0yrLmgLXwAZEqt
Yv5HDzdT9XE9Dz5iXiyOrBxwqdKoR4euy3jYjtrv6YKODA1RlWraWt3pUPBtvKj8H4fhv+e52A2g
j0r0IQmW3EItU/wFY+6EqmWwyuGomBRYqsjYD8mArYTH0zxsg1nHlEtt2+XoCo0Gixx42WLmE7B7
rtt1vsz6QRirSD7kmCDhCiU8Kl7XxRn5OQG9EIqWuJxVU8xKXIRMWhoAmmR76/k+R/NMJ7QSTq2B
DoVGtBy7HRLii7HdrjJgoF3upsCUYFJRbQo4Nb8xHX42d/JO8ZGVyzRbv5JmP8YNtVGcJ/Ls15yF
gaQDw212pakVZcnKF3HVMxomizlFaRjsVPkklT1p16ue85iua5TCSlLexTSh8YvSY+yyfSFNSzkz
XmZQeteIhXIMcXRO7/1IOwUIg4BjPscfbtr7e9NWB2o6/0LIIDIoTIrUOlHWbSeZqUJlPUphj3da
LLazTLL5OwYJ9tZAiSnuunsZgflU+UeogQMPrbbWlra7eF+baBmMxQ82XWk54jXuhd6/lO4fUJyV
XRGSPYUx/NSf3/2ilKpSfcOIzI4MUEVe4LDk+r5TgWd4Ce9T8/R9H9Xy8wswIx6V7vPZ17GbsRYU
cpoL8KZs3xcc1avWZ/sEq4BYf4ZbdLoPmRGCEGKeqWsPtjVGbt2X6up0C1Q7Gw1L2aUxmwHSGfkA
KBtsQOadmDaxL7f8YHN61fa/+5EnvhM8LncaVffIu9p6tbXZMN+bnkn7nDD9s49VX1NgbRXkKJ0l
A1+3pA0sPiwXySEBrqS5xlQmmGwb7HdXWclcE5e6/doyk2aACPiXQbVA3hQsBoGHV53hjM+G01gY
y5lZPLmFvPi1HcUmoyM0yle+4Eqi8YFrYhHtttvzW083Iu/Eu/nP1PPHtesxiGwausBrBjrMDGJu
3gy6yP4ODaYI2UkF5ZSVR2/GP9+CZgbcjZ2VTY6cs9UJnzGpWc4JOl/hkcoZOHVLwswJgfU5rcWd
PF/n88j3R0oB/0ko8QdQh7f4pKWVs4JvDscYB7Y3YZuG4I+DLlf6Y1JlWebThQWTEBcANo8A7UgX
g2JYOHYvt2PRLI8Zwki756iUylp9rLhK1znIQBce1iO/yiYFTAFQBzOi4nRgg41TA8F5Z30Lzzxx
dh959h/ipOQn1Su9rKdX+MeErA8d3F1JzINONg1GZL5ZpZ83ZDLBMp0R/H2Dv1cRB3Q1rr5LENSC
CV2yZNCPkZOOXcczKRsORCs1Q7glb8N1JSkSAjImcAJO7QFEFXiiaT3r/h+yCnDhGND4ltS2xx6n
dl1CMLk+bglyUm+/vdjm/uOCxGUBDaRJLoqRkqyYpAFfQPf00C8TvVVQpb85TWRxCpNuu/gqg5D5
rXdvS1gH+VrsCDqm8F7CCW8tlP8X3YoauL40gx8lLBdGfppJzfe52pBQAC9VEkQg7rstWSQVwyO5
tbB5UJ00PIxe1Gr+PeTQ2i4X3gaGbtET2ZJsAkEGBr/Xd3syG6D2ltCD6Zf1EmIBSdKKR8aKTmFz
bM83zfi2OiGp+/ZKaCeVVL2ZvVsAiZrPG41lCma2Ca0ukMbdHCCEn5RNM2cB634Wd0b0CGIlIL0U
XO/ZFb0QXGFcCocZZet/ksu3+JZsnWa227RVh5TfLQ1OtIOP+ZQaQj/6UNYA9F5EsOG7UH3FqvoA
Kn7Gu6mXj0ETt/r1+93mMtOPbKaU8WtBVU2ywjnBevcIm+Ha6VR7KTYHcjODNK6g2Ku1Pt0oTHtb
33yxuyaCMwGXU9NuCfLHHMRMRDS6EMKRVPvKnFmVb5jCi6d8DjxfFv/sMUuR4r8W/swcP5nUt4vW
5h4AynDm2oROjiH9+Ud1QMibdfDf1ke/Uqsef8KYfbjEc3eMKQMzHuPMC0WnKM2Lyqsk1qdPj5qT
wsGBgBpyriNeMocsi4R1xyRp/hEVSE0MASLOcNPzvvS8PTClbl5r7Sq++BPOQM/piGTTuuZ6UrCJ
QflaOSFVakbOVpt4kLGiB+AktkXu20h/E5CU2CWnE0dKLJGpUx0LME6rxnU9sHyhy6JeDkp8LjwZ
PGYUvt7zp90XbCNo1S5wUT18pkBTfEcSEC2aarXXIq//+BEK90xs4vxnzNUNIZETtMID1pE7SqJ+
tD8BaFVIyrZkl0p4rm67iQbPnOPNC5C5P9Zjflx4Py/SiEZxtxTE8OVx/T5jPpYWo68r1ysCR2pL
3pWzCSc9/ogg0IGJr3D12l3fv6CaZ4X1sVNaJh8OLAGNJ/3VI9aZMEH/t1XrJOzJ4bbkAH5vS7gk
Migl+2FTHp/M/nlA01c1ZQWYJ/IzCwBTQXrnCb+wD0cyaG+iKawN/HXNecxzGCn3Wy0QVxErtrz8
Qu+nbTN+29lAqkh1GDYNslgBDqA/CgqVV+NgXFsHR66xq9ZoWlNgzHgVIvRNQoGePr5E6JvKxbdB
G4xsf3xNGRmWWCmJWFPeYv42lynR+hoXFNfV8T6d7GuJjVG08tuwiKibh2jBDt1Cn6Mii75V4eet
YczdRNGHMpxWm4vZa69SX/nHZUNmwW6mYFa/qpKdMpOmyU6B6qzy35Aq/r0UqWCK0Be06cIRiya1
Qbpm6rayZ+LTq/GZLYGK8gpj4fqXBTMaRS3RGyCfwWZ/tlaVdX1H4I/qwcynD3xBBmceb2IHbOnF
/serrb7JRGC0fmJJnslxkle23zWOS9X9VakHS+W4p+ooFgCdziFrsuzZuYskm45cXRPfPz94KTFO
0PV/UFFDSvz9h9C/5qVKLODkCwkMVz+3XHxXsUxNTPWH9gx+hD9+pCOEUGVRtINuO0FREEgZZb7w
ypmF0N883NHOhFmofqw42EPh0pq/e9Sgn+p8QrkfJey2H3w3TBUO0ohIv7oCDkzBnrHGXuI4zrfl
eHqVRCdU/XsFDG/Z0juWktNNNKKg92qr9vX6r+rD1br5A/qEsPTk+QmBn20ZDw6xhRQw2P4wOTz5
AndZ/G5W+W/vNL61YU6nCe2L4Q3JWFsmBwYFVe04RdNjxMo051jQ88OspNGgMB7AVqhKYlVTg53g
PtqKFvX2ulAytjlwcP+pPKJwcBXSfOBgIAHpfgAGFKdcp3OcpwMmi5zaOdprSbsPHcmxkoywCqvU
j63VRm4+uToni0Gl8hWbPFG8j7itqx3B0rzG99ck7flo2aVrB6ExYpSnkezeMTV+1JDcb2J3uPkw
dwmlhMvILGfxLO0kSRUbEG2rZ5jK3q/fV37v2J+Y/57nxoqc43lFgkTSYscP6WxqPRlwox7IUAZ4
oDYOYdKmzNuaNi7LcFzLsiRbJp9sqSHni/EA7mCU1hnFcunJQsnlaaJ+mlrpOFhFCqfAWMOGpHP6
77yiGgtqJz5HqnsF46mqBzsFj+E8A6LLd30LcwWQ51I8BncxwgeyID6S1CI66aZrSHP/zxvHoKqG
8EVISL11Tr0pbWZJ2EyEbP5Wog2/51bb44QPHJLQqWEQA6IbI60HUtYAn8zWhik3YZkZ7L8Smyg9
k9LkndOKH2ulZ+k36/QLAvD1Z4rPxPRNihxBKaiV6MTaJUtKbSJNOqAWi1YMjHNpANzidWGriUTr
w6iDTq5qDoA2ko04baAAxy7o507XpdE61ltNwo866PuPnV+iRKmle7bUfsOX8pUGK30iCjsjGMyE
O1vtDk/hW9wDAMISwZomYuJH56kd59BPRI3GBa0fbo6uV/ISOQU9Y2J1uZX4BlPDqSrc1EhUeDQM
Hr1cAWBIpYUhjOd9WHoDISUgmdwxo4NaM1QAMB+ZIJOYaCpNR+oatSPyby2Wcht5f9uVlKKGNAdm
QTpwD/YotBYX5FzKKwLT/2RKw5xnZErz33APEzR+o358evrcdNlhQyNPr6ih20qC9o+4+GCb23sE
QTA0m8tsZETnhIaJecyvx7E6/Fdf9ovXlY1L2/RfqWB7DL2RkiOKBoCc77Y4B977RE4QSbmdHrgS
o3EuzMg7wzpI3ivVtpZJnH32u9v2wguDI3bSiPU3pLhATR8puuBegM/8GMRRiTQsUr+Nz35/uzrF
m6qOyWssL1JOC6GeFSWVGWG2aafivKZIQ6gtQ2yLGd2IxQbH07bnMsafpUhoXXNBd6WxLGSYwSFZ
bKgbg5v0t5wMNrs4A2w9+vkQeRlbHcr6XTBBOJGwtG5FDwaEdLgla+lkYnMwiUIt0KWFJhLBPptk
GMxt3rS9KOzdkKlOzLekxfqvVOhQNgMrgq7ebdOHMKk0bjT+TEwUHG6t2D8IzDtrc3LMMyWq1Ul1
dBIkTC1rvQP24cI6gHDVgC/qcueY1fqTat58GI1gxFqYKyF3muFSVy0ZJwWJKFA1dzI9o1pOLtSY
GJZQPjj2P6qrFYaWKFYbVgQCw9N7/eGmtChKR81XGWGe83QPL0gPAZ1alhZgQbGbxqf/+v/+WzMH
GnYeHTGLMoJYeK+pZowXQ0gy3oDj+IEfrk8ziT1+rf2MabPhhHjRx13ixqaW6ldoBF/uScYh2BFH
yLy+wgvCjSZ4HqXrGfmO5VVmH1+DyuvOtccX5fSt6l/T4KUWPU31gu8HsXVD1AG0jQvOdtVfqtyf
qhphiNhKyFYddooXuUVNVnd98MvdChxE97/4ZQv111uWBIb20FhDMFuNUVGRkGZmbyFyE6ZTXR/H
2pxdxCh6xxG4b0qlmbSqZZ1lOFFF/9MyDEnY0Ywt7rJIvmmjNwgriIY8SgIJIGsrj7JBc0W05g+c
DtA6XiUuXVqTW/5hhF0cI0TBu8VMruzivo3Nz5IVk6A39LW1Lmr7mKB2Cy47yYYI7Nv/ojFSvYdl
lX39JPAP7zyn3na81XjOEMJGR2poqZnyVy9MwKYifmkgMtldSnAXUHMNKSiiSNXtd9A8N52EKotl
2bKtjpOQj8g1YLV+Gs39nF+9Nfai3hWgQVjwqs+pxzYu7dP5RChVE+ZS2LZaUgKr9gu3tyJIBGBl
Ffj5VTbtubEsAmGkBaBY/XbPbqu+DYYEEn4EvKaantBDQtDiXb0jM9RftAMld9rgj7kAd5My5231
2QHPHQlMhtvAK4PLDESyyeCo92XGsmUS0IY2d8zINHjh/V3PxZMkbfQpmHzNvnECfqdmvvLKslaP
v2hXeAd8L1ECCYuEBX4w4kx+kYSPJqNbISxcbCTL3s09KZ25dsQ7SfxeDIYCzLoYJUiS0xg77L+m
CBq0Py/qiluLYHYC/mIHOzp471DmPBSXEBRYuBr7gfNonJ+rO/wRjYv5vEgUkzqoVuA3RGbBOHvq
wvq/3jFQc5KnhkLrj4avbHEaDde6lJS/y7/TNeygTv8h4PUd8jPtiCKdIq9jcFsogEVUlt7hWc89
IPa4NQ8tPwzmKzEvSl+kqPjuZCuuYuHibYIP1wwsACKCcBRt2N88n6g7tVK9/xqq3xUDK0tkOucl
nuV0StsRqhNDwCopAw5t5nYrfSIExiKBdVszV0MmxafDvTDSaxZjthNSKmh10f4dYOOVkHpLH5Er
BMgUpSM3wf1pa3fi+Ql8VRIMOc+6M6Q4OD9mbzTD4UOPjgMD5O1Z6MY2VdCrOy9rt9pTqCEmwqe/
YOrUKMGkZVMvpnWPOJ0C8EX0rMi5i/g+3+Yr9aceyxe4zaR+kbTodp3omDS2ZTCXHCFHJNeKDz2q
3vagfWn8h4tLNDVdVEOQsy/QChgXyHqg0uzI9/Mr4R3vUmUx1wLoQ36IphaFlpeEn/C2Mx1m7cXq
p3nmxcjNvcm0GAR4hSU+diMTMTuiKVvEp589h1hD7ElZ6lVYa1g58uzRvehTFU4LXFdNqlzmdDMk
RtNHB1SCM+bEuCdEWWITmqKOaTk9MKv9KaJFaW0PF2JmloRwrA/hRP26v5DmiEAT1DCUhpP6R2TT
qkwiVCr8r6nBoV4s+M1WDSmf5BfXi9UqiOWfjIdV+sddVnqM1tFIcLLqum4fmIOZtXNdH/Wo6Ae/
0HJOhwOYu7gtx4KPtHphp0HrqTDrG7ZhD9Jh3EUjNG6wvbptEecDZZWCdwkTT8RcW5XHsMnuh3R4
eTG7Ko3iCFoErhxRiQClzrSRiIDrl4ZSSvQGqY7KW8ZxA7cDwEzZFCJU6CpgBKp/Aay37+jsQqp9
D520FPutMyQBaMxx47TiVrFmFrnrO8vTc73LMsfSKBIL3jV1X1T5uQ+FTlnNDFcErUaUd+L8FwVY
SRKPPbB/g+2In+3IVaeqpt5tyXGvNwcYHVs8qIjotNwZAfdMPDkoZcrbVQqDhA1La5XDD/gXT9A2
Zs9MOgGlPr+RwBptiRdWwJ1ICMdsCFI1kV+SBIoyEe0MYHeAmNAvpT1Hp2c0Zz3rMfww0IOSUnqR
4iyRMJbjdmv53OdJJa7d1mSWWSm3kjd8B8hIPFCCaFi7ShTiBx/te3nLzs4EXDcTDH3vtow/wGzc
IsIVljg5oGjqGq0AvDV08Fn4AtBGfQs7rpCWyZgojVEueUCAWrF/KAkjQ2oi592fENkR+MUr46qZ
VqKuHjj4TRp1Fm8Ghkvzog++cCxEYz7nK8LVNepWPoX/9kIXywZdDUPDFy/nYZaIchonVaK833dL
sDwNG3QS5Ud5L3TFSRijQswGGPKgNka1tRFFBYiOlXQo3kx7A4koo5s17tJ4p6Ljc7PTdizhRuVG
+jW2vPEEyagy0sEstWXUO47O8OnwbFIrysdZbuFs3ME4m17uG59LIRiIOcEcII+++VJToZtlEj/D
IYqYjvvpuqMK0ifXUeKwZnmfU00isUZxLrDOB7H084m/91aH9ytBxfxqrglU0sq73YDMiXrS08JE
432R7uYUH3LPYHJcZ8u1In8IG02JYesfXJVxDHBkxus/1ylLIPSrdV7o8sY+djCjbTmqmoMxBXIc
T6yMHyHcGyoomBBfirHiIDmJwE8V/TiFU6+Ntt0JOAhdsWZBUVjfXeUdeet+W0qZ/w1kAY/UaxGF
6kwbosJjGy8xh/YXLhKLFq175LjhP6DKOBpm23Sg0fueXWEjXklT+AgVRWaf+gpYTez1SzmeiryZ
4EMiMG3Dlj1Ny27CXg9PI1dtct0Mv+xQidCSWzvup5yOFTNBUawETDX7WT1saNJkNo41cYe1vlKN
9ofavUciAWxnnN5VgACHfuY5jy8IW9GfgUzuK2nNtSG9UNPsx6+puwS8jactsSevRDRn8m5Y+isu
cwCKlzfCxDzg/W+sA4R0CW9CjzJzbbzOKsro3yo4dFc5yOhZPcZyBweMfbNb10oDuq7lmZO8tQ3y
XFtCh1SOm0yx8ZNPBnEQ+DRdifMaw7qcb2BSMLAkpOzRf3u3UMNCqsbWeQr6++P2En31UQjjSGBE
YDy0UBTIoVFRsoNDe1cxm+SVg5dEBgjGzXqcL/OuFWzgOjOOxIy9zndJK4UdTeT7kE7uoNB8TIjs
rhdxexV2EA0yeT01dsWfTi3s5wz4FQS6/Sx2pFZHWBiZvT+tnRwxPAZlBPfV7ocWehNGvm6gdze0
6GCD9qPG8rEk2vfEPcscaxYBM2L85jZq3lQwM5uvQ94WVCAUzWHQmTewRViXWQ/G2+/0gSYF2Hsi
kGY662Sc5vr9HqJ/ag6rnUJTTC2OAEdjximJk0xVG3DAwx376g2Ez6E1fmoKXYdS64GsdYmUykl1
x7eTub69AGv8+FGAuNBHjK7BIW2A4eXHp6J3KXHHuulKsA8ubbOChOW/kK+m9f/XHg9OEU763rYa
AGNhLmeUi6zdIjkGEVBBdXeLQBe1fXv+MY131iW4j3XrLo1MPluFz5MylcI6qD+v6BUuDPX/mE+9
3X5CKROMIfBIV8kuAwM7iOOYv6kPC7hbq27xK3oL3QBatpw5ADt8UCVrFbCloP1eqlZA/LUAHSJP
XKFfhmvnpMK3fS/3zF2tUNh9TbRbnStY2bwuCpChIf4n2ZcUFm0YLuYxy68OrI7Ld00KpOcdFgHE
gzgg6duZl0IAZLlGekaxC8/ynI8KZmnIdwrGY/h/yU8NP6GjZDY9eXUVyDc5ZXe3a1p/OAlnvJOu
OY4s5I96WZSqKBLW6WBdcoZF//R2u5ak35X4YU1smBkroGAWo1vVJyP6aoqbAhcVkbuxH1T668BV
ibhsx3c1xNO8VTDALK8fYudPILOPknj3f8bELwq6gN6pQ5mV+VhYnetieSauXU2MOxjvuGmO8gPi
/yA9jFyE5O+oUA9dta84Jmbc7kTPMVevajjgOrhjf6tPA9BGFz/wdtppLGokIFBDDXYVSd9vs1k9
oZzE4N8RBv3CAz7TpKFRshfMMFa9trGIjhv+WKCTTiA8qlKJDnYKhl4zVxqs4lTC7drjjfaOmrFY
HzBh1XHKyKOyThXOC8KBMd9Bb1QbF6w4dOpmLybkfAr/gPh1BmMrAttpf1WOi7AtIBpf5OurGHDs
FlIW3ryiAX+Ib5zNUJ06YlqgUC5TF7sVYe7DvWpjhoOEqw4VZwsmpjJKMbB4TwAY2SBffJNoQTAU
EHGSRdmTnkNOQ6e0ydkbviLkzVwYHJZpGzmeEC8egeqxTKIjsrcF410QjvOWd7g/3SQOFWYngNGp
0aF8WACHmX1Z9G9Xh28LoBRZEk18fN/2VswH0DTcBMvRwLNSLU6auFs+d4isjHSDCG3HgaBi2ki6
V5/d/9cisJCksZi5u3o61EHCGEyhmTQSK6x9+fTO1N908K3bQLYXC0/Axaj8XW7iLEvLrCjajU4v
VRdaiDMX0gdHvgEvYB9y5oJY4I7QTpJ9/04snkMnQf0wggzLVVMppZmUxpXjguTwd7ypNgGot8fJ
O6NDhNN8By04bsOUdMGC0qyPnSytyaSJgfM6to1WjVGMy9k8VxeBi1JEAjJuGHT2Vch2Q/nYvnCk
Uw8DcoIsZCditifOZu1JYQx5+UbZXyIqW54mKiQEnKnEI9kum9UcU7GrPAllsZKr0r4TJ8RKhweQ
jPwnfgm8mRPynf/eo2FlvcsmIXCiC/sU6bYDx1Dv1SLWCoMWqJUKXa/MigV/VqXFc9qipdG/CmMR
D7ivbXUoqqLJPIkWvctCAOxGi+Xwec8OnVaiFcCgMO255SLbkgs/j/1GhNj+beBKMQ/5GIpnp9+c
NORL5DANF+cmiDZLmz3txfk9114uMh1TB9WtChP65Gs5i0yRCfNBYKgrolpWCRZhLnNAWAclwSJr
9W34Nrj3SpnV5TzLSsi1igx3Xm87H5oaAutMN539qzjuB7RCqzxEOoOpI37bgrHnv3GUorMpuTeE
+d+lJkNYNcDGA1pRVKzuXMZ8CPDuxF0aSZOIu0qf51nIIlrVFl8Z+tF5DDjHsRBXHdGsx0jjdcOI
0S8dom1dlZBInecMoDvca1xDIY/p2swg4UY/97uCshXAbOJ8AcmB4oG/6pGrCYzPT0pm5Wru9Rjx
AppohLmcjfZ1MnuOYL2AV2zbPq0s4AVTTJind51LXgR1pJBsRnJlwxkJTr4MHYjlm8Q7Cl1kjIAP
xk9OwoktR0LrqAX+tPM4Avo0Vno84j4R8F807ERW6LJfLUTL3FOzfpe7oSz2xzm4YsRIxgZDX1Jr
nDOdVssiASJk/mzYPTE978C4+sNkiXg1mLhhbLVkTmcQmOINPCbZYsUA88ihd6+VrH2IoBnG27We
uHfqnBFGqw/10AkCWX56r7rBygnY2HBpE988j7PmZH+epLgc26IncBIAiBOczzqwb+Zb8YRGexN1
XXmXv2JbZuXwB9n9rNIT118beysqgxf6tuhcn6LWJoFSgk2i7swi6XEhW3Q8ek3R5i6MiZwLZyWs
+CgWGZ5GnZ8uvsZa2RhLb8OGrpUN6NCJWOJJhSyThUEvO/8w1yGV1e11beFA+nVi9oZtCxY8IyKJ
OeJsPyU6GuOTUqs7GwAP854tkDB2u59CGfbUZBnNILcl9JeIzj+1ydlwVHIX+VwgbF/e0ZzvmyfZ
a2C4oRX6bkYsI6APqunvzdOqWkarWEVptkraGjNJuY8349C6fqWq1ebSkNQTRjwdBg53HKUDxK1K
3Ijut3h60fWFOAiO9CrGCDrAuR7K6NpjdhsPq9MlaQUBEYoxf5L+6xYMP5+oS/akZJlNugW37vdP
2bdK5ZUwxiqzIbEosKIwkcVzNSC+iCVyb9TuuQS8V1MHcseV8mmwFmc/J8gyHr2NfuT5kLTNQ26/
JAT35EjkjMpAzM71njWhMejZZ/nK6R7NvcpdikfoXse+Op/HRHVOhBBF4kdOLubwXKPf72/xEDoL
lilZQzEybYGn6s1ea2Nwutmup7a4rpcjjClZfsKqEGGY2CwzYa668dr7bCO/7xriMw+rzOUhDnMo
pPCskg4ijx2CIzsKFRPAgdepegexEE5fC6rkS4mKtWofHDe9Z9rjTZK/WYI6yj4i5j++Ymu2Q+Hl
oY7pVwwlzqr+8WrTcAiNQopWjK6k+XoyTuxYN1TSLScElUt1rUyJAGeNOTpaLCHoRi1cJj/BlipF
DeC/lcFmCC/kArcYKhbymY99dPSvgyWbMkeObU7Nr4jbt11SP43+PALkkGkfyuoAFtUgNJVmZJ/Y
NmYXHW0h4vOimOLPZkyFuz+c/oOUNot8XpKpKsGUlGoF0GJ+t3ITOfC7ayXH+w/+p4fNbonsXi7W
box0TKDfZmu5y3FhVXrrcQbUYj0lYHhBzExoyRkxZqY4U6py8zMtSe2roiULoxrj1TresCyORZMm
LIWz9aKR+ngwbqbYdyOryRLsaaNsnjP4Ay7choiL8mQ1KsNfoWDDKo0b+UYYzYDef61OSH8+Aup1
nECcKLIY72CtjE1+jAFCqIo9ZNeM7Q1uQM1EVXVuV9d3d5d0rlRrxXl+Uozta8WUU5r4vFTU1joB
XsonZP4CqhiUrwX9l/mUBT2dQ0VbV+TaZs5ar8j2Z1dJAxwv2BwFEiTzW2dGJrzoTTu5rxbWquiz
ZfvI4le82lEGe+y64MMvaEGajqq9SxcPJn4hWpFt33xzy/DVoaQ5pZhrp3e2ZTeAzRzJQXbZ0U1q
pdeN9HhLI8j5d5eQUesNDPn3N2YRdRcoyX+r5EG20UrHOWuUTzdjdpW2z/KQpdBms1C753CGHDrW
rIqxeVNVaZLzXwnbpl4teUx57PPI7jNJlnIPi8dhJdFkBRxl1oTA+Si3b7e8D4p8iGRgXhYOW9Zs
RIhxhsr7BSLzX8J8HSKm6tMHb8eMC6HGHw6aFZpA1lG+FuD3XYQS2mxmoWyDbaVS63YXTZQ3k87s
8xEVgyamGVfRiw0FJydwR0iqiugme/GoLc7w5IH6QVyP3SJXe4s+CQMO0E1OfrlhOGuBFakl9Nh0
j+OWdkx9UcEqERQSY67mpce3lxVQWE0kEHOkntilHStVA/gmskx3UuLX12cFKTw9YtwPvj0SGGa+
urwCXbCFBwtjjhj221C7Kb3BeMgMSRyHyTRdX94v1+yMSxAhdbN2Dx3KMrZ9AtB9X7m27NWrTYY0
SpiPaKMQUrmFvXG6N/gkDZlqVNag2Y7UhkWZ2Mj2NAt9oXaFs1uCAPAeBsBpxJOlQ0J0PJgneB1e
AtUjJMQ8dAnJoeo2YyGafHy1M5e9vkOQaHz4VD3jA8jg06qpPRtOiwuV4YmA01D48vogW8ytpolJ
laNT278b/SZYiDYQY3SISHzZ7lw8nLZXNoK1tCoPD4JXM7UlFjNkL+S1pRNuMX7RdHFIABV7XZNv
XMHXjFm3ayAeie1UrWxww8nKsLhwt7u+BlwG0ZFsCgMljzQtFu1Ivd0ljQQDQrLJMvebGnHLxyMp
DAZ/qMXv2gN8R1YNK+XRHP8wmdLFh/qI30VT094AdKDdL/jeMx2wKb0KoeczqOGPCTnxwbJUCwW4
PzzioJZph+Gv5r8xOntnRiXJerPNBaGBuFK46vPLBCkk86+27pVOjmty9l6LiPXcR2xX8uVDgRF2
5x/2KDJ6q878xX2F8qXn+ipdhgmgCsKvGRe9kIqjQBVz2q+vpzEpEe9OF/uBTu1qZbPN8l8mkmY0
LifkuDXj3cMcs7TLN/HFIMrsIDopNpSYlHpUOMP7KDikaBj+5wgmOHWg7fAxXCd5J1997+7NKT4c
4yVs7z0zYThcEmdyuN5UaqWeNxOqaVn/kauNVkPxfh4j8xwyPU9cnqbOVsLdNSPSp9pr3E9auNNV
riY4fRwHq657rFAH/VpXxoSqIpoyfcRUOGdlPXPJfPahsMF6H/9k1zzidmJ49GpOJUNNSfGzTh36
IajeDBpkbeBDCQSJzRK+AuEIk+S2r47oOL76dRTJXsjNVla1BRcPU8NkP6owKHVsYoqrfME0/Vfp
du4KCZ5d1gHS1hTPxA0n6i3N6WYvTadC/aRkNd5Gxl3fexq8xmVKSGXd9K+vtjl6XDep7p3t6Aa/
UzV09OW1yJ+IatuZIZ41ilnRzhcrD+AsRQywnIWmJ/w67K3QHY4XekhJxN4SssDdmG4jvqVQbvGi
745CEmZd72neihgS9Wb89TyRMzakf9m8r3/HyIdRa9DypTINrZAKWwBWEEn+HhiQxk5WkYsp0LO6
/r34tLN/2gMWFoBl/wb0FCvZDrdEM/3Lpij4B6g9yX3JJyZfV8MGeryjEECkADa7hTfvpSub8+vH
q/mGugnyj4IIQSuBZUipJ5FuLIdaufrAZTAN3a7BXyCy/GsjhHzxUVepqsh2rAq1BZAoc4ilryJ1
e+EjmoQQ2pGT5eiUbCPR5lFAFJ0geJp3liJ+r26BgFmPLi0r4YE48f5dgpe3N4ACxDwIMNtWNLMV
4Fr4XuTn2RQU6J2iPGgBKgDKzcHMwCwX8RrsE62mnnLMV279W9A+dZ+i4XSzUrVXyOipP9l/SRCV
yxnv4uENHJev4p4uOE1bURVPd9ITANS/6Ve+vqQT4BUC0B+FX/TzG5el2zTgNbXgpVJ4zU/f/IRe
WBwx3ZmVOCzHT6VnMM5T9RpnmTAwwDSsXaJICewpmLtjspLPzL76gledadeGozbqJggUzdNxPv4A
Imz7ES4+1G8LxstdOgCHGzlclTU/NLOROujx1MGSlFjL9qN2TZ8j/iL/Jr5T0cRfKwlbSTO76QDK
/b/zh97eAprdxgRg8dTutUalzQhXXdAI7Oyp2DFQgkaXVfVYdwccmlzZ/tanktug0vqsC51JkdL9
CsmEsp+Cg6yA+qxut/uo+SL0c69pRkBSmp1T2zm/KCJdI0AVKNZFVPDnO/mWgYTXlxC2/o7r4xL2
0zNMjegWrN/RY3zAF//mUC8VxvWTgLViDwoAwQM9SolYvIuLSl4iulXxXWwEWi3wDHRubjvf1+pY
6q5Skz4EMx2F/EwO8qfElnXpPyWP7OstSYfT9Ck+oVDPGVpxr7+UDuU+lCxT9kt/SetUeOdzBH/1
pmnmFdtccNi9CDtWVfSfiXL5sBx8z1r87S1jUKS50NzL3dQckOeGQbEg0EKl78FOUq87t6XXKy00
t2uxgbj1Dq1fWjBHqtHTGI916kWX9PIzes2oEbcyAKPWEFoNLy+0kcKEP3+DOItxVTzU+i5QwRBQ
yZBpjovHUCsXFE+gVSJ/oA/xKHSnsj6kqu5+jM6G4X5O/9bnQ/cscKJZBwEFx/KIyqe8oUbVqonr
6FekX1VXAFrhp4yv3B7M5c7udpT17dAGZtGy3ekCDdWOcFPkQ/YA773hAZINOJ+6vrDMKw3nywOk
+A46E9bRkzPzx5Za4XtN6xAVZpCquWp/uh+0wt/TAZvSMiOQPrz26uz2UDI8OZS7LdPmBVfk633m
lr6EhuQgq+01naWHLSNMRcYK+QT+sBI+JtlNyqZ51mBHujkkm3vvNCZp40LyFQfyTHs1Ttmxr3UQ
N6alFTrai+FfKdNsfG4Q5fjZiqNxke+0mX5c1RwJBMVyXvsleXDowm2OEkWY1I9zGfDww8PQu5I7
zdFewktSdsJZHhHqVhsAmsciEocwxwLqIXO88QJAQlgtKmWDNdK89yURk8X8MyVHzFVDxu2mMs6O
mZ7vkzVzS2Gpg59el9ltPh/sDUgZahwI77LEJ3yHMVtETVtZk4mB1Epw3CR2EPscxk2ZNgfzJv+y
k2x4fQ29wA9FZiiDPqlu7nDmnbbkOHwbcjw1P7vGyWQJWOr8pIz+/cJ0En/MrrktLEV7/RTLkNQl
+nupTC/xI5WmypTMt1CyDLE4wRz4ctRVfMMhcXIUN8oir3zgiXY2UhyWzLxp+EHdiwihdIXq/EgE
dhufnWq3SRuAKoDbxU4cWg1k4qmVWi58h1LWhEQg/LbIL+j29r7TH7SaLpruFrk1JDBZ7bwSK6UL
md8CR6Jrdrl+pjjf5Zt7yzZqQCe0mV6RQjwOZr+z8Zni0kHuMw3vr8Dn7Mcji3Kp6YnwWNSt2mPT
Jk/Ht6BOjxqEZNBPoOM5lyGidkbc/2NlOrUS4hu8YztbOWLD/6lLAmmp2QFHMYHw5yMfzz4Vw6vN
lER3uQwE1++a/ocLaq0l0/3rF7acG0B9CZBzLRKRE21ybnUNEPTt3hk79kDS9iABnoXv5e+8x/or
iBGGXFcJ3LjDNcQcmoklONioEyCnCHSZr3A8Pvu8lbZsXcJNYSynUg6GJiX/C2q9KeujJqaRqRfz
x6Zn+gIXGU2DO2diETwxGoldgTKgFtbXxP1GwTKyW6sQnn+0K91GaxBjCMSG5jwLxJQBCgbZBcyd
jUON24MVNumy3+FBjiXvgTXaFYYdTK87Hqh+ILPygHpFIukcsT3mjNp8DiZts9iUMxzrHO6ny8XG
WtySAlbJ+teUW/+D0EYBSz6pl56qXLaWAHCUa0YuupS3M+mYG3tPmfAGBcX6U/RaIC5bStHskPkR
6ZPNXTrCgjZ5nQyrqlKyAsFjRuFBWfk/lpOEZgsb69zajAbLclQa8ZMtZcKKZtnXSnU3r4xQhJ4w
ST1VX++qo2Mb5OKofW+hHMMlWz1l990XZbX9CA4QJ5NT/y1VZk47jIpzWebTQr5I/XLmxk0lzybr
nERDa3WE+Mm2OJxZEzWbX5BXihXNXdC976Zm5NOqFdJI/BOBFdjAiNZ5tWmSjO2XMZq9lHMVRX1y
mun2st62BpJTBUPSF16jjb7JWbM6mxItQHVYLC7VcmSrutCjFX5NrHokLzLJBDVhSsZOyPnWXdNK
N44DExzGgJ10GtFUGRjbzxyC+r4VyUJGXagzyeGKAUaIaZmVJXJ3jOIbYoA7BnLSzQd9AReY3EK1
j0bCDoyTozkSRmr0m6GYgVHfduE/MEZUn57VN2qLlcRvv3GXsF4gKduYzWHgxpOFYNGVJEiMQidE
tg5aMQMMR3zas2BdYs4Mk0pqX/EN5Gq4DZul+dOVxc5AkyYAqNBtKMQ3OHFHZvKg3FBa3509dWZS
l6Ah7dJDAz0Y7KGJFDj2uWpCLLFuc72UP7QcrjdYrDlJCKYTdU4z4OiNk0V7Y2WT1AUi5OCNLC8q
kU8Dzwu/i+Ch9Tb5/ahPBv5G5sVwH2Br8GbZteJT+oxDYDZOVLIxRKqAeudwhKi48QanZpCfVedx
BCT8cTXP8LbS7NUbG0Y0vJ4E8Hg6cFH+qzTZFP7Nc99S5RIsYpBhMgcm1tmasIxKcspCbl1Z8fRH
bAV2leLBCFwZdGG4Tz59lu3se1cuXtBwyyAvIzJKswvO6/K2XIHGWSpYwXCG+0ClxwgqKmZVjL0W
9d2AnY/YAhIeiZqBs+LavwuFwJ3AVF1KQlJZwxIqXd4SZidGjWDApgPThKTJhvlk917zbHgR05yV
m6rWYJo8uWDIXZHyrHFLryTNCiq3X0PB0ryHjU3/erQJzJfuYvHvCUG0L6EkZIIw4uj4i8Qq7rrV
PTXeD8027er8AmnN9kLEx4QXex2UOAvjM4os+cHxQX21fZ6VN6QkEov7pVztHt71Yi/v6cKWvL8g
gM+RP9tz1uRVuiQqvL3gAhwMPrLwxrwFZBv2JZ8rmLISjQoul3OFg8s9noLImKFTdSAuYX70g6uj
2OvQSty4keL8sWN+rpI06xK9j+OtWMoggcilOuAmT2E1SEqY6h86GJ81VQOyuFV1ZynbasxxeKJw
FLnnCIos63JjPCJKZaIhm6c26MXEnqnp8e2ocAXvysz9hWJ8uHezL3EJqwMGeJvQOe7n55j/a8t4
g529bZgg4og4xvl50cfHVItA++rGceubKjf7+Fuc+f09tT+9jreWGPbDAOKkDXfBcIMXCfJ5nyOB
IrvMhf9507zw1mcb5D6bRTHB7S+dtLOz5wuCcPmJGQvRbzjQoK+aDJeaEGDi15JY0RsQtLtV7FkG
5Kqti4QPJW9YDqaIXE6YEI4UzonO7N9dUEpJwrnm+ib/jl8Vrx2tHBybdo1fZG9ooDqtxfKRUv5H
48QVC5e1aI/Gee5pGkiyw37kC/ggHMjMgXiyV/asjtJTu36sOjzpSNsvoq+bij86BfVJpA1ZvEOn
W5PTBBWdNzwxSg61MNc6BK/jBPAmurvUR8IknYwI3s/jJhGhIfTdQjkSBun+6oCC/ejCPCNYkxFA
fBg+uz2utm+egLDUxCIpbgKYXe2YCzuf79Jxh9m4kbJ97QmM8QRfcWHSVEUZZMEaDnR4N/TBu+f3
llc7P1c7ksFatfJfENM04IHPv8W7wje8NEgb8QjXZPzMmLvUnQsqwNUADayAnH0QgRBUlI7cikRO
QhmoBxSg8S1pG18IVZGCahBA6hMoOPbecXX/N85L2vP5jqaonpeCla1THwBDEWtGgNg69UyCg5yg
PRCxWc/DNrdRvF+Q+8LwHZOQk1LXINpITqEIGkp+VqtNUI50f9GoNOIcp52Gn33LpBgDMYjhZES3
a5cV+DwCM5B0eVlGoWF2RAhNUELV9za+v1vTT/knXX8EH0ax1TNaqKORfyyRCCiGXggpc0vKq4zM
atqeongkpygbz6s0GDfYUFIS1bMs1G1VwsXEjHJRGa8Keumz/Y4DViBUesNmTFndL1/ST/yGvjLI
DidXR+6tg9DQnKHM8aINvLAxlnHRMRtFF71AHfIDE/Q3zDkWacEX46YeDYoF98zTc2L6QK89f7Rh
lvTrZcWt2VHLDB++TpAe3nxSGAeIxgB5iymT2pnHYQBxkTysBfKZQyiqjsKEXcvBr+I/C/mWpf1d
v/cmu/N78xUBhVyFv4go4hfIgpTMSIcM8AfP6GPTTBxE9zT8yXi0jRchBnK6Hbkf6ZiUiU447y1Y
b/67OKGhS3b+MbOyGKh/sdsygk0OMB9YJHlo0vQ02o9iLEYiErffe72HaQJQAn6Gf0wlO32HULHG
QDVta3yiQfuqDaK9ixEqtA5Ok7zfprBc83kIJUM9synxjIb5x4c6IYY0M8VTNTOFpXylFPcyNjIO
O4KJizTcUGrc00/Qjxmbvqxcch3gmMMLetuqqySTfRpGFPEE0p52g8GWi1fCJYWlhSAywfJ010jl
jiZjS7Nn9AM+uJsiaf0xZHIO6DoyHAN+nFh9zCl9ZYKrCUCZPP3TyiUxYbnAiOILUkZA5LLaEKGa
WlU9ZtwiPjZObb8WNQoiiEeK/hDAuXIs1SBtez1aK+q60lQSkeraHKAPn7FXzJZV3azXID4CdTN+
8GaE5yX0F91Svjs1nFp+cjSvAl2eWCi3oyIkq1PPeY8g/kKi40ZLjNXR12ttQT/AqJUkPX0qy2PQ
pMyphOtRCqj+Edfer2VpDQUJ+8TOIyHe9/wAlOKW01GkrlOFnVDejfgn80wk2tM4F39mnYAqHNyt
30AvnatzU4UJnBwH4h/clDHVw2dnl0050ckRsZyFy0tkP7ijNsS/wjGQTjzbE/n8y7Ql1xr9bgN8
3a6mO1PqhjODcM0IfILu3TSDyLS+NeGdERmNc6wsudyVoj3pvgA9xPWlFFtAQuA8/NKCmqjOVK/9
2VVaXGbWtSKw6qjbZy/1Jbjn8BicfqJpf36e93rQBvww5quJxDftnQbm1KVHeKlIOC1HOWfDEAnB
nigIA9YLHmfUJwU8tQNXKHQ34CN9+k48we2JU/01Tu1ZmuwPrQm7PDSBtDPS2jjrWXtB6CRhEkyc
EycyNuGjvmydFwIz6maVPZcpOoDHdGLfa7PcavjJI589hqcOR/QzVMD2uns1S8BxSN6tuTHjvCCx
jNo1XtfklYs8ypI7mZB0gpDis8Ez7pOmxdevYVY9FpH0erk0hacm8lkDK45gGSq4106+en8qmCmo
kfsfIz+xhx67FUnORxZ3IuddhBbeFpZJ0IHQHcIMKZ+iMeTMwaaKfq8Tx1Uig6jb4UJsnpml/xRz
OUC69ji83QKh/tPeXHUUpzDh1KBXpW+aq5UIyfRL0flicz6fOEvXI+9jWaPuQZUYz68hojCiG+/L
j5iSTGxUcaCRoU7BI6axi18o12W3idO3UFaY3YljPIj4qILTlTg8lmtkM8y469vHoQMIy5RqpZzL
f2vQ07UtFvMM6HCH0GqJPPTbMAj4TFoE36T3CvHvTXf69+juR7M7TwjgSwziXZZe3Is0Rk5ZMTUP
5g93C+SHrunRW444oJxv9LSAXCmcbarSxKqOP9LqLbtHgkDImmOaOiquom+1wPFcpXvfWalvl8jH
ktgUUqbu0kFLQk/K7uh/LoL4cxi5CHC6h1KGH4T3o0hy+dj0aAF7v5Cq5WrM4bVlmU3kSCqo9bGS
mGU1A5Bv4GfYSizBaDCXzTl2LmFNbRjltOCm7ELD98MMqdFKT5sox6Jiq8rrouemlFifqBZJjwBK
EWl2EbhblMRkb0krXAencdCp4AvWL5c4YGddnjBuOEuyEsfGDdqrgjjDfruT/yonKEMCmFC6/5LY
hDULDvBNyu50HjGLv1L5ytO8TMlKJnKUzK8CRAx5/PTL3Mrq9tD3V0FUrtskumIhS/b8X/HI3FRU
1ZtDNIem3aqWwt+l4eCTOwPazUY38E3m/kMxzez7IE0SjkLayMT0P4vjAoJg8kswpm8ZKYcVoA4C
/kwSYA4Leos29I+jgKHI98MDZslprw98tsYcdfGdITsBhp5p0Kr8XkpQY+XqhB9LmKHvkGMSl8bo
0eSGK1M7Q9rjZNOjuFmYpxdLwKpaSbcldgZTyupNgQ7qjO0mzenKWCR95ZaD4JQEf/9fhjW6Fkw4
+K2oL0th4JNiTV77SAvpUH4AaZlj/Ix58/fIqpPPZBznzZ8HswJTMwTRPM4aVhtjhiCN7WH26kox
sTcurEm2p3eJGUz2sntM90hA1bdEBw5jpy8LF6Wn+GRCMITF3xIYSBAbODtpnViO0N1Uyf7vxFcK
QKTtCvlqlZ4bqsP2ohUrUkx/SRyWvQi/RVU5o/XA6CVwPmdwBQkorG6X1ilLfOfPsxg8ejVLA9F1
mQWBXrdsH1VNNzKEsYfPrD7O7HhVBYaM9jfZWWJm7WuitLH/jiPy8IkfayXFI3+LE/qlQLZHrzBP
tC62rNcs9TVtSiFrUutntIOcbwM1Rg2zlA8CTZJgmcMwH77PZHBIWkh5WvPMbmbXB1NcngeBR9Pg
Qq3SDwubceDghtOncPs+KJ55G3smquxNeb2HkWzPH02xk96tnA2fdzpzRyOzDPGMwotfThloC692
sPeUjzqOhbTeuKFjdLnZGkRx3rXnTGOS658S4X8GGw/X7NbYLznmLtZjObV8SejMXuiSrmqxgiD5
mv0wQGfq0a2XjJ+gttHi1CEBNJYGqAShFgkljKKYzPzpMu8NEUq0rwfybYzKGl78NDZLsAnvqqYQ
O0LVan7tZEykilE667U15ZO959RJPidn/iqrOT03qrnJYEZFsE6WWw/0EdQUn937DQJAJqLickgV
p3S68KR2UR1Le46uIINqpGPgfYuT3DeLq0ySMrD+xqKUN9SNgjwPYqmJ1Bhfg9Bf8zRJNXEmA4Wd
tIUJIyDx+ZF7oVCaaslWxN8sxVzyP8JcSX43GDCRa9N4CT8LQwWmKfW3i9cXBnPVZXS7nPtcSgRX
w/S606btEXIdv3KCS1lJEtGvFAoN79gxJSi/L1Gga9puvLJDn8U48pHqAYcQ754jF3WwKx/J9qvn
2hDDG0f4KpHL3zx4fl2iZODj50z1DoT1aOEONRTIbNcRAZ2btoRc2o19VqiyqN7SOnhjufGar3oc
+g5CQAN3A+i6NOXV4MwbEnJuyLUy7UmG1z/9eAdD+gXaSXZMkYVYcN0Or//La+ga4Epci3nrpoeb
bB/HthIVBiyoLPfA7gP9W7pzopjh7FGv2SVKCM1AciNv5WA/pPTOiUN4yZCV3KLGtMelU+uVj7LP
9Juef6f9VfM/61XSSwXNdkN5HFnTXKMF0fBPs7538r4F1kpAFchwPlCUonDeGpw2kwMdtVS/KaGI
TRQ6BVv0els2GNQh61S4uMRbNFOOHO+d7VE8AirbWslqQyFyiDY57+8tcG6bjXr88NDz8DE/ep21
fbaefcAjVHPiWDk/ngWAG/OhNq8APd2cNlanrWYOF3V2bLfNZWMsg28fBwf13lavSOSleQF6GOih
4XTcpLhzRLXnMYsaLUM3IfiagtESH2E3mE1hT/+FSU4sjAkA9mxHFVXejWByJAanUUrm26x4DBik
2N+/hkHgrox80uPFefoF1x88ePGfFAjVUb1c3U/YH27ox23vkf9+nUUgG3EodBES81MDjE0rp490
H/r81Gj9ZINJhNO1ED0FujOL5tQ2MFUk30uFw1LsoIn93x8FjCK80cLySnlc7Iw8IPEJukyrEDGL
tAoA9c24axD0gMG+hG101QOuDT+MrvOhKl4R//nIZCrmCceZBBE5mWV8zkDGWoFBM0ds6x47SzOx
D4ob70L06vQ6BYsfr53Rod7fSWecRjXerblHOCoC20qG+KmQDc8wa/9Qs3SioDVxw8WEgleFscAp
A/GJ0w4llr87fiID1ZFF3lB1Jfd7Tt78poG9wXZW4Gf1G7CXuvZZfgnVF+I+SLWWCuUBbHIFpNJD
9XOMOzWvYrOB2EYQYstzMvQiNlxZ53bX9LRAWkWyZ4y2ncFzQ7haichZJ/OHDmFIqFUkANK8JTqe
Y5cZdznMyLno4G4nBKtRJnHMSxiiLFvcNqzeKNA7zHIxPWWCUn1+5roki2sYQHu6kSYDHBEcVryM
clP+p1Juu80JOpu3pX9R1awK77evJVNujD2y+usoHSGLqeKvC7O5fT8Sex5PttKran7sh18qCUQg
2m5TaDi/xnrL8DsVdHBEFWFyBMgRS1lObGJqama779I8pjFTyl+D7zuTf2zmBOIgKjESARLn1zbN
wkso47HgUNiJDWmkhJBOeVMns5PAeot3wG13A5X3eyPgWPNI2BRyKWLlcn080WIMe30b5lVQMP1n
aw50loJ6eXTNhuBr9I28tbGhq6iDjFfBOWjXBTq70DgaQPCMue+UhmUM/SLSiWCKRVzJre29w01Q
GLXM9rvCvWUwtP8hzpa5F1gWSG0V+g67niT8QneF8ZKw9CnRPpgVk06QW+phG7Kc6+LIZATwdAvu
w/PVjyAAsOEC1U53B/mf/3SXM/DKR+CsmGXG/Sfdt8ogBVi9XyUJp4JXCXAYto0Ahhziw14W4lZZ
LOWDvIhxeT/0wU8bN+nK8hRUSgf3OjuXBxGNrQIUkxcEvzT8A4YQ+S5sXxJevJLMVVuLhImY7tUd
RXjIpCGfGpjbUb5khheH/D2lkJz+0OPfp9WeL0h274a2/Z8kRwlo3ljCUJ6SqeS9WbU19jESRdBx
8mvQX0pL3J+d2NDT24TK9i7oD54UNJorshAodWFx4y6lYj647eHVivhEgcWsHIdk3itgqRZsfwz+
JMeSGIVczRM3aMRKA0EMJrDU/QgcPueC0FO3o4rqklgTzSHXHBXh7KUXLhdZn1GpJStp759ukVDq
+SG/NhQ2BmzXWORj/cQJk9RWgn4ePpNV0XeKq+IwBGlw6qZhHcagY2shO7R8AE7iuJ1KK7Qi/Muq
RzURbDzL/kChsDc5GHqfo/CzuX2a46Nf5+zQ2ZfZIWWGekmvfdb3GQezc3T4gTEE7OIx8lzhzfGv
nptruuhzJ5CRYllGWBW9NxnIg4lj8FSGqox3QbpY2oWmks75PgF55P6dqk1lFeWzfSiRWvOou8Lb
MRjLYy3hFRdfQ4kCFcg0C9EXhXC+plbCN1q/Wtr7/GewUDIW4+Ys4PdR8fhWbGU3TBBxtuOm22Ym
BYcBhsD+qujnPAQo8RAFFbyodjXYKvUOd8eRFxTGMO0hfPpvyifl7Ft36SF+Ocr63vQ9/+at+ddP
ghjSmrJACoTqNqfxNRhw9rkl5hnWPZ1UjDwAGwIGDds+j/ZxRLTqs+6dMwFEu1SjYEZTtJxNy3Ob
WQ0sZD2rR3C1gQwgjfeXD9RcJ5asPWeHAABCquixdc8H64h0DE+dBpE1vi0p5SZ3Rmla4fnur51O
dmB9vOpbBtQU3j9YCgeIAbUueK0PR/Wxyi09zLerECtQnYQI1S9jrkQziAkBfwhrIN8MDNHaS6aq
0Knd80f3HzNQMoMLXCUZUD423HvRW7yfOb1vxpal6vvTi2+bLogVnu1CUs6Q2+XAaNs6gYOWLJ70
pYcO9kJOuposZ9GzUl3b4p3QP7FqazFLBvBGu/oJXFBnSblHbt7lIxiKtBU5X2p+7+zqui5Gc2Wd
sRsv1lvRbxjSriQ5PEDBzCTcVvTRjfhLy1M/I2s7Hd+F+yMHEcg+UnWgRb7U/z7P0mDuBF6OIb4N
KOARJQzrPPZABu4CaIkzvm/NSzNU5zB9MJ5I1YQH96RHqLXy5wvjJav1ZLtYZqwwqXral2KKDVsV
PMLEEasAgY5FhuIfYER1nDiAGdmNIbRrsiaJ2j6NayOrepzMsjNfWfiH/LY2vE99L9PSoQxo4Pn0
HYE7dyjQdJ6SXZ9QX/PFsTH/JvlhVmnkJ+VbTqb/TojS+XX6IwVSFk+5KSNyhfLAbifw1+WNccyh
TVzbqLnDEhU8oDpcdh2IykbonPeFfbhELi5QPNvjdFgJLosqsXDRII2WH3lnusAPZ5Tv7Xr6ZMgx
4mmBgkGt4UFCsBKzUbOovWCR/kBysepszpkW+jtshOqz07TQfPzvAyjbUl6yGSsf6YWWDqHbzX3m
Kw/RLoh02kkE5tdltWppMkAhMOoX8triDfrnB/Uz8GRYDdtaWVKLTn/ue7PKXKhRO4RlxamEFFGn
kklQOC250C/dRBBIXoMlUEU2d+bmwBQV/hPpjBOHXZ4WezooCyLDFDhV0j4fKiHwJ/Qqu//MX5ZN
mhEFTrh6dbM41TtmNbXIJ/xq6J9KzK2kJvOBEgu6W7sHlgZjkbQdlhVepdFixQl/4OhMdsrNGyMO
56CDaiWYHY1h6Kp3SqUbgm/zrKtsoexJnPpIug1TQ81nQ5pZHk9aPfXx5KEM3rv8WysrRVHyFrv0
fiaqQnNHYn0M1dhmW+vikOdkq92q2rvMOmuOd639YMUIYgikX4xXEG6n3YODiahZf0JE43haVxRQ
2jxll5s4i+68qBkAn8sNLfYSNBFUlgt8uf1d9s+z6l74INnBBbutUNAdUOak+e9vewfWFfhI7gp0
Z7x+/GMEUBydipNq8pM2sENzRQBZk1rvRT1c51dDydMmJlVR3VBon3XmbHJKX5D8/f+kTVeJ0sTZ
P9veVoGHMb8YzFI5Yxh5Yy4WhS1Hfqi81aok5yzk1DRFaYwCRWIkbNOL51GF8ag1+9eAO3Y5mlB/
MIX5XnbL+5983mdwQql2xnn7t7ak9Nhtyg/YHTP+KaAyiBc7931yxfCMTBF5dhxBfmir+8hR4jF3
fSR2cltFa5yQ8uLysRCRM2HCIsqb5taWj9esf6AZA7/TIBtzi3O6TyU3CnBLLRtv80NGxmoWpJXD
+VZwqmQSG1LZo5Db9R+55SLU3+QxGMJIjPRAg1g2JL3ZE1ryda+Sp8s5/XpDeabKmKd/L5MNWoM3
qKd7RfdbnkAijgGYbNgkuFIMmIh+HjbpjYHY/ESZ1tvvzF94cIOSmYx6EtvqmSnzsvtuN+SUNwfa
FOlL4RzB4fMQ7VYwqKNsmj84JAcvSs6B0//RATQnUT0aZVC4DIJTCWQGvuBYi478Ndm+kuHze8c/
PoMiTu6EJvCS7Ye3ssD7V7FnxZHy+//jv9VsR8cGBXNmAkMACiWK6TN11Fb/nlni5Szimt4Lnvv1
i7/ow+rRo7LCvF2c96SvZyOpMYmPxfMTDXwMaUMI92sUyeW3dKjBIRpnrYSLOXjwsUuWBVAlbjNK
cBnhQAyY3/8/MEICPhPbQpmLpoheZDup3gEjkgm+qq37yvSIPJ0dyO+ihp8UgTrr1Cx3FcFOnMY/
tuPeOtEUPM+nRKOR372zCNoijB9nQHoNAo43RJKoW7FdgVlyFpSQoS8JmKxZ9/j3Mu9qLrDNg0vA
3ZrqwWC9AptuKtb2U3YDefmSzoCYCnTJwqEZUtAJegChHPMI0YttwYsB+RPAUfydj7mefWpHO/He
xf6jMKp56ekMFH9S2NYKZixI9e05y/QckiUeLcrOBXPhvvZull2+XQZKvpJPCNcVJk1LdycKK7vr
aN9JVy1IW5/pLaAr8KdZhocMZ2kSagIbifc0MR+TfY8jZtNGCJYWjx+99OFfgxD8ZFSl/GUXSqqO
1zUuDw1HnRyW0b3LqCK8vy9EpC2vTHEQ10G0GenYG5mWPr1ut2xF1PFOUyTUUhbYuRyr54bmkV7V
inSlTD5WNyMR/LnRyou1YNPAGy+qCGpCvcX14Y4sAgN+r0TZKqYB7rCjPBmy7uZkNewLXMLSLtiC
GyEiBj4I84gZScN6oN2dtkSCQy7p36Zpt2m0jwgu8EBTPvYsY74CR+0HbE30vhsMIQJMUe0eV1xD
8yaWCdJBlMEkCtOiVdGfGZ6tq09jNhKXezikmRyGkAlGysfN/u8Wc23hE5exc4xR1xQ1vRvXR36v
i8pPEqqn170erwOzjJmBk5hN7xLXFVsUoEWLXQGIcm05FtpwT/SPuyzJ1XlnM78Y1zDDdjFYFW2n
baAZO0MBwdnM+gbckNcOOHBP6MsQIYl/qeDl8ic1kNe5o0uKk69Jxw61pqjdjoOpUtSBch+sphpB
u/F0kLoRZA6u4TXH9PhQoUnVkHenjOXpFP1JMtcQYSme4aMB7Cslb+b1otZMikr7Jfvzrvdu9R5A
fWXdJLU5uPYw3Axye9njbhzbWBr+L3rR3CH+sc66Pix0WADuZc8uF2AnpjDY+mINyEFwkqiUgHU1
yCzP3s2FO6DNLkNKdwzRoNdi1Bu5N61X16K/z9nfgoxAMKAVcjaCgR8KjAX34IdHR0z+i+u3yrOS
So2Q/atIwOE4DLCyP92EWLWDUUX7fMjUpArWv2tPCQuDAvsJ0aX6BywEwfaIlobchxqxZG4GK6r3
7OiY7zIkW/pClUDIT3cVvg2Jpgnolu+TxnvexIbNDnGYvx31hrxEiaLA7aZ51ucPxhwNYmHycILN
pdZWXjsBaoJM0p7nvL+VBrOsn2k946BofyPf+OI4eCpS2qlfp/Cvn0QHlPZuUsLNslNgW1AfMA04
zamKrDWJIGbQ0R/NRpUOxRcC1i193PZBs/+omT/X+TfMVlPYRcOUibsocGoXveiGPwXHE4epak+6
+2sKK7j5ZrnPfwBn4K9OccsNXmIxBc4wM/NOJcrJYPKlRsFtT4TH6mzqPK9eQHNCQzg1/XzxSHCn
2meEbvoXwKxJVzmltjTUcXYO09HEDOqTMT0rUaJWqmqxlme0vCBqLmMcskB//IV9kg1gpmVxCA0x
pIXwmJoBHWntbroW9ZJegUioUnWxkM3BqOJWYU8BkZ78GtcN3DKc25qALYJPTSL3QQw6C6RTDSJe
NH7Scmcztoop3KBVMzXF0ERgLNQFOijivQahEWIjlqivl++XvHey+JOgWQYfZ1bFqqRMVyVJnxF5
SNe7eKBvPCIbL8V4+Ckh7sHoIxRZCZC8m4ZvFdG4j2H2JyBOdhv9LNP+Mf1Ku78R504ibavcm1gh
epba4cO8KIi++4bh3352fzaeQAdwSXnzjJFswVQooZx2Zwx9qtoZNH8VtXnNyPMggjG7WaaYZHMu
d0S9ryLWPyxVSWR0NQTY2lhl0g7LXzDO+552DdvIkIM+VXlOlkUOVWoa76FhesWp0HK1c7A5MesJ
rD/SD9kvDMdPObutBufoXQGLVq4RXAdwZGtaHmIE6u9RdeVZjnrFoSWj0Xk623vpTToiqQWBSatr
vwp2WrEUYtWxrwttSlkU/cY6MpUX7G92bP+hXS27/S4PEjYqz6CO0UYu/bcJGMZBmNzkwEZtfMsa
yKE1JVCP5clorjP+Oa96zJHgNoBItpIeCa0QZd+sV33ZlCuGKjyMoSO9skcRvxrbVg48uWQDe4y3
mJEejZbryktnmojN/ArCAEkLaEji8PEotCu2gUBIVMWRLd+1O3gZpSpTjGUJiabXwbPfL36DL/G+
Gvjj/HEnreep+U5j5/bhZEOGBk4TNoaw7FfeuNR6NxKgvPq2/4PSGk4w43vXpVKQJU2CO/HRYBmU
NleubQIGUm1GlbdSjaYodjXdCPf95JjBflqgmwFG07UCufii4VQeszbakYOqfor1E+bkvCyiN6Zh
fSJgLNh6cJzMi3f7ag2S07cQFoNYwlkefAttnwNCPYH0t6F7ENyst89k3dYgn1KnQcU21IHl90Ao
4c6Edg5prhSZ5heep4xfngGVx2aHKI6IvtfhIRDYcpk8O024IHi4bgqAIsGdo2sJENgpjCbYjkoC
tmRNdxdz2p5AxdPKKgaYg30+xoH/Jvbdl+IGUjoGaviuqfOAVd+yABSqTB8umswugYWYEMKDqDyw
8uI7IxJgEDunjTdAkxc0zj6rXi7rxupLsVLco/vkTODQurLJj77Vukv0WQDJbzybifho+B4Mdmjn
shlAZCoLpuWIGX1j/QpFFfg5zaPOD6nkHLSxfgegSEvtbr1ClNNNvwULhW9dnN1DVvn/LKRZ1MXa
WD4zZjs+YKev5ey1nMLo4HQetD/Mp/nggLSSl/TPyhHeg+QTDYRcipV+G5X1zP0d1cP6Y4uGFm9o
fHg6sFP0cyF/U7mc3MjUBmR4YVTQ5q61IwNkxRvLd6TyVNLcAZFiP52V9EAippnZOz6w71zexAj8
AKiGctQbfnmv7VtOxF8JYshYdh1Lftqv48iMVME3ZEb3c8vugPGawwj+jp4dIBo+J2tegbICC9Q7
nBncC36WiSxf9Vl4IBUvL6757JdIxzfrGivaAq1j01AyxEnGou7WSxo+yEv8ZJrnxcvWgCCpdZtI
+kJyOFfi1n813PhuJH7z87UZEyQiibuzf0F05QS6Y+L6Z7LPqZOSHggsviFgvlf9//1aH/3G3LPw
R/qHowrJYAaRTyUyBrGfOlUzer7WYXVBlVsZkshSWNB7AEgH83Mfkr/MQexamjBXEl0HGlvImdWX
/UspTffxjMcC1CB7g+4R124LzlijYFGx0malG6cZi77dJLDDJhXw4cUZxnWRmG9acGYDiASeBSoI
EnGdNIcwn6JNrraAYeD//Sllq3tZ3FkbyyedwdRTPYk2ZxrFoNV/87DPNggGdOqke5sGEodgN5Qi
P7/T9O9auh1pvEsLeBXrbcbGujK9ho4PXU744PgqNP2j7+LsR6HEYz6f0LtkIzxJ7Qr07IZuhCS/
EhRXfXVhtJfO0V7CVOvmeStMLnUO/LIW7qGXYSGGbqCd4hMiI3DI+8rIG+gGbQP3yyEQHgE+wQpw
bhFYG0QNG+FXrWJRF40wWeNHWLMoF4pr1etABurO37Y4oIrdBYRyTzbosJZmzQI8OPKeG0cWRTel
teBKAXAY32HxjNkFEPJZ0kdu6IKyJe2Imftt5Gmq7kH1BtuAU+vdhyhly68iB5HCLWg5n/lZpf/T
/4LktfgFZtCJL1gt+A7/rEtSCDZfZBeN2/idWdVwYSj0nFTHLg/F1/UgCHBfMq0k93rKc7wR4y1d
/UdGLUYp9myVLqdWqdmXibJfII6EMcNOdMeERJAI8pWJuK8+f1T8rdayPq435oxPMmpmq/JiAwva
8PY/UtPEd3ga1TyfIqhdIww0SoQIJiB3feBamovW6fWAqQEuLrhZMsQTbzSgQLU26XQRO5hAMBBV
bC+BG9UsShhJChWnet33hmmEhSk/KI3jTzDTNy+IXly834SQykvMTICZh01yPOkSxAdJTFCPE2RD
Z433VbF81i2Ylvn4KjuS5PXeUn3K3/lzOc6Lgkb7rKUVaNSkDOn72eLclysa65fGqQPKX9ZJ5k3D
RfaLP9Nc8t261yiXbdILcmALmQkeTAAbW29irGp4a2X2PI9eq4bBPJ8Flk0Q8r22ekt3WsJ63MhK
pFac4ELMmwqdidEQKCNhzHq7M7OMTkR3VQta0yt+gUUbV6DDxvoDy1SgxKvLsznjT00nznt2XFeE
MeFWe4H7N55U2I8CtVm/zyYesoYIrIl6eakAhBK+7fr7triwct4X2ca/O7o9o2EGBqYf5FFg4ggQ
3bk6hyaLgdTLbSqYmTOo2N8iLcFXbDGv/Ks+DZ+enbc/8A2bYWDWQh0NHeErzlhY2E3uxIKfElWr
UjDZOguVD7t6iFpfg4c/zM/Yqec76qj8gNiRDO9bKWXGEUM2zKj8gpWHzaYQSz6G0miqZFcVVqNK
oR/pWZ3qw7pArDYYVxfQNW6hCHlCdRfyftzT0PHOyRcDuzSA6H9ZVBxgKrTMV7lSiKSVAGsqCiIT
pKtZplC5oP5C+3aC2dV/zIjequ2W4eyJIC5jQVUfqDgMJwIH5XVzCqieqrgddQNcAo5qDKnLYLe7
9/WaJKur5B79UtMM+DkICEexFfPPVJ9F/rQZ2eNDpT39Y7QUKk8CvSDwIxwpu/SNXS/JQ6ipKGjL
bauMzhP6ZpvqbkhIRI+OeRivrym2StMKe5zhh0qzKiVd8xeaBPmGSyMKJMYFnAxy3hT3IeZgYIpq
zBwTkU/SODc/mXpyaTB1VG7kotNmR89CG+HeKK4XbnpXJpH25ktC7l3i/5P4lKJCrVHMAraEWFdt
rBqvvfAK+qcud7aE/nui5/KI0V8CbVRfFhDHuMZI3WAgiDHExIKuH60TMsklZQ4V7Tw7W/zsej7m
n82V9CPG2mRLjHD2dcxebcL/TljGQbGIIOIK95SDCv6RN+XArZm0EIVTWkAxna7PJw2n59LnZw9/
JA6qisoDqqeTJQZIReQf/wdvqR1eeidem58nufF8d2IZSxHhu5tRdMTHHR+OtZvtVVNTIvNxbVtI
DIYj2Brawik5XpQxCiws9eSE48ttjBEdHTpufUmFv3CTIVRNnMyTFxuDgfs+3FjI0XIIUFUCCV1o
OwgLSnz/F4jk0Cn8OEhShNeOccFl6U4iD2YlSMg3UN4QT5s2U4W+zbpp48sbkvGwYnPLXPdAX6FF
2zho5TkHh/Q61frIvr+e4kAjbFQu7dyGU7Tt2PhfKyXqxp/CJD3ikWK1bUh3MX0OX3GU/NbW4oes
1yEH8Z2QQD5s4WdDj245weXXzytoTzJh17eQd0G97uHFvBjdE1SieB2+CUioFlKeJD2A2l04S81N
xUjEdJco2BlPiALpx2YOo4J5C2Rb9Hh02eRDYT5hdBLOI7PTB6rYagziKMi1/E69tMPommjPE5hj
w4sLjudmRk162jDbOTjVuBhNqqqkAI6Ff/1nmuaaUrFcwYgu3MlCyaRnsxDxMM1CLavwbuKUCAVN
RT/sTgrIHhvQo/+OHjfgU4gelgryBws70rdGA5drrOsS1tCWX13zn53Udgzk3LgLCIXnudqCctBh
ar0JeeZhmq+7S0iPQY8qtdnllTfCvhVk4lISq+sPEMlX3akfpg+xGpBHniLRGlaOv3b7uANa8Hdr
8yUUgzX1PRp8tJBTc9797EvHZTTYRFnScGKF3Le130MLveKu00vWF4VJA+D0PPas4vI0yM07SGIH
f0hmgJ5ujRAR6Gg6ij5pOQOY20yAWPLHiMIlW8grsfrwQxmNRsxIYuUkAv32vuqwbFB3N5uGzhVg
l50dWnDhpmpMPi2PgghkkPmF+dIivlrkEGPlspdMvmSYa2ehWQ7tlPkfBTZDaW+O/OxqOJYmYeK6
Ts5bi2rZIPUCUUgz/K+36546gomccMioeRKI/YFX165k7CK1bOKG3sZ4i8TmeyvAAlX0hv0bI5Y9
QKJrIyNLIZxWQSFHzUEShN8eE8WiDyERPDTT6wKlB9i1QpOrLk5ooBIunkaMlePMlPeTe8HVDgp0
8B2L7cDrYuqzFewAdxmUzNodZFaJa9+UTeQhJzCCrVOADxQM1VgaNKqiqpnCm2V0q9pDbP3yVLMD
3mG4qZ6Z9AT2x2Xht3uYydVp9PcEtI9kPldmyOQlJxLYMVu6TB6weiGQhMdd7XbApiAi3cvbx5ay
BIF4tDriRFB0kFr1v/gLXrJd1XQw0t0ZUqoMUvzKNa11uOf1LnzPXDOGeaapawMSi4dAhYeKSLXF
EljB3sXpeLY+3Bx2TY4W2RRfjeOFRaN2yd5uXyPZ2gS0TnuuD1dTzCae53isaca3uK/k8lPBM/2N
LepdIPOnar6sZaf9JSZ4Ht6DCIeUQJ6YLxDkm+SIN6DDgMFFR9lhBsCxNVT8I7D4PXBfRNYIPTus
OwQvcoBh303okcgdcp6GS1P4+t4mjCrW2MvGuCCO8N4fyiQhx58oRTVsjVesR3iiaJGMcfcIBhat
tGlccMtvcrCkJT8YMNbcE6JcPqaABePru0M7X/MjtxrQy027clBrulvjdw29IkQ3VIXwcRBBZW2e
vitTFNcHbp8oT92QWZVuscrj7QXmEeP9M+QxV/zCfyaQJTbPXqP5BIf3PDPNQCBaLfEzHlGRlYqH
QRyBUxg3dtRNSxQaQ9cFtuoK/zQk48SeD3iaQDVai1Q/rs51Xd+7wT/UihIgVWB8IfKcbuDJeWQS
gBp9T/X0zR/funa+hRiBA/py4PsiISO2A/9O9MKMgkLS+w6/kLigo2XndACWNeZGi+YR0qnuB3hH
eaOx5GrIRaTP/QC7Rz47DxS7+go8kikR35hBXMtOB6oXrRqaNNdxHh7BJu0lAXrEyYMTWz24U9pR
2Twn1BgmduaWzygJqCA3bJKO+Rz+ZdxKqpz8Sr/JeIyi3zg+1/AGtOGB7SmmNepeVv+o7uKxK9Nl
4NygV/5x/ZPdNSZSaA6uGabHtY92uxZa6N2ThLp8kcmfPuwC+fbfvoQ5ZiysOcK1L4oaq0JK7OnX
SpwmmS7UNBGWcaSznKQl8NfLQ1GqJXmabzBlD6IqNjIbeeYXJ+w1zbgpILlwgu/kiBrDnLJm0/94
2Nu5ljQ+3RF8EQhztcVkdG9xtKXu55hkYLzB83u9y4SIWXVZB0eCTxrKetlrVOIfqPL2PzBmJCna
5HGzEZzrWwVYSbOxnEm7sav+pfcc+nsCcFAnoQf2ph9iqIAkQBrmYuFLknIJle0T6/IzU2gDTUa9
ponx7e/86Q0ARnxVKhAComj2u3LIHdHEEXHY5UnYJ5gPSF8BUToph51QS90xadEmn6JR1fAQekQW
BcSVxJW9WG4kOZPDhgjZghJKcj1grdJWrZSJ73XOvZrMXIcXwgynyVGpGns8L+C+kDAN5kUXL5qA
VSq9f+Sxfoc+Xrd7ZvLXlK7rVnGOouS5bvFKYvvboWZHbcRpYPj1x5yHfC3u/KmupZ+gNSnUfqSc
Qv9D84ArhnWyy3uUnhd7ARH0a5fdILGU+pb4l/Dsvr6f9Hl38cQ3L2qFaw/gGvoi1dxIOfO6CIPT
2wM7jwvrUaZHJZnPe1XBpB0WPX8MR5TzgCj/KnIr7HbE54ZW1sVAH4ck6g+i3l1lu+83knSFDCAJ
yAd879++afmNmd8vORlqKUSEgPpRE76vpkfe09fOfipbv9xB6lJTQDrEOMdkjjJPrpMJ874lyHS6
BI9EP9Vr+rpsxpC1GjZZkWyfMgBWNy0E3wZu7CNbo0Td/VjxPp+LIFskci9dxbJ0E5Ds0A8+8H2R
qMbsB3uJJ97iZHjQAVm812/phXQogpJyk4q7UOkeFlEGGyC0SLAhmB3l4CXXW2g3ZZwhUM8R8rhv
UtR7dZZrcDMonLO2F6k0Nbh/hqWzosHwUvQyEWpNDfKoeDbA7bRlfqVqm6zv47Wewqs8eL0GzgDV
AtAWXH1pqfWvFLY+2fw8NYm3Humet/xHSEtNx35l8K1jfJgrnUfz+cxUuMyVB+PPbqcVMCwiEdLi
tXKpnrA7kIxA5bDiQ8VAkdn1SMUsTXVRP1AILahUCv3RHjCUpVFC7UnXAbM9lW0lFOzWZ34Q5MdV
PFUZZ5G6QzFQgt1yjcMre4pomDFYvG1Q7m7JvwuWqGiwzdePUDJZMC+m9XOInxPz89YRMbLOqPMz
WV+DHH/hBW7Dok5xB7DN0RXJLBimhvZZgbyaD9CcUnxyp+HXr73LcQEhQvbJZ7sHmpwR0ZzMAmSW
jG49n1boT191SjqGqCOGQ2j8V2DtLbj5yGbOQBR7UxX2ClEVE8sVBMcI+QPmq2+TxpGZclJtg0Ws
ALmEc1Iaa3kky5Ppr6oXAxZACFGRWz5/XIWTLw5eScTEOcfo0/fEEaZ+2S+WbFGfj5SdQEgrvjd+
FjJuhwBlp0V6yK+gWG9mgYQkEzlpJeGnE+n8szhuL1fimDGT65Y/aJ05avu4A+kqgGdDYI2jLkt0
5pFQyA+9R9MmX/Nex6r4mBGhC1S2By0fZ2d+N8qh5LwX97u/wbVB+duMLG4NMlk5WkjP6ok9vGyX
+pGvVMMliFqV/ZSGfRf9rm1qsLUhn4gfuMynzBIybH1oG2tfhy+RwuavcGYryIkjc72K18KlKtsK
7p0e8HW/U3RFk1V8Cll3tVyfQhPrHH+ydT+3DGdGrwOQZqQLqapr9rBL+14Rr5ClKcqCOCwCnEBz
xJS2m5K5NSifrwiAonnehbUlbK8CNbx56qaBGUk66Qd+6s9afBUhaiSC3l4qy0b1sSl8cnyc/zHk
qIBjxTDysZZ5nRXoCoGz9JVNSYuhsVTzE2b+61e21jLXv4cXUm9qF01hXkqxeYhjp/Cet7pwiYB4
vGOVd5hZ3FvRP6gF8FnRcxFKgmwzGKd9d7/ib/toVb1pPHPjuiGud3NpIX7pMri4AVfc3XW7t5jL
1PcQd+8FqRPAH5C+1hTLz2PevyYXABeX7D0JYJMsJYE8JsAPX4H1+djE4l03uDF6Y1nloM6SYc8J
UbaRJ8aNQpcFvJYJY0pixbv2DUBwTiU4msf/oDF9WhPGACxaokWaXN3Auy1o2BDLzVJ6K6ciopI1
yFnqCATECdw0HThkQseltOcQRtnktAdlbug9pJmjBql91nI/i6abCZSWQrJm0Bml4oVqSCfbfqgV
qnC0yRjpQ7LjpHaKdNqlIIvP+SJbmW6vx3/O0uc8+sRz6uVAxGd0FdF4J0hvaLr89t5d9fD4Zmez
c4eGZ8uu7RVb2SuUpTJxGd7BfCVb5Ezyxt7tyzw/eh0fLNR/pDoyoErR3LDltia3a8dU9xhKJ7bO
ogWhkWmxEPKXsWybvOsIhOsGB1iInVBGyYBPnSowQTByazh2i7doBv+ybqPWGhjB2K5WyFhKEBK1
G4o10Z8SUpgKeTo6dJdAaSfhfh+SNytoDlFKspGHFBHZG536RfIEO8yXlrPPM0DvF9j9ZcCE7A3R
npMW8Sq5dCe6oA1Z9Vvc1hVPXKljqUMniMSVcvms3HE9Iy/MesIJR/NMqUemPnkwEWOmk4Pvrlp6
DJbFQYN5fWKB/AfB+TkmmaaWSwGOARKVzDHebUtZydzWauOxV2XnQvvg9PQoNyC72DVbMPf8SLyu
n9eSTdqPJsRWJJACb7+fhFf1Yd1VtpgHgk7yHBZ+37DfEilarsSLQ1/MnKdVO7+NMNfbf8p5sFVK
FQ3OWlI/WvJwYHAm8FhiG5wWFUgjPHf3Dv1G8+5CXphDPHTOVvGrTJeazPe15xiJYhZWP1tHUY6U
p04AvgwcQVePHdyMnXqcNLtrpmgwdCUPOp7LdiSNXbu+rVJxRzHr+ecZ+cYMZCa5/Qu9vKT7ZwQO
o8tpkdaKWQXAJRtiG4mbkPKNTDq5FhbxlT68SrKVcHqtmCoHtoGf7OHYkgQvMJ6iuO2kJXqsie3+
D3mE7w73h1x3lKBOrYcK7yMQXfbK7DljQGva2ELG6edowuc8gzHXASIOJyTzJdiJ9/hGzJT9E+2q
FFgasU4hZzlq3t1tg74jzKTdY2GEgmwI/sTuQhU93IP7rw4aTIlBAcoG7Rf2huEvrjOjuTZO6/32
+vHyban8OPuFEaGxUMdhxzo37g1h/nM/cRtIwN8nl0k37E5qOHwy0nwLFXp20Ktpv7nOUMpfMNoK
ySksozeT77/vonELhZ8/oTlxgkdu51vW+HE2yEgpG390Dj31n7IcEX2K2oSbBqK6KyifV358DNh6
xynrPtK+kVmiy4CmXcVTvgkNmG7O/dKOiwFoKBnwdF7lGfaTlhGDbT+cal5MB53C6yNRn/9GjqAL
u9HwyxdWCCUrAgt8zg4FaUYc0VUHXxlIsbPSLVyBymZj66S5/ttQpTyuYqE+Vn/I12ro9A2UYYAR
RWHK8mcnXaO3vSMxuLeKl28UdSZaEUPa5QVOlbFDFTrVcjxxXG5BJvqoyOVTWM4MVEq3xViEL2On
2lV0b4n6oYwAMvIF45M/Myy1iYgQ3/S2XUtnARb9c2l6jbrlyPVLiefRj7GbX+fScWpB56dVVUaz
4Fl1U/3CWv5ebRurWhxPysxvqUPUKHdekr+XwE1wRd36n+aFtOHsROKtGJ3BDbgz8Dphb/iXyYso
rh9axGP0nQ1NZsPQq6VCL5sQIHONWDcCi7+KsHbdPUu9ZgKzJdvy+Vf5ceLESU1GdRF4D1iZCIlH
rtz21HsxWp8WWgGA7pqwpiMl9PBtyRAwYZfgb2Xc7L1ujFBGvL/qxJMhNSB7Ox12fcEXWmTizAah
W+FttV8nLjm8GN9BfxLIrEHAGoRjpd9KtfomOpUhd4xhxtlYmBvkEXKk4qbJzlXR7txQocpkKtbw
yAkL6YbX+baFAzyCIx/HsG+U5FhwW2fqCk9SIb0KTkUnUNNW8BRSsSkIyatFIgVEhJIIxNtOMr4Q
AnJuhBrb34hokwBPMzpQegpW2ESCCJ8ebFL4BpoQEndAjHctcsc0d9nUsChFo6lU29hjCbJq+suM
Gh/UStOvYYZCuDhEHMoS2FQor3SKL/THcacw1gPf+8oCyNUOWLNK5yST919heSVFLWIrUbAvC2sd
rllotKXIpUStQ0oUiI6TASPKQtViB/GppfHSjgIei1Qyiey5u05CddvgTfgAlV/SIG3Zck6gKkMJ
aSKP9W8/CJsRVTZ09rNdRrGIJkgRJtBpcCFDizdxwdlNT3YyEXvZce/v9iVXIYSfdtDiyNAB7Muw
qvgm1mW/ixSjm/rI8k6KeNNHrHhse71WUqPYVtIvrlYrW5T3gknpJiGQXwkImoCh1dB3NVBkIjAx
Awr2QKn036p0Zlw4S4hg+dDWy2jNg1uOTGENxxM0b16Msx35E7rOo6ZH9jlEMBnB0N2i+1DuVk7J
Iq9rJxEWKC7cdY1FbrrpSdk58baRJf4lkK+xo3knmNdF8xt6PQLFGHpyuGaaFzWk9OXlCyy3JoJc
RM0NLbnPQWC+9m3a2GHbpf20pxQ0eVNzKt3MRHUo7WEjSFL5UpCffcdQudUCuMOdABZtUKSQRNIB
YyxZzVx4GoTJ5jP/IPOgIZGrSvHPS1m+bC98MORkx4FVRyr5IalQgXjqNjzkdqlDtG0ld4WolWqn
4NbDDC4PxDXSrBh32iQpIhhPF3VdWQNm8bHgXCdAbK5zxN1DAP+7EPS4njR6UYRowWEN53wGyf3H
UpUwdSY2QuiJ4177qiF5B+znX9EPeLIH0SVcJ86uO4smoHM0m/h0TGypVhGFfHXRECQrcSoTHSCC
BYPfeFBbaQ0ljputHvVbMtJLgQOZxnEpKZAFuYkilV0nCY4VC42B1tylz9ej9QP7C7yq3Y7BLRL4
e7ArVtG+n0BX2hfSQOtHHN4uFJdbtFPErbce6soStuevWeONx5scby4+lxKHvo3RfhEB+20a74SM
OAdaa0VeXBlwuy2h4Zp4BL1OqdqNii6iEhY2LQyYjudZgOtor2u4rvO6XJWWVCaF8bAizzgX7yox
n1ivi2h4KBR4cl2OAZ7/WEPks4Rg4BFQmk96+jGjW9zKwyhIPfiJP/KLhubz7PrYReZSgZBEdNfb
e89Sy62usQ26soNZqbgFPSYHqWpjpx3NbE5G89XxZhFac3t1XvS7vZ9Ymgi+sNwMAvIyeEZBWjD8
RtpTlCuMiCLwjP43i2D4OlLNGgzEikIvdT60NAl+h2svGwkcsHM1EZ4W2M+x5Lj2olOxov6n9tKj
ML1Io93siJSheiQTutW41zIp1Tk+Ol5dOf63NOJLFGGsxAHhYbk8/8GwWiCWoT6DUzmwl8CGrggB
GX3i1R6t+f67i4vLdQMBm8iFpOkNVpxQWHdOulo8ReDE9QarRRbGCmU/+4E2ChG/xR6oEhce7cNa
Aq24nVcPd1wzyZ5em4dP4onTo0gh5kwmJhVDWghBZEySShBkW0P44Ne/EgwzGd/5VfHu2AW5DeEJ
FLQk914yG11duLSkWiFWeIwWiTAMSSucpHh0UjyaajWRuSOGhf6sa6C9XMKI16fg12KfGGd4kOEI
aMTOYLS9l18/piIQYGhYOEfnIgRCgqmCR7agQs+jffFXukpKtwzYZh5yXnz7518gN9anIIyrvLME
2fLqh+20YHkUKhXgABljrzWfTmpTKX21eZ2+gLK8RDQiYWajpI7b63D10qGILbhK3o2nOxtFIyJc
i1L20LpmypjHUx0FeIS/XSBtWWPzw4mysxhZ5LQooxAkTJ+WUkwCGcfAHdu+OaXCnQg5UZLqhMZ1
xNvVufpAPgcD+cZnAMTNynX4isUNjehBE94Ncg7LUHrMEYTGDSRQPp7eoV++KAqLFj7PkxjPsEhH
TSv34WejURBb8oScRy0CTcfDVmxifLHtyjnrdGLNA+0BvmU3KilduinLFfdyBnSp3W+HfilYNw14
wQH03hO/gZ8sZbZNdJk2Cgu9AVosOU+x61eR8gNsUbYo957iAZYHdrz5aMeMJyis4dbgOqh0QJeE
uxADrtmBchAwelDgaFJ7okoUNNzNAsaQeOR6M0BJED4f9lD031HaoSxaOjlp2YTQJfUWYXbbLhJ7
qJ4nxnRkJsZMBc9OUA9Dfr3b9c4SS/g586PMC8M3eb60YABbLtbAj0daxzDRrXvzT30KPWqUTUTK
9ORW6G0oezkQRuxnzmq8BX5FKtP9stPEc/my9eVGZMiWtvUBvC3QPzgKwdJOPAlrekhm8F+oakO+
+sxbw+3QSHjI10pN4OR9X1TzcNjloLKC+CgNCDQ9icByno1/XoMo80q5t2xhUXGuD3RnswwbkrkV
7LWaFb74zBSsKlp2DG4YhCGeYWSCWsZogA4jV9kJsPE4GHZV7ugD9qYhiV107Jx0eq7ky1kwIFJ4
8zdFIWG9h4z2cD3ZxZKH0bnTWb3QeGTBWbaFIxvQs8Fp4XgwYhsCDTqnI+CIIZb074rQNpa4E52t
K/dWwDXNafX0dwnpVbT7QlrxhKOYTXICHyIENniq877S6STIRlC9d2h1a9Row09Va5WjgjBYF1t7
p8Ob/6X5KEr5lgDFJ//zdse51Q9gTSaTkmSHIRjNsYlxSnvXqlzSdHHwfdfn5liw/MxvV0xQagVW
DeNwdbzOOh6VQmcSKo2IryXpY8mfC+vgw90Fb8UuuRjMiGGRccylKiD51p1bKNhye3Z8mm2ley4E
8sQ1T8/QpAL20IZuCTbwmdpXy2R+24v74Ep53Eazl2QrCGwYmNgJL8FCOdv3ASx0ToBfaN+b5Kj2
1FqtyE1GR4nwNyGjw0Buhx/Ys7gDwLOi98u/o22IemTR8BOYxCZHXfj2h9A396zKq4pe7clnPMgL
DptFZHI3bWIuoShdTSGjy7l45xDaey4pFciS+UD4J+esGuyZWR8Wvj0Cv2SlXks4ExhaQ0s1TJCN
QehECNhWE7m7j+hFPeqhZuyoUEJGaK2ir25QLuR7d8efC9yVxFYpFkXGe2aJPfdSmghNegVdQTLE
tcIwgzTmCWL77LbzPft5on3bqmRJ7RCiOIJYrooiJ9+sUny5EcLCiqW10FyOxinGeHDvRIDVQ49g
PWlgKM3vtESeG8gkTGQT3LlRsU7Sp3B86skkRk1H2/H+k86omiP0ZvXa62Eyddt5JGFAVIHTJIbq
UJLAyNofv3wvqPJ1JDd/oVB5gP3MvT4nVMe+1oeJL2sSbD4GM03AAsTFi2fTS5Bi8pQTeozXza3j
IcM1ALW+o1c8M9K/quAE9G1lo21XnDRuWS/Is5S1Bu/0vR3Dyl+zdTxlazPYK4ySWSd0XTc8kva7
HBqqGI68lVBqT5xo2YXNlS4xfdSiV6nPLvbcGceblR96CGI7vzhNqRF7nJbj5oOkJYSenoxpEjur
yOr2+/W34ta2r+x5x+nTql2ir1eIUzDivsFFdgORHx6g6DxCE4R/KabkagwDn7P1mb4FpOV/N7hu
PgNWtPoxy03WBYQwyyWSBBvsVw+HAGcxzTwOZV1i/yCcopFabh+RhG+LjSYrmnmlaA+NLpeEVlNy
0eNj74KBueJpTTnMOoU0gzofqnk2KRNiOEMZlNi/xyt52FAJ4+y2zMZGrUaYe4zLWyHbWanowhfz
wT+hToBGhdFBVP1erZhA43e/ngqXgRwmAG8v4FPRSYqZuESCUusEvXjIe7ER8nu7e5gDrWU21cBE
nnkzqwRovO/OSYYBniixszK5p86wOlELT+SAEHQ+DNqFPjpeJu02FE+E6O9lPwbcQB54nB/uVsou
BPYH567mP63ndQvJRvNEzJ69MIMHBTgnbmyWPWhyqx1yhTUL66siYHuc84MxedOG95vyAobGgbhU
FauUaohal2n5p3eXduu+BOqQraXaNHJGiUqYyC/3EKS+6Zjl7XedfXMpRofs0HjESgqUiPD+k8dn
hnDTVynqWkMAeo5HgFjHcH2ETpQHaoRnG7CiO/h1EAHkLgeNljY1Fqz5xrIwPH53ObHYy6vc2Mra
QbRjALPlICioQ8QIaTvApOrFgCeRFJOzvYjXSYd/61EnxXAk8M1UlDesWXCiDqiX1BMv5k1X1kt9
DQG6KqggsGIsBsocMtzrA1MfEx2HAEjaYDEkWyid4LJ7h4hho4RzrF+wduDhq0Hn+UP1RVQpk4Cb
BGA3nz/gl0W4kWyx5Or7xcQJpHRyEoYHmkONzplxWpbrZYSpWIv9K2M6LS2UasCdY1HgZtg9HxS3
aPj6Ju7pNiXp9FkCUoo2yCwhuUV1d+SxadcwqbqAKGwBwlNfyyNgbsQA6D52paDwiVQ2uTDX5G6S
0TV2vA3V/Jj8pG5QNuEbgAk5+kulY5JEVhbrguTaK3uojGJpTJY8kUGdegikvlxMyqNWaOI3Z/ak
JymYzIjFhQFYqmxk9dCQ42VijgDC3nqzZn0sHaZ6C4v48/aprb2y1sQc0G7zSk+VOrIdtyP11/IL
6xRoWxNNV9amG1wrlYNd4PiEVUP/Cn3eeao7Hh28ps9LSD+tbFloSzcFtbZOt/0r+8gKJ5o5r4bZ
qwEfwMXSvPJggBrWzthKldpl2lzEVP3TwtSghx6BVrJUvSOfoXiOtbGRh8MzE0/3LHdiyHlsmecs
Nc3bkkCelffOGofQ4m8lRT3ABR3rB7DLd1HZtD93/tR39N8u+PCAUy6WapzoMpMFr+5m9CXrgsnm
ABO+VtFV3N/EFA8htPBaH3RfKamEf0tW9CiXly145aFS6BRzyfgAdZG+C5av5EFnx61AfGJVqHWd
BPZqr/zXSOSsgDu9cMPC4c4VjPWEVU7UiYdG8t+ei6pFTUK8pygCplY3kUO/9z1D6TkTdt+bZ+nS
fwTBBwIvksj057/FFQEYyiis11t6hGn8lJQTvOiCpMCvzsbO2LXrsOvdl/ChCgFDz57P4Ac525qy
qnetnLx4mst7VPmRXyLvg5vvD/GJBPIHuQK6DMDRwlSdH3N/vxHBy3hJT30zzq9eRRfNT0aob2Ao
hMruTM8xBj/fgiW9lg9WH5wB5NwQrUUyPGtwhV1r7t5g1I28AYoTSmCp1MHjMPRJ8Qg7jQeViTHK
bcdSAnuBez9QCXjjlNFityME0DxTk+ewDs3/LDCuH78OFkbqiPgTNNP09XsiRfiD4KMEU+KHFk7z
cEAQV7suvoe9r9mO0rk0RopjKGF4sHgTHtfk97fDKJ+WvJwnQNTGRHOOxljUB0DRl4Ty3B0Ud3Wq
QBxhWR6ueZKZaS54n0yT0fsrOeHgKauuxbZFpu3sfIwMa2ny7BWpcuhWSEGE+2J6OjUmlLJJ+hz2
hSmmH2yz6duj20lr/fSM16qczbwp2qgLzkb+I18SgbO90goceV4/vHXzrfW+YokGnXz3n/I4JEa8
EsEkKMtQKIFAQBgdbe7TE4uFy52kwpm+3LgMKgaaumJZRHCQlXS+Q7D9SFtoxvMt4EB0/P+iZoGk
0u8q5rEZNHbSldHtyn24T7kxEM1JmWIEO+s57bsV6yG8dZ+Wp9oStmH+LZIpMqWm90PaGNG4wv/q
/WfkWdzj77SC+PugEc7VlSu9kpzugTKCC6zcwh4XKFbRrWHBlrv+VhUo4sL/rCtSnQrdjP+5XUBC
+J94Mmy3iomL7IkmEDcMfmsatrbxWrarGlSNyKe2JtJq19zYdzvG5L/jj4AMIEvujI163WCD0LUQ
dS1fvi4pDUxkuU1/HhXpMbgiS/XgeAx9yeRboKXzr7EBeg2GqkF6eCXmB/XR6h42YMUFSSt3wiNu
cu1C7IO6eZpQSEThy1bwiPcOBCEfUzT95EHXMeYyhSRmEaTlYppDzEpDzWYAWBDGWDhuKMzX8IKG
W5tQrbhvnWm4H8QpqMYyFGMApV1eEsQHHvjrlS/NUYHARcig1Y8UyjaH8/naKWf2o3gbelWYMhWU
HPyFiFX7lWAhIwHKeBZGmI/xj0FXd0jbf1SRbpH1ZsiyeYcRY9hrTtnwh1qlWISfCJlFmlkPH0wY
TtiDjoDse7z9mo9Zzf8fNfTVyPGWIs4qETagBpI6alwcam3gl4B/4J8VNsDbQNjOPcJaa6kVd4z9
dmXjp0JuGEg7EPFWkxpQ4laPxju7baLdHDdwlc9mJnhm2wwHLRfVAH8n0TZvv/cxGgnuAFFNzCi3
xm4IPbkQGov0whz2Fh/BhSBoBeWq1hINFg5GscjtQSB8G9F5U/1ZF0eBRCXHhqSy0xUMS4JvZuGh
T7Go9EJoq4vmZRNL2tjyP0PEPFkN/6LrhYa/D8V7U5+d3AON6Tgvct8T1Oko+lFFd8w/agbq36wM
XiV8p8SNWIQw39q4odHXdjHrd1LgcbRAV8lCPAK1GePQ/c9yqvjgGbTHqaBVa8TcHxlxiXCSit6Z
W+xNM3zPmJtIMZpR3Sbqd6iXrKHPgRATFjVapJRr9UGMlNGu90vwHUHDhLFhusTTk0URAmC/Q38D
e4kSsvLple1+A7fsvTzj8gZsfXXFWzan1oSDKXF1khNphdun47jh/Mt6A2Ay60mCsYhK63TE13Q3
xHCKGv32Ldg+UjB/bWWC1roNIAn57D+i3zsSrhe6avyrdsCXQvTaa/SI3eS8+X1/r9YutNLwHMjg
zIzhk/4we+zL5GFv/7aYEJqYfKeeU/bcnHBvdSzzsh9J6j0NuVL0jz9vf12Wwx9xOsLu0xn1PQsF
+YtB3oiQL3T2Vob+PIRDMUcRbt/ldyMtQHKoYjO+w6zrzMlPMvfjPPcXaz/Q5UsT7bGKcQdomfNZ
yhRWDjQhnUN9gKk+aGtzZsmsygWnu59lXmuXpoT550bT4BfDUOx+1uhwvKmyiVhF4sxHZdKV8g0S
UeAuLxxbsusL5pflgCbBW1837HWW5U6uIR+75ICTos9dzSw89dzqw7M6jKXbz8X89JPKhDbuCaqz
7V8T9REnrYTtDzck1ExG0zCD6MA2sWwAMpzO/h7NK1OJsl9smwc0dcNkQiraKeoFkzRmt5eopIlw
uYUSpzztKVzo3kRHM6AyoqlVP8ZwooAUbByGIXi0aakW1hsg6zPnBtFgwVb1Oq3Q9HjfMTKoRlRc
2lS5+4Kwc0CZhWv+i9zBJ7k2UDcMEpCzXadK06utNwue7RXs7L8uY2wk9h4LmAblxBI88WzvkmU0
Asg9mtTOz62Au0l2Fr6A44WcX7WehtIa8Piqy9VTYgVsxLuK37iW3c6ZOiGZaBTYBEmesbvhnwfg
Odd6KSJ5Um7N5NcZNFh1PZgRDmcCvYCDcHMoi9Jux+DKNKfUDzOMmunscjlVNCMzkR8IiAavq9QW
Xr1rRLD85asOYsKmpR/291g0WzxGXiDgEsiZerNpvMgiLD6XnX3On9IWLcSjWKeCnz+9qGUDHuFC
LHfROOEhGjTxGbj1hQNCKBktwfQbhqesbaMQREAs6/Z37g2puRIoDaji7sd9sDOYXfQ06Q6mAIk9
fHTjUMJkl/493n52kAfPIJSwCnqVxXaAb+xneGhD038BAqh/lOVbKdzTKSHofKhq4p/oB+6bmwow
eRrePdGgFkv5/axcDIrk+KumGQXd5D0Sb6+hYCgpUz/aBBGxlfqltMEKdtwHTyR/9bANedH6F+3v
81eShjgPDsmaXKHWpoEm7fAG7vxTC3+fdaYlPf2qp3LboGnt1T0d7b9c2pTPp8O0v/EQWH5RE7yb
8FcvG1r7LFVxbrXXo3A2UJrH9tJDhk6fR+WRDXXknKfxk+aQGdadLBM1aFHBKbA8d8m0v5yeG/9b
bX1sgvZIe2RcIzicWxMOF0aqeLpUooHkKDGCt8thlQH2WBBSf6VOgGaQv9m/UD7E9AtXH+B02mEh
poak1Lva0afyQ5kiKy1d5HW99B9JEmNuRkFX12cIhk+nJaff2Mn9CZHj5edFSmIuokpmsqnaG2XP
+OHJlg4qqW5wLqoTq5QH/dEF7jtqivXlFFyY8BXuq5cI2l1kNtlXmytfVafgFeq4XayxuO9Y0415
/+BX9NNW0gNBwkMzf+Kf+OznJC1YIYJfahZspgyuYx8oK/Wt41EgWeQ+ea8P58Hl3cNDlIXNki+v
os+umFLX7bM7aduGh6XOsLFr9pBMCBsNh/7pd7vLXn95Z0HLm9oOgQC4xcvHphiQjRx1onlXIi6n
WYl1GY8Kb9KfXdEVnLRhAfLw458MHgD9dcdOmFcoJzr5hekqHXO4bZPMnlLzTdKrU8yY8Zp71TuP
WH6TmDW73vwZt66ggW+NqdmU9R+susxaBheug5EJKPWI/eKjGBls3S+cFK5am5EMSCJ5pDf+eTqo
r/VVO4EEFaer2SN3jN0YqexL4Bh44Rr6ZFb7yMn/RxEvrT5yW6bexIakd3nW7VED3U06qFa33JbZ
MZ7cl9avKSN2nfXOnKZw7KkqTXhkFpfdGhknSg8U8hLLq+rfNfTJmb9MpISFGh0FZ0bhMwID0li5
F4dCgkNnOFl6bSIERqkXoHjxXzVoF6YETgSd73qwinV4StD3cDGG/C1+zBck7stSBPVYgfAQ8rU0
fqCM+OZxj5s/dgj/7OjVg0zcHjge6T2u9C+U092PK9/KfttRDBjwztfSxA/arbfMC+4SGQ8g/d3D
0lBl7Qi3D7oHT8GeR5edz6ErnjLf2Jqvi3S8hD6g0JbnbMoJr3Yh5xIypv0/MNs3zmLcE3XbcLV7
cOU4dUdrT08JILgiu1ib0KefPX1JPBvacz0E5uG5ImVxZ/0Of5CVb8Mw9PUSKIRwY4sIPU8/crLz
ESlCFNoqWXtXyvYETiXs9fk5PUvHln/PiOHS6kX7a5LIxgHsd9GYny5e/sUP9BEy86ysw+8AD6FV
tcDYFcb7+drpyy9IaCKAP/DmywzErhot9a0LM9xcfmMfxb2Zi9fV/TqMU7VX1e1oTy7N5iM/2RnJ
fP46nyDB+2z6kJe4FhnkE5mK2va0btJzD/PHYd3a+y5GhHIfb7MqqzgFdpcqaxhIh0CpIOcuEE+G
3gZG3zT0+nf6CpH2rbylo3hv/Owwj8I1mFXQGl7IC4oKtlVHSBhv8ntfDF+aCU8g2JAch+/91bq0
kemm2IAUtM51oKWp0jqX2WBj+1/kn9GWOXPW/15rllQJ0GAOd7lwJjdRj3ShQsXI0dQp76u63LSu
uCtiwMYSR6C8mbPElCYuZjGiL79Hz7Ux4ltuf7oSWJOGAKIU8VsLVjkRfpA0MRwyl0qtMkcI7IsK
vLUOg1OQ3UzF42PtKowmnY8BqMrknySIM9y9mGOb7hegUJGAG/U0jaJv09mYThhs3YaJOGd0QWK7
kU6hmCyyu3LP1nB3OZ1g1mrGE7dbFSBkc3fn6V5AxeYzFOdqLr5fpTMQXgmXfjXVxGerC6Ab1XUG
AbRewtsZYxK4rot8krmA3P0SOe6kQkVApGacoe+kWmbwN26+xYPphpKxRe4dOzAcwZbIqElMOdoq
1zJlcObE+PJscC8H6oElsa48rb2gnjyh4rYNPsEWIRQLkZLp+db9U2jbMTEc6p5gGZ71VW/JCouh
2v4NRlYiG+2hBzffUULljgsCAD+XMZr0oVfQ3V1/ogXsX0TBEDTWJPViplrpP8BYF+QhXaOgIlCP
cNRphQ9Dzj/wQCHyZ8xZ9EHajJLWSEMdWTxZDdUFA0tZnUmcSKq+mRC2uxS6IaTdBwKD6HjrjwkI
cVLMuOKc91y+FVlsS3wmHVdPC2n6RgvaF3eSSzeIQ/UtLVNiioiUxtY1+WFFJ+bmVY55c5yzMjCi
u0X3vk2V3yUfzyQ6O61Q0zy8EyJ9sr/aa3p/qNd9+EK9JCEkQy+jaLbkV918fZpsy9DC4L98helH
2fyaw93Y2Q0RctHQKjc8HAI/HKKLuktZf5/sqvP8cPgXpDQ70ZuRxou5xGtcu8eCPYD0unOEOmAG
OtEo4JRDHfav+kU9jOiVnsQbNvb7QNtLqLNd66v8Q2LvOsUkeLTyD+xBPdiKX+wSgCmmFYDq3wpN
UB1Lnmx9P+g73FPKdIuhwP7eOmyOev8GFh99nQ+2MJUfjJnenghlxvw8UrV6ARvKUoNcmd28/vLL
n+D0vX3NO/2Wso/y1bn4c5PN4EXhsx3PuCTEhWCF+4esJSmL3wAlyo+sM97QSIRwd8XfwMknqO73
RUo/i20wTTWu9bnwYuv0Q9qJXSDdPzhm/u8ReR2JnJV09PWaUMZThyFvD+GzezElEl1SnukjA+R4
qYkkcntEtCBzt2NZ/SQ77V6Z41ph2YQ/ClLLMNUVkTrsyla6HqICAEEn3R+5Eb4cxIhmp2/mCvWn
U6RaiXeL8Em6tMQczZmJQBkBlkNLMw4xxZpW113J/8XJa3FnHQenA5C6vQtJtGCohOEtFQ/afavs
KQfQCTe0G+gVAua/6fX1yWtJ7HWJ81n39KAo46s07ExREyXQIeYzsYV9b8D8JV1Z9Kp+nCVtG0lJ
50hS9xm78TiLarcqFz1xzt+6APJfxnB+Aqan1O91OUjlrD++//lAhlBp9oqaR9cWdPGM/b3MMh84
h9m9OQcCjJ/VOWRmpCETFZDauOi4dHrQ/FNOoxsHr209bf+7y2BYnpoBwSfhbg5oNxwqkG6skN6m
rX1gbQv3+psZgMU4nmm43vcuidye2C4+8Val217exzx+rRvRPqSRXeQzLISTMB+IreQAitTubBMI
mT4UtxAMh1gafF/+PO8JUYlvFd0saG1wwbjRSnMY1a2NYtUCJR6+M27XLtmky5fAJBgzHnsYhtSz
aoLvsugFZtKhIGDLnlC58W6QP3tyxJOlSqytBQQVZOucKawP4TwxvbC6p83knnORgtBLeGBkXF3B
+NDAIswsjg4/BaNzdmopHzx1napS0mkDXcqIUqNG0VDJ9QhVUAGZ9cPHjbamS/DuwqRAtcBNvXRS
oQEL1v1TbCiB9ReVyB2Pvxmc0RKXl2oQckEYOvDcCMzdcjv7Le+AAeH75czybboWHfzEjML2mQ5s
WW62Vt6tqipw1baQ3KOD237vcLCg2cP1Mg0ACxtMA1s68OmOaEO7D99cwXP/8wvduvzVcV+YGl+l
NOxq0scLpvB6exaECB+0tPcDhxuv4MhUsSES6jnvC7UIfxKwOgThLISrcgn0jiKgXeGN77ELbls4
G2yhdgUW8PsysqGbpSMoIbOE6CDIyl8JtlkdL4yKhkz4D4M0shsY6NBnnnqei/s0rfP4S65tZF93
/393WKBfYXr8V90Hz3MxGeThtGs3AKWYIv4x0WmPVCckij36oDnECucdEv+XPI9sDfhgHE4n4jcp
cUrnjgK/fjofQuzaIMinp94Xj7QSNBhFwXW6/8oPWl4qcLETtvDm7AtirJT4YveiWK0KpZrh55QW
zCJSzlaRG+yeTKrCY1IkCTsBdVudJw72EM6rUmmj07+itcCInBREKiGDJlVCkyARFq1W+jXcepME
g68rPYITvBFP9d4/TZGzmcnHnKWGawDm124vYXFEmx8ZYU9LUMbJ3jI8vMDcXPeJH2c5tR90eIb4
tgEhp/On917B3t5iSyFhd6cdMXeCA0BncKkt65SRwU6MolhQqmcq8ojvPJGD71O8L3ge7Zjy/PMC
YjYcFsDjjF8OQFPbffdxAMUhVFmhSfRlVihYqJN8xSKoODUnvLp3nul5TfUBQhedukKaEYm5M397
OlUn7DPume7d5wl4Ne0vrWBoNZZf2IFAi2uEGwyoj5k2W+nXsKP4LZdDRX+xCQxPsdtmgxxm4j4u
B+MA+ykLUnmfnUsiG7Tv9D6MfWzrgbTW+JRuKP4UpQw7KvEXiks+muVDPeeMXXDizQn7N6SWeovs
KFGcicxIJPDkPhQRBVdRicD7R8EsiSyS8GOwwq8L+2f/svPYsTo57GY1JHdlAnxhLd5nS+pwSxfF
vBMOp6XQF+ZET11Wv43gUtcVcICfGNkPgPljvC2CuqJ07ENGkdaHowP2CYNXE3tf4horY4N4bG8j
47OoVTaEoz9QQrUhcS55iElgRwnaqU+S5dJ/OMoV49VtXRZ5ccu6GxqQvJQ8KMwMZN7Ie4ma9qs2
rzgLL6NLRzglDBEj+Sn0RYTow0gQnHsMpvfofxrp/Q9u4eAENjDRCvF7SuosYj1yTVt0SGkmTudV
CjJlaLH1j1cLsmZ1/YJDI1I6C/worrw4saMkwU+Gop0QFdZHLHstytaq2zjQB6NEeDhnmizrTEFB
nRQgyQONDM/+3+F31epOYt3p61knQVyFznjEbS0xfR0daa5XsNMY4ht9Hue8hlE4RmJeWT9blkql
XuoK/LJ9L3sYsazXxePlAD4InsoMzhyU8t29hTZbTQ1wtQEFGsCQo2+yOSe5hKU4716fxdK/6/+8
aRNYMviMCAuSiIwbxWN9tkY8CAP1VR/yIIlw/eP3bzE6cQgtINNyugAV5/pXG53apKaTdwACv5XO
nXqazFxdUJtK6LynpdrE7ohwtW6M4u3/ILd9L+MmjLyJrxw/+PUd7ccngYvRgAHtLcu2mPZaGdmH
7rj5qPHaaXh5EQSNwVURJN2AiVYT9/eHuA9fC6vhx+5AhJfWTLq7M8wsA9F65pDWYlmDG+wsjJRY
UM7+xssS+g/h03ARGWLVEds6n3qxB5C17cDhiHcVe979t7PCjBWfybLmFBJsHX+f7LYdxh1Kn42q
0QCL7qgBIUCNzQqZWYUA+yaqsrg61QLdC0BbOtjWV4CbG4Et/S7hzY3FHbi4bM72SJ8OxvZETsie
OlJ9Mr8f+/Jo+j6YRujz1RSVnGGWF/l8moh9nN8qHDMDMaPNiyimgR7m/zP+MwFxTqr2DDnlgIp3
csF9BvRxg8TPuWBUEUaME10Bnw0M9oDeodKzt2bZzU5RLueniI4IcG8itdGVrEljL5Z/8cK/mkHU
92Z49TH83emMGW/mFDQ7WMCwHqhrrAjHIsaG8pmAdAMyPBoQqz5aN5bWgbPuBRGMk4Tm6qQOoyx0
TN9YNz8G6S8Igk4E6wodhKoMMvNHiTLNzoyMp78lGZs4cp9RYn07F418EgRTfDqXlrIoOmb5PsS/
OS9mGvGaMXMNRjoKKiWXIg3442YtqTntY3Rg6Ln90wojnk7TO1igQELrrwjr0KlWEHOJoYGyzm3p
a5wIjrZYqDtkyv4tPmZFvZzHorBzqF76O+bavoNHx19DkLCRKHu6wWCdOwPeReCG0L9OI6oowe3K
FJONPpg4eht2vO+BAyGJkWjGNFKYbO6Gg6Pqm9/lR1oQyA4lUUuw+bogTP3J6omwc8erXXU0jaFV
teRTbpLHlDjJ/5n6Bshk6QlhxUWpB+ybfMK3ztMqXipXTT8Ssj0Z/iOXyHoOGXfVDmTe8VOrlbyn
6yXANobbpBXe723G2qvTWn/fnpk0OB/BFTWH8j78dxmCh86Of9WUibrSoz19sQS76h3Mz+UXHT+4
vMP60mGMGtkOoZHLj+fRIwMfPDbpHKpQfviS1p9FpYAy1ML50eVssGd+srTPoRhcy10nFA5QawHo
gLZAZ+7QEfaz2Y8YJFdbMihMAZVNHoDw0SP9h9RNhuyaSBQtluc95gCi6seP0DrUW6pUt6VtN8uN
O1z8ZK6ii6jaCIP4eOzsEk7fo+LQaq/Uy5qua+rXVasE+Bs6HaABwImup9H5J5rixmoiPPWbj876
EOHGPfoth1tAIoDH/1Zsq2/wlCEvtGv3Up384NK5GO4j+Tc1FQehq51Ciipht9BVXd3wb9f/F91g
pg+/dqnCcU/nhTVXyS5+Kn1pHifbFj56MzH/KOdSliCQEHMSBnqQR9LHgER+ibd1VACB7z6aSSGa
ZNBvhEtnHfI3Qiiho/4ts9xCuyUiYwpTheOhR60Dw/eOvaDy4c75NeJOFLixghwDi9akBDxNVHa9
LFPQcT4JJpY9C45MVLnqBgMfVaLuzRiwPfvdsWpkKcbqpS+/guCDJPX7EJ9TIoQmgBmGLOS2ike9
p1cFVWwQCSytGKviJSnoZk4ZeDKkrpbwO5fne5NFdT8RkVuMtlOyRHZ1lZeEkv7jEw3F5qQl1QO1
AJI5yjljVh2BhbTrj3jEXDsQeMA/Zib6TiVYmGvRwwURIvHvRZ5fiPwAzTUw+HFHRrXLziRRcqrH
UdlhRP40YOg9Fq1j9mwXzt7qou9hyv+HYHzvLgH5THCB+4BW9IWzlpj966ypwn7zPHWlhUtmzePF
dhiZjYnW584BEvvXZGtdTYOQamb3x4KyDilci5E900ZxlVNoXwceNvIox1dJKjJNwz3QzAnnm96L
L5eyizZpGw3m7p/UZHBnfIINw6GWW8fXbcmrN9V/3u3aFX6AyqbrXT7RHSM9VxkulvcKY74sVQRw
Vds+PYSxdB8YHUGyua3DYSYvOZOtBU+Irw6KtBy8z4A4/Ga+PHbzvIHrMcet/+eDw0MuEdiFzBlx
RTrnJ38OCK7A7+sO7Vv9i/jIqMVMcFBc4f4rtKiEgeqlEsoyTZUN+KNSShsTlYsozu93Y2NAgevV
QVNv/CRs1ExzuzJG1jYk2gH3OKSDIzWN33NmY5+CYlzbcAamiH5zYm5UYtEyrPr1WOUb7gYq6FE1
YYXbMvOhFHrJpxM1ofJQ159ftSArWfz8PgL5cj/NY5BzisyPSyY/fZikD2CqU0hEYerD7/GWD8wP
EcvptQQtQUf05/qUiTmvznrGpc9TYyBNmP8rNtY9081HfqBVFM1ds1FPtZbvyKMNYmOfP2bG3Xir
w0+NcIHenJ78lIHCr3s3QmRip76SbdI2qJZzmvPcFpRhiGDlWl0628dAxsTxixVD8VJ75H4T2JKx
PPIkOuF+HZRjMrZ+cA+9+KpDVf4jIPLnOqMhr9i8ltKM3h6weqxVEe9L2UeXLoT4EZ5z65fHEJS+
hp4fjcced537PZragxaE8aB2k5W9Alzf79xiiRcMYv1YSMRGZTkm/cU4ujcfXPPZe8WvIGEuPxYb
4T9MYto7IhvfsGrfN7XJfKPgNLawHh0u8a/QhVxz9nth8uNF7LE+tJ4hKuLS3jvxlgKcZRNdm9os
W3/eS0lmN24fe/IbDtJFbSwd+IW1NRsssHtmyxH/7j/WAX6Sw7orij7bIDIi2qrlGjcLnpdJULDw
I1o87k3fIc8fTg4WzenXHh/Q29EdDqzZ1D5tBGPozKne/y3QSJUw26tts8uBBY59iy6+b6BMk6sy
BzjItSi7KDMNWy6aILAZ9FFcGlkCqSk2X/uMfVzrsSR9WmkOwiGGbhgc4vf/Mrcw2thteH4tbqXC
5HRcm5mJyhzEJYtHW7gsIrPuVoKmR1wT+m23HUbQzoZ2svUCXdDzF1B6G7iLhc3p7oESD5Kzr2Py
8gKcBn7fMMz2XFMvveyKqKbV+TJliol7gqAh4wQkElw8F+G9OIUpojyCaArs24b4vqRbui1JeAJ7
tWsJD7oD2to1H9Zcr90QlKYOkrRTmENmWU+P+sOMu81KsxSk
`protect end_protected
