`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22384)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/yKOvhbch4frXkIkj4l1RsEuN
Nf1rx/+PQ6jdt9bFrulpmVY9v7MKDA+8KT4GvgXrVVrRBrggWvJ+Bwu8tN9yFlCUrP9yrrt+riqZ
nTUpx43L1buJC5aJjty/nr+m/mlE35SZ11Qh4Yo1TGdE2dS9EOOyBKSFUOgGyRCZjw5MzgvPzB3e
tQs2awhymVobN3gdG1otHrYV71rE7bKVZVZvWnnvo10dK1itKsVIyo4sjw3+CuTlE+Y8JHd/Ze7B
8qQZL2/9N5jr5AofBPaaqiL/8mQDHDM4O6BZsmTQm4EDAyk8dLuuF7HHCc7Tc3X62s+vxm5YGMTr
MOgpDSRsuYDsmekBAKAaRq2F8BB4GonrolvIAPng4jxJ4HT9j00HHcOJ9JQKRUKMMOuh30T8H2eF
HE4VxxouilYBJ1YWAcGxxdIiRKr4kBDN2z5Z2/wUmr7oHaZITMtfG1uTyZGdJae6CtCCYvQ/SblM
D9wG4ZuaRbI5AfB5LUYFx+zQt9NWhmNrlhLwx6e9+hx4VITFrrHPxx8XC1gDQ7ieqQ9QRUa5e4lY
xiJqda9VRdTQLaWeTkuq7DocCLjZYg20qMxCf/k00euL+4MGIlgvXRSUsvXHzaKeRNU+JNvL+g/0
9plb329O0yrAWTOwmDT0eKmi9KEM63Ct/cMxbAElGXz3CIVuUj64K6901DhbnyebbMALFtqTKsPQ
VQRBeFH3rugIbtkAeuJc2LvWMcjvotdh8TJOzT0+GxsVdNtsIdmsQyltpstXfWdNU6+8QWTmuoHH
4ni50v6641WE4UYYhWcXuy0KfS9+V0NJfgbEeVGtv96w06AvQigHVDYmocXA302M3DUryUXjraqT
DP7yGRiD+i82gForDU7h08Dq8A9sO/8dAhjCHP+wChGbeKsHnrIu6pIwDyw2t60hQj2j1MSDYEBI
cploOowc3Nqp8KtTPhQNKaMeKDXYF8Ub3zBpqxxcJZkf64NA48jU1zdgRvkbwJ6L0v0yAHsLKi/Q
tPd3+Gw2MQUHcb7a847dkfXfQkXyqCL7Xuckw/yVoWFk7MIqCky34D0AtLeF3cz/3O89gg3nisKy
Q5zff82S2mwKWAhls2oGEq86blCKbyRC04nLWa+U9Gl99RFdDVUrqrknqcAFQUMe1IjHaWNqeLbl
ewSzobhnRktsOF/expWB8ycVOHqRY/ZtZEkjFR7Nt9nKR06T7DTdTYmV2E6dodwDtONBL5Wxg4+P
80ARA7HYly+MC33L1HalbhXMPPOdfxmy9Au4Tqp1CXg1JgfyRgV7wB1xy6N9u3WvQAyGAM9hwShU
9ilJR3J3GqroP9/do1sbvwxOqDbZ6FuhJhJymDs9u+eZZY7AATdeGTKEbBj1nFiv9WS6ep0RaQHO
m8ZUm+QP4nTnpFWjqOk8MjDqbQjKrVZLykriXEMfAqmfL3HnU+sHLDpx+JO0hoJ1ROLt9SUEje8e
Yyvn0YOanzs+68gtCkDPSgcAnOsqbn6BkDe0/yS4yoII3H2h1Z52WiqvQl8F1qcmNWY42Mn5e2hB
4MqBfM7+zkzSGl129MBRNkQGZ984M6z7Li0HvzZc1VYB5ITOQKwYpbfWSQdm3I+MkHbTz4TijXNE
eoCXqYJFHt0f1db5MOIP/CQV/MaqqYV+4jNGR360shjvmQXDneYEyW5vOrdWbzVVjp6Gz8zgdwki
W0S1yIR1hxvoHFIIDFmk3d3IfmzseKkZWiN7wiXgHhsxsg8ttEcvG61nnvl1jH0WMJYPdquVeAxo
ekGJaOD3K4K/esX0qItz+vS/RTlZf4R/VGRqVhgz1bI+G6oCOj15kCJNMiWwhlXoP+4mB7oluDYA
M4tjdU0Qe3xKkzvlXjIilxD/ZIJWkMZjGOPU0ClUkzek8Shf1+6zgBxwHsVKHOFodmJ19C2870Wj
oe5s9q9P7GMXv2cjtPrZ/3tgbBfIPoJBjm+GEGfpJY4lrHGUSm8jeEkOZtuS94Aj/coLFxB4jKun
E6ktbK9zMnRIc5oEOhwDcOabhOXQmSonBCFw6dsTqJllNx+H6NIFfF1YRvL+zMwsdZ2DMCIBLRiD
q98Aeqf4dRwaZoDSqaJAuxKHoFXj3qLhcmDwvxMiE2OZQyJMuMCmvTJOPeHDdCX58SYz1CJhA3Gx
txy+fNUeIEgMBkUoRPSsEZixz38t6L1V4hg9hjKcu9a79eMug7NWJ/XyZX4/sgXmCJ5jzLjxHYFq
F7cGrXf2YBR/AxJeGrfn81mySYJBSiOAbRzjIFip7w6Q3DEjjsYVAfy59XHs9yLxLMncW5Ulf68m
XiOXp7ugLKJe85baSzQrPJjSVYsEW2xI/HmSBrJL/cARlUON/NxxIwcDO1skZo4DfGGHGUKUYF8p
sBJQrGV8CJs2r0Ahx7o/ON5ZxHVlDbij9z25UBBKqdHs9Beh1JzTR0B1DorAZC8L5knsFF0B+RZq
yjuLIFRNrJfibM7RPTCct0ytvXM+6DmpQXlWCYKM/zK2CQqovYu8gOF1QFZA72bP4jkGkm/lagIS
eeuPKMhNI7/qD7JhvyOKk0LBFwUp0NmsNAyAm2aNN3tDNt9n3SfSemO8RIHH6VcWfZfv4sXjNQot
PQpb4lu44gxnp9MN9Db+kIbn86s1Vg4QKnAurWJADrmY40CU2DNCbJ+YF81o5yI1J43YHJlXmIiD
NQoJafuoMxo0EKK6Ojo0g7pu9KFOzgDofj6rfWzwQU03HWk12Orr26i/MJO6XWEGc//ce6jru+PX
ExRkaiClRsR66bJPNe8fKOwEn/Lr5DHiuIqSP6loC0afKyXX73zW4RY+Vug+6nAfHdjAcUUiQ4zU
I7Cvag1XcC7AnKvKeIT5D0QpL2XUhql1YquBN5VKrQmtnkxa3wwHgx1q6f744CIspMsUhKLuLVQT
StWOTfrHVjhuu08uKKhVRno90ag7Oxro6AaQKv4mNt5ekQkQq5Y8eGw5KryEnFMQWXwyTsMS0Ghp
p/hjmcJkFOhuiDOaUp3J9g3ivDGY/tw03dzOHMTwTKvNsyJ1IOpAQVXhQUuk6ZOv9Je8d6cg/b5e
XIIGLHEUlC7dscNqUahYd6Kg4JtnjiAKozptA/92XKiYI3vGwRu/EE/DmkWfH849Ahrs+Hy5UuDY
smQM8yDuXH1QH5uh2sffHhOAzmH9MRCOI74NufqcNgcC41sfjWsjdpahu+mRFS+2gHRoVWngC+JZ
g9WSiE4z+f22i6oOMMSaicXzAVwLyLPQkdpaKcp/6cUUFZrv4Ok81YggNRE8mB/qfG4vR5PrnxvT
52ccjtzvhrACkxz3DUmvlni9Po7W6K1sbO+owCYK5iriT+n23+7uzlj4a3zR7JQFjGu8ObwzJHEI
DUKplltl7pPbdSowiTLRv3WwzyRVaJW0NI+I3ySiPdxo4Km8fWTwturNV2ZJ68u6gpp4z0ukKr1g
HMJhVN5XA5th5FWxvn6jiPDCFTmGTAn3sIYS8c8yVggR3td0jYwDAdjleh6dwodVlDd4tvFpYY1B
getiujA4HZLKkJs2wDiJLMo6VYVyRrieRMk3lwF6/sY0dEhpA1bkiBZVOKM3RXI3W+zYCTWCkCCv
u83mkLxdccQ+5OshInZORrUno8piwEiKDGubK5GrylhD0o1qET3pRfBNY89GOLqAKsxjQ5CqK9sB
8u2C+VGTYL/fVfxkBOINC66KKzGtpHypEXeaHFnHqCsgjnxvylWympr4aTN6fLOkgLyIBd+s2Sn5
VfU4aZrxF3/jnc/vkl+KFAD6M4vmBdD5vO1u/vT3P/865f8kEMWUkKAiblehbg5DmGw9vJsd4VBd
2TXnPpFmqA2Vt/5dumNJhEkfMfCYCsrKql/wcKBD90J3hFuigQUzmTKZWZBRfzz1IukN9TZoksDC
3wfRfOBnK/uPTDeqTXKI8yOOpwv4bw9T7oxrTvP02H1db3cv4cd4EjxlAxQ9r4Bod1CZQXGS8+xO
FQAHOsJgX9HC82553f6IvYyWmjMaBdk+p9S49j78/DqSf29i+FD1ytUhzxLSykvFDoFBiaJMvOE/
vROjsVcjMuY23sKg0NYXWj4bD+WqJqjHbSuWk+oKfqrT6XWikCq43bSwOmaJRr/70XOrRqBndk+3
s6BYgY3ipsrCn3yFgrcdWxl2ThA4Du+2Fs2BorQ9y1ES6BUTx/S+mBSzfIZ95c/hm+9lFckpQKz9
76gloyejl0rVoFq545Ao+mlraylSKcCvqA7WU56gUC4jCqTY55m3XnPTaIbT2xxlnN0Q9F/5NgmA
Bx0YUOcjXmdEMJ79P1LnUqwqRcqxyZ7NNxBSyGO8ga4NUPZ46GZGplnhCAqIdkeZKO3RuwUQsdw2
9dXxAcj6segBEXcHaec20m8qWPM6yyVvnpnsix1Qe8zIi3Ur2322GNeg7vKwprWonQXrypPvO2Q6
hMpUauBioC/lZ8jDkwxZ9GtscBmbilok/r0ku2wZClYQ4ngW/b7hXo7RU9JDEXWT5u/twjxo055y
4fih3uzxxPfpzSzpZ81J44VVtMWE435rDpm7Aunwe9FLMgzvrtblQQBu/Ty8fYZUBeO4P9w0/fsd
IryY+yMl4GJHHxEY9sRh/ubrQgaffGiS1dbzRGRq37O9LFNVVqFdLttQ4teChJ8qkQGtYsmqtgFq
iksEku2bdNNUkiuh4ZnF6lbeIESh1bDhmLzL2i+INBbvQ1IAEbcOPw52qHrWxO8bLbo2V8tTyeBm
x36cp7lYqdv/E6ClO2LDOsrZ4BVjc2qtFXCKU4VcYCDjzkxMLt78/0xaU7N6dyzGZqZXkOQX9jTj
eekao1XOwFa/kNRt+NK4AmVZbzTo0CRNC5rG3uWEFyS4bpfW6oJW7bM1G4KotuBWIuKcAbwUh6bs
JYxxmpMjDFq5wxsgIOE8uzTsekd9/pI3WqAo8tyepusTiyXM4qT8aq9/Pi4MeQs81EJBik73TB58
jTP2ztFa0y0L1GcrePFcYwngtBJaYE4sBVpqX8vmlKRw5sUDgnrLMtd5igTn6vZOjEnj40ZH+x+u
MVU9nq04bYTzuiqvr1o/HecS4yRt0g11uMEZIX4v6RetmfS39qeZ9RGyMj3KdVeIadquAlyFynv9
enXDlM86/5nNBGZYMYOeKyo8lde/RKYqsWeZu6XBo33gqUYlMzyD++tapLfIxdASsoRc0Tycfu95
Pg4EoESstp3Y3+jrO+AmIFIYiqcKdIeqH6zKp6wv6H3VZkQIlPqXYbAKp0CZeIj1kFwh1nzwRBlR
K+FY9KZZnRYTQiS2SkAEVqye2d9X1NGIBKLS7I7oQ/O5C2Xx8N0D9tnGHukJIS6VC4fNxIe/p4A3
qLw1gRp4pedZzZ9uhYtm4ZhD1ejSSldPX9SNDl4KKVxw0MqZrrxvar+evXIE0lBkEqoIcUB1I6mz
AwoRoqL7Xzq9/CKgYLfF0K+rTuTh2u/+Pa9UTgu8gWWePkE2Pi5NnAXTqlDGgmClwQFIOlrLYbIE
CdSZ2fEoNoCiTKnkoRfZMv3np/5Lq7TwtNnXblk67uROdsZbPXsmW0jmNAJ1lR74G0YhdiaepfXr
T8LbXoh+SWp6dnQwFM6rMbNc3kpU+WZJQJqmgrjJPpRU6bT5JpQYNsH8VnLXYC7kpxqxPcO0+zk2
JyU2ixUC5u6VQQg4KohtHjeFF7nA4wZweit2BqNDC1YP6C6doeUb5gOLtjdlKpTtIWahOmNGaJOV
73yaoFlgnwoRtMMS0TYWLfc0YdgcfPSqIxR+UykO4V23sYjPCHYUxaqA62FfTG2nj8T4db8rjMEb
nKSZbUhSGybvBcBuWi5VJzqFtEndbJn8+hzM9a1+LegS0YhmzHKcb9voSQDMq2lHKHx5+cuzxXaa
1tOaGTWypN4iB0WLYsFvWJ/MM/665J338/m0g9uMXTHRITOabbw7MN7jMeH81QfvNhqS7vOQTilQ
+BU7hlGPz4Bq1C5aIFnSlxrVdFG/AjK0VwPEOLvWw208xPppEZ6cSNb3YXwsyjMQrldYwBv6LwIo
2udtitmIfGEuZifjh+Raj+5GlQme7l2qEkNGpr7OEXXr35AO3PhyrQAIsGDccfqxI4H7IPuT89xw
Hv6EEgsBF4yuf9bu1KjLLwaqC701ruP084COz7TYf7E8nLiTJNCfnnINzJLd43q9etwy7loZLj/G
fSvdWnj+ZmDci9Gi3xqEyf/8WR8KA89JXqLyW5fdi5u/ylkPrzWLP+mX11wG0qTW3UDTJJyszFl8
AVrZ2MJ0ks4f6dUj/UoX5D70JjZYy0ZUZvADa0jZYH4O10WwG+AjtBb1kkOq5rlOdSCG1szrdoM1
u6Jy7dsV6bPLNYC3O5EsU/8YBLGEGWwjKbG/+8pxmUBfJuY53F2WtcxgP9wgh9Xmlo2D2PHdj1M+
3AqvO1igp3IadDbAq4nHvVpdumqXz2h/RkJZ/GX1A8cL3KjK4+KYbWj+NTVFj9iBvGcovNMVNbf3
Tt13nwTnC8X7LWnahX7milRoaRuGMiBWrPLGTYbH/cBdwhQdk2i91jb06Ht6I8jZpKIP53qdfZr5
YyEq6odC8YvtmSRwsVza7OOC08p+wFl//aV0J7tD98hkJEVtOeya/N+sFWx+fwl9A4uHr45ZOqDy
FlaVkTG3bal3sV1P9KIrmG9NDatXzlBXE5rvEcPsh5DpSBisC3gDMyjCt2ZjrHtgQQoTVhKgCOsJ
tSvPAKYAkfQklVMCkxUBgSg8KdI/YdDWGp6pS7ASERpWnjhmJ6nkD7jLDQNraTAY+fvXVgZUhpKd
jhwmDcN/XD6cl9jWnfmJ5Sgq+eGpXOgK9JQG0phcCRTlaGh12DZmdynkBgkGYU6aZAohNFKttHx2
F38wjeE7YBBFHHuajXVN+7+eZQXkHplb8OAsQrWnXnSlQ8ff9EdKpPWZXjzN+6G7I1aNQUgRPSgU
eafxPVwcsh94eQkZULb9+89kudku9uPZyRaLst0Q2cxGURzDE6uBo30NE0a7WPFoAfpdk9/+mjbp
R3kKXobQeQt0lsPxH7kc6j1HHVscydqbBDNwu3Ec5iyAqgcYJil7cTBs35eJ5rWh1yhohBeH+KXK
pez4so6TJOaivntSeu7NIBptFQXGUoPXdK580Lm71aHgbyY00F1VvALZZBDoINtRTMztaAFsZJ30
izFxxPKXwtBmY135uTq47C4KBjkU+VM7z6gb6KtA6izKJOzUjFS+zStxi5SRnt0MpO3bt3tBopV6
GPh9akNF3VcWrAELGQAww44NLiu6hBlWM3driSeeSBX8HwdnMVYpGLw5dclsMAc2VorQlrqbjvlh
5rXSiituHYGXg6pdd/IV3S/9FR4wsqypcACFgLoXS39/XJeczWidIj0KSa1SYUs3Nix3H+3AVmAI
wXe+MUJokognZZ9i38nj1uuk+X05g3JXTibvyPgPQzcVDNzf+YJj+Q4C7n9y+fouzs2wdVTKh0aX
5EK0d3Bkx+RtnemTCdd9aFRv8mE0EDZDeGnTU/T6bEOBCsAribAEZuoS1YHL5hpYZPNF4FDAn2Wr
vop6SvKMPM17zT0cUEWFYndcsU1vcTgDqyH3Xu19ry1p3GIg5egIJyAFbzaSevjOJ0wLV+ku/Y9h
H2PesQ3dcdNOBH3FLUuMloxM1QwP2NBsXJ1ag7+FqIderNaY5HHH/sUmGi8aXfNgRDNKLqfRY8BN
FePi79flwjqrgtHa7LfekIfVdkSdkfGrqGRHc2S4DJLgkb0Cq8azMuVRykv5U4wrjS9NwHe2klHZ
agLYKpbml3S6spBSvX5Lp4iwbQOASIh8aXAoPtUXC8qee825I5t/l3I85VVj6sBz+7T/wOVY67xm
P6b487dy655Xm9/97zKnaxbeQih5yu7k445fXd86sMuPk4/f/n9fitObREtRCvKd8FK63Fz1Zgyc
5eP69SG37u5D/dSMQUa+GK7ulcnw+aHrbs4Oibj3vWC0sSesLJE+XNVTI3inzfeioNliQNJty/eu
rEtZ5yUi1Xe/DEgaNDQvy4dnGXa0/XkPQ/6FyxWriqYVMQwu5oANotc1ttIO4ECSRrX40RUPz4kB
McwF4JbjYsw/Xmy8j4X4ZoMZjlRQHaY+ZwoYiH+JyS5a7aqoPR6lB3l9T98aRXLhUNVH66YN0aoE
NDPeAtTYPQ3ZOhTs53Rm4hTs/6+yQ6ILzJofoYAK1OctjumDgIltg9JYaPHXie6GaokbY/Io+rBS
yKfsCqttTa910AShtsiwi8QtyuZFLiS0aRmvcPRrwO9DW1K7qXfLNsIhbtdH7jD90nV4+G7mDq9P
nEShYnlUJRWM1wVuzlGf+9N6M/ncI5XELtckLN31+yzX/DfZawNI2rWOHW4zx73CKnL0mTD2xC2K
z3VJSWSZKe+EEe6cxc7KJ1in9dbAsYVIEi2s2qrS1ST6vK3GfxIkqhUF5SQwol70g5d7LTz+KtRD
YBWeEl8hTAIn2+N8y0kt1GZIv2S7ICHEXr3e6CsaeklGopAfO1UiIifTqZjettak8oz6i0NUMrXg
kGdBb+u/sngZyD2iPWJS7A+lwVwvQzQkCo4J4Fct+uNjf19QcCKn1g7cbZbp8GrOzaGtuk1/tTAK
eFVRKJs/kMsRjYuSozleYHejl0m8xArEBKAjkjnEEFSSEbDGiXA7HzOEf2+kPE8w8t63v3bSjJO2
pvaE1TIhqWxx0ghklVtiv8j/HSaLVzd5WJguobcC/6l3Y99UsEtF2OAP2wJHuTTjrKHyPA5vfTkk
eGWhaL1i4+bDNjHu1X7hhc5mNOH/KmYl5aY4mgfDSJB3k5MtLZYI9w8gVO1SK0xU/6IDsWIAhFbV
pZCR4mDL3zO2qXTOGeWOsFyQa1ASQM6DWwJs9AjOF3OHShHQb3ZZsfzQHNhOGiW0Ardyw3zwL619
84RTxuZV7wjF0dRf3s+mcObt3K5+LjDalEJH7R77lqMCr6Zdrpkut/TPkyuAuCG3hV4BXPYo+5uT
xWEEBgMiTlAz5jkQ5dFBHXOLafOO/fpHeA5VwTiY/quDC2kDcZQyng7KMIJzk3kjoulhJBViAlxP
Ug180dOZT8t0e4/Pe3vPhKqocXCEkZ1LydH9cNGq5qbB68iQd+CO8XimuFkrGwIkTf1YS6sFs82Y
JbKB/jn96Q7cmhudhRrcgAFXE2Am1OTodnFfE5scl2abzwAm2V/l5zCfy65ynXzUdZSIGyYz4Bx7
qZ0FQzz4AJzqReoZ50q+wYI66eWimfnN+DtVyyimmiv1Aks5VpNUuB2ZWK4U08N5KUyOfZ+UAjPr
iYNdK5V2m1SdhXWuR8zL6XAq6767fTyNwhJCEoO1byIxmN9Bdy9+tz/JWlYk7e7N1BDXIhMWEQHB
is0WUq9a5kDHJbPraYVvi1Zl77V8weyuYNfgUsS5HmfdMQyym9zahQV5MRnNynv3v79QOrW3Fwyl
7eI9y63wOLmZhjtRjfNDCQZ5bJUbzpX0hUwxPlEdORZyOtDye0VVUhK0tiDlg/3oDHpE6qV9Wz7L
01HBpb8szzc0kdtFk5dm7v/kxFrEWNQl+nqy0LWjVdL835zq6wsJX5vvdEItEoNYsb6JyVPGLrEB
QDOu8AO54y+hy/HT5xWpAWzSIbC6do/IjjFaKc6CLWdkCWml2nrUM2eV+4ZTq4IfTp83Kvs9cNmy
OlmV5Jz22J4DI0FzwyktgJjZS6BRVpcxRNbCfFgfzpCC4EMybk7Au3gLTjXUgN6Wf7wG0WvNWbKR
HOyluGJTzl0aqBZw/6k4NrYMeu/X25uV5Ao8R7W/adDVhNf8WxZlV0RHClmSOHBTKNA82lTKmQ9h
upya0fL/0R+0/des7JB66Q4hBQOqpUqV5I1XwYzmtCPHaiiM7/dqrizB9A8Nd/mp8qhelHoeP/ug
15ymAdc+3jT6HmDXUWGrfpDYLx0RjtfsPhs7hyjIhSXQebg/JxQaanhGnxA6bWrqT/KUYVBy0qhv
PUPL3/fUPlwrTlghWIvW3MrDcufPLT6FYUqkXW5NQOuV1WxXPPzzC47PFXs4Smg1x9NJvVbq5b55
Fj/rKBCSUqBs03a82qg9TO6IaWF4KQBUxvIYBtNwehzBp9LRTjYH8LmQvCLPKn6nv/ibnwvK9F3l
ErQd8J6iVhqDycVLlo43zRBNLz/z/gVIG4GxS5n8MCuGdzDl8rXDEBQ2mfAUhDED/AmZqIuVentq
slagOBXaAA4InYwWIR7BClKfH16yqhTSKDOX97pXaUbWi1M+sVmIN6dq/rSSaWUiyu7iARiQ+9Sk
ou9Zwb05UKuuy5//G8DZE/xx8zC+i1kpLZ4pZ5sfgLzI/U+mEfv4nGQJWE3+v5gA53X2Kp3FmBrX
+EYUq8H3YsIPUf3I4ErkH3eYVArtgoPuVuBm0Ce99eL52eJsjmX6sQjERxwNKUbHbwKMtU69ReeM
oimOkM1mquCIx45qoAsguTFIgrhqgjrmxGRqLd9jvX40HrAr2Sda7BM/1+SRvXUgnqfpvJRnhNCk
/GnVJxoTkAV3J7vQ6OBhIFOhqGA3/wc1fPGrzE0AND70JxjLQy6ZXTdzek6Pk95876Yb9Rd3Bw/k
L5+5YP846tLVGwzCq+NWU5c6boxoqUM+mNGUFC24A+Kz7xjYuuy/93iBcOGrzW96HCDdAF/DW+mR
h9paogKwvyYegY0DNxFu7D3jvhZigI3nJykvcTA7fTZMMcREA7qRTDpgK8JhGmiHVSE6NdpQ+Jk+
xrPKe/v3fgtga9caDhMdfNYyx065fhvpyF1JSCpo8h5fW+1Ozxjvhqnryag2/d+SGJ+maYplsFuk
Pjh7na0CZTCL9Lsap6cm2RvikXFPr46IGghrusRAIbq66m5Mo+i33SvOR6ivW7146NP1Yw5Bmps5
qQV0fe0NOqbpnEdSapfcPd4sv1ZixYzZqbhrtkMGJNDstsMujr196GY9F/5EhdXdOBCwTJsfJMEx
HGxcpAN9GTrEABUrdcNOJVlqS1Ddwcqz74FVE651BQIEytXR8ezOb+sRAn4OalcEX3L9oqpjQjUc
3ULvDY4xncCFwR13ZaF8DPOYsVvnrQxpvx+N/MpWOf5R6/jcl+aXB9dV8cTeSQrNwdOwx3J1vazN
PVcx9YxJiOahq+PI83I+c/g9ZuheOqtK+2lXuPzfkxfhc5QXiBM1xjxKqQnq6wxCb1wkJ0mWO0GJ
IfO8zfIAPRjmqM27oatiDs+2knbIP49NrbG8K6QtxDiQPRn1S/jFfS/enpoju18LLn7hpIV+e2GV
950pSmwsssOANf//5KhCpiBokANryAquR3uSqwtYIJMewmJXFDRCnmUVVOdoRUGpDLflNTC7KqiJ
2B3qs/tpCWaGRIcoUfLfJ+Kva2oZnGlykh0yCFj6QcJqOlLzSmVp5NdhPxDQ/ylFcYUHaD00q9fX
ZnXLoqiB9eHVaLlGHMs0H/u7uxECV+yNypwFT7csPHe0qKKZ8LLbP8wC7YAz4aLKijdZUbAcIbKm
cEqTAbcsFCdjR3n9brjwpCzGhh/YWchDXDayUNAK8BWBkvpjtxyEBxHH4zSddi8V712SkkFDJTkv
tW2aZ/Ge1W2/E14jfM2+FFz19YK2FNHcbw6xugDFtBGmrmOCqzskKWMR4dUXnLjh8FN9wMhaegGO
jzzn0dWLhmyq1C6H5M05q73DV11qPQp+yrRdyoeMukBejg7h4VisE4KWmgW7O4Wwc87vLt/j0HBc
CHxEx+Vj9vljpbx1x6ZFYBAhDBh5GdxWnj8ulta65VHEp/THZZSv7yRWuDOFcArzwaRPI+aFpRxy
LA2bt45/uQTDYPGZKBAlc5DohLBnZxOnf0WGvqGTzziHkdtvcE13bppAqUGbuGydSYvoWhYCIxYk
4s3hffh54DRALsBHmxREyqd43IjUjLepTYAaVhee0FxksSv1WbE0lRGDcGgyXGMnxYfgTPHA3oJN
9TGAsDnRH+zuhL4beHu/3gGDW5TldurqdwCD/Rj/RU4hs3c7/+QXRKU7mekyhHsfczKasfaBnrtm
htswMzk55OVubMBlLpzEit+hTNVi9ANYNkH0261LPdbXUPA8sa1E8cRwihlCPE8hcZQYdGw4gfPh
nUTtZPlV+uv3C0+gHBXjT42z1rTga6KbaPB3qMpJ8sdz73RAXY6Lqc2Gjvr9F+8FXt5WDqdW8Tiy
31nySN0a2W6CWUD1ozs3pX4ugMxytxxqUhVechWqOs0xARPHUTh0U79W8dut1Jz5gbyUMi9ftSxh
6feqT5azZhRlQDgesgQNurZbbNEK2hcsapJlMe7ISn2rJ+F0P/cMcBfOYoEfOyaAtzIeAQte4wXu
sk8CB298MydPULCF9ZtakVKu4AtCA04f+RqjSOtAm8xhIlqp1xfJAyj2ttj0RtkJVUse0qMm+myL
/WWCyR8mTs5WXLZz8sJrsHT9Jy+cIuSHLn9v9mjoVcZs7aEGM5Vq0nUVsx6FGkNIlZpBrOf4bkjn
Yf0sjqK8PnTLAMoOA2f/TofvMCwlvsktlom2MXpRvfco/SUACReVWgI3kVFoMgFbEY8iB48vAzLZ
uQYIbAQprn6F6P430bvMULBxku0Gg92hOZasGEN3KXoQ82MXEMHOZ96iS1mY0DfZretcrk/5PVXN
eRT1P6KzqE7XkpHiYjJe/LnQBhGT7oZDI15Yl6ZcA2k+OYIVcfegWlRI0GGmakPE7G/klluSt5Iq
1gPTXs3BjMwpREIW7Ura2m4SpNFAlqgB4dm6SNupu2/vzAlkNEAKiS/U5Kpc6SjXu/lxd1TgbfqG
XTh/PUvASOKAd9aJDdgHwwGGcyif07W3Dngs+2SMaphVJDz6PXRN2gyPFrJMPSU8riZnVE0dSdJ+
YQgfqyEsBP43uEnMZ7eju7ErItVCrbry1X2C2mJ2RhG+SmPNYLfAduB4ovZMCJhegXuIssiP6ysx
g5yLDYdMOwp8jOD+4XhfGiMdwEDphqn3jldPzeHnxNGfgcf7um4DLmlFBirkjmGF67pIbWKqKsln
51ieQQJxNt8dC1rfg44OO91cPZB53Z2XmBP2Q4NJEN4JQCjp0TlKA02Q5M0cozRBvgAqj7cmY5gQ
CAN5v1PYaconEZI+myYTxJVKZ/mSflOWoHKSYqrHMH/5Vxt0wF1TLjt2ph/Uw4k6RudialeZSmuO
zXGTy82P7758ZrWSxTTechn2sE25VKtN9cs7hAmRV7QTDKdhBAsSt+1CJh3ocKVyejFX8nkVlgF6
zxz3YtOfemBGVdbUgwJbogegWFY5hive4Rmik2jq50zxAJBiNU3A2dU07/PCgzJ7GJVMPl4og5c5
plUyAOihSWmhuCd9qOb7i3e2K2PKvpEBV9nokuD8zn0swTCKBtUemPLOPyC5iMqRE6NJ4tvGbjL3
PLA3Mkf9GrQsk7Sl/sd2WZylFhxIRwP060uL/qYVPXdCBWfB3DSQiQl5WG80vlViQ966lTS6gJrq
Kkx6W5QWWIN2BTcpSy/NM07UJn23B91aM35VqPLW/0rgSpz/pZ4SLCS8qb4kkPO5CiCxws/uOgcF
nus6cEPztS/Mbriy4PrVLNs+4zbHWNNiI30KTghHJK1s7/ddolVC3Cvorrd/dS+0ce/xYreKFP0x
DaVl1hMa9f+XQ+UyRdWw0MlHHj6jTcW6o+PRhOYQB1/ZXimlLgOMyvX+/b1ktKxAbXOZB2lTfJX2
nF9rrLzQb9tVPWQ83LMt18NqGbvfLva2Mla01svScUzvUocZrh6aGEz5nOj3eHHqeH48oyiiPQtB
4DDDZxL+ziF8uhTRoG1cgi0JzoSnG5RMdAMgA7r5yyAy4Cyr6AdLk4CY2zORRorm17+mlqBe/KhF
qFklSoBfizLquwLYEtaWiFiiUNT1c0EaLOtWAuAkesiQUU+9nRf0ae4lcCsThG3e97Eyew6StNV2
M2wB7003X3tlW2pZt5XLuZPVT0OF+lP51d8JVv54ZpoHn6xqjnQyyGS0txW7Q7UNMAQJLVel2GWH
lEk+Mi+8jkwja4ln3eR+lkMGw1j8b5ad3txHrMqJlE1gixbj5eO++9GudQCcLnecF9ilJwiqPDpB
0A/Z3gF3IacbTKsJ2vV4uleURjX0A9BbsEGZwscucJZluishvYHPkCun6z52Yfw8jh1W2HjFdsls
0GgnEGqz6Vjs5iD+DQCjY00deD1gXaJNM+joTKC0w394oPsgw9QFmg2zMjxQu/x1P9m90E10dy4k
cRiDEyaZ2ks45mxqTqK/rzUXdFyAphqZ+EFalK98EE/p3oU6JB6HSTeh3QDVKDVHQtasj2jnMIrt
7IrOZaJGeURyNelsNnLj1rXiCqOKQn1f2H9Z+s7Kac2uWTFZnZaiek0jbdRBRgMB/P9ww8MnZjU9
a6N4hrhcRz+tTaOjARWNpm+uNZpL/9rLlKLjOMUAsbM0mFBdR28yF1tRokaG7v2wlp71M//Mp6B4
4mct/KbK3oC6wO3rYyWC8NOXaUBEfoSKp0WzUjjYDHzHjbDYOlGkswCvDQEID1OoQov0YNdiZoY5
OJqWq2x0ZJxNJr0VUHJZh6JzLLS7YtAYXQ6m2HIVox3ca1mpomuKvJ0nTZMZl8XHPDwr0kiU6M9t
yO+L2l/Kf/UUHiyzPSx3rEY4DGkBRqLZgZlow8+DfiXfiYNhcqw/2DiVGRGTeUfQki0btr5ipDkU
eZPP/YsikBh5Ij10xT7WEXRJONMShdJHfpvBfM0y4NMufh13pkNvRmUBr0Z2BWWAMXk5HA5+QzVs
IjRAqq4BH0njLew0AIZ8ehDfKGftcq4k3MMvRuoLJHx9luB3EtaOEo2uMJlNEZoIWDOufuW/hS6C
hIJNyHk5XyrNMMCTW+84nVWew7P3wmvKIPYej3/Bvn7LX55d0Aw4PR2xBXSYwUmx9/JUkr3uEsDs
z1YELg6+ldaQwbcJRcqaHAUTWpfufZ1F8eolqp1X9TCted8nEbuvuQW7Ux8n1HQshcWaArDecs44
/cug3FhElNMw6pfEMYrHs82mkR+NDTrdbpo5f8KKP3Ao968kLLhVnzQKucC0Ty1JrKoIchvn8ZvY
CieIPFsBr126GSgpb7rifHnSg7h5NFrGmxHkSRtUmG5P3k+TBQRQ+TbuKaj1Vw+cjUBego8pfOaU
BYZDx9McTgPTpEhbZTmXFs5TCyXnYnqyRjvT0iFAnjP5quyBwuCmA9BL0MJ3YNfwuhYSnxPEceWg
+3FYhpft4rMcbh3SmwmlfRMZL2G3AP9CUJqlERd0hwqak0BK0m8ak9YBELCsMzrdE8eHCGFUOryO
nUQMW6zHjkU0bkua2QbmUJEsAAP0y1Fbou9iu7nJzzNS6duXcyXPtCr6OuwHoPpaEJRS0MQpfXK/
zkRtvUtVE49tLOiiPR0y9NZ5eDGmX5Uu+jptjGQIveb2dBGAO/u+ktS1EMYrQNXPrKj6CWuODtWh
sTIyh8EIIYnoHzzC7QN597FA2q5AfNwvNFjzIRmYNOCvXKCLb3LWfnxSK4cYSFoyLLrhUmT5vPgV
JCxKOVWCQcoi5ry80PCzTEDE/jRlKRpsh6hBU/OrmT8NWELPrKDHBYPbXpGzurH2D7lOaNMp/60c
f0/hDiXTCQcwjKXMfO6SorgMKCYPl+eWtTycCaU8Lyse7d9MJG9EdKwmu3nx3MLTfK+SIqC8JMxY
Inv2kGQFWO1ACBifTeMl/2/Bd2cUQ4g6RTrnMKeZMrhp3AY29TmcA4GN331PxSblMmvUEUh5s+do
pcEpzxyZkNoadBolM1rSUgBRJFa4eUrb029d2qpyL+a/yAHKMcaUDLijsP1YGaJZ+2Wnfsmkhdj/
WMgmvklnlr+FSQM/ae/iEU1lexVE0DZj6zIPXgOcS0P7DzPRVjYWvZWtXHGI+hXq2SlLGUxqo8V8
ox84thn8m4t0pIdVe+TbRUDMklms0B1JTjKdbgeKrvT/445jxY8f9yk8HffRMQCyVaZtmFOaW303
K3no2FQ1sJcMyOwezjqbXPZA2C1yDi3sEFZOqKoeXMz5fA1ZPcLAiCkRPc2MES+sKIPQZJGBhAYO
Id6/7DydjjfihZIEwtHongl80isVuH1QlwTpvb4XYkzUIY/0JMeHMggK0qfhMfvpXX0RuYdVvrPn
IeOyR5cl8r0s00SQDBJ97XW/mB3R//Lk9Z7idCfd6sVWLlAemCy/eHqpSekVoDimJCxlC+tr1YZI
riTO1xdbTeuetMq1wVCY3rvC+2v1JKThmguhxTEUiHUtppZYn5jJW6l9JHi93xve9LWrl/QfIpN9
3EnTCKr3pSNi47lrqdnIj9bMopwU8Vvhyc+hYq5G1jR/TvnsYod2j8LsfkeUsTa36dmc2O94AFGB
PtBxivdf5r9Uxb7uf2tLiUYFejFzugZ/+i66ft3iVVKCioX4sQfFlb9woeWGaCLwCM4wtgAC/lVJ
O0bPkvwx+eukc3DKfz2nF7bnSnD37H308ZSEKibokDh5QQppv1NycpK0vywKTxQr7G/5Tuh4zHtQ
kFIDbG31TZ9dTnm8vU40XUKJrDFjkgpOxdvqOOeCsxYtICM32NMuNZhuqAl5sKkc3Z7NETXp/W4x
0fKB3++PSqwVFBiEqCvzU6muV+p1xqGe3KYfUNz+KJvFAxruBJPf+ZMPxjs1Dfydu7fP5lhJIsEn
+/t1+p1XwXtV242SiOxFMlxb1nfEk89qSkfplJmVjP9H2uvHVpQzHRxUWUDnHvigtm0Po0DiIsLw
xjdJFcq3dh+ewYVR/3QWhVor2AD7edbgNQYrJmBrN1EKoqTdHCBAhgSKYJO/jb+ORf4cOyANIKDA
zQjcpVgIu5VYHyXEpgKKR25Yc48KFMRNVEeRrv8Q8P30BMlgNjlLgUS1O/nzkDoZAthBXZISE8c3
/OQHOviNX7V6ug1NLZpZBy8JK1g+Ilv7s5vaaWIPS56jBlqBuizFEZqfgtcI1bmQ1oS990ytmm5P
FOCInbrPHRrCFM4mxhwuNemJs8KL3aMkXU3O6dYn6N/55h/jl1Vrzt6Q/LwZFffNdDPL+pP8Bzlc
r6s+EhKFXX+sFLmKZu0Cs9AQdAGsM5jer55w+G68tpx+vnUTuyCs/zjTZ6CGf3qU+VMvqw58ruGW
aXpmSp0W7PbA9ALBoVYp2cvQRyJXo0QpkaItYIfBC70ffraLIACbsaV1BOFKuL2JpwAx/P2HM2J5
QA58R1AwdOrqlhNA5SvjgA0hBvMk91N7UtVWmVLd1xDvlAzPaFw6+Eiruw221BNlfOH+VWqVm9LP
5ltZM8RmkBLX1v2d4nHsLji4pAPg46IFzsdtiwOSKMNNmviFDlzkPuUQhoe4M9WliJl1Ns1Ss5JT
FTcsWCViUH4NfDBsY/aPZ+qyTnmxhdagXd0b8xIIVRbX9jOUALIFW7gpFanpnIwbKCoHxp46UDpV
Izu8KqQPqtfAP2jsvZ/qjS6mYcDzv3g6crEMqUU1QCxFJB46s90ngc5I5C/tYhd6fOtSSVKRY8jC
y+CZK/YMAWlKD7d0h/JAJNxpQwXd+h2qrlhmaC1QroPHhvebVADBT6SlLz6orxRBmHwt+UriPd4B
N2Ev14EKTkcfLm6Hs7EuO/vKnShGM/xT4ZIjIgFoBCP3mudslG4NZ0MqxiZOs/kLs+rWNWRwg5Wz
zvXH/pWSTB0uYaO/y8bOmwuAtNs4EtO2ggfPZZ5gaWkNTbL2gwP6zzYCn6w82FnrAR3rI0CmDuGr
0LZtqAtZnjq8KKqhcFi2XMygaRBnVEyeYSE8sP0H8arPs612l9+HNZc37QXueKf72e/QBUOxU9b3
g7LzNIp24J59S4qYtqS+1vSOnsW3NuuFIGiK9iS+Anifb6Xlo8MB/6XCHRjYqjcNVggZ6fyz87iA
ZtV91GkQIlPD9vX68UJehHudaeH3mX8FCeGGKC/q8SAbCtQ3ByQ1GQOOBg2ha1324UnnpsWQDIrU
8AB15KOUYZR8qWNG338uo1BU8Gf6O7NoL8rX7iM3zXLr0W2Ph1/2D1VhVEXZODbDrabZZl85T+NS
dKGqyi+lmSj/AnqXhMn3XXi5iJWM786NfPVHvcx736a85BrK4zCk5kyl1c/2vFQ1nGtWhWI4pFAI
RlQFbjX8+q4VY9onm5KoGLFEAkj/FDiWfVxCD2ggkV4xqZFH2Jdn266T9P/7dsxdMSHu4hdzU9qc
H16ROJKXZX9647uT9kec5JRi5BTAevytF9+OovRuLlPD2EIMkE6eXDYh3D9vmWiJ2JTlzQlV2OJr
nFwKfQNS9BtFTMT/lnL0GQM23arW8aCazOrEFf49z1bHpEtXvNHoGCg2q85lAMRTiUWlLKTKczo4
1g92TKKdJ/UQdnnPhTkXyaJSWq3kNQnmbeTlCv56O2RnOjusjVqpMwunoVndm9SiM6qx7eEkXzjW
7y8xMFpdrXvZJ0whmp7LMwTtsFIFkyF5U9bGYsXunJMCoreAffRyTfxLMZfA3F12eWF9a0v/bJ4R
LwansfsTqzg/SDLYtmrpOyBI7SVHC9SO6VxZl3AqDBW/ySnV8w/pt+OX/4/36b67bQPl15vIo+ZM
fEwXVxqOiJ80MAWf+Ud13L00uLpmfc9mFjBZhIWyzHbPtIROyq1eC3nVhU4tGuzt3w08ygTUwVfG
7iwe3nrrRgVmXjzualYTOHt9S9gsCpjH2zBA1X815bKAJMVZU3MEEXNvdJQPdBwrYXueqWVhbdnY
cErFUs0h+L9VLWAA/R8hNqodkhXz0roSqIcWEfs/a5lel5QIFoxjTG1hg6fDrrLoKot/YEUiK0MC
KnzzPQbCIZSQsT4PUuOwAXSR2jOPM53tyG8KTigIcMgeRZAn0vlpCI5448HXpUXZ2kYiXn8rur+5
JqCLInqb6tj+/WLWwHgkh15Iugkogx1xpyNbAURRfIGSYKDoBXSi4qdWHCvi5jHQKlq0sh6rpIdu
PO0mFyNwKu6NH55gV2yBO4ryTnQJ7uRHhtEfGXGNtgraABbg0WmtahhhvDZfXK7rOcWY1Y6Jf7Vi
m3pUNtfY+WSGuKsh6B6IzdrN0bBtTz9Uae3zuT1o2ftfHbnSdZ6k/isni1sl3umCLKjhyoemuuP+
SFvAB9VsQZnBCvvaBrkP7XpjRb5gdaF+cEQ6rzBIg5CqmT4WfX+CjSJ2URVeAPnKBvRgDNvccYFo
uSXgOT7fHEZxUbehQn2P9PNpdSj+MXUYm6dpBbVXE0QkmyYAcbZHzoyhFTSaOwD+pSg7jWQeLt3D
fT7JjAoahY4Qdo1ZVAVwrU1Au3m6AgBOdB9b2qlcG9Its+hTtG4Oe9QskZiQeDFQhwNPhaSRWLHK
APWsMisiL/iz6aHW988Mc2/jW/5WdrOjYeTBTfgH7lQFoEKPD/RVX/FG5o2DaCNuXdgSAFv2PNJE
Iqefc1Ih+POvuWmr+JG+s3w1AcJi2bUSghpCN3Z2rCVRyl1/r0qSrJUhJ3RAbEdEdXtkwuI1cmHf
mZQqry/4QS1B3HsAueaR5R8Oc7YnoQOOxJB0VekSckppE/REIlfYdM/iG++fgIV4T2Wuvu7sWVHx
08C2B+odYXyefED45Rlp3v6XPU8NJwyfguR4V/mS6r9TkX7Kwfqk46HaCynToNgE5Zm4rIqzU8BR
PJdkYM74V6+iCrld0KuEmy6WN5Hmyvu5dC5+BpT5obOxjfp6U7Urejy83zozL5eoeDb8Ll+83pDl
Xc52hZCnPOXU7aQlJ+ooZE6LSoLraOvZLHkPBBk9EwssfrSCp4Uhx9SCSgta+gKl0hVxofqB6gUQ
2RxHlHt2/AhS/rvzPxyVCfkphmBNRTU9o3+SgywYYX90f0NsVdyoBA4X6pDk5u6OI3j3UN6hNrDi
RE/6Z8owa2/8cL2AClHHWM1/7AJEhYW3CVo+VcgUgNZFDOvART0SzGc2KofA+u35mjBDxMeTZTV5
NZn+rTY5wKIELhW/f4dz9W+InwEzwXgyTsH34THJRe74YoSrKjIG8r1O7fBFEiRSRkFlC5GGXlIb
kRzjHUmX1nUj6QqDmzHXUkcIAdJ0pNjt/RIFzNOO+BhydnPtEWYgGXUn3WHM03r8GhSq1hYNOAQ+
NTeJ6B6Fn1bP6IVkh53WmbcTeE5368F6P51YYfaIBEVGMjf2y344rhXpV8KFzNde+oc4TH/m/vrN
6dv7mbWfsA9Lhzph2OxHwDinyJD3UIFtVmOPUSsriC14SRdXtrdgEl+tLDt9LLz7TCaJ3VVdglmZ
K1IlAonE+g03f+sMcDS3BL/ol0I8+Vrbu6jiwtDpypxT+eGZt1+DSNcNsJATCV+qbDSS/0JTIj4k
NYWDXqhHfHRGdQNZyJcbbDWi23QJvVJ7TmBPAcPD7Ct2HLBOs/5Cz4htOB48pIkmglFeqcm58Y6o
7acSI2bQJKZoaEKtoRq5ZtwoqhHpuWIieQSDssDPT3c2cK8+/wPkzBDxPFkFnk7r6DSiP0/uFjS/
QOs59uD1FhLi5DXG6+bGv4VncG4VnnoVKu7scL2T7Li+iS1BrHqWmeIfFAkt5bOartdt5jvF4Col
6hlPC0NhLg+rXqf0cex/FvnQpE5BoE+PI1f99V0udCKIakuOTAB06Fam9K5IP3kq8UPAWOVjT2dp
xKAuvBMQM9luttv9Tg7zsvfY1f76AzK/yqhp2gMPTpwZUkfTVSjtEHnlbF3+lOH+vpHoLWjn0/Kp
otxrz9Q61p7MnrDXzOhmJfnEV9dw5ZT4bR1RiHpMeomxnG+ecUvPpsMN366UkYXnzqvDSJkFOnjf
zgVsCya2Y+RbCTShchyg/QBv+22OPcTNMcp7tTXi2CqGZuqCC0092zY0UthAGbdcFNhN19ZHgCaI
xk6fjRkZVSFlLTNp2PvLUkt2bO+HHrnP6Z8CARThc9PwxUzgVWywys9RHuGbw7sNFI/rgC02OYPE
Py/rQWiLMmc6rc3ofU1B6XAEpdISaXQdXa+RPIoLe7mT4pGY1152b26OtTo3rg4Cf++3IE4ZNlXs
vHDhExkGbDI7INIU5km+DyIys4EMnIZ+Ei0DKVtgKlbB/Xi5lFqVyl5247y0Zpjqm9/iMy++KNQ9
ci9x5JLpv7F5DmesloJ7Ar0BSFpyhtXHCgoX9A79XLAz02LKsQNLdaFCNfRfl8Prw/LhRy8XYnuw
ZU1/vLK+cXr2S+MiQSN3gqF7qn3yUXvfQff0qwjo1FFyjYb85oyVfRuoazhk9y65dBfNoydxLfki
SeaP2EIGTmRoEh+G/0ogucbV4WECLqnBDiClytoSZY+l4rQtyj+Ls0AoWum8oRzZ6XoG4kVrFILi
Ufyklhiffwvp9r9ZrXE0uWALsa1KM+OKdZ6SQ6TbmDqtR6zwUvDczf3j3RsPcxYw5nQlKsJ4RJVo
qxjkpZqPqsBGsfjzKAHJGeSw59Ho58ipR+WwXpuUwNtsWWVJ7dZhT5isrsJg8BTEye/8Zpq5FJgb
mvJf53GDEX5tnAc2C2RulL9LQ+oRbiefTIcM7p25K8f0DqkaAu1uGZgbEuXevoBVTReaAEP1Kesa
4bFtrBkfGjf3pvzy/GVZMWOhGrb+uCoEvWKFq3Khavarfq66j5todXHpkxisMya+kozVdet6OdbW
ywIufwuSeCCSETITMeW0LbZoGEn88278nkEVtagDCpBOH7zIC2OTIoPDUWJ0V1ks+SzypPVQyMMo
8NyiSncLoX4uALvokWAYFUX0vUXiU4+1+g4uXn/RVWzXG7r9jeAWvyDSzduNQ2uYIwuAQStQfKWe
Ej9pY0OBlL0YcTxCdEBvCRDfPQgODrofTiyGdsvCXx9uJ303Uwv6zbinifme+2hwYVb1SC+u/w8S
sjIDygbOlJjQqNpkvaxm9sst3mLCn+/sVgzi9eZXU8Cu6E8oa6QA3ld19vDwYmV/tFAjVEG9CyS9
rTBiSHtBCEMtcf4QIB4AJlCsQPMAcoFAYuLfcAYyVCxXVq47IMVz+azQ7NbMyplRaflwRESzUnDe
RgQdZ4Dpo2E9hC1Hihfp9b/+YZ8nMAMVQm0AGLUXmkshRWeT1ikobFZF1RzF06vX0sY42/rfBC+d
sl5Ku4Es83dZrfiOoGKhyT98r0FcDy/yh8fIaR/l+iaTwvUBUFD78otm9sPBNT0/LILMB9quq2Zb
ukHiOMl8bFO+iD8ioIb3KT1Ikqv/bpXnkpnU9rxx6MgvdEhWjszJZSt9hpokWbNvWGfAXiPct8Cz
EQqjaespjr9NlibyfdkD9EortPvT3ysr2++LwOBx0obNPTirxnjlkT0PmSchcLcf8vOHWkXQpj2v
JfFImRBiRNq5IY63Hryu5JfOCCd7CngrtD8phBEVjCnBTnSJDEIR4tA7PUMTmP18dGirE+bfEmA8
d+KJB6AoHDGSkHhx1IPm9Mwncrvrq/57DS8XmdZuP3P0kpoWlxkiqMcwO/Gn7TS9kaXEhYYXBnNM
Fvygp0w0VLdOkP9JQYUZNA8EmYe54uBJ/ggC9KbQj0uz6iZCsYdV4NZzN5cO7QWhAkWZ+nQxzQeg
lrplq/hv4mznACYFo0s0WKq78Xb7m6mX8KnzUX36F4XOJ/Q88GkC5F+xA+Re87yfrhtPI1WpK6Dz
HljeAtbqbEXyj9JDOnVxKwOYiIPAMiVf16F8ncx94xwwoDEgL+0brbCEQu9e0P5lVAuqNm2TwOiK
RWV+qNqDEfWPkiN3JF3yWgNPCP4g2oj/nTSKQ5FNcqkwuGsXvxg8eyYzkCbU5OpkhnDPfZn9ddRc
PJBFWra1VR4UrrBIZJFrqmXCbDEfbfyONT+PYyneXjkCEvOqBfo5GOi6dvFF6Zw0hanh2wwVdXyd
0RIz63SHf+dfKut/AyTVQEDVLquCq28nDeSza085A2TECv3Lz8GV1UwzJQdGOQBdaBiSk0SVqAha
uv7uSUmWJX4OBzE2y3Crje83WVbtyxc3W+AMkIdM2yqgKEcqJFRzCVTHA31SmGuH8Tr6pL7Wo9Zq
NAgWRxbX+fXZXa+QHGwEolO9wy5KN/RM9sMyjBRDz/JHIrzZlcQ7aFHDMBgROnRf1uKWcyjwUebv
rdJiVK8cK1IfrFfdLlC1tdOrHwzN6fdItMjKkmB+fjNadLvvrIQJOydZYF4aMRuMLeYeVC9sq2/T
r+9ZNmGvLg4PY10B5OiGfO+Bpl4UgNLeYJUcXbu1PhIgwEPzAkMjMu4/KYC+M+2GJZwpTZVjAFoO
xS4Yl8j1paIw9Txo93e9FQJxM2kU8oJ7+LTI67SnKNxplkiM1fOO03zN9lh0ZbjEchfq+bQFI9QY
h2aTaI9R+3/H8qTSTJFe4HAfex+eM0LetjXDJE7IYDUXFAnQyMynwx0jvk/rmNuTLYpD09BPC/1T
bI7RIQhqms/xCjCk1Kh7STXMUhAu0T6MkCZhQ6zeuducMWkjKi5JLT083Vk1vbVzDwlEsGRoW37O
o/BAcpZ+LKIsKwrlfmAF64B7UPvmXzFR6l1wu8pBAEpdkypoyase1OLa2dgIQYlJJGgwhXVanOVL
bf9m1bSLM0hey66Z75807x46ir9rS6R4IGYuxu4VJpW6tFlDeOSj238+eQDHOQok3kaIwZRUpRbM
roaBRpXBAdplfx4OUhdqOdIEahl5llKkPpOoAi8pnwhxUKatq7BvNud9BX29qpkoe4YptaYC7kRA
+zC3IxFoHdmIi/MAYCbSNsXN7By6SkFox5FBh5OcEW0AV5Mvf4HdBajlG0qYmxqQMqk6MsDib00f
+PuYdWtvpBbQj5prZnbx6m9usX6p+1WKOL80OjW4glWCkwSC9FdCx5I46SiFsrpfI95i6K3g1dFC
jHco65YYH9rMgCGiOAQacAFijRc0+Moekx39ZhdqzfWqB0CwKfNa3aGYawPqf+fP+Htu3O/AMKaq
bLIBbWo/6sRqvE8l1Lh+d4lsNqp0R8+wV8gO2hwSdfzs2tX5Q2m/5CIglQwjTIedhDVz+58/hQ82
lA7b5YTsSXyuEIaNC448YT3tsQPvGJ8etI037jHW92C1lxkPgxx5isR7q6X1wr3S79eV636TvfLv
17Wk9yc1WlfZK2oN0GAa+kRvLIT6lNVV30sAIiozvA0SQvFmcskZA6e5jWDmW7xCIyvSqDr8dlFa
QXU3eDcXo/0DmQeQvPUzPRnNc32XmT7WxI3uHASL4bO2YBUXFjzTTjZsfeYzap9qhLymlUJTbmVH
IA3kjdMwvI1C9YVD7GlwbpFbNayaZutS2jCCZx0xuhEVovDibdbiVvrLZYG5h9t7rNiMCOIL0WKE
Vyl9p/m8emVi2DukP+y9pmmaN/rHCn1tf7I7bkUYxl5RyeMDY5g5Pc9iQRRh4DK+EPequ6WEk2QV
B3lAafN24KCa276p/ZVyjine213MRjPr1uzsCG3+y0WCGTfpEWjIgi+o3klX9DK9bgiaYoRw1yGk
h2EpEmr0EE0l6BLAYAL2Gy8XI47ALawrLRFVPue9/GHQvTKX3EUPbaGH8cSOqwEQieuMtXLHm2Pk
s2z2b0d6SGYKV+yCtZqPgdjkqigx3WkYhdzDmj0oTPkF3i38TUuII5sCWa2Q8UEhQ7h82N/9vG4E
+3JOPSXSbEqTrHv7Htla6ST6Ge2GPHHWWEyTmr2yr8y3RFKES7T2Oq9ykalLym73w/n2zK2L+r1Z
/gFUPU/Cy5n4uEiZSrjR4cmQobOum2OvUfp1Vt0CfOR8i14133mbjjiWHf1C62fRHpCnitP6iXQB
BZTDz5n8WJgEPAJHB/CPvIJN+Pigpngyt02ePQJe97pu8wspkF9xIupOy8X0Eu2MGQiL8d3pJP4g
DGp69NExdB7V4verUnrkeJiG+yxWOI2Hr9TFswWVYQvfqLJtVTspnqUV3JGPpiV3Yz00Cd1/VaDd
Zn2qfTVQTw9tkv8nQA/a2KB0aU07PfwfC7cse7ZhUxyJHDMctyf+D6IhaXIdrp/PYjmZChbaElf9
OZvnSwhOoGQAtn9/hfADywZyV/VNYKljLl3bCU4r1U4Lh8Te5kPqSRyyIIJZrxpXes8cQWxZHaJ3
prtuqePVi56WqXYOuvgSlxLC7kKy6WMFcxNUdiGwMsg76Eh4hRTS+lJlm22E1wlA5a9inz42T668
FVITfsp9Yi2cHuKxZvjS8+WJNKrncVqeNITBercZbBMewaTBD8Z+3VV4ZqxlRKThLE2+qFEJTMGP
XJ56En/NsGVO9YtT91tjOX213G3QSc4Sc8C76JpKfITHQffZ23jbd0OuGwI0jHJbJqzt+5x+A+5c
t5LAtPb+xEcgV9mPaDeIl9riQyAmAbGMx2NHtHjEqngdUblGSDIjKnFnlyMvvsPf+0UajwZYEmd0
yFkEEUCexjlECJTSe0hWZF3zKiH8sS5Eg3mVcDvl4pFdo6Ez0tlir2gVRbLv7aTr0lnpSZoi87AT
lm/netTO8HUdp7UFbQkTYUN562ohCDKj1BvYQY0DyaCMPJZCAGSkqC5YPx2v7Ov8Nfxfj7Vyi0MU
pDtUdgWETaauA5jNTMinbTB7zVSSZEdTEERP7L6faUrlgDRkMI4vHPBP6PGrwQbsiTvPulvCE5Cb
hRcMRftJmk+BZD5Dmig1yOE1GXWYnynfzJ8NowytBaHtZPm7uJ6cSAhnAHJjN7zbsAiQtOhMVKRY
pHk9csoKczbA5oX/4/RqrQPzPhz9l+BvBj4uGHpeZWrEvpiVmuTczoPJaEU8w7+KJwfVYtiGh68q
5PPR6gj6xLq2Orw5qHNUqV3LqpVRmqj07kT4gRfTmhDwS3N/pUTLK7H7FSb8mm783/r45LTQ5uZI
lzIxenw+bhXj40IF+rNlShSty5Hmc6U9kD8/w8+668EQgHSx2ToXXGnuJMHh/fpFT7022mWoyNwR
gL2tu8IbsEiCLana30FcNDFZN2pLifdFM8s82HD6s2eVNKfdMGPpZ8bqhJj7U8yiz20hN8OI2S/f
rVeUaoAgAlbpaKJopZkUYTi2RI48dd0c8bT+ScRu90X4QM+fEMUgEP78bwpE5amigQXsnk/ym6Zv
reYaYiDOGpsyEUyuWojvjPLipnATDCgaqSmJHv2Ga9E5bz+qi97lkfbj/d0F1lDZNSShfkdocbAy
nXYv4favLUBWeCwMEb+rndjQek58odnR3SevhJdPWLWZDxMgr6nrNkLhW14QhPImcKojS8VrJH+8
E/Ij4ShYfeVp4DpLbK3nrwqhN2OJVmHguydTa9xgwtAGWXsDheX/xFFl6NToFlKp0Q6HvCh4hKOr
sXnYPcM5eCDlCBJkdTNcHCYOwY87VB4F3k4KwVxqjfM64djMUZsV6Jt0U9CwYoQ2a4axeuOdZSo8
F2iAFTDnyrgKA9SYP/7nx4P4k20p3RNCGqwf3dbaUb6DqF5ePGK04EtHwdqUZYfhNkGPQDfW4pNa
ZLbItrz3qKudQ74W0rsU/4f1KQsnNtA8sZ/0v/VI0myU1b0SqHkbxQyadpr53+yO0BUH98hGG+kv
3ncB5k+y5I1Lv0VB8mdMHdaVS/1RT5MksAwITLYsAsbuyTufUJFOuwc02OhI9RMn++JsAXHEcwVY
nw9sZ7xUtn+Xd5bXDIE8DfSys5XR8SQlu5UGo7RyGA6hH7oHRXGSasWE0vOaSgxba2NkoJZT3woJ
RhP2vyzffY7LvjqPZm0fms4VeklarOXPv+7VNJbY3wkRS4ifSLU0SumGecCYUwJ7rIxbT5nM3OSE
BtDWQVodNJVE6R9y5zFgveyOekf+cfc9a70dIdtOq2wH3w1t3VddYv606dqQzGjyxBoW5hjfDBTu
dPWtZHhRwekhyaz1uWSj6sOiXjOyGKqUWE3tr9PyKQjCTGE50SxVI/P925dtR66B2MFIvEeAM56w
ccIFP+VSC7qRtmhASNGnk7PJ4TpqK872iWRGwP9y98KcX6FOKE73siBXv/IbsozHagY1byikalf8
SyzJ80V2zXdgRmPRTImgqwaod4JZV/oU0QOCK46toA0VJ+0lHIIrIMeOI+wfnRQFvbDJnIyw+LxN
Y0DBEE0T+z92STRZ2ppvKFYdBWXsNpp+oVTLXpSPe0jFdpdFw0UkoIDG784f9xiXbl5ENdfZyPHO
bD71kMqgLuu/bFBHVTuN7Lkydk74O1w/5BsSrNrbO/q0lIKE+Qua0ADd3UDZNA+tAuWpIGbfz1Km
F9Z58mZxWxgkt59fgAxEqP2my+Cf2XV6GLcBe+hDJNRGLXx9qWQHgbY/6EzeKIuBjNSbmFT7Dezd
0DEPOes9x2+2hHhaJPi3QzWJUnAI8bInPDfW5wV0s/e5yQzAaKWVubB+GD1ZqNOsBhDIo41mVucv
xxOE43KiMJx4s5SqhIAjOfXhPdcYdco1l95bAsFp3Ng4pD/DSZCdMN0fSodYiaVCSJwQWLYD7263
6UFrFE3hApprqWyPs9fEBsOnaA6Lip6b055vmDK7EMbhPKsLf4+yH7XNgM60keCoIdqcwBJMHjNj
arRcgMBEHZa73D2Bqzxdtz+zyrbRYCNgpSuIWaH7piO5fs4wpZCDgdou0ExaWTgl+q0HPEbDOKxI
RpiynKOi+HWN5zPgbI/M+XwC6alt6OEz97TVxR1ERsptPHSoNjuwSFZvVHNMRkqwXdUTbSFVDs/k
tYykPEYcVBGTysGlOJFKHg8BIa3jRyg7nTgeT52CHA6JA8oboiJ0YZq837ZazbVXq5t4EbPiSzLh
+Nz8DHzWMFEWqwyxV/Nw3Zr57HAJFS4VjrNQNNTKwI2Enht9dExIFsIEPsCqDVIv0+O7yLakLHWh
fdaGXdO+hE9mJigRXZlmACHm6qBV6gq/LCLk27Tsb2YWLcFi+uGyZL5ARot9XgI11IFns3Pc8jnU
YiDAyAvuL7590uAFsVikGFO2eHv6zJeIFORnfgygrr4j43ppgZkeCAUcPnR0IFINTMmysEp6CziS
oDuMS5cQ70zRM+PzlN0d5MBINrNM71Z+HfwyyM/8rLDnREfZerDpNLFSUofc3OJ+5mCAbv8b+i7x
psKc40q5/C1whpHICGUeSVueB18SW0BVYAP/ZAsTcEnCvZwcykD53LwBVCBZ2oBLGfHkcsPc/xxk
Hr6h+DRvk7pzpmE98fB5HeTbUx9M5BEZHIOuQf7T6uXT0D1+SpI2YYMUMD+TlKArbfYpYS9bzhG8
Qb4gKzmRoLUQRwsOditsiU4TAyl6oJZBVvHWCb1DYCXtHCBinsjj6pofJjjj+1+VLZWger2iEoD8
Eajqv2nsvvmw5ZNMyhK/+2rCMQQYYGOouZFOBDRx917YT/PD3Q6Cg7UxZ3fiyxPLFeyUjhjr90mY
0V6JBQRZ3gFh2uN4BfjoGbP28H8bvI7GqJ+0GlrUSfJlklIcS7fCHCO6+LKLIloqQFjtF53t2T6Y
VE9i/TA5s671ajJB7Zl5s4QbgxWcumDm14U2gluYsW+5jUP8KfQVdkeAj48/iud5h5LIL0JPaVs9
0YSn9q/M5nk/tqZuJVjdgD9PDTXP9XejteDY6wNL1IPHIGoyPLXa68956NITji0K1WhrrXdgRZN1
S4YlYrvOBaxe0g25a7R3OYZGDS8C7ez1AEIjWGV1uxIto5P9feH0QDqhilkJbCiR084dy6bGE2x8
7/G07cGcwbLMixtSGL/FgRr7LNpds3SvKqNQhPv0IR8ewfdFoiaThm1wz1Blk5u13BECjI+YkU3Y
eVmtHMBxUjWyhiGG6Ng548yleB5zvC5KQWnQRsPvjyRs2pQKk49saLWes759W8ZCmGWkB/jYR8cb
F9bPUnFrNBgZoq1qMYU4JolxwfE+7miXGrKitUjGCWlgqPhi7oP458a9Rax5bsrfLjFfQPlsI9vv
7n1JK8xoAf/G3SDp/ha1j7lp81TGJ7eie+4f3XNuIw+qhuvuy8wGBCyGHGTfvazlECFLcL2vlwgF
ZIHI3LtP9KELktzoQJR8BHQpPl2MvOgBRHp6bQfAc2ts7keBPPMrDO0ymBVItE7W/p1+Cn52Kpw5
iTdwW+PIyumK0Z6E7AYvYKsBI7Zu5YgwOYOzIjY7flUWTT0nGHh8oeogtScCphapA6QJStOxOM1s
B8Zw1o99+yqu4CsV4jhqYLf9S/Kh2W1zlgfvmNt5S3jelSyX1zM+Qx4/m9Y0I/oNhyvRm5RCQ2qR
dhWSD/HH4rENuYj2DkUD5/LHLC6rZ0Qqt2+J6hA3qIfx5aAe3cD84wkuEwqa/Tjwq0E8peTAwFg6
7gEMpiJhx2DSBrtX1pPBoZCbBlGPGqPC/t4grxVS3IcmFIVnmfUX/jEYvSAXp9W0yP8uAVOL8yLs
TjmJjRRRmNmh3q/BI3VyPCManGAztU6Hupz8zeta5zkh3hR31FLDpsVvtNf+F/0jp5MO+XVbR/dP
n97L2fvA+mWBovrOk2jmk+DbD8w9qd9GfUPwb5yOULzzFsqvV1j75uQ3iBL/bjDn+tF7hZYLnUHU
PFLmRdG1eB/83+NTHMUaKLbFI57GUPywULx00eFiSP0FUdT3AEfZg4+Tg9Ujmdq7aqvx2bexxGqR
NTEsWR9WRZKxybW6UzrviPVCuBfYXfaomQN+UZJHQvQJCB3ZNxen1jZp+VXW02lL9hLgHvNVgCQe
pk5ox0kQFgIhsqTwTixytTEUUq7nvcvA/D9AysnfOJeXitfqfiEfDs22yyCud3wZyliGXpOjzImJ
/sZY6n9poxu03tqvLdMnUEtbP9lEjphvNyw7Qn+2HL41r4sSjC8Qtg==
`protect end_protected
