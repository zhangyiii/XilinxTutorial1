`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13296)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMK/PgSU3QY91fBkoay9fSdIXCM
AO2YSxjwjCCa4kjZ6EHPcdcS91g4JnxrIce+wgiy+F0yDfCFR/l8LEMbQwShR1f5tCcIuBN2aiNX
9l+q3c70+3q2FvtIEUa0HWEALsMfo6LD6XZJIo01CpXkNpwtyDuMqy/hcKpknHBK+8rgD73eQpXH
5BAoRkpyEqTGn9FB02+clZaxy3DoGHjao3tsf/lYshWoubzLglfjCdH5TjbiT9CWdIgVQa/00KlA
gh/vwF9lEo+2Oj+zF20VQBDrLjGo+YAfsS3Svfo33npzYApZCJDPgrX4OgJsd2ozLiJuOQsOt1yU
1vUbUdfJp8BgAF7R4uOmbvbDgC6rDggGqb5bo06QP7OuQ9rxtgbnFUpjlKigefmn4jEvUrWIbCGu
y0r3+decpKJrew2EQlEDxpF+WjqZgaT21hFCg5AAUkt+GSDNCBNC1TFjS8oGgHMcr/HaR2hvo8vC
c7U8d0QMsNgbua0Xr59MLohp2JM+u073vgX4+6ANOxM7FyXSgPzklkFRF8B3eu37p5gN/FNFxaDL
5DjSpKYzRPf4psYmePTIpCDXa4vyX1WXj/cqRNB40AUG637ttbLHB9OF7YUFnpOMnGlMxrexN7t3
k9+SFCmr0YirfiNK2/QygLxkYuj/gaggpABGZI9sZXT/eomJphYxGCSqqzCpJBRQFvwi8lovV/up
+O6hsu5BNelPbTTp+46l9Vu9Y3AJ5QBEWqqt5v4K4D4rOFSz6VjAZ0BNiWR2sYHTRLeCDy+O697u
9439qttpvyG2jf0Zq2Wblh9p/x2PdV4f1x8oZmJdEXURVGOPxgtt+2dDfus69U0pIoNOtV/jrtlf
ZAGk8QqRiXNUjglFclDpbS0uTYCkCUFM8i3cvSw6LdlNWFAPyrOnsCTYbQ5/sziisLMXgb+hUPs0
e7I2G6hYqmHWAs6kQJAHjhAPL8XS6qshQDXl6UQdaksK96cgGQM6vW/6+1MxUiHbbHAfYlBqi9SQ
pzwBz/PB/14XrLHQ8nepNkrXZqES35h1Fws8YAYlg/mtRmSX9ugat7nU1yZ6X018wruFuSxmD8Pe
W+Uemnu8P9QKjO99gNLKgQP5553OAqJRzOrlXjnougiA9NxkUYN/ljuBOt8C+E9JgLkAI4MdTM32
Yt7Wd13fRv/SK0U9Xo7tTN7yYUB9DmikYkyZbmL+MhaOQHyp93sFZBpxxeGVS8JFT4NuK3DA7HNh
+lS+0WvMko6CfMAXQWv979u+CFFbCO+Ad3ELlVDt0SIF8vwGd0oVJSTdmDBDDehvwVqYhyKftJAd
uRHcS9a7eCcUtY3d0LK1SE9H6vpCRccsdiy4WeRP9B/IhisGq6PwcCvFRn1VmwBANHVkhKBkhSFU
BL+1g28J6Yd4IYJ1lFiQQN6zUK7CLnxJEdTOyrwQnii02KzZ/nybFxv6/ZqLZj04ruePygE/COfc
bqISfb5i4+T0wj/dZaig+qJfZVAxfhCuhhstE2MlMUR33owvays+q7RC9wK5vYh0RJY8PtnHaeQl
odJcQpMGLMadawDPu0SwVOLKF1vWmdgRp2YYH3QDj/gLrXYlm39IxTRNTV94CRYL6TfBg1K22N8Q
GcZYfV+LER5XZi/rhfvyHw/oEVTZDDrtvVyV0Z7ic5cfylBnlPSelKMjh7Zd5HBQxsqQBJrq8WnH
smbq/a8PwPRjs+3WAttzKcp2fWyXBRcIwAT0LRvSXdfMKPer9pW5ganhJMKxa2zf8PfSdF2oxJhz
Kkx1g+R9MUz5c8SN11g0r+jkxdJ4hWLcFK9pmRoNTBsFn7klEMr3REEPtvRJSbbXAOtut1rcudkS
e0CsH3yzy+k4+BEO6kuQzWmGRU6x8+9iRiIVcvM7OomklpsQgpsC/Y5XISoutZa4VuzsN/Kt2odH
6YYc5jVM1+DH5B/sVk+tl+YeNZeDzrb9e05G2rmgAP4A9mhOV56Ds7UjBfosq5mn5wWYMiKOgT+P
f7Swt2XWQiRZgTRTCNsrf/3UAQ2H28lfjHGabs10372F8qEP+gsc8qoc3YaBYVUecKiwY77OhTFT
9YQo2N84XNkIT/PoP3/gJ2B9kJm6nhFKjMJPXcyS6Or/2nQ/sFw69PYh2/Oq35ueFT17rxymfQ50
Mu08EpOUPFjoaKZzqrBGkZLipi07bbwdGYMnjywDpYjX4+/vk+2c477J4xJNUZMw+sJGDiqAN51u
XJMwxIk0z4kLmLvKwDFl2AnmCvWi08mkk+H6oty1j63+RF/p83EOW0fxB13M86hAquq75qov4F+h
jF7Isi/BoqhVNz3QZFK8KueeYMcJjORRzBawP1MVomZsZFzRe7dovIN7K9CU2Iwed7AcdzVwR73X
rx6yxeCLtJzaJFycdaoF62Jk2T0jY6EWEWiwZIQOjGamU1srfhv8su11vQIqHPPtOSzYR+t3iqu3
8gJFKAl3st9dWN+wonycW1ccF3eLfmdhIsrBkRnrNbpUTnegaZkgySPswla6EtYmA6B2Wvs7ytsK
NuLTTqo114aQ6nwrurRCkFkXwMvqSaXtZYLbYYQm6GgkYnehXj7EJdvfrrD7eaZuLU41ZfuMeWiB
/Jz9kXFXsAw3CowxT5TdC7WolZ3WSqSRuDavzFoD1v55s6O3eG8g0sWv5dltPTJ5gl+d99eBZz5d
tmUlOrJRWvMIUbycA6Aa8JmrMMxFZ5MvZotSdOX80Zz1aozIT1Cl+zMoTOAWUE4nvnBizxkBIfFB
mmH46qAyENzl4YNcVzKSUAMN1SjKD9cMT8gpzcAhlY7OYQOmsQ7o9Qn4nE/eX2Jojj9Lt9R3aBez
W+sTXplYbgFUqVH0a+ldoqIBBxQMs4Ly5GU0FuM0WQ4V2KKFX598AXMhxaS21+mivwm1yzgjiVms
F+Ezvy8BemXjMV01Y/67CeJ+eVpVQSk+WXqoYk1SfBOOFJzZyfFIKyBY8pe4ZeLqi5oGetXoPRDv
eBN1lT3kFxn+Q5AhiW/7eC3oRS2jzQnELxgWP+qnAMCqSOC1MMola0bdepKzFtZKARtMAalUplL7
yum8B7aYywVEyTi55BNw6kxwiOH5vmRGYEXo8I32Ilm5QP3Rw7Oc5j2CSEdiV7vnMmS5V9eeeGQP
gLlLeokxuEgRJC2w4B3swDEADCqHTpdh8ITv9U040qFFDk6eqY/pn6vFRQUlOudgXBYrblBWWJUQ
WZISN74oy3MUlYQzNcVyv8GEgq4ppxK3acjCXlOO+p6ywFP152JcNc+eqOCmg/bGiAI+rcwrBWEV
nQQVXeMMozf/uVKG1Ox/Y9boMEI1+HX1IHUBkGkEfd6raEs64siy0Q2MLSYTMkbKq9qEKwwWtfQf
WJTdmIBcc8LV5sMuDPz08nFO7i3Lp/oRikOIvipA2F3AKIbmCZTqlJWJwI1s/Egyy9c2g3chNcUf
4Vxj2/LeKWvdYqLv5gd87nMjGSATVMx5YoGtFii1tbM/M9h5g2aq7FWguDoHU+bW3sbfbsZE+AHK
ZSVtWoFkGboSY3WcKHzHmFQhm8pgPT1zb1BQzKsT2/RDuBPQgdkQUPWi1ePdAP92Wj51O4TVds83
9dI90n5qkhVgT39+lVmSW8IgYjsjAxdyGMgMw4btZcU25lcSYwefPWBvL3DgshVdx3T5cmW7Ih9u
iA2h90oIW22FiA2yHz2N919bXxzhMJwxI4J8o3cRXpCf0IBYMhGqccZ58zM2Cb/yDtQ1AHz6aLm2
kPMMkuUNfwMTBy7bxrBIKav2ijb2ntCwj/IgWpdiiauE7yBuou/mnZ0NfCMuUUcGGMT9iouB+3QC
srhv46o2XRFX8LLoYxe/HKn2/z+smC6nzWZRLPC/MRTdp6ykFuhizTnu0r3FgRtqD0hu8Xl9iboB
ZqKOg9QfoV91LmSgpvLz0A2V7G9OXI94dKE6Vv/vkLeJu3U33LnFU9Hy8WrpH5jIRZLBw/yJ8ILk
YBK85JGGZ2PF7v7s6qk1Um57YiSUzc9i9O7fCimCbU3tOd2wTrlFNEqznA3TilktuVy9bJRqEoKf
/1SQH4IV3DL+qaiOBFnDsiAgrI9g0BjBTr+JFsVuq80yQDQWNN7S8DJWvtvvSazc14WQeBI5muLD
z/1HsVdVq+X4+QxfLMKMoCM3mESZmH07ATMocy++nNLMzCFDLwylPUDUpYq2OcV1FZoCLYyV8gbv
VihSU/D2j5EhPbEI5rNAJ8rz03w8ITBFFVfYayM2GtxkB1o3CakUjZrf8zBiOsdFADLw6E8o8JI/
vu9VJuxBsl+dWPFSPnaXMAJQvC0Z7zYceZRqST8yDpCU2rnYbOLqwLwUGlKtvBz9vLUjrahBa7h1
Y02EDEaH2zbQ129r8F9lqnd2HqCSF24WO0qB+XlpAtuKhHk4Jww0ZYJj/2oPWe0SCNsQ4/kz/oYd
bn/oARZ1evW74uVXBeFU+enw0gQhkUHmLs/WnIPbbyUqgPzllyfnXfuaZ4FfPlvjm3H9FLn00BTS
pp1EksUNcmXLwlK9sFp0AVH1Y6AOLt4+XnUm/Z/Z6dSWwxPWwKmcxf1qWRuHfonGlCfLKsl0M8IW
J11VRdKiVtG7ujpujaLFe63J8GDtJjJtnlJ/wmjaeBkDTCSwtK2Q2K6WJF6ACoXM86nZTaq2h431
2jkp7jzFW823Tg4SLL89QSpUHJA2ds7Lg/m3azfMa6vnoGflQ42NDpdbQz68VrHddaOog0DYyMww
ef2nprftNOC2OkHukcIAuxJ1OicZovSPdvl25G5CaapZKmzSKBIEcOOnu5MxDdGEH75cA2oEkRgq
qdTXdKqQ38NzEo7hcJ4ltm1ux6+FjMXx2Dg3oHPmNYShc3l5PVRv0ct1jIAa/OyBNCWDOaCGBdGN
sPvZwoxbj+GA776PcO4WkYanPoDz72THZj5LYwzIdU7ZgFkVJi3f+803Wp2h90pEFG6y4H8nS62d
wLvV2+QyMa9LkKOXxg+lKHvH1bMYCPnmK0qo2v2twIw8atd3cNolI4q1vh2ohNJxFLycu0HqvGhL
R7aovO6kemAXUCiP1QOESJsMDN0vcn4EcArcUqHbDWxoOQZIydifzhUwCXmoolFniychB2SBzc/I
aeX5lDMgAOjUr3h2jd4JkqJ+84BlfBNgyXfiGmz5GlYTqQV5jWcMJG/nfZwSwgN7dQhGBzfeTRFm
uiNqHY5bnZBgDruKiUy+X27RiXHel7pV1n0IS1nEcRWQdWhRmkSf1H21lvl0gHVMRDZOdakUDr1n
6PBhlXLwSj0Vc/4Cw1gcUzHfES9z9KaqUygylxFGpXPCimTnedWzEjbxpeiwzGh4PrDmHHZE5Dgc
CJOA/R6ncJ1c5DtszzJnr6PwxmcNS12UUVg4aYwGos1x1gzTajWaGCXAu8I1YJH8CLNIoZFcFCVr
kenmurLAX4My/Z8coiQBX4zScU1/5yLqFVKz9iWFowCTHJzudKcbLRVhD+u16HF6n8XrC4QsX/m3
qLRSGI9Bebh9/q1vkBFFgjirp0qJuRA8o52S1uaE9Z97SphVKp8IP0jFon5ms2IO5kRHRLsg0+vs
AYHDsQHzWOI6q57zBrt9FGA3EQ4yPQWQSXPfw0StNOrmyDnthedXeVxkB+RWUSUtfjFU0uTLjV0+
YQUKh0nhzQvW8TLcM7D3/RyGx5FtyAZGeo+yG/TM+EOIF0GPOqllDjgh9UBRWeFZ9dMcrPEFsbpn
NdWsbFQUXnhKfxEk1R7CyS0E8OVXLjvaggCSzxbvTvsetMEPIjm9wK6tMOdLmrKMacnde2bxY3te
HqP7UTgiTcJgDg7ljdzubJkkJwoOwsqF1PFwGhR52KcOTNcICNvOoTc+Ix7iBM3n5goBBQUp1F7G
h4CH6fDDRD+bRnVL+HAlXbTM9uMUhGuFIu4kiMyIp9Q1nq2JboibcWAtc1tNVoSoKOqV3p9/SsAY
RK323Bj2AQV0GCGKnD4UUpDjJ2D6mu+hstjdPA6MiYg0Y+DlGhuzvuFks+4BGi2PNr+ZmkGhKp6I
eNaSH1t9PAKNaVnBAfxQhJlPcpYCLCjPex9Jcp+fw39gHYBRbccxeZvN1NULaQ3N3inEv7tOLsM1
GagXbVg8Y8jnbmCS5pp2Ao/Q4blwxk3v8ye/Uk9G/MwgqVOLK6xjX6F/Q7Lx/IIRzfxRw5kf56Wx
/CClBUXSp2YNDebEsZJcBimklKwOqVnOt7Vs5E4ezvp3zrl5nlGgwSEAM/QAhZUNvbvWJlLrI81H
OgNrKQ1T0e8R60Ud/Cc7FlEb5HGMt9uYX3f49nyEVMDtPQlUHX2f9sM8ZU+VTC9ZmYbEsk79ZZL+
l9pK1lneqa1Z6+JNWJzhqpLaN0hTHbGOgR1xrijMg3UqUysT5mbLyAUcmG1QF2HyMFeaZiyMMJkm
A5hofWTdtC6aecYvoMVkfjb6HOMveAlzyEhPSuTptiabKl5CTh8QaqDDIrhfdJL05q1NGgqyu5Vg
tw9e3/KTTl6bi+jZHcaSWwdzhG7vt6O2Qs3ID9eNrjymT6AecHss8D6jLeRb6rge+SVXBeKZgjDd
kVBp++DfnfcleVOX6nYR6o9pzFnCF1sATp1NUdISf5NEBn0wmVelFcCCLlCSkIfXaF5ZKW4ZUnAz
ZMXPjbo5nOmq/tGn6mMgqyLfRsVaNTC2rZPpKyj1SDConWIiLTJKYTeoqQuNEFcZguzfJyTPPdap
dpZRGN4PCdFvwqKIxTWlq/XVmx8OWkY7lg7M24JRW2DB2hz0qQeN2RVHuFyb1rhsEgBjFihd4Eqy
QbAIT5iD4UqQVsqkMnydTgO5bgXdwVEotr/3jAerxrP95SzuikMnD0tQrBV4yPYoLZ5Ko3tJUkAE
jBpr5OQYk+2Z34Y7AFJR4VD3LqtLfecefDyG3zYkQBn0ey5i7t/mKj2iibVj9y0DNQJE92lMbUl/
gng1HP5LUr2nkDnnzkIpmYG7yQhtEvlqWjbhdpaYGg1B+/FEdAII4ELlQUOxepWYjEUrNZvYdyrR
m1vUSMR5vnDtizYp3Icy2OHtwtQdrRL8fLVZKcKi2j9hpmNcppJKLGXBSgjAKiYRi9TX8m5IFkth
LM0gv10vGLNkpYB0eJ0HDL0r7D3YCMeV4t8dQH7gEaYu2l7Pt0GDzp/R/b6vgxX2+MAc/4oghFma
cYZ2A+shB9HmO12/yBlYocu9FtlVk9/oGKdEaEqqA49oICdCWRhBMQkSk6jNsh3fTmVGpupQIPxq
KXN5U8P/PAaaZd1TuYTpPoGyLjEp8jkQ7zmKnkd5DhxuBsYIJBO/29NxfEvieEX2IyIFyLlAm62z
Vj8uIy0EihnbyxCgi84ueLrqse8X/7jtNEFbIovENS/NuoYihtJaCAp/2OX/GwHIda4AsmRtOnxW
loRvXQs/r8f85qHtfj6bz28Gd1zI3VWrLjerZvXggoD9c7w85tjsu6lVzviTjD959O1bGDdnCZmu
PSX/7mJOToigxBPWMQE+Ha+LTEICin4NWoD0scrVv9FyiI57CNbRXknujiAM3+Lsay4HoXJyVdij
RwQ/NBlqCBKLQMdMuzxBaIi4jaxMAnpDGemid+4JUryQ+Dd+t8s3p0CwC76mDOdYkiTi4DBEcd7D
a13TdzUnxCCWtX83pqJknG5PiDLhXb8FHMS90NN03Pm8ySOrRd7E8aEPP9A/FNHGiOGohOD6dNbt
m7MPEwnATCFDBwckfW5Tn7jM+g2MMPzcLGhHDxzh/RoQia0AiFhfVEKTXNZsZDiW3Ur/oNCAiMzc
i8HK7b3eOaVmLVKL2mqZacNk4TwcgyjCwhi2/++EuDQ6osPhWi6CbMZ8jQj7o10BQMU6ZezoRnI1
qE3heUxGyoGHnGmur9ueVc0ruTAGpso24zgZUQbbWP51lrwMq4IoOrGgFDvdS+tn9RSfLItFXCo7
5XglNwV5w7qOeo8uuhM6SoNt5EVl3HFky4mgnUKG/eKcQY3xDwR+IQjJ2Cn4codvXgYhcMks290y
rIlvnB4/bCqOXYNH1T2GnqlbW+y7dazaOcz9hWU3HQDhgn3inTWE4Ox6bg/BYGvcWQS8ynWZ1bFc
cdIGJZ4z/P5nKhTmk5hj1j+WC+XfmkGAVANAF8GOLiXjl33lSKjMcB3bHyZigQnWHnL7cAPXfmCY
CUoTE0ixHyuVToyWa44pIDyDV+Lm+URpeahcEc1kNDnGdrYc/g3oApMuLlCBm6lki7zew8FHu60w
zcKoD58OsDZt9SfYbhFzzC5n2kVIS9yI6sYnAz7PRO6a7vHGkAk5mKhTDGIgRqLKMQWuRQ1lgOYj
LeILhwY7SbUR+sfAyyre1cdDB9xeFVMEr2ylHA3i/yUrbAvSml9jzqohSxINMMc67sgIfQr4LJT5
tqBT9Dtbyo2/kLIMDYHedNctqViwY5C94r4kPqrGKbVivGmOtG2s4hU2R4KrnUtf7fJIs0Bjmn/C
/AzyLjQMqfW0SoDGOMnliVK/BvdtSzXPqQ5JsC+CHyd2FZexbY5gyjiYDlOgSKQ5E/ASEfrFtSSo
q2ktNWsiXXT+vicvZt2Z3TEgjcFwJxWSMIGNWSUho8c4ilFwEt434da1pO9HXqIjv8mfmqDElx7y
JtlINHl9BeIS2QdpdgZ+wzsvvzK4R9BGQ/1aGzPUNN0PTbESVTOL3T5fOZn3aflgquVgctlY8RiY
AtgTbBpzdLxWPR7BJ9LKqR2qA31wMEKQQWSDIv5i0aWOKbT70KokA5xsclLHYqbMfhe4G7pb/Sb1
MnixKiRzeRXdDOLh8vz2TwxEmNSsRLzEwRKRqR+nyYuGehtD/ggP0G7eb0A6k/BwWVK9L7bBs9R6
rOdXJPyRoigFEJkfJlUIa7lAnJasNcKDz8wXccBezG/5kWRz0t5zC6KFCgp5O9f+43o8r5i20aSM
eI68VjxMlmiG4JEBxUt6qz7S7moumlIlvzoQ2xnoQQpvVweXNC6Uz1Fi5hsdmaJ6Umvx5N8OkTXj
u8fQ/DGaogjaiPG2wxcc03gUlhHB4Hpi7NVlsSmToZ2mjZoDjigc0JZXosfuy47ibHc8mNIoe1qm
JBjKMsB0kKqoQ7iZ6NOv+iepd/nyFoMM8p11S38WSA6UxqZWOK7VL4qm7LG0YOq4NX+576ihUFwc
Wia9ZzO8vdvNFZiSEtDRISrxNhCwLf9ANQNBKmBzSEmzSC7piDHWv5S985PfaxWqRzSh8AlZjFNt
LRos+1Y+3+KhjWkd79VT38VYkBl8IVqdwS0ifmjhbRfniz2a1bAgyX02cRBe6nbxrJKbVv+kwIDK
/Gytw5uEGLsUc2fxsNrQQRv6sACeFxLIkLKwziSwyRAe69NXkcUGPGn0ayrD+H/Hl+IiRnS/1ZkQ
/AtAq+MCmMW2RQ0gzSmjNBlsML1dAIUE8dak4HFWBfHWZKkS89ISr6wkRBr7JwHjmKCW6KoFVq5O
FF0yKDjwadJt84Ny07cduuwRXk7Ec2k2g10G4DThdlJGehjYJhZos4kDvV/y8D9WrssRJi1WfZXm
jUi+NZm4p/iufVQ38mEZMmnHswHG27eWYSoJNMZd/Jv/7nNWIFXgEzF1Np2aJoMyLZiln1+6bWvZ
fht7g0o1VNJgXZI3ey3JPqmqX5MW/l36hvX0CZlKvVJYrgE1bzZgz4OQ77jqYirsoTfdnRtV/viD
yRwCTQYZ6sTaPRoc5vlnTkrIpSKAEa757WbV0k8jp4l47ic9ijIaX14zR7PpN3QBqFV2lw7rtds0
b4QQYAMYzVLCR0PP6jfdRXVI/HidOGIWZb8efg2oc/rxfVQB/QNNIzwMqBRi/rzTKGN83gh8o7Qc
/uRFeQ9ORBIkoBbNG6D51gcQAmQL4mfUGZo3v0bJFRzcRfNM0uRiDGWUCStvwIdYkdUhSrNuqvvo
MHDDG4yYXMsLLQYVILzOHEEpQ3khTDz7EABrkPfEADSpyh3P7pCKC8rLEaHqFVSTrtJBj3itzr5f
nHm5BmvwM7tTzywdaRQhA88aiYDPyqvCcR+ySd9yMFE5Hb2zTzfjyvFYi9pZ9c1YiYyEeASHr9on
XXBzqmarnnNuCpaHGJ2WegJ220UoqoLPZBuQBBRa92hKa8Fplmc5f4yxJ8UAlwoIneTwUxtw/AUE
bj9BpI71gVlRrrKyPODr2HpICsQkozyMJkyEM2tcGtPUefhDI1QboVe407CXmNXo1ix3MjXfyxQ9
X/JlccQlbxN5Q6hvgqf04Yh9mny2O15UC59m0T2Lglhi/GK0XwnRzcXTmbS1srfgYeDZEoOHdFKS
OO7g0K7hswVVvJKFZMBvYb7awXNPWjzdlgoPLfNUVTrSUht3jqfbYvUP4Vl/sKpgM8K7lYVxXSIJ
W2mDDstK8MmWyd3CscmB7eqNog5Jwc2o4dJVXpgbUVeftKo54ZpkTafKOVivLL6wGWFjKShPJGDt
LNALO0BN7iPXhNjwXDVrzSV8nW4XdhztH3zqByH6U+QOEpjp+KpLzeSMoQ+AF9YmLL89wONWJzL3
b8Iq4TUi+wr4yVM7w7IlzWm3ceFJTut88NkoRCDShVxZqVnHfs3cAMVbINv8YKnfLfv5o16fbVbH
45vakiR1nezZW6UVzAmleABs0enxaz7pb0ck0TVdu1glNZvA3fdQraG2djnBXmua9pJTLN6NvPpI
2qR8ETAZ19Q6YQLgyy7RnLNuyTyshy95g60OZmTcpi30JtufFYgSrr73iVfWNanP/cfi6H8Le9AR
kzkbTDy7QCNEIS9jsVhPP9CdO1Dgohh1MEhvS0+WmXg1Z5J6wnHje8nUOx7kywvzAGEgG9rjxdCQ
PdRnhv2ObvoTUwvs7hmuM07q/GpZoJkpNW57F9Fz1NW81EB6gdLx3Tx0Jr1Tl4pvIZWUhmjRDWic
bbXiUubzlI+2IrxpDV14vdChb+dvXESuVgkxIxbw192AwAkaMlt5YIPgwIwPg9qgzwL007UHJD2Q
dvdyC7unXs84vBIn8oY8nvPtUyorYgoGQd2voH3k1ateGZPZ7KAqrUETEk0qHletYthgJnu1g3ro
frY/IoafSfaZq9Se/VyBY6W0KcHkIQothlaFekUDXFXWnnBx4usXtTKMOKMRIOTFZmZj0hO5TUze
YNQ1JKbO6beQ7qaKoJRcCslnIT03gSN7/z4NnozMLpPcnRtA7BoP+FBJ7V6wmiAJ/cmCEW6L0VHk
OvtDoX3oinROCFSH69n/S6H7+l2PeKdI4n0HdJVATC2M3LNHEw/sxmYt5o7co/zxP0DpFhPD8k1O
o6AGwBcoyG/a3owdYupv2axIfq7U6rz+ajFwlhy/w2tbTpvODIWmMeW7p5zXvu4qW4iDKHfzGH2F
GK5sfPvq8U1uIhRgKMXG++BFctGl4IfQf615kyoKCmrc0u0Raw2RRdG+13wr2Q7C6goUcc4FBTLB
FUJCrhtDTtsNSr1N5CliY04HBLG4PqgajCEkqqYTwZ/witSs5kO5707qm2FV0wWXLl0IQCt/TBJx
Y2W2YkH0dEGiVBL9sdQY6rLO9oGTrtc0GjubWdBw5xnncH0hytCqi7ZXIxXud3LGd/ZtWOHG8yyA
1ttI6JAtmiJxwZs9Idk+usPUfAAfudZS1/gO5UzqBaEJT6UjKnDdp0dmbQJYWUyNHwn46Wu+IDig
f7Mvl3CeYsRssD9Q2j9w9Znzkoc5MTpGnJCKXRq1m1GdoLIxaDEsAP2dwGD4TONdkszQTEx/0B+v
76+YUFHHG89X6M2YYEi1cmTG4fqPnKHYQCoVbCwAR/roJmZ9MbOhV5rOHRP1zs0S6yjOn6KL+kYE
xYDSMzevdkR6WpOp++Mwx7Paov10ERLN8Y+8Rl/6cbOWkE+u7dvWX6VZ4kHrl8HETmJa+/kdpJ8l
Yn8alINXTFZDXupBa+X3PdqxGyhAd+KHeR6saVMI/ljdJ1AhV24/Ntt3bUU1DzO/71VzZcKfLzjL
02mpqFdqKvWEDEWAN6QBc89z23TRmxnN/Wlka80E8fpvqCccMUr6RTy5TKeReKCG/278ODjSpYgt
bwmfVY5XeWVhXmdvazTH3AVcXLJ5vYoQPfi7IhZ65dH5rGRuyyYPlkKYdxva5Q03pLy7926nRXFN
SzRB4SGIygSwcovRLnkYaPxZJC9DYUnmvDt/Mr/kKgspaedU4yIoD3uR8E8WrhZSQiXk/E8gEFZW
p8bqYzh2ricfxoZdX/V1uw6DBx+EbZq7//hBbiA3LMVNSxqaRgjycW1zrv6+4AhfP2VEAPi7wUNb
0maxfmGo/tfsvyObcTZjyVMCbmxDiTRxCE+1iEp6kDzd/jKMvRFVzAZaWpX4VcebZlrXV7rU2wR1
Xldkjj/P9Eu1ktM6rhJCQbfMj3nsuvrKYLGr7qX7Jf4hQKCH3BOhJ+UD+i/N+vI70C0TmypHiy3/
g8WMWePXgqXTxeYEVcMLoqOgsZPM8kN/WqWBJsfS5q7xqVV7OFK2BA6wdTwWhE06B8Wd7D+BrDcz
AA6EWuppMSAUjmEXm7PtGu+xf6yyqTc1CEXTXYeTz1JruLDQFvIOZWJsICNoRPqfQJX1AZiObUqo
ObLLZzNJ2FNjIAjSiHjCS1b+I6GjFscZ2yP0PRVAYRdbjM+AYv/JtzcDRHJGOKcA+XprLCKx62wU
WRbc8LrgoXHYRaw2b7L0ptxEj15u8T62iFxLFoDUxUPLIL0r6MtBbkOCW5N8peDj272KlFjmvhnt
rt+BDLE0oP9wxHj8lO4HFdT4SaAEndfMJ5fof+EXtrPi7d/QXA+TMBNecLy0NbIfGtqkcI6Zp40s
EkEG5bSYvUPPu0O1BKKZbpYNh7NMMAycE+Nsfd3s2CTqQaKIE6f4WLarxODgubVDau4gIhE8PGqE
4XdS32S3DrselEpVikZTM/yp15trAhSl/18UErMl4fy98jwAS/z5boiGkSRk3Iwa8Pi+1H2ULwJB
J5Q3LB35EoaRRx3u4zeu2HuOd0ZFhyt1uDQjS4FhIbJvid9D9xOrdfKb6cVugSmMmM0HgJLpAYOR
Bl+1xB08ryXDpL3YhwbsjHnYC8TCqNucaXGJ/OLgo1mayo2g5K2G3to42+6G6IZrOgLWflE1qZ3K
r3mMgrgLurGoIZw6sRkD7D4gFv8ioBEcmiFV3/yu2LvRxoWrbJlKZpEOc1NZ+KEcAp2DlFc4R/u5
rU1DMzYwLThXpvBI61mEdYngdjsza6cmEvMwdGGpvRKqHzQCueGSBQsBWSP4YO9vsl2RpnwHDLxM
GEexkyGCwNgbNEQY5SYjnLM91C06EZRJ4FpUrSZoXk46hbBkLASc3Myst867+l0jfrw5w0f0mgx4
gNPC4Bqic/D7MFWqXI2aCeL/DNv4vakBV3e8sL7Ad61rgAJLUoRmDAHlyxrY80QS4rCgP2JucTNK
2WRL0hP7tl3Q5LNkethzZg5LvUMpznwEYZ5B4bTfK14O0VpqUvkIFrtzH738PKJuoz7dGJU5p0Pm
Wba/mp6WMJouyviMROnQ1eCco54Aq7p0JOOUOX0n2H7nQXK9HjJRMy0ykklgufLNwd4c4S+uo61Z
B7h+XUcDUsmuoMpNfrHP4fI7ccI2vE5EXfCm2La6/fM/vsa3TDp3KGdmMkyHFRJ5aMMjl+1CCU01
+ysVhdMys/9TZFb6sjOl03bKvAuqyPUMTrIDSN1GqSNy1Aw7rLAsSZ6eZCHFfaB2B+esOEPMJ2c0
u1sF2ktEFun+UFjQajzV3DzsqNdqu/uCLJiWry07SGoNqncYu4q85z7PKw3cjB7Kc4kF1665Mps+
79GlPTraltzUS/Wj7m1qnG/2RyrapR1hlZ5Yo7PZY3r+OtjsiJnQ2ITy07jsfMaM280BvjzuhG6k
+gEWqyTHBpndZhhat75tLfTihVfMeKF7OAbJrv3E47Z/+MfSvBQ4pU7Jhm7nAacp1z6KaJmAu7Uf
THT64UV0TuGHoWp9J3vu8fHO4r+jpxxQLQLyVkZXS9rcbsxV3Y3ATrh7O3INAj/KOmtCMGec08ms
IH0dtQviqtnviExjYgCch+yznyBH9K+BzJwCJkgEGH92yW7Tqq9RgISaXkbI4Lyi0ON7iwSVHFcz
qM3jHH30rp+9agGUnEOHWxiAPgnNasY8dStsBbCIJWxmoKox3kvUZW1Yn1VtU4q2MhKu5LVVQ4Kr
rTplirTP0c9QBUVtm5Lm++B8jOhE7gr2xgVZpQAF4FVT/jVWkhhZZqMgNCvwoxiX8mFuGzFvbR6z
RajiKVvFK8+9y59iXWoVNV9FaHNB4qBMi1DlHBILl6D9WUGn+AdlIhc1OkDxqgQsciLBGW0YzZoC
RP8mCxw2Ijz75+3cumcFsrzsAJTtq+EJ1BEYdMBcNp84m8qWhVBYBfx8D1fx89BFViO39rmetoME
VgzKZeo47R1+S6AWIeNtNivGOt8vuyOqtgD/lPjW94avbIOtkhjlRGqsiPIy2h4N8gzDuiDKpIQ4
KKe3zpO4OmNlc9RGVYk8g17DW9r/eBMmaw8ESaJw/wqW7UEf2ctikl61Qidj9Lzz+WtlmB0soZlX
/4rvLlUgJQ+sKxnxf6MdbriuDT61W/Ez2bE+TO/lOeDgy3Og3NkNe4u6bZ+etl6JmCmLk1DgGOxa
SRg/if2jsTOKAf2sz8csvBLRh5t5rTXTpidkByp5wKsSfnMLgGMjuWyNBqUCxpifbrYLYlnEhDMp
MLFL4YVMzp3XOdt3vtG5QuU+NumUkbhHZ8YeZyhr7bMHNDmyJZBoS17B7edbITFIEOA9daxhEouL
zzH/pBM6B39jhWq/YJY0GBcXqnwi0Qjy/Y8poXW8dFMf3rJ6KIYqFw3jgAsY2cnGV/RNl+6SQZ/k
DZ7mDvTRRTlYWiRntwyaAuZai2uGeWCnmvsBDWOcH8EwKQjkHODCfAIlxbh+XRY6eBAfu1rWAvEG
0fNe9jTcu3DgtUzmXev+1ow3XE+q3oDhpJam9s60iHkQCvqBRGnyHCwvER0IfE8SK3FqYwBZswer
Hi9nllpooAA09MHsUe2F6oEqKAdeDllzxFyr+D1Gt6Y07B3cxcWhQZV2cMvnklsszdjIcq7aRsqf
ERdIwRvdUGe1DmiZfm4G0JVIzD6b8Wo7ugGGX8wPDXFjdvUxEm5BkYODaX4wLxxRU3TJaz9abeuc
stmnj+/OjEd0qRgDjzpiYdY+0qpJYvgJ58qxswCMTEMK2G5AWyNqZ1gK6e0e0JldaBQXzWC/btnz
BiOYNBKyV6CQnZ4epqMvqvVeYvgC6pshDuLgdasyPpq90zKSRMslnkIalUr4EXbU4ZAWSZLRsbNj
jMuRn3MkcnFjMBAk1FUpfukr0F1beupFDRw9M8QKXmQOfbRVG8PVzRkTvzk+tih+tV9F4S3Uv2LH
/KZvdvmErCkLlZHXnRrIGXCHRrISYzuubpiKk6BeC9Jl904P5hBDeKFKmKGJQHs9+z++VBYv3CQT
UdwoNiAVHnUfNVls5C8xPwPLq2gWfO44LgJdPEOqBr0a806+7evWuvcltVQNQOV3KLW4QGCwu93N
k+Z5S/todbjlDS7uJj0B4MBQkgr8u2wdyRT1vEY1iVDAvM2NA3jXYJcIBlr2wn+r2/XhbXi2aC/0
ijDsclDjoaoH1TdO/Ox7n1hF/P6IVmTS0GdzFbMPVLB/9DjT8CHveQRFyaLgM2S8TAs2sdszi8y9
rKzT3QVS4FUcO4lFkreBk9/Oks0kfiBVEXlrRtPPTZhqYkwtrj9p3/a4zN7VHRPfS9yBZASnOK9I
wxAenyEisNDXYhdTewPDcpUlWkf74yNJafynm+4nXBgoooVoXaK09ap0P4iKxgBbg02UvjVyrRgw
lvN4CHfBwPMpjmKur9x2fA/Ykv2/j3EhAvhbTa005vVZqbj8+eJc9e8htdIue2ZNvDeHiAUVwgCB
MxrbNkK170thsoGSR4ITxMFLcN6vPKWdEeB8wU8+Gs3DSw20qWjcDN+lHwh9xPAMbqZQzGr57Fpi
slLe8cC+l+aAG0SszwXnPygl1hDo4NmOb9zMiRwcoe/ibLvhD/IPt0dy3Xy+TARp5nB0qkhYEpee
zjKxK/wZcOuDsb+DJF47xQGwaNwiHaFJy9dM6O4YaBUL5KrLNTxOmIepdWN+rTl7tclGpQey68YF
VyPtT1vfcBgVGkeTA78qoQPP+1zb+Pz/qqeyIdXUEmwMtSDDOnPFMRNxnrCwLf6bJ+oKMWpAGMQe
04azDti92izVs/JWx2wqrOe3uRacD+GSgSlYfGlFR7nKCWZhLf6PlrNPZ8IsYfQPcJGrQ0Xvk4Eg
0ev/EsS+1ILSobinbbbWhCXRzF7lXKvr2d+3ChzIq2Xh0o+kYGeX9RNoclIk9dB209g2Wk5/yVp/
l1zQHxKyTsAApqepsuIoAQN2OuV430fC7XHZvVT8SWTVSXNfI101YJCvQsFosEBsgELYZRk1v0uO
yhOGOhpYiNj1FTUR0ytCyfVdQW7FG3/6nS9t+AAZ0EnmhL+Eyp+ISN2IyKZEKP8yWlNCku0eYc+I
8WUsgivn7Df+NHP60p99gJZD+X5RJGHOySV7A4kNZjWl3CDeNCqY0fdSS1a5a2+opmPsFl/1h8jw
OVwdKQW3D9lbduhYiTrSYamWylrYCAQg88QIRG7vIJMF6XiXu3O+UJ8c2puU9Nv3dko9t1TyMZ5z
8mMfLPMw2ikmHK0/PfiOWF4KEyshUcmhnGvAnJb2Pcw3ViIkKtoSiCsY7FuOJRWtsDZju7bFfe/U
QyR9yGK5JJ8uOG2/jC/uNt4sFmiU/W2pzLVlMOnrXpKTtxks8V4DP78KPCvQ8nvj5o9bsbebbGGZ
z1FkuLWZagqeOJ8ugujbpTZhF0Fcae+7wZXkT1GUJA50muQj3AH8AgWYibC7JE5GD9MQ0g80IzS3
VYQzgTUkMI7A6O9B5OFRqKvAjTHeCCXwd9m+sOubGMqURwikbjV5zkoWf3m/quupPislCKXc7+1P
lf2UKV/8vw6KZrvyBQGWraZ7zxluZjp3NoBIrW17nJMvnNiEHrRQxJgsT7IFsK0JOUgHkI5gpD6J
K1ZUTVx6hPw9SA0g+8z31xE8VMB/yoPD2K7fY6en902E/V6sbCFlqwnxQmntDca2fwpAWe3nV0Fn
vaOdZxrmF1+pot2dQc9Lzypw6G3FV0mAzWJF0eb0oqoR9JmpzGXbm6WhOPWNM/Nb+CoeDBrO0jgi
kIZaLHdmn3Xh722mjog/Ydz3vE7B0pgXRkg3G50UlRfe7ARBXijfNX35OUMnvDZcrKetUssv59/G
nL1y6xWbPuv/ZNhbNOCgzvQx6dD8f6qbjgaLIqMUEglOZrpsZp4IUqPji1Q0WD9m9dXL2Eqmm94D
L9Cg78CB/4ext0gbx5BglNBbRS5gvb5L3DBY6+wxAIFzIiXcZZCNjs81z+sERBoz2LP11X9Mi8RH
9zNa+Ik4ninLIIqFkDDgLmEo5sUsgjruOgnaB/dsDl/jLuZjnwXfLsEanBmySpwUEmf0U0JhFB/U
nAXkOaaSctPSsCAkQxkdPMEObQ/YwkHzpgD6rn2GHQw8kPdrgO2OjtRKinYnLDgehm2c13Z7rXL1
KuxgJOXXt+15bLPOTU6K
`protect end_protected
