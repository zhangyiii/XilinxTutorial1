`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5408)
`protect data_block
hTX64IeLyHzfa3tJyS5Dfu7W58OMH7owjA+xaI0LFp3aXNyg/WgFR8UzwM1yxxpfSMxMLurv/pZl
MKFlgt/ZlX2hcyFiwMGgRgwKsTH5UTE1FAonciR721mJ6qT3Og6sAO2HXKuvAyylBmNK7C9EiD2I
7UcyfE/vTfUlAvUxm7kqrF1jFYKU3zSXu2kCqyg4buM+WwonwpfnTqu3ESdT4Ce0i7iQg6Ja3WXS
bA/Aq7XMwyr4z/C5Dkprg9zTPAX3Y56sUxpi7zxb5jqNe7CdUNefkSOw7ss8wWgauKMIQgn8vRAY
zTloQgY3lkA2pArlzWCukV3efPAzKfowk+hLDXP2Do+uJoGnwTwiv4Ta3NPkWoO+nQLSJ9/tyHzj
F6zvp2hvoup2ZybRoaIqbHmqAOkjT3o0ou9WQ672JcSoDF/4Gk8Olk2c+E+ghaswATOpM+T6nLxY
v87m9AYzpxizbCIR+wj4+ONBGapzQyFt69O4pThH6VmVJnHNobD4cylBwcp8Ldt2jK+MAK3dHCtq
1UfiSd6OfevvCGEnFO3BzdMqbCtvYa9klS6nX6DoSaa2qonA9ttsow7eTvFdO7DNT3UPVI2DkaUE
M/tR1AzFh6OL18rAWelTVuhqTFyWTWIx27LMaYePMJV6mQAL8tud2QLpSVFDdp7yEzZdHmGsygfM
wvCBtcvJMM8X9msVB40A3kVxi4sySJ1Y4l+x0P+9WC2K/4cfh1KWZPNjKfg1xIcUIvM/IoU2sjpB
h0so2sCp8kBTKDj78UHDVtCd98RQC/Ug1LZkz/KI0cFK4gh3APIaaojGDlCzVpoGkN/FzRE8AtXv
iNBz5sgiyIOAH0AVgUShxImM0mXpTg+TZwTAx1AVy2Svcp89jK2z/DslVlodh7NPyEzWmKC176Jq
rltJpAvzidfXu5ZJN9afHAMtzwzYHTug/qWsMMNo/Cb409FaTQfAQpraPAzRuveTDjD4NaBprwrB
UAgB+6LiDw+8s848s+O8a7tN1SNDIvTG5zg3IE36amcpECRPMnSQr3Otda6T9qGitskDaNyShs81
a98WgWRogi9uugncdl3EdqXyOBQrqmVAytvg/akorH/bWto6R4TQZt9hjnen5VULghlmET7aeRZP
PD7+qBV1g4dlu49MZ1M3boA0z0OwXSlVye1s9XxCvczJe+sbAXgzBWUFgRZTMfJ2efVZFSsZGEel
SgDrlV+ZEcP3Yx0IJC9Ww0gsKLagskRL+ud0SJ83eLE7uq8pBTnAy9wxtkG/sz1mOSjFcoUy8A5e
Nbqhzck2sb3puJc4kVuZc61VY5dGyPr1SpVxKgmgbKc/FZ0dMoyo1IyMJ8IH29yd+zwLxrG6B4RZ
jhoON2Jzxl+qBEWmG4y1UmVFYKN2zqRe8Gm2drqFGEAC1GflBJPTeD2v2nFRHUdwvo7i5/7Y2dr2
g4ZUrTR6cfPDgAkgGzscFGlSG/0wQU2y3JmGj/iZWfZnCbUdYkqn6WFUJCo2assisY2AZzC3ZjsV
Tn8Yq0hvPfqZXYkLNcZqSuB7shC+7wCW7d6IeDtxlcF1VPdA7nEYu3dFmQK9oOXxWNIZz+vRg0W1
SykzZ9RidwpVA2RbjvbWj6dXp5yG52pMCBBDhZNDi4iFcfhWzhpmWrvcFb9BW9B52LYEs33/ivz7
882CicXRtcJdDcxo4XIzfvLAQKv5Dhg1divVe9L5BMx2F1/xgAmD5KrTZxbHiE6WV3suCGgL8YqE
KDYbEPgiRdwNn/XiVm7ZOPFOhz+FvjoHPp0JEiClNoycg7MD4L2WTi6aY3LSWD6PuEd0BA/JptsA
yygibp7mksLoA9bgAW2x7t0BOtC/KRMNgqFqldTILgW8Lo1OmulRgmS3zfgUnaBJJdEIgVdbMxFC
DR8cNTKg2e6+3KKdVliSGGbmK4AdOPv2ReQmdEIhMPCXyZHKvRzyVYTe2I40Cy10qyhaJa2Oxapl
xG/MO7owi0tiK+w9otjlIuyjgz9J2bL1Y5jhNLNhtQqL6aCfC5K4bYOQCITw4J36Xdd7YCCmi+Tl
fO/V10F0moSQp/B6Sm/a7FgJF306OD9CJ1N085jb6pT9jK8+auIlgbn4HsJCzk+G5qvCRsCVJRct
8TAJ7RWTjxFHEmW5+quRxhTFpkKNrZIrtO81cPhtfWLC6mLVAz8FwWuq3d4gAD8kIspKWT8RtuuR
ebQnuEXkYka+axZYbvO3xu+5eXMVzXwYCmx1oMz0nfg6G18vlRz5VyW+tVVSFdpk4lg4lKZ8owFi
5FNSvZMIXKaVW6XD4nWpsh7Q7KE4x3OsaBE3f+4KqX9sWs+3nKsKtBxu6TLXKMMDQUvP6fLz3HLQ
t7j6GF7McA0/OOXoq0F/tXQQV7D4n8TZ6AD28H/t5HhquVb2/SlXWNp61zerFgkRoJXMPKPYQlzZ
2kRE8YICDsCE8xSePguuEFHj3+vX/FHGJqFlwCznH5vhcF4lSGNW220Zu6ngQdjnS1bVpP2F2AyS
w37L/72XS8156GfSbxjg6fO3llIMnuHwQR6oiauzRIN4pFTTmNJOdl7nfJiVU8ufZfB3AW8j1nEX
N8u9BB9rpNz5vWlPMNusDp1idqDa3UAhfO+DwtJ3QSBxV7AdbUKxtpBa0uIcZRoko0dm4r6owslz
1qMONELul86nsVw8e1O3NZ0wLpE0RROTi7k/dNIk8vtirM5XIBBdRl5aj2LPkoC+CBkFDzMslmjM
oZJ4PCbBlXNOQ/aCd7L4TIBv4nNSxsHG1T2bm+kk39GJ7OXufZG733Jg6Jsqraa+4iIIDFkWcKiP
XxSNb3AvaYpASuWcK9t3i5kpcUoAEptoE9pFZ40ozbWy4WjnPDbq7laD/kLLLCt9qxP2fknl8MXB
IMCELT/0Xv7k53V6oSBsD5rXK8RrB9NKV/dZG70yFo+BEBoUZGXuMkUMOk/8T14eDz79qB88gpyl
LSF8Fz9WoAohtUOnGE9aCFmf3yc6HWoLZMU6/IJfF+v1HuO2BJShZrGvf7zlw/kO5fXpwpNanCbI
RUg+XKH77Ex+bbrlFKi7e5+5p11MQ9R68pVe89txFHd4pt68s7SfQoUwQp8ATVcl8L3ewaagKozW
aDTjcpLIACT95fHWkY3aNzowk6us/YvAv4oD52CnFNptSfEFlsnAHyTVW000AGXJlt7A00e8mQtF
ZTO7nevAqUoemSKdX1DzOmnmzVs4R2nvsNpH6B17ydF3dMXn/VnR/kj9mI0Te86H0m8Jlse4Z+GT
yGUp56qCeMuKJTW8HjFG6FqA5wSEiWPZY2u0JYK9c/EIDPxCDWcs5gwNtkFUk8DTPifsznJ3TyOD
Dm2YWnnX/SEPPYH5OCwSgxfYhlX0sZFdlG7A7ysxf6YXpC2VK2fRkRhjUtNFHt0odJtVvs4rlQua
i+J0cxlWU/NyMF0z0SLX8ZXvdO4/f33UqZ8lhURyheVwXEXez4b5J+pSNIdPw8xvO4T4QU30mXcz
9t36X2DxwZiJeNNG2f4kGmbl6u4YLRK1Eykw8ifN/mgrkLiw9CHNgwIfy2YW92GknpEQRQ8FAtsf
TE3ZSpy9vNWLn+qi3fumj9UCiCsjzAWC2IwECFf/TAAYs4CI6BZSG/oOMZyH758L7tCr6UzMys1A
eM6C2Pt8HZCiyn4hCoyU/rJ1Q+wKAPll33jChITqI67hxSfU/NYaWm4JYdV3HqWEpsge7c2zR02C
EiYIkStbJ9d7JoocYpO9ToycMBUheBSkrJdtdeS6j8Jjjv5t06JCgFJdrVgBqaP5XK8feUx+3pkj
QB4tv3ONJ6kvGneEZYI/ayQEB/TlBSR0puB8U3LIP1ANKWUgNKb9cMFlJO4CMV6btzZcmybZSnB7
U220SP851SDxCN52pNkKIg9BaZQWXx/ACmUuIDaonWfqzh8OX2wkst90BjoRjo1jg1GVMJRz+OdO
dogwIRquztBph0HBz5pB07rbRneHd28S/rMLmWUMlM24lHtNszfammcUatoVPG1BSv/wK9lQJ6M8
YajO4++//aUzJCF/lgtrANVNmZR+JWnN9F+5+Ps2KB1mXsbuX2rKJ3oWiE5A5SnzVH9J3b8fQiEp
jcIg/bU/9O/g8rFIkIFGYwk5cQWigp+OiBzTdw9QWvxCinf+px5yTZxoZwN4KRjQ8ZnXab11Ela6
KhE0qKGPoPtSLjr4Ty/mZlNIGcLaaGVL5zCU+FDWJtkuk18pvk0YTp+0+IYIAHdSlFbUrp0Y6l58
Fz4LkhqogtvkLlzuuF5uE+Mbdc46z9I1PQaLdx3Xg7jQXYQik1/SuPOinB/7DulKxCy0CvAylsgz
seqGGfMO6QJ3MxKHvXJlTVKW+AiopaL7cSOcRbftBdO8aarbexClxKHrdaNOZYGDWmBqZaklsh98
tS+62b6LJqw9XjhC4nl6pSKJLIDiILOIH/2+ovHzE9Q4W6UBeYg1qpftYU8be1pQFLIwaNXWSlx0
c52uP1mJLIBXyfXMl8cj9fnwn07fIQFqbBlqgjGu7hmIUATCzAyX54hLYmaIfnTXOoG4bpImJkdl
iNTEoLutMnw3bVWfI6TVAJ/puvVMYrYTPeh8573MPiBczjGyL6/zgWZO9TPeF6mWMjmz8k1m8i/T
wHnmJdOnxMW5c6MBVeS2NWuFHrcqmOG3jdWVf2sqgvBQbwlHvML4qGFLBTJUNucDrLtfUWN+Lrju
R8W6XwGbpL/fXZLdIiLCpfb4BT4bTI/xRbogxAPjfTEH+tYQ0lshx9fHeu97iVBnAqCnnmNrehOq
ta1wTkvTvkwCsgCiD9ggnn09sG+qmIvi4wqZfTcaZVPQpbWSWECP/unEDyR1z0McaerK+TAdpHR2
CF2hltjjG1nTMqtSBbw/75lUH/zSLG61W16v9jdXeTivArwrsNdhFmjGeeIl19SSsza1C/iGGA+A
RLZ1WhhYNo4U1HYsEvIo9YNOJzyQ9p8WlKnDqoHikn++14+W5MOlD93uFucpE/nabmTNJcnum7Qp
nYoYYeVTjl4eG0K2FhxgtXsYUrEtRWYNfU02nyIytZvYXyAkj/gDdoJzcCqSumcpgC6GrH1hylrW
6rPKAaK6+o1vbAZZuQYswhcsnM+SXnGR4GhcRs9uC7TDmz3s/fuu1+GeLgi4TAvfPSvpnjxa0teD
HIZiyKdFZVbuXzSHMjfOHGK2MYhoorYF8VpDs9IjOB2ga7VIvCF792COC4iR6kZgPC9T34qj5CXk
x7WsQ/xWrwvZAiWzdxcJ79L84eKG5Dh7nX9uFRu9cHoqBDfFlyUGu1tvogXohvaCTdtVAZz1e+Nn
xe7GRBberlOOZI4n+HyBFdPH3YAWwNtekw9ckAryj/1N9nXe7HoCAd/KNLY6QMnU+yJkuhDpOfDS
nzTHOEyx6WXiGqam3MfWSRBtea9RUJ1gvtQ/d1Zv7NY48Ew2UXjGtMOj+lTgiOgXkRR8zxRmlo/x
rJeq86ED8FoSQyF5n4o4jlQZTFWQoRa1VitFHrucj4BCK0E05GrvTDxtclxL8r9ARAI4UOSEi5lM
DUq3tZk9BXT9tySOu7r6GGJ+YH/LveEUWbtB9NuOVLyW1x1mHxpcmYJyssqe18K2nIpbSjcNRtD0
Hc9qAszBz41Cj+XlA36IloRihYLUvgRpxUdMmW3ODahdYvdQstA1wMZJHVvvE9nIR+SBWBs4jOwt
dNGLFyIEfXczjsK5jiPnOFlxeHmJpQ0Fk+UnDFdF8IkvrtFiLLuiuCEIA23E9QXRbBA4ehEylhF7
59ymokgpn5QWIsw9WlBjq1Z24aeYtqf+GcVks6eDW0hUj+cKCH22a4YWpwKBh4wZvEc/8MatZLr4
ArpR0Mld+LlaPFDP3ArMcGSjDCIld929IhDu2ABvn8jQIBqoUq9tnUfnDMo93X8zh9c7rMKX2eJq
PxFUz6PH4B0ElvfhznRL6mHwQK3OIhbRleuljFrlag7wZsFAZGChVY0JnAC0QOiuXHI4I8i5oVLt
PEPq7GLYKELQxYPU1b0yBEtaRbGi5xGAmojdpZSTGenLfJCF7BY0RVRP2kPgfh6Qo/soQ8YCnhyP
Dxf9srxcgOJOJio0OCizRi/v9vUosNXqjGaTzCTcoPsD/ilB8KVip9HFvbX6TthlFH6AUT5+eLU4
9XhMF+pU2ElNkrm3lcWwYyQEFQO0AAXAa+9078xdXcaM1ZKVokV7LzlZkDrkuHhtMEhfmwMkHaIZ
23sztsubRuOdYzOi4snc3A+nosHiKEf1Qb4s+FhEe35oCDEB/xTTP+vu0urrX2p/1YBz71tMBT0a
2myvETgnGLzQ64MeFoWD8FwmJtM1eYPZonqgh61eXHhfeHwFop7Od0oeFvsVDkYsqC8JTYvJx6Oq
Zzp9LZTJ68CCu+C6uMgHVf8iHPD7m3+M7qvdylbhpDAyz6STGuUIGeaT4GOCqkE4kO+5kBu6zVkv
ChTcloUD7BFlp5XyhUPmn4v/fP9C4gNoIbViuJIYjcr3NCTZ7z9BtNBc5O/P17r3k9ce75pLu92I
Ad2t3sIk0ykERIytoZ3GaJY8lR61k7G0PmtWq1QTzKNUn/U9QsbQ2sAT6QqhXPL708B3MK3pYDti
fpWFVzaa/nqdA4G4bf638s9wJr05DMMfl6QzjtDvzEKL+kjXVa+vq82h9vtB35JXUqtqvvou7xER
VciyNhPQ+9i7Nj94l5kZK8g9XZFOgDMlkg+kgPgGyx81KR7YHDj9BbJFK6L2Wl0WQlS7c+Gu+mNd
+MkoZeEHdvjcVcsIspP12KRzzBjnPZKquUgq7lx9OR/p+RGEnT5FePz/IifJbHTXL7XSpVAXNfXB
KZCzmXeGZzwcmc2Ba7+HEhodiNxCTjyBsB3XSXPZOqLlUaietqD2R7e1WTI1k2u11uI6F/oLfDHV
AqP2UC1/oal1d+K4I2sdwvmuZWfEBsZjeLPZjvs9XBO3sfkjKS8ul5h5SrA66sXzzcAIJ8Kv+Xob
e8eq6lky/VGr/6lYTooC9lSb2uDV9wIKIMQUpxVU0/59dtInmvWXUxKWq5QzOBJr0sV6RbpTD/ov
gtszmS0dqw3i0jR6lekTE98MDeIldP/jYf5dr2XliqOpaAR7v6+k+NW2KO7O++Y5TJZmhWUKQaLp
dVzKeZaAcNAro2CFLu2Tmy6t0smZGhGlhDld1nYJDANoTBqK7Lc86BO36N4SJ0edvEU=
`protect end_protected
