`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZT7+RCzMGpoBYSuObDu7GHIWP4wbG2z0+NZPy5ctMvSzcpDtYTeVa9Rt2jwWGft47o5EJP3ckUaz
ga/PA8jA7w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nez6Bl347nb6+rwYEAGUgNCAGAzNmFU5MeAC9+3K2UzYt8qxPFrJ/SFJLhvmq05ak2WdPG0DC6DY
KQm2he2dsLt5QsRiFYmj2xAL1KdqCGiHsVFY+u/PuU8GEcfn2GTMt2pBI+06udHlKRy3Gt2+icT+
Rzwp56VKG96Z/MuGTf4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bJ23shOZkE3PVggRHLeGJ2PbG8xrPMkBPZCJ8ZYfdCaWhZ4ZYd1C1zb43X+ojqULL2oHyUgAMgSj
ecIJtiACC+HQhYS9ZAedcNObDtyg4oslk+vfdk+TM2FZF2Etrw/yAEbq1f/PH0Kn+mbNEo33Zwe5
Rm8FZ1wDWOyOXh016tcp0RwCvdj2XR1Kw/zAigz9XUFsy0aJtcUXIJIlKcvvsjSATgFtlJhxEDo0
pnsWRjWP0UYdXkfmSQNXFz8qVRQRGSAtue/7tEuKBK7i+2io/Fn8ReAkkGJiWskeE9nOr9dx+4DE
9tfPWFjj0ZgyCy6JPKhTrEZyje87nH/0x9mcFA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dilSTjuujT5h2DrLDbS/v0rUBHgSqc1odhqH2k0dTfIZcb7N2jGBdTrXFekiehlmoGDjU9sGGdlh
yFg/bT9j8pTdVb3lIkuOyMiLP0CoFYVl1z2IegKN7b9yFR+7EZbxn0N/B1ycLjS4ssnQq+SGbWl2
k2N7LLrQtkLu5td7xjU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pVPXt9t5C8qS/9IP6M6Y37REfDMW0SGfG45oP1DNSuCggimX25Htte0JNMgNJo8ar+6qTjWsopD4
IXOQzxTzbzczkdAIs6+pl9RpNOeJpa0bvybm+uwfWb8+Rcnz3NLflVxnmjLM1ayKKYARNVh7gQb9
C4SQt1FdooQ2JWlTXbp3V2aZpvw5F49u06L9Z5ayEEDdOQE/HQgnVfIryQKYB8stQTSh++L7A6Hi
fnnwsPjJQ2SynIHMSopYLmrhF02KU9HJ3WVKZ+nUrhCKV9djJvyWE9gZFn3X/nfyIkmo23lpYTgC
rYvCI0W4K/uiiwV05xGsCFhMYz37LiZv5/YMUw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8720)
`protect data_block
6Wo5rjfCVuPcU2g0iGcqP/dt+/zYcvdDLKJI5x/fzK0akg8Wb054KDhqA0eCD/jGGam/LDP7pAGQ
GW+/wztIrNMl7c+4j4E8ZCpndF/Az7yoOCGlAPFb+tfkqYdThtyL3Pqww9R/jbu4J8LNCXZshzYk
mApyiYtGEvBYITVGqWl+cmy/KDcIFOy0NJJKCl9WoIOEqfrOpxHhri6AcdncqNL1OGZhvUxgFiXC
KE3q6FNewNx8GCn8mib1LCdckdtj5ua3KXg9inhChVhIxk32BRwX7BhyhHxB/L9X8vHwOWuSLDq2
aqtykyyx7UG5qfwHE2Xj4co6pOpL1FkGkqbrySAtadT0vy+/2cIZp4oesSeruIkVg9KPoYG/MpSj
dosY5GsYoCDtG5/Re0obaTd1CSUmS755VS9qHMDdM5D/sjP+luSE1s29T+cYpgwhtmENOElVsEJd
wTmc+fhAL4VhebIMX27K3XfUkMGDYeH4kZP5uyJ1hupLWpmwiisFPjtwEJ7u346bUYQaWWq679y9
H+WSq21AxPbQHwLSF0tSgEYc+nRs1eWDE49UCY2z+aQOBrr4o4FC3dHmoIONjuJUjry/7xCAmVO8
GyiY6Y1xvaxCMX7kXxux+NErUJSb30eADzc9MWUei0SjFtuEMXPV+p0q87iMKppClZcjeGdM/mJT
fSp5Mg6j1mXvw9/4GRMfrVCz2tGCKsnARCVT06xU9tdkMEBE+5GVzxrUD9+hE9q0luBl4duCy1sa
PDdYr1pfLncWO9uW+OiFMULDaLS7nb/TeHPHH2stosmrM3CjTO2KSXY64T2D85LLKGh71IvdaWTd
gtHWpzNPz/FQgEv6ILLUirAzVjpOzUflgJuMyq00g/fgNzWW2mUJs4I8yc8Ka/jr/lQVt2uiDLIT
gJDfadJ/WRpAFc+Jd/tCdgK1p7Anica+u8ZgRxwLhOdD9vY/+s55zyrbaWrix3z7pb4xm+6sRPQd
8U1XcLMqRFhBmmVuyJYAe4S5AvWew/+bf7kg0L2ng8TmY7gQYl6mD1QmWTTW6jzPlEpb3Pv8f6pg
OxahuvobGoFsCKG06+ARZLus3wCbSgFaC8lu7BIIRU0f7kRTae7OAnGEltKCS++F0EBKxljm4EQM
ixDgSpOQlko02jH+JeIkYA7qDFTZTOshCKf/prw0SyS3f1IvsLk4RNbfegrQk8usMO9NhCF6+24w
lfcmoDiHofpbpH+jl5d9SKgb8lD36JX+3tFIFBE2LXIk15X5ounPizG9x6F7yrnxLeAXKc3I55lZ
1M0YDfybfkWNJZ0+hEL2DCWpnPBq+9oyctHc21Bqims2Jco4oNM8h2hJxK0QQVWwCHLIfXyQ5nar
6h7RklUjNxWAnJiVLpgOMu5pPY3qBIf/E4snmHVgNumrwbT74AyfIdJx7WdunQGvhHJ/vHI6g4o6
pd6WuhIPD4WQNDdD/KM1cxL6aLyQEMQy/6lFUbQnKEzr8lk+zjt/+1n5LhZfgC6pb+sLQPIPbQkl
+/MJihJZ8VNnN3thilkWhU+z+5b0uWmEBs4HYE0lJy8HWuRdj5gLkP/vg1rjBQigtAKg4K2O2xAI
g5BXChQtkHzXFUauDFAxlR0aOtlFT7wrju3i8Sb/1yJGLZq+F7jg1g1jglO1RLp7bZ9L/0t4dMPX
U4/+bZaMqbm8inpyVU7Ow7nCjdeBR3PPG5KCL67QbnJUnYiq078ZRuGVkAKj2zduChZk41fCt4hi
jPWhsn/73NiZ8Yrq/0h8dSjEynUmTT+e3GYVDCU+6r7x10kSkwz+4NXSBg8FmoFmpk1XDiEeTgPN
0SK5MrbdS9vjDOlk/rh9ORNt4Wa0QgKJLGAId5BLJWpiXRjkrNi2FgOV0Y40ehBpcVbQpJNkBTqR
fznk/WqaYRiD0ekUyajcxOpAm2VEFr/BcMj8pukQX8Yc038iexVU4KmFi/cq8mFCLn2nSAWi5FXh
coYx2e+TGKilnzuDaXAA7IQEbC1rYA6BM4dQqgszNhgc8FvjcQWYTmC15Db+s6himzDmt0bhFM8a
owqpxtNKzCrFr3r5+Js9uAZ87zvzYgMxujdpoNZKwqrkJZXdFBqEfwoNTDXGJcAeOiBNArUuLZ3v
PKDUYcz9ZdMbzRCizg3EyUXRQV7XqfldBABKQfkVJEdZGpA2PLW2eDyKvCz5AXtla0r9Mkmrlfgm
Bz1oJhQyQW1dSpxsJALqiUQMmvOaKh6kSsSzIHNfjrvA33xH/AXOCrnGfT0Ylv6sG7oSJoE5A/0e
5F61sEM+xpQaB3kV8Oo7oawaDFsHk17631fSQgQULTrO90KZv3K+UvF+W2Eip/TOITI1ZTMM62nA
FiN02dAC04e9leIzYHjaeQnZQMWq93V4k949ymGCGqH0lKPhGLMwk0inkjDQjkAGjVVtKON+JxjW
z1aAjl1FUUjVyt6PXl6ZFRrGXlQtbrCYQy/JuKnsey7y3Dwr+5t7xr9WbP2MuuhC9I8uNZNc3szP
GR7zpnbUMr8cyhRYQF+eLBOO6oEjBzYDdlRIv3LaHXYKfL/nUQhX0L9tMzC24ntH9kPngREvrDZn
y8M+frT7scrZpnzXShRDMNR/YlJKma7Pb0fSO9g667zWePyIh8ASaQ8Pd+UudPQGcxSG/UvhRdw4
XVdJo3BWWTakUiCO9db5w93I9Y/EwE80G/R5SpJ19isL0oihw2O3XM7fMim6M1RGJhZBZxOgRRJv
bJvb14ql0TH4uTh2ysbvLX5cE/MByRH1UVkkFcVDMyv94gpsohHiuzlc02cvedg7E7r3U/1E/GTO
WYuSbQTk/JvB5lDYTXCmpunYk7Zu7kLkYIGGDxsIumMv3aD8JQ3V9B+aWmttioI3ZgxRH5UDt5Is
6/7+pX2tmiJBel5EuHTs9rIdxKZb/EXprF9ccNl7TnJC5vAUYg1klsWYVmMni1pENgtO2fSkXSOz
n+TWxXZIxFcHQnSdiZ6h47uO9uMrGhT5VZT7IAJrMIPoEbOTj8A2Ym5zw23Lzy5pGJI1hJnin3DL
mEgZfOdxb7mE5nY5vDFYZmhiIPOeql+PQbtDqXjKAkV3ENHtP/n7H7ZtYE4qYu2Qy0jnwPuE0Ozp
A2h3U+q0Lon4rKN2Q/G491yCg4ZiVX8r05icw6XQ2plfKdQZ5q/vjBo0Xz/mMnfG2dH1IfQZAaEh
63Em+oW3R5gNP9O82MkXDiLBgR2uRK7UQuw+aND0LduA5NVMqKy3r26nj4rl3pWXwNt1G1PuImOB
6CGBt76qUqGwjMd6W5Zh/UxNRrbCPas4w/7GXiKNBGBkjFt2T0fo92pJ5dgNna2qyUtexnAR9D+E
2/1vtvHBpAATY59uqgrTfqLtwa0WJWRbcPBzF5YLo7XV6KnFFHwZknpSDP700+ZODzdc0Zn5CLtL
o1UpN0qStOQz0FeUGZh4Y4GlaUUHFh4+UOYPSshJHoBggJLI8EhlS4ovdoic0wfdmTXV+90Ws2nN
ygWwSHgjggpbKlQ0wj3hD3WQX0+GP2rXyjzlSl2WY84CTkNkBJEUlLoJotpJc1KOjhCNFW0SVkHy
gLFiImusfPAMHSNadCoUPEbWcWHPdCrpIhu9LyCPjj5xajlfDLxsamJKJdBxVK9/2AQur2h78Vc1
3nTG41kjxer/sthdkrr2eUEVmXmgu4gg2XQZLxehJjeRAl5uYuGBiJvBQIiaC/PxnemYGPNNgGTB
wAujPb6TbBzyl+SF1rlE49Tm862F7fcJH8CHo0hNMP7zdWsPjjUIo5IrBPPxFHlYH+U5Bvrqx/TT
EfO7TL5fEbdCSEHe3uVjyT6wNw7w5oFAVdZ8LlBSbR17wFrUrDToSK5ZVVGwmQPHcZCRWvyYO+pf
irQ2nH9CQrOFfKBqYQr2kv/nwKL/IuThxY5woIMQYYSHYtgHSjmN1lZx6r/UF7cwz9FlG0o8oCcy
fA9N4c7mihNKhumY7PC/8e5mfBQPQ8SlbtUT3fpgXKToB7qISJoe5SnLYOECkfh4qXPyIBiC6A+w
1FFQCdjxxD0R0qfxBjtcZvFRUoQtXydhHs4KWAyNH7I2Vrqcm6SxHshDeDbJSjOIX3Sudv4EIWMZ
YtQYlEvjRRvgBtI9E2pvnYadQ4rednWtOgSNQdsFjpwXLQClZw313BpQs78a3PxT3hDmZykbjYL7
le1Um0wB03NVNoTZJM92Tb1B/Vgi102YPtl23vvhA63befHEze8Ic9H/dQ+BAX75J8a/aENZGrgl
tpc17S1gbIOyNe/S/8DtQnrV5BMcuIfM7AKyqK2hxURh5lSnAs3dfDAg/lvgm4ecDqcfAivptgyu
DtZbB9hseovi29XHfew86rRw6Uz3Qgyx2BcRxrfHlHlhzLoaKeaZAXxVMQO5gAGCW+zYH/sRDD0L
ye2MIqbdqt068jnU+u2usBYkQfToG5UeRoQEcNaagokPQBSsEd9BU52WZl6BtDDbPqJAETs5xTBt
tjyiqAUwbnx4xKfq6gcYs1JW0w342cUb7QE+Spw539ytUuI0+cbnMoblTHAjTGLE/yaVFJKHwAit
R+cE8aHnZizgxFf1CWDAEIcka9s0GbFvNNA8D9/I7RkDJH7t0RVhP0EShmDdkCxRcYSEj9VE3a1Z
RBzV3fxqDBzXc9CI8yNKJx84Mmtk3G+42FmlEJq4YrU28+5u+0wS94lO8DI2hq2qHoWMyyDjYjdo
bXaCSUkFGp52SPtMUoCEEumP2ksdPA2UEKPxBIWtHsAwneNb2Q497XXBF0WcxE6yBCWbOtplG+J8
79vojzU+kELtmY7fC5qpH1kV4fFhDQCN9euQGwKQAuJegvu8+wFAlPsRUOLUcXPWlFGwnjhqzQmy
O4eXK30KjhZL6W5PP0+KCnjfk0/tenm27CMMcR5hA0mmGGrOnUX4b5Bz6flk/DJ0EfoyOxDIzMkb
TRD4tHgnVxdMjbtolciE6SlJuwGedXGxQIJ9Pm5LdKt57Zk69yca56cqNJ3zb8vIn4hwWzGBVAfg
sXzPVvlxv5zqBgvlk5Sstb8j0yUery9jin08kEWru4+DRNOijVnVB6dcFGpHvQzlc5Z8ZkFEbsQV
m2JYrNksktvBpOw8PQ/foYLMXJ3eAE3+N85Dim/i8XaIlBPuDv9tH3ww9Nd7+B5WPVBnI3cu72my
gOf9kwt4k83rcw6zh2jkvgbRKxoYdrwBy3xSIUAuPue3ykr4T7959egLSKKbCmt+S4LnmsSFZjoQ
k9vp8qM87Pig8EXBJYOZxng7RWmZlyuP0Xfw5XEWymSKmQnIwHfI/pT8484BxdwyHNtefa0KQa0n
FG2R8nA1mHnXTWgxe805nlMpGtCtEWZgLTds8gNXu1/iiq6AA2c6YUKmj8WLn9mTTWImpt6okpnE
VK+KBsFqjSZsBk4KRRyHH3cDRC2quSoYMSyWv3FnRGc4DenY4tBFEMRM+f4tEFEtVcMrV+lXdmoy
adQndFvLM4VpGQ5mNWU806gfmijg6Q/l94rryUnxsFxgLIr/VxBLvB4j33q88TCsZvD3vYH032fO
Xjl59K/eDakhcKgs2rhkZTYTq2PEB0X1HBWNq2WUYf2MaopyNY1tUpvbzUlXNmtizMLhBbZbG+2K
j8+iJkBX8w9dFNkIiVQuuar1NvT4LIy06YQgAqkb6VrIgICQm+F4JFfXFGHRksdOW8YuCYOo+Gu/
+GCM1mLWoXXSWbQZ8YFiu0TlgLv4rJcrSO1u/kJM1wQzsiHNtuls9SQyFQQu5nFWvx0paY1wqgZy
igf57I7VyC8v/Y1qepX3UJRiII423x+g5tHN7JGDB2V5tnFLz83i03zDFoQMHEnVDcxWs5pKco9m
mb617W0Vlhs5SXDZpj/QcgbI5AoUBq0DmWsNmpujV45ItZj/ibpPWTbqCKnQKmM8HXeVoddsgM31
NrHW2/gw73lXWh7k6D/jqp9APBXvYjsQTsbbxmphNYLcedqqZQ6eKR3duA7XiS8Pn5C+dGgwHZQ9
4XhoqV5O04Ip2ZQ/fvQRfpscqyKTuTGL127pt7gDjemSGn8voD+hQ4A59PlIsARRaoyQBK5xe3IN
7if55gHLjlnH/j63v2jUgDrzX2kn4ubME+WH0rYT0nrq24+kCG1lJ7gz8K36a5TPdQZcEbtNb8mo
13Vq/GS0BY+T4wixg1lP6DxBIA2eBjqBOLAXHc6GMchciorJwSd6gBdMOksmtzEdBc9PcWsI8rKn
llYRKUhZPTd/q6ITRUTPH4q5D7q9GW9EXftBtmg+S57+9zX+11wrI3I906gP89NtytxPqqsCWjii
s+zL+VAJuOrTj+Nn6TQJ8ehems5BvqbgAVnwIwft0UdMhE3bZ2CV6nIrpa3vCrkxQqcwHggyIBy/
1ucRI+uPAztAtp9qCh4DXG36HynIJDYdSzsTjrPBNJ69Ga81VOGI+UtMdKudnHlpbU/B2iMHIu9I
0Jcarf6jCA3pR/pb3vaClFQ3wketkLbKEWcT3umESStju/xspbHHhU7y6ExYybhIpnfhKJqsmh1e
4Ygy6HPO+14GjC21DmUwF8M/a3WA5YOxeRj1Eg0NwF0pbladovy2S0p3fl/UuhOz+dGXXhuK0JU/
ggRd4rDq0U77MZduf98fq6YP7MIW0bJ8nzx4GQ+t5PFrT3HBDZCE9nyxbqfaEJWzZ0tzxSpK/xZk
qu5T86KLLrTyB7JENh+5byWhG3aO0/nshzgBULXp3nOL9lIYYElwpEOP9WNdH1owEtG1QoHsZMj6
Ddtd3mMsoWiy734GsZSsIN9a3j6xqoF/k2RFFSCckK3rL4JS5FEiyIC8bNxgA6JG2Zx02cBTtGX/
HtiEB/AnXCrsl8/hzKj6XHYiX9rI7EiwP8veh0/IT3Ox52cC1fgSSYtcG//8QNamyLXbaZ9miV1x
5W0tMjpFwmDedJcRhtNDbcGs3Ao/Jh1WODW/UoQBzA4ryo9vL09096fOrCeW12TEL88J+PNmzT2S
c5ltyT87JPUxR59VzZ8vydAn1SsGSKzPddg2CoAt4e94WZoLO4j1SOb/y/bXyiHIdapJ3qPkwPmL
OdkxXJzV/OVZY722p3SLsOYvRYHk9Y2D/s6Jw2LqH9w57d/aox+2kahiN0c01+ppMDkXUYM4iAIy
ahhoLeO9pbvVQ300h1K9AVpO2J4c7j+fz0uDFShta4eRJbV7NpssTAb3cOXMXpCU7A9vsOg4QIPo
Pco+Tg76lB6UjoSFxVDlIV9WtOWsId2qQoQpzlY+vHnhOadAwx/y2/cAV7OvpkZds+l1940aDXcQ
7mbvUIxZeI+xXvsimsXzufyR+//oPuNdCj0QQtpOOqzc4J4A18xU/Y6v44q1O2aDngjd0I4xZL3d
n01DOF3SMVeLoZqX32zKXZhAWFYS4t4XM45hQKwhMdOpY28/m1rYGnptSFGYPrVwcSbt4Tbj4atC
Ws0cQN4BcJiPbNQ6Imq0NLmOfzX9yMC9jNLSxmAVs/BdUeR3O3gWlE2rPFQ+So3XsQSpxFMtPnIm
EQFLVEHZrpjMzXfcrfxAk8+H09bS5Y1EW7sRAhL2A0WsS3o/i75kou85/9zam+c5CUTrbbnIHymG
hLwdyl2oxXs9FZH0P2uG1o7TL4Db4vdYy8CJpsO5uoxEbb+aKg/q5iphwgfI4G18DgR1RnWHEUye
eLv9jUaPzrld0OWtbbi4d2OMR9nSn0I6T/uyF/4N25+os90KvixO8UnImgQEuK3DTvDV6PMkV4JJ
B+8XzdPoxWVwTDqWW8uC8Uu8GrtKLlXxmT9+U9iZCjAfAmUKzmuj6CrKrEq1CCx5hDZqq7tDWEqk
Qtk5TMZOB6TLI/UEs2STk4RUBfJFOrnkO+Y1LN57wgHESfRDjdv6nZT6S70g1n2e6VtaRCll4rmB
OASEQarG0CU+n7UHpmynUG+/o81wGSSnMM3YwNb/LZgsOYMkHVl9V4WzaPMzLRqvy1c5jva5YgCA
bX0UI9YYarpHJZWCPbSCOGva/J4G3BhnDBkKeY7LthVxKTWgLR2DXI/ShjQGu+TmHc4v1zdMVpSO
LsKebW9WZU8ThMAD4lkTriPcn3zrRomOy+s8ZPMITY3h1tFLP0/5K//yMliHZMz9rxxPBSP23Emc
KAKBZCtQP/iYPFhnKKF8Rxog3YjL5i93sUxu3ZgFJ94aP4KOMfjFYYvNMparzwyAP8lM7q8z0JBv
F6E9CHVZyoqlJNaDYJjwUL4XV2IHwK60SYx8IeV9SNUiSJgSZQ/cMWD0HWsKTu+ha+kiwn6XXU2u
nd8yrXDx9x1woGs2aHauO3/Aa4OKtw2jtuofjAqQ71gB7/IMc77irdkJ+JmcmGYxnRZ7U66eiYam
Rxgsnrw2+boqvtJ1RXytnpBOpSbgVm+nGNu5f/6811AgJ2JlCE+0cK/83ShvRbCXqWlHKz1ZdoNe
qMDqQCkE/VboTOBEkXw1VEmSSMjx+igJGw0pD+t2ekWcJEyefs0I2XEJn4L4UjjZtexvCx9hlBOx
yHIaoGdNrRYHus8mjyzG+fll+GI331BZuoVG8zz9rfsldE5oe5mwCLqnaN/q4OB2GF7dEbWNAouw
CJI0WmgBVN2HQ5wYXWWymPM3FWwF2ZylgPlzLXDGK8CRZh4fmQXEumGtUgdZ5/SswPGg2m5idZbo
DVK+GDFbDECIshL+aa6l1TVU/nBygsdb2GqW6Wh9Dc/LQ8XuWuvbfLlW3PUrLmZ3IbAFcrHIcPSH
A6G4XYo/9Gl0tKzI1ow+8pN1MlPDRBdl9PJxWSsAJEeGAmNPZ1axA0dYaklxwaYZ0AOliF8Ojlzl
INGmDJjcLhZBzHgTk3NJaQ/DiP6GXXJNgZ/heZFNJD7gNKoaT94iuJIykFGNtHVQq20KWCBRzL4D
4lpIeeeTgTC1Tsg6XlF2QbzW58BY7QMEx+7c39cusdEMRtgfw9nGNVCMAGHsduq6QE6juC9jA4OJ
qzJIIRpqSgAj0kCSzYcEV82dYdwVmPZNQwee2/vIgSiB98xe7lctWtVpVD7C4Zf5Z5c7uqo5B1W/
go5ceLMB+1aQr1sBKfVPTtFSHbQBivNUF1I4hM5OvWfqi2YqQwANGtXjTeTpyAWZb8oK8WUtyetj
iuL9j+E46ZutAz+eFPZBYVj47iPhYSUX+Uk+EK5+gIdGEKVYC1a/XfzJrYI+C5qtuhodXTBjGMAp
YrH10xaWbnJ9K+7Hhzq/OxNPkeKv6EVDTZAwTnNqwedaSbbCG16Z776S3qaNt5YrDZq98ell8bJf
z7k9Gui35mY+GeyF4b+nRe9dKnwme6mgcxuaBOURA0vjZqGajrtEMt17CIDWERkhxVOyX+D/lzDn
VwoLn0f8q7A82vVmErN/1RQ/8P9soXVkXac8rpPRYAxD2sKE89D1kbQ+z1p6nThJSA6Ryrjxcy5H
OCgZiJ/iYAZ6DAt7NcK069FVUp6ebox57sWKq/urFZeyUbggmbrE6XIfA92rH/bEbvhN49Ps0/Oq
G/jUFmjPuBgWwmCr1fJ1nGAHFiahCoFpGydw94oRRdSLYnb7KKQIb344OanSOpxJ2orlAkNnF47Z
tV9oViL4XgPVQMD+UmDNFNFVxgKK9zLKEN5044Yv578LVGGPPLzoku6pYki323vCzQ8k7Jq0OEE1
cPLmMcTvTb9MF//SSlX9khxEqt9+NbPFuUURMYwBnSmkraGiNA9wBbavzlaFy5aJfmOUt36lQkcm
647f0Y4GHxwIGxnz3V1pLrofdqEqjbyg5Sag8MjCEnPrwZS7H3X6qnowaupJ7ArH6Ypi1xFzDLFp
gv9/4AmPXJgWIv1KBuVT0pj3dEnjUTFpwGfKDRYm17uiW4fv34XQAkparmVrbgL+ZwYz9tQ/1RIg
DP9pzLAc3BOXZBP5yYeL4b+X4SvJXdWF7SlAAb5guL0Lw/vQ4Y3nzTKET71RxX9XXUuaWyfP7sRv
SXC0XOaot0QuVG/NA5aaxQ1rd+im84t1VvYcYu9Z0z1GvPg8z5+/EvMCrb3cmEbJWUw7Fc+dn8NJ
pqyFlW4a/Is5hZbAPreENzMvYD6npt0zbEzqBKbAhvHs136iTmZqHzRPmqrxAE69g5DPxRPLuYQt
37PixSkh6dDfWn9LMY3srB+nYj4dg/L07X6EYb5V8icFxYh6Euq8cRbVboXC6dgoGNyVR/3VwvBr
hvbPxYY0of0OabwiB6Vm3hgeQTMKFly4o9RQ952oh9Xk+WsVI+qbbg6xLu0XKEnxduttefqRbk+X
faHaF32aHUQo9rOEE7TEnxPFRSH1t97x+LgM0rJzAl9HUzwVgmbmYDrX/xoNteFk9n1owQ0f874n
4StFQk5b8gRC3SKBXC8p1CNW6yWy43VOeoN5oWLQ8Ros3qU3l60Sk4mtPx6GppVYwZqHmGKYCBNz
1BZPQtByzYzgj59IlKTS+XXuu3Ne28NTzytpSMEYRejxTr/oViyAhu6sCbWZPWc9aUMcwQcJHtv+
wishE3pipR9OskaTXjg9XXgoE1SciPjbEBPrOmXx1TV64ntSCocgz91iTx32c7IeFxAr+uqpxtYM
HCWLtTJ0oetU6Te0mc3v0YIbAbgJQWyc79hzynhtoJhSG3w3s03ErRT9kW/ReqacgTQeV7UdOED4
n1MjIrkditCp0r9u7xoiJeR9wjzdt1Q6v0Wf2nasTWebg/eA5SuDfw0UAqGp9v+wNH/tjKIfDp9k
M6f1NYCi1jCkmudzEQCHA3+8oc28F0b0ngOcpeUDdoy9Wp9dN+XCXZmbWCYWm+NK6MYiEUzcRcWI
7hhH+pMlmLZYhagB2MkzPS5g+MD2w4YMIhfOm1edwXH1P8rQwo5MkopwYvLxQ6nR1UcwYfu2fnSx
0agapJMMMJykNIhEy+1+jnA4tzjFKIm5MY1ERB2LjABd9JV5/9wRyBQ9+HwI4M6PwcC+FFEcLzyL
6+bCPyb4cnq6Um4IOn6yxf0Wckk1HkMvJwcf9oZm31PP58PF+1/BXm+hrpIKyXeL5tMVaARB93LA
Eo8LXWsR9rSGBvSVUKVwsiQnVrNfKnT6JjWJNdeP97dCPSlHP9g6q2kZcu+JQwxdSxLU7Fazpvnn
w++LLi+VrlKruvJTvafORd66ff9fRIv0iGZlapNmwOxc0EWrD8gvfVHZZ1nzGhDJfx+PzFB0f1rE
fIqzlSk8M4RwLmT6qVFGaPb22qMUVTDYyLtpY6c0ESyiTjj5JvloThI+VVv9lG0nvHoerlc8TAs3
U3tar4CiEi1H94nk9X/ha1FXOoxUAnF7b4iWEJfb9u46BkcnHNaN+g0JAl0uURk3jQM7ZJ3jkazM
40vtmCF4irkhDGV2+hEB6ZDNLTcZ23bLpV1xA/BVVv8CiP18P8HQGUH6nQIx094qLXlpC387u5ge
hDemZje1n8aiQfX0Q5rmX++K2iYcNEbe0kiOqKNrLiXXLOMj5ZwZh9TTfUtBKBaE8mLH6nKUd8Bc
Stnb/e7noOJL9yOT1p4tlx2Illh/HJ4pbr9mTD9Y4hAIRcKJzSelWf5Qk5O1EcaMJ0grD3RlJRYG
GBuDsDutfI1Isox//1kireI2suU4iKbOGXattZUo5cVNRiRneF5UFL7U0utUlFgs/bcfqyPe4Sw=
`protect end_protected
