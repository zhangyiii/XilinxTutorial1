`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
crsuNbGKr2+HGjsnrWAO3ApjaENLE5lmTkmDpqy6wXOqFQIJnrktoh4R9l/TVlY/BEwSOhFtvEbq
RKvf5np1ZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfoL36fNI5DjzIQX15YYPTK98uQI+Z0aMjl+hiAVWq0lzClrfpDjXWaPyQGiPvnYkkUnnCNmSyGP
qGrNm7GOsjezCGzMgQVr0792OKktWuV2kt0zVP1RUZuHk/37eznwh8N2o5rw+1YzW4dGzl1QbJom
tmB1UpBcp868gDBGaIo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nZKDyxkYA9uy2Xb3FwpEri9edMFM6SqsP4Aed0tRsVeeX445M1QANBu8GOl8sJ4QNxr6T3VU33/s
FK93SNbe96iXZq7rd0ZTftDGFn/wlb+m7r0WSjfp5pkNrLXaYMROFr5Y+cSF68dabG3s3COIhufS
z6LjxtxffkVZFl10/p5NYIyhVlCgj28/qTLowb5EYe1tZ0WPUAxBFuTyFKtX6X8Ha+x+nETiYK6i
PAhbV564AhzWOG1ohxDJJcn/sq1JfdeuDFdYSbNKycH1TqhYGY4rODz7EB10q4+UCVziUOr4Tv4R
NCotWnw5vu+fF2mIxu+vVyyYTSX+rhEfPs2iXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZ2XWhB75BM0Dt/9VMCHTjvBqUtECoyfIkFt8UyDN1IrerieLUkQavGMJnAyOgfgB2F9GkPnzVQV
7H9tsdZ87Y+A3ybRmsawN7gt2tqx/GGsvZlikuuSepi3sHN1vWxch8VpcI/SFn7CnlCh0jupM6VR
707+yLDj5AJkQVyH1LA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S4eCKuneguafnmn96ntdnponlGVTmyJu6zrxyF34ICbqsowM9Vhvgm6poU8XDQ/BrjS+RNPc37Fg
G4CZX64FNy0IB8M93ARmuOVvrGN2bYMf3jNRnVO/z1hOqr23u4iXXLcNjJcX+q+ntygTqDn+dkJa
tNf5JDJd7KcZbafDC5iOu1RcjafQnwlpqyaxuvNRdQkJM7f5tDyB/fmqWMaeSiYSf6cbwC2Jk6x0
7wUP2rAkEzcYQjkJqSGT74QQ9ZxpJuO1xNUbfsJDlmWbSmEyg55J46Q3XRBw9O4UV1TNB2XnSxvt
0rRnDIzS8sn75CDPR31VCmG8K+PwSCayofA3ZA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11888)
`protect data_block
HGwVbJA7sypyD5yh/+WUmYczAUp9Ilw63ul2foAahIAqxWWNlG860q1IJCvcDi+ST5/TvxcuzPir
qt27wGW80Ur84JcU1ohvXeBLj7wUxE4SSH0YZIS2OeLGptmd6Woim7TdjDB1wNiDwHfHGuSA2jrC
ifMC7SRntdZinO1r7CXarWiYPpYWw9HzluLqzIY8u9DvzsQC+rfD4VPTkrV9Ql19KgGDppmRaSTT
+2K/pYRQWW6V3MRdnme7cjQFjSRy23klUwqMpp58rYI9r7XwFFt/XdKcyTBJag8YyVjneyIIFFXE
KJikmd7o/bawp0hKjUXzDgj7O8O5KsM+QmB/rXrShFc6DTET6fHhq2iovhiEDFMLwC2hWLaZxQ+m
qmqlY1zH0k284T8L19prUmtW93MJfJSnScLOR4hgeJBZKugWKEGvViK7MaMh7QNqfJJhc6fgb7TJ
Lj6SVQQKtvyDvpnj8bW1Ln7agI62DiiVIK9V9Hmn25b3I/banczqWWaBBEoDcRoW1AyLKKLhqAuG
AkTqR2iqxJlUn+SNv0XndGq2d6zmmBDGvfdYcRVCgZvC5iREXPH1XRh5+KnbkXUV4KkWm4FY9x9W
+yzBq+vDOOh0kRSrhUXy35dUEt6nyqrgq5ClPCg5ATG5ahk7y2O+PWAAtSu3lHQmvO4eJf9PVRk1
xJ+qNJBjp9qwSVUF0CB5moh204QIyZJbk7GFW4h43NW/QvlittKeHeZ6QioqhMjyZ6siwgeSWg+K
l0UUJa6KJnlEQkAjSv30gg7bcw8kPKay9SLy/71uzoxCJiRB0K8b6a2mP/Zftk9QTJaMMqkxV/Yt
YEa18yrcSOQEbI/UOYdTQlIUjQy+45eXsx/x/8l2ssFV0aJtJsj8F4JrsQyOCSvDap/tBA3FlUGM
udjBHhS17uWDffo7yPMV2sHDwL9UjQErmRRdbBr5Z79wpsRYCEVUY6pPjgyNItR46Nq/RuX7WHiy
XXGTbyrFzPIkWwg380xt+7W9JImCQb/wIeb/anQnRLbKC/q/cL4/+LUl0lccCrfl72JgjJNiCPy2
UhA53ML5prIZNcZ+FdZDeEF7yi7YVFptICpDNUg6Hnfps5EP+couHKX77gJkpNGaw+aZ/0oWYiMf
H0leUvUeTFk8la2hc1NCDmR2pO5HQx5hqrPiI53CWrKa+dI86ZEbQhtfPP9Zs6PlqU85j/q8iTuv
hl2CRFyPOAWS8RvBtoBJwC+UYKb4XM478TjHmU+n0cMEjlxT241GDq+2t2avf2VGclb5FSPhVOY/
QctelLrW1B+pMh2mNMqjeBkGCh+LsvRwNRA5JWXCI0ydPNvk67XtJ+WtBCmQacMEFYure812JzJS
e+s1BeZRTFVaKgcQmvpgt+/6IrOlY7cokILQqUAgF15dop7awKug46pDJE3UYV37pan2Uwf4LtMJ
TXCLDPM+lE2c18Vd4dG81Ecv6w8tduhj6ibAZNKkIIs9J2cctBM7Vq3baFqDgRsaWw7rUsBvX7oi
Koe6uXL6SfU/xItPEXzUAaz+o93/JMrKOkzH7G2+/S2UFc58zz4cTqmEA/mFo2/8uYIa3lmy6XWl
L5Ddb/xBFyBauSLnQAuyFomkTIWwVXKSxGUUqmMT2We62c18TFeC9l1+ZkXkbiFrqLrOVseuUFaK
HJKC4r7ze4EJV8n08wMJPMQQHLccbdUFZbGBbg1fMgtDj+jPucJX5zaUPlkCnHJB59R97R+KnwA2
WYuxD9vbTP8CFmDXcy1auHrvitPOIVcRsZXAPHAbuGW6bZwWiEhRlzDhIZtyd0DDk4MssRbCA4Q5
cNeS3/qM8BdTO3pb+cZYfg4Yf0YLteD2uk7ZZipW2fxmxu1XTEI9YU/wsLWCHG3e626Y2jYur78F
umIokNfX1ExXtUdSDAuArMHPBmrUH9rtIwntuP7CM96UhZsVdd4XMACO6g5+UohdxkMpqnbEY2PZ
/dJkZrTxysSMnYGVHcI/D4grzy1bknVOe4Gd0SgRip/dcghmV1YCWJ2F1+1Dlxyu+pGI3RpKYntG
uENOkzwg2R/47pBUoyIJtk9U51LjrDhXrtpkirrdOsPZIfXZOJmMFQZDIMDqJSvKNRGmwxyvKLzv
3XcGRXg5VBu4BTgqGEeJdu6cPGaZui0rHTUXxD1mTfWVjfIvSdMzsdyYB6pcDEA9X4AWNLgRk1K2
l4Zy3IFwySm0vcZwugVz8ovSn+s0S/hV7nc2Jh1k+QfCpC+pxg4FrEgrdq4KF8hhW0cQk8cBw14/
pjtujB3O0gL2a0WrlnuACx/ItCJz9f691VY3C52L3J9TvBApaHV7w3+dN1zJCobZuSIMUGYEC5KF
UHGrZ48i1nfbMv4rcEYPIFGTg7F2sfW35Kr7+RnTJ/rZV1211cvAbmowEBi8XcwuvI+N1S/bDVPB
65PqSkZlKMfc6z9MTj7+S4en5/dTXmttKjl3RaFJha+17arevaJ1zXmeFSw18ZeGEuqdllwXfhfg
H/5GDzmDTqqhkgDWjSTizg2nSER1TqVBFqkMurA3nDckzYO33G1N4Q3uyVT6UQ03QOZQYZByFLZy
yD5MW+PMYy/uaFLBB+FFy/z5uOAIx6rVXoRc5WFj1lOGGSMl2LSRNViSu2IjlmCaBh3Wxnlqo/7H
YqVJW2OZxuQTODbwlxlbGOAXMI4duw3GhcgCMGjOYPMSzkEZwradpgMBRvXGWjhelmlyggYPzy9x
yvnRujoJcbRMeWu9mEmPVNRAAozskUYv/bZgwxOMHJ08tqsccK32wKyfXWPZ4gn3ja4lmJN/4Fc9
zuHLn5Ia6SeaLXirnqNu9VeV4V9/Ilc+nWG9z/Mzz5cI0hULuNd/Ok/vyRTbSrHHoXxnIi0H8MlC
YcX3s/vEW3xlhFOLqCLYiiF++QLKx84sYn5aseENp1aOXiZcvsytJUWPfxe/fq6IjKMBNAwDWkbM
sxl8pL3kCcZ+RzdEhLUYA96Ya/T9NYc5PsNLLb3EtjhneJjntQIx1zMLauQa8Mo4dOX2pZeKQzgt
0eope1soM/oT90p1X9UnNBYN18YknlwaTUtyyAWAZAe32mpXdihJPvptZqx1AbSjaZuCFQKqg4SU
RaaDxukWX7WlSS0qlNGPZzV40iZRWoaYdIgOcF+RV0/2katM6CNNfLC4Quh+XB2tRD379kTm/Xsl
9PWOBiXF29+93tVd1pm5fapzS4v2d6gXDv7rB7wO47K2t4h/8R1UF3OB+DS1GjLSCOJqCyT4Beje
iRUnv7RuG81vXs0dbder8TW/tqGejMf1xMKtZ32rFALkRghiprIRsiybFku8G+RQ0thNZCO4eL53
Eg/TPNAj7L0UV1WjMzr05nd+QIflSFt2feBoinZiFqL6vQPOSnn7XnQ2FMZW0dvkmEb65RNOBX9/
tyn0rYetkHjGuK0w66vqcQdoLDjEM21n8DcrVSTqpG0Arp4nU2I6T4rt1aoYmG4Y2LX63ieNxfQC
23dPPfIT9zIxPXhhDCTMeITREGZwtqKi9jrbYBObrewQiVRux97d0Ra4LgxH7cnkuM7y/GpxfP2c
SIEo7NKNsbpH0rgnWPqwxj1JiNTKTZ6S1ftCZyTxB8E66ZRRul8BDc1lvXVCjTD5B75fvQklxyFl
ELFQjj3Kv/4xh2lyoVQeJoBXaesJPrw4FQK17fca4vQmtfK/TUPap1Yke4weQZWVo+ii1xc45hRK
TITxDGP1/KK9lWsdmzVV9YFnfjt5ojn7amRHJL3Z6zNS0tAysE9AZGkacZLaxOhbj5CpQ1UXj+q8
ff4Yyy6hYl7AIDY/xkrKWrPpK2fHo5uEvwUjwVnX3hW9yGg3eV62SV8K2DLMFsi5EFZq2jkVmrRe
4St4XsFbvs87m6ffPIySlRDybg2EfORRgHqAB3xi+MfniWJWfEsuXhmkeEDTYU3kme8lPo7fCl03
z8O8mEvASGrZD0cVb0ogkB/yiMMog5KCMnqeUCPjh+VnyUA4Tm+JwoF4AyFFIJZL+2D10yPDIzBv
4X5ltFpMmt2XQNRN3ap4Sn/EcvYxKn/dCV15Vh6bWg0XwSKeq/0b0dM2nVxRiBetlCqFhBmVLWK9
HtlBe7/mt4eG5woz8NHE2amNY+81JIi/+Ll9NxfOhslXcA4NnYRXvXJVijakF2/h3SLFTF05Ch1e
qIqc5rinoGB24njqgOfcJRncczAJUsFTyrk786HHhaz5ZygMwmKbktwp+wUxmiJbCnsx3+EtwjtT
UpLncfH9d2SabcR3tmcdvr4DH2WAVZWb+M4B6NU0KbE0SVb22OUc3xmpK6GfhSYZDSMFmWWp7/sD
zq9cAjl+Kdw8qGsdDSpo+0PkNlaCarpvCyzo1NoxkiJfmckylNJSQtiPGe+ioAF0DZnAFtbTo2og
oNpeILRDykx1q08sqg2eXfOHYA8nQw7d3lb3tWdnEmEXL7nrOQiRINHxmPoSeplS3NHo4lo5BTDJ
tC+HDnbFBUf8NBXCq3el7r/8/9ktcVx9CzlWtPTIlOpjVk64HcyAHqhW8RXuWtoZTifg9atVy+l0
FatLJk98QWg8r0505CNw6SQ55w4MHXhBiW8MhPR9qWE3CqAfSHE9JKQsfVijw80FFDjAOMUF4qU+
ds7DZc/QlkRmvIS1vVX3x5036JlnOnEnUj225J9vmSBz4dpH5JToeXzkj1OkASwp4DHsHr0cWJXY
oUZggDAMr9gXDiWoRjZY9s5+tSFDGl6Y8zg7IL9dHr80U+owUr64IKyjiVeBj96VYACNx4ESQmy+
FciZpkacSfVSa7b5z/Woh8X8xHMa2vm0IUxthBqcM5uCIQ4EnR+ZjYtdH8yVrE695ocxphCSfmQ/
Hp3yj0YtFXbf+t6JAPdmO9DwCssUVl9ncQg9LqWPz1sXP7nizhxXuRf3gZYhqnSbhyVE3MulJVOB
MtfZ7I7g5j4KJU6ZETqGGKL1x7WPMKjjLxJ0xX2TI2LbQRQRiC19+QCLLsDFeORzdA4G69Mkqi5i
oc/3uAGzUfgQhJQa4flikaRyL43AYDmPIU9bhLiYfiBg+PqEUe3iOesbZRG+A5ThqFyVSXysNFyu
u1aWmWoMiVvhjPQ5h/aEV4VijieJLy+jvBKivdRzgovp6l6yDxaiuqaNj6x5pRV69Ug7O78BWoJO
wzOv2tLnZoudxkvcIvZzbpoWbmWOlFrFPF/1nGuNOYe6mWoE03dkgLhvW58pummPTn8JrFvdnWfi
xaaCLOPmMbmuAoTjawv9FgVvpXmEbq7hvM0eQpbYWqyzGsOQI+q0dtAV09EKTbeLPm7is0lQbOkw
Ng6HTlrLdYmCAB1VuV5hcjUeUQdu05Uw64ic1cPNRpewOtqNqx4k9JFfWMAF3duEcsG1ouDNNwrK
mPQpHLGCizV1Nb/X0i+wUUqHiohE10mieIjSLHz/daG8OqbDSIcESiNygum+YcktMY27PPnpBW6j
wP8QFvOvha/xghbKOqHMNEsfDHRtiw6ZLVvpGZ7SRJxm/KdGNIAYsba9oTBpZ+f7ARAYEnTcZ6l0
d12EMR1YX4mK3NFp1zHAV8SZ/vSY4zZsV8H4L9klw+dp3/LIy0IBH5l71HxCsTUWpLMasFSM0eCD
ke8mGta7dXifcnRQtScmxdZBG0hInNS1QCdecvVeOZ0vdeBD6MPNSm0Cz30QohL4at5Kic4phqp3
VIPr/PNXZrFdT6/34WuClXBA/Cake3OsB33UbV3TCOz0SMvrR23ZHvGA7+fjpQ94Q7iChjoSeClq
xKtL81aSegUYxPq3wFNrhhGk02LW3mP+CZFT/yyOWT1xHvEMJHGj2Qoq8lkwB1peRbsqGG7oVcGZ
7NoTP0h9K80a/re8VbJcjDyDgwY8jaqmfWlrJmXfpsRaF/PSxBrSPi9ONsFu1PAJ/frPOAnOJNuN
55nr/MwLZzuX3nhbAbuGLVl4YT+CFmPzDuUKShTnKMhO75f2Q6f/45b/S6/bAbre6ZfOI+1FZNl2
1mldrS3hau+tMgxNvCXv9i1ZfOUSk10Q5eyZOianKPWNCTtNAVnTQ6on8J9m25y4FGquh7B2ErCI
LzjQXPzs3iaH2LlxZX1NhoEyofJsQtMrI2N9NPZ0iVYar9EmAhfBXKY8Yh0jpa7UFLyoHzFNIjiB
97rkAiggMnaNOcCwZXb1fhhXAAbtbWTm/Jf9wexWvLqCGhOGXp7+/Huc5etJwPuR2Pr18IBpctZ7
mhlkkUD4/dML9xp7KdFXiyAsDmFTBFy58ilJi2YuTZs6lyafANHWB+26L9Txx6okSBpy7ozkWhvA
CdPUcSVKIaDmhyG3ZIKkwm6B8lVKw4m6SaDUni4ARsCiklzjAbrqTOJaLFlv8THl9KA+ggQWLHDR
Ewc9ymbGDH7ZOGnJYH4l6BqmmDGqPAMXUSzPC8FKO9qya7oVOMKKiQx33WFTdgFcMlFgvfEa49Hr
orOwQ7wu8r8xqGbdx9VrFor43KZ407RX4N9LXACCZjJHFg/slhbekjdp10rHi58DLlP4yZTVlyVJ
+aF4YDLa1ErAUDX/0r6wH/UX/A2fk6274Ik8RjBrxVw99cIapjga6rEzejBa+xC2GZs+wa0nrRFT
g9pOAS2gRzdJt+3ifpjqEOMF2ldgmhPM6XcLHcycki+y9NYpoKsiYmnkgOhjFQrfV8QTlPwM6Z70
FKBsweewlOggvIAiZFqyc0EtPLAUXVJsu448Qovz34b1vX+47NhfLVbTpPZlo7lK8yDnqugGiAiA
TZwsKZkh4kwxrGh/Wi/KXwJOUJZ0RsqgfAzWapRyjC6kyePp5L99rhMUTQBNb6vL3hg59BkYwXHa
MJM+7DFFDL2tlUP3yx7GOgFP7uSUbxCUy57PZ5IS9eMoWdxjmktzNLBybcUfgPx+/j4ESqqnVYnw
EdaGuB1P7vahOFedQvNfcmFH15SOpqIEdkmiCSuOsrVqjY9s0LvYrxf1wZusXjvooOt4TMY1IaSJ
uHWVKCe2ZN0BBWwCj8Si7n3DKho+b7pqpf9s96WYhuciMEJ3H+0cUti5sCrgcC6Yy9wOPFqm5w2y
iepilQR0m2uk+Yi6b+k/AyDeUvFU6lvv8Q3wU8Z9n3CDELdRW8ZZV8CuVwMA/5uBgJEfh/9ljMM7
+XP0/6LK/5bjImjhIGXguQcbW3JIei3O+HfZZCYYB3om48XT0dWA8FjunZzpeyzv4REJs2a2qnL2
xIp6Umrp4XXdE9wG40u5OJWS3kQmM3L+RGj0GHrb9jzn/Co31nlwXcqEdAOQuh4Yucg7xH/J1fup
JMVOOy6AdQ8DOoONSxCLGayHhP8hAH/rAOCj/ftkEJXbnqcldVut0eN9MbzsGnwb3CQ9bLaN8WL3
NFJZw+nB0StmyHByAjKGLE2NListP48KereuIem/IBNyuTJL2dKjpx+9BH+mbHdHnfen0dfSOdTE
aObJSGq2JkP36ETKaX086w7jyLrO6pTG9zp/d8b964Tb0ULYoJgYTP0QyCwHkCcfFCURlMIeq8Rs
hfCRs2qyFFWe3q8g87TYu6gWDdOIF4y3ic8sHXoCnT+MN7zL5+GQqbK510OOMZl58LLV619A0KGv
mj1YAJ648Xh0omdcx51bDMHhn4wnMgRcu1+HqTsdFUXT2a0/zLON5mrk92mrw4UjC7ejgWYkfrm/
AUvxxT2st96mbLHx1i/z02ADA8OvTAjlpllHsiChVEZLLw6i7PeKQV+GBaTGdfUSwyjJp9amv5VV
6zGWvR5lQgRh9bdRZE/ULhrKsCoBj7EQ9d9Ft3UF5q8m1dTthcH9w1tzJsX5eI4qw0cGP25jAS40
zUfKLnlArG9EuT8eO/c3LpCSFwTlf2y6P4AMpaYSiMFuRDFq/z8zb9+Xcom2MrFHsSU5+WrK7BUc
ZDx8O3U2JZW//fS7Sg1Udrh/8foShgg/RviAn4by3oJyuzx/KB9B8zVXdc+XyL1HH8R2I9zsVnQt
9G+WmxgCsoN/MvrEtJ5E6U0/OujZQJMyyYkMLCyl50ch9DvRzB6RcG7UWaPDLJj2tjQw5b/iCvCh
v96ID6ozmu2cTJJA6/EEfaewapjXmSXY9UcOFRBclo1BwK0C8WF7Gn3n0qx1AEI3nzVdaOTAOQ7O
W2AWwausg+tkw//PJNXewSCjSdeZMRURXJ70GHfiW9x6jdN5TiO68XWlsDG3YEzlwsv9bae5hNIy
LldoGPW4j4mHsAhHScM9qGFLZxhnD7696EwqX/KDQfCPTyv5uE9HdrBgdxrnCLgLElVC2PkZrkNo
3P4FAprKL0lbCRApPfDx5gV6ypMN5HH4NqciEo7iRQ934pQS5md9e61fWhVgx1oWw8VEek9ifYiF
qtDhIJ0IMGt9QrxUfBj2fr57RiySeBp4n+5juiwNP/gGfcprc8PNtLyuBdlZwGDgBi57EnCh8fGj
HSvUeal4ibZyXIqITH3t2C10wl1Ntl5WCj4fovaJV2ROGXrhYuJ1K5zNor3PBNNSGiUIBE+rtb6Y
sRDP1/O+rmC1jsbO4XON4kcOvMj8GgAIIOH2jVuIc7nHjhrBqzKDz30zqF9swD35fnHiNv1LuVbQ
XlgiTOlK3jQR/kTjDwSuatVUh76M9l6iUHXhSCMdp2USXOoBOonx10RxvkNfHnlg+RGBC6WgMMvw
I18uAIfcMVzSAkPdCuVioPjk69Ft+naj+Y8XHYJTn2v1Xhdv8yroaX9GA2YF75iPwN1bRWsYvgev
usWfpyvIM4z2S4SiQDyUjzREclThVm/E9E2wyo9f1GmNwBtgZu4eWvgGQbAjqsyPZOeCKpNxY5as
yGqT1LuxizA10H/nDqCfs5pyjdbvSZ9v7BE335a6HEs2MhExWVIVoH7KJMN0LDetDPhjllGywCrC
UOj0wm12ZQkRj4pGOdWCCYzd1sAjEwr0BchLKWORCtuP8XUs6CHcJHfeCmUXP+gzK/PYwPwNmm92
kBfwsNatYpXD6tn25rH2EsRg0aUIAJIVjoS3JD2YGhmx+GRCkLCxy5VLs/4d0RvHc+BYMHuLevHm
HFW1qMJMzpesrw6pM1KRsI08Cq0DbkaKHzpG7/73ekpa8AyslFQ8JUFTVTnmUwgB6tYeUHoybVo1
sNvKEGhnVgqCsXikUxmnFtTI6blH7gNzxloCjIu7m/Hr7K4U/YRNbibqVjAnzEtMtXoEBe3OyLbd
z/drif9ryHcQThClJqc30wNEiynPrn3iinJPhqXhkmRfSVoXlz3v2v/9XrLvqF0xeuCIJn4+UPc8
V6vgHIRGezkUZV0cQcZs1PRwkyIowmF/nY1YFuB9zpvzoMleNB/JHU/M2z2rNIe4U9BZ8VGY9SSq
DsqzMw/c5xR9UZz+GHK/bslYllPe7xG1lzF1dl955m730iHsJDG1mOjJl+4x/VufKvp6QrNcsK5C
yNQCxts7U8GntyC5uiY9aws5J5v6tXk5/gTD5erLgQTovjP408mXj7M9G+F7+vw27KvPpfs/tYhq
n4P17kx04HX4C9yWF//a7tRR5vGvsm/C+HLBPHohZOJvn7BO076gOd2bzLN2v8MQRH0GBN81NILZ
N7e8fpC6g8WRe0rAsnLXU7uMoKfKOk90731AU7Krs2oA+MId/7id5mi83YTQsJDMIgY9osl3c2Xg
f0Jifavw3hKnImZ5m691wWuH8fKnMZfFl3XETHHuKqfVq7VKXYu5MmMNLu7HKl2Pq3xcyNpjbKc2
IugCUw0WHemmaN6fIoTLcx2S1vgsnVednRF6iqp8pMKDmk4nZpvlYV3pAwTbZ9JeyNkwg4tVOBh5
D3WzVptmljp8OFIc7zBpqr1swebnrc6xF3hJxDf9C5E2ytCY7c3yYSfX1guPDeExXgqoqfhE7OfN
j3dzRM1YGSbFiy56DPo0cbgZre8KKm1+h87h7AtDApYfkpJvhXKMjD3pg4WXnRMBtpypzLU6JDAd
eC3aWF5zkF/MKITsFmriig6nKa8w1MNNPTIW42pCUPs1gJ30yn4VXTLdmaLeapHhJLIoSyFPfXKQ
7VOG5owIQlyXTpJ5iClTj7vp9vcs961wpHanFTyEGQCo+pgskwHnHmjzj9FWOvd2XfBEFxFvzUhZ
Dkr+l/l7ELvolLjHeXkxdi3Ulu3bydYEBybXGNa0wR7o1J4oAhxX0FZ/rEq2wAtwWVWyaSElosGX
tJAvahhjBhJgqC0PaHFa0mPoB3EOMsaIjrl7J5bbRlwpvkSa/S/u5AJ0xEj2YjXbQjZDUXDYDdxB
K2Q4x5xdqY7IJ3ciuyji7iBLwJGc5icFo/90uEH/e1G6VrrN8+NlJASirffPS7BXjDB/be0gaLGf
R+rajktl7oor0z4O3yIXJtNyqtWL33YUupezcJoB8NWv/LLvxU5UZmvnQ7m5xt2O47tAP97WG/x6
LCzQN0V+V+WRa6u2hBn0BUPk+jrBpfrfyiRNW2Ac/FfLtOPmhR3du+P1lKuWJsBRkKxxlgC8P6V7
zeJokhzcbHorIiLWCJlGQvFImrDCHWZ6QZaoLZcRWqK0WDPZbBEmFW5Yf+VmrdY2H2Wu8FOiCRGO
YQlYf4FXBh7Mq5erkBGQ2Y4Vw2gTp87zKcnhA59A0qtbJi8V+WgnLLJGAvfB85q4zMB/OISuxVtn
3IDjFaxnKF+GQ8BqqAv/7t98Qcl3yjfUu2M6dbNc2Fg+QlSPU4L2YXpu7A+JKPLAe04NVdH3UFrO
BP0qkh/LMYqsb/cPCISZEkTdkmhOJd+GJHKBfaEDXTCuxaxWLiF8qm3oQTzmZVV+22AxSjbv6jja
Jky23Lu9NooqSVxPiyftJ0ZeM1ypgHF2nR7393MSZLRuKAuXup6Xh18QC3pOqaXagex/CS3AnY87
MUc7Nd3w2zxy5OEmvsZQTDlFGnyKIVN+X04SFmqzozvnHAdmvs5edsopQd0dPJcSIzW/f1A8Q6Ps
s2NHOcepYw3y+dwLFdlx191ZUiQdEi+ZUL+O6sjEdy3ehNo6FSAijjQk5US6zqv8Y0dJ5z4eBs8a
eyh1iut7TN+Twaqbtt0pO34WWCTzRuvGPiUDO/mPe+yJNM0GUnnxVrhTQI5BHEWR+l8bdJ5gMMMc
uU9dIGOPxqqgQlMILobFDaf+bY9hDi1zWvX4fuUJzSZ76pviGBFzYPxGehChd4JqE0oG/nL6Svqk
nBNiGRHw4x+akx4H7RMUrHzxp9OtaOLv488b/eawMhO61r8iUDkSBJWhcMaS57INvmloCQHmuq1z
BKNHgPsjDEYgZSVQok7qlZ+Tb0UUoGyB6hN/f9cCMdddIzwZ38gj3sqcNi8p7M02y31/leFTDnIa
cydmu5isGiG5NkXEQ9tPTGRU6BL5shNOEgabCGf0d1kUh4b0kCHSiedFcj608uHuxLNl3r/ImxpZ
037Hzh+bkMqOmUXBSUKG5ilHspiL6x6C0hrIVR0nDAizlMJ65ApcEGu5PLy6iC/b5rRQwJNMXKWl
OqB90Q+pQ2jdnXds4TEddhhq0yogU/yq0MfgA6C6fdapcprRDPk7LVQaM5p9Mfdua2YT3eeN92r6
KsGA6Rm8jlxVZ8eid0XqrmNHBEVOUjFpP8pqtOzcoWocFsoSNrQVZ/JP7t8EREU5xH6B7wYm4qHU
ZI8AZDBlgHyWBfKBtCqB/73e/gGYXFw1Rpjm+cy7KPsDQke8qG3pzT3Bd12fErmuwfz8jNg2udAJ
rEnlXTld+DxpHHm5ZVE8NVEF8yYbfbAsZ98oHysz2/tO39pLujoV99ntCU0jhiljtStzwLYy8QHW
9GiI6OjGkvCjOUHon9/+z9hUhH5DJfcmyhIyiW914utK4fkSM/D19taoda1waB+fXZlPryiaqe9Q
rmeXDzhR/VvCJK8kfsn2UMHcldBllSZvU57/B6iT4fVq9IjKDZ8vdHd79YuS6lEokpz4g3zm7zVa
PFsLUyvv9fui/orxAoGrfPZHUyFLFB0ztBX5kR0ByE7A0wenbj/qbXzv6jwtUfke6rYEdkufJiIT
XeX7LVG19wmKeRCgAV5lh1LcSeK+12GiJsdDJhnP6T7+ozkPKhE97l2Ry6O/gG1ZbBO4qwSDUshm
B1Ppv9JjtoCQgSH7zwT8WudOyaRJX6XF4x8GDtZSIdM4ABQNHfHzaupgQpSSQF+ZP4CUyVX9VWKe
DvuuIiwNvhhnJebRmBWYnR4oACYZSSvxDezANJhJnbW+xOrlKGHmPw0+GpYZtlEmARV33a7Nur0I
ixmvC2GxHQVMtZfa1x967CDO9DXJ2Nt0PrdK2MAY8u7Pn80t6jT/mIwpSihVXz242wgDdni5Ekfh
lT3NKhbhfg0Gf1nGY+UNOmhzed6bpIPHGiXfmPMDJuWnLhdlSO1gIMy3d6l6kNDHr+VyimspjiL7
mVyUFzf/wmDou6WSNH1GDZIEp7EU1vuPxLJjLsrkhjg2SQ1v5hjg5Vfup1cVUIDHtqAhBwUF786J
DlElXYi3IhBcO/NKxyE0ITVH03U/c83Qkh/7Id6anqHA4F6tOt+KdCgcCZBp4gf7FTeS+qVTi2hQ
QvEvqYJvkJSCNE0t/WdBoDxmzIc2avBxwW/wmK6ioQoAEmpH0WPEjaWjYoOXo5aJgRfdSd5gEJyh
WQZhhizXgyMjTeCGiT7w0snYg4YMx1AHnbNcGISu6X+eq/U5vKxW3JSFvnZxuuWWPMQXN4Fj9saY
S7XI6iV7XjNHskra9jJ03iC3aTGnFoCVKqaR+Ge+Kjwtj2wCv8Dzmv6E7J/Fj30lm1kfKgWHoxrM
jy/gsqZtEeTB3BS8dP+Da6h+B8JxFVox447lqQ7WgIvb9pIRuVGZFwlMkF/sYKxANk2ceMiRcGj3
NnMNEkNRcN+hfJsurRjTQJEi31Y7BP5FcAs02CPYRjigbhuzB/VxolFU6E07K8BolQtFe9O48JZw
2ugkE3dmCehH7Ocwr3kgszztBeED4CEqqMFHmTuNXDbpXonTehETiqTUWF/L6m2i/oEVWCYPMVY1
kqYyoNvR3jM8NwU8KItbwyJF8faw+9UXvVUQqCYLbe3BQLmf1g/gejFIn+MpyS8Fg2yMWdydPGzx
d2AiXZYsD0nPmuDD+pzZ0Ujz+19z/ztkYWb31BZNOzgS1YSeSCWQZqCfBdtxWtEMF+ORSSpnto7U
Xl6BWHD1++mgpD1rGadiXGhifAuShQs5dVw1X9Mrvn4kLHvOydrZU5ze5ndnpwyzMcYvJ3vqTD45
ajDZ9hJnN2OXMNJ33qn7p4ZwQL+Z8apUHtlyOclONgR1k9B2eT8jSi98hNW7SL41S1V9s2vYmCtD
t8yckcnWd1/pk+yWVwvRXEOgpPzLzYfRGGHe3qsb9okkUv3Y35IKoev9fpVC9wV8/xnPTdi+traA
zNFMkPHH8HY5rLwU0XCi5BE7K1Av/S7dd1bEIJelS6SxMVyr1kklVXJUmg71uNJ9Uc/NgBKeLNbP
nIU72yrzx1iqj96UqGVMdjvYCP077RaMhRIOFd7uBgsSxybz4R5YbzXuNPKTnnoQ8k9TB4mQkb3G
KEHz04EHIfeUJsZwU8hP8emnUrE+/f7dTjCKGQFhS+z+4TUc3/N3Zqgaq3YPdYgDA+jUJRS12BML
aSGxGuiLajjPQV71Kph0xu8gVFzuk28gwL5Ke5H5XASUnDVJkWTv4colVmcyTPux+5Q6OlRXmgQL
QUWnXg7T9+JIxqq8CK9ees9GMagu6gloqS57Dr3JvHtJblV1dZBmvR/2J+axS1IEVhgKB3KKOPrb
0j3mE7AJHOFGiB2hmZsLghDlLqb896V/+GASmOnNX2AdZnGRMnU0ltk8/9Y4rBcs24Jl/i4qiB64
KmmzfXbI3liaEfo/YSvJgAyAj1lzU0HYEEnIr3Ixa5OfFiu2RkgstDvafk0W+iT3BSeIGFhbQ2jP
c2GKuwpLxii2k9T7DCYUyK5e/TyiUoiPxWWiUc5Z637cM54VQLlpLfHHuxr//ddogh2P0t9OtVgL
Oo7tfEhPR3ozErlUufjeXy+66VVdCX1etWVYPT+ogMwgY75acsvk7/1I2mdTGSsrNQ3+yjgH3Ii8
mnTuoI0xwDt3731neicW335vVBfxg/PaKGqNpvHDDgKPf5AG+VgMiQbIgYYzChxJ18WOoxhO5zxp
Fgv1zn61dFr6P2u962StzZ3Wl1VdcIEqAiNCxMMG8pqGZFyAn1fszdJCDVexQF86idNiBZ6aFlkS
Tbdbr4UUBW++CmIfaiBOUoABi3AZkxtv/zvrZ3YBefIOHeAdFLgF9hqb/Ke7VCAn70vqgF1lQ7N6
JOUXw239dLpnOUupyPwpiSsFwZveF6yuROI31J0OHqzF3gg/2Q12NJwBX6Zjuplcp7HlUKAL9Ro4
Z507PwqU01n6WgMQ9kQEvay5ZubODGKypbYFTbELAlDF580XV90VVrTXfOZZ5nu82OnFXqAdwyIh
pCVh2VW4kC6ay942YywLdIolILb0XdItMQP+0YA3PxYKvLwVodICbvcC5G0IJp5TeeZqs7IKvcXb
L3DgHjF0OR+e+dbRG6Sp9QxL3BbmrZXNHPuohXgp6ODyZV2lsMI/WpNHjhjrxlfkIBydRzL1rxLg
0WCDFOHbO3nKVDi+ONzbB7nCz32UtL0YOPKrYVXkl+3ReSXifA9Jp/XnQ3hklj/OyK7QJS269040
bkYPS9t2l7sUI+EIpz1IUTDAxMYaw6/3vNaEbHUJiNuSKpwehpWcvXwFACAEZ+XXX+bWmK6qq82m
l2OWviLv7WXc1SU0SjlrOzYwlU0IfbQvGdr1phdQsCW3EUZ2KrZELruQ5ZJRQj0NtVZtcdJ/q6nf
uKKCyjeERcLua7FXkqUPw3ytxC6ockqAbgyL5GXXQDnOo8X/byPqI+8U2ia+2GXwFXW7DRZAp4Nc
ZXOMKj+HrEA/CGOpcjW7Ij9KV3DWyLQM/QZUxwoR6EhdAlEDcd8O4o6J9rGQSjdDq2iTOHvvKMoG
/uh3x0XEDCPGntjkuadukgy6+LxGjEqUB0h1L7TnNAxFgbZoi4NwpXOMnpx5aOEqSrzWuCl8v/+E
SOF7H3XNyITE8+75B08j4XQLsNXcMmJGeocnLSOtK/FlEm3BKr2uZk7jwsy7Xp1WQsSkGgjQf+1C
VvJBtdFDPa/FkCWm8hu3MOgvkj1ndldhSUJEt1MDGboXueb3HdlpT6bJX1VykPJbgPIiAzofrp2l
JPuaiRMK48gLg9kMGbQsFsFYWwshOsaS47W21aDV0LNy0mrEr5AQiWKVKjREuRpWf5vVcxhku5Uo
8Xohhyr8FX7MptKJlvy2ZPHtsYE/uwnw28WR+0iZEkNrtnknaaUi5qBwf+Iwu12Gw8XThwkv6OfM
lKl3W+Fs7TmbTWduCQxpHy7rn/iXwAlguCJvThJleWBWgqmD14nNHj67vMXmOqQIJErlVDt9EGLy
L+9krZGNRsJ9QB1iVi5JfGw0SV68fqk71afpF2sSTNm/UMtDx0sGjrp8HddFFoxCDuZPI5LEKt/l
/jpdGdgvKBKwKcCWGQZaIMRA3owW+3Zm2IA7mTdFTtPH/rZVgwJLJhvmhvagCVWp+hNTEb7BWuIN
hiGBofk5NrMWxN42iMurPGh3/shQMEbr9vSE2HIFrO2YJSes9bVkh7Xs2+7PAuBuEXvoJLi8eHgh
1QGTKizrEcq6TjinlUoO2NEPLFiEFNoOKYFXZlBpfoylGAqIKwgq1BImcUMEE0uZ/e+v8cY8jG1d
Arz7u3ijFKsaatAcyob3Gb05PIR5GbKqRYK9nJtCEp0+aZnAxHv553R8o+M9FUx9PrYXBdxn4CRX
SrvoM3nXwWXTEj1v3XE8Kp/xV95onV3Ce4fq+WhlOLg=
`protect end_protected
