`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jNvGKMNtWEUNKagzcg2Z6WIUWv9gWJV7my4RvssH/ux/cX8RktigUyw+RYrzrXJGrNW7g1x/nBwF
74yzP41Y4A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cve4pj2EfLuhqfhnGnOz5iUJuIGWUldTY5TKWZtU1S3TPZ4r9ymlKXit4YnjR9S0JtAX1GoFuudL
h/jZOj05rTC9CmxzpO6a4qp621eKZhXdyOHyWMf8jPXE24P9V+aRttTL8nXifMfo/UFfsvRfUHHL
a0V7II16UbNY0z/aQ74=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FK+UvGaeunWTo0SP2EhgyPGTZaNb+A6fyrB0Pb4mabhgLBujusE/NHHToooQsIrVtG+iA4L6uoFa
xZk2qbFfIXLgeHkE73Jf9tkvOVSfNHKkwE4Tk/zJ3hux51whzpeHeM/jgYHXV/AGxAjK7wYmqNEp
cavJsaWgLnwe3yjG331MbcwzkmgERAfcBrC1i6iTT7oe42Z8bgt2QuADWtJa6+y6yzc95b43/J72
7JqV+DovmhlKbNR1biVaDlEMoR8wVeDr0xj6PecXn0O/DCkFw3POXJoaMT+xrRj1LksGsCY+qMlG
IfvdA3kKCxIRZxGcAPvET4wf6cGXK4CAVBa7IA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
z2wDansBNwtedB12HDIWNrI0jJ9Of4AnAAv+qKssr7e7NujivlJDkMFVu15DOLNgNtFvyO0niOHn
/kdDAjIwQtt+ugBkFsRzbHtzg25iwcWgxIDasTP9xLaasNHS5B2OfeSNk+sAZRujgTnv16OLLpuj
xCVg+ocyScQyJTN2fY0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dHaEE44368Lqz+gkjyTg7OMF1sLix1urvVlzCGNFKkIp5zxC5Hb5ei+82XYKqaRz661xkzrxnXIz
CLpQVXEZh1wM12r8fA1f5G/ZuHgSsoz7RWoNbHd4G2GQJUG7WVKCnogPJmbAQZpXthW3KW14NIsi
E34leEwjyTjx/frRrPczvVKGoZSH0tKOZiCD2ER5SRLpYvlTJUkcUEXx3CipAjm/wVGV6SSyQJeO
CTF45Rt8GOFQIMhL/GO7xMB3lpMvQg6M9+8i4GbdQOAk3MmCg7nCiIL/ptz2eDE+txQ7xQlXt4Cv
Iz7BX+6KUqHhfTCrqRi9bRB7HwJgifi1MzfmqA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14208)
`protect data_block
dBSVDAWiIsOQDtztSiCUKR3HLs/5iSD8Ul+4l8GtKXiMuBaQmgXwjEfrqHVcXssRVfUJauoA9C/s
YcK/Ggp1hrdr1QY6TSUUGSNg1rqOGLqhHmTpDGkpCcnPuuoAQP4UK+u895eDDUSuWWQjDlFvoO46
rtkOUQQWyeZM4Ocu9OwwVwizQviNxBvZPYNI3kEwIbFp/SPz+cY8+kx3p8++6GV7rrZfkSy+qrVe
/aTpyVeEY1rtesXLIYgkJqLO+/uZVSQnTVIEbC1VVAG1JfAGFxpu3DBL5bfnu0VZmOrGBgokb7WU
DXpUPTc5cSfJ9Kaxal/nHrPQKoNldOLihS+3d/fjirGxQcs+lXkUDfuaJ9KWLuggD+UOHo6y7kKT
DyHWOTNcjtjtTridrou4cQ4GMuLcCmRDlPNnFyIa1Myq0zmYpmujMixtXTNUYM8FKKV5cWS59FEI
aDtXlzfRork85KTWtNmrWDD5PbsufsVdVan85nM4GJ+sMDVGj4ZDwLx/PUX6ZovYfAuozqOpgqve
TgCSLIRrbKmBslcA6XUm2qnx7uZB3z03198nuD/n3mi+qyU5n/tbW8OiP9bEDV1m7pzgxVttJUgZ
H220Vix1Dd5Ju7fq1EeOzhfGnfWjMt2Qd6Yq9KTRO1AfH9qYPBRAg97Ktvns7manT2A8hOeuWieW
IbUkb8GXqN/MmRohrDS+cHUeN141kC7jk0FMhkeS+cL1Vn8b3GPFJ25gxMmMBFqJV5Cb+WR+BiiL
zKWO7CFrYgqI1/+riD2oiyWf8rSuthiw+EVaUKYhAg1bF+lR5blFBTmifLCNwW1fiDbVURNARWOM
Vx6ZcOjvXNBAsFGLWGfibWdpmU6/EB7uYXDPfDZDtlhjq3QS0dTAB22oVWXRp4SPt81AZLvHimnd
J4l2m4pcAICQ+lZ7xwFly3X+3SJFZbW0IeZ7Z/LQJ64atsQHUxbQ1el5tzML3UafvOv0UIDYdCdI
zMhqS7BDMb1upg2VNPBVmUFs79LyBMV2aSanCJtF7hPrUIcNPoRYCpdXDIE1hVXyatixzrRp4o2V
2El8NIy9tEURXyohBJAVBjaCdldPTx+4QdzrEJK+Ewd1/CCKwEp/7fEQIp4XPI37ExXsiqbT0RGu
m8hNVkNUv8aaQ+MHCSjkntqhpeMlvtTYr6X9kQvN4GjXqA2IGym+PS0zbVoSXmCENTmapcLChG0/
0wUwxL6aw+RWJ9HopezSr0EF1Z+bdUARnt1jhs+69fNm1mrTprY6HlA22WKUD3kJXzFAJYL29sx/
WcBUBp6KmDgq6nprBMcrSTMwBtdVfXrZhnIc2qwzjCW3ncgSEXlJ/365ZYlhOS5WBcNTZaqDNOlp
ZGYOcZeT4/5TAjNSU5axw1QTqMPrnPHOK8OpU3pWN/1EmIhR8KB1Lx/jOEkEhszA2KsFZ4KEp0re
4OwCJ2IaO8JZGjanOjggX506TMRV3InDMwATmK/dqWQVSjIVDChJhF196NHnwWjIDXVh6GJ0eg6y
fxvm8yIRPLtFFXC6Cuo+lj3utRnDUjVG+0AjiiO4v+Hmfwpx3+6G5UbADL4RPT+cX326S4JQQRYJ
mSTuuKwAYancGi7GK9T7qRbkSIXIlreo/BdZP809BrCEV0MwWntKJt1V29bsja1X1CrMJu1qmwhu
BZPHufiusdsjt0BkvgFY2Ee4eDMieX+POUvmbV8Bdt8WF1zQpfEvDGj/8JpCvF8Ijd5LnVtsgZxN
J8PG8Pk9kgQbgYI24qDzFehmZ2BTKk5h2E2QEGONRNXkYoQ6Vge9zhf6AB3vViATHAbnRhEBhyGR
vHPFOEWu0muo0nj99yaewfgxReNrnB6Fe74HQtQb6+hJWSo/wZq29DYLB7spULTf0sJzHo0tKKGh
jgd8kbnTJeTlscZh3zgYW4qMNWzpf+3ndbig1o1uUX+/KSjH46yt1IhoBbjbqPYTTTHKKXQIl8AM
g4NLBr5vaZs3SHHDea/At8X8HwuomzUaLBzOtQRwW4pwdNI4haeugnziTHeEfB68QpIc/ngZvvDv
ZfTb2HPcflwZvguO4YslVwXBoi0+OMkzZJkgZALoIq4vFKKHYw9i59j4XzJtXJgETvmiW2hiSOZi
TOKdrD0Po1xGT8yMgtzLHT7ski/tZsu0dhkNuIKDIr77fYEq31F8Aq1Ov9zL2EFVEvtg/+xrShCj
3phRWGXen/vdfoRPx/NIR6IzAsxEI4MEyyrJbH6DL2oud1FLEA3N3Jmo/CMndAouTppF0WZGZ4wl
l1u0yNfQIG68JlVu7ZmCv/KZ89n5uIn+c2cwqE9leBZTSAt4U4g48DMSojI6dfgoaGxHOWpIOBJi
p4RhqSahxXuEQrVbBxMut8vbk3/xUWGF9qBgMnuDDC44+0WXxhBcMMfcyylLbF9kIjCJVBCV96d1
wua9LLBlKNj9n2hYKvw+CpXID2Zk+rR2xyqj9aQ+2gEYEY95BS2YvyjNiPllyzF7muST+oO+vA/a
qYuVBprzMsFKLdBcbcob0nDrgW5hVRTL3O3z9RjmjmB8V7FWSZ3r341gmyTfNXcYfiGvDYpXfEuc
UN65LdN0ronfOvrbKnnLaP7Eplz7cn+LCKc8OXZpzZQ8Rai5qquLwcpnV0G5F180gwAYD57TcGxi
YaxYHQnZ1QoXTS+a+7QBeCKU1BeEnfKvriKpm+vezSJW+vil/LWTmZvD6KvJugvHZo74iD5qteSb
Do/gYQHLnxHAFSwfWTG04sR4YupaHjDDDrqq37fxy1R/zTT5nyvVsg5GBjrraj/HAmxtv8pYIPVn
ZmA9Ldz/wUKNwpKKCun7FhKvCxXNO3uj24a98RwtGBrqfnfWGqc333R5qDC0DOTSFX8O3ugCwSWl
B6gtR02XzwO5pNwqEqtiDv6yAd21cX+wp29TDJeTcShtqVGRoOjvGGY159FsZPUgd+nIC/nb8YQc
Agz/iGOmy2HnlPoT325y+dWbsITC2mXtZJKm6q+WfSB8/9CQHFidH7y7KIj6GHPRP4TPyQNGivz/
KSuNktHotZ0m92p0zq0l+FRqi+cGLcRVwV6d4ZAA0IgT82iOhsAaFKitHfkuhi1N+9LWfUO8mIdG
GF3Cp7MGMZDlkjaHZJjrKgj5SMNZy/QZ+k37hQ90GnEy9c+kWhclrZGMcAj8xUN1QQ+kuxlWCkVh
AxWHYwcHivlR8im6fA0BrIkpEkCy7DdtqH7nOrmXIwRnczNEES/qsb0jUhZffIo5a+ubvGjLe+f6
qawVlaHn7VLar0rITsbyCvWfSoNcjuaT/zK+3qEDAHmDxOdWxJMxyeO8wBFH6yL4jH3UCT7TbuaV
TjsiAEx3u40Z88VQp3lSAQMTkGzSkEqIUdMAFNJQAL0NV6SsYXnYDzH1JGJjZgGlt2KWvbCLCeBL
wchNwmnNIPq3D2D1k8YFSxaswYgqP+U7kBbWQD7u1idZqPuVxTrmSn493ySdbA79P/JL2JdKR9uj
Qndv/eHC3JrqZef8QrLiJ0hfX/VL8px1uB9m9AY+OOM+iTmMQI58JJbHCA2fvD4bXxi1fcEZutVD
6A4lJxBq0I2DLb3pSdKkdaNVf85YQkAqSSil0/KDjd/QBnO09v4yS2YfkWo5q1C6N7j7554o/LhG
PNsRkcMuT2jfWIk8y52+qOeP8nLjX8nWGaLc14q6okH3yiwvLVh/cwuc9esEinMkv4TIUHdMLOsq
OrrcYYzEiYnZBl50x1/sQeevuKSQR2eF9apLv8uWry7sLz86G8EoWzsoxxblTnBhB1mpHVvGQS8Y
A6QPNB7jaylTCaF/CyqpT86pBCAZDs9B23jllzGY1R0apB2CqL7nUTTcFs1QgRdll9SHH09cN/lv
QgCQQ+jyndiexJh0BOqichAbNRt4EfEqgbClIssC+eGPoB08Bn8eNOm7SxJgD287RyLlHP53kOVm
g/bP6R90sYlogALMaZr8Khb3QVfFgHAJj/C4GLUG81ivS4KnOO5xuE1KwJT7zjptAD0ZSdeXVyfU
har+ACR6XFBVsqMQBQoEuOlvfzee8VoNFFSu5+gEleKLsC/P9ppxw/WcBFRsxCs9bbUQ0ap65XSq
cTa3Zv3fMN9zDgQ6HMCLlItTcFzhzdJxJddEYQwTdWgBQvgdGGOCfiFVw7VdFdPg77AVn2f0XeYO
YqRoB2+I1XBmgjDKj0j291KsHddX9J/bfHzv4+nXFMoiH3BgP+AfKwmFl874876wWBVrB79Z3HFU
+DKRCEcLER8cEpy8nbvYYQ+KoNhck82JTYUQBJPLHzFcAEbLL908+MFnfjEU+qWVxBXWbg5f/n5m
RLrrEOVIbnN+moiNz/+E1XZWqb2uN6SUGXZKnoZFwtyiEpx6UhywM/u1w5Bu+2UK3Q/NkbMtODSp
JzBQPKOBCbd+z/Q4Iizdila+oCXAGFmh2U5SnojU+x3Sh3EC2ajSMrRI7WyjCY6jbWdJHUk8og9H
V63qBFAgJ9/aLDdMXOa1omsFLz5IYOzdtSprTdth7nIEN0cN5tWNf8CwFrxEw8xUfEtac20icWCO
iczpkz0ZUjuxIYf5eU4oWc46hFkeDOsbEdC+C4/p9mSMAXH44Qxwhw8iC4Y/JP+SWIHJ2zMiJwoA
7GWrIuS0+3rIthBLbEGll8e6eRUvDUE2YgYV62qkjdEkrLmX8VFp50AUKvql3A45VZfTqmgZwVFl
b1lh6fYnw9ps/2TWPcTiMTTs0irN9TAArT83gn6a7PUU7btd9ac5u3/lKefkM7Ki8iXNgui9PgSc
HepxPvpovuyWj289dVTkHftoUJhzKLq/Og7AVqQBDyAipojpY7UXkk2ZI4cHlGsUHWYtlwRnKU7c
GVGcwhyX1HLHDmp0OV9dg15K01GgsHvRUHWQ6532mQQ0OTHsiohXUTzmGH10khWhjzASPrEF/VBG
GDdRlvIu14+5EsQ575w5ObTTIDajw2fndB1hlBFXmlBPCY1L5NdTknF4+E2NUK+NOxSBlvp9R1uY
00TySx+kOU0nMdW2Y/BjHP++fyTGZPDI4sXdrlo3lrx/2TFtrQbskZBzL/KSuxkO0dwIasoBq0eH
7mL1SSnNPs73vkMMVyPE1HLhIPvCBGPX6AxXc8YmpFujkGT8Z9cYilBslYgh7qX/ReISsC78f46V
SMtD69+al/9awuULSB6FDXsodI0QZo9iXMB3YnLzCwxk4GIH9Oz0ci61mxhq6qGeTPQOGffAAYLj
FYKdEVoxho9fy1zUwPUiilkl8PbnUI2N+2/MqMibSeyASHXkKhFE4uFX+L3nTLVMQpT1G2XMQEkP
SzdoRDTpPHOPLSI8QJ6LtDURCiK2YhFtWrm/oO1luFXVUpQ2LTNMLUpIjaMwrt1EEgo9d+hKNuU5
HZ5JjhUFuIDaed8BjXeLxGAuCSfD/EjPOyS/JFbf2grluZ6vIQn+Q8cp2MOFdlJUjMngtdVfodUW
WtiDW/zeqqg7M2+pHFAbY5es76Zk2oz6NDL6TDBANO/Up6glaoyDof3wttWYj1Zpdy23s93EudyL
e1ii8lhkZGf58aBNSwuUroBMauVPrKIZG5oQ/Fo9ew50IwQMtIrFx1FNSAgmHARkESj+G4J7bL+B
rxPYmlosbUceFwrfsAdY33G6p1jIMXasPph4HSVUnJbFyWLFCSieA6wwUjYz0CPy9Jxn5mgek2/I
jSqXLMYylvO9C0vpv3cAGclXhAJdS6vtK5bocTaSjw6KMNG4JSfThUGXB8SykM/D1fXjUd0ACgRg
BGeMy+jYIgYeboXm3onH7Y1lzATLJcxiKRD6WIG/RIpe3Qxnx2Ug7yo/97/rrqFsH/zoZeypPyKC
S1AEZ4TEcz5jhSsHfXZOFlCzZhJ2rCufyXurWLNxiezmeXW/ONKWygx4qIrruDRf7JMWN21ncAKf
AlyqxrSvccll2vBVwsaAa+vs9EE91ByyQ3sUAottGmTs+bJaUuauJRb2pw8hdf7lxfoNBy90hhdv
YeWb9aMdPdY8wDyp25H2MgKm+tWyTG/bvSSmQ3oNb6VZ/6g1hFEGolVY0dAtPXhmJ3XHbsUxh182
PIYAdNj2pLkMaEWe/70scN1RmwcQCaJAtN7rEDet0+Fl+/1dZUgY1jIaq+FvOa8R3KxhTjJ0sRax
4zYjYzuAy8PFlTxEp0tcWJcjxHQyPh69Nz2X/60snJhDxLR9/RXwwa8pB84DlwOxv6ajAMc8jO2F
P9QfvviDOqZ62U45K4pVGsopgj2XtuZ/iKnMNEbf0BGZX46/LffvSTC1MdrJrNNgex5eOzXAth+R
qucB+Vv2I2kEYMctSNzwIYO/lRephSa0vfGCLUS+uE+NRZgvzyGchhBymaEQzUcw4edKwLepDPrO
F1PauiWD08Fl9vMOGD+fWvQG4srcH4b1+p1zCat7T4/bl5gRSZYnEPptonn4moQA7a7ZpD0SyUu3
/2h4g/VxJ7ioQSeX7rcJeZjmrgXbrTC2enXKXRl/Aj+txTSCU2/s+WMhTlTTohcOwiJZ/UeDP+Va
iWYMTQ310+rSeQrSoHsQZFb3FUbjCQZthi/goffVDLSoqXwjIiCL6c++qYY7OEhoiCqldgoqFY6I
u4JznZjRA3+e+8BMCzq6ZinTf4uVufRIB8Mwc+1acYETflMHExMTwEbsoHhjXgXWcv8Eeiidyc3L
psXuAlVQXu5pe/556nVIjS4Gvu7Emil/Rx3T/Ej5CB2wF1xjv8XEVPQ0BpjwT7dEoCLqyzST3TXS
A50fTrzq8KWr+so7RDPmZ/mc5f6jvXQL5zGoMmU2jCkclVf2MIcFa1ZIzWqn3Sp1kp6oWKbMEwsZ
QDZaXGRyn0KJUaFEGmfvuIiUzR3xY84VPszFniysUiJKSbYAxwUGFbWl+a/SEvu86Ur7jfa/fl6E
U8bZNBVjv19fonS4Da5wGwSAh4T3OVkLo0XvZdo1q7+I9Qb3opoBdZz1gjMd6N052ENbdZbsir18
sboADf+mIsOIUGbrMu48gtQcMXdDEPOHMWyLUgbVZfKbAyPUDMOOxd39h5D8dGFmRT7L+snLUzuG
iMsgpBm1ioAYaP2O0UGplIBJ2yHgBNI91TZeNiSal7u3FE/e0ipao7mnRPHEgW0WxV3jnCNgY+KG
0wcHqWUKzb1Yd3OiDtD/pGeDPeJmPGImLRwRdDMW8tR2mMQ1uDrns0d3dwIYb/Crd+MmiuLG1qWK
qtuMYnlo0l+kyJpJeT56EThtM9hz+dmDdJUMwh2kE9PUc66gHhwaPPWBfm5FZgPpVGwL7bNFE3YH
zXCkfWB0Quh/nVVyPVZq6S2oUQ0quIlrqVwEbWjT7aTYdpB+gRjt/iYk+MlPrRQtJVq/hSgP0tew
htcTrsesk2/XNk10awRAqDE8zYFJrQEeXWv/Iw/0dlaHeXm7nb3rrMXCEvNVv5k04BRkKEil/HBe
9oQLAbiRugSAH3tcH4sVhxwfme+dSH3tEMr9+HOz28KdxuS0JoX9YjnuTRR+xw+DE3Zz4Whx8w1M
C7RY4pmTauonyb10D2clldIRoROxEfYHP9LjU+1RHO+LbWE47eNae606YDLxySQooUB0px2nRCM4
T6oV4QyM3LDvX5+uI9R2Vl5IA6sZmGXv3fiRM6aRe/PuCkWu0GqW8fEtnFX/4PEauaumZpy5zJOb
lfU2u1IYXYHMvCGzlzmC6hrBoMHBUUUJtojkvhUV0DNRIzMTZfy2BKs/74PrQv+vLP3HXLVN71Pi
opmIWyR2ZK3h79CXezi1ckuqBMRbI9cq5VEtnRCLtc8YPwC9pYQv83m4gg8fm3NrkPJX/Bg1c3G/
eFruVeEEdbal7vvjv5ESO5tXRaudBREYt3w54ytNBnOwUOs+5RCCgEVBZu3YePTaWK7x3lEGPgpe
IUGOwh8TqtIW5YSHxWQKIuJuPu9NFZwjoNsm3GY27bMMYgRaVYZFX6lwITh8DRHHGu/45EBwX3Zz
bV+7tvMLztA3O+5JtBuqJnhv1X8muADL8/WTjKkwql3y47TvxVoDaDZa1Q3gGqGvQKDNFSccG1lL
FqFc7EB2fYiMh3GXZZDgynhnpyUT+6Q1TsAGaKh3wEoH+EFfMdOyAjmuNMgwOQgWtM7rTKi2Ztjb
edq80H/Gefk9E2WuEiZCe58aDCIN3fo3478Mtr/tymsXLdcgJlXUQNe5SoiVG4wCyWsxn0ai7vz/
bn1M7md5oO4iu+ANplL22aDybvex9NfoJ6lMoQARxqFaPF0Xy9B3N/FvmGeXdxAyBIYUg1vX/F7X
nbNblNDrt/76oB6zoa3M93i77otZBe9GUqbE0gc6nHp3hlIA684Ygwbu8e8lJ7WJjou4KoIiEwtF
UEReezVx+FFOWO3zQZHmOxTR8zk2kLfBSsjVKy7miaPwNu415GGmEssnUP0CuSsdB1X34SOe6OSZ
3i1LmqN5U0ZAom2bNXXqGMMG61mudITZ4fuBXioiJ39K63lcLcoh6aiTyQSnmPDOTcP+g/uMr/a+
R6+RN5lm8BRxmYigCLsHvkA6LIic2hcjdNUMYAGLvVjk2NA4OIJB2iHZXW5S2HuzB0qXH49APwfY
aW2LTQuTia+byVgz0ah48iY8RCnTutOA+1stW6VcujE7s5XT9pT2VHIHJeuwv1IPcZtIC/HEvLHq
AHsqjLNIHGPW3uBiQj04Z09oG2q1SWttnHHmlxh3aRS7Fp/htCaAqAuTOX0qZiM0aG6jv2BMb3TD
1Efay0+B8uBRncUkvzlQ6EONBuc7bDZA5f3znd51dur2sWG9VPo1jT+IfBe0wHV2699J3alQb+CB
BFJ2SWdghjpIti0h01qbSaficlub37B+tXQUVpvICSlssVqxRJXjrKvADAw/ftBKtCT7U9IpxkT8
0RpKSqwmRCK2XeYglUvihoMZr1kpNZg+F1E6nNJps49VTlLZNLl5g6mP8+/cOGEmKNoU95RQGssH
tF1FP4PvS1G4S27KBPa2ueccLznHvu24yrZHn4hRVTgST8OkRLqPcGpPD1ZdUqQkvOsm4tKfpzzi
4ug2xhMGDWl2/2apBofZk9dV+vz2/mMHcFTf+wOvCs7au0gXBtlIlFemfekbpzCHTPPs6R+Hl3A4
whbEY2iarsFrFnE2Y4ikc3JzWn0rt2yPfYOQ++LLtTBLgbINOqyooEIaPzSRvk4y3XeNjZ/nteQ5
14of6ifHnWh6nTTKyPlyFSkbvQ3DMseFd2loFxk5ySSFjC2inoL3fLxgUdjuOd7G2Qvn8Bf7JTd1
1REDOC66tgBoD4CA8R0fdh9Yx7lKWp9I2ezok70xciDSR+R1FaKz9U0uYSEPvtAZj9aJL7JTRwLB
/poJKb8CCRIflO7kLpH7uSLYaKTT9kJYVZf88aSRYKpeFtGfNwCbvXX7aSdmXZx6NT4YmyAVvsyT
94Zj/EtlhA/eK+ksXFrHA/MxaF82u5Gdehmw9XI4FYIcWepBikM+nw1pCXEI7fwJ5kA/M+QFYRf5
omoeDitMKR4M7z1c+Wg1Upzrl7LtS3yFKdWz7r9OtrBH1/bvpgWiCJJqR0MPTYZ/p6grm8py/CYX
kCDWaR87B49uRO2XAsxyExJhBRGe3QvXiScToVziyw5xUS3bjF5Sf1qR+0WFEvaFK3rChinJQAcs
gOox3S7I73AbDrkx3OSdTagR6vl2ahhh/MlYMzaP+DmTTfiWXsC67/6amEOG9v9rA0RZIJ7KiorK
GK/vWtlhXAXcTahHvWiEwSuJyaN+odl53EEFaSLLWufHb1McgGUjdCgLwbwKYRheEcz0OjNg++CU
41yzzCdWp6Ru29f+6vR3K7opN7AeO76OdIGrOGwUzeDd15OjjwoG3x6GlpY66OPpW39mE1yADjs4
sgvSbFedLhX1LHm1id05ry6xi7WXbJ8YUCyTJWmyxyUeuDmDHteQ9zT1gGnLvA2O/+b2I1H53Q4V
5clPwNKyJTttzADuiV66eMNhYnvTO3jhgGEmyQm+H5bmW1XNCyDnJ3fjpdtatBUPhyIbnIaFSTaC
2njcJPgB6Mq10Q/wMwRFYwz3xRfkkc7JYqWKBMNWW1TOU0PNKcdHyda0WtbCYL7upSezN8UMVWjv
BktVelEIdKbAqvXbDkbL/RpGUQvxm2qV7+fahDCnCrcm4XweTsulbfVUTP1XOwcaf7gNdHIW4tX5
+9gFdWIuGa8DN0SI2gaeJGwB9s/b/bA3WPJu1zNgWZT8/3f556TlOMBgAl9MMuuYqY3bmguOag4X
YoOLFnepTm+RaLpnBlYDoeRrz0tJvJPSSJrzCMLPC7BmIG3BZJaT7Dlr72Y76iuQyF4R37IWeTlG
r0OoxO70UDMm+mZZf7E/hh9RaLTBczluu1Thc//9GvxKuHp31ipk0VPPsLQRJ+9u0J6mBgd1PUa3
g3ttzQW5aJrkHZcVFeNfogb8VaC8T3kMPAKMTpATFg8Y1t8mk8xlyo/NEEYyxI7OSpR7pwJA/zMt
rAUhRmcSfgpmHxyuyaJbwqIQqSpV9ozLfeYb8/sH5JTgLFw70kQDhJY8cJ6w3muF6zbboNmVzkp8
/9NfUxRCPVPiI1s5JLJaGL1KU4sGcMEU3pXlq0mw4wVBeonwZ0/eWQ2wEMxRD3yTLeI9BiKfU/k5
wyrqH1rxmeztuyyoRHXLxH9bu7dSwE06XnS8mcY4ymwogmQQmK1Lm8od7cb5NoD3wKN/GbkUKrgM
+CyV9KO6Ue0hnIp4u6Ng1S+xLGvVJ6GtHfy8KykQ/V8nlGy9v4jFAzP3n9jtZzPSJt9Q+nnbYMpD
3U3qpncvb6vSHnN+0sqTNTGl6K+rj5QNJFWGzDdprCwHrr7d8AlVc5yYHpYqtS8CV/WYQ0AcTv5f
AoalNZJLRzSAmzQA8aMBVGa6nWU29omOGBTINK00pY4mxuTJ+ZR/B7NqBA10emUcHJ80VZPqWkQB
axHzzHcxKZzPEAFoMKnd1J1/dUsy4sZ+y6rSq0f4fp9M5xKrjvUBr9N7Y8GYvpae8ALtiubd9Gl2
a/WzMPS8SnUj7geUZcjf/RZlzwPnQeXG5wbNoZaZUiydxMilOoZBVtnbwOlirfhqoOMJiTMuiiJ1
cGA3ugR1E/mhaSjF9Cgg/7HdsZhM7gfZ+aFnGICq3HzlCVDBSeG+YPMlqAQjq49c4Xi+CrfUgPP2
UCRKsqw3wUeRHXJxjuMJnG3yjiDfEJUCoYLS2WFbrm56tQalcD0ZUbVGwi89FqotrPI0nM8YQrQv
ppKgC4IEDsAwtKJvEKu8X8ZG5rL7Z1ihIhwSEQ6yPWtAdSQEnepwP4PRwMnTQGvzcUvadbY6IyuJ
q4bZrXxGV+yg1kEMYzUmXCojHs0vaimZR0Q7AwQIK4Js+6zUbRa+bTpqkWKVutBmmrNc7NUmpr82
65LdacS9NQ0kwjwFpr7thoXNXeC66OQRm0vJEEr+jMeAh75nBwStARK7dyRxL61Pn5YbCmbEv9hz
Px0quBYyZsd+P1toT4m/Ofdv0hC2JtlswRkgLHovEnso93RI9tiE6R4sXyHbU/b/f0korcfxVz1K
dWzKwYtwiUG6FumSR253IA8LIzWawIqMeyu8eVlXstnu5s8VaRM1uB1fn97MJEO/TyT7aISru0Z0
XaaPx/rqNll7kq9MLLJVmRTURbtKzWKlwqn3SKnKZTDMZSlOq1T9/XOUcFpstOYIFH0ahmelU2HE
iLJ0CUgE2VmqR24kiMYEIgIdfRck4SNweoFsxgLBXgcovCywx/mQUECp3Mp0KzyVKW327y6vkk1C
lNLZMoyqXb153x6AzntRfDfJ9pxtZhlyzKBi+LAOh1RzNiqU2x2a6SVtyEP/VBvua0g/sKwqpN+K
QWccETbR7mpjt0JKX4Q44KhaEFj4R/RYXFLYXrL8KX3E/nKvW6vMZlV8OqwsCge/RgdPI8C150MW
IqbJGnSyD/c6vAmOgB7hYsMW4BRb0rnBDX/uQa4MgLuAeWf7+V7ALWhBzgFzJ9QtvZQh427fIjLw
Zb6G0weI0t50JBnH9Z+jA7neZVWaqgs5DgCrA9X/QLF1PftK0403q6uDBvgN8j2VW5vb+FV1IHKU
apkPSQciy20Ll++6um0VPVi1ux1b3pJQWl3L+xuNc4bvBXPcN6li1yGnwPrckCgPXW8PqdiFmLro
C/YsL7aZen2BLGKC7zOwmx8KJZZz86Ab0KaBDC4i+EV4ZzAR3ZAMnugxg9uPi1GAO2Ry4RPvKsNF
YHYVQPbD0lxrxN2Ns42KXV07kdk89U3Eehku7eSi28LrCWPfBG/Hc34FE2LGgdp4oowAHp+b+T4i
8NCee6w3nKccCxOd/gNatdX00pTYYhOqI12Y0FtDmAWmjDtjhyOtvxtKD4YhQXzlIc2310/BMZ63
Hjp1sR5g23jhY6+iJThxtvup5PI11QMPri2wgAfmTuxzo2qqMfOphaCiYzLNuwBFTWVrGf//qW+H
MoVBQeOvo7Pjvc4Et0fCm0bmm+ZMiXtbYB6J71QcUVyHHzLvXdyMruMT8LekC/4ES30RzDmU3v9x
PW2Z4lvXmFdetp6RRTR8uX1o1twKPKs9B0pLsND5id5SJG1gG+1Bc20oxIs+wV7XICvr0bq8aH/t
DMMK5FBcG2sWFgl8RR5OH//QDN6pXxnuTurXZBgE7pMrpCQTiX1YGZo1Razs/ZgdXpfKxwprLhpb
DUQ9CoTpKYsFHT+izjtAf6s+1xLTnGCiR7+czz9CAj5jjXnK+volhqy/BioTpfbwWWCw50/OCnYu
II3bIQwyjicB2N9SlOaF6zBHddDmsB7RCL11KL/w9JhLGBU/uInbLlD1npNBJdiG4ak7Gun6GTon
E8mHi1fQnmzsbEUYEPEh/fsHY6QfejutBxp8vHTCgfZnzz2hMnVzXByEMdtxZ0c/Dlmq0PE3i8xd
sJojaylW4ko8ACtGG+Pl282gpH4N5MDiWIGKO39ZMV/7OiDJJPUWrsC1GZa8pSq71e0weTqacmZz
qZpQC4Aw0/Y2/HyEcjIyyLlUzogF4pilnUdFmFacpldpqQNZjSNDPnVoGg70m7xBAzxC5nOxuf++
fz6aVsI/ZOWF1IdzpZHDgbSG5i2YBq70rWU45mfMtuadorw7EaEtNef2xAhrAoFYgcahDEF4nohP
paunU346HSM6P3P0YQABfajyU1Mo26lttRI0Nm1hEwJl0HNh/PnltiDY4FzNnMN3V9d/wLlzn1PI
P5rfj4GrRSHIdvrJfc2TsvvI7uW8zf7ALeSuhwBV32idb1RUer2sZ+pSjtek6NtuBMPrJkrznby6
ZOxbLG2YOs3j7hOASHshuZLhnsS8rtzEkf0fLnB2Gx2LtlWFFLfdcoEhhBgkJi4LvKRVR9edxDjA
Wh4jGeXoeL2S1v0Y4Qs99TLgbfzzX2HY/+IOmAXg3QVDp+xHvjJsS7ZxTZ8BwA2XlFGdrXhlWhbO
vQEhmBtFCntvKd7Se9wlzsxcKjukoz3kiursHz5f8OTmZLRs5/39rsrNM+pdBwZODdRzWAzlmCiU
4kg7UI+W+588pz4Y2POZMEkpoRh65ST3Q1Ie/+SjbXzSIo10qHPX7XZJePv8NXvjatxCjh9dn7yH
gG51KtOoKo4Ruq8drjMEBUk169Ug34C92FyG7nfREWrK/BxCcKr1tDus/y5OEfaoD/2JmKUmHJPH
p1mIcTnClWIxSVUBH2zR4BrC3IBBBEcd3gO9ZyrdoEWyKSR+y2Q5X3grnwB/elwRpm30b9NsnhLt
+Nnsbu94Amp2KrF1xDYGgdUkOJGwmZqqn3OdHd2d9GL/A+iD1QCNcinNKu+NnNIiCBsPC199YSYU
lnZI2cV71ihrRHh4nUlEDDPcDECV5RQoJnHJ9Obkr/VexV3YiJpflcN1dwXVVYvYFuzw+1J1goUd
MS8j6GDOBIW9fdV2ihEYsuiwlWhHSHOXn4tldQOjVxFDSdSkbEt+cDAX+GYKuQEeQfd3ZaMCFJSv
SWDpZGxg2Z2raSYRhV0reQx8eZbvP3tZfvXAd2G7zKkKPAbF5KqjeYV46tAnoPz+I0kv4SaOeN3k
0tVBr73DeG32cEEHM6oNk8UckPZHvnN+DZTfthK1purmduwe4IMQTQZCbLt21Dh3L/8aZLjTa/Jp
maTRt/8eiZ8qIkZTgU100uSIDJCrrRRWL87JeLi5NPN544hTMf/gL8lrsrUEIicI/gPGG3PgoY1i
Qt+fTTcyb157imypVt/vpeyM58wLHCeYkHmbIlubN6QllH3FmG9aIr0humgZbwxYjNDK2D2hVk9H
ZBudBqqwfDr7R8uYWF7my0wglz3X6P79cR5Usb9mRkOfhW16aDrRsOICBu/dQCk/jsCGnq3rWKxg
oO4dnaQM0ODOOOk/JwZYJEwR5Uf23g1TLS9RoQuFkaX8p+bZf9TeEK9ewEOjro7SA71TkK4hJRWX
KCPhazsJvD2c7ddZYoAqBCx9Au7Cv7Wya/lt7PH161o8ZGXHDcGSITNiAIUC3qUqygUyKA7djsQD
G7d4Dl0OLxJkCbl9z4lmoxss6S8oASwyRY46oCw9hnC4/vY5vcQIGgC/bCWgtHQEX/MBEWGWIF6J
76wU1JpIbNBMQ1TVWBVYcgdn1AmwaJt2O4Fpk69GY2H0OZeUTTE7gSDt2lVNonQjm0pwKvmzcxjC
fEvgzayyVgkN9NOY7s+qAXefB4cTfbAIGvKKmMcxLZV0uh9CIhyxjHDiW17QllHQwlMVU/V8UFbJ
RdteJh/50rYu2uP9AoGELLbQfN8OeA1/T34F/wO1DgVhc+gBMu8cb6mIK8gQt8Pw5fmtjBzf+gUf
HXxG8O+d4bLp1Jzte9KBKavrPLH+nZfP6zT/wEp8nYzYY6qcwLaxhgxgxqSQHo4VpIu3eX3B5fc3
UGa/qK+aPuz533LuNklZZS8RLPNMnaL0+4E9kuH2aMCd689cCE2mtprbWU2IIvkc8xDsuMb2noa3
muxGowbRMMrJB3ya4mLtNMl/UniYomDbeV2zAkdx69CXsG1SzDXrHyyk74Onhz9d7DkOQ0TH4IEe
U9Nz4S9VEnh5YapOEVlQrM/Gge+BynQF/t1d2YgQuUxDRF2wVi+ohyA3bR7yF2Fuef/56R49f1FX
PbcFM0qvGmqO52/ZVcSB8No0SX/GK2UIEKu4N+kvIqyTqnwDKgmFODFdLEeQYIAgTxu6mBIRzbMr
QfApHrGcuQVQkZXgWg161jbmrhIqwEflxeFFT7dXO33IMds/4X2or1LlrfLODgqERIQ92YwYFYlp
87BEbL5UNMkJ+OWZm/gUnBO90qncftpKmxqg144GMhZE22KsHkoPho0mqGcMWc2QzuDyQPcS6gxa
TbL8O88XvtaVnvMErSYq7NPX/+2vAUu6FYwETjPpiWxiebuv+IzBh4/im2eN8Pf8SmnvGjCZZacV
5HSi5FCTWXiJUmLRE47LyyUnefBRZDWiLduXN3R4O1Y0wm9kAk85vy0Zoo0pQ7WhMaHtL8ae/5Eg
j7lXFSncQrg8srCpj2JSRMWyG/2dMqM42XOPrRX1Jcat4y+r5bsC+NInLOIZZ6FaFHxKH3sTBHnY
gzdnQG7rKnL3LhMmhQT3SGMyXD5SGJiyqa63TK64l2M5Lwx3IL0LvKS7J7F7FcftPwS6OY0QFXrM
S0GvqkgLqJkp+yP744bNLkkGs7WkciMldOISW5Voed8qbyLu4p7BDE4njbfvLpylzN1188HVQUdn
VykHdxVYhouK5pWQDvtdkkO8KIzbTbyu5IEETUfEBRdHMvlOpOGK5CxtNWVig1HLqCKjkFFyBbAy
37C+/AiqKs2f/7+h5yjtD79FZtPZ6yaD8QLr8gB/VhDfcWi2uIrdOSY0HGZ4yfrYO8LeLJELgBfS
de5OFGEOiKwdrlRSb7NFisHn/A4Gqd1VGYEIWLy2dvt24yFIFFdeYNeFLOS3VCXb8PH9kBFNg0Dk
+WzAv29P+z+oVQ2YUzddLg9uujXFH+K745XQjiLXNXmRDkM239hYNXzOAL6x2KBuVIc5Mh8M1XDc
AZyRdowuvDIFPtoOjZcZGTHHl9Gp5hqrtpeeIIPT8PvuSP54Eh2e7SqGZ5WpfILQUHvK7Hof9zC3
LRbk4fY/XaAYC3XHeNLVEL3O2gZXZ5Ye/6uda2ptBTypJ1htSJ3HqduHQmkkYRtBqEdxCmbCutkI
oYJYeyM4r+aBUGmnzq0gKBiemeuHLGbvYDv3cHT6DFjZHzMuDWhlUeeXmYC1cu17PFTvYk/oOgWd
A1k8/FCWRGTOdb/a/u/mmxOmnyBieQgS8Zg5ux0WnzI6muPXPyNvm4USjoIOCGasxHbDNzKj9Kl3
MStRPGwWyuBQLSeeS1ZMSTPwSNPrpDKCcbdZ63/pGu/GPObS9fWKjUJmCDh2d9y9hK02HuKZvcrV
4a5qIvlRf4YGHMnpVLSNx+gEB9aTY3Igoe9+PP66+NaykZpVF307SrhygrWQJW1t+8A92rUw8U1B
diSUS0XPcLP2seiU1v1hSuNf90zT2X2P6zlnCIxRsee4AXAyBEzix6WSHfpbs1u7gZqqKzw9uT5T
bEe4q4M9JF2zodVu0aCKYfMWpkJ4qDIqj3T92AAFJ95UPQi+B4j7ZmVBGHUnwDWc2vKRJ6s1dOjz
Lkps7dtiwpqpkK0RiTl2GKUJbZpkk+om42vbRoaZ8E9VLDDjR32o0ID9Tn3gAJKLeGpb6k8aP5P8
3qdP2fC2+51EidUO/tFqFUkN47Y1kYS9akd34aizykW78m9ioFo1ktxMboQYlsj5cb514M1uwcBm
KImQ/3Y1WO+iGpQ0S4bj8iFSfe8EVirdZDh8gZmY7zHsBz2Ddbirosei4sQa9m/5n+C9FRYNAAcE
OlNGqE1A3AdWkw33+Sl9uh6G4dUlQj/RZYZ/kPnd4d2mrEVI08aV/0OvjxIuOV0LLqHbz7Je7iDz
JMLqnPGe/mEx0Vs6Gpqdoq+FkeI/9ZA9qG+aIn7ZTEaFT2QqUSXuGpP4Nv57y4QnuuYDvYazHZRp
SeangpU/nuqWETlM2tR7ozcdqpXacNX+HdONq7glkqHC6KPQ8ZTII+RWNY64epZo+r8NhOJ4cem1
VHdUXUPF/NwnjWv/m+Dl2SyWK5CQlLzCCgvn6XlWhuvvnM3jpC3DjNo5VPOB2hf3SVb3hP3J+WVC
hKZAlWA5ehm+1hKwL9iLE955GTqc9vSuOlmt0qhvhxXa70k/n/c1GBpzH/HiavwLu7EwzUl5ZzXD
IIP+goZnM6YDI0qDn7sqjvMzW/zKmzdbgqOrJa/kpxIrlk+rKHY/tyWB+ScNLhThFF2didc26lCC
0CkPDD+GXqyMyHKtHXhNaTsoW6Aoo86EEkZDuta/bAwi3WSbxo8o382MJuv7NKQC+AVSF8iiXxGt
EnSjP6+B7bnQ4XGe7NNGEwS46lGa1Mu9ZzIJJMJuCNPnkrKP7Il+xqcCtPBkpHq8fLib+b8wNRxq
qMUN97ZleQn042IJmvTPIvb8mOXjOpaBS6ZGR04s//OQCSKGxojz2QYEctvmTF3HaJvDrpF+RyZh
uVeNHrM3N8dXqwLhPOgffe3ftSZnfejf0DXU52S5VsCETZuBwZADWzoy1VNPzUzsyv8y3/U3rkWo
k4S2OyoP2yyd/rtZ43chGAvmuqUhb7VQzfY8N3fCk779BEbIFRT1899JKUJ9P/kq7nU01XGgd7n6
tc7mPhlWsA66iWOJZBoZv4ECD8UmvHv7OT92du3DGK3MIJjnVZhhRfXVQoBuM0RzM8X9ovqNG/Mo
FByHtZtu7tpDYTbPRjCdoNWoPZx8bbldk3XFPyPRsbuZdeGBoxvwwNPu0kbtOBj3AbfAZj6nIe5u
sjPIbTgH8qfqZH5NZroMUPwKDo5Lr+UGxXaCUWfRGsQdq6DbG9QGOG5WwMVpRffivfBuwZ0t3S4t
H85MjsJeu9WkmWlq+cxP4SdTyzQSZ9dlA5JRijJ6ywkuvGs7ymO2NjggmeLdZO2IlAG/xmHnlJgm
FLMLEWchkLwiSN2XpkEAxhezRltLOohL6F0mOU5HxgTX1pTnW6aCSUoC6vzo+LQjQbnda6jdrDsJ
M6Ot/eB1dfqyEmQvcu0gczJ/zxKra951butybheIo0IYOjNXfjRulMiBIfxd7iIRj+qYlUW0D7ar
qRhhipm8DV7VZcZf4ZMGLHSBT9DkIkSB+Ez6v9Vxbx+GJjbCAtFU52IY7UhXaY7wFvcy1QKzMI5c
XdhVDcFwqDzfztKSQuIhd8zT+7y7WLuo3VJI7g3JYIkrvUIhKGi26UPcmbUl8mvJ+C6ImStcWW6D
iT5+5dev3diJnCmXfiN0IroXSSYbp7AYUrA3ulD2fbxgJ/8edNq+/3r8wmtN6icz8JKlP1vCczvn
5vJEOhUggjtApI6OheDqsoUntXFr1rWPCGy2WkDKMIK807yaSMTNOkwvmfOgLjR5NtZ7EHB4+/JI
ZILWl1sXYE9K6SXCWQwa2FjfLcZIuTnpmdZrgyQfbgY7z3hXOcf7YAToNQuZTzsyI5O+9MiM7bka
emhq4oILwfHB+LOkR2YjcmGktHA0HOHy/kLzG8iYwMi0vRqlWMERELf4qZ7Meys2N5GvqKWsHZJl
hTQQFhycuz2rF4J/h3ed8YWd27xnni9wmR9eNAM+74kRONsyWzdJ5wVc6iQDksqR1gqAiJzKj03O
NFjvgW+U4wgI/QW60KEz2I0LMVKzXJbSVOEUw8xbe90nnn9nalJwmLk02BSyLkBJwjDVuDf7JyU+
vgmxjfg/Gr6e9vy9669PreKG1LmX9JutfBDHbI0+MAZdNqRmk52AqO5K7weMTH+fK4mBIoFj0MVc
oE5cazTx6HvCTMMqiM+FRj4TjCIKnoBtYT5M9fh/gatCdVjBZcRse0gF1V0oKb6NcczjVbLCXWES
HbffMck/weo8Io3s+SO5
`protect end_protected
