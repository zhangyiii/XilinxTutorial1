`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45152)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aPkk/LZprZljgyNzZTGF6gcxBz
LkEl/7f+3dcASD/i/KjOQr8a/fv4/JgFmu/jpTurJnqQGicyJIWJv/Fz27LYYmvHoRCkOGUkLqLp
51FhcmORyH0ErTiypVzJy3jsR2PtzmL8HZbfymaplrY0MWw31+7fszk2SydpGwkBeo7ZHfxrfZmG
asogOHza2J1qyBSgIdmClafB2XfopWgviC9L/MYTgY4Q9cWwugIV16oNnEcbRNla3Yfa2ljj8m6Z
QLTgvNl1wfOh6EOVKykDaTAaSOUKHRDz2JmR+JdnsOm7+JEwfgmo7LO2lmGxH/0Vq9VOlDjr2KEG
6IqAUx+lUzHAg6pgF8BB5RmQpuO/RhNfJRi+i6VI/5JCeY7HAIpDgStxpVwHKqa9yzcC92OWaqk4
ko1ADgTbpupB+yo+JWU80SdCbmPGwDXXeUzQERCuiK8SRWuuWf65Y9Qe5r3RJmJDmvDe4hj+4Av6
oP0bNp7LqZO1HAWCH2ALmKBHuRaQCwgpgJvW4vUnwUqMjGIhOOsookvgurYOoyHyIswRDTTgD+YO
USMZPmp5iZmiEG+HcZPbJV380+KgwqP/qk9DN1ESvsjWE0XOex/8oc5DqfPnIFMvkyDLB5E+ErC6
E4jijtEVpaVMKA0hNYxhBnYbLKgPg9sQS38tcYxWFMMKMl/5w5fLbh1wThYD9MTtXbRzc3od2SjV
DaHa+i9sj/TSKpmy/GXR/45sDg7uKtATd0we70psq0ohf1cQRGVx9kp58EC/OGoHCOUnsocjwPkV
gIh0TeeiIjzd2IpIvXaCTenXAwxOD+cU3XH4XSZMDDazdb1vg4Fr3yf8dszouFpnKFNoTP8J7tkw
E7vob4MhN7UgD3Y7N4KKgnSjVu6O7zYaGIeQnp0+Xw9ZwOK871a6zze1suAPnudB505cqbvsy8VD
Q2CvCDjDTHofZ1eUXMVuA9kVictuYJ2jP6R0Il+r8Sw9tZHyQJfCdqCGD9pTNRQC+l0Ba7SRoWhS
toDlUNZEzR8owc06dnriuzRUcDnl6//fa9XxjRYfO/GYSMz4K2gHQgnHCS4iLDjLrKnnekki7xBq
Oqo3pxGjLbDwigUofHesKgkxBk0W2TOpdBgnRfUeepUlIUpoDX7kHNWKNnO2Ugt/2KSugfDFDyBy
YEtALNffpvQtm0ahqV7SLXu6wWrsGZePChWwVCo/4J0MgUJdc80NZZY+zuKg/dIfPDDHTI8uNzYA
mpYYqXTHiDmqawZkKWPcy3yqaAoxJvb79prePAXgjv7omHkOGVDow4lQUzLVNvPZPQo2yXca/2LT
msYqOh5iz0UGuUrPc6wUfZhWmeCzkdk3bEbqv1hhmvFwaanShML1Vmhf5egpbaimiP4S4eLt1rKC
ZB4jSImcpvzadZ28VhpSuqhpAiJAY28Cr/yA0ZXyy92RbDDl4kyNoxyMjrNAUSMe8EdwleHlnhl+
tlVL+yfrPWZbI6tT8RIh+ulj/UwsJt4wus5DESf3Y63yzQpcbRdcEHky93TL9IoWUix+7LkwjgnS
eNyCYMtufxjuItd7DRmmWdLOEWZYBiwvfObm3k1vQW6SqAYrqRDvddhz8szuVehWoAZkks3FUzSu
BylWUeJaDWRVDmRYFptoD3lIK5rOTtUMsWmVvoDAgwnCBQjkxJwjeHXYOoVR327YlhasU1dhaUrU
HE4Abo9zyIVYcMvsyALtSgDuN3ImR/VqV2fFCZ0UjVLcgcbrQ/m0D8FSEPJNHzooevoonpBENIqs
Xaxc8XXWe3LHXIrQcemrPxnyLFSsDU5P+JtVXc4+qc6LlYXTJRkCqt/OmUMK2h/6sbtDInmJDrrW
5XSR+zQsN1XC/2v+36vG4ZICYU3s0cg5XgcNWEiekdAHaQy/OVTdFPeFRTWJQQRpgEF8M0y3jsrX
XVV11cVcAZI3KFB5Qetqj9279OQverDMmtr2ALrhwOMb9gNuepFRY63PcyMN1S4iz/DGa9cETrTu
i6CHDnnZEJmtz4+KBlNG8Px8Zq/lnjqTj8igsNYFl7bKTWVvLqz1f5/CUK8lVNx3mtONtoxWXEu6
lVCpwh7juEd5goSKJ3HdvIg2SB2U9W+KjMfFdbwjxrpXfvUf2SYHV/dE8QGJ5LLcAoAFmNttSEFQ
8pd/CpK0L64shnhYyycC4r7JUxS1JptVnp64JKXaZ9bDVhYOtNZ7WbHS2gLoStpVovSx3woHf5j7
vxsOS1KZvH+Fp2+AYtOFWqyV92ma6KK/bHBnlwgv8PG+3LxvTiwo+xJ37vb5dESnHoSvfXWvV9RS
FneL9JRhKoLMXGnRClf06631HjodFu/bAuqJTUZuzEAEMDwd9iPNwzyzcoej+dC9rtV0PApeYXWA
3UMvzqt8v8ik0VOMk+bhrgGvxbLt7H0E9Z/SiYqdV/4OKR6uQWnnaYnpA8/AdDb1+M3kVvX3w1L9
ZSvg6S/oZk1wgf6E5kOSAMtXDSXndZJNL2Qngj0Y81myYs2yCWb7m4WltvMkCLv084kReYd125ln
9kiPfUt3XOE+ftWbgk54wRb46ULoEG/pyUJDv9xFfnFntngALGiSUtUQqTTApkMgwEomTgT8t97s
VTY3ogjQAS98LJlwKHQFZbFRBw+69awv1tYGIhmPr6qFJfI9WSl+atmitp7f4FiJ8Tq0A2+4V82x
gjiRLXxmQnedABP+01J4NgYkhnw5SkJRTkve1o6WgGgZZYau9s8eLDAiQd7oA5QWEs5qnhrzoewN
PXFlYtSKDfWuqGu07LBt8KfsNf2MYZGcpePKlv7eYpJtoYw6Rn3f+CRzb5ZkH7swgdG1+On65gzd
gWju/bFjoUuEOLB8earEJam6bWc3uD7Xvak8p0MFHtlNdWjgHRY3N10cpPIklrx0PrZGTfRnjvB1
JwWKQuILX/Z6pYVeUALjdNC8m8tdOHbnv+/yoRB4k1N0O0dGEVYQRKgpSZzxiPq0dj4hDNH3Eqoz
kO+41KIy2Fwgd6qSpfuHzrVqfEOE9tKyx5c3Ux4A03Wzq56i2LazdFzV5beS3csdL0DCzzGlqwDs
A3wR2ZOKUuztuodDJVcrc4QnvDM/ZjcJHBeazEoc/XOO6NM+v76ctrNTjMDjbs0wdWG4mBSttlGg
h0K1oI55xqfhPQGyjgzBJKCPFBDfTocYlxrX98bw/YPqBQllE/C09gL9De2ui/AoJqfTOWGNwGPY
EPUGrjrRQZCHt0X/Abt3/rQK1cUBedvxyq5A8tFpjdR8KwnwNQjl+xtV9lZi1z620f42ec6AMJv9
bwzCg8HDFbj0r6VqXDIZIzXBCytsHeCDafS7C4MkTyoMVzVT9JncEYSMsmoWFB5BKqv50wMCQfZF
527oVtc75IYi+SEF959lr4gpQzdPCdCTOm0MJ2lElZsZnCBaE8Ar13lTUgTPu6bkn6D/Jtl+9kQo
dpQH6fc/LvP9mE1/m4tLrwszw3rPo2Mh1sm/9B2n1osYv/dAe/bEkTWTeIMf3Wb5UuA+N0dzW7i+
YctpnVFYFePfhG2hnDdi3fBxS4vaBpTHUiqWgIZL82qp862XRNLWK9B8X1qHeyVjyK/Je8hywqus
0r4ynyoewpvABvhEQtTiAVu4w03kaX9IJxdd5KRFOr952YVqiq7zKlCsoya7GZ4Csa2DfZ+qiIIR
OsbiUvbsFpQapE6APYgyG0TVWVIM9LlzsSgV9R74KiVzz34uSBikI+IPmZ23dS1gUYc6X5/AHQZk
XH+o0CoiNVMV3Z7NCyDbVvhKnlKog8HcXh8OrXLtYXxPq9HPMNZ1EgOQV3n7WoYvumlESGH/RDSC
syGI6kM1MXlSWN8EvH7dfb0hubqZ8KuBnm5/BxGJh+vD9SPfukUnDAlJKW/T8Z+nE5Tr9J5oc4tx
Ok8FobWUMEd+yLV2OfJbfDGsfTNtWlAtAHinN4Lii0JBqL6aormbTy51oF6Gs4vljpNymzZjdK8r
AkCXJhJSTwe2q0n6CPBWD8k6JsFylKyRnoiJ9IBigZGLGgHvqBGHLX4Vupla17YsInSo5Yrv9S/3
IMBS7XfMG9Ivts5S9ckmGqm0yfNGHSKLr/pc5oCAI8nxL9TCC+Cx6jr3mCg7BVqB3C0vijVJkm+9
BOrRuHbIJBGzhoQG2gGkXI0hxooRFYrxtkjASuVplZDmS+r3hwZqfapX+QSUdtCnA7v3FjFJyf9/
Pb7iOqq0bW+AhsK4zZn915S1o4V0kTVNv2cHvCBiF9oOMbSHradfCo74mFQM5LFQj30R+i+uqL8m
xlS77giRFJ2Db11AVUEqv8c7W6AemWvf/ka52SfS7YziPu9hVUdLL1KCYpaDvN1u22aPPdgyh5h5
YIR2KNitCFCpLa+pEEMLFat7EDMXu0Q/juADhmIZP50J2YHAua4eh/xErkqtnAvNAYr2rA7zjl+5
kaFs91hRpflw+X1o6X06Orxw2obtFOBg/LVFnroUlrqwO2n6D2KULVQ7r0GU5vCnnBfN9gY/EJiq
c4CqJG7i1Bmf1SoJTvbzcGLjepvSI7+Ox7U/0W2Me6wGbK6NRpB701BP9K1+I3g8+A04MAhKAI7w
1szu8s41iEySRQeQHGwHsYP/MtbMjVigRyIMpJVVGuuvQf/+ZsR4rn187PgtnrCxLV/IJxXp2Bfo
8/SQZtC2zZtJjz5DT7t6LyF9f83bb6kMWobsOo7WEEE1BuFnCZh4YazcjC3PnTIKEYR75qydOu+1
C3SiyJyZc4sUbVbrKpyIuQzMAAD+/tpzbOdknGRrGkSKx9T6dAIu+2khoGdZeSTkSRx0TkH+L6pD
2iVLCJv5kOcyf05ccHc+iymhrfr8kZQfnBE+KD3Im9+STBKmax1TxXItH5b9RaAq5mjNnVAh4Qa2
59WQkXZ7WEJAqcHjiRvWdgJf83OJ3fxgXuSlmJRTneK1XBzVVuiF8E2TY0Wm5W+AwvbOsiREBWMT
2Rssi7fUVg5qdPCaG8hVWgSO/JgV154KqVeTHXlXLhP9MYcT7fSWZDxu1DjxWigvQryYhdWLdwuK
S05d0DDunXvi837/6H0yJ9LaCbZseydcb8uBWOLt4OzV5YubV6uHI9wikSRO79OzZcwyoy9ckBJ0
RJ26re1b7h7Cv+hlrU9V69RJ5+H1iLhJcIJULCPwtpXU2xjpx+GD3X1arZ9dypvAsqJ+edDN7k1j
Of42c8Jv3L0xaid7iuUFp6b9KcEZwlzeEjL7ZrnZWJzQlMM03YJGZHIrNFXWroLpIH7mSZdWGris
FEG54oc4y+FgVwnrEKNUPqcYFvvEE8OB1isnrVCgjCpcfgcudMVSATwbeU6IOCIZO1UvWQP8ybD0
iQoeE3u1DMjltyU9WXDJVrLFCE/XfSstEyY3nOuuSu3q5n+NuaqQq4zXfDDvOARAxnPouHLG/lLw
7t+U+hlCS0oTRo1kRIEBIDDhP9iVCqablsmYfH6NQqX6WQtG/ZVKbqkANjwKewimBUX3+A22qKIc
CykRlnJLv5ZZvP9fxjM/Ek+EI/dkXeNTHfMWjGoi8Cc7r+OQilxJYR60jiBPsuXTIiGVd9/N6ihe
w2cHVQCRAOi86qK40baYegxF5TXnBeFnrWbMauXMIMDzKrIZDV12SIkL7Sgf0yjzu9e7oQ7xCek5
Zf6JoLvZ3YsYBI9fph0I6jde2HkViJ6M6dQpADnPL1xIxdgkmFjsmP5oU0fWyNNBEuCnOgbqJE9t
IslDP3YY+2lOd+jI4a7Cg9YyG/YeGrAmyrVBEigZKS2X2bPyXy+CZiMbOa1Qu69+s3RGPaHOn6zG
fZKYgEfn0U4GTlreFcyy4WHGxkd5KT3c8c9QRuNLqxBw9LGPqEB2eg1IV4xl89ok46OJfO9rxYKC
HQkwblqgWeJ25OOgNi3ou6N5Ru9nmjssJ+707L5M1vRh06kuA72ZyF74auSwKoTVWZeln+TgRa9q
1vDznuhnv/jRfby7d9urPSQHpWHn/YXOQjuYO1MwfrBxAlmyPYV8LyEa1j0Ea/TJva82N6ZZkmtd
9GvvsNKL/u1KCNVoQqpspP19uhLrlSKVcJ+xk3fygnGauKlRUjuE/o0cmUZDCycMFT9UfRvHQCtJ
hmeAKXq125M7LfpcdBQeS5wEUSwUTXjywstYD8Gxk5fcM6LkG5oGArlnFVnu9l41GMYyeWFYc+Zb
GANQyfDtNsiv0pNBqQ9tA/SE+faedlUuIXFWUhUra4l3+Lz1KufxCD0bKOWaZ5hhoxQhnlAm9p9p
Ft/tKBsGS4tY+aG184xI3L3AZzFl0DX7RDpmCciUs9XJjWIl7ffkLiwLbKZehInBZmJGw4ulXIDs
LNUUT0A6c7gavNv74XJghQFCZ2VjeFTkl8AZaJFrh+WWNy2+V0jtN9h/sBB99wGtWJlS7EzlZQRB
IN5tPl/PmWrwPgxnL5A9nF5NZ/M+Ij81L+bueNkeleqP7wfCh3j0+PFJWIA+AULtV11R35unE4Ru
fn1917KyDBdIAzPBGOHjfcm9200BF8noQqhtiS5kZ2Dcp6/xfOfF4nZy69dbzAw4JS9FtHkhAH5R
8KjcvJl/moPIrf3QYuMH2GYBb3sKqkuEuVjzt8qufN8DqIiVJhVWQoVIIyuKJMSnVXKDSehDE+t5
ZuKaTsEB6rdB3vgI1PykDLO0K3WI1siUI1lrNqx9WXrW6+aUTv3Fj4D1B14F8oJb2g4c1W/Hr77R
lz95wfd6ybSqDJN03sFLfrVE4Lq2LzXcxB7BH1TLfCg8AnBxqxZLONKxmH3jzhWvVMn1yTStbI3/
Erj2sfSUPc7wpeWCWL98O8IWSIqfmqHhEjAQoMjr2R0ARK/GZzMFb5LI3PV7CAK8R5NNMMcyj3sb
oFFjA81atgm8Wv7A8rqZUPKC1efItv/1Zfcys+r3vTwFTwE7Fu8h8Le0WHOk7lvAx1Ea8SOLm0yO
dgRiDojLOpGm+JIlwB19EVFsVXazW3nqJ5paGVjTqSe3VR3+T4Orvs6vjta7xLgQk5ST81BIrRGk
k0x707tDNiEC43J7AhPKI9VXvAlwM64jKw+YyaAw77/bgti1bmuGmorHhCimU4n46u7uCFP6239g
L+JGmLvAzVeecuPPgWWOnOFnKMkMh2Jn5FIigpZux+PpPKqsYc+IrGOpQJ+Ny53H+u+EE3KYdLqe
g22Q6fsWy8o/bPeW8RzhZb/JpAKRNO2uta7JggDCCMl4e91TrxEURd5TyMsz6l3p++lFT8g6i5+U
4WEUjT1xGKql6liBnJQ0OGNy/RhGymWN2s49Ovbq0G2vk5Fknc5vYoSs2ArjST0vVDde3F0CXb6R
66E5DKSVf6cgx5z5juq7teMqSNdyd39qp2pMGR8BZMiTG0f8mOD3AdSjVz1r+5xZ7Wogr72/uz0v
cCKE1q3QVXrrc9nZw15W5hf4zMNnnXZVgLxRsfpRCeCPX5F9e1qYy5lFnSN3H9a0mRYTFC/ySXt1
07uwQ3qGh1/695QSVRZ2nSu18E7+9lDUrsQyyIbjaQiSV8f0wxqyTwogCvyY5l1/SCjwoMTr1EQY
yYYJ3zXhiX8WmB08xNq8GpKnWAUETEzsOr+gC4CLm7KjYGQg7/TAPFQxVr9xNCeSMyWRVR5F0sk2
X+Y9k+4MRBkNUKBw9BeIOljgbBC6J/FXSz3Ps9rZYeOD0zX2ByoHPLn0h3g8UV1Y4Kl33/wKowu3
aoG8prjKUVb2IDP1MXFknj3v4fzGGvC9TKaB1wl90De5v9ltHRgmdswI7TbSL4e+PGPHUgM1pA6n
9BjbE1xtR2TzwDerAIrk1Jj2jIzU6XSLqyNf+BYjK5vzAqsh2pWDBfI7+4bO1VdJZtd7GLGaVpLl
Z49fds4x89KShKLcI1YJJkbCETjDU4fc6oIhXIBI54gRzE8GPbOQwziDtuvzOk8C1K9clfyAYsy1
aElGLsNdiodOrE+dmWXHQe8EsfxpZaEjEW/reTDae/rOFnkpxgbLNpWeN2lIE9LHwq+mP8HzIRN7
OuBxkc+tUYyhwOTMNLEjDpJuoTtxRQKGvFbyhpBzTU9wJWzK9JWKxXd3Xj3gQCsNJ74lxOVKLraj
7lKPjGkJ62/+1tBAwXk4QTzcImNcsEw2qt9hK3hZ8pewOefp2E64CuNMEcfoxbqusl2/TpLZhlR+
+SOf2o6wnnQ+MXpq8qkncWHsKGIcFc53aiN0b/yzNbnfH15bGDIEV2wnEq7li6T8s29sPR48uYj4
V3RkDaE1GFRnAjN6ScRla2UvYahUp9+fCRlv3Dw+olSSWZhlmagMe4HeCbEaS9ww2+2JKNqJkTa7
82cVRigDGNJDw0TuTlTKD5/ye7/QARSmj7vY9SXBHqAGKKkiWjpVoqtOXM64oNZ+4WV/hNKUo4aK
6bp8GISSMtHPlCNvnO78EQb65oshqbeKGDpNGZlphycEJzjCRMnDbzdUJZex5QrZI7zemRpqj9IE
KiR7Cs9P7fP1a9oIzA5oMaRfTs7u81gT0kXVc3LlqCULvRUTsq05EcIlt3LeWrpQKMq8w1w4p4Sx
+wGp48OmYstAPyxlRCcd7OJ9H5P4sJeAw0ApATCINy4RlbBhP8xcN1CMBUw8ZoJ2VPWQCzmOk/hW
GMwkx+Bvnon2+heTB5XnU02Lpw/tIqvvplAz0YcAgXdHO0ydVdGWjuHC+5utWpUv9bEKbIatgrDy
bW6wfRiAruDbPA9PP7lKgVP/y51uH+WJShSFa1gT+rYWaKCvrSxCOkg1SfC3SRABfr3Ivlgr9HwO
H6IGiHA+T2o9apXwPdI+pvPj2BcywaQ/cdWdIvI8X5U7NJ1lQFzRTJir+lczk4FWnlmOB3SnspWy
BqLDy53Iu8IvFtYFypbDjlX30rh7eMmIVilzBdRjmD84hFPtqA/UR4TrzhGWM1moZa8kEpjmeWL/
tNAcqMYO4cmyh+STrLFdA8dE496ybiY0QK4PUGWf+ZDBop3PDM/FoM9DQKuZSypxRKizoHyOS7gX
7RngKkYkFHwHvyrNwkRXiUN+Qbv8/TmcdQ4v1VvHaGet+IMO/pXq8SWFuxtyWQ/qjyLbIjheZjJJ
qHsjKOh/y3P83nI7tALREYHlBWT0CVJ7PXhDNfuj6HyBHqZysBtjDAw6dIUPcpoA4QJd9pzvvX5U
PksOPKUuOnS/SLiocG7EoazGjkixTwYi5VewrtL+2H16cVSETLNtxeusaWpZl9elxybCmkyQfq95
lM8eAStRvx+clgA+mYVJumPR6gOXghHOo0iiHjEdrCC2ZfAcrsLzPdDkESjYSA7fWK4oJZvWJ7Ks
d5CTUnOOYLQtX1608VInbj3MFoa1UUW9Wui6jznptX0bz98G2/6Cxu2xADDg0GmEJIRVKOmGCUmm
3FOHBqc/cszN3q5ZN5jJjTUo/31+rfTgYDluC2fzF0dfU5VTalf8gv8hcNwSILu6c5xTYkOJ5xWd
RtJCGQtYKLZ/SKA/VQHKCJQCOHiLov4VM0DMKqmTC8A81XOF7h1aEeAuWpdEOrKaa5XXv4/sBvRd
T0DWNo5/KxVGdMUa7orba/QpV2Vk9l/riYX/RTHMutVOnkpGbx951kvdSnIYKaz4nBvke0gFafSW
Q4AzpSPMnibn5CashhMnAaRrtWkfrhxCsSMp5eFagzbwMY7q6g7VKqTAZIRSgwBOLGNF0dvaN+5G
V7klLRFeH4sq2l6TRZ5EtPcrvE9JaDJJcbPWWpWvu9jUVyFs1avHCUTFfZGo7yT6EVcq4Rg4HS+Z
tOkUW/oVk1h7RRs6WQiJvXHSB8zPiwIfRAsquOtAIKNbFoPUWa9+biazoi63xdBlr5TkZuY2cJy7
01ZcTTHaRRGArUp0jSCR8WEexs4tRKf2e0X6XOS0W44vgPhDdvQkXMtta+FrZTnhrBcPHMvVc6do
HbqmffB+T1RtPmVc3ozBBLzPJYlBZ4GgCdB0nsVPCDx5i9HWgNO7NaV5ZM2w6QLyT9mtwMuJeJvx
8ghjYIwsnWsjMtKz/8tMnVaAmCfBqLubGyEqfOQrvUKQ9RlBBs2rXJlf+CZDdynkSpAJkvCGvZUI
Svix5AILy7u+IAK6337YHy3wzpYFCExWXe2+YGJ6p8WEIaiIXCpOC86AgCzPz2LQAZ41OojqIC1q
TvB+AQaUAaPmV+nV9qL8CMKo93nhBKZPs0WAeJG9urH6htMT6n/D7aZuBqm7lTp3YHHGzlY0tLMV
k1RiVn3dJHIAWpo0cwxbJqE93TJwuqRjewm6BQad1Pw7nJ0P3DsfvtnBKPkzbHt34yyCskRxo2vO
UHy+KLIS3dSZT7g3KwJ+G0wbItJqTeFCMm+U2UGjgSBaiWkYLmjdofcFrDJe+k3hXWXX8BfCR3QQ
DFBh58sqz09lgRyArudyI7ZYhbZ2jaustmb1k29tPx74J7v5dic7JgIuQkVNfKdm+Z6V8oF0miXe
4v5z73uUa4vuRSNNi+32eRKmYiuMzl8SsRs1R9ZyVS3aHETSdN26+fXQAyWO6nlE8uBhCFlFaBu9
BY4oFIyUJzuTBjAgiiOsMjXbkrJwgC93JVBJryqMpug55YMsNn/pUf/rycZFWfIPxbTWgOft0W7h
a+XuvbryQLThhuyUpDiObfWtJVWDG2OReb30dKzwiVNM+tdXriEhflcyPKtq7kfGNKnnucm9h1gh
sTeZW0ar/T+9lILx/t/HO0M+dvOhaQCOklwdm9Z6yGfITWvPx4BVtIDO5+SzAJeZPTHLC0Cu5Vav
3zj1tFUFLmbstQ9gHlddw7JMoDbgY2cKocBDTBY1R30FdALENEGQ1H7QIsbdTpVmYNTpHZAQvYzJ
ynMvBDPQPjsxM4fP8uok7vSWZkf23DthXpXHLpZbM7oMms3sLLODinxwtwp1jcu+fqzsNQqTOU+G
1kAXYY7+S6GYq6eSwa9XWmC58ZhMwpr/1uyCucI1e8yGJ72cCryKDYZbu+vMUYViukqk07oafUt6
AB3ZYs1UEYJTxiRK8DytQ9E1YFGvQGZWDrIVMhP71LJIdOoU5WoGT1fmUHn8DKfSOqwnFnrX0aD2
PerHxiGVduKgVGySrj8fVs4dxUheAt6TwHqx67tY6D2J35mInAI7ntH0quetXXQ9AVeqQdL68euM
xzo0e28Fi7SpgTozF8OlF69sVLSYFj7gUKJqPjZ/mgPFQxseNWKnttF6fHp5M0FT4d5e32tja+e1
LmQPML1Mye9G5G9Qq8/IYEYR90cG2MEM8Qhg69OTnZpFTMQK6vv7euQjZct++ptp8E/PrV2ApY5Z
cLHJgi+FpwQVOdzuhzRGsJvKImkpyfIN5toYbMUiKxHhrlEvt8dshRD+vrXaQ0VDpMxpJRnEcI6F
dzr5t+SfsSoxpu5ssspyQc2qTc8+qPNhq9ZQEuyJUDgiDYKEIf9fGksEkCpfh7fl9afoTg5ujQyu
5LKzyFH39rALzVdno0fos37AN42gIGR1c0QKXpt66vhjDYN94rXEbtCR937E3BAwrlb6EypJPaTu
f6JpoRSMy9HrseZW2Wzr4QF6IRen6JfOYcGbuVa/sj+AHJsUn4RcbciVruywkSkFnnsAV7ZZ4N7J
+fi52gKwflIKK0AP7RVhvV/ucn6MelrKO//myo+B5dJeM/2ccjWGQG8F2Yqgd5jN/QgLH5eU87+3
OBe39hAqgiKzw50c/Xh+2Tgc5+6K9SR+2iIVB7zEIip2swBOV/zscLzodjBjb/YY4HU4YKtARNch
DGYcEdQtUVsJmpcHxg56OZbqM32K+Akpe4wQRd+N9DuLn1e9GzdtVIPfgdwCpYIG6pq7dot21ZWw
hiCbX2Fmu0tjXHLZ7Et7xuTk12hMdSbWp5fWNG+wA9GVq2RB30RNyiZJW/0mNatxgqTOFPV1lg+l
aWi6NBmF/fOB6my92PUhiQgdMxzuzlquzmlwJFFBFoCZ6mnOy+qZ/uklBWsxyv88517EblomMkya
5dzrSfHt1G8gpFApMuHJNIZLeGkl5x7C8U/VSz7gimVqbbX9fQZXlyLf9FwnGxWG5VZEJFAXzEUz
fZAexqVh9/sPZwfFCMjAhf+rHpbrdSPpAZSSBwj4LSFyXtXM+hrETaRuY/r4ZahkJjNWCX7xgGj4
lUgOQgTtCH62a0Yq2/+KWhy2AFOI8LClEQX/XQPJAx4N/hTSSpuDgUNg7A3Tpcz3NA1sWrQBN/Rr
3FCL013Db21L3OQooBnH1nCg4U/0b5GvGsT7q0gOX5BWw8gTbGV0R6LaY7J+IRQ2GIgxq7QXAu+a
it38Q/oGWF8IHXVbeM4FGH2O7Tna4TsnzLgsRMN2NMdzexEotEoit/LIb6Q81GqMAzD0zLwd0lKE
DQ3XqKF7VaPUqx+eLq0Mg2DwLxJflvs8l7JtkegMsN609LVwUR69CAEew/eyC0OFb1JmexoynDu2
ZWtIdSSOPug33h1hpkP6frQHkbf8aB/BMBK/FTrqwSuDKXYScOzp0NsCf1iCYTTcvxCaZ4BbNpDh
gn47WBafzPtDnmE8xxGATTGhlE5SWuzp3EIR89L15YYxOBirP40uenXJ+++Chhp/zgtdk7SAbcu+
lNGIqr3s3pNhTJAZ0MqMwZ9uyYSZ3AlbfEXfC4f88QCSJvOv0h/r1wZxLW9HOmSWSg5u+aKcqXo1
JOldZxfM5gqMqzVHp0hyrj92CW9FfzdgU6XTXhDqut1xyIFe4jhGDWf/puypvELDB/NDzVZWhoH4
wETz5ACugsDVr45fXcqMDExNRrOgkNilGNjHqRj8BmcABsfm1plfjJ1n7r5f5MCRDwjZ/5UuoW9N
C3lv3926ZeeieQ2SX6+Kafsc1SPOLlzCn7CPRPMD9l3GQHtPn0vSwvnXBhJqggv6K3hMlczwXBdI
i2vcCtcoVUqknXvysQs7jOPlnLHDGORl+0rUygc9a/lLt/z88oPZE8pwdic5HerbrFgbL0Urhk97
UQoeh6NVQKg9TN8uNF6h+FS6Bjq/o1soFeXwrs+08de4JDp3RVwWyzc6qqDThMTkrEPk8WkVpO90
SgQYEvqqoqiD3tJeOsf1UUhFDXz9UakrqoGmylPWi7TbdSGaxTqSkpaTe+JE50Kb5n8b/zqBzOpm
emu4etSUQMT2MbAH2ATN2uOqLOCUs78G+YAPmtjtDOeHJ+8yzO3eKSdgxs1lub+WoUCWks6S9L3n
0JUs1ELFtWOeePg0aD2oOKZ70bgf71eSpFAgW3ksVARv5pr/mW1tgMjZIsrLilqsK+XjemYgLfbg
fZ8HHQMDx5q/YrAXYiEXrwo3wK4ZGlAM96CRaEiFexGzdA6Lkwq2QeCq2KjK4c2HqTPEIkR4mDVJ
hh++OiCJmA5jgBUbasphZafkoPMDiSFxlA3zHA2rpm3hJT7dCSZzh27oDALNN2xji5QpCei103va
UsErH8wtXZH8EDDkK7zuZAuXO1ReE6ZtLbyYcZVI6gMmLbUgFkRJ4jTGUNdiA5X6942tQFqOwupH
u8dQLAMROIgA/LSrn+bjkQcaLDo7Lu4ZoiGSxWZq9hJpFkS4rX5vv0exS247cQxdoh+gx+Pqaxvd
+vC+o9R3xGEr0vTTvcYWfFW6+3J6/MAMa1/PizXwpViWsoJtpOU/x19cCWiAnSFY4L70gVuqZ9aO
yW3Q6gFP4yq8QCo5KbQ/UlEHA1J1NAuvm5zn0iNULU8V9byFU2iaZnG/tRK9EiwDoNtaZIgz468j
bcccJfySxkqDGYUcdX1Smfn0U1goq98aONRSk7D5JPThUCOGxJ7YxPcxDbaQaQU0cOny6SFaU8KI
9dldmEB7R5+MghlRpz+O1nGNtC/3gg7SgJJrHRKw0xHdmIoL9mHylTyoyzh8b1pTPfzCUgjEExn7
LWxOjNYAoCIeu11k/FJPkwg2YZ6s/A0kEaLqaUvkSv4mCzKzxoFkNYeq4XpPvnMtgCcjPnMQQ1n8
62dQ9F1OwzNL0GhiE9gRGTNGkCIlvMzsZbYBmVjERd4ZebJYlGUR7ADI57CM7QAgpdZDN3M5aghr
vs4D4+NQ4mi/SrvvftBZGqf6+jC1iFFHuCU/61d735BvLc+XJ7iyzxqZc9lPsG7pt3DJGGJJ7PJ8
mL8xx/Fy1dmOunhnczHtGEF2C5DD5QgfFPODZyv/qSoG1QxRHhJRP0ZXkDw7bzaKor131v96dNTB
07j+ee0Q5YCMAkSpp0RaDdF4gYdk7uAAv1GSrVf9pWX0oKD2Tn3GEMfsVCYrXQez7eEKOlEnTAmG
DXfVAMV0sQ1Go/DpuyXDpLUxOtM+WEnYsLhc2F2Nk0oNpuMAIbMpmDN4p8ACwE9JyrNp/MoLXOE1
bvUkYC3HRkEK/7uAZf995ckYGuy2vrt3OPPjvMN9NEPnmvI03I7ZrqLsuEcWry3ebJ+wsDiSqxlC
PLT7Kv7vOS2r92hlx0Ss8Sl/1elHL03Sc2YwyZpBHZUZ/w96KGxuz/f4jMrpkJTN4fIeKs8PS2qN
zoGmTvRF/S+PeIQCul/aXQjlrOW1u+Xd7YwWZS7nR5Pyej0V3JkWUeKpgivYx9TPW9ltR0awK7iB
95X+Io1xsykn+2e+AKU5ZxfnRABwkHuwKU+01/mQTXRZNr9QP4m6Z2JvqaYIS4Aw5exkoYxW1ae5
LXPjH3B9BjIo8Go22Ssyi9fOvIfClszmRizw2Vc+KWISc0QrMOXYKScHsm/jU7NGlCPLrWs3VhnF
bhE9i/nh93ZL+3q2RKZayVC15pDwaYU8+S7U3JXboiNZPRPmcKDpwDAJFNzzhw4E7YzxyivjfXVS
Le7JoarnuoHWVMwfj4nSQvW2fGi+kP1awyz109UFSlmpdpQlBaIQVofKvWA80iTMa5j1pLubW2CD
rEQrQSx1E8pPAj/DZcfAk8Rn2KREYl3YPrPnbgBRnm4MUMSwbOe2GwBiX8z2TS51jB86X7rZjU5t
jHm04+SkOPwjYcsn8On+NgpIwr4uoOv9EK584Jx2XL0qVYt27SiTPzr0fxF22X19mKkfrl4ih3dD
6j1CJy+NYdT6GbXbaMae5HphzwSoexeBXNKCtJb7BmyF4u0dkUKwedNlrAJzsBXJ9R21pKNBFJZT
ljxRejrlSXVm8wHO3mEK95YPUL4iYBIF/g3GR48lWOD6E7yo3SkY04iH4bOZ+plrzpXZXUyJC9Bl
GIfGezzz7HqpaU7/Bt0xTA3CKvagyZwPfJ4q1BM3yOCpsUTGlx5IBZtDNJyAHv0JGjpb7w8Tyn/B
wGE1gItajVGBAkD6Atnmu+dVuYiiB4C3VJw3m1w0/BWizdPkeHExnwChsYsYNcKMTC4A2Wudyd6a
cbQzfHLrwbDr/iJTUAbubzlCpvM9M44e67b2wkwvdUwLfsxnkJAaVPAompyAnHbiJp1qPaH7ZXam
yL+J7BB7/oDpWGonFea1GhhiCLa/Kvd/GCnguM82sLSI1QfqT713gQ5x+J2W/JEbjC4m2xzaXTZz
mYCVeHASwyIYQyK6sS2jBrNcUMlqc7G5GnlmnJrXF3Pbdc0ucdLnwOckcxmatZzbsMBfgn0DAdJk
SzFRSqBjp+muhHVvjRRvsDmV8x0V+XhchOqFeNBu1Jtp/N22Vq7vkbQr1VMZlpH4h1TZahhhDZgp
Ch4vFrCTx/LD43+a3Kzr9+Fo3Jh7MNOIFAuo9/9XiUsG1eNZ1i+1ptLS6LI4Ju75l8tmiL33qNS5
OLUD7RbGfYY9GlWTzc8b+5YDPede+FIrIiNLzn0KXfHDYYlZ0peJmo5mv5oRP1CMrMHmpV6mAKKp
wfc0XEA11algStfGf9pgtlSe85tEGscpc+JjM5RaFKZOOfVjjy6sJYSDa6WZ/4jQqCeBEu8jSpn4
bFUiroyIcbhmzPQ5CE8Lp7nSHYxBE4S605zjQXvDg40qoZPlxLn4CRqFt2zrscdIUqARmub/2BLJ
r84IZLf1FpssLLzh0CihE/ous1HC2wpXtcN4rjYk+noUms2ntNR/u69b4KNgepageF6KMwKL1XxL
9XVcza4mPUSky3yx6Shr/vcDca3OcsFZZDX1UFBYww0fJ2IUDSgT06Tx6zRA8N4AvPEQMjN6LX/E
0MaOueXS6aQguYkjVDAPkpEWT6sSxuer3TZU+zpRHObitrwzc6ABYyfVmKxcqtqMmkynhIkj8qN9
7SsJ3oOzgyV0vzJTZfhYGcpdTVK+X8nqRtoNQDAp/xYct/f+xbXGzrIcSmXwRNPSrP2uENLmmabr
wlZP4VRdSuHN7ByRD47NGz8glBQt25XXCXjZD915PTNIaC0h9zmM742L1GSg7DYSBhMbB0qWWNYg
D2nJ2BCMdexbRkiegtjy9Ei6qi0NmYFbH7OWQ9IdlMbTdsVvMbVIgbB0mEgflOh98HJ5aIZSiLYW
HW2f8fJYKdTNzro6Bm147bOmAXmtHDKitdwyBWvTTIqC7Htv8uDgWLrP853yC+Sftov/3EB+XDJt
nfV0hjRx6Jrxb9PHbKfSSWwwb9xTcaKq+lUHLLcZjEa5YgAn+0MxS7s+8jYN+s89RpflaLJGZ8wv
xJIpqCkLf1PY+VsISVUuRrxHUTFWH8Nefg9Fg5cL+h/wJJB5bCPR2QMQxN+M1zkZfuYKypmBtqKu
DQ2QX1CHEsnchz44i+nKjeHbsw4YaYMSuUb32v32yshlZ74tcksy7lCKefRw+3Yl6cIcUsQjkPhJ
ulvDlgMrn08gTpaqq1/wB7w3pjwUGWiIToUC0dekcK9xxiPpaoCz1b6vTyZehReqb05lq/XeOlJR
faRqC0BNBf7ReVT9qtpibhZO1XBt/vag9t9lNSK7n+h/7ux6bNgsaqn6s70BpCrd3bSIN1T9C6kp
RFaixDCtqQhfoHtIBcUlFio1CQr5XAHaLZNXl4GE4mGkGJOGVQLAxEBH3YBt3kNgFfMJ87ucJevb
kl7lvnWDXDrx+QSQabawfbAe0M1Dy5HrXeY/Tg7ZveeQnqRtSiv7ux84lgw7TkD2JhxIVHjuBM3e
eVABJmOCMpJIBBUYvhlMtY+6kn3YTrRSi80HMn3Vyh/QEewDWu22cTV3FkZdEfYbYQAjthvBTBBn
s69LhPOhj3qJb2jIJ9ntpLEep1Y9vGBGaxh6reBLqLEdlMXzhuDK6SX8wYfnM7/OsseJ2Ah4APO6
K9lKX6HHmQ9jb0Lum+Pyw7csf7YfJkSG81a3f3ahwaxZutXiK8tgQRXKb00v4XeboSudZF/0uYX6
LpwypbD8cBcwKexlYcAr8fEDnOTArRR1pnNo5A+YR+iaIDJEHbyjiB8OPbeKimSdaoirqSdN79yr
O0iJmqPEaEqUSQoLWunhVlItig9YMoJkiiCsCJU3A8hCqh5yjxgnUBeGUSa2Z9lEAsYxWuTVsNJB
5ajxDIRXtquc62rdl4L/scI6EG/FvQzUuKwNNnei/zObEytyTaQoN9/FjWNAdSqy26s4VsYu0mLW
h/AWnXDLb1ayFKSwHlNbud+QrU/JLYTFtpS4oVqBF6sRZNrdGbPpv2qYTYw/TVZSRSbSYnkkOex7
XAFQT/6bcnvcoeG9GIPR6XHgAg/+V1M/j+iPDBODGI7hakfG28SAj9m9GCk6piKU3v+lYMHifwct
hNCxRjT4n6icKdpyeVxTz7eLMOitroGRzPgFtI71b08hJdWVnuEgurBSneldWxiRfQKAEDtdaJwK
Cj8iyJIjp8rGf9JdPY2kCkY6XkKkd2AyNfjHkE1nnAYhpHvo4KdDaxZlYipxmBV/wJcaA+ceWAyl
h6XcjqAuCb6BymJ9EFgTiJCSeOOu5gTAPxPV77tOaWQGYZhrSk8LrEKMaWJtALxTBU9sK6iCuIOj
S+StFyg8KBEstU/dUVDd/sDFUK785EvWPOmLK36cPUZF4aD4WwtFdan/ia4AP80jqEAGHjAYlg9l
Foh+yjk2naiidZyzz/O7380Mpip6pEgobOyJMr/omXXjop5qSe1uNiT0qE980uXhEu4Z91sK6PcT
FBGDSXcbTAgzLrRXe11M75QicChFfrgGLBZgrdZ3OD7oo6jPGFnQUnJaSzktoMxzE6hVZ2IzUQwU
O91u9b6qtn8KCQockKIleM3IHap3bE8JYtSeFdqFGhdoUN5lGh40h+RXOaL7zbStZqSi2l7u1mqO
FwIMOw5OYnqp+CiRFl/u0UnUXFR+FVXff/gN/Q1zpzUh8D7Zl1VLEcmXgwELIcH7lr0LoD58fWUT
aLv10ucwpwrSExumKjA3ogT4oZ1WnjIAxaZe/tYyHyIBgfPDF9YqmLsn6dMqPfNbuT/XPK8vXs5Z
8k76rdY+WKU050COeJVq7qhZ7XB5kEAdbzo/b9kNxPfnx3dAjrZeGlwCBULfOzx9QA8c+x2vmbyH
IXYs3RLxarCqfNOelbBmHM7zGcTaHJw2TUwRzmC4kh9CHU9PmrePzAWJWh73Rjj1/pfNtepWneNh
GXSSCXoh8H5lnQ5hK1+4Gjgu7he5U5arsrRFOthSKn+lNyN/eI2PxM5KeillTGcA5V5hJqtl6FpF
vYI+u+nwmHEcfl69Puqkw8ukKYXMq5wdHjqK+QYTCTb+41zFjDdGwwD7zkdD3wZ/pgvJHFld+S5g
tkvY7+9fa24bMTtF+G7mrqUdDK/9eeTGzlfvR8S03FZiXnlv+1a03le+nMqljlpYgVyLTDQMRszq
etV2NKEwQD0yBjZfjiWtjpBhyGUPGPCWj5UGQhSZBKJu+V/diiMRfLO7QJGn2Jkr1pFZW2KEi+Ps
KAdjE0HxhbXB1dDTdi0MQyoezzDoIfo69JG/Yg9GaBUzFK7nkO/yHB+XUzSFGI5MJzRAjnNkM/3n
/1yRilyi6UpGRP8r7Ali2lLa8u/jeKHjNi0LGALqBK+ML0hs0n1mP1rKmD2vPJeEemwZBmg2b5TG
miLQqvUtJJP/xdKNnMR/PXmHg53TQrgSakQKiAYx9AofdcTTr0mUp1RKYSBpKjWrPXh73ai61lI5
+VWF6l0C9mwEfHu2+yZZrShOGZqpHCtU6OgH7YNMi11eg4VT7YPGcku2ZiyH0oT5gQKRw6Iow0x3
Q1Ruv4JIKY1Nov03BtDRNvaWIGTVs0Lgqot89DCuGWgQwLZLWmXZcC5+7YOWfIdG5JqXAiteAu63
5gBWfs7OepN58ur23Is4+wfvPzcn684Kt7j9DIdEEFzOZWxOuuBqQko6TKFG1sawIj50G1RVe/pJ
H0qAItOxjkCuz2wzMyMVMneAygbNlWWkZSDuCJJhjPy52yt+klwa/rUA5Usylj2DufZZZ/S65WNo
nJ6damH5R03yBR7JPRwaLohSTlrJTZiKLAjsCEoM0hjIrK7VinykN6mtV7XWTlmdKWmxaN0MjYMA
sZK1PZKE0/pAsGGwMOycWljSLxksq8/7z9hOZmPpbVI+9VT3CNBibsluv2DhgqbyDcGYtu0B4zbX
bYVG+BohpadJmGEWTT6eXOlkR/y2LChgDXxH39jIfT+7rL2JYRfPVPYwf09OWflcN+8n327Ld/Pm
6R8+FsXrSPeP/G4L2oCZnaVzGQDxbIN7jrh71nRxavyQILtIdhqvcywYBi5EmV7uwpo1H9z9bER6
hwxGx+93Qm6SMhhRWJYcT4z3IeLzmGV+ozdy57TzdkrlxGubXcT2k0MjQHwpQtzBEsKzoTQK5o0D
/ipzDCs5jH0ehSwUafUpNwSxtzntyMjH7HiRKmsJf0hEVVd9jtC1hKOI1PsyId8jC/aWCWCiiccA
1KpBotQQ8ffHHb/IogxG2XY4M7z/hhKSqYJfruLERa4XByBL+EYLsmCxgeI8whHHXLp1S+S7GnIQ
XhKSobmNiLh299O/1E0l2KXDBUt11AsK2LvOo40AaomX60j51Tm8LHrOntEtBXM86c8aFhvlICMx
ja7sb4/bcZ7+Xq9Dd0OkV41zTothj5xWZJ6caOsikWh/BUM+NqmfXL9emDHVDjdfeZCEg/AhPvch
ljp0dr2vFpejZFOJdqpdRMnnll/D8MEycQN5y9jlb/hfFEQO4QGThb1udYtmheal2Qiz/MhQ1fO3
Twz0IYKOiVOQskpjX8Gn96GFqf6ZtvaEzl07IUfJUQja7a70nLNKHQOi2Hsw4ka0O0ZSUgit6lL6
xumxAOi2uQv0I7ah/Boc24hcV7BFRRuA9gMUkssEPwQUpMtwnwdTgVpwO6AgjkbhNQnmnw8RiqPi
TnqV7vUM1BPg0VCWSzSJf84Or5Ne8C9ZtQ4j5Zpx9+u/OLcntlbQDEwBfKvKi/W6LX6S1y1RQXL8
DWtySOyPU6RYDRm3vyAlgSWqQBc7znO06BL6wHgtpjMvoFYecUnC3wpG1KCFdaGpt6e6q4j/0ul9
0AIvK8rfTCyAT/+6qes6mo9wbCyVFfyGDWwbSvAB9G4t+DihUhazKvftxADatY7t0wfqIKz/qb1/
hIau8N2MPWVcmEUHgYbOc9f8ol8RTweQvQvswv22S3BfQABzKm3R+oUtkhu8B0q8p1UW9oMPE+w1
2nZUPizSihxaZV5FWCbfNCSpoUim+xNjy32lBPJigBBjnrozsgUM5BjpXmUKQ07lSr5NkKgDEzhQ
h+3NzoCV1oN7wZvWSf43rmF8749SRo+FJumhj8BKrn0GupVRxLfAgwFdVZFqJWDCB0g7MS1XL9Da
3ZZslkyPQeephS22+PRJMHB1u1PBrLz01iLzOgM80CiSMdLa1+vXEFn6WgkWgsyT2ukPqSfNtTHi
dyiZjhRu/VyIM8Lyed74SNS0/Yg3rWTpgffML9ii8OOhMhTTPlA/cVuJS6urLi9yRhkXLKiM5mwR
jhrO8CnCLnUNwPDqIZHz8qv+yBhQ/t4asMvORfrBms09RubnWcP98+RORlyabFCnE/c9guXZUHf6
zaCOi8RrWI6hD5rTM25c7OZr8/fbgxdh+PcOY8YRGOti2scohPdkr+hUvplG6BIvGi8aVQccqxAV
mPIWeuc33+llOX8nYLdWEg3DEh1TjiMWRfa7vhU0QJeh91taMTj/jCOxexs7+2I8w+dEq2XhLfKL
q11aS7lUj6SlGb0l+1UOpuXKPsbv4vCAI1QEENm2kFpeM9SGtJJXXUJqC64QYVtXKM/xkgxwDfFX
fXKJtlCozBUYEA4MAsLFFpZJYzPQSMQErj73CeeXVIi3ISPWfg/J1xex6Q6F2J2YD1G/PDki/zer
w4f7MyvFC9Ppk0X1OnPuS5plktaa3Cqi/tUk6gEjdM+2f63FhRHXVMR3Mj8pLFesczOgiljEP9HH
U5byOiRAM16WpCovUU4hRKLsO1F5qgsD9uQbd+dfX4Dr+j1vRW0/oQGusgeYByyRD7oY96kG9e3V
OiEOX/tuHtahE4mmQzuoF1EeAcZaU6CDgWzgzmn3/c69/q2VHMh8oCjU6JInSObr8tDeZ2UwS5AC
/9lPAbMI+EbJNPhDIvtKjf3mT8HR653U2hIyOFwKwDqcu/PTdkkUX7eOWaqFlMF24PadeHYUrdXZ
ajSiGDyz8BmvxzsiGcUXEG6CePBWS9giYR7nLWsMWHbOBjFGWCQM60kS1oxVgUlOt7A5ECt89DN8
1hw8jpFWBCPmmuEAzuwPldacoIGTHnhtc1I2aEGMOkUuTMBI0tbhybrPcqNPcoY60mnURtqBlwx9
ANjyYeGtoYBg554E1UWIr98RjVCoIXeq1qqD/Jylsd+YErznU1bkW6TP0n1TSTcNTjEMzinK5t0T
ZZVY2QLVhuZfcD7qSqbyh+c8VWIB90KiDHfwR9YnuTjekPtQMw55m5YefT+xLwAbu+Wr/Jb89vei
JzGB+2rcLZDPwshcc+O7aw7gDpvlbLg/Cq9QtcbSiNCiTb3ddEtc2P/QmTSQbHsz2V58ZLwKHzni
YMUaKwI63QVsS+95q8FXsvUabRn6htdJnynsCU/PRsDPs3pnQd27Y/OLNNjRDVy3xuQeOcm4owN4
pgkmA/YIwbEL/iJvoG1feud7MgQe+NcwzIOTUJADYB0ImDQAHPUpdIGKDPgmiAbF2JT/fMs/LPjE
eDRb3zyceQNa2BdVo6J568//4urm+nvBnErzrDMmVSLXT4IbYUl9nYC8TMF1OA4HC34ITyuJzlSo
q62x8ozz2WZNAVsbb6C12P6zEi21oGn9TkihcGHccVA9IZDK5yOGHpkat8w5+/WY8Pr+GSsJ+eTf
cmt9qAtM+IKblya3aYxt/bM+boVHJTMVaHAx+HzKu+uySUybzjgdn8kv43Zq1SD9q3XeGInboU0r
oSuXftdAyK/iDKITnEJkJKT5k7S/Zc8EvuRwXqQkahYMhY8b5wapzXoveUza2yU5v2IR7/iupOFy
+4PSk7hzQFQJKAAVeDsDM0oBFWJRh//TT6TO4geOiXcQ9XITmSBPYXUU4xeJuzWgDaA/0r5kQXld
+LMCpRO53Lmjd1giXNo+o9NnDnP1fU4yTLbnENIfDeIr1xUlZY4icoeOgdAHwl0JduFLH0leQjpz
eH8gBfQBFHUqXdjR6m0Z8u5s3gf/yDrn148fimnyZclPZEILh7EniSYb8zG6M2J6lwWIHddV5voC
HlgwZHxs+lBDIiuZxnzbfLgIiCoq5KuRQCeLqHkw2cF+FqSuoQ4ht3+Z6q1ORKV64JkMIA/3znkM
uqGUJbMCsDp+Fj+20RDU8sXpJ0M9KJKKgf3Ndy7HEYxiNcs3wfUOJ3wgIibDIpfuLxB4WWiJJkbP
6xc7oN6WInJ4bdUAa1ZF5MbbxWbcsBVToQWEX7U5+gDnyxB9LgWcGnOCM2NSy5tDMIHdcZzsUGW5
Q/PGcqTLSGWL1V/RzzGOicr+HJ90PpK/KEffPFKIPE2CzUk209vLtLumGdrN6XpNjzVoiRFVndwP
sSQppIV1RHooFtmBn/T3l0qUOxjzu2Kz+o5IGwTuKzaWSXuIJY/mf/Y/J95ZhYH2mTMTr24x2pxB
TDpQ4niEX0q3gfkqqHKvLrgsjp3yUZ+poD65pcNq9fTN37Mx0JqEIxvMaUs3qh9PWrV351DuSKa1
wcp3v9PAJeQT5rcTa/y5+bMP1tt6haCnvUesJ1huXRqTwYuanYjRu4Fja35/LNMJTCp0HHAIrYD7
cFmPqoL1evQq7SJkL2J8ftWSlV3gnsk84lJolxq8oFAXlQmhzmmEZKnCs+VT2IKkG087tw8apM7s
ksD72IuKJ3EjmCI80kAMUfH6BZ5FSwpyBc4JVc2kBc1h9XW2iIZbWO9mHLqCkJPbzUR/SRkOmEjE
kpnO6rPxfvpY0YWhUEJJUAkBrNWYqayMJdb8orbpb30vmfjgQgVfkCUoGraNd/MdJg/8HJMlAoF8
sMX8IQ6BZ72ZDidf9EL5E2Cw5sNUVRlUxL7PQts3monprjYVZhg7VV1TrBvi135UO2pq5Ssj6uvR
9L1MJEuO9tGwDuiqtn1PvyF9qw7F5+qU2yi11O4iHR3xl8Yeo1WMA0vNLgVLsxNsK8/aCAdsUzyj
x74OgSM5obKPnXxN6puPKb8/hdMrd649VklZwj2Ea8JIequ2H8rWHo6YtnecqDZA2tq22Ta97WLR
wAGnZz1NiPkZ47LrPTUA+uIyp7LSH6X+BO9m/JvWGChuhfRVNBZkAkkdSdnvgDm6E0w/MQ2PGMS+
8GnjGRwc1YjkTC46+RUp64kQNTOUxVkqXR7hyiw+wzsSpLDPF6RVtq12uht6IFw0SMLhSvUD052q
S8srFmKFDflS1Qdht4sjOgrR6XFYJDcpMlOVDxmvSqw5cMMpQqE4KQz5bkQT8O6O63aDmSyCnAe3
BFD+OkDuh6EDQx7GzhshXd6MIG917hkdf+lhjHFFe2uEWUIQ6CDfTFaHvbuwPB8my2l8F/z1r9kr
bvbFrJxlMUa8HGyAMG6PvYA76wN/c4waHNQkvZZadvDpkWyoQxkKFkTwOnHIpMf2ZqthOA7c143h
ko338MtCw6MMUK71xA51b4rnad3WXwepmSqSsejpdhxs741EW0BMsXKRa8hkTjuWwPU1HRxvGJJb
KTW+zBAHyM+ucaafZTVOEAR0/eSWoKiJd0E+OsXa4xraBl0sVRc77zpLuEiiPX+nAEqJCrZ4FV9O
Jaupb8vRxh36O3cdNwMxnvm+Lci5KJGLWsTIRfMFopdtcn4A9Tth0QE9pKOOT4lwv7chqiJo79Tb
3Nthmn53UQrfNpkDHpeVeGWyL3wLJPGGHg6HYrko90qlQUQe73e9g28pW+v9theKvv2crSagmYv5
p0zCSj+nkPtQTvRHfqueGxZfkwe3yJS81Am9FdcLcvbW9OEihmsSBOMxa0cWuuzROAamVEvcYNgQ
h2Ik7Ndp3s3BTXajRNqzay6DsnEsfdIQxpliS0zhmOauzZtbdMiJoE4/IYDoIT0icutGZznD+E20
BPdWkQSWfjrU+IRNles0VDqImqInsCFj3AeIVGEy+KTPMBbiKynwcb92pNACGZyZERR4GjuqLaWs
YXoAgDL9MYHrBuog9ANLWznqgp5Dh3mMGSWNmyOD33jyD0swOZLuP04N0my5I/VMPULlWBPGkNPB
Cp1Bf/Qjn91d9jUBZcWUki0a5yrVZXsYfc8m2wwbEtd+dsXkxtcRcLkObshHaDAOBHXK3xCE0ofJ
P9N2EzP/xgi4Px9eX+l+r2ZilsSpdHafmDuJSg3RhdxDT6i00MriCiycihiw16HJKQ0MUIjzI8RS
XPhdwrw7XIZMxX6J7CZCwozgg/so7jKZy/jKIuJBFScasKfsRO6cRx62uV6OULmQy3aRlil4eadg
MP1iKdb+hMMXSz9hQPuDBfBvlFFze792amNX0naijAKaN9cXlBpWgzOEGmTlY1mC2f/xImaJjp/d
NOWTjxJAgRG9c3FC0uIbuU8xvI4MXU04Ff0J1OWSM0Qv36Cz0c7LOER8SSyvOtjP0nMn1B3Q7F9/
1LXqT1DUWh/cziwey7GIilKMpJI5zwQv1JPDGrz6DUcvKQZfJzzkc9CfRltm+ryE2G9/tl4fhzzj
16B1WjMk2YSNA6/Rq1COPmHvqLnYvs4EmAKxI/hTrmroU8JIx+UXBnWpR3tOKCdXIbpqOz+VSAPr
Kmo/e8ThKY3lCPU/UAW8HhSBMY1m47GDPfw56RpV+YO2Aj7X1usG02ET+2mnh5VSJpqBCA/3NSdt
ofOqJH5zqlWbvPUFa+Z1V4yqfnXgM8Wj7VYtPN+x3pzt5zRiNvccKyjfZVd0xS6MqU4iTu7HKTvp
L83jBl54pz7KUsPUq26zOMmFTocnbCyu8hZUka3z9pxAd8UU+WToQx/p7fHDrA22vCCRY1nHLJxF
NXVZXlYxomWjfs9MtWFJ1ESCDubbubuvFeg+gBm+ksOvPyKfK3HcrLrVXNHdxNXLoriIjWCtVOVc
B1iUYS0Pm848CeEO5AkThkub4EVwZdbCsUJejwhtrg3TM7YNEWMPcbzw31INNphYSqb8GiNueoX3
Hxku5igMfaRjKk20e1gxl5xYv7RRdFqVigSoiZB3b8XwQqapdM8kQnYIqj1LIVs7So6yTI2YdEjp
iiZq5l8NsNvx9io6CcQFhM8HCRaa7zG9rRqYP+apZ93eVmv+uE4JsLLNAGl1DSih8c+PMmZMOvys
JIcbZf9byrRphhHVwpR2CFIP9EIk/APAAeluIsDK1FA4raUwmxwY9njnI0ME4o2RurFUNvN4LyFJ
d1MqbOGb1APEAriDxWsxtcBN9PrStvlRzjA+TpZ9UvbHz6Kj7eaS+GgJfYo0ixPR/YFldK/jJfL0
c9UeMEdSabWENtqThO3rsYhAjWQNzNwdh1hHDxtPsaB7lDRzXc15xeNH9DKRWEThW7KedAsP7xSL
kEVrjsGprjVZffvDRtGLrdeLZbULOBsLwS4LBmmIzCi8NLSbTzjDREMsqCJ7SB52Xhz80aaCEevj
gqp35O7wiuBflXaBfgcG+BFpuJGN8pTCZ+yPHtHlaut6XPIDvEyNIMUVa6LR880XaQW2BLj6vXSp
raYJEkpgaWP37svkyNcuU5XwOX3SzpX3i0slYewKrvlPTAEnQOBvfu5TKJRqmRL914PQyHd0rwD7
40Pg7G38TDHoov/PaBPurwPdWUPOzT8UWmEM2y92hxQNRr1G5FZ5OGyUFBtHwvD3a8mbIG6vHRZT
WWUmg9fhM42fGh1eoO3Tny6Y6xkb2JUX8O9UWtBiJLyZvFHkL1P/u9ieP84sdrbahjrv/UuWYk3A
drabRMLm4xJMPwdOZ9ZtrHkEeM8r2QJL+tXSjFgvHeBLJjWo8f+bbHV1rhbbmeq9ILu33vDm+Dnn
90qJBgcGGYWw0B2y+ha4ttVdbjZ0YucAli3XFppQ4IQu6MU/68dSeCdcvNqWukt0eMusM8ozkgkE
FfLt4eQHBacF5ajfwbgiZQ2PBhJMCm0ju+nNy9LmvAuL4kfB98zzC9MAOHs6BsE6aGNJzSY4WR0w
lzYW6yWIp+YxgbMIxVXW9kpP9UiwjGtrpgKBSZNm53ECo/PF0XmX0H8l23W7tfD1vfWmg9zmyuxJ
89xpclL0E8h+IqCjc0UyKhxho9l+6ML1eUr8HSPKwaz/vDBQ208r83xQHTbr1y4EfL2OvyWOodlr
gDcJePcztIDCRg1eUU5U6lmnS8rMddqBSRFhqx7y717C1x6rHJKp8aHCXbAwio/RcsG5a+hpi5Y/
Gud/t8qwcNU5JluLSCOEpw65+vrH4zHmbk9SluWv16O3ApTefHnw7LfvU9qbrpfcuCzPcr93RJ6V
Bch3y+qb0uxdEVl4MXKt87T3EgmfGRU9RqNxjgBmitt78TwU9asWDVaKGwlPa6DA/X5MWum6pSNw
Z1Op4zuIyFOc9sOgXBC0Up0XuAAjBqlfr47MGzOw8C+iC8HNk3SXRHmE0WVtdF/6hp+gHhxEjVlj
vyj7wgYUl1OnDJ2lWrAbna9wpKhGeJWZ0oeBsLk4TDIymtANrqilPAuETLJSZ5kNSxS3O6E8mgkH
WojlYDn0zHi6Cm/X6vnwfd631Qi3ChIU0C2tmNHSNecuaCMKn/+3vYvjt5h3YEUD6RwM2QpQRWt7
s6v/JSYCIewZgjcHWH+KrUeG/0zQ/+NN1PV5mfgpUTKsPLkPjiNSMXjQS8yhMicNZvBEiKX+dcYU
5KF1MmfqH+gZiWXDVgH8AdatGIo2AD+jh7UYg8Geg7To/afC01J5XbDmsTwTfmahPRutMJpWqukU
fgGifZLnAnn1//q5b6Wxv1Dr6Y3GULXNj+rOVvcBWB1OWf47PZoHBH8thz5ux0NcxEJeXZVyIn6k
GhmAOa0O+kjFpTrLaSTSCgCs2CtWPA/11HaDguHUBvAZGQTGWXbKCZA8QNduMl4L70jzKdepmUkG
/RaTmFGX5duR1rsOC/YWG2SubnKZIGSJLndUGmh1zJ16DwwiH3UUmOGg5KGDH6TPxV15d/We4blH
a3K/xfNjPCgIB1wUl/1pPC6lnfU/DCimcfsZN52GtFjyq9+e+1CtecB21GReEv1nBMNsUF7Yp7eI
pS0KC9ubTQcybgcCUY0suCm90nxsxaTRnutvcDnly48i8C+iET48B+jm20Rr0aoeCIs5q38cN3t0
6S7Y2v58Kde74MqdKtUuwzAdZLhuFRnhCMdvJppn2VVTEdTgS3he0slUY8wLUYw6ipbpYQbj6Zia
C9jP8WlBGrOYBcsmQLIyLA1X2kpNG/mADU9ZpDx/xk8BZdI9foqXRnEoDUL5wQgmu+1Ubbyol5Gf
XJzk9WdKQlidCQJnbnrtjDe7/cbkGY/Yz0KLW+zX7mluqB28SbFza5Icew5Tsg1MTfmYBpg9EF4Q
Udgn8zoBKAQV0I1tzb7QRyHHLkFYo9ajg4j/G5AclPtomOgm944DNxnSM6I4l744ei7zS40V+vk0
kBiJIIokybTY46cUmG9IS81mqjvJK/LYPf+U4Ue2kzs4lesfq8PD0fVb6nNK4inaTOz/CRO09Kw4
UuCA/4AY08OiDJ1hhFbvadTPu6Q0gw/lQob0z3gflkduzPC+FWQGogzm03Uo6YB7RieMXF4Y1Zwi
JZw1lgNkX7glXRFNWBRSNp2MLeAlRlueyo0Xdkm918FImMh2uhemFuFUhy3xeggcl7dz8KAf9Xl/
HwqfQMKXSJmRQk+pT1eqg8kmWwpThQFSnMQhUgfbTQsZgac0wdxvOOTNsUonO0mXIk6UJZiRkML4
Xs3pXF1QyAYeMEvBqc9/Hg9vtPPQt3N1lVEaB2G5adU82p2RcLyOXofuchlCPXApMIHJiQ/xBvbs
2wcArpumrBofjyUwQ7TZzNzFXxHC1KuYyUC2SxJO80nMgjlTc09rVIePFI6skjLVZAKwgwKnYTrv
K7cbshuREgvNk5wRJcKMT5is8lW1coJz30BSsIHZ7G0jglJdoOPOmLN/sEobwaXzlIvclz0wWpB3
WwOOgJq59tGzVhqtbqXAmDYqDQYFwTJV0Sht2XGhQ8JNaMUt5Tgr/eB73Pmd75DQdcBMWfk2NcQk
KRE3Zc3UnEIMRPFpWpnEph+mdzFVKAWnWaxk3LD3HX5eVG2jeyc+1or5xI34dFc78X6vRG3yKLT6
4hJbfWexb5AFunG4QZ70mWlJkEs0qzomAJP6anoBo9r/ce0ly4q1+qDu78Mj6AqnLFk9GDizipnv
QJy3p8Lug52fslADHpMAuGIMO3Fll90cUW6E04IkxAvz/08COydzkIdcXL9Su91gVUqNdIwJTSOC
GzHN1zMDBq7uIRFM2ugIXVLynmrVQiO3/IX/IDTCyWy2XTLJRDqQJYXFmnD4n/1xFvBBeSssi92W
triyVwT9/GBkE21GzWq4t3sN/4yqvicd0u9NUXjbTNg1E9qebhp9KSWcYswcPfde3NA3BTSPBIvZ
PWlr5wOO+lj2oP9RruePseSVpiM8ievpZa3b8akCoaVETvk6GCmokK386p3yvEEFmlsmJBMJrMR6
ZkxB+EPOh1EPMVzCggd8XTFNYrN5MWi6Y4HBZI32dxT4hsK8wh3XvhiUaO6YruKQc8Byhd+Ykfni
qBjrJyALHIqNUZYDQl2mkNQw4VZTKHbbaJrCN9+YB+smMwz4Rc6dqa6fOhWJljv2lti/a6IZrliy
RuRw1KeWr5vWxoRRf6YkTlJZ7UKXm7E38cUjtW8oJVaKUZMfu+mmgM0sdpXL/GnMYUyM4SnkQArr
JK4IpA+2L+ilrb99SY56+zECYOU/3tpCxj++9dZUIy9uSzD0Xo8U8+jelQ+SDHhC1npCeC5zoAx7
b3Uissf66XgDSP1IpvD4KEs6igZchHXn0KmRfTGcCxjcJ1wLmIs1SCmAlsinS/1DxK9DexRb4UiO
jZDGa7dsvOoGz4WX/88kBpyTBTf824mo4S+aUHk8arqpZ9yCW3yz8v92TlDOuz6RNdxiJWmWO3Pk
+8VnHZ9BW3uh42hC3F5cAiUGlYuJIA1QnUUPbtsZiGkiXEUTbIYG7a0sfDHB8x9xDVYlQAXtiTGK
GNeBiHYSd3c6Aim4xOmKVpYBkIG1ZWlO1VDWk5MRutHWKzCgvaJuUESkmxWyicYDWpMSqna1XSfc
NlqXMS5E2VkfCrTPriheIAtWrwPsYnHr4rE+Hzdk34YjLNW12TA+ecxDVU2hLPW8agPXMojKIoOE
ITIFO9McaIkUoabJ26ouuaunwahi2vz5vcrpb85+UWkSVTCeqS/aL/AlD426eyir3wTql1Z2Gvi6
QA/XVpiDoyXABHv5AWScTfEkt0JALxX2vOB1G34TrxYujO7ATX5fjdZOAVv292FcYmIF9v7BbFQb
iuZlehKmYYuVuGPy194iDQPzI5HDxEkSW/MuK0lp9v0gCjAoXpIN5BUvxf5OVWjLMlqdzh1jY8ga
7lA2n5SuFEw0WpgolAYoBHdow8sOa9dBK3AHKKHiUJvXq7OFnuRKWwaXDGqAUI/CV1F6jufSFdr3
eOoV6JU3HEHeneWjaeLcKCyHkl851O4DsTtzrN2vRgotrqPC/A1XgGkP+r0R2AvNCpfRwdJxKUNk
1J1hTMD5E8RQEeeXSSo7cenko/LfwAvjzBZnNmf+VgzjTpfYr0+0I13Zb3nFufV4Ple6YH/UJFMC
7l1JIfgRG3mZLKbfSXS03ULDULn+tvt9zVElM62ykJilJw+2adA76MMrM6XuDV3w2j66ka04prpk
nadVy/anazz36WsqOgRqtmdh8BmfOSZQnUGzNgaqcWZDtHZuUz6gJYTa+RYvZ+IEXrqVw8bXrrFc
iU0k4225Udq/87Gif1boDsufRXNNbziRMIIlyM8DyTEBcUF7RfLujhVANPRffs03bpEZv/OTVnLi
p0jsx9fA0fKOUFBMLHymTfy2MMZVyknStYG0b0+K6RhDywDIocKgwK1xQsisMC6H5xE/XF+CC4SK
Vgpn0v87P+ULt3A5YJyoyUKtk7s2Xr96+dJZkYHewOwVR7LSUllZC3I25MawAMqOPpsir7ibwCzJ
uq155eogdW6LyBTAvt5hHScBNRQFw8zRYTd8Lb3W5icX8j2XMJI7o89TGolsKBpd2JK/nf9dATJw
c5134axU04NJGqFvIkzmt1BNGCQF5HHdtdO5F5BXoKwK/64FdiRrG2GePbsZzJ4PCrzwRVwYnB7C
qZSuicL1r0nOKn1/34d+ctxaKfuHGDCMpFjSjuGhBGWrm4u+rCpvyS/9WwdHOBQr/9tgo/guf5sk
CRuNKuMGsgVftPqHRGOriAVnI6bqA809j4fEc+RZ5XlURB/cs9ppyh/T3BQLxQESJvXQxjqLgzsp
hIOy2E8JQoxhhZP2oZvFWKuO6UTlo+5+HP3qOK7ec+JHX0vlIJtohN7ZFVzh2kxyjJMI+SueGKAG
mAY1LCUg4ShC5yeAATNDIZZvp3ke9kDu+kgFIbnuBuh3Lyusbmv/AW6JdQl2Srv25LUaq6qT2Bjp
BQ5qISmWUPMiPB1pdZlfM5knyDoHDokAFPVLeqdCl3YyfojPpPV6i4l7VCXPC9C/tZJyt7EqGyGO
QU5ObegZReF/FgA1ImAHbQXwc7Wl0Kk4Tb++XbuqoLNXJshORzkchzEVRcYi77h/x9xRKP+E2A+h
bPHZz1Qs8u2IJf+Jc+iadsUx2k4rclB8GbIw9+59CrL8AQm7RpCA7sqdB0huqbiC9+VWopOL8i/E
/kFzSK6QNA2dcZgrhwbxJ8Egl/gYtgQ+EplNlxroFLlNzSiUUwnp0wuQem5g74+k7+Ta4Lud0zk/
XVi9DBi87U8TFyF7Yp96JHuqm92nWes0tANxjqdhtAY7ZFxU60We80vrhFBVzRYVIcAmbHNXX0Iz
7AngWgpIKqJKsUgzg84K6YzGJRuuPpeU5Q8eqSc4z3Yb6cnxh3CKFmW25ldti7ssjrpCqmFL2Im6
FOPol1naNLdPCw52t3lNTAmg0lCCnosQ0wjnkgbvVu88GC6K+/TUjqFlZd2OKyNuL8nr7wpjHi7Y
MK1pMuzTkcVgrH2qrs+So2np1PVPFNXry0H/DqfbP5yM3ID/kJnj+sKL2+u/hSx7HcJOyrrTGbFJ
OWD6T+9GZsSGNP0bHaiweiqlbmyMx3wz3dmnZMHZMyV2XTKj49uYfWjxFsVcr9jAJsuuxRbxtjRe
8nnodXBpDZj6dXrZOoQ9Exuo3JvkUEuN8m65dJpfETZOLewRq06CcSIRXRSgZsJbvCt/FesmABq9
pAeC9elmhz3VwMCYpnQVwL+PzBmLN5MJQ6QHR5ya1lvRUXknk9OoVbTXDwkNPME216AwsWZYo7xU
vvIC6l1iss79lqIDbYomS0Nyimr7BFYslKne02dN42isQ5r/T0fnOclbB+tH/bzJUBqswEOXAvTu
TP+phjQS1a21Ab44Y/weJ9c6vAEas19GdImL86XHZ6CK2QDSJBypDpFXKQbQwvjXtENF7cVi9MRe
Aww5ddd/MoF9RdtkVRjctBV//SOReMEe1VUcOuwAyOBw/A/kYgjlVrIP2ykuDHff3m5DjwZNr7i5
fUGvzqXjTnkFRHILJAnAEBZIcS1ate8AG7k3VNSDtUYbAr3oG6YHl4MGYar95+N02k7qkAnDSuSV
cNfIyQZnxzm9E3q1o0IbqYPwmTKHk2mpuQrs+MsPidhoOtSFH4MyOv+RzxA8IPrqYL4GxDEEvwxX
58hOriFOMxciHqqa53s9ZYkCDUgJeYvepz47yEtI7qZad70ZPewrgFlQBnibuqhC95SjHGwLN3Ck
kFSXEzJiHq/S52dZm2/2Rm5Plw4PgIpQVRI4QtyVm9byk7Uorm2p1phNraCg4JCVsCKfoBVYPTrk
2fED64gVRYGEn2ifLDgMU9ssgfRjybnRZpaAOKJF0c7edt8v/1TOH2MJ07EGb8hp3+ZUJs44sGzh
Vl3t64+Yi4iNfeqDhXv3pZzJfGXLdFiegqIW02eCb1+WIMofxm4S3bbJiWlLVi9YSfdlaXtfy/tZ
FNj9P8dUYghfC36UnQZ7n2pprdU/v6qy43f0/K9qVKNJDCKy0rhBBuDMJczK+fJPgbeUO5ZqXlJz
Y5p0AGF79Lsyinyi6pPsc2gap/Ui1/VAf1Jft44B6+6dc2tcZH/885tEo3MboezveP2w87PQt45I
cRR+eXHfVdzJ1Dso3Ww5uhvqQcAwzlaazlYXFNEt+AAAcbemhlG7ucC0jLgIlnmnSwiNYnwSqZS9
Ya3NDJZuBRtsGSHj6rkQyDsCajJmGPx2KsJ/Do1iHKQQWfQnAzAqqe34Wnv0aU7zWPL6AXM/chpS
6Rzv/W96R4RvQFoudNa6oVzuybDwI78UQ8pkLdenYB5UpAfIZh89icLcHUNKOY6ILx+mJ099jLZB
EHPKTB4Gg1dqfnA4tuqX7DzCFaTZeqHkzY8tsr1pUKlRw0T14D/gNEazVR7gunPW8S9x1pY5PYUQ
OawrWGkjzEzB0mfpCfjPchYyxLnBiru7oDqVJv/6Etw56KrK+r+D01ibU5o9xPE5yCn/B/d46dzK
KDKpFLN97mQamNqJlhuSZAYtWs1hsF3Ah+gF/UNG8tjy2dAkcYS5Sz8H0Pum7Oh1ssf+jfT9SZam
QUl6byBLZLbjOy7okgjbUtffWTv/dShnjOvViIoaiMfBrjJXYC/hWmfOumhOgfTeAdBqV7t8JAbw
hQV//OpXE3Qtreugb2Zna0muxBbiUcIkb8+p1W1pz0x3nb3IQjMKVVm2/rYaQutjzXWM8P/3JMzr
UTkHLEXtaWyng3pwltCpUhwX8iXaBFUjGO1oMZjukKSB4Qddy83wenhUwsiWU3fHQhFsS3ZOojzA
onbhApA7jgayvVxBB3INtRmr1PUDQMmQuVDX2KNgzo08flQPfaOpoHlRCk1OX671c5dPiOyXWJkj
k2B4wQosOo53Ox/SVDdlMza3Xmr9/AzpIzHjTglgHRt8j2G5SHpRPOOVrID8757CZMKAnoKTlB+P
DdQaW5dYe45TYmyaBALYmgeQy5trn5XdidvKsZntY2tUREU0948ueEmkgcen/Yer0zMF3a9J8Aw0
khb9tEYUYqPk0Z5ekf9Lkys7E5J7gVkv1puvtnjS4c1gFyf+D/NqGXJ/Vd6fHs6ehsi7iuE1pvh5
44ow7inH9fj5HuzDcHCv5MXgu1TUthm5LN+N705Y0y76qOkkK+Awqa54UuafdWeoJEFt7HttLiNC
3U4WUPMvYXggeUm4jqtVqHjy0U3Gx9a40k32lhByoWa5AGK0BDmsjL0KkHi7bTeOAdvKEod6RQrr
jQwEvhd8jShUY3Nhg6q9oFNg8EgLfvDYk/g56groJXU2OFetU4xuPgD7K0/DRkPouFeo69QIHk/n
KO/OdzkXFTk35/+wXZs06Vqby0gA++t4jzvDODCm76mxnVIuYcyfpLbkuvTrc+3FQhJjStT/Es6g
n0yF5S3hjteiImrSFi1goQ+o6iuHCL2BejC+hHmLXlA2LHeytDspCll2MIrL7QE7U8EbQiMyHZPo
iDlC6yfiblSvYATtCLrV/JfUNAUAUeN6q74R3C9kgUbBShr3OszjJbF836pn/mkidqRZ/fyYoF8x
2HdCByWilGXSIFW91tVrfHrzMI+BVLd7hy5D69+zndOY9jAEdShfTJh7j9bwFuBXWeOdLBEIyLEy
idCRIa2EtPs+YfXIieoQL9bkrwSmILmkvlWrns9tGQdmCNwyOO8EkQrkVtTLPYVj8F98pykJf4ge
5LSksTAsa1bzFlbtkerAxTWUuzwCzhmlcZYVtPzF0h3gYu6qcOqMIC6kCIlLBkzX4+hnp0qXLySM
ptPGQjIYZ0XMbMKdKiEIozlrfDnNO/2CherIK5Ycwnis1u5lPGvcVngG5eF/DGwsgdUZ+3qXu+Uh
hrabqqqfMePL8xSqlpq8a+naGT9nYlUuYoa6LFOoWXiSXDwaWoPjgFx/7sjnvDPfozDY9zRzlmQZ
jGdOm8Y9fLxkCgvj2xhmiARmHb54q4QPagZJYHyFU0N8mfcq7b5iqiF2P5W15J0Qe1SpQ+lHqyyi
3EgS3xKs+SkViUGhFskkx9errl4asK2hAUzVt/8wZ6hG8iFRRnnXBmkZPo8YTQCOJ/nlRLr6fyu8
KPWfPWqIH8pztZLha46mVH8/4YfmUwve0xF5i15u4mRR1zM6na2cIDp7+oe1zipGbeN77WLusRWG
ImjE7t98o8jRH29cZ8hrAiYmBCPM+AYHfBKGRsDCW4SPYerGn02iai9RM0DUv05x5fN15kmtRNeJ
OHqL18k4wU0mPTotMoR53iIlzl5w+gQ+i80pqXchSYGUxE3PQ5lDGZixIm7KRzfkUCFVfeNh+4LL
ZA0P11GSEq339Mr2tXEhY1NxdUWn8c58FvCAW4aqXx+ygVCvjCswKq+EX7jtrqGpWMRMse0kHqLa
OuGriCIyGFAqmtuHvBpumK9gMp5mDOiRnW/dJBrqrBr+mz1HA7k/6RpEMT7mvOpobW/tmlK7To+t
vWdjuHmTlKqKSZV5Rwmwm0jS3d/LkqioFQ/yHC2l8x7csuXMOmRYuM07dGI4zB8JLoHYFW1QKHtd
5GX3OghzGCCoyqTpAnts5ZnZ575TKvEDMEzwS8f416jjsNk8THxgHzlqQ/ll+iCXrzhCzn6IxVLe
wFjCD+gBy/aRZIHLhv7pVLuqBN66W/iizDF1r4bi2Hws8sLyeyAnqlb+YoySQZENqsMypp2dzPcc
dIIxuY63DqqqBneaurKfadmabe6RtAU1V2rRT9B/3kijXyp4EgDhcf2UOp1ij2kNxGS90jOu2dNJ
8lNp/fFhiiQ3/QymmPSIHA9KgbBJ7zhtUdMiWnai9UjsVyqi2nrqNd8cGqAJ/w7bMFF/p0EcBWzn
TjfgQ8MgpnXiC4L8YkmQoiaVHsiYARb0MtoktpEt163aEoun/EsY3uGCnO/4m8RcAnOtX/Uycj1x
feZ2fd0GZQu2kaawe57LtcZa9/D14zo/JByISkIj7WQE9zHAttIPBOzRmxWRLbyUeIDwgBjta+WT
uMRz5lXwYrR1nrcI8W0Xh6EJ6SI4eqN6uh8+2EKHn4j+GB3V73J3yFHSlsvPTxKRj4dHn69SI8d4
PTy9/FaUzy0iK52Zqpwgl5eZI/pdTAYCucM+YiHQ4EV6I+biYmNHSjm1+6NuwgLpyzy0m1xlLCOx
nc0FVH4gvUvKLVDC81n/n6l9i+BasB859s5vOlGpo+NX/QUL5yhhB5q6vjBs8uk9oXr+O5WW7Pkl
xpuXt7y6EKCWLw8E3fEctkChyI48AQV1+7YuWA2XYRcbP5UYW10sieR8fBzpZSf4Zsmf+SvAZo2R
ChcWuLfpQmgVX8Qscc3gVJHuRwae9N+lJeTBSxJybRjciGjEz8QcMW6xgpuPpeG+oGUSE3iUYfIy
AtMJs+KbjV6VDSmMB6OeQgWggojX87BljD/+fNqDntWdQMuNG390W2hYNgfMyHi7Rqal1bj86YMD
p5TK2h0nH9K000ROx4ayRZbT8U4xD07D/EvPFdCVcfJO7FtuSeCJR1xc7PZkX/4R4R8NCeJDEWZJ
InzvrnxxvXWL7uREiP2maoYCIywVx8VXdCYJ5djStUTlACgvrwXGBL4GSb78RUe9SqHWMf65ONsq
TrvsbI52sdywjy0lJ1iqUOxEe88u5Kv2P4FLrvxncpI+NuzYPqX8ZQkWelb2XmfCDD4CTbXvNeRO
5czNLrVTJ8IgxOD4s/oVsDnHtlZJYcn2tWW2VeHZN+8xVcX1vf17pQnzQyQUBeHgl9PqLzSoJmrv
z8NK8xH5Am0PekPSAm1AZUYF2BZO63GD/grp+ivWMpYgwDq+J3yr6SoRZG7b2T2mtuLtlRrTncML
RiypxKP7K6fCMErAXy/XpSTCR2l0q9jmgRiJTvymi7pGa1m5kl7RV8jrMQtaw/JMYXEKH/TM4LG7
07dURX6Tot64cVfDSfO5PsqENGaIuNUBW3k6eJtE/jHOWHCp2/5rYhJOKb+l3o55Cc5dyI7EjDQr
1K3HtDdnxoiPteOhrSSk4pA3+kpH76/T6eXeu309nHMmJ6RO/IUyaC1XGiKTfal3/jtisKmMyoaG
GMC0Cd6RuVVcjtAWHneBseyXF7dFIW2hMtTtvz84HVYb1fZHjK4fpYrFEcjkaP3oTzdt4Q8wSElk
an20TAyO6JtTziwpgnK8D/bR/7J5m90rCObhBMoOJPjjXwrRmIbEXOW7byBGgEOfCnjvet2G90Dr
xR4q+yNiXtY8XJETaAOPAxPb4Rsz5KefFHrt2CQdH25aUJ6LHgLVECyfVHiuGIWNqx1LJmdh564L
pziO3HxYZyND/ygpSvkjBkW070dbTJ6g2dVOEA/vxhvnwio6fSGzSbKWYryEYfOJPzYDbYgaZzU+
FXREuqkHPFolnbEXuyg4Qsu2g57J5CBNZecFEUnVRq+sR32C21Qn4CczIWsp0pYpb82iqAoi+GX0
xqt6nCHNhnnoIZjCKkWWfiTawZdTjlHylfYEdJpn7dmMlpUa7PeHkrN/+J19iW/dtxlAP4BfV8t9
oN0xsG0yfjVY8HM/ymJbb73iycMb+PkhRj5RH3pi7xeELVit825Vi2568YWDlIAlxTSmbYy6QdDV
bDAsDH8HnC60DJZixllyO+VKgkHHlVxvVf/+/zaiJvE8BeY4w/J4Ew1DfyKiCa9qjSEojoBp86Q6
hYv0rRMH3xIxowWPvBVcDQd0JdaGPOMjtHSlhBhyfWTkWiE1ODQUW0pILB/wtTeaTeOnp3EwI2Go
nV5ZK9w+BQ0KH1pRaGHrJv0fMXBVgi+3z6y0jnkqBValxxGu06yKGE9qQgJW/0sP4q9thHkoS8OO
f/fuKjA7XloOjHSKa5F95fczLBXuEt2H/XD969qwgYPgIdtjDQGWkJsIPE8s5rhTKRD46y//cFyq
NkmGeOhNTxUUIbCH0lA0S/8FX8uyn6veYyEaRv5om8ZsRAUF7m7iQAcBBN1lLyunQT72cug9J//7
oKRwRTrkeXo6ZZ+vgi+fvqsjkHp2XNeJGSDzi/90mrwOSYL6h750Jhtc1oSdHeG8rRwlLmWezwhe
K0B5eP70WDav1VfMpp2GzC+EAzS2Xo9lE1ElvogGo2UY0iRYlBemg3ASrrhBqK9tKrSFFuQBNsvO
8e3hjPskZ4FzMTpu/z7ByO2Gl6FA8J5H7JRC17tLV2/mAP+GQW0aWdE8IZdI3okb58OsHpkzJ1mx
Z4LwF892gaVS72ZhLzGtf9RzTxMwpqds6hfa2YkR59fKWc4ZtWHClvd64OisZszhs7m7mGTlsSHQ
BYkvuyo0hQCiDIs/4ju8h1ohgdkodF/FtYOgwgPgxY78kmUlJK/jE4gY1DS6K5oh/IkL4bhyGHIY
pFRChHXeqxENItbd4EZhpSsYDMiXyzuSyeEBwsl3zbUwRoCbBNuJFrACpf6ZJVghS8QDHLasNJQd
0jQ3l/1cF/edxL8b9RnIxBL0J1xvSiFyvdJvvNOjwn+nOIzi2n2+0ArTdnQlgIdLlu8+yshGT0vd
Vs0DSD3HGTmOVBQYXiLijMH5RTkO7xP2R1AgwZ+Z1J75rQafL/69fF6qYJ4qZRwn2QXysq01Vdz2
7bstJi/hV9mM9LeWqNi2e7uGVAhISNvWKXDH2Lom3FvJvjs6BVfUYnp8miHg19tz2bgH+Vbrk9rN
xLNklI9tsclT2YqyebmvjHBzcE1n0FGnKYVvJuQbeconz6tnAIDHjlG3VYgsu3GzRYcl3LCYB2P8
hS7e/cFj3omj5R36pZgOMoD6HPcsOCyCEHibgx56Aqxi0xFzSw1z4K/4kcLAxsLBE1kx4Y1N6PGE
sTk1ukKSi4EIcNg9PFuAlFTFl7YMfJRT07TGx77TCdR1RhqnaAVJwjjW+7egSeK0CfkT0XIvrDN9
D9XL42U9K3AdedYZhIfwCbGMFiUWaXEZkvfa1mH3BlF8rvlu/HlsPdI+oq0rNcMW0KOXERdn/jz9
Aub/EPJImiWPiD18ktRyGbl3wt+ZAYWb+En0/6BVzrINVujCggteVn7cEM1JgPH+dEXyJcdwQA9Z
1NSXJ3FL/VDjvno9lT1gia0bZhWweoLkdqtsWosBEtA8w+14iPVAHmygHbSydMrXAyrxSm6c25SE
7RAQisx+6j+oCquM8Aj9KhLA1smN1qxbHMqb+ZEa5hfT3MhD8kF0P67AiLMImzOmb9nF3r7RMubH
F0MwMirqTFqWP4TfDT8qLVeZZwSEg3UZtTQ8+KTS7eflq4sw6IjcnoOwcTK1QkwMl03sKUOhNs/c
EeuD9s9PT3OqYAwBzcE7KEX+rrnY5Xo+90gsYWM/Ik+txWfoiOFS5IKzYLaPh3eiFowuo0aTZpCt
b5KCK2OAqBIGUYMhIOtt+6/jHZ0Bjr4plmBwiVrBkWHQLdD2MALm0Wv2IRSJi7OsXZqmyhl9LnsE
ufpfBRNwe9nmVdPIn2SSidRLZ7zw+TwEzAO0G0/EGubLtksT72xcugD08os5T+ANUk53pPCAx6yt
JugNPqVslU+ispUAxAss8uZaygWz8eXV6EeLjojPfhIVGz7ydd0oLnFBs2aRbFgx57Hc075Sz+cO
pmKfG5tZu5cdwnq8JL6PO+9r3OSZmK7ylyAPaFpQ4W+W87KgtxyZq+jnusR6gM5wV5R6bphGFh/3
Q2KN6vK/KxEQ9m8AEpzr+y/7oCqSfFBP7LXiofoVU9qBzdYqyMO7HdjMBBXkXo3sGAytHunUuYyX
5TLUjdB9YmbvXhlRMyYs9gi2b5cq5BKfqTk9R1gK/5lU/gNClu/NvsNlmvABLZZbaXWl5xhQxugr
/LeDdMiw5X3lxYGu7I3d/tL1PFttaDdSJQ80Lf77C97eswwVbQxl3w+qLGKCfY+xaas3ElJWV4RZ
ml8INUKec5eVGLfuMf5meT9eDwp3fnG+EQIWrkJ1P11Ty6iC4mGt7/rm6UTcpfWH/iZ0F2c7z3+P
fZTod/xLE03PL6dQjp+8gdFXmGBcbFL9u9P9T0WLOQRzzoR4PzAMx81SlgNI8pWx83C4U8aM0aOT
n3nHd7dQzoxJPuhQqAIBQ9UQ4vXO8NMJqbXa+clzDrtf7Sj9Z8/0AXJEWz/VDsJ8AOgz8A2yPUoE
sPb+Sy6NxICuw2HZt6xOVRDinualU8Oq6iTlNjJieC/AsnezMBz8uVeNqFPPtbHrBYRg//iAS5hs
/Ay5tppao3mWkua9xlCESWWI4f2d77A7ycHgaUwGznhMahQc/1X72pOER28EUnXFEQXPZRlh2WVo
6ciVE6HwGn2s84X96AMF8VD9d9osEzz+5izlMJlj35RGaGrFRj5e9pUh8SH0z9l0zyqltrhBJeBs
qQbXoooI7RukQQ+reZNffGejnJYYkQVcSM3XYDMNwmwc0kwEBzJG/sfErbJISRXMFAOxkK9RH1l9
0V/JyxkOQaI35M5+C56EXBE66RwkpNN/OtKgXlG/OJeY86M3LEVpO+lcQygS8/4q4iUkSYpHdOxY
juyAIMFpVaxPzg4lTohZLdDs9E0YshVhdO6+8EiHZBToEJrXLCZJUruIxOmoak6ILgg7ljFnfvC2
tVY+E/wYr+Ci8u6hOZvSRn/5sxxDnCXedbQ5K7iwtX+n6yltWwnxLWmaycsCNIVT9HWv+yn0os9N
ttmDVzSGKUeccZYEuaFRDX8DbOQ/tDW0zbb0aYvIpA9YkGKtLUGJrnczONZflYj86C1jHjfDHYVS
TRZhoHMaD6PwMrWQIWA0ljsAk4PH+pHNOO7fZg0PUa91Ztr8AJ4c2AQ4o06DsOErj69Gs/sJSKPz
wDxXKvQVpxYujnbzFJxFSA+bWK6kjNF7klZSEp+14pfSzmVyrkAehMLuT3kdJrWGup1sCnNCpfEV
QFe9Egu4kskUDDQHrusAtW921piWkVTQdIMHBnuY7SUDzY6aCIcoGN6qbndF61mwKKoE/XMl4qi7
NSZtQpAKNs+tNY4i7LMP9pTygLqOoK6xXzQXBwKhbfqupvaI6BxOkI3z7NeNA4QNPssSBu5x3N5Z
y/FQ8+/G0oC8kuvl2++sWbVHF6M1/rE4SrcMKjDSXEUSgEvSWRqeQagnMFsciAXAbEP3FutziC5I
2DMSKCD2ZRwvZgPc/K1L3XiwIe2HkzZkwqWpdq3nQj52tYZVNe/mcVVnYHzJNFNs8cq4zf7h3PAq
ySY/uwkj/zNn8I6oEMD9ALB4i/VE3jd2006JRj9goGD/VeKADMt72lgFUYiJvv4Nr+N9EhJJYogO
alxUo3Z3dZAP2MDL8XvP5ug2DK4twUydErJEdMutuxcIEKBNyvw95TwArEHKCJFdP2F+/D2glcYB
zW9vOHcZNosWStWcc+1qqznNyBWZHPRQ/lCZirshB+ZM2kTrVRF8Aqu+Dt1cXcz9AFZr7ZsWaLKy
18iUxKZfLgheYz+FdNYjBZqyo0cw4SJJY4neNX7gEHZ9M5hy3ffWLtEmM4t2rzt9Y/ibq9db9pz3
bhjhZtezlfZncfdzqQSzwPrUDCtLmJaT0W0lsnMzqd66/rtXQKn1DBye53bZRCg3bXfwpPFiFdTr
sKvPgtgU+wWjrMt+VQQ91uo6g8Rb4RHFUwjhClbxl35bxAtpRrFA319yl1rLnWTyz0Jv0/zxOSVk
RWIbp724ogEX/uh1Hh9xiOTdTUKePgsM2bB+p350f75A+K7TEbu7aCktQ3DkiEg9Keo7m3MePmLi
J43aWjum8DzshtgNHw8efzjbEo+ELpn3t+0Tg2cEVbKSrIfG4Y2ZJCXnZ9q+SbpcXmpNP1jnnYMP
FAUCC6PSHQCHViexEreD5112Ja+1X0gWJlr3HgfRr6yaImwHrfcN5zkwh4JombAQDlNSE+Ye6rLs
QhrZSrante/aRWnhGICtsBbZsN1wVC2B3jQ6V2Rr+kxQj4yRjdAzacejCx5rmiSmjN+BmFAEb8R8
ll8gskHfEw/wyqAcUZarUcxMZc688xxVnrvlVBwxsaev0x4+17DPH6CbwZUW54f9h/P4Z2EIqcxG
qlzkGYLxOsLNmNCEHjmfWlUS7hSGMQPlwdKWCcHfUlBsiDYczaujshWJqO6pDeKVVC7EOc7uMqNR
ceyokzxCRbVDEJqjN9jnrv0NlC02OIChvqkcMJfc1VXv404Q5qxGGDMxai/gs0Sov39Fv2vLefzd
2BeMOnLbY97jhmc4fAuyTcR401ORG6kZbNGFOhgFL+ICEghI0p8Vv+e/4V3EwsHiCnxK0TDfrFCP
+ebc1wrg+GmRzvcvR1dqOLI59vaUn8bK9jkjNbcHsA4+z5DV+ycjTb6IR2udrVJDSdRHQ8JrwcOn
nP4nJ3KMqpFOnxPpmMtIULFSIaAx4ykffy/8tuBauqL10SXmc3V4yveze42s+i0f6E8JaHNBYbPa
avOyBqg1XZk0/ST5Pj0hUKzQCEjpTruWP06b32N4mwUHBLij5knbw4vS4bx1NyT341XtSGQ78QxU
bFHbFGuL14+4wtp2J7X7JwH0xZPOV5M05plKzEWujSDBl6J8MaaAX4GEvBPgObkhKRFM6JfYE9mb
I1rLVdtFwC8Z7C2dVn33+aWjfdQF5uQchImItpDghbEUOm4beAOHWzhPblcV2lKCYZu0hclTe/VH
jplAXuGEa8cDkc7OHpqFp3aFt5cC8eLVOde26W7R8v4RjKRrhAqVUUSec7C4m0Xmx8qqn0gvRQK8
AJfJGojY7vyO1qF7smcIICZb5v9VrmnZVa0IcXW0NXknsGj5NZmJd1LZWyx6Wy3Gqk0q3oys5tTD
Fp7maJPZ4YVaBAKBJ3HIFJYPXWin7eKYgfTjkOPLKcTbEwEcrTBy2eMt95Y6wcnrWzic88I6DuyW
6YNFBJwSHoyZhpG9hDuvCGo3OAlErqTsXoTF9EHKkXGXUC8CTgPDZOqnQEeQKgdxecxm/jvQGUGS
uuItKYHq/iELGX323zP5KOXdT7ZK8Ao3dUE3RDFMYuvfGiHoFrt8Ue8v0qmltarVMof5KR6TAH+U
iHSNN3jJLTZjTHP/Rr5+rFE53cNnznRhKG4ojo2yG5JirNoHpT46dg5h8dCjHfdo9LVH6uj2Wr5w
sr7wKweXmE9y1kMMSkQhgmhwUNIH25zrFOM/wZrTtvwUfp5Q2A8b+Mz55C4mqeBHUTPluowRug1E
F0k8BIABurd3VGnnM2F7Rg6V+Gr4ZQC5zoTgSW5YmWRBcHzoiGupfkqncHUqe0RRfs7TQ6Betinl
B482UHdGxkW7NQtoU5B0vFI5mbyCeqiiLFshu5vIK5NYT8bCEG1wiq//iSLZpQFGsOBxbVkmFiIm
/t+yV7NIewALq1Osw4gGn1kFFlkxMQo3COsi4PoADvyNiz7yZhNqUQnGVsPxpFAY0RqkPDCP7YGJ
95r2w60W08MqLdIvfzHdl3IVOikqYq0Bge+82w6HLiiN4EXtHcBqAlMkP3x2GG1KAvxIiXyEX58p
7uAFR5U7DQFC4jkzaZO7VkPmDESGSCFiF5Z3gCKThsQargvJ44lkeCIb1Yc9NqGmumJ+HId8dz14
QYiqEvvWoT5zzrDbjKt7vnRNS4IfTRyvfHfaW5xLlFkrOxfNIAYqiOBbzX7EXrODxL+XcB0rRCMG
Hu/znM40T0R1Wm1oBXsWlHMIB0bJejhKDly/N1pNqWE4mjTriFBK2PSxpXiqoLLRrFuTK/TEZAPD
lZToz/ZrBkaFaZ8pr5G7DJZ64FzSzOmHT/GNWSw8H08pWtJ63r8Iv6pa5FRkD03JGs/yuvfL2eEt
Ua7kZFU9ZeS09TnOj2+MgHUldw8EFvY2EhT2MYTyVS5yIjTkOH5jnEreE7Fo8xEHI8iTqYkm5PHf
ub5P41gw8clOJnhcRuos71pIzPZM4CFnHYESkqo+3ZeL2mOfwiNFMNa6vjXhR+JTPgC1WJwXU4Yk
paqPKY96zwDKDRV3s9hrdqE9UHPaMWnfH4GO29cu6iykOwBS6+LU/mYFOoSP/bGLPBgfIIKUdka1
QunX60l7pNqxJ3I2OyKEvoFE8y9go/Ue9e3RAtI7eQdFFNSJhfXJ4s8ZdbPra8raJYlscCvEKVEI
opzWK7LJgwovdyxqxTEGYrQUfA217fRUN2EdBW2nEE9AUZrxhuKx4XU6LppSm+8FyTndZBkYCcmF
fbCPH1WH70GfzO9YqRlf01WHXRBhEd9J12uyqhgoOitLIbf91nhwIMEdB/NIuU1FBmgVNIQF9WPF
L3ocURotO1OHwcg2i6TAYgdKYib0QNp2VbUAdmEgqJ++wEqfazPRC0Ol6dwk5SgfmnQn/GKpFglQ
E0mM+GBuiyHGmKGDfgEqudH/yj5FRttHbzlBZ994Q5I8LAZPXgOV86ng2tJnVXkuaaRKKPdCniDT
nXHosuqUmDBCBWSs+Rwbb9eamkY5GydrX7urpmyQzIRLtoapO7k7zGWgeAraqmHUWUfjj+16Phre
Hm3nPGBMUJAPdkXeMcYrYLuLjeAooIsl0ROqA0VoMdx/KV+qskYr8PhPBxu99jAV9/4cXJ+5Y53o
g3pI4tSF8NamuaV2azxDYNlDWAqtO88M7rSga5XkZDucGBjP2PCpO4wZb7AO7TJW2lGvIpg9I+ZH
WfCqEFRTp+xRuYbn7siq9nG1H5XbzFCltpJS3jbffdTcxxpygYUJONYXAWaPPGAxjzcFPmkm1v1s
YwZPLiSbI79/6MmzjTbj+QsT5chaE1K1EmvcyWCphOkEwa52MN0HyJdnw0y7yr4guuNZiIdO5LFJ
WYMLyzYUAy+0nMp+fKTQHSqXc/Q1EEqOCf37Ch5LxtgX7FetyTtHlQOBwZFHi1npTamQhJfKabzM
qCii2gfxE2gQfwj5zhIv87xVOKNh2npCugf7gTYwOWYyUMnGWbNTMa9sy9NzHAuq9Lz1nzIWkiM0
025oBjKWC7TH6SF4BA8FdaAr+EIRfk8WlKu+I0HbCgpfV+RxtSnFpROk1t5XG0dv8IIFNg/bhSOD
BBhVAv/OdsFwuHbBPVZV1kqlG0KjZe80tfbLCTLdwIjRoZ8aVpU7ZW73u0joKbrXPx0tLFsIhw5u
zU12dZMBl92mqUo5GUOpAj1BrTlYXEVNTKbtlUWZfxLcmE9umv/FyhkOsY5pCNev2UTN3CC+foYh
MwI1l5RhELwK6eg0/bV6Woo+0N2ZKzL20vzIIIeJ9dsTP9Go9/g/zIEDzWfbEH7L5HThPu5rrp9U
Ehz3qL1M01teN8y0a24fBEGsQlGBfCGusz6v1PCQeYlxlrixtx9mmgI2B4hus1aY1vJTdV7kwGS4
eJ3/m5NZNK13M1lVji9Cgqla5FSmQFQyF8m4JxxDuvJ8kMduWp2JpY4enbN6tu5hFnTeZjUYAU18
Y5muywnkLo7+IA3ha24+yNy7TiheFvD7SSuicHki17RDBaPCgWCgM0xm3jdpMGfu7Uw0GFHXVvXS
FurCncGWAnaAhTj+JozSaBDeX0fHZb/S5ppmmXGPKLFtONcc3wmAXETjVHh5HI01rmbgYujtzHcm
3tY0g8OBZq9CoH9YuWedQ41Y/vqZlqT3fU31C8sDfvsQqN283lh1d+h/fdicuW+/578jtJsmUOvP
lOGAjre8+kdjsGWicXN4Kh274AvwtCwP5Btyy7cGqUkwO+cGKjBGovvXztM6M5u1tIK15qvu9s3x
RPvFEiLdkKgp2NUUmptUREO3eQY/bg31wwKCfqReXAhUW6zpGYwfWRnENS5tXfSL5/iWcs2MBv5x
/MTAvaZiBkyVJQ9j4uQVKt2HKhSTqKN6+NtcXvVugKr0FJTz8Ci3MspLyi6SXEFDZ47w9/qWVF50
3wzyht7onhw9aB/pnfzz/AdMBHov3DBujUWZvHjvaHr38PseI+ef+EEkYdvHYBFZ2n3+CvgcqWPr
wFrrTLnKlWvBUABIoHUU9Mvsg54yjFViYn28pGXj12s2iQEWcwn+rcE39jE+F3uL0kJM02ffGDaS
adgQSmmGMFkibiAAA4ojrfMJGus4stnhkR/4MznWuBPxeg+TGP3xNL3/tOcWKiSgwtFV0lj4vogx
QAnoX3ViyZXvbr1r8ZwXKwlhoSxktGDoMPKh5tB3dT2hU7/gjcDhxLxfsXieAYjSZ/pBpRyvtkeD
WFVzaP5AetTce4+8ON5hbo3FTJZH7bNIUhbddz9h6cBN313RodX1QhGyDB0PvqqfvZVBNsQ+6v6y
tmXW1GX96bqHboI/9upcolLeaDd7+ddSlcDhQwbalotDF3gRozOpQbBBKDZh7CgXVJHAb/h1W53e
RcyT4cnCQCaV70ttUHP0hyfnKz7DeKu4wvr/pf4efb7pWAVd78rZ+So7zL4ZLDYMZ0dWHwvoSgi7
hP0rO/h3IkR8YozgVtju0rb5Tn6S7PRMeA3fGkLjEUYwILVYXbZUbszvlYiD3INh8JA/nMY9O4Ny
hZI/CglSEsbTwCVpDgAFcUbbaU6X/fnos9188Qvc4Kvj2U76o5+NkXSjDu7bwXVCHQ9FFX4MsIZX
uWALEPtReQuylw+Xfmw1Ih+2ygVi+lexcoOJRT6BuC21WjxOB/CSpipg2gVcAmaCLCIj7I+xkftv
ZRGEmwMvZBF1ju9GyJ2APxTAv9pR8XVnqj2mfBFzLhQVKb5OMU2xlpOo/WSWxVwHLp+CkBXKWKCg
HaCazyWtrk3IaMnYfomajlMarT9afBHpC5r3kVBcLMwn5eWVl2QIpdeROmL47I5dOUnbphS/A+bs
NZSAZeOvHur1BELzbL//MJWTfXtHWCoyD1ZLQvTs48Ng5Wdhp0PIOcG3OI1ykEiMvGpTFjkrxvM/
kJ/ccGJ4SqQusfeZsOZ2MrJT9tQdUF5pDfgBnl4VMyT1cq1YujQlx7k1CuzN7mRU5ZKQ2ONpGImK
od7n4CFtGAaKUwpADL7ATrpug0RFlDTUdNNIx9/mYbF5kFJo/ezYuyNOHCEAD8xIERzJX0FRCLV0
kn2VynYjfzSBHM4nY0FgKdhWVVKM/2tF9r0g9Aulv0WWtV4J5UQNEUes6c3MBE4ZJywNBPCt9a0K
WF7PNj63eBc6XQxnoFKTSb2hoZAOVQr0r/LXbwyX39pnc+D5co1HRsfdS9Tu6t1OsF7KYAkMHkXf
cJxVJ/K3Hq9P2JcumBfkPFqV2K/bKPxCMms6G0D3M45qyWyyMKIyjuM2mbD7L5Ey+46YGHxm6X2I
MxDkqAx30aGkAQnRp6HqLun/pSRhTPGcZNT0DczDCLpoV2iAK1IwpQ6zrbJ+Az8JN0+kDCwZR2Rd
wvV1y4gTJ3Mz8aWefSwxyI3qlO1e6kJmvAxBiHimM/15emcPJg/lKD60ObhztA+j+0j/wtVGUGxG
AP+Gab8dTri7L5E8xw+o/hSnaPnjsoPmlFgEqR93riBhQl34fX4KfeX0KRug155vGWR6iq3RZFh3
o6CGHX87SJaYMDQXcc0R2HtK2Dwb7gd62DhrdgCZNgMbP/d+trpr4BJE79BfjQBPullNslBYGyG5
JkJ1T3IPsEonT4B7UqvOzNXeW214kDY0IF2hpszQBKxpjbXs6ShbeTZMZUvdn8LHocWn4udSB44C
2QUiuRJffZikJGIWvqXK5moB9YqMOoe1NJc9NoksjNlM1Rrc13z3jIN6c4qh2gqX/xhEuYrl8lNN
xwg6+ZKF8GgoUvHDWyzMI1Kj8WqlgKtmhsWiYz1p7LxglwURtOFaP1gCpO2WVCcEox7yDZh+QsNU
Ci2GalOttCSpgVDAueHjfye/rszlk+2aC8bpCD7rAu8mgHrDfFOUF3lcFbPjFAQwyO0C9paXsq1d
cI2lRHpeJZ/jwVUHJi8BK4Z8RRA4Na1H1KkctWAdWzWMbx1/eYyIgFqPp8Ez1NFyTMqoMQFYiGiq
3YrI+woJ+rlwSW2IzDudmuttiuJNnP+f7XCy5L2FhN6TqB0ojM05vHoYoeduloyLeLZ8iKeCozHP
UOgP9y2fsf1/wAvAoUO2XcuAyXjusVg1gCO4fAynWHHrNJUEwUhp2YmAiYbGXjNH3L074WxVDOhF
7LnKImNcFl+iCDRNJYRZWSQLoBj56ecZoUg+o/pgIt4SdLpA9MhuZWLuZJocx0RZ4g1syCKWRXuZ
yUHFgkZnImrG+tbxlXhRqzZi+3tiRhBS2Bf4UZ/5xxi/iaKNtA95VUKirLzImzZtxm6D4THTnUE8
/7J/d+H5doZ2xeq0WpXcxAzcyli0g9mlkvj8KaGA5JEqPgmDfqiOiMDeEdk9UHCLZjCo6HpopkcU
2fNnv/h6yzFB+1u+rNgwFDJKsjCPeep3yBth4CcDWTKHGCEGqc8d+fl4nCPv8X4Qn/bH2M1x5VU3
JKiXF/8ScnJm9Wp7WVT+JbKz0p2zIFcPfSSrxsh6UIFmo7j3ima5I0wetcpxxYaG4kKprdLVbLP2
HlfzbTk00y2meN31q15GlkwGYWUYnTfLInbzeB5dH8GA3pFbtlNW1+xPGJpWXRcA54vpnHCSRYCh
mvk24e32JoRxa8E1EBuxWg2RQsJLJ7hH0XvNS4LsZzaCCevQlswt6aspqgsB+3fyDHjU5fljUyRL
ShXt55U43+AaW1GSEw2+jxyY3BS0azk5K8p2hBs5haKxwtIFPvIAISYObNzppNpgMKLFIwV7lXBB
Zr7J5Bl/v79vzpCcx2ZyB3Cwm+fSEB0yTQBPEQuPpPt9TTE24Gx1eQJtVbOz3WF1wsIKtTn9zgS2
nl294wKirQ2fFE6dZWx8OUClUQ/RCje/Qv/iE758tkwlN7ZW2brRVB+Msw2Ty1+YQgcyFI9NMyhQ
4kNWDdhdxXGwrsrx58iO5sWbuP8IKN32FxsZDlI4tDc2VWKQw/hz0Cx8DD6hcwzFSHoDz6L7kk1a
XbrziuwroKnXKfN6r55rldmdlvq6pBr7B+8j2XlEsd5LvP/4ljmkl7svfOMpJqRT+s7gCllz8/5S
xH95U7YzwtVnlypHDHilk6GkQtFC7Y2rYFsCntYl6mmNp2PGtM7K0J37el3AhttvxjBhNOYprvh6
7IOVQdL11j5T02l2C7CvKBmY0hwSXimtN20nFJNnxwVYm8WLNQms8Xp9v6/s+rFgO/WcsM0x6ftJ
YO2r1MHtgRSw9bxW2JAsNDdopzPRCrwBPVQw0ZjjNiJcMtzk9nelACQoV/2+/z/WwVYclOFMPUx4
HBe8UOpL9FrJB6UQ35+41eWgDF7JK7eoJyL3XEGnBYm6F5aAL3c23dUUCfT9caXI5uOb8Rw/3tKW
W/vy6ou1UPoVrTec82pkU8lbNH0bxGgASEiZ5FfS7adGNCJemkG1AMUrbE9pTLkT97mSbFYYGKAU
ptMtu8grJ7bqTtCMwlG59Ca117lpJOGqClupAFwsQsVYZBEgomc80JfhjLsSuaoJaXRJ68y+nW/D
uOB7L+mALPhfBAgP7cz8vrgGEB/GYSGYmXvrUcALRrWX27jcpjb5CZaJYfYqQKH0HFO/Dr10P8bo
V0BRVSdQXPD3Y2O7jOk900RYk28UCze1T3J0xF0+ECuB4wKnv6cr0QbxLE/0mk7bCdkPYOUA/cQG
wRUfLJoZfhwKbeSjxvbHOatihdhMmPCwvZjz4BEezATMOnzTAKJmUHruDCR6QjLP9WW+sFKC9xXg
PgoABKPrO+hDDzL7fk2ZpQ16TSWwZON0P7K5p8HJvko8KtuIVb1ye8ZI5x9+rplN3v6gVEXL8F0d
LH91TfvxxDvU+qn3c/e5boazDU9/U6N8h+3L3aoRwUN9AzeoC6/ECQl235VWWJ51hTo01C/sw/v/
fE1EHRSd8i1f/Rkif0i5ub9JYOPNGEG96p7MMv+RLaVrnzG3xQOMh37toFKEMqTHA1l9GhRn4/Il
sfAbr7tzNqxd/LbhJ73n7ZNiN7NBX0qu9gCkFhb9YVlX2iKGTNfUbyss/lQTHed/YslqJIU+Sm5l
UzSj/zsBJxctozDDrFJPXUAmVNd9BcL7YgYgPwfMwiCxGHtflpXbirMeApdRpQ82ERuYn9VWUY6X
ei8znkRKuh6sh9JkMAwbcW3AOIMm6R9uPwYU8VI1fydhaGYlqXe+IiMct50iVXPI2IDScyRFzuNP
FgGCg20XIpZ+cptanJ41ZNncnwRrAwThMSiuxFcXcg3gGFj+p8XE+UOvSrKwmy5N5c28BASQ4VUu
UpbkP3nyBY4wUA2bJlRwmNY1GlCeADdzUiOJcFdvUDdB442iwq/kanKjh/h1zCDNwzKbnGLjNTvs
Mj9OkQAA85KkdoE333UYj/uNEIXKtIF4fTIk/o8tsjRPNmef7bzmWLUAM4SIC7Xqg+ZCKewDh1F9
M9u+e3Ad8+EaQ0qhhFqeW5vtCy6BjyRJy2Yx6ZIYEiqFIdms5JXulRFNs13nn8Sl7t9Lcmrw+Oji
q5eW5bQSxv1MPOhAQjYHGDWLrwmMKzYDoHizW4RXgQc3QptXXhHD/Bp8geou5aTND5+YeTMbFrcC
Du3etuULwHbmvn5/S/E2MuiVELbGgiw9kptLH9cC/43gCapWwNdm/9d74l7QG200pJlQQx1MKg7E
kgqtbxF/c5YvUBgziACWZSOnMb5TsGYGinqK0fsG4KUeX/djLIHO/8cpO+yHZ3BHN2YInkbNIkXk
YooaKxz9nZcfH1NDRxgGTG0rnYPb+8nYoxtGTpwJ66P2WtS9dYQEezfa47LO+nqwp8xopY50ku8I
/qds9yMa9FwFsthigGrBuwKZEQ5cjd/gms1BCFTIlaX7aC7urVM8kqhAKDAu67mBn2HYUb8kZCQ+
Ap6i4CxmcNLpI1qMyibqDwjrf9ZDBJVvWyqnKZfWFQJDJDa3IcJk5e8C6htqfPn/zL7uloV6Pf22
Stts15zNN24OGxUDcQGrMkPyhgfAPXqa8bEQrZoSLUXOT6AnNUyZlKotlLlqdq9fI+umDP0dG5h9
tQo8wABj2DNmVwiCHIcyeTrb51zi9hw/20DDuVmaGsQDF6PSwGWd5cuyP7Z7Kft7mKftMXmL4Ggk
vegHqqATy4/G7vdVt7c6BnrRNaZYsPQ8U/1t38kypnliKQHUV2HbfJpgucf4zglxtXOhCc0oFBvO
ypii8SvGjpjVKX1XYT0Bmw7aaueXRyC+LJCJMMFL/A6isfca5UVJRLnjhbabtqKdsednKbn932RN
AqpsxoyO7T/67AOGpbemgvMlsxQ/QjB2UXsraC1XfqtFDSB83NAgwC4HzQXYqxYb/OvcZOMTCHls
AZP6k4+KoDCMKrCVa+45TQoanmv5WvA5rebXDW7wO7v5XRHr7YtR6YGGZzQySo0/OyDafQSteus4
zzlBl/zsTb35ojbSY5YZ+ZDmneFtGFmoC8HX5GTnElCoaVyzIyxX35NP7NAJy6oG7JftWANU3Se3
QVgxCyOAjqjnWaMsebPBSRMQr51Rwhxo2s2HJR7miH+JMxn6Ju+gdd8vFgBPAMYuwRP4G0KJSwB6
e3UcuM+cnQHrgNJ2cwjSHNx9UCfVE7l9j3Wf888+6ePapWeekSLrU10YmkBZ/H1MeAI6xsZToz+T
7/7IxIymxFiTYT3U0ayk35Zr/l6zThImNfYbePiLIiDuoJYLvGw4sGTgyqEe5EAFGeUXDXAld7Lw
QrECgllORpYxyQEkNp0l9hkingRFLFKhNdnhZxEGT2bFaZEMkjgLpYLCoWhBiYLitoeQgvWZHeLf
+tyE2KTHR96HIilyYViX/n7oPTQXl/zp+tKni8Jdqb7GJKM9WkceYY2j0uI/C9XGD/mCbqI3vZIv
DyULkW/L356jJEh+MEXydo4Mv9OxonhJZDR6UOhFraqR65I4qKH/9DhHn8UVCMsu8NU+pzKsmUYc
hNBM4JFq1R+zoG+kv6W6f4pfA1QZ+8IisvDDcYbex8ttaT0b8AebGC0tNdGZbJGd7WJX4e449ShK
j/yzdCyB/0SRYDl+29QrVBYG8rGsqxt1JLudZMEwxeFKllUhJevYWvS/SpVWpbwdMqVXXkJfrZ+m
IyEva//q2nq1RbKfSrWgNVds2qzrpT4k0B0LeGCbyDzuoSkOsYZ3iSZNAsBoy2t7p+XXzLr/Bq3W
K+1Yi3kJ+VeiCkuiyysMYPBJvUdkPZqroQQmu4tScOlSTPhBE6pdZGO0wKXzbqPin0hR5hs5w7Od
mqVYv+qdfwRk9O/g9N//1sgyTFjcidW4hq+dqIx8wOV5D6PpaklO1N2cYWtALCbEeEzneRC3H1qK
2bZNL2s7dg4aU678h8cvlcxOm5/q0KuccGDxfGo63X+Bv5z9agdKz//eQpfE/p+8QDNf6vAEJaMu
XsljUFVk0drSsoW2KGYNJPChbg8TPRVaNRGNLHWPio2vDFMuZFHkLY28eQcY0e8SaMg4dypJCNEs
cvmqODR6QIykrJUmgRwOXWeHpqMVksYTVXksy3jtnRevLDNVencWM770dsM6KGVheSD0g4odCGbD
7AQM6b2i1LmwPkInbUXno7ZwTtoImzFDDtEggNSxPB2aaD9iMEOwtIt/DcZNTSyrZoG/jCcRFEfN
BzAStNe7vjUkNbqEv02UtOcTM8iQ8IzqN1rwCnemc/w9ERyu3j+fTX7D19aJGJeneP6fDBbjJATE
OmJxaRruPTPi5cyuvzONCHgEHVgv6cftxSpNqUSoH9ixOdTrOQt74BKDpF4I5qZnO3g27t4Co7PG
0VFa8a9sCiRWkG00GyynDazH3dTEKZaposKiDa7O/tDS1BNpbY607mnTFQqP8UqHiVd5eXNYAiBJ
GL5br5NLdRRcKnaeoiL9l0q+xDvbEtyThwn+1yru7s+HGP7mWPqhbiJZ8nm+18E/kI4mGrUAupKU
7fB0MIzOI6JYQKYHS2EhF5feA/VZlc4xttSgaldXYu2l8NE85biZGTa8vPs6GGk8JER1b+uZ8bvu
9TNPcr83AWzd2SSwl6AFeES0pKuNRod0MqzR4WjXWXAgjPZ8DACThPMa0Uq7hQC5cT9SxpBwHcyn
xsHjOwC9p8SukePNnGOLe3j7eBnrXBI/1imOjQ7hXgTEfQmlMambwhAHjht27MqqC7nDQlorwmvC
lW7vBd4ZMo4xWiySr8hzz2lFhr4RT97tpkGNPxQG9rg/mkybcPI64NGheIqrTu9N0KHUYenmF1ol
3A6y0ZCMsvCDTjf9xBPRCkHTaqcLc6rRY2dJJry2el0/oNss6Q/2JgRKZKxtOs/GicsiINoYGzlu
6Cv4QuIKxMuMY+oVrIYSHWEeWWUWCTp1FCIZ9mgcER49i1OAi1W8AKh775al1Z+CGebM1ug2uNYQ
wbmhkFWCfMdc47FesDU2c79a8mMESRxWUO++187Gk1VLgfQnc3Ao3xVw6xn6+d+0sy5UgoqEiKYZ
sM2LABfPGOT7sByYkHbuiUh3Nkgq9V7s2uvquFL12mFw7T9B75VmXXLTNkdCoJZjYHOfb/pPdNKH
RtZbT2/WcU+mkeqsU16S8IbjinvJKuuWkigCpUNszYiLIOxNOddXSn+1dP03n02hftnmTYgiEA7w
xDFOBVUVOPvemArRJDcAOGJvPHS7CDVfGL0OYVazitBTaIwJGpgqnZWWkGX9i9KV+VQymAnpg6fm
wU4ep6T0UaMkhZ8jDcj5R1FZGvJAjrc/+/3O6rBocQjdrkXqN0Pn9q47ic/9yOdH1j6AhqVB69Pz
eX2xYtS83QKWg7NPvpQ94gxY77hfT2qsJ0QN5Cs2tpAeN6WUdSc4GRo93fBhWv2TDmW8wZj4JOFO
7ZMdnPjauAzIXlkauEqnaCL497oV8V8OwDXgeFz5e10wlxPe3ob68D/EPZd+UqPLoiYEh3+W7XP0
ff6EqR+ollv/xSDvRnG8rG45CtizKoxtYKwk0sDSGvJO/7JJMGSn9T8/9D3NC265nGkMog9ZOqer
evN17Ujh0LIV6ss49/h8cWUIgKGJD03FSOc1rKn2sSSRRFmzQRdvyOgXEQBRk9613huGEleIQVp7
PIVDsRkj0O1eZSCJkDZSp3Dh2683cqLAUEAx8snbWXfNQ2ErMVzc7G7jwoal5pTfeFxwlMzvXq3Q
XOcQd5v2XFSdADpBets+otflhSExUbG7Btge5FgenA3EDcil4v2+Ey/jnEsT5EJZ2B9n/DfUb7rB
KVK3vheiIW+Slr6rabZ/bqK9tqwV9P2gE3JKsVeqIg6FTuWd+UwernNWS5CStNUROjlphMyWoGG4
wvrWmsDWx/Z+iaaxfZ5JT0RFk2N3btBkfN0kjrHrzRl1hqBzDCykXIFbTUEmHHhTWwQDrcRL6f1B
JB91TDTvZtn8ir52JusG6bHeVdsk+T9Esf2iuaMjzvLMUquBvZQZJXAIDijKligfwsXsb2Kd2b24
sz9xUAmyWfVgU0l2pZEV7n4bqSLYnFckYcbFyf4ZAfi1ytZECDhl3rP3yuAckwzg8NhY8zjib8De
OaLXn916kqlhv7S4r6koXQzJPogJfSI7c1SchGN+C35suRIyJ8c7YIWCXH+gUy24Lk/YlWPAdbdL
yKR48TG8g0rCiG4NAPAO0j9Myg08W0R9S6sTmL++hS65ifGTs74h7xGlpnXH3rYrJc0rsTphN9b1
WaDMApyIFAIl5ipe0zX2bbTH8AO4KjFKNGs8w3ZQGKZGVIqLIXmPWPZ2v+Z81uE5iMToohNJCXkn
B7CvqMyF3o+9Jz0y4f/0OExFNm+9KHkgeIpNijfWbudC1qJ2pUKB7t8uPtFInuPbaK9vT9CcfBge
sqfoTC/lQR+5x+gQqu1mEGVd9oTSe6g8TtWM/rHUmfqA3xgxVVxJXPHi/QWnZSjAYWIB+/Zxqeem
E0zgbbz/QNkaQaOAyh2Z9Oo+37EDJBLXbJ06qolpbSgj5fYP/0B5ubnMfR7iQb1W4chNYdlpIiFQ
pCy24+M1vn+XloHmyPgHIYArkBLbfGCFOQ1kz2B23Gj8dX9JypYypYIEIh+WakVowkhUXMwQeFvd
AiGEIiPB6sfAF+AI3OvdBNzxKiuno96fZ1NbQeMwGnWyL+Ff4LN8zU6PyUB6rHjaCZ6SiBY2NpCt
u0DKMvDzf77rcrpgfR2X1kGFWrGdxCMjW99XuAs9x8BInpVTlgLDn5sZ2kTjLDU/zJqrTEE9jd4e
ZL9FOF6/Fd1abPuymhPRJy2+hGCnpDzwQvEMj9ecwhrqc3aoAqjuKPn1CQJHU/oNRMrLDLhqVXSp
4T3e7XS0/BQJkvYA6sAReo5XvrJ11xqxFUZttaATQQxlUop4/7vVCCvqLinXnVt+CpCwpbB6P1zU
+AKDFNG2OcezW+HrHFhmSy0tJ3JyGFcEdPhIXMmk77bEwEiggfUCgD18INA0XkWt4idLSsiO9CS3
nEU0OWkilI6EQRuXRc0fFZczhupm4mw76MoKPt3wMwRvdv0xN9lX4z4EL9oPicMyJhqklpyHEfqi
SES38OWpKW0IPFe2HjAuQHaYDizr8Go+j74c22AIMAVZs1pvVGqNiAj5sq4w2cXj4CItX2Ashtby
W6twxXZko4/rW4iDRdssilMOmHBn7ssV3rDYu/rtbifoGc9IlrZbw1QFBDcEcwuerHa14j2kqTj9
SsB+0UrdubycCuGQND0+BMhI0HFDmj4PcO3Aro57bQobDR3ULRhGVxOieKXOBc6YlXMyD3VNgLSv
poRjporLzZ6tV1mQOjLnOFtNZNSgScJeBFTPPDmckZ9pNsU8qy4vW9/IUjMv7UKx3JYQGSqPOeNb
B8Lvwzbz31wEsiCC4E6OCmaQKGBLfbVoM5/SN5IsBIX54cBdJaRQaHP/9G71KbcpiIHjeo7Ryn8Y
0gd5xPcudLEyL2MeKMAURT8UTPX2ZpCGAkNVzBVj31/0BumosAfxK2nIfLJYWareZuye5MEPy4/M
u8xgzaB/kPOqAQpdLBsrCt/MG5iKisqciyCRP7XVJItekZ/h2rotS5Lc8CoRVHUeaXc5LXV1CEwX
cnkkRBBiRbkh/rnQSi2+uZIk2I2J2Jcg+4P1PZxUlWR1qeH3UO4q6JJ6A5+auxLNWpdEghLhr/5y
PuBehpzRmjPTVuBQUfTbJAyEC3Ftipc2+xs8EIeR1VMksTaM7ULaBkxSq5EEw48+gpA2/IIBNGni
nHbebrNFq/0oIB1sla+nY91FdqGIHWTierPgkIj7totESJd6+x8aSIyLcZNa5SMRymv7P2fxVeJh
EsS2cfx+Z5ouf7CYu8pRhDvxd1zFkoKKv+4CmLoB4kWuJbW6offcFxvOpup+Z5AuAPopfpro6agV
CGiyziHawo4qCFdICFJofKmamMkJKeDaPSUITqhqpEr9O33RqCTY3yEaHH1R+lN8LLGNSh/VbDJ/
lHkxnwONp07JxxlILovgCuY1MsEshEtwUPCBxe7XeZQ0XvZ3jf5ADZ1mA+OgiRBUHlaxC5wvyVQB
mZfKcNgxgLbTBdlRHKRTDWAqYXBD3OqRwPJRU+R3TGUT2G4Dw2z0YLAU47IHndc1vFhaJ2q0Kynv
duF0bUtcp0VfjT9kNoEv1/bcZ2GNQSeiJnbVD/w882OZ1HUcYLju56R3wBQukkPxvnk/NZvUVR/b
zMr9PNUCrozOFesgoZ1Qcp/fGpfXfd3V8QOK549FAbcZKRQJtGrfKY3qbN7lhcYwBqrt64HQ35V6
f0hBQp4Hj88L3mFx6EkP81Nxm/isOUToPFu9kQLl781MuoFWNDa1IlMRZbhcVLlx4PXnCC2tvhJU
1ZraFWlkKgdTZa1Hv1K4kDGPhmVv8hL5osYS7X+ERIRgHesBc5NTs/DEUfh4s8R0XUIoUKrY5fqQ
Lno2i+2NkyQ9OZ/DhmXH4p08rN8rQxTS7pr25BhflSN+H9r2Zx34bhvMi/8xY5Uuetkpbrp0lFvb
deU13K1prpAkzmDmj5wvAoSOzBxEPQQkTDY+K+vasoiiweXpSbkivuthpPHNI8ee6RjLZi+4vXuQ
OESzSmgh/VYtJcxqSSkbAVYhJAmS0uhzXVAwASqBc4V1RvyR/wy7F+2qMYR5BcPMvQaymZPGmMQW
Dxp8ddIw4115GlL4Z0PycHlbxt4lrcsY3O3Lg8C8YwmvRfKEJdtSOX1RBaAXVA2L+JiIYhMUpKhE
9rEOtiJ69lN/2ryGKpxnaaXyQKm5hkrmEtm0uIdtfwBN7EM2rorukOQR5+EPdhSpBEFFlz8zrXe3
ERsi3hibBJ7fPo22RW2pvLgG1+0ESk5Ohfn/mkQYudLuOkPZtyXgb2D/wZYyNZ0YoaEaB6srmkHR
sphs4BPWRhvW2sMdDX3jBKncHo1vsxWWC6FnvHxAHO3WkevDPlARYvzmGP4HAXd02eHA4vXMhdNV
7PN5JCNi5/4TE0KyQLvNfu90zUjuN5SweOTc5YXs7ItLg1Ztj11zuJfO6Ifwwpc0CWKrwKon0kcc
2skYKBYshHTWJnYhiUm36vWJOMvVVW/vtjp1iwkTYKcKH9GRBCWT+2x6Tus4k98MdCeuIbZYOFhJ
yMn8RJ55ccyh04IkWG0DKrE9vArQDCDe8t0ZM54j7WXxPGaHt4M3RZcTws2dRUbTDH85vjvkGkBO
bfOWVFHr64jeuhQlQ9Zrx1qpGQNIsXhwtyatT3bBYWjnCFS6SB+l1OuQGOw2p4S5zQe8cYT60iP/
CzWzOxtr1/WMPxWG3Cd25L4h2QjIWImLkizeECtfULSfvQJnXFvM1v25BlcYQYhmj9W5vOSrrsD6
if38guhY1/tru8OocuzSw2pcggv2Sjvj1yvy/55u/qimKqs28biMH5WsjdByq3eU3g+0CDqRxLA+
869saEfgnYyONhyzBpKTGK4SrccuRz7Iuy0NQWc4ZEoVmQrxlNhHeS/70yFLtB6/U81HdBlyJ9dI
BNNnEYz1+PWDCfV2BTFMl2dBLooXEwl/vqx2ihpZ8flgBphfYXYtqBDRJHsmT824P3G3nLa/8tyC
R/mYXmvgFimSF518ZRI11Eb8KIFuMbRV+n5nqhoc6B1zTpaZ5VqsPHaSa4wkqogCEmG5eUytygYm
pz6eJArvKS2ZB4SIPK61JvSviBz0/+kC/xmUZiWyLgz/8UkUWBtvmCP8af6/81u0HWbsFbASIr6U
PFwsNsn4wkWInb5as6oJioMY5tUvl3Rf+o9wIMunVo5EVbwvLJCs+/guNJmiLW6UwaaIX8/3sNfn
ELT5R3tarD1pGxCl04lU23xZuRbCEIIkBnkK6fVrGonK1oshvk3pP2sztN6cDllMfXKvdnFBydAd
RCo1Q9GgN67wy6fIXFYlBiXVYHNAUBxEYwyC5oB2nb4YIrBmmhH1mLHssfxMpY0UqtTIikDTbY8+
v7dz119CyfPUpRcpw0YotOPJzYI9QoW1zhOO6IEiriZtLIo8L1rsrkM4fVBuWVHidWCm5w9/WJ1l
tGQm/LKn6ThyLY2/Mp6zP32Fa/vGloVLOg2RMsF6k4zXvmhhUipUUx1JRTO7On4+IYL14yB0r1Pv
UdAjFQ3PasmyHdUSw55p88FIkqo9QITA1rn6lnOQdXKZQ87p2Gbu1M2ZMGETmfkT2mXPjqAtDH7L
4ut43F3kwk3fKziANYK0miTsfb+FlXmx94FaJFB5ZzBtaDmwhSMGbhMeDBWGpZ2yVbDdZgHDO6D+
HsU/Zzj4/teqSYijuKxv+hVQ1bpwPoziGI18d1og5eBdM7YhEED4//qEk58fbZ7rz+7uj/Y8AgOE
UD+H3t7HCKMXZKngkm1XI7bPvbDvpf+s3KwOve7p1ls/pUmaCE/900Al4XzCieqeerVwMnoYNwNh
iN9uQAq24RLp7MfdJSMBUWOGBhvncK32WM34CPdbNi1ctCvHdTrOp48BLoLnzqlCuhS1x366A+pY
og2U5yb/6qZFue3mWrl3RNMI1X6RVRaqvCpmRn5WcmE66n1rqRJ7jL1nKEYvccRKIcglq0FgVWnp
eaoqLk876wcvEM58aJFACCwA75VV0iB07up0rePkJ1ziDw24JO8gQChZGg9kmtL/PbfP1H+hEb4+
WAaAy+5k/RMj8utZtQyNuyNuSMIkAC2mrBel6u+RJYbPnEKyGS0g/RKTe9mEZQyrhsttVQf3Ddl6
Sd2r9qglgDxajHe3yqs1JgR5burvLu2DJZZAeVU/qC2guFKEij5xI6IW26GlZOM3oM8AZPVBpbH1
gIBQdwDDnJ+S1omvW3rVbk/Or0Acz4srofhY0TrGnAVD8hFzq6TE/tSNCxP09zOM9/6bu6JTvNyL
2LCkn8pXliN08/I5sKQQL5cpZMTHXZszLjxrC7bkcoApMB2b7/yNC3pY+LtWms7lq7YOITRBbqPi
dmkpIzrLY4HSFKPZdWFPw3njFDkjw7J9SdBkcTjU3pU9kPvHEItVO7lhaXUO6O3OEPZlklcCy1/C
058AqaVuZUN6XTu/qQcPetwhBCJHCkeJR3bqmcHK3QKuo7CZIzsl1div4i1QBLTsPmEq9LEx7mfq
v+CKJcXL2wm0US54H7v27rHeqpj2GxaYUCMPYyWpIkHWcRhjOLzynIgHFGJieu0fioXLBZSx1sWD
05+JdbIv2CHnPVQjK1Qacs86+BEexeu9hkvIOIvIoIR8Fph8KHXWwqL4Q9iEKyoqcJSEqho/Agku
eexYAZLO7X//R6x5OOPtTX3691F7z7dKdjtp3DOEwnyK9GrCFMGeQy8ivghHYrwJIFAFpI5MeG3o
7dFqHREZqpZwza4boYaFYJjJkrgbbsdOjiQH2lYx5jt1HE3b0o10JGY9xK0ffGypvjgCilT1LUok
9hEJykK0mAzgmMiF3RumP0zuvx0rdYX5JBmGApy2TH7ZPBx44X28cXD+vtixPAOPhK8dIsgoQMmN
TxXirgD0HxG6cNalpWHIPGe0CHcQlgHOg53U1hZJmhtkL645pildFboHuY2+QL4/8UhSHAHcZe+Z
wcvZ6/KuZl/wNF0tGDSW6yAoEse+N/HDrKZKJeqrb8dOQJgkqt8RNK44KvP3GtCjwTb9JvXFLvA+
3iA1slpxsLlRkfbk2GaR+TLbDBYuIT2dsWhVjIN7vnb8BtUV0rShiQyGj548CbAfv1fitvODVv/4
wGWn1B0ip7f6fLrjCObgsa4PAYFlp5/KgTU4azJRFz/j27bPnmNkLNE2AS55jPNYHU5CcbGA0Ost
GFnKj3/Nw8aSq1oXa7hSbG4HzIyfdkd5YLW8KEfiZnLmgqUCQJwFdhwVilZjrtPGB22MD2dgjgEE
lSEwYYX1p3kydfzrW7t3i8bG6lo61up0v94TmkjfCM/M3Fe82ora5Jq3NeFbm8E+rBPKf3b4+ixh
rh53l5pjpo0A48y68N34MH0QToER+9mi/R1ghVEYaowN05lHYiTX+Xg4ytT+0iPFADoK60r6tqqj
4wv10iBZc5RzYLPgT976+eTLdP5rUC09S8ZfKaApeaKkJvXbQxjIyTtNu4xiCXduf71+h9XBmSgP
emc1gOXrTvXleZ60ArlXgVede9zl/qAQp6IdSkhfSzW7zu2NMNB/FoDenCVZG9QSithZW+6JFzfW
MIAoqjFfbDpnUp3MLbmZIUYl29+8IJY8Lp/zprR72S+dw6XkTwMBRaKQigdJ3mDOn0UqIUgEZXsv
YU186REgA18b8NIxvV0TdH1/UN5X7jIFTKCXrj9IDHSUaMZJDrI0z9vxyUdkCHyemmp7Di4egeAV
D7S6yQcKLIA=
`protect end_protected
