`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cI66OANCJw8fIIQbdpCG1eUZiUrVUYlTNQ823416CUh5RU0Z0lUSscJg0VdsbyeOG0GIlqnKKDcJ
g+441OyZKQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UgqPJ9i9WiJwgzx9hA1QFTAyJQbYygHQhueZLDtbtfbgNYIe9Vf6qQf08t96mKA1gKActJ7BeV+K
6uNMiJfx/3aUXCSX1zJ6wf3n++OQDmqvxVVq3gnHpb+740+sx3yxZnt+NIQn5YfqgmEXSODHM65H
T6IlCQG0Rk76FUmssyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JffVUoJGoNenA9JkXMLk3KS8XcomfWAzcMGUl6pS4bKWUvYmY13D3pemGWR5ICLizj6/IEASX4qM
MrcOHNOZ78VNNGbrwydnmhep2T8HUJ/34A8F6RlIg3EPqaoJseDBIuA+1YYmvMYUPXWmDmWnG1uq
4OVHNHuSMmViCS9G0XZMw9OZMd079W0WWlGjxgCIsCbTxgr5NySjw/l7QR6gLw2PWlOAIibLSL/6
FYbf9Pq748eBFOa73RMaFJULQdNMNcUKu7XbHElWwAbBAEQETSA5PY/T0Ovuh5VWjxfKceXk9gE2
s16k5nL5jvgzFecQSuS2lSlURIB4qY5hje3ZOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6n3r5uCHMurGEnMpYNf4UX/MkeElsrXqvd4MQdfthvZDOuXHZxcs4tSf3laM+WPFVbsOKpN2K9r
vOlcg4pO3R/XBxH8buk6fx/j1Txb83yD004eikrbAzhD/XMeJoB+vwnOXVjryL4Tq7ewJGiuFj3j
3aajz5Netn79SPqpagQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ux6EQpdIiEpdxg0F62ecUw7+0Os42ovKYC5a4J5nt6L0NXwWYNruQn6thnH20HG3CkZMjYPVsVdV
6fsAhKiqralBKaBG/Ej9eLWDO0kqJYBDBHDr1KxCmmsfP7tgcSeensV8aAfsf43ITwJDMIO8VHys
LbnRxuW/uncBTBd8BpuuF6FOlCwImGuVwEh0SYaZjLlAA/zvuQGePlYAraOXp22pKz1CICW9YEbL
RHIga+6SQ98q3/eoFGq1j3ZXVJuLYcvW94K/kJlph+VD6UU5Kix62jbW5vyq5E8KMpqmJr9NNRFn
j81j5XKXBOZlfp+VVqMs7Hlviysaj593wan5HQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4320)
`protect data_block
td5QFuuLITbKOtkE3oI0mKF0qX1YlG0qJOuKpYVLALIRgK2tKeqDqhqWx84hsVYe6J/VgYm1Ulub
f+2CD7mu6C9xJWqD/pIW50Q+pwWHAcoizUsNWlWv/cdEkd96ghXZL8XkY9vTSxkNgxfJ7B88AiA7
hxrZbat9Xl8heEne31vI3pA6Rb3n8TlfUBrKz3DJhn1Rh3mU5N+FxpCC3/rXLr+roUDS/0uwia9+
8N4JHjJsML5xdOCkLysmHKISphIC3QWc6whUQJBh+LDAE2dteTRAhiMNkdrSuY+SElLwGkmyJt5q
sfHqOPxJgVD5eM7qSM6wnIusx4VAkeSWM778AC72TjNVCgJkQkWOioYVELBg1xnEvftRWgZtbAPC
iX2SzqU/y6JcEj0x0eVKxBJfOzMbtlDyy0uA+5rjSYxRlr6o6lunBi75klPhmpY/jQw0ZO6F8+gw
7Dg/r+dIYVCrgtYA/MTfGDcCZiF8o7IDVwDHb1m20RJTgMTP95eLOx77U9KQ4SOIb6EWQRy3tNtz
13HV8I5ZFTw69rjKQg1XpL9zolJzq4yPqMW768ZAXgJKQW/q103s9bNeQpPgV1njlED3kwhs14mj
YN+y/pU8CgwMLPfghKzPQOvwUDIFbxLIscy0cOMc8Pgr/l9/eg+WKiT4MojWCsUAIhHO1F2Pf6PC
DBM+UB0QzhgrLa5vp1Ci0i3SAbiSD8Lbk1uJ1kfthNsdME8jVLT4LVN/CStTFI9cO3Y5r9B8H3wM
gBaSnYzo4GiEGzCyCzJsCa/58fsfQK8ziU6ZsOx673aDEjleRvC9U2LDF9Ry+D9idp2jM3ztj4d3
UffnRAJRLC3b51e/9u1Sxw16TND0LYqsOLhMj9ZF4denDwcbFwjwXnNurHmqiyJVsOpxqHQn8bXS
x5uuVBOHiJfb5McHEXTwU2YdSzUdQ1Z9XQ9CO2F39O9FPXumE6N2AobFhDs2XT3XU2XeVqkDZtd3
AFvAwLdXRHG6tXIDVbw8P7RTdikAnHGgDIMSZvoj0HaPOnnGa055+1GeZ7c1ukvMaZUjLhpXwnmp
2N9ZLGdtkimgD/RG1tUsEFSz4fCOFMW0KdIrqLlH8Hp2yeuX5ugLPKh8iDengRt7/GMYWLpRcBrr
PzHpKPwVF1IAFTS6tv689zS84RzWwp75n+2UeQKx8zk4fKRiiSjs/S1eWYLvQ/lpOlGErv5azHiX
XT8957pcPnKd5m6wZ3outNDVIKxVRbP5sPyshiD8uZUHA1c3MMCGU+p91Oe9Xguoi1Yv10AQtIRW
PqhY7DijE0szRTZon7h35Dsaf8SooyN95GN06P5mwOAlrDQj/d97d+39fvVfC3GsJXy0Hph3IDLd
1XKzsGMFJlc8U9Bgmm6NcbdgUjTGECZnx47i9M3snDZFOg1UHfw0Xo+XWacJO8udvK3+EZap0NAe
fJx/HYcAvSk6iDnMOhOLJUFr3UxYpdhzVkpIENtBRqG/jNiuPMjaxbJB3nsQttSrPzPDifMvkGyu
b3RMyR7585oAZqQeWMQSKMORk8DdPWBgyNPgOh5w6TLO8OM/FuoXvomX9k79bOtpPOtlfyiNuVCV
63j+8xm98ZPcJPz+HezvB+WR2L4edTG0lPKJyTB+pbAEBWWtx9Dkpf9U9rc+LgZuYuh9J2xPG8Tw
Vym99516/NuWTLK5Bmjw+oJtfJvZGutN/gJJkU/+xCvVTWRibfGzk41szDp8U91Odf7Mt7d7Xd10
ymjvjIIRUiTYMkIoqAA/mI4vAJ++TjzoI0ANK+Kzgr9PUndpXX5UttWM4gvAWIs8K3E1oq6m4kGt
WOsquAWbVK715hI5LTkg8SBxh+P/e+4rT46Ygp4A3pHyNN+Ay9UU+j99KSsiUaBtWcBUWZEgnjI5
e+4UjJZzAzP+C5o3++m1kUmVK4xsAQz5d3bnwfnOM0fYrbcGPkljbcIlhsg5BtzmpaeSxhyK1CLY
VocpGh3XvRilgX18k/DbwXjLE2/WsEofnGCIHlZVOBnv207S9wq4Gn4TBgfLvErJKqEgQtVPrJL3
WYGlYj0ViC037Q6nz5NuWLP0wjEx/LbOmvnu4INR03d0xnfBNrePBHRlWBWuOzkRhkAHAG2xefxj
8SF5skwGAZ1OKSKOl7qQQxjXTWwSi4MmA+vijj06mL2Gwr0KG38563FrPweJ5v40Bn0qdCFWUWOY
mZEAUon1fc1XrgIKISPdYuq45q4dZQMkKSnsgrAcp3YPAT+Y6zKgr4qYEJMk/ix1udSCwD99EGca
xYYPkR+CC8AbzE3S2HAgxvMLwFNyO4OcQBiBfZ74r/tUTZmmyENacfUXZ5G08wjdGkw5CRolT78A
dtcLHnRWCArDh2jf+pjZuYVXu7ig/yrHEd1J5+6B0o7Qjf5vYFOK86sHQNvOjCNSxcv0Cxxb54yI
17QT0EqzszxAcap9gt4vxuigGgdJmyd0DHBJE8vT+8d3tYSpGr0DPkNfaQ/qlZzNqdeZQmH+T2mq
lRyamnJ73rocFmAfjsZg52bmD1L4h3HiDoYlA5ZMCPypWXddUlr6RxLNDMU2yE61VX5ce2zoHOUf
GgMij/e3U7+GngH8ALYrbWqAzd/GAUZ9JfY/eJMWhY21hZVM2gMqY9u7TFkGhSWPP+tpK4WiiLB2
thb+v0IhJrVLZ/30YgFsMaaxbP3BrVY7TPGgRcp+6Ihgo5ev/CGUfugUDw+7UsedXb0DyedesFiZ
hqP97DmMghZSRgpD4uSkYecOWmR3blU1YSw2KWshF3eRc/kZ1Yo5NpGtAj6fLxi5fkyQZeGtD31s
0XDYBdn0mYmXKd8USA8HDVs0SjI9yI7QQMOB5vmAZcfdRItyKmbKCeIwr2N/lMo0f/3vh9Dc3/r3
3XiMpFD7IX6eahtM7ex2I40ScWJVEK60hyM7En4Qyg95XUWs0kDeCwo2A6lmGFc+Jzvzagxzxmhi
qTFIj3E5Oxrrdpl3koC46FirUDQQ+bnUZYMYiqu/FrT4okeyNkbgOodoudpMfm7h5Q+BeZCAEoEm
Fwx/jw0PZ95eCYxf8mEbwVDYDoCmdd2/zTXIFS7u6qe/wyZDt7cqe17cmEF+LPfEu7Og/F5/6Odm
spXWLJEYjv0bUcATwTNGFwPx+ect84dichqVQcVw91Ek+9Pe5DM4iqKndX+vrGr/THrTjmxlxtsD
PBcedSroplh8kNInXdccQxeudJPYyh1VUtOmR8fUvS9r06mitJKmvNtjDaMHtOQAJ9MaJA1m1tLE
KcQv4xBYVh/GgUWXyUt4i1jFbbBFK+dUqFIAY2Sv6jfGYhAF40BByJLf4ddhbd7M9vjmXy2kw+Jh
YPhCUS8YquxQaPfpoGH2npQOGDTPR1DgZhtAZNV985v2lG221KCKoiTAwp7MdRb6ICLfwIttSff7
YlJol0MglpdAc3j4PiV89L0YKXbpvwBG8AZ/BSc7OeOHCi/+fdke05LAim7mjxMJ8gW8InkIyGj3
4745G744OSwmmpGPf1UwZRoafIXwftZzJU7HVUvwfFh1lUJ/uUyUKePXCAfRdjfVwUKM85yRemqg
2XIhrFu4yaWMIumE/d2vm5YigA2+LJY9RGjnhFjzLJvIJw4ScgdTKpGYjgQITFK3E/0VqVOouCUy
IDy6hECRGij/irht94sSCdifk3wZW83U0GO59aU9Raxs6WOm2NxHIqZhlCB3n4FxfdD6TaZ2htky
+WfIw0IJ8lq3g7PZLZG27XHlo4Zy86V2zyK6Y72Y8DdARtD5i+LquGbOVrmWJlBqdn7Dpq1KOycU
fm5bH7aBxyyoxIpt/b2MC3Xpy1aAzc1kUEwYEzMJ4I4+CeDdMM7MVo0ZjWNyQr+QMSfxDocUGbgQ
8+a6TOnRj69ATCiEpCkU1L4P1ytgDlkbvhmCoGhiUZoz/W/tb32dd3dNiITvDIr1XdN6rE8HGVDs
H41MRAZTLWuFii1HObq1VvSMj04VMjoC53VTiO6B058kX2DNsRiBEgHJWv8imVhMjLu4UHuF4c7S
ysoU0ckGSludbG2A9CZ5XabUMFBi35s8IMbCzqUVjWgzy9RWRtSZG0uUkb5Hmf+UhWle8lJ2IU3b
Pl+CAkh2hAnZusqeP4C6ZXqZL8DxS1suBiwZBkOyu2xosTStjXSKx8+qC51cIrnvVrsD429dtS74
6ywhAu5S4QKBmZ8z7pe382CfM3QvL1K0C0cHHvpbpev9UF64hFZLIR/unT3T46aPASR8wqVOnZ3v
QgRGen4Sdou7pUwMDY0sR39uSge+GWCAa75yVPa2EhqeATv0G9DfRth8GBDosCo9ssTYWKkMfW7Q
lNDPeZ77rTBnAKXxHyQJr14g60/AQPWX1jz0uhMxmIMhD5PmpWWttJSzhQNJI38zjKuDCibjzdMN
EdhbngCa9P13IipSY6c+bxvwywmGuw8nLe7kWCAlKMy4+Fo5Ml3XyotJANrxOf3VyTVoKN5cqEIu
HgHkZgViBxbIpTJv9xAEMBX2ajqHZyD0wU49odyvL4q9Lre5eN5MUCH+HDwugqFb4QNMFdlfBXDs
LCAhQh8rKo7tQfgBwuBA9Jp7N37Fq4ucGTisL6HcpxUAJwG7+uI7HJACruJC59xoakFA9hFXz8sq
yPWNHUOcqCuk19KS2mKw3QSofkTEHTuCHVUyEizZC2dDICun+fXwgLoGy9Hao+03YMt39UO2+nll
iJAvGte58gEBhudA0CVnNp7i9TujzNEViWR9/7iQuOO6Dt6ZDXjWALIPB2osQN5S4mpxlzCP7Mo4
opQCol1UwST1ul6ajoEpx0cXpYBHu0xjXk07LjSC57KvE1YwQCLrNHFQVPMePPnbLLal/MwWtQN0
QiIzx16IicCG6naU92V9n5axhJYRz5iyBxwXeOTJ7LbceWuIXYE1kIU5eyD6jHyoi+L25b9nIwAt
BOcxFw2AaRB1lYWExArOdDFab1BRRz0KPvRYGoEbCS4/SJbn6+yUl9tIcME4WgfZnCpd0aCpnYUU
cEmVkkMMzxRds4tXp8YVdWqp2PCt132mUnvZ/RNYnNkBIJNOizcLFLZ3LUBZXi7NVypxRnDlQdj9
0vF7UIbhEQ1zwQZ9ozikuz7SrCvyvOz2N6ku95aKE35kH6LeZMAyWT9GTVnaPPdhp69HjAPfOsPV
69gYob6pq6fvGjd8/FjsZFNs5cqP/sZryAWgKh50wYhaZ8gPnkMiNXU/eRpD/mBJ1e8Uu2lMf0Dg
Vuvy7HeaNoCxcq5jDV5kv4lqId0P2V+ilIUmANYt8RHFihNuNlGRdA3++PRuHgE02gE8UIvFQTy6
oG5dCqiwXXadHSksL1yIBnXIDTMNCqAS6Frs7vkyPLi1bO+CsJ8UxYbzgu9GnH5+Pn2+2cpR7g6m
TpjrEFGetKYKsdciG9PSPuwDYsystNyseEDkXtFTsJH/bG6yKAZJAKEfcO17IL/bZUhbNTmlGxSv
Wv3bYGjyC5E/mo4MMF9LAgPUKlHIUWtbjqbcvzD6UzOrwAS3n2pfrkSUiHjA/WUe8G0reLcyG1fi
pdVlYflmjbNY5zj2LR2gN4ycTvqHkETCGFDxIVtg6wSJ374BHvJMWsVQt+gO6MWRr3r9c5RHZzy5
A7g8dcO963BjQN3d5yQVGHN4E/A7Sb60JjKICrpjc/oHwUfhAcO8RJlnDkS6mjh/ynzURFNI7Sqa
umSlYlfSDz7Ej+ZO397/qhy2mmNrh5ShMgGIk/XxBASh7E+/MhTLoZk3flsK
`protect end_protected
