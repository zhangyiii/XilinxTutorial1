`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56384)
`protect data_block
0eB40Voek3XE4QOCP93RnVPhUSFs7gsuZImk0NukmPcoVsXmJhe+9mR0Rh/ZKFkpRupwtPjB+wzq
+iq+QETzGXL/kNGqH9zYkK6pKHrLQqb4XRrIGrPis+mpo0dqIE9Uoct8g8HMTYvEszQQYEBNSgT5
ECf8EDTqrvTtYzBQDOt07EYU7jAtbQ95YspE/r9Afm03a2xP2pXV7xxY2fc7HS0yQGPuLogLx3Ww
XJO5PXp5GN+92vBgC/Y3C1MR+jAR7rQV5XtMaUkd1IkO6sfmj1wyu+QI6d+5z9SSzPev+WuxYUmZ
LqdQOKGEmCnjdp8s6IBITYXjdHBcg57EeRNikeW7qehthYUd4Ur/ia26kwBeZsW+ubMMewcl4e54
UmEzsfnGusrWnRU1yFlYOnFo1pWsZLAK1f3qlQ5qbPKFmx5XVQpyFGtQNqBGj4vC4EAvHvyUKnEm
M4C/GmJx7VGCtgec4ZMzcCXJoPb8QXDOcBgPSTgqxX7gdKLn7klTdSeSJPJ+9laRZShYzY8/cHyC
jTC/cfW3/vxCHv4W7uR4s3UY/+DctanVHkQh0kCpnbQMYLF0T2NUcf0jj/l1V/ks4HesbmFkQiWd
4mqabqnEvOU9xqFJvoy09yWYrw8tTiQdUlEf0BS3k36XSH3O3UiMvjRLEFfqoXassuWEcm9/IXP3
JWsTgXyBSlVvhW55pa1H3rqCsX3dKB8ZQyn5LXoVXri5r6mj2JwRFRphtYCbb6Yh60jXJ7V8MFn5
REO8wILNKHKMNEY5EtX3iz8YWrVCdlGKyPMmIIE0BHOvv+JZdxTrUzp0Ypo2RsbxHT/DbqmUxA2H
5DREmOP0uErGE0AeX0FVnJaQcYdOPG1paH4FY02UD6YLgJPy3LJo6K3MoxOWvzO468z30AbyMbOt
WO+NPvZHG+dgGWTH+KlQ9kZY7RTMPq3tivnWtGqTmCD+RZpe1hxftW1YjepvuWlCz8KiJPbhTAza
ax9Ol9qvLqcKBmrGmUK7FQL5YQkdQoHiedsQ1VEMjbCpdsRMydpZyiZO7J2rl4n8CcKLGdI4GonW
9CJNFf5INgIZdFSoBki1fD0MVQTv7l+wp63HplYtB6CvRfc/bkCDDrgnB6v+KYtCsOYFBcK21JpP
N0FGgekuoB8w5l3k3k9UOwfB2lCNpZCYy8EcbCgEHtl011NU5q/vUqkvvGaR76KCDl5EMeJTeDIk
GS8Kw8VlZCefnA4Os8tnfV/RVOgWhVfW3y7vB4Tcxr8WtGIxLOckI+G59BMWqyq/n90x2fc4RUZx
CBM9rHI8kCaxiBeSAUSacR819CbIrbmrz+Z8pdJi8zDyj9tBcLbId+vD3f4ipDdbNlRqAexGcumj
xTSUH/s6nfP8L0mB8ycGKgoLFf0nFZol9kdEMyhBFRbZA+BawQMhWGrTWUTwfRQbN/lqtuXYw/F3
Ubm1jNlSm6/+ZYPht4UN7hCvREEKec4DwhGcQzdQtt+p+AToB15FYvTF+4JOzAjaccziYa3jvMDc
eHftvL6Td9qPZ2c0+A9BPKlIAhLgGm6SV2Ai0gJ7e6erDdCrxxyawVzBPOTtdwkX+a0Gn4vnXRYf
TPuWePhCOEmBs85dLkWVQVY78XilFcr3C91K4V0dRShXRtzzzHazwgpplUWYAhKcPLHmMydai0zm
Cq+df4DL5r/+fy95TMlUu6AkYgXSFAp2xasgoFwZuI84fQgIG8HQCueQbxYTGWj9LVOk6vzG3kTh
iPZPhPOQ4Gd/qOAeTCBq4paGeGqwV3H24eANnDR0nHbH9JI+L84aYmU9etcQNEBbTz99d6km2JkC
u9LwdQHDOzPHOO2FJP+2CIQ40/91tIgSodLAJnrAScvtPWsIfIcIO2T2ifDv1mx1DFXzPX37ab5x
oRq6SbOGDmBJFsXxFW5ZW8SpaoXAV7xjvpDC6HUIA9PlyYuTGWNcdHtUF1ZU+IcH1Ws+25w2Z0Xo
Vjfdb4pdvAamsb0/pDJ46oEYSF/J4ZWUaQe+RZQlU3sqO1jkMrMieLsoiRSo/qRo0VOjOTRSjc/f
BSwyw+wvKPq6JkDqC2PzoFC/ZLbTTPr4L0mrnpPweRJAyq0yUK7W3rdjlTybQsdtXBqmQaKQtz8W
4PdnFNM6eFqWSy5w0CDOELEQlkB1T5yFSx9ZdOaPldBrPF9TIn6y65N+gnNA9Iz+ReAHkNnvb77t
iAToQKNmLG1hNltC7VR0SF4Igvv3LcDMSn+ZishN9SqUxTLYqzxwyd8G3jv59RkLADfUOj2fGZGJ
IfmhfoinlSZxkLNmMg2KN0Le7DlFCeT5/Ch9hEklloPnTiqe6sHzrAn0kCpshgGEk6BGHc66n9wd
2vRZqyKHMjrbFpfhRmc1CeY6he0EaOZZSMSHQe0IObilKCYUix2lpOWE9qxeau7+TWZ7m704SUtg
7AKmB8InWMZvULUt3cudYbsAeKJhHGQED3WUfmv/qogbM4uR4J7nhN2UKKSV6B9DQdaPO7GLCTgW
ipgzdnwxXDKfzyZD1+a35sS4RMbK+yQtHAO9TsKvbjjPevlk+dfhCddgO9noWZXpoMcRjCUdM454
dS2S+u2XxK78iCE2UJaYHRSR8u39C4V/i6TeaKgVqCwvaXz8rC4pWrrUFNsRjQSdWRfWdx49t2dK
9ExE2UMadsiEFm0IUe6xN+t/RsW5PO+jliQt3L315/8ftDHGFQS53v5Cg3y2REkwfJxj0lAgoeMy
uWFiT4cYvED14Pgd4YeU0oG/qQHH1DU3CqedokEvBq337dXHO6fGYeSD2FB9vm+TrOJyqgpeENWq
QYy2owOWfRGH9atHIhq6hBHZ1VG7ypvKcvUzaua/QNEJ3SJz01DkB2XKwj+3yS4uiJSSXPSJ2CTL
WDiXp5tOUQySoOWVN/HNi2OSbTR/seDyV4BWPTF2umNMLOkclFUEi7Uc1OPg9DSO5hkkR6CybhDD
tBE+Hm4qBmLoQB1YQOkx19urd4bxgRxO66LEAZrJbtXw2StEuCNhWzh0NQqMgoHd7F6XuITLRYoX
WvY0dV2bBWLfeX1XhpGT0PmbLbkuo7hOfxAKfdqFaoykIbsSac1O5bXpKCRiHC47VuKIdm+nuk4i
SCJUZ2lfsxwC81cgBqgbg6r1ghsqzp428EvOP/AGmaihV6rL6fnqY1gkbP3aUZ/a5saGUa3gNjF3
z2KZTnVlNw+YoyIGuAWEI543+JqzsahMk9Uxnhs1qgIYFrDYk+ds5W5tVFADjyVLUYrvalQKsFQO
7i3+pms20kxZpy15lYBNUh+POQ751whSe0bffXU/oxm3wg8bDfpgvhqlTCfuYlu5ejN7/xm8H8KD
71l5GeiuoaujYysuQpW17SISMG/A+dUIgflMx+LGt0Xw0fnSYdz27kulENDJ0CxuePDBWuw5EBdG
zSSHD3/xRHmBOH+UPU3PZVkkraWXM+G4Ce5IELd4MWcpEZ+Z4UkKczYVUumAJlm5y04VDSwIk2Ki
FYvseQvtbEmMsMwoFvn1Q3PJn4YqgyYj8FSr2Yjgqyt3niqEzPvoxo0gWWsYiTRMKlHzCZPmlvuP
JQZ+Jsovg3EcQHblwJLkI5ke2ipyYGLM2xANMOr9EVYZYcIQauAJfDYRuayDRo6sb3KbLBycjuA9
GXQzuyp43tgy4jHAhONgjp65mDNIWucP+H6q4ikljndQq7gErL8xuNRwobYxLp40hDKHjhOYVBL1
RCFMdpR6mXcLA1SYiU4zVfioMyLi4tQC8HDvy2U3yQFPXHX2mUCw4jP1FiBA/ADB3AmPZpOMzv/B
E2RHIdw7/5S0uWm49ln3v0cUqM8IkQcEkXTgapy76E4zOczG5yVMGUyUmhOoXieWAhCJ3+3yI9tH
9ZSwlhZDFA8nccgw1sdS7t3zanCvE4H6joWLAm0B2BGbIF7O408mcVdVmxXa8HQLoiky705if59B
lvMaHXX92UqdnECPb+DdKWlHcIgSIYop+xwEwYmWZYKYAVHYxQz7ex3APBFnBjRF2RsOXUoLkCmw
P5lYhWTar4GMBV/vdZY+o3udigNKe5a7/2SEq3XHuyi1sApa5WQU7zijG5G/sF/8tu5GNwtgIUCG
XWn5apbisMoGTZSoSQi36fQgDrOeKs6pbBpAX+vSGkXqtwuEzLTbTFrda0JxW+CCywg9F0KcfPCe
1+YAEv8G8J4NB64q9+vLf0691QMCxcjkSgxfr0hV0+QsQR48/NyCrdMdi8nFebN0gTTZ9KQTC6+9
aEInzF5F6Ph24bp6mRGx11cg4fDXl2LNPVe/veGv+komo9Mhkhvhb3823vS7iTrTiWWKlaZeIh5W
XaDpQXhM5JS3+Q4NvLoBXEChzJ97X3XQAZ2sJJ7LSmhhb71SCiJ3Wt/LBZREho2ylwGuN4ZuUOzt
lJkOuu2fmhPWovkY5lQH377G4hYwjwAxYWKtZTrLvN2ma0Yk1kzFOVpe0KwaI4Ygwpj+4Tp4jsGI
AXWVigh8sfqtDzRhtGFq8eQlQvSQr/PZ8Mo3lyM7DrHY5eFWZ5ysH9bhHc5PCOS4/ScD2w0rX8Lt
EfVgIoz2lU2C3Q4jE3j/vaB0nCQY1q7sCmnhMCjXac57Pw9jRws75dH37icwvqjtEAcsLjDfZpyj
szOFVeXxyuc7eT9Nmsjg0MyMcIttwzxXfZHtwtVgrkiljNVvh7/02RNzGjsJhptR10LrlQ0Miv35
ynOX8qCeyS/OeF/qTq03NLGNqEoPcc85t4dlAGDX87VuE64wAaKNgoPiChhwqUYrSXpvbDIvUCbG
oSUt4xXEfX24/fPqtgxT3DhRIOYEJpIpaWpogo8MS/ug0MT8IQzob7HyR0lfadZt92YD1py132DE
R4XhAA/+SNsxtibgb+X09PPOhptkNzRsyQl6nm+nYpaksCmtJbaDpmQfPcTZvYjV0pjk9YEeyBGu
OXy7XwOHAmqm7pL+2hmK3kLpeLFq9tb0trC9f9V3mauK/Y/l3icH1YpGhY+f5k2HcbaJLTB58kta
d/hjCUw366XC0I7zqlv3SoUG9YyY8AiPKtjqYK6uc7/NEM1f0N+Zumvt+ht5uhmjOv5CCd3OSWCg
/QB/UAn55RlgVfPz+Wy55rJlBW+KkLpm8Q49s4yEwZQ49AfkVQZ4AbrtZpDsH7qvFD5od4dRB9Pz
A0YIHF7oz6rLkcyNjkBzG5R5+GW0KqktINFDzghaZX3PFdDbFGFYXV2uBqaemqCG4A05rdehNpEE
awlErhvuSAj3NlVhH7Pz9yMw/hFIXlKOVYSl7i45oxui/sCMhHkQhHJ3e69LBHjlfEfkPh9mNtXt
v8fAhmFN3ryftmqJMyXiGMFFG12IN5fLvH58ZEmbb3cQ0n1RYMCgEtadMKT1kSt9mBXCQHFfovJW
VCNDkNxGFm6OWGVlvXWZ5HqoXYwliOaCw7kuKDmA6+smFf1VZK0+uKy6+YjH9p3o0sAmYGsPfGgH
4swA59g9F/+rEYiUiCPMqXUJHmnen/a9worPYNx5c0D306svwBK9cOy28zRk9ZrFcOUG5rpMuYzo
56kEyri8F1o5XU6V9+uuCCwtMRi9t43/Oannve2MpD0bYF/r+YCSErgOc7SkTzgfD7AJAXQsgpG0
Pus1PmsISvr/B8F4rHd44Lmxz7WMFDu0SlWXu6CD8TUQY3C+iMZVWJG2knRd9De26zWYNm2+hPqm
BEVbtkxflc5aDDQpUbw3ZgEb5z/BHkD7FCzKPdJ58IsW/AAD5fipMdehIjfSBTIrrAqGML/zhlep
K7PwuRvQn4rR+lp5I5t+86i8jty10gVAOXkU09hWLDch2qCVX8rphiuz7p+iuHF4/YJOJ9zrJM78
k1+VePRHnIMoNSzkwMMWRCHiZ0P+21G3/LR67UWdPca1UrHYtp4xFi9akIenHvbWutKmV1ZqN/ly
OZYPs18ZvX7C1G92mOqOcuMy7fYl4zBzhD1i0E5WperINrmNaXWgqTy2UmDIQmDMUtTcDg2s3aSI
fv8JxQsHjMYghLRblVU3aZYD3XJOqcePzBCmp2C78E653D2eoe3qHuaT5hv/aLxgFqMxtpLlbKeF
pwrUyBtk2jl0qSc6ugb/ynwIgMLIFo60/WQgm+wryPA+rxJWwg2AZGdvDN+pgrvMixmie+VjGdzD
jjChtBmdq71fiZdhMrJmsaC0RhYE1MsQp8oFdD9+qu4gPb4UhhM6qf4+GUGGdt6Uxj9AMB9Qgmgl
QiTWAI1+PZBWKFENkXqK9pMDG5nGZKlRbVYB2+GWfkMbirA8Jf1rFAxOfM4cNjurw7Bg29Hk1D/g
SsBToTMIxcN4y1SujK9n7+5n5KdD2CX4GjAIsq9yL7oYJXelvqgjJHC34BiMgogFqFJZpFILeCcD
jaABRtnIjBGicAyyc/3nEO1MNyO4TXqws5oAkvyVKo47dBAkPkjvsvOLULoWwyJD/khAexoY9QdD
Z16BYcmqIzLU8wWOpsQwMyNpWwsGr3UTOl1qs2whUkWtkH3Xl+LQOXLGF1FPXKbIzNfJ5skzbg0Z
HS7+4hbTwiyEOEUa83cFkxOM349hiOnIJ5dWnamB0RJLiRGKTCswJ9tpHrsQn81nUc3dycs1EJC6
Q2/RmJrtMGq/dK+XxNAZpl7lYTjDqL5vHX1pUlD4XkTzBnk7qjtVwTno6IPLXaZFRh8LOwVEebZK
dFFNsOMX9PLpBpnR2s3cCtlFo1W4D93L5MhnOAe32kZdiOQNiKOs4Y9wMK8AeOXRHTOxpdjmkKxg
ACQwhxHmqn2RoB0Gr2+BMHiEH1owWhnWvS2Dc6JxWVe2x048IBIPLs0K5nCTnnaCBZMdXxgxznHl
yZjUTfkzXvu3w5y3DoyL2pOHL3LcjmUEpr2RQmg6A8VxHKbFocP02rtx6RWl0CGthkIUFXqztFPK
tKcixKZp28Uy5InJNhP9/D2DmZArucoeWcD2zut8rt8Wz2uZwvKBeZG5TNC8lESxIP2DHysa0xq0
MXewRqdayUf/dOoNCaeJ4dTB2E3QUjBJ58iCEHgbgDz0SAF5mpbL5W/5JU4pVIh8/cq4hztnZGE7
MalaVrlsUEXs5mBsoD0psUn9aVTsILa3uvRhHfsOLvXPr3dmhzdRcNfazxKExBoDaen8MvaScqoU
Fqfbsa+gD7VGhjes1aBTi7wHObZEJr7BJo5EIvcOYJw3BY/xodKmL3flBxWy5GntiW2CRA8Cc8h2
t9VELPy2ZulT57yLF4tScnlw6pV68J6KxrpWZjEH+4kO6wvgxqhMJPcFw28frc5PYeRXsWZHkGm1
BuW+eM0QWhepZiOJDn1XTmIiZK64MXybjwor0CjQS5NTO4qZeGIj5YXV42QOiRvioo+IbX4viUb2
FdlED2CW1yIU7RG2tUYiuHzyv+tDNvWzwcfFHkA6X4p5z6gzgy7WUGwz1TwDYi2vDIR4pLWygI8B
xmhV3iji85NGPFc5Zt0UWOAOQaX52ADCwlbyIvNVOMbEcA4y74AU78USvjYivM10DGTAmZZfRA5R
cap+dyvZmSxSS9vXr5rSydYRcCA9UwWWquZgyMbZL8jn++yoaTGd6C/YV/PhrRpEDvL/kLFtsaK7
9NZDY0104lsK3S03wLmkqf7OBb+Z8F05G1dVy7s8oWk5MO5nPtkvXocsmkohrAhQpEWyTy7mYHOB
n3sfeNw2a6XAVQc6iZtmu9o6EE6P9XdE7/CoZwgZBD4KxcexRWHFLzbNfN5lGXW7IoZtqUhsdlme
ksPLa9OhjBNtrIkjtIphWCEmCQwd9fdLb2Ya+KL4EWtd0zNMH/ewhj0emigIsAEhj/aOxSCEfyOD
UqkWHmdCPdXbY4soRnNPu7/XRuZSOuGLUPnZyErXkuPI5XGwjiKBcZSyCVs9nUZB5WaGIF7Gm8gZ
2CLEKfzgYEhlnH2ysNMWQTA5giqW78QJWUjkvqWJDAjSORLEZyxdqKi2mTjU7eNmB7vox/fTVGV2
1U2ePIb3ZJAfHCr4BkKMSA8ooacX2HBrZuCllTD8t3toXwbcsqxXsXQ6IctVZUZpzHTjh6JxmS00
pMAISr3mBlq2144WzFvKmMItJkXdA2Kpmi/SOpvxEiiJTN7/MfKK+AMm4H/P/YzbqboiPizu5vSi
6HznWzbM3ljgdhmTTj36Bxq1jhxA7dU1ynONjWKG1D/cZ4EFiFMQYVOOSY1tsQIGLE9Ri+illcKa
OfJ8qda90fxpNlRSY1PizucFjJCEcnV2ho3ZdUYWoU7/NpLLQnsB7iT9Wxi7cgDtEbrvGDPVUon6
xWQa14N3otWAh3/miV3eClknk4FDCzm3nZ0HpZc8S1yV/Q0/aoRcjlNER6o9O5nVBi0ngmIB8A9O
ycRmQ3TrLFbj3H0L3HyInzxOgrsdCb/Od1CxYRu4hxB25WS5snkDCXXKuDwPJDGMPBO8W2nU7uOu
xwrTH2e4Tqju56OXmgZHyVkfAM5joQ2442XXyIiBpH7QNeFRGP3VH4559GGjiISfDdfriees4HIS
4q/L7bc210vl0xoFtOgcJ+gm7OLaX10DR7g9JeLf150ZTft0gUNmIR5/lqT6vq46BDgMFpJ6CcV+
epy9UvWdv64eFULlBRP0tqdjTJVlk3PBadOS48qkO9FrNox8d1tqPAzsjTYKPJxPCDhByQJ9i5aR
l2rLjQEK4+bAL8Obnb+/uQcHG+L9duxwXDDB4LUN/OGL3VbA7+U9diC99UuUZJtSprmffUpHlbhx
2B5w/mQwuDVhBgIjp5+0Sj1FWjnokmpnp8be/w/0Z5eYJOQjyghuW8l3I21fvMBn0rxiStj+W+o3
GuG7W4NOKQo1lUXAjc8S1kEknRkDERup+mSDBeN3JwSDba+r/LRW/gq3iKZLEypXtKVBCuDgK8mA
Zz1ww49DdA5Ur1b210fnGemo3R7tMBlOoPBcidUR25XSLhZxpP3sXOC8BgmhORZ/KuSqGGaGb0MY
U3KPfCtBbU7oSbCic/OsAN4WmprQQPhIRRLG4p/YFPkpYXJRDjO8ieLjpjaPGjyQm7HJolVVffn1
F2GthtITRBX4zMqUnpRl7gi5XjEksoqM0OMvMM8UP0zpXGjn76ktwESJQj7PW33/HEyLkbrMpdYf
p7M9LtIRy2plE9xNUJ2AEPj5T07crKztaprhOoI07Og7J8ASo1FurmzA9XeB+16+MnTzjON4iZTk
d6nErczqAHdPANo4KmPKnuh7e9Rd3y5OfcENnh0CksEdc+V0WZbAjI9CvKLePTcFagBlLpmxGFuy
62r37ziNYmn2ufTFsZ0PD8nRXk5SIqRosa7Y/ZqXTAc/iBovBvmeMAxzE305M46ofAmYkXhTRUcg
8rbMbPyr5xeYMzUSPWeZK1lzaNZS8V/8Rv2uTTdvnSIXTkVaYjrUoeS5jeIwfTH+Wd9XsereCT1H
2OXqELJp+hDoPU+Ftj7S8D2mjKgx7wnrqjfAxjPhGLOyi4HQD/iU63Hyx/Uzdm0B0ywHOQOK22TV
Li7aYQM2S59NzVuyQXCH39Lm5Uu3FYNzqNCf4IITqUyCKdaK9PvrD8X7SqtfZdqzkLUNA73xtbJx
4wEljsoqiyybAfOiITwfddqZgVsjsnV0/B+AwkAFbwyLEtHd+EzAhWCc/QqeXkkuX3SgJAwYgubg
5u3cH7GNq5dwKvHUWv8Ss5UgzPw2gKpXjS+Hqu23Bbkyq1+F7cgXl56fTaSeITG8ovpQrAMOfiZK
A0TLahdJiP3NkuhcN1Hy/Ii3H4LeF0v4mQPzJ9s8gWO5EVO6OyX3JldJdZT4g6PdTLjPakShpMIy
SioTBTD3MAQ/ciPYCJ23ElhK4rNEdc7NXCbucETXd2jpge6h3F/Nq4OLxtVr5iY1gVURb9JFCqha
150I8OsrY7ewpsuKrGtO0zJWovvrTbkNeJZtGtsticjIMZE7gMGlv/p9PV1lxoFAafCPFofA7lNn
3EACBVBLJiBPU/wUnQNZTkG4U4wpagpSnfoPVsCwVirdePlep5C6OaH2G3vMttzSqKbVq5s4wIaw
cKWims7Zq27cht2UzUlb9Po6Vrqu7LaxQzki5VDSZJP94WVJ3G7mRS7HMSGl9ZUrbEP0xSs+cNtB
ru92eh/mvC85LfvrL3sbBBID3nbe7mSGunxMBsviQn3kJofZNOAY2xoxmIdOiEZDI3jBtOvwiEa4
2bv+VuoBM9pObASE2h4CbqQkRsWypx1KMOk01u5W+m7XBKo+QZHORt/dvWXEjadcsQ4DlkMyAZ7K
0uQ/hJEM4lDqUDvoHaKuMCcmx+48A767X4lIVm05pvadAuFTAwF5t9D3m/2ZJP0bqZ4XLPvJD9yQ
XC6cb89dcUW61eI/7ikNPxJoh4XiHChxELHbPWd3ISez+FtD+sMeUNZ2YOiUMcgptBymccWL1Krq
8CHXM0BUjGQloMkZbvGIXUoTPbVMrnZ0BVjE0jHw36Q6Ntkcu50TVJg0GlEM4uwHhP26a3DhPPoz
GWoubokU6GEguyxTf7+p0ywIaTuEqTiAK0GCg2o/wq4eG1XTqGIZ1zL5xujwdXBwSSDGL6Umz0zx
7H2gpifLbs1fpjEBYsBobqXTDtVFrYnUVym8ZTiqXolfGjnqwq/JvgbDWc+Kw8DJqv0alJ9SQ5iS
Yq65gP4E0xwP4NGCjrsTHVu3PQNt2cYwsJbxRND0Ii/bFOaq3Xp58qTzvlgRXz7VKU4Pn05Eb8Zw
uKI3CIXM9ui1PXHhYUeg4bIcCz1yFucE12qvg1CU+5KSiAjScLhwBfWpN9xQwEH1kTb4qTgv3q+c
ssWNJaZ+h5sbVRCEvsubBxliGOL06oj1U04Dv+sowuQW8QQLDlxg2+iiGmtBU5ElIuZc+5L41fdM
0fVllvV5yPPuJsJbLRJlE8plMrT4WiBOz2ysJSGEXjdg7j3aV42e2SPIsM3Jrg39pzt6UU7on6bk
A4T+NpjT3O0Y2Hmfc8lcVB5BH73biS37/awkzEcb+YHXXuznSJWOsH9N0aXBmScFf+YnwcYkIQqk
z0A6mKSyjyopLYhWbiLZuQBYpm3tIOHSukdDTLy6QiX6qf3UZ00vBLDWXk5AJCEBzQaM1YTd2fiU
Pug0aatNMLcMcF+Oj9TZbyEceFWxlnHmerPNNkcK1fcq3fquIf2UOTI190mQy/twVlJPLpIPwM43
7UqFY4Qb+d5Yxzh/AmEot4o5A6lTXxe9ZInSeghXMrJev0mm1qifm0gLrUE1GMZ61ysVvk49/YtB
MNj/U+qvnieCXTBjD+6O8BS4e0bnpgBb+qm4TLsVCnSHD1nZhYkruAhjk6X6dMsIxbz1Nkk9bEqL
zDumIhhEFl9jp529OWrvJG4yiWIft1arUOxdVneNBMwzqnTrnyEUYbqPKhL6HkgMmJrclmNfkQEV
o4BXy+iOTqGwdD0/0y9WY5SoSZ3SmV8XaUjh92PpcvNz1kLlVg9ehWbIhrG2fr6O2vI8dQxbWcm6
rYjGRpMTqyJUZaFtQjMs5Qlomjr/l785jONTY/uINcpxu06R/62OFFdRV0VeD+TbyIGXOb1KLScH
vJyHUHygvKXYYhb4Uc6EeCviE9jLDQFCDs1ecutbfqGlkFlE7jrdiAC7LPrvqvSW7rwVixfXn4Yh
RoK9Q2MugBytbcRyQigp+JBVcfbjmzBqjIbPSmirYmGorr3PxOCcYIMNrIiH3tJssXwYRVX+KfcE
bjzgtTg4RZLtyedeKlS/EjnpGqCDfKyO6rlUprO9WsjVj3KffYGgXRIFT5I4Q9SfchI3DR7J4keV
UMTt7KkS47t+IOdoYDnIflAang1TO0e0HMjsnwABt67eUFwAIW28Mbk0+q17+XkLXj5wBStSZxDa
Rp8ur0N45KGL6gAxLeYWioiF2tGf4xn+h6icp76jh0pjD9n5giyX8gV3CI0T7o32TRyAB758orX7
0Gla1ZE2aDvWcnamQz3AOvZFm6c/XoQrLuBS0ZsIwMMMBVoALCPMLupvdiMuFUotHg3V43HF7jJ9
yYHst+K+bvpTj6J8ZMZGNsJHTTqaEgCACZStQhKDqxf5xRM4tQcpzPgcXuVkg5aX0AkPuG3WHpv5
cYMw6YWaLqsWfrm0EVQ6ffDbtwFEbnQxDCvrc5LZO+8ecAe4qSu1O3Wv3rR3t8c9lbCNh1d/aPTK
fsJkFh42N8cCB82gPPoML5LggIb/Tgh/NbYwkdCFTlnj2nzdxME3egl7a+GmIfY58/cjHi2wgiRh
7yFEkxChvYp5i3FfnRkJ//RSMR1pHz0YLIwnyiVlD3kgW/P60xSHSpD9hYfiuHUCBvuFQhtiEuX6
/1k0oEJE3AzQE4FWjoC1X4Dh0y4zkz+uqxnfQI9AWKs9P26FQXkN98zCC3joNzxeUF6J635iCAaz
k8Z7vhCl0JnNGQyBRJOearuevLhmP8vZBkQCIJf1avPK22jJgGMIJopjp6WyESrEKr7vJcT/dekg
yTBlw5Vh53SI6uBf9Dpfwwn0dLc2n/AAoY0CL2S7wvPswqT5GLas012UJoM8WV1aHZ3ggIYeAG1M
LqyjDMwCFCJX0/nlfKRsgmeP3KqvXfEQDf5rvDmCRBUQAOzoKzfLCV2oBUrpa77QijqnBIPDJ3V2
FxZV7ZmQZ+UWao1EuQb+ldVL7Zvb+rqLNt2LgnQSGbuhrwVxGWehdx3a4ZQWh8ihlgQcfTVl3CHy
Xi3Xv4jp+aF9CWN02abF1e7G8ruRa9ubi4JgC70CWDXD3atXgroPU04jWE2zXsq1phvQsty46KDS
3TC+uQkflfRH5GV6/hehOQhI8eDMtPpxmVS54VqUOrpB+L3JhmQrGSHlUfCo6ynKle4QqL3SMzIu
o1WBPQALsWr+6QJBwwJL4HPoLD68WjzEUirsGLBsLjQad8l6Jd5dmOZIFGLSeNGRHZd4ajn6ciB2
bAFAA0F3KvhP0m0oMxzdCvbMjB/lsJ3DRGkDi+UQmRB63AK2vUVhSONf+slc0udx1j/9ZMkLWngo
siO3lHiS4x8U8JxttBzgPLrkTKrl/iDYSnOLPDf+0T0n4onJuN/gtdAtUAfb+FD4ndUNyUCD0H41
FvjLfqeLCicd5OXwCXYtCvtg0BZkeuy6cJBCTqPvSCfGrxkmCx2eIT/O3WINeY0zsj3bS4FKheDh
nteme5i+a4G3DFCvj7JsqIGd0XhsC6AEOSD2TdW+d2zBIvbOxoDEaEC1avJDyzgf+xur9SASrVIQ
9xYcftqvEV8jcS/ZN6h9Kp3wRX/kgORGpaCMWFU6m6PcNS+BvfpI7XCWoY52lGJKrriWvtdGCSSs
yWnUZRqDzQx/w+072CQsEuWbju0cI6PO3m+PgNRK2+AgoQO3L6H0PYpogQlA6lIZCrp2DNtoCR+A
zarYJ+2uwolM3Kyk/y5Qy7//ArvqW+oMJtW7uIwhDrEnP6WAIZ/baRDbpuyTtM38X+KiQvyowMob
KBdjkZolzvmvL8zONIe3z1Wv9W9z27YeK+n3llGVLQ6wHaIJ7NOGpo4JV8bNg8Vpa5XBVPSEhZsS
2nEbTFi4kDl3Y3M3pMaSrihgzPJbx7QxGnt6D6PCqy3X2YLfBEGksm0iR1SD8cnZENiu2UifDKg1
o3YGT980yT3LbVknxhqVyTGS/yrYSj0O8vSdJCPgcRO7cIYkHT4Ti3RUgXXb7lv04JFloSULbNAd
bMzEa/S8Da5KZkCSYegv6LfgW4Iofe4R6OL0QXNi1geA6nSZRVVNT/mf+GsGHrzs1p1hKRpqxNhO
texEVIPhytmz1yd5Htwsjc2oQ1Azg6pvX7ysiRDlfGuj/iiPk/HniJJu/916mPuZivpol9RofdKZ
sGJE7MmVCrpywf2xyU6ADHJZqAQrosrU121RRJ43kUaDoDbknM/i42/JkwCq5oEBUWTBs6FbXSrY
bFJcYVScZJ/g5G+qS6v0xnsVKtmdOn1CFb37q7NWlRxmPH/t+wI+OGBNo0C9NPtOlWXksZjI1Xlq
CeMAnuzkqiaDDwMQzEwCsKlCDYnd40/oWn5SZ9375QIgR2CoVs9YtdJvV/4KzKkx6Ry/pG+Nai2n
i1gPTec1V6iVcCGFQAu7vgEd0iFPNJzx9Y9i5ZlJW1o/bl//tf833WLU9TUoLwbpr/2XfEL7mwZk
n4vgvhWLtXcJG5uSS4SXdErtqvVP5MI8IQTdqSOjCvURmA3WZxdq26DFXpB2qMTE7pOkqiIDsUv+
UYa8Trqi7nGXUS2w118Euh+nEGEa+Ya9Yo+7s5sfQe2ROm213kzPtzaYdQqdSg6tnsgFoavVIk4e
IM24zFCU9LaRt8/Rq7zadl/aUK/1qnnWP5TnPuBEAMMfj3JACXXEcSDw76DKHr8BXCJNBvPLwobb
BdHi0SALSub/MO8JthEfRoWqVFXwrZDzJQzPUypURgPjLeTN4Zgfza2NM4gcT8yOPqpx9dU+CYQn
1/jiJTWkYyRf8YkzLJktfk955uqpe0uGjy5PYvwv1owWmZ3jT2uOtKF0z/2SQxaN/z+Fx1fAQwmP
zP5wKxmpgeNiPpIS62WHdMN/VG03PKzav+vbLTGtODKLbPSO8n3rRaqD385Lldvm9vGxkUE4aHkY
dOXhhlZw2xgvoA9B9+/yc3FYwuo1qM+u3IrCCYf8yb7paoDtNj+6V1zhYaSrXTeSz4yJxRdjGUC7
DBXXpy7uwPluK9OxkOezuLbej8GhYEzraESNogW7GVqpHoE0/e6KNOrbIGp9RbDN8cTp/kko8ADb
Oj2DNQjvNiggW0M+wwKY70GWW9Ns/A9SP+EPZKMQVZyw2ygweXbqRQqECaJGqEqQhWek5FkUn/BU
GbQl5fn0cmV1F8TiTXQ/6cwZRSPxMurVb+Pq5swn2BqhyhzxgHqE0UImfMhIXcRc/mpgVHacOybl
E59WqIlFyVYNaRnH9W+AmRJG1L4D5lUa+jHlYrp7umAG/50yPaGA1tDSA/zrB2rQEE3VvbhMpXLJ
xNBqbfJQKROrSDQbZuzoZjak9qztPIoK4tjc33FG2BPI/FTMNMOtXNMBq6jIDLLZmHbl88uR5mjF
rmh/9bAAoYkLW+t6wpZH+VEOSC5XPyuLGVqH7iKpZu9k3+a4nbHbWUZ2xH8Qe+3J+573K7h+JpSO
xGf3Zh+cYjttF+8UfOVCoFcZ+Add32ZAWotVQx/8z5g2eRCzXFUg7r5+4RFJKam2lEepXHqkyu6l
N6DHUBlOhOWe/VzJJFEAUIDXgFZU8fIqj76absSD1qBW2mj/TMujyqGQqTZHL8zZHUctBduCr69K
+03ktxsMBrX3kBDaFCSoIGFuKau1QyMFzu5xusavcYGVgClHU39BYkKTUrG/3qUhXbSDC50CMPqh
N3VovGvO+SD9gZNTskc3IiMMQMuLsy7NkzRt4eWXs4pOGCTE9Rqce3L+A3toGUKVgsr/sokX6HSl
6gSIPjiU5iZkOHcbO1qDO1IwFYuozi9vIKuxErGrVGP7bHEQ53OaUxuVywJEWZZZX6d6AERE9MZK
W95zaqi+fJYYbmxmX/3M9owteOv5AB0wEoktpvJb3sczk03sCX+wA2K9ZLaErOyCsVED3DOQ3whE
pr9v3sT8GfOy9XhWrETCxWxkThj984F/rNPjJGA9I5Rcz5+VTLy1z5nuV21/lZJxBeBtT5J0nKmq
uoTbAkru2SUoT0jgUn3zQCtznjAPcvqAdQHm1HdWYL3r8XcDhLNSRrtIQd7QSjyijS2mLkq9spy4
IjoJr/VhKIEO4Wrg4B4wiflNzPi09jlak/SzD8vBSHxbFVa6UMCOZILV7sUkxIPiwoYrhw92i1i7
UdBs77MHy62b8pOrnflG388hZe8IVb+8Go/gkdJ5n5P99fFZ1m3SwlkeQgZzGmpLuvJFhhzJfFYV
G7l8PwZbYikcv9qAKc1KO3Jk/V/zu31J0S+bDrNTS6vAYgWM2UVGazSHnpo9D2ZcdhoTSznDnl4Q
W52lH+LGmij1nwKC9bctmUxJzSQ9sG/DMnOQRRx+61dRfcC28ZjOYwCTY2FGnFuj3qGOh53lRXV9
13PbVa7dRPcSWuU30YcSP3nVkptCIu2071jbsi4ZFjrVkF2m3lJcW7bitcg9lSidQwrcCSGwc4Hf
TP07hAisLKffUKS9DbgYWG6bICYv8Q+CF7fwq4hdVV3ZKYV6GMDu5ENRMoUNciirPTaPwdBpH7jR
cgmeSkcW/uvVbwwB+iZDeUqqXXkxlDUprvSjAXIV/9eVN0I5sWPH3DgiA67DNdTCUm8TUutzjQyf
aOn9NWUckgddo11JFd+F8JwNIFGlt4yaLX7Hrm6LF5/1s1159aFnkGrOVlLhOpZ5P3ebwunhReaC
Sd/aVNUxZTOvOrWqxvY4IeF6vaoNiMtV6cHjBbDFzDAr+nfsbqcboNy+U1Ml+tkUiN9KSAwA07g1
ImKgPhup1XtvrjmXeqbK77QUeQh0rlm88Kteoi/8Ie1vAxQSG+uf+4oOzGpXSBaTkfCNKbq8py3n
leWAmotZ7vb2Tg74OpFo0Ns4Clx+wk7WAcOLjjBJcJN8D7TWA+puM91IZ5SzDhhBBvL9zzkoSPg6
pnyvkSvJ6wAvrrz1cjlhWBOz6gSsM+Sgfb36gH977rByuVqGwqYzmzuzM97qDrIKmUj1grmESd0b
hTDtRST1RlUP2Gh1nYpXq5eO8ngEnRNKZeP86Rb0Xs95ayNtM6uRDBdKyCWKRhJp9Qc2kJwxQLr6
aNbDjD1H4m+hI7vMg1GXr1sh8ZdZNHKP3WmOVzoxVZg9FYZBdjhSQSq3qr0C5DK3wo47ko99Fbbn
hFz6zLWvbK2j3njpZwO0qTyWByPyqWgoRh9DLdBDF7pfdIoH8xp4AajepGEjz3LRFe1jr/hSMwB3
SFgtyDq2ootfcSUEgiiIifNyR8acPVAfSCoMj4ZT4x/eM3i77F4a634qv74SMBEkkbWNjZqIFvoP
E4GHP83mLhbYhOv6TlYsCC4tirPLJDRjNoPQG8UiJfMCZGDbnhugUH81xgyObhSkAoy6KqZLOhGT
do4l1mgYvO8PuYH8tSOSH377VsfN8TC3AZ4rr8bs3GRAsZW7d/p9/Lq0UzxSfiliz1PD1H43aFAH
DYvnQ+R6xgWw/od1oZbdJnegAM/1n7IyLbVRHGIy1XBKkah0i1qgkv5m3FKJpu2xo43XUkqs7pKJ
v+NaGSbF+QHk2t/OhFsekB/Zq7TiYKLnEWcChaxScHBMZaz6ApMq5Xpj08bj/ZY7ut3ZvP4TInTa
45Gs/GcwUS7CVEmPtyPyGcBa4YMB/VCyxn51ViO4ekVpK3+kUoX32ulmUPuoHvF2+Vb0Q2hRwpE1
x74tec9pxxMj5HI1xszNPUHBzSYMUMC6n9Ph6vwh7C6DvGKYBC18QnrRcX19WE9m8J3tKu72r/cC
uPf4kDNeOkXTYggM44nznpqPBfamkRj30njOUdU1RRLfFTeSctWL9uLF+eCFEzF1egzoy0LEdx9f
1JGZm99/SXEHiFEwoVD5IM3KpjDKyOgxIU1uU7ySmdUQWZN8YXdWtmtfR5gbqe+3HBRbjETuGVqP
ABTlMTRiEYrC/qbpiRilLAHlwFrdTkOAjzxC7IICfpNIKps8uYP3hlNLwnOK1fp6hxiWyIfvecBx
n/v6ottMrB0kdHBnIbK6iyxfSqbqN+1Iub4xuzGXBo4au+Vj2h9S7/l7E+eSHn7eE2vxGUAMopdH
MIVUduPIWoZu0X/1FBZnfUtaemFTDQdThnqp1ZS2anZHC8c5Fm8DJYZg7HldKxaHqsevxygHPP2p
NF5u4+jxde26PbJ9t9QrS58FDXHLFdQ+xRoca1lK6PwnphgI4Sjwl1ckwg7hfY8rqkrcPS+uGTUM
mv6p6tvKYo7U9rRDaWxo7U/XU1B5/11gIvO5PekUfMWPF4k21U2IPEz7feWWkAhw0CGn7O1lsM8T
hr05ZUXfn965WEky3WWmsiugRBh4lZKGJRKEj5zkTHQgnMZdEFiHm8ot9bTRHy/sJOlsyvrCW2+1
azVIF1LJAO0+w+Q0Ihtf7pURiEhMtnNxgZ3Ik/UZ+1U/QYQlpW/dmGLMqYLJ4jHFNCv2vJ3OJLby
n6LwsMNsHnkkG9k5k71Ip61jv+5yse+cy9SuiYamID9CYDC0nr5FKKkkIFL76/CSR8wqcMCexzrc
keGmJ0U55XlCzMWdB607/jbNcwvtA0Bzowhj8QBW+ez6s54SIBBb7KYpD+pOqJN83BuWkvvIOaNT
mDdBRYgry4ZQnVJKMYAHMeVNj1+XkvjExg+KpT9DCSQFZqpJfZqZAQ73/Cwy+AFmgdoG+ASISKWo
3fVSY+n0C5UDG1SJKrTcS9jiMDyC3zTD2CBNy/2CLmf5I7OoTFmFsqykL8ia6nQU594wqPjCpIso
+p9EIQNwZJ61TIWn1+yaD4a5SP1mQti4BB0Q7N7E1RDt2VXTgCOhjubvxxXe1P4eAd/lz9vUyaK2
QXrv9CKAdG/5u3EgRHC+uqbtZjBKd39k14Df2v9pMfcAgpK2M/PnUEICOcWBSl3oFgy+Y3QauWPQ
s/ewfa1vVRzd1i51aWvY3/k/VHegoOP+wn4NrluVbhSLXGIdc4LVpyP6NLM6VDJem6bCMCK9DtJf
Zh7Vn+B0OXQ7D5QCeKlPjMtr4FK//KUmPIBV/Qcmvhnvs+83W7xwh2bTecTnVbG7cR1VwvNgdzDP
TXBaTJp4IHdC9IQ6f0cRv3YJgm/KFH/FxIqW/6PtuvfK3MtzltJVQSL0iMSPDJOhRSpRSprzW0sl
9ovp96eCWnSZfEqoATL91/M96PHam7brz7shvzL1Em2Xyy1W+akgpghPtaxzJeVBAybFzaZ7qyrC
Urs+mYAJoDHTlI6WDWhK4DYTZmC0a9dZSDQNHawHReHJj+Kj+UgT7fXDpgfuDYAAOX+bV6gm1KUK
v5PD7b5Qjh9Rxqg6Bqd11BWVhV8dZmBmBtYrh0JU5yVZmuI+lbYBnbxcBXJoywicZsOpzSCQxUxQ
LKKxopgjIEBQNrHxyH3nb3+3lCwFqBKg9BSzKjnB04SNfdDbjqFnGovBVPWS3WZkoRFNr2i8zuHh
A+teuyItUgbIrUwy/nbxuxE5G1Qwg0v8aGs+qSlj47u+LNF83cqc/YmYpMs+KJuHpnuMwRhQvS38
MQsEJYqq3MG9uE752f3EcUx+uN96TiiWzOL81riAmQtOFAYHsSAUEJVBw+vgD0Ww3Zh6UR8+tZVp
rHtjog0bFqpiKh100CckFBIWmMcVl3U1bhMDhtYsZcE3rBlnlbEjj5/N5wUBD5r5KB7Q1hIz9EXB
gpBmJjkCuIMQESxw2zqpeNHama1d+PkfwYxrXHiutJLzGv2yRk7ZbePcvAmxtu68p0+9gSH0atML
CdYZrPos00Uxm+U8gJctBjJdiBxRO2Rj/3fp+FKDhJjvYQvJ6aCZ9RWx4F5m4EGi+U81X6hTy6Am
f+2CorLXd9KYVKI/GGQB7rHkP+t/Y3JFJGsVDwctOL5F1qaFLD4ydRhE5qTNlvpK298FiQ53lMk5
7Pn/49uSUQvTjxuYF14YoIegrq8hXQ+eI5y4HjBwCQ5Qacxuc4fwuvTlnT3pchu2tGDBQ5scGyZQ
P8lz/hTFp8EPwiA6sAm2d9I9fKwYJIBxc87NEhiJXtr5NV4zP28OQa31pXPx0LWw7UkJic9CVP+A
351ei8rkLymWrZQcXtA28TJgZp2bVslrPIC3Z3STd3d5cZPLK3FLe9GPUl1IlqwgKxvQI+tiEIdG
0KBmHAi79lThUW9+ew1mU1uJd+DTgE+QV+Dx3ENtd+fD8fv4/13iBJid0mHgQ43ZIXg0kHumr7Nk
PBAkvEvASDog2SZV4P+FFYH3FCXwQ0xYN3lsV4Eg9jQuGO+z++Y21gw9gejBKU1Yaq1dV2PyvM9u
s4tQImauJ0M0EHD991mMbZMmCkgPy4DMhBI/OY2guqWcFhmx7Qo9d2I6jnByN1SNGxUKn/Z94hZ0
VsCdKinm8mPdLPF7x3hpYn+AI9gEecKroHaOagjfaH+v0MFvMfQUa9Qq40BY7WsPpkiHFMyKLTqA
Tv+2o0+MSdqf6Otpg1wsC7S/zcxWsrunAnD8GkK+nFeQPxTftObthuKgJlfy3p50a93w9XDmKaWG
Lkb52lP2O4HlUhw7Pk6EoRTzcPgSwxQBafO75Ek5lbuPOhaKNqzZSjv1vM4jcfXEaCTmm+Nh2Ffa
sPv1DL9fVe2nY5VdtkNQxDWQ6D/6EbQRDtC1GZV2SyQ6pCcSIWAd9pLG8mT1S07E/hRoJyunz6Zh
YB93/Kaxo1sRr/RIZ8Ew+C3pomRgjqgbnK2mAc7b0qaURTMsUGIxCzPx6sH7145aER5S0bDViYZW
uzagIeEC4idJ9AhfewqMoQGveJbPcgT0LUexvby/b2s0mptwNfghc7D3YMire7YscGP66Fp9IKkz
s6T7QARLdtiNYGf+FJY/mCH72B4ieXy0vW8jgjp++uLQY0PCbXPgsaj7tESj1GFTmTUG2Fi+k69w
QXBsC6HDWQyzJdIN1KWlA0P34voUm+tsA3WVEXFyuZmbi1o5pVOHyeRMbTmjV1U2e5qzWfY8TqRd
ykhXvGq/iwEwV2xUI2IThj8RzkHQvpMXpJ6wiaLq8NjfOST2PeJGfjitQ/GrAdF23FmnbSDwFhPx
9rbOfxtt11mX1JQf731EapsIk8Kwz58dQJ2DYhYTJmtkukTrlwQtrvpXzJTA36EKBoND3y5PztmO
TZoZ2AqPW2UUa7qp76FqBqjLHzCL+rbLWrc4g/CmrHbj7yBUWNsLwNy4+xa+n8ll5CbzgkLCcteh
5n8Ixg5lBdkOOKYyjudPRqyGhvCkiv6Y7mDjcwKLRupjm9EdWCfrLCzWZyAK9+UJ0AmNkTWkixSa
2pzOWdJagGMd5cnIBretOe8YtsBUiQoXFXK4L5ljjWN+FdFIrRz27rUzBkuPEGMeYMzMIUBrExEY
VxXVKHiAZiQSgS78jmENsDr3EdgStU2RV92yH/W7OZedFlDK5+bLhNqZRFVZ6Gfyfbv0YBZsMZaP
xAj8/GS2Cx0PVpJv/KrFwLrGthmajSUvy0KUewZ3xeIp3Ozv+vvj0jK8OGvym9IYFENj818HVkxS
3nYb6nVQ2pFwl+8BTSftXBBZfaksgPfrXvLkVz5wwB3WkJw2WQQXUL3UuYjx3K2x1Zdfu3e1xlie
oRXS+QHTCvFl8UlKrPHGoxWxHBaSxaPfjVEjG20nGbElfI5WoqeRGqpwW+T53ZcqW4n+HujPXC/R
mFBt7qK+Nwv6R0hCv8/sxKcEiO0IwT0kTO6ytdiQrFdEsAL+WR8ynCFaQ5z1uDW4O/uzOos/eSTq
adPFS81T3PKRXDSfP8RLX8dIDwZJMJ1o2FUj9IOl80eFqxZLozOuC6ke8nsHpFG8w7I9l8016Xu9
mbEVQn5bZ7+ticg0y+AyostzuBcphntAtbmQPEWLAWq0BBUMf4lMdPM7O7+XilMpKlfFEyB6Vg5C
r+lFdYgmCwfZ80AAwpFCL+mmwcNHMzDxnyodmnW8BY3IJ1NTaZ8/QPj5zkM2SB7QJCPeThjXceHV
PoRdco7s1mN/tM+VdmsLxHsB290cQYzwBAXMirKJVzayibwJVC5CFpsMa41A2z4RCOhrhk6NqAVO
drIG1/+2yCzPW803UFNyg8mSzSBxY0Ie4BAqMrGn0KFZkzdjFA2cPu/KjXRyzAMAFUJ4p7uJ7f5O
1dWUBtxfuRFAwF2E7e6E+R+JcEfDMPJFPD3pmd6bF036BXyIueHMIMYvu4SdmNrpdHrDzSEQr38g
xGP1axLuhkd4aCLsDPNnSY8qPhTv/8NvAAxnaqKkQlEqJ+3EP0zC6f5RPDBsvVfi4wv/MadnyVwI
jkTZsAf6WNm7WEUl6MHo/21mpKuFXopi/memefKW1DrAgfQFDU1qOowuuyQ0jSGQmwvWjDfBFHNI
ApttjxlDbDdu3cDhYg6+3pD1E7l3z8sQTXQiRV/Wt4IhWK5P0m76sAKu823DAK+68awuzSU/VKJz
cPm9J9rgVr5are8uc00YRhk+W9RwLM1MToNQfUEN4K9nVouBpzyV4ugAwRkZHM0KzlVbL3vUc6/Q
K70AQZw1Y6lSoJ8/3u5PJCdwt1Ki1Li/TRGY9jgqIHliOhrzjmDKupOApjhgd6Znma4SFdOoXA8m
j9hs4+UhQ9mbVTv97I+N1QbkrsZXUQZaZzk/P6t5dERaS0pskU+cxhXAvkf7W0q0nb0qrLt0J4+1
0aBQkHjbEQU0YWZdS0CK9Vs2BkwWaHlxNq1EoewOmA6s1yV4edf7xT3seIKrf8pWvvT+RFIbMR1i
GU5HojCOM6UKDyx96h4F9s1yAxiWAR562D3KCisPibfPPds4harxRRFbVOge0WxKQtJcrptccAPv
6kGZMxzLiczra8QnicGo9z6gppxsSzJoquuWuD4l1LbirJbuBCdbt27vxBrj9tFP6XwFCWtPCH7g
1V4NWctCiOXypyrov4F8nQ1iF4D/GWxgI+LycDIKBZMkhw93OjRvd2qel5q6P5W+u09MyrgHLFlt
9WHmb0L+IKMdA3UU0VZN5829NxnMXgkEW8skm5nLLcwNtvJApG4vN1y+eha9/Mzf+4Ek7xXQYp4N
AoNCB9Hm4wxJT7X8KGdUzhvmCL29GyOuYo2f/3t4yHgGi8T9z9eAMWWVGIq+FXvEf9VqwsFMm9EA
smT4De5dZ/XMP7XW/w79cgc985ONwW3jxNL+Vt4+wS6etGIUc+g5/dhnZeh8ow0DutugJfUP/MUa
fAPd2I0yVz3YhAqJ5xjSfeOpPcZhfiRGqVA05v95yunX/ns5fzTxkr5R4XdRJC/kAe93NElHZXTG
wXQRgFLM+BXZ7Dm/i0N2n+kq07/0SHMCFtrF2/pc3TNpBawEAMvVWoKQNr52oQz1QszD1fZKPM6e
psNHUouHuSJkJdkFyWvvkmhavvVf/mh9pJNjNJqHofb8ljw6sWEP+ndAZYJ702FHGyNLCXKBPk0D
jZGQm8l1U6oecPt9BZKYqoXARYRgQ65AteudUelUWv2eLEFkU9plkmK5xyys5WMOEPrcmACue4Nn
PziIUW3iBjjFQcAHKhuZYhqKUYaRTrDPbTz1q8nop05azSIeq0awQvXoeGy5hf+rO03Y6YjoJK8y
1NdiLjwSxPIwMSQYf3EFLST6gMc+aNk1cP0weTUVvNS7YkYMu/x6aiArrObseEE/aig1+Fa2LExp
7wjG+PfpgrGx4pZWz1cBI5gHYuam41aYbswBDI0GghP0z87spPvJ8oTJGV3Bf5WqC7T9yEayG4TX
fwqkMkk2bGoUow8kfRosScHFEhYKptLbtH11pxnq2wLesRok2XHZhEiyNxOuiNY+rKjR7n5mLhi5
kCHM+kHB/sSQHBN75w6rDdDkXp7TeIia/g40jacucLcO1EjpA3Xta4JKtICWk/VoVUx3LuhVP/Lm
jh3C6/o/ZRt3cYSYLOyFV9f9QQfpl9dh52otzPeviBYUWWeOXQPRh0OA/3ogpEv22oy/JKnyv76H
f8FzXUa6ImK8Q9i7X/XcFHmtsrMCvB6ZcHGJX7lMj4cwDDWucmyJOAPcmfEaDQT5oi2aC0KXXUG3
Y02U4ti+NEcbF3kGwqP+nXuI2Nlz0ZcIZhGTWtX5EJ9ZpZkM+dO9gNfbwPm+z9Mw554AL0bCcz06
OLhl39HAmzXaX91/69gtpZeWFULS6i0PCbjMaQ1bUyICz5VjmKJ09fVp16jJfSnKMtzCk7W1Q5ty
k2qgsLjuaZFqeunsmLh8Udei5bt6XSihd7rX54l18ukxFpxXWm0609vKYHzbjjwqKpJ/By3GGn6W
Puy8whof8H64R+Flstf+OjjIHV7x2ipvXGFJegof9/yg3j01+73uVwRh1wXmzZu1o3xJc9yaE9l2
sUdLswcRqbeyskCxHxilak3gIX0qFfGdp941EJN8xdNBFMs8ug/DriOMDqbvzO0HdLSnW5ijwaE9
KhT8iuUrOEGGed7Yz4vsXpIfTGWYeCxOdxRMCYHdUStyazcST5g7gFutzAIlYZEldj/Lb5Z6AA4l
ogBF8LMg4mJ6C0yKEPZ4XEZfimn7+Js21P97C1JzsK9etvE3rIQpb9SFQxbhnVKJtYQpij7jGr7+
tjc312gBDO/kQLAo8Zz9ortjF0noqz5ONcuqHIdwvaZyZ9z6qusoD+KGmzjjaXea+4rcItWSx/Te
nqW/Y8XbRu7yEiRYQkqMue19HGSy1ZNR/ynqThfX3z3GB9gPJaBx9vWDc69/pXuwg/Ffk8hz9B0b
/fj7DnE+cY70mA+FJ4J3JmBRZ4Dc63h3UDplMpVrEHpeTy5Pj9nYOK4uFWHWkIwcNeXaQsnH5JEZ
kILyRUeAxSfMNnf/wq+GNqcQC4kRbdrhRMPvk9HqDRtxc+9A3c957e5WmcIg/trEUMbTO5BNbIo4
4vTxlae5HOsDuhHOv+39LQbq+XdwztxrezWsHC66Yhdr878Ofe94m4NAM+94P8GBFhjn+L9PzCy+
1LQxdIiO/qxk3+m3uykz1sJdKdox5By3JUefXgZyp1+Xc6u+A3AnsL9ZvMEmdOCSyydkHP3er/oi
UNdafyd+D0BnvsuOufOKgsmRWlV4rfile7IXbAaopJbxlnHvqs7bC9IxU4UdS9maq5PE1RReD0Ls
HcxDWJhUggBI5kMhMnJXvbyNRk8HQr3jANm2H+f7XyoJX2K7JGxzGhXAsG0+n9f8WaaIIVmxXwvt
3rRWtZ0Sxb4HrLFTEYta12zAhZJZVxwIUHwwbB6FuuYs0QYHcbPp5Up26Y2r0OuxGEobdNpm+y+F
sLCB6TbX0Nk7UeLSEjE2+MR8vkByjXdA/l1CLiZZ1xOZfSBrEz+dpdsjrVg+/5xumQpkiVogETzM
DBTIW1nkhvBDPW5DfM5NnWMSbraW3l6hqo0zeSP1g584fAufUtmdDrrNZvRcvQk70BBOqUV+TYm1
VSIBbbYOYJf9LgtfvpEdH1KdITnWtIsCWz30EiUvuC6lnHHU14N7GfJ15GFQ6IxHc3c17amd+hdd
HfnP1UkLwcw698pZ/JR063SevYFSoMhWfaY/KJXNEGU7tkTskCksuOCievxHkLDe8KMHbhRuhjHf
odXzrytXRrXbEPBK9nAD597IVKirpLLS6OkdGkCH9WnOjl/q2Pe8IQ3cHWjM7mJItWn/wsUP/NVP
Uyh44sDP/f73st6nt3tTpTdHTYD5lyN232jOuEWaCt0ApaDEtGiG9vKdH9CQGRRwTfG2+zehA1Og
aUqbyo961wPF0urSHF5ccM/REoJVYtHlHqu4ThVcb+61wcML/opyr9hsZi2xYH8QorP+Cf//Qj96
797KDor8SEUP/L0jxaqOrY5xPDGGnIJr3sodCDS2Zz2NwdD6A6foah6ymyD/pje+TS7wLvS8NnpI
c7PzurJ3s6T2shSsb/svPXXu0EH+sPFpjmzCRtc/cKEcKoQz0LdyhWDh2MZlbLGhUelddF2KzIy8
jZN+dXTLvipfCZ7bSdtfGn0dEhyzojazURhWX4D1PGBDyd3WRJbR3fsDlD5XpAoKn2w/5sruWtS0
VC7nmRr7qd1HKhO72v4QPIw7enkd+/3g8SOCT/6d6FS/hQa2h6NsvCv1p1wx/0eCk7n5kyrQXxfD
ndUnqo2qQqAx2bKXolXrMl4Uz3d7eK4SXdEuzwqRUSEXTxlKeiB6mSUis1BJEZkDG6kLvwvBOWJk
RQqED9lZogw0T9iiJb1MUWmypD24hI8A/KrHkI0bNdGPC4wuBXpr16XI55G0rGKJxNbhAKXB4k+g
j/2gbi/TNPIgx17mrObfp3DmAGETHU/jAaVc7RMRP1BbaIZeHbh/kA3bPS9AERb0e+5inbWLLIuz
7iS5ynHS9qSVcsPDm5tdxwhD2jFhSJkRMNxyPpxCZOKSFx3vEfrCtPkt6lnN0f64GDvidTn2Q/5J
ODXCE2WOn5wW4XdDNzjWEa7Sp1eTDbZSztazvmsjwQoBgVZ9qS7dN+vai9mvtfE2Tug0ffCHYzGT
R8BOyMrvk4fJ0/3keFUV/xNnx4RkLjukC2A12B23Gr1rILxuw+sfLraJRXyjsy3C8nFfMy6L5DnL
aM4UQlTTojCjbTeL72CdwWkzrcdImVHKbZIFPDuGmnkJE7fGa+MO7PLShk1ANvbeRzyYEn+fNWEo
noVf+wl4ScytBqO8heQN1aNk20+fZ9u1IhIg0+xv1q6D0udZBhlGMLuUplXV73+ZcnwSVA76JsiD
RKHPF8bs5m9hxDn5wOc1IYwD5JvuVGcLUd+MIsOfHNGcfz8stUIyV+jT3CycKAcMBhqT0vdEFmh3
RSYdPbGl5ASbJl19mdOT8xW0JrL3W+GIGF+vXoqdpndY1P0+VX85NZH2qg43p0ewWoJi4QR3TlTF
1Pv1er70qD7JPSzcL8IVnlkdaBMzmDSpQh73muGrsfHvqWGU94HYUxakS/ctbe6wKwTFTwg/XxrY
aiF37iA147OVNLoB4UEEg3IO3Kab483S7NHjOtkbU4kaVWHGtiZ2g6xOl67qeg3EPFiCkvDjcxl9
xEY0OLhvW2E/jCAcAIWTnZgR5p5owv9mlG7XJXhUJxbobsll+tfJkSU0yndup5/LZvlPoSFJmtn+
QkPfqx0hT5us38ZXWJfTf8i2dhn3T2AD79AHLYPv9/4S1c8O4qcQiVWh7jLwxWC7vLcEvC0w4ilx
Hr6SJWrjWcyvErG67DYUYQPpa02BEaPSc6XnGCbMtyo1SeTOUnB6bm+iZIhLwZZqv7MhKOuomVJO
wdsEa3WedFPBKJ+UBJ6OXlSLB3HV/xgK9S8dSkJVKenrHbLXMcTcOVHNPPW/fpD2uGBHILI7iV4W
ZXOEtNLXLCGq9cD+1fdbFjoxJ2FCbhyY+k4mzW87h3RtBVYbunoEC7Gb6/XeVhrCQc/6XnHa04M/
kI8C5/lmPgChN1N4rNXtOi0KnXYKCDI7FdtC9GMP3sQGuuUAjZCXTg+a7sXmGWbU/572bLN9b816
y7cw47VgHFL8fSj83kA4TRs/uJDIfHw+6uIZqKMKE3Yhn76w6HKNm50fIYXfG2isBpUevr0yUTG8
j1Gvkxli3j+6y+Wi0CfqK5iOM8ajzAVJdH5vRVcJglLCWt+XC0QcJUnIDf/JTY4LeJ5JdooShwQ2
MfUyXaWQTos+1EvE+oJ0p1+m0cZcf7swDvJ0BCL9JDYY/cLd6Ps6Bn3p//FcFyy2vqDv0lR3uy0A
1ZS+Q5hX+bA/vQ96htiWhaP50YJwsyfgcTsRmuSWyCUkArhONib4BsjNOzpxTiJnQ/v6TuXYSAUN
2jlivx7Kk7Z1cecq4AA+CSDCyHZa24cOTYQQxelT9AXXaDwm9nQ60CZJFYPixyKV9YVZPnfeO5Lh
0hcWUmc5CB7A3nDW22W2cqaUOOQccxc4DT4cRO/S1/RyyrNmrU4R372T9UI9EwvZB6qZsJl6bRtC
HReVPMFQEz4opaEtE8BjpNLrnW64po536P5JDrEz3lqPjVKbC1GkETwUHVTG4rUbEeN70BzR8i/b
69od9YMOo+6HwD7PU8nrwzuroOZyWJ9/CJLuSYJqjEDPQx+99kEybEhMK7MLd4Y4UqPaJqtLfXk8
u4AObVdpxXvTYn3w4UeQZX6a2U0g9+8x/4hhHoueZ0yjOfSAhHmoXsQPJoN83hqgb/P4evLcPu3T
C/Bh87vS8oxFZp9SQDjLQnoPXttjj45QfQBhX0jiVOr2rBOV7huJWAmM59hLLEEVW4ZFPoKNw3xr
nk73kAjsDSVH2v+JtO5Pk/feqyquZB2jHcUpwhZ9s7o1mpvXlpZE+RyiURLdDh+U0G/h5mxkeSNe
JAJwHl0HNZa1oKdp9H+7XCgj0PD3XwBxqBMkWeIgIW5lHwo+vUDJO1IQmFsspYRHWgSKOKVMp95R
tqeIoCOEFkxBPaSXpu4j0byGm8QP0QFQv2MX08x1oRRXrMMzFvf7HRHnvdHAxwEq9sNndvYOvVAO
rXsH9/fBdRDz8QcogmTCnZh6m4bpnNvV4tSEfjfAdwZSGTlQ+y9i73tJUd8FT0M7rbZNrBUYnAVn
JG3mhHAfQ3x7jdhooGsIaV7ue8Z51ON4oQm4TQA4mziGKMVlAN/jGlGfZmn9ibsuwl8Q8unaygz9
V0y1USx9gvg5Afd4KIhH+mBxNPut+7Tuzumw2KW/YUh+3MsoDSuLwJIM2wOE2IF8SzTGX/0BA95E
UcEFqcaaoMdck18i/Xd2SOcnt78cTFV32aST2dMERXyEl33PTFKwuty5SDZTAJxX2NluxHLX/M/L
L1HHoAp9Dbj7c3NYZigkKrPTQV1bMMOMP5nLSxyfltpKTXiBxIFbnu/aAf/JtSmATduyRBjSsdNE
rkCMSICLrAtEXNj007T/GTvVkZP8gP0Gt3M2wXS8+TpngnTrGFRSi7kl1D/BfWeKn9YfrxpPyENq
dtBiIm2KLWqvJEGlz4VXz8BCWCd6XPaWSZV6CawhtESXwGpe4+HRsizzXulEOOQm5f70C6KfzeCS
nsj8wgxzp6bATQ9Io/lJoY8gX5SWT4CB49nSrzmVr+/sRbwWLp01rGZ8CPVnmg1JwlwOK2Lp4jRp
xfNF3G+lEH+MBzu1T/BMAJR/FXeoi1ShiQ7SXiPzLifRkqpjmKUmRIe1njd6G+MopganwdW3ub1X
tJgnjTZuHkkeiAgke4fp03ZE5cPW/w1XR2/lIIPEK2J30N19BhWRPxkzSGnzFfgkdUiq5r1HMxtJ
avvTnpF8a3Co43xbSH08pl2RKiQ+2jFGiStnWVarPP2x4hUl8QVIyD22+ijRw2BNGifIXCXJrnp1
iUzaOsT0g1icXSvnjlzo3k4H2YpOc4b/u7gqTXuZPUtNN4tMp2dfy1r9vquAnjH15lqYFwelCWPb
4iGCIO5W0nnRJolBPKPeLgWlRpAsHGuOF5Ol/SxxtwQ7f54RKLDzckfpp5jLZw7Pq8Q8LJm0EIxl
eKv9qO1UFiomAQ8GSKK7MFyl9tstbqLDzLT6Gdqwo52WmMp9NXTnhxPl7yV3lEDFFIwZdZzSutP3
FgAcioo8sOrU4fr6vvej5W5qLy6mKxCHr3bSsssNdiVsWKKVPMNTB/gByzvnKIc6lgdE6s2RSEZ1
2eiwAFVzExn0cDPRvzQ4HJeCRO6Sd4QfMXkhSdBYmdei96AMLx+UZ64sU6UlGHy/q9fEZb0nsJz+
uT3qr/yzeZEaqI1w2/oqaG3hK5oSxVGwt4ev27slv9Kk8jMXP5BWQRjc2HK09wA6++0orZFb08Xw
xbFNZHtQUtI1tQDVAnDlljpKSt5Dn8Dew/EvaQ4vsqFia0o5CL7oCVEc2kbtEI/US8YSRQ5oDQBN
jsHKiViJLZifl7q4AWTPgAkmzjcd9z73lmA7ojp9IkA13BOcjhvxZiaLCLzdJCnED36ah9kDs1z7
4Ly1rj9u8Yi52kuqjACkpCOS/JRUPZpP5GtxQftHSGvfg/JqVJS1+x9zErwGQtTVasbxSpWeS7/d
s7ofhIs/GENHrAjwoOWElczwp1o42IZ2a2oDVpg2WNBEelb5G+wXjoLmColakNSLtqY3D9hc/q/7
r3yacanRC0iEKQS1s2XmyBVnFAx3pJW1A0GFF4AuxsinoyKDS3q+IU3Xl16W+9kfz0R46mgsdNVT
SK9QBQ8BgfyRc8xsLGrMpsp8acVI4K6a1IygueUS/GtnDgbB4bY/d8nfOzsiLGRNYcqMKwYpXz3d
g4jrbt6Jn3Hay9TJoPfhruUnFxkudlELzqgQDA1b8cB382SyW98rU0J4A9J1oqFBLXKRJoUId0sB
4p9gM9hL4EqkkTuGz5ssHxrWOw0sB7VTR8j5JhZQQGSk4h9BKQaguLN6vzigv1PDufY+1z2yL3WG
6jfJ/P3dIZEXH90ORwX9SJe2gcaD+DLg8aPSQRAt/d4hDfCWO/qTUwlmsXlMoXaSzEN2bEkFiOBI
ZZ8Kfj1z9qxfz1ZtP3weDCG/phBDuHq1uqMzt4rk7OhAxicdqoqRarHkaVs/eywJmLFCFkvWVfND
t1Tal6jOSksunmo+uhBFstcfIswbsC6SnDs2fodMBC8zOTTx2zHn1CNG+mhakiVO0/WUrPKeEJ5v
nHsw4fx0SNNTa+JHiTidl1Tcb8dztknCG+fTCEjosdZ80S9RMjw345XRPoXXCV4cz8M/ay5hSLVO
8Aq8evOF+7MRSwkk7wIh6tDsMlUE0506dfu+KtcGL8y99YOl0IZFx5NYZtfnk6aVk2JglJvPrttM
K+aXg2KfhanR1+FH+X3XzkVAPJ/OngtLr5c3pJmyHlmakyS9QP5l3iqlopo2goeUDgqJsWpqmQei
KLCj7sow/PYFpmRoi+sRBDcEJNMXzrRtZ0Q+2fjm2koeWUWktsYyWUyKGIyM/7B3NdXqygBZmI76
rezbaayy0ULG/qjbTeIP/6w/nAEYaSOuT/wKTQxeytvTA4AfigRBNMLGy8/jGInNzMIYbOoVLna7
gJpa4VQuTPTNYfgwWdePRlDWXb/yWYLoVguselPj0Irnt9jJWxMJWHsvnYpvHjQFKhdcyfvl6vvU
B3jypnXSqwj+ocZlDyRTt6G4Y/+5ikaZW6wl+24SLKXzhn68bOsmEJiXV2jhNaCv0DpbLpLTD7MI
IjWwpQA8OhaNL463vHGw84E38Ef+dZzaXVq3EFC5CuPrAxRq9ZyEo9/cBoV3DRR95tpDqhl6F0cq
yjLV9hySeDAARxIV6hWw6kNIF0uvTK1wEaEL+xLuR+lxeoWZH6mXJc+iHyPDsz/n0qUwhNUJMO6c
CXALahIEgCEs8O1jiRg6RBUsUJMfC7bNUdgW09xI8gUlu6S4d4hXLl7TDB2NkAmd7dXtfH1nT4At
c7vy3lqBun869TPM5xmjcx596zLz8FgANPkxUwKt1Q1toALWh9E9maaxpVhjCqS0Rx7Gr256JKoy
0TvjaHhMyF8Z4DfiRJg2Wb3bYwXTGASJFyKYu6G8Ig5wuk4+r1TEvFaFaOmrfBsk0scpkr1qGn3T
FnXJapbK7COQN555TbPC3N6JydV9cXk9mUqvApWYSyNMpxk4jCCcW9glTcd0KmUSLJWa1t5t26uo
+O6Sp7NjCODifOzBCD6AxmriUkyaa4/sbnP9GeAM8ZGAFne2OIKFukfsA/TyftuT71/WqCfhUGeS
/8HhfR+dwzvXFKNz1PxL4NQZJYhrSIvbAMclczFxWgDEAQpcNlifzRdtLlPhDPClBc2Bc76Dhee6
jGIVgrnC2uOGq4ahl25khMOUWaFKkkrSXGUTq/WBIKN3NDTmuE7gXmfOXrNgkTeMZWazoTbmW4/0
Q7Z/qsR4XioQ5fIT2vPDsH/ArGFISTXhZQZ/KcAai9FCsH34bHhB+etOrc9IfM2apYDsFdvf04tN
z7H5xKZkPLr2YQJ04lzfrglFwGtddP1+PJTExi3Xu+bFOeypKgZnPh47/greEgGbK/GXdlKNnaDn
XPZCKYx0+5gVHp2vd0DBGYThnB1LBCfCFHEG72cRHJHWPKOafT3w5vrhZehbEYKTi19xjAlcf5ca
1eJwY70nJwUhoQ+n3TFL2drq6bTDlmJl9qsyORuqk5A1As2nvCB4zlaqHwAdXhFGFk5wSyGdTs44
PPpYpC5MnU/kV20pnM6Svc6NxPxDBktzp+g6JJ9G3jN5tK1hMHMGNPqUH3z7diBrat5/fY4ZWVaK
Fqg3MwsqPi2PUkRbe+6alDTsq+M7yQUdJsTKVn1EcLto0E/ZVpXg7Fvz14donhizZYje6CX/flHA
l8DwXhadLn/4j5llCYw0ywaYMU8KoXSTKAaQHLI2R8ctsQygiJHc+8R2rhChinD4OqxveUMrk/2O
x9Bl2aOqd07BHVJEciG518s6Z2CObjBGLx5b/sNfsnAIt67+TCRBt+IkxunUPm2KQesXmhjcnKPg
avPPvtdA7PY07u6sjnPZCVuDaVgo1d6KD3xRQj+2vaLWSlFW7e4FaYvoDc+haqqfan/xd3YgIOBX
/f0nCofK+PyHbPo7JjJhpVAE4bu6OH2x+r0snHzIazXyGX7AiH72ixsMGFTQ/auQE1C9V60QWEkh
YMVGKzNVPYOJOw85Jjb6HfyLCvRSUduPS8G+cF2LzT4/q36IRciZXVsyW3a7ARjcJ+F14F6HArnn
CfKKSel4H/J3oUXiFLObic1Qhl3a7wlJ+0R6l0NtSuaCtrLDDd5IWkiGijf2bbdMQ0AsovRknCkA
Y7Ul6bisLI32htaYKMVwK713ur/yTrnbVNoG/iRKHlEjoSEfPyVzJzQ5y0sbnvqIDuo+OjNZOEHy
dDeqa9BLARUOxaezqowem6QLq1uDIGjQYMLo2hwbDGyRFNKn4cY7H03v9H2r+Lfj2UOQ4udrZ93b
o+R15y1NIIMwBO9dDLxQCzBssnen1hqCwPYTW/lZYlv7DUCxTgdmKBWzCGFHdlYZBKjAQP83ZPbi
BXK0vGCf4PL65GtNqWXCGoQVnollAZgRnNUIx/izMewx0DV+WcW7zU2R86olmn/toYzF/S9xNGyQ
XX/WcrcnwRqkd6rKtSbaFKtHD4PJ1bAzNcUhU4EKcFG6nLeNzk+cDkRgzePN2YqwpzNzHyI4RL/N
q6Ig6mTIaN7kIPlFa+BlHRHzyY8YTeRmuJVGSLZZkPCgXjGcIqRlZtcdUDTB47pTl5a/lfEoC9AX
RGVfHA+gtZV2LBx4IZfmdJxGjhq/N/Q1CuN+pf9Ecxdn6H6w7fUAQe9EzIMPKY5voD+VBb8SI8da
rtp+gzIca6e/SFf9uqjgL6bClGVrYW6lKahoiJ//oqOh/WDylu/aC8kB+aGL75eImVbNEVjQJ7SP
wDT+aGX5l/L5YgX8sWwFHEwifkEqsF8Ro2TnLMWBY8Hh998tA8nWXgDEUXzXOYBQBWCSlzY6Hzac
6kH+6JWDd2kSgvhGojKNEQPrclJp28Ah4h0KbHzJlvKDhNtuCoWO+HqHvSXGwKm2R29pRB7Rv3gF
DWmDFV/OJycf+EmxC4DI2bQKAwTwu1DaOwPTPspYzogg1KdxVQ3/uc0Ap6DoG4fkrt4MYlFaKjRf
qQMIE9ptF+5XghsmiE75lqwmc7MdJB60elJGN03DyLjaNyj9vW2b74SY4WzN085o0nBnxCc0hioa
gmRikSAy3UjXP9OoUUVO8HdF1/g3PhoMw49QCfzqe7eVdwaRRTeM4Bf3YybSwAO+rrX6/iHjzd14
yOT5v8kDjZXKRf6QGR/E33N4Y/7H9EbrdxbYWL7D+B+1U3jlUtNKo3ldN/BHzqA4jgakzbG2nJQf
lksSxCi8PblWWYLCIYqBBKNivu2aohX4FYZOzd1U/frElSK60zR0+r3behT6T8sPB8PKEELkS7GO
G6rbwqTgySg9/ksYJgVT2K3TJDeHbiDAMUJjnEsJqm7edK1fI58acoKPo6tj8cL+N/947YMJo/r4
9HSF8Hj4pdiW6ewHojYaxv1ni3dkr2b2Yh9p8MqsU3VUs1EyezB+MMfJ0xRz91g2dQolFYF0c5FY
JQihES4rjFAOSIvaRdKf9NYb7Y3JH/0xjtjXgboVHtRfGEaWemnDWP4fFXlumLUmKt925nBTl5nG
paqrWBT2DVCsoofr391WYYvX4p1CYx6mVxPwt8sqWZP1lvh6p42hFeXy+/coYVmNUXn0eF+6N7eI
W2N5P8xIdvaObJC7m2TmJUi4BRR7Z4KXNht+4/HFXrKspLwl4FGajF+IitkKjTC4rcCPvOInjYta
d7S+UcaXJmjX3zVDWyr4rdFmA+o8uiv+umEoOb11wKaohkCe7RHZnJ0PF3vZDRmpEvUU5YSekH2X
GWfQ1OdYcJvjBlf8ExcT1B0EYo+nCytBwyGTM/g3ArZ2ggnCJm3x1nIysr3a5fWq3xcgFoJ47e7b
w/uioOM+UIft80VnnfdBuWEZ7aSqjSUjuoI6a8o5XMl7DE1D7J8WPxhSwAtWMNYxJTX1BsfT3rGT
/1CfgJTjB0Rv3rcUEuyEgLUhMzEP85Jf53HwHiP2Dkis/wVh4ToSz6kIFHLzgQW0pS7hRJmWSWwb
5iK48dF4b0XOpKkY286V/0lFhCVhVig/xjGA97kTHVYIMrM6NBJoKX4vJbCmfSVnsZzpEJxGAgmQ
/4C7SYW+2niJ7tzCrEHIDmt7Es1ERnwMQfi5wY1pcxPALofp6FVZzT9FYJXjsnFPsqyxAZHzMH6y
+h0duCtKLhPvfihw3LVuVxvg5U/IiCJouLvd+91/nXPok/tiudaRd/HjNL+J5FLXAtcjE6r0MjNW
Kn4a8S0tfjVPzY+LTU/ampeYYj+O4lr6OEo53Sc6lCh0ADuuVFt8+oQp2R8CFyOM511pkPrtszIR
Aj2Gm1rQTVVgk78bNEYlWkswcaWi1yA02XmMlyUK6U8TDFYTKbRVNghmq7lElOg5MtMfFJexsi4k
7jXtQbt/D4667Cprw9q2gnWLGAZaJHtdFPPuoOYLLCm+6F3VpBJ/0upCrPguPbr3zwxC62ydmB42
R88H+rslmzfqs+vikL/KYBASYCYJq1cYxCjTUYiWh4su3zpE3/X4EDfoxSWUJ6C0jhibTvn+HlZ4
eG2zHYYfVIm6BluTczzQfaquEruKqYqFJg7DbUc6siPqQ+mJxETRf2iFetNqv1wJZCSSnCo5SQgr
uKcD8j+fiqFcOKPg8gf71ZCNYlx/49QMVA1Qaj/N6A9qMwW6GPept48NCcee+hJp3WjTlTDZFNQ3
8w6AnDhJnXnRs3q7lC00NBWuXSuyjd0urUFy3MiIzrr2TGFnAxqqClmbTEoe/0fWfJ8B6F/E+LV2
1q2tW4DFWhbP6MMMWC1xFjff0mpRn1o5fB79obnkGadWpmZdPlJISfVV5q+a2oeLOzVw2WE1fYq1
FdtTlMzcDXZyonfUK8X5WfMm9KILbSAN7A3UuH1EloE6uhBFpsqsqHVmD4eesCaDi97zzqyrdqtn
aYSNCDEc2mFq2+krlAGobQUTh2QZCqR7vLfMX0nP9ETu/OdfpXRK1ruh2jeZpEOtJ/bDU3b09ri9
NU5tC45WmW3lriA07xdK6QP6vf7vozLhjHZ7PRtORDtzRYKqfzkd+eIosQ+x3R5w+OCNpbVLIIn3
lyFaXnsdxJBzhMgqzsjcbSnVYdLrkbzNv5c3mKRWUoONGWxV41WRByOe0dvWwbWWVxZnlPlbN6R9
lDqzyvrEOdybHZW6SSEpr+vZWUxG0wta1moaDlSNaItmpV1N4hkOUYEC6dWp7GtI7EFkX8HWz5D7
iCHRXSp0PbqZcHALI1I4izTW25H5GePKzOuCOvw5VUFGVB9114B63ROe1C4wXoHllw8o+/rv5SoU
p00SOCALBZxiFbZjUuoqa1fze66goz+EpJgLmI2603nrCe/RDZPDQc0QBkidajpL0NkR3t5ON2Pz
BM1rseRdFSA6hiCmiRU+Mm1txlconZwPYd5S/W5gCPIwmvfbKS+FbP55J6D5+a/Rw/bG8/5qU3ne
9U723Ik9ym5KwdiS/dvMgvLBAYxgJNJzHOHkg5Oveu9Jk0KSwwTUBLxxJnGI8esBDir0ywiiO+yt
5xs6i4Y3XJzhTCFpjh4HHh3t98ztKtCZMua2/elk01kS24SG6rqL/bzf9BK17jRCq2+YQMliUtPk
Uxki0sqtRg0qqIhOwQvZjjvo9UfTIqTQPF7v7kuBc63NYsrvwvpvfw+48MZpUcV/HnS1pK4Fp8Gz
WRoJ301T4cuNExNYWnRUQ763RuTsY5FEkoc9vH2UKo0UGxPy1zaG2LmcdyxDOdIJOwbESNwnW8E0
m9V6d1DJW/p9dEz8TwbnkvmuRmlq+Tt2Broa50UhDLxIBKLJwqRkYd4RCz4OyeSg1EYnXGQr1Xan
kVQ0uNK7HBpZQuCqIqNASSextdoC0tp/HPamNGG4EVuf6qO1XHy5iLUEvH+8rMTKbH/9IqN2wieO
vzNu4qERphVJMthYqJL6unhMvZp2AyZGcDKu9KRtLNLLsXsgtmDK2JgeqvWIcxgkPlmsBxBY/pUF
5NvDkXKnSi64k3HWaoEyVN6ptPwqm/sCefda+KgJ3UgesbY4uiat+5w61f8drIUHIKkwtH/1XyjY
SnuHJWJcefZq+WwmmGkw5wCp9RSzA100T7BR1W6n4VsCTOZmBCP9eaOiLAqrPOaBxxFT4Y1Xp91R
EuyK2JMhO764CFBCDlyCSmAMXCnsQg8VCPz6i7vsMz3KlNWQpewiJYGvjWhFVeif23tnHXBeK7eu
j7zFhQ1tvDQh9D5eWpRXlOFPMT36WtMr+qN2GRuErma1ZI8Z3PjscKvneuvo89uUn7wBbNkzLxqO
Ih+unWGAsRUjio66lnnBxjy3u2hlI5EimztYhg4jc1p19mpaN5GocOWttFdnuHlD40CLond8zKOM
MEpabfSDsg0lMv4ly2Ybt4WrxklP8LaStPhclFohCkUR8zUnmCDjDD3YlPKbN/gbIuwrMzvHv0JJ
1yDPXbEEDUBiI156Y5Fm0pgo5n/9S1EGBMrly3cw+y4/geD9a2e0ldrYdRRWdv6iRSw0Ipmn2a0x
7WbvLNkvYCkuBCriMrZ+aEZb+E+r9rKaYiIznOTXTt/DGGHRDVp6ofmo3dZOfLYbfgfynTE6eRUK
9bG4rJZ94e+AtFnk3kBvzWzJnQAVXiug14dYxvNDgOr3JwPRznEDDCXNF2mXdFkRwuNSy8knIl5Z
Prh4rV4k2KLRlQMb3r5lQDewZvIIxFGxc/QBEkGdPwN4npSpbDmSmU/pa8I7iSdKHbTD7gFiv0m/
PrQQzmTJE+gZY0LPZP9wHDWv7yc/wJ+jtPBQvIjJjoMqtUPnJbYlQJucrhylBWKDttN+Dxb9POkr
yrGpOiFrHhvrpdBay7FXaEJ9PQYqghNZYJyhW+oQexUzoOIJMar23L+kp6ONnLY9QXim3K7wHXmS
CZH5ohscRc7lYlNaSYhFvLWMrgoctky4qFKK6G4zsdR+nXVZIIrDpR1hfpIfJMGPbK+ICITKeiSi
A/JzumHgiRl/p4W9Hwa26lvnAGN8DYfVydd28tB291yZkpcBscm2zwX7U2AtOEdwPq6HURMh8sB0
nPaiaOk0MSER2ceq4hx0RU9yDJXBACxC84fS1gN1JC2IBiC7W3SCLslBdZxY7fcNOdheBA6SucAF
Hr3CbehCvEC0eTWYEQkxcp6cu+n+8ZbCRLT94Ud9QCpj1j+XY3fBbs4tCd7ZTQ+1kJhpUq8zpMf+
4EswqN0nku3rxXQZvHvH+wqYjFoTI3L7cGFko57OjfGuSICQSY+k/0hnVcoHWox3SpX6OeLvTiag
LPRRU4G6ySx4NipOCyqyYrNbrDf3yHp1f4qFN7i3+rnO1/ximoOlM+QgdUYgwQMy+2DOd+mT3Ih0
4pZCeCZ3iFV8v0bhbB6tcJWeWVmbvpJgf+W2CXMmmwUNYDyY6UmT8o6cpW+9tNPfkEnRX99gnM+p
5PoW2OswvfhkoYzad4U/aVghimF6Gz0KHlj6HQRPLJkpVFqbufqPjbJCSP3Kz2gmZSgiF6EJ1YEP
nLeJZtYa2/u14+oT1za5u8lKNewvfsuNh7+hcXBcm9pai4WRongpxbs1FuewyiCNEOhoO6HJZHcn
XXezBFiN6fpgOZmoznt/Iu/vxm8v+5OBA97YbkpIASGl/Gy446jM8kzqJ+wmKZCvYK1HorCwOzfd
jflYNIj13uIabjFI/ZrPdVHq9x94qq/2tMosmnl6z/DbghM2E1HEMjc3vpLK9EPc6XCyfil+/FpM
m4mEI6GWFGCsIsndEyThUlAIRsxRjbLrta41bITUK7dMb7LUR8DrUisiVYVbHmYD7rfEaAqPBuIS
wggRP/5vCA0fbbkw7v28bRMQrusgi/gGUCH1nCmgKGUB9HE9Heb6OlhsSytq+Tvl0+4LibaYQXFQ
oZIoeXvA7II17ki/iaHUveOLYKo8vP7ux85BUMCJU01HfGOy6sL7ZhSKqjH2DP7ejsCZY4Tb68lz
bzyfkPAWuL3NfNXVPo2FZWfm3XDdcrqnhThLRN9Q47968jmo/q8/FU3Lwl4QLcmT+ilP2Dj4GGom
rQ+i63xXUQVvPAGHiZXYO5rMjOI/fsMA7mE4qQgvOZmGB6D4W7bDYzp+MeSWboJhM9VxVpk9C3CS
ccQw4AMdPXZ0wPUuqaBP1afa43KJZ1Xxev5UOdGd9oAyWY2J+/TFJY1qd//TxoTtuGs5VkGQS3Pw
xFVSpYVWWV7pZLIFpvuipuFWPPiKOYtxhUVEPN0XjErhcQF5QCCfA4ibO7AzJr9bJWuyimjskphY
W/Jm2skXGQyQMgAoQi1jmW68GlYUeUrvExc8qSeBJH98yyNhp2qx6ExmoxPVg2YvGn53uPymRdck
igX7CAjHWK7vzOaJn0wxl7+X59Jb/9546z3Z8LRPamHqnn/jyJ2jCYJn0w0S+TJxRfwo7Y/u0x7v
LAJZ5B1PH7QJs9/AqQQzLiHZqkQ46QRHHxdSQj4bT1ouZa7JLT2rrms+rHoR0OCxxBc7OBBw8gL2
ds16ClTsF/GIIR8GMpInhyv1aLuJ9/uQgLJEQ9cRrxcEtrKsXQKItUdJEf/ISdDDTKK2vUG6wEYa
wve/AhzdqiG2HlUSqIitTEXcuXKqg7Fm0iX6NMbo0z8Ij1FbxHZ5/53HPS7/fFaFTYQWgKKWSWTL
Jo0U/2BxDjxDfo60sJAxMc2zwgAA59pAAUFkwj2HjfF+ewxhSy0N2NuGuTcD78otOjIMAe8mtEba
RRGnZtYB9UsIpFUHOOESK3ljWDC1Tg2RGugK2iugK/nbAvCCmaYslGzUdx8K70qBlllTxcuOWwIN
kNh559BgUjS8i/+82mhD3pIO95APEJ8wxTRc7raxDFrQoWKRgHvABl9dgBgQ/gs3fseXFxrOJgpR
HiNv0ELb0Iz13jmYQ5u/80w0p9QjYhAbx1JH3wpLP2ZwAQkl9DBNqbdznx2lunnllTx3+WoRs1+4
ULU3gwyCQqKbSzTtuHYZNuGGFm9uhV87olh0t4QBJQlg4ncu0vwnLGEQkBmdG/naS+tAi1RTQXnY
+f8wJ+uV8cVEBwsYsvZXPuMeWI0s0GwzPKo7oAaFJR/F+192t6KAwLuYOF9Vy+ibLn1eKQpARE/e
IyNizFlhC9+hb9bPysebX/zqPnf/AhHzPexYJ0pSGMGW8Acy24+dvqWzj0CgpCqKlfIF2XmLuLBt
11T+PuqLppM7mVVXgoLbqJ+diZ4ZKKFntAGlU3pOyK5OLHLlKHMwBpMYAImTVLAFkGUdtib4GVov
K/+cmMUidZZe5xPbF+uj/UMEC61vMeM4/X6r366ukxxYBqA68Pm/0nSirE23RGo8tNC1qn/+lzgq
fsM1Rt3ivGkVV4iJKa+tynDjB8499XxC113ldWWVSouFFNs52d7Px0WvcYiw871qFCKiHzN0kI70
Dcm/oLvSZfmwlgYWaTtpSPYDRIopjy09KUk77L3P2/z4Ph1/nD3ORhtGU30k34aha7/Fd29Szzu5
wgN62CLayV/Bea9OE6a7RTVi2zRDkUIPZjgWqhyxJ19rUktjybGFmn8XI54Sgl+a5poRIWtVYi6i
xzPMd1hzofM2h842ueKDkYKfSm1bHVr5SqL1oGbtOBf4uFnkd+EFun+O4hS7O4HWycjwSYpFTg22
aiR91hwQg9XH/BSyJEJtKhiW5zg902HlfJl9UfPFLxYUOGo6OzE1nOMEQVqathtNbsw5t+LerJ3h
8oMsxNI0QwxnZxQBmZxl3TWwWiZpFN1KFbM81g5YK6ahHv1jjG4KhL0tQwzvIk2g1Z5cdnJlH+yO
SO/oj8obfvaEZ5hg7QqlhjwU/zG5LMeY+qW9O/TllVE2S1oeb+od0fNrpAMXAwl5dd8PLWtiPD0b
DNVnLSxJACDQFiRpcR25lUZ2C+N4smmOyBw6Ooym0W9muYnb26cObf0rBjFSmFfIJzF9rBErMNYQ
aOezJIR8w4Vto/K75qpTEstidkuzxJvkFspua4nheEXfUO79WYxd0oXraQHiTm5VxLygmNFZnlPm
/Qv1NuVar69f6rOd2Gw1T92DHvODUzhfca8OJGT4ZuPGkI/b2ZHZVbC4hhgadnshm67Vl2Ov6Fix
xBCC+WLHV9Yrp98LmsGoLgyBh1fpIdgNJ8fDvk2S8u0+pYUlaChfMAaS9o1hjB7NrxX42Yp02h8I
Cfx1ogHbna2ka6aPtV9Op0fBASK39M/cWFve4GqRCkAZami8AOJ0MZfSbkhPkCtJz6kTjSzWoIQX
EJIXApQAm4BcJgIVFFSL0z57Lylp+mNwLn9i+2NL4HNCQpG6OCRtdxkZLYWSK+khcAOcbYgJm4IN
V+PNQ3XdfA9nj7LmN1FldJVQ+lBR9iPVB76Na7yu+nJyuqpEdbBkD/CegfZSwHrVCe0Ej84UBYgq
Svvnu0pN48CndMpozIlP1NSaAeb/2Fti+bo7XpKR8Sjqo/OS5rU8dA/AMqF4SqPVHFjw1BIl5SKx
XR8JHe5gPECowcqFbd0N7ucTfDUo2QoMj/qLoFYvaYTsyT9w8m/Z4CHFb/AW1DrnJ+XGtCvWk0op
cuWj/BV3yDQcmz76UhKyVsCdkiCfIHEv1LDQ9irb3YP2UL7JRe6XD3UT/k/mHD9B2EZOCCKr4gQ1
SAE6FAR6WAGDY6iTpel8qn1592irTRKlh/Dm7tp/iocLAFEqJDZC4mJSe/CX0LbikqogLsQ50wu6
SDPyMTZ6RYNpuItxoItx5bliI+Sl1OhJyFoqYOpcLrdFk5WbligNI2S4RYw04SkbVvYB1TcFtRkL
qO0DbrFoYEubJrI6e6yBzaBDxMzVp+d5iiy8KxeNkfG8NvavmFFD72wtJn7bZwKgNQr+R+nH+E9Y
KUpViLL4gr1W8g0bf/MlL8C8dXImuzikolVB/mrDRCQhGx+Fj+geI3MYADa2icp/UL/KZ0OzKC0q
SPGNIXq4VjZrHAHR0suAl7G98GY1lIp/bp1zGjjCYVcy0CYCJqmep3H1tXKIR0E1SihSNFf+T0Ql
5Iv2seYbjjA+0SAto96QhjElvXEB9fvlfLvblSVqQ2l0uZ2F4hIdZo90UOJ1Wj2Hw6c0PQ1aDOpV
46vKD7aRZoDBAC2BhKC3pxrVGciTRRYlf2CHNCRxQrHp+PJ+BYvoI93P1s2hJzuo22ldPAxxwJ/9
wOrdfaafyDQKG/Z6sgINFuEF3TgaUd0jvJVY08DBzgbrGw/R4eIeM1wDP9hIw2IgNISV9mlTaQun
CD8wS7AWb8XkF/8WRWqn4FRz54JpC8mfXccSRKOPlUkTCL4FLH0Ff8Gx6+mfHFvzQccg0bPW5RuZ
mgh/GlLHqrchVfeR0rB0zAdoJj1uAHOfT5ZU8NZVNwWs4P9C0JPR5ayUkCeuqsVtdGrWtwV/2lyp
GINQSz6rW1K55VTWQ8O5mH7waqd2Jh8KU0VXz0iQNAzcsrYE7KE5MJVKevYi6Eg6+supB0RlVROt
OmmI7cr4Ju2NXMHwnyIb4iS57Vgr63KIqNPeJjwOEXVvc6J7nfZqyPybYeKAH44G/z7OeYahUvhv
/d5S4ni8iNx9bKNKpCv/CYyBLti/JSwB/+8TGCf+9gq5ntK6VdOZx/HkbgQOOZd2WDG34UsCwlLc
xCHM7Zr1Ynzh6WVOIW3FQsPPue6rmVIs7zLRVH2k++n78ljTmlVqg7bEjYlbmdyC5DRMGRX6Pn0X
QEX+T+nJXG3KKDwcrn+Zb5brVPLOi2GwZ6UleJe5BvsUM4tjloFIBGa1nAOvlWyPEv1oBsv6KOS6
Cp755kHsNCyCizGVQOPRWWTSlKcFiejklRuGKPdsWXdY+MpbcUIUHGDtCz4CS91NJ0pThT0vBMij
LwbDOb79cp9s7NgH9o+ZmC9CEwDaOGzTTcTjlP+0mKRHota+6o9lo97zhdQUMTn2ZjOyKX9b6C3o
aVJeYE6+ldOB/pFcg5XlTH0TjUvMgJvGRR95vypNsYfpHsUY+un+1CH0z/bnWNRYdF6DfbMvTRGi
l/gqZv0bvjvM6XmoOa4gTM+uh8YMg2oVEaOXDFs12AGg8GEmABeeggvKi8GKoxRrNXGWvKWgpv/4
8x11skI+GicwHBEK3qcMoLnHiW+ykdmmgTCos/37BBIZswM+wBDMamDXCdzULnPGgeTPEBXCrocb
7k+6XcZKgI35p9+vmEN+kP0/b+roPd90RAfEodYIWwHEUweqtdmmuMleo9bND61f0j+hsCQXBDWH
/oOOh2AysXhYXkjEvGTKUFk2vfX5+ov+fIE1LNckqHHUeLcpvpX0ltBs3ka0dFBT7R+5xAhaQFxM
qh3d4NsTDsT6+2Lmg9REAOntmQvtwiN7Ha78+gigm0CZap3ZW/AwuJN3Xd/3uzPLEk8XZLh3K1os
JwoTnBMGg4XzzW1j7am87nlkV7tQmV1rG711M9pK238AYU5oQfRWydbl5ajdf4cS7HcC8253Ia0C
NGbyh61kh5g8ZleQkRjN0U/ZL9HAhMX1q4GsotYeg36DjdGcrpbhJlalrQ5b9KsNz7QmUT1NiJyi
bZJ20cvPCyULEzIumArl24qCMjTcmg1C8Vgk9FUYsUgaVd3ipdiYnVgKpORe+uuwYIsNaOiSboeJ
ikFjD6b3+Tt9rz8yjPSWYBC4KqfHNsjnsUCuqXJ6OKvr8JitgNxtbShK36672GhEb41QrE4aJcwq
TYwJTS7+HB6F9NEbSTqrzhz4iMM+2W3TJRGjJaiZ+xy0SokUP5LPcHln0K7Hm5tkqP3iO49PHmnd
AhsXaF75go+SEryFu6TlD6AxFw+PzPRaHeQV49fx+mPa6vKDXI1eGyZdx9GY3DZyq+dpX5tCRAlS
/oUYsiWspG5NYhz6M1i1MrAYxiIlrsHkqWl4aCfrr26bBtpd2Xx3hhpCZ5WcySF04GmEwN6xERZb
36dySGs35dvP0USH3Wx0oaSC1WbdAO9/BEcmIFbucTk1CxthYL2FU5XiKu0iyyqmQ0V40FKEHgp0
5dxi5cSOWV/VXMebpRqQ3clmLsDD0ddcb4fD1T3ooEqICRmdB66SfaXMhNOY349JKzZheJfMbKK6
OPG96X3x+kQ02syOIvNWEn3ir6HgQLuS1aKb7MgHRhkNDhWvR9WXB4wmXOvjyCs65Ivnl1e6zGwo
yi15w9weBhAtigrCyi8frqw73VARSF63ubNNTvi7gbqvRYG4Whdjz6pW5IDl/1JStAGvUqkljGTw
9CgMvuOOKSIrX/XyMeObe/5aaq6vIoYNuRv6yZgSUpA03Foa/P4AGU0TEzC23MZKMH+EM9SDdGEC
LMWcZYOeIwFoonF/fnFP9UGA4UoLEolou9BtXyUYKTP9jmUCHeqMYNDduzrxJHYKSurCtXiFVcFJ
MzEVBlOR73X6h1QuhnB2opuWntOPObMlg9ZGFGhB4+83ySyVzp1Hu7lb2/HZP2o+sEZAzhX1HP/D
8CM7GFDvY87fMEsRHlIibHYeXD4vA0+Qq5uM4WnMpdUe6oI8/RND/xk2dGudR2GHgh1qGM17YN0I
vbYI3BX06X7wlyC79ixfy03MdSIb0pySCDAoWiCY0U3Io16NTWBYJAEyO5xtrvCbWD7AoJVmXJCO
hotBVR2wX+emsK6Muo++B6BWyVcBslPVaDxHox3M3BK/iPhT5KzDOI2Y1ZNxvE4tgwon7qj5zENO
9glXO5vuZkIbvtR1kJ8hez/b5xnJayoYHI4wgO4wzyK9G21EVD1WQX6pFVwB4LfFyghxtNrdhtit
ocv81KjLgUquLHia/h0VfFXFVbFMoqSNk2mOnqe7CkMu0o6xmJA1SwJs1bRsYityGvMRy1k1NY9J
fHQe7HSb6W/fk6+XliY+sMbkaNqpTWbB7CQKu0SFMKW6yo7HxSd5lUvtoT0Zw1FTwB8QNaGEjnsF
F/3zpAezo7TKp9gKg/qwddtBZ9lthk7AksyxdvIqQS5UKkJ3cB9BmeKtrGMDRn6WLGUopXmA9235
b6xPwh10StBZZh8vm5L/YwuerQheT1gxl9CzxGub40hD6nAUHD6v0Hd5E2nC4p2i9JIyosOtMmLB
GUmDoeTSnQDM+iIMMslGSzFO1+FARQ4ct85oGBmlvFjKp5x2IJzn+Ig4u8Ouo54C1VpgKyOTF0ut
BRSMt+5Xik33b0eswT3ndGiWX2tih9RjFdpsqLV5fZ5F7DYqz01hLuqVy8UNq2+U+e4U0dBJFL63
dc4Wc2OZ2BXywFVTN77J0TJlAT3/pHvllKibPKiv47XHmd8zAQ1WTJGVzGQ57KUrjCBeEFtCFxxE
t6FlfYUB0Zg3POX8s4ixvvEawA1pxbzjuBQ3j8dAAY8c/3hTHc0Fb0beUNo7LePq/KUoJVvmS5X/
OOZVAW6mDC0mYyvKosFAPiiKsoWF/yxJLlXrjEnEDAPmOcNJYEQJ3Hl+Z2HAgaF8aflD29NzYKX6
mQIcKCMbw/3QsCyjBbqjDpFqoBrN5giN6Hwj7jmiDzNMwCGDO72f3w4fZamcz+/i+H2Zhb/SUwf1
asKeii3YB12AHcp07tSzK73tb76PI4RpSE/r29dlz/xNFD2zMhZia87DcGooctyTMQoKFSNFHMWE
Xg3vyPwkdsUGR+5UOIaxxybpyErsaAT8QwGHUbiikDRl6F/e0j+pdQ4wwO1FDkGLdZ1JML9w+ipG
pe4z3AQ1Cb8tFvVn8wiznkwz8cHkJv8BbdAEZCQ34l6gW3+Nz8WlD/XoDKJQ61TBW9FqzBKRmqXa
izoTO1zK4hyjYxJ2cmscZkirJZ6UU3KnNFhOieVsv9mh1zJk/eRbiQ0KsE4qkiHtuByI9f8zx6xv
FpNJfouSQYNxUNvWxjKvYe6HiUuon04cTsdgCZdVcoR6MD24mZfg0Ufbe0w/qTKzQezmcVTanYJ1
sMWBdjH0Ekf2udVHmH24cyLO0FiONFUTtnuLoGqD7HAMzjH7TmkPHFWs82d63aw6F0w1q+6kMY1C
HnwOf0hxITshTEF4fyjJ5dEMNlm7XkkT0R+xdnyD4Wrj6blFohagj2GB0OjhzXSZa4Y+nGeejrIS
a6IXEo4iajekpCAG3ztmgTEnWLR2mHV5nYiXuWhYjwPy11Zv4rBJMOYKHTFZr3wcO+0tIIlr84ZX
mzf0VWYQFncIByE8Pg9h1OWfr36QQNJhE4dl8rEaAkQXOvX/B1SEFoSeBYEKby4suE8/ri30KohH
0kC/Ze/d3L9nNMVsyBvW1QoQDw/qxZ7Hd7sySDHiRmZjpVvaNQ8VIq4jrZcxplTdisnVJEjFUbKg
NzzYNP9q+JFnZlYeNH6QhosMfk/ZMf45EJv6YMYLQA8gG8zIN9cbQA2G8QIOtJXDvlbcuftW2a3d
dlHOnhexUi4T/j1YgWvUHR6mNuSwk1IUBCY0k/ZTFKlZArp3cSzCZLLXoxbDvvQq2E4L+lnRjqS4
LfvHES6ooBHsZ/bhtbk2vUd4SFLXXlZJghtXHZnHymvyjtj04JESRsTl+QJ7PfTU8EZXO8N4l26+
tR6RQKPfKcYGkKCjh1kaFC9yizo8ikScUoluw3/rJWTKSitF1WlenMAUeEwwQZLfqSLruoXKHaGE
ibtmnFBsK092PNaxfYgT0ljTDwRs/G8j+8D4aDQxmxDDNcLi3sXjLrDSMyNrH8v4fO8+L1960iyz
VfjpsX2M5XHGDgTWMpaJIACb+kwyQZC2pTN9jgoxFbwJX/S1iC64VRsMUaNAr/meVvIaZwEnPVwV
iWZnKAS1kUleHitVZIAsT2ofjZ+RD8NKmf3VO2gBBRtNzqQ1D4W1LVnxGPKD05iV1Ta+GoUAzBje
i/L2iFrZyb6vU+W73lrlY4keBZ2gjLOPpBtjQOQql7qWViU8pkifoO9nzkSE8WyFT8HZRzCSk5ca
LoeT9uno+LXrSpKVEjZQk3Yo7PtfN0DJYvoL58HgNuqq3HMMZomtDiJHxkMqEo0lG5rEZCLnNxMr
7a/bNWOkFcVbFn/VSbl5Ag1RbigZOXpTR7Ux9AcBVl0SkATMga+NjhKZHVOo724FXK29cKLNZTHz
mYtdDcRY9l5w4gEhtwasm1LZC83nl/2F1+TsSRp2c6ISlzaTCZLfRkzMKxfZUapKAfXMzirMRlRr
kVBeb5ukW3IRQovcK2J4WZHs1/WYPdHEzPwf/o0YvoID0iJNvyYA9T+eXQiaElF+KrSCSnRnFuuX
AXXLodT4frr+6DfbrjXZJ69OgKK64bCjg+UXxgacBnHXtiPxqvYkVV7X7qjikrw6Vz8Bi57g6pgr
J1Zej5TcJnaG0FFVjJh2mBag5h/dcOo46bJh4HCZgiDvP9RiUSZJHjIslOe3ZrySxUEFaBF4k8tM
EmIG732bN6bXoSjhQ0PizbOrGcQQG8scL8Bf/+vtecttDvzsUD3txLOZqo53at8gUbi3jhTG+7xL
3lA3sONFoFac2uafiJ/sxpzDD0QT1esGyDx6+/J+vclfdkJDqqzz9DPSGYp2RXoTsoFhzlR7kKlP
yOagje96SiLc3v5lG0YhRSPo1DMfkHpC6bETUS348pryul4PgZJrx7TOQ5Ti59o2avcNVlLwp32R
gBttg+dc8h+HCf+ZVzL5TrEOs9B/GA715HtoA8PxKSouE9GAHGRDWDeUIwHTvJXNAD9hO25mFeft
VouT+dpVe0RE3Mdcho6G/SZ0SsuE/0PElqkxuNhSszSr53aEsAlzXVu4qSLvqTvU31akjrvPYY7w
7I9qm/ov9OCFFa+gv9yz9E57ccQLw+4aoxLkqH+52w6fPqGbpIcl1f5HY4b85PD5SkbxAXEpCrIJ
U+GEVuw/LqUd7f4eWVREcmXYTOkW4GllLwspLc6iCroh8lFPd54Fff/2p+D9jlDv8pplA+IKOsJE
05pb3tDJGNolsw7gw7NbHZ57F+iPpKsQGsEVb5jUOqW9tEc+LM4N4M57zu5bDVFb2l3PJXkRpl6f
1yAs7lkJcFKbkpwhjXJwARY8GEJMtruGBKLgaSIPDTIm5ybyPTAv0UuUDmZxNSRz9wfL2qM03SYu
lx9Aj1g3abq2yTHKlaNeu5a7eqexs94aQ6cQNP96gL6IQYlXaBxoqTH4xKz7K+yYMPUMraGCfJlb
48r0Qs2e1NmOLTBk1PY+C3czranM9xQQrWlyGPzpEIDMQZnzPbk/PI2q0oQbZejtDvz4LfNdHf66
Rf7CrRocuO+2sRE2TbNmnzmZ8CMz+rptT34Bihohjtiqz87hnPVPmWjP22rpgD+yjDiibbIcrIyB
GYhQXsGD5jgwAbqDXVvsMIdbPckaRz7h/jAeyE+sz604WtWAjd3iZrsLMAzOKID9fk+Y/gMr4Utb
eJTukbaefPZoPcQM11zdErAgW38/3oe73nTTqfzyjYl1aNsk5KycmU8AH7CJH2EzC3xIB8qx9wBg
J3DZmi1Ber/vcXTqTWg7wudKAR24ZQRoV9BTYnertSHCq99PeCHR43vggHCPyLH8Xdvy0lCPOqEy
3vL4bT2QVOmf4La+qvS7m6MbFeJ1+OJyKuN6ik+TpliwCGVoGW6h7slTCYl24eB6SetpomMiCR53
NBFxlHJypp6Mn4Yvi+skzFSkszS+WbIwkCkhIys6jXCIdm5g7NaQ6xYhpo5XNoNezrTahGgnNFaI
2eTQyP7ThkDQVP7EVRbFw2tHawNg785N0nZiWeZSXetlVphEH6r+a0Tukh5vzu2UfNzl7Dv9skgn
1HWKFhTK/QLI5Te+LBfivH1M1DRy+MhruUpv+bZ8Ich3Nwmao4u43POusCvWFG8ZDhNvxp7ObHLV
TGOhSorCFZ36obM1AzrWhH4KwBoMBoLsjN/fYzwmrBUTOstUpfxoHcB4y2YjG9j+TZLnbgvQ2J8z
XE/DxSn7AGphQdV3EPtVdXSCZ7bKMhsjf8aWMWDU50aghR9WoXS9B0J+prb3g93WGTm4lrOkhthT
3HjKtJmhM2MMUrPUfLgSbhhLPPrkP+ehmy/+ebQT7QIJi/hjxfZ99Nqe6tnQlVsmzHL/nqJZKEbW
wlb8yinkfFUcd7vUCSOtwcN4rjZlIcyG7r9RpsULtOKI9O9E4swKjj5yWw9672Mp3n+Axv8mM6aU
QqC7casW5NQMynQvmI1lisakwKOn40jO29yKZrp3IoLOVPhWXfF9wVPFfO4uEpAiSUGOTj7UAupX
0+7F0SI86ratdDixsVUX8awy/2C0ZMpRJgcwlnPLqE4XRKTyCEwsrm/nHIhkSCfAvWJQE+FOUu4i
/84Qo9O/yC/5l2w5mJUfwySqyR/s/lCbqVJk5nRmPlfwWbPFWVpXkl/bkN1kKaEA5GKXcih65puz
cSENhV6Hjniv5dEY/FpFvvFPLW/FagYMUZR/XBD9hf9zreU5NJ2DgEkEsB9HPGwDB7ZTkBmb2C7f
QzXYUSdrzvVwsvcygQPsj3FZZxRHH9mIM7wr+op+/Pyaa31tqqjUUpbkbnLk54bnUV84PaunVLog
3e+CswUN1cQmVRUcqAw+uwss3LaEnWXp6MQ84x2pFalbp1Ee7O2loE8krDzmjRWkUptkDklmx8JF
r54O8VtnQ5d3gFd5AOBBKZvfzPvrVt6haRwcqrQzIJXwZdioKOl/p0ixL48UDPXToIM6rt6NQYSL
FnFp41x9iwGVDzRBRRCBvuQkL21N6NbWqDELCrvY9z4ksqnrwz0B50n4khJLFFTYrAsfAljHIiUa
hW3DQe04sMN4MGLT7Ml1k/NZVcsyK174rC3Vh1l2AVeFWRlvj2g7E1og0qL8UmqJhpO0V2OBPemI
CChCoaD2k5/xOFNV5DcotnrPpC3/ZnKcq12f3kYJrArUgBHDQ/UB2QmQSt//8/YhNSUEitP0P68n
yjJ/IbwWc5BlloQ+PJ9KL/xn8UeVnwSJUxckGbxLyWuRJYgynjJ7AHU2eEy6HdPqq4zAZygDdg6F
J0SAjWdycAlSt2XuPUYM1phoYNt2rAHs6RgYRLp7HOMzP+X0iBpuXl2W2GYA1GpWuh8/7c3FaLtY
HEYTz52qA9k7FUCp7jFa7vY/V7a+a7Dd+Gwlec9slkkwgumk09rnk7MUshe5KnkCcN3MgJ8zz0Rs
FX1a80eRASsHZyoPK1cBfY6AJKaxI+QKUFX24cO2v97gycfKTlqF4HzW6bllOk0N+Pshs+P8BqgP
1Gq+ywrdvyrgpT74mbQK+sEc3lpynPkugwMsbOrt9Sr4yoleKUIDimymck0U8fgT7n2FvjLsv6gH
m5swcXGmDWRI9eKI5bZsvwFBOCG0MtiHxyiQmrwUczXBXmlRmpMcwYsc0QeKcXubL9t6+50MZgzy
0T5He+38c+RAJT2kWD584cnSGX/5aROVDCamtPMOtMgFjdIGktEURFGNk85G4Bp4ffyVXHC0yRMm
4S1jAnsQ6YwdFuDFiTh5CAwrQKAbm2hUVrALp9wwoD44e3T7xEptlc6lgAe5fuzo7iNsUf8XICkf
nWXTLAcmus7RJ03NN8HxEh8cSuPhpQ6Bi6v9Xa6ojf3oXRgEpIU+MTktrD6/4KD0on0FmlMB25Ab
asGkMBgyUP3feXpnFA+lCHwO/H8DpZnWkiF65PmqyxOBFQtjCaQTG1PCJc2lAFNOgKIALOjygWi/
PFwwWkkb35YwuzAubRNuVlqJ1A/VCAG3+auoRKMywRlsU64NU1aOaROVyH38L3E7IJW1JNgHG9/+
ja3VmuzvDHwGA9v9dQpyS/wf44Gw8UhKdRlLpCRTNZdMjXXXel8X6mWFWYPToKaZ0wjd51EQxISh
NtIutrb+uI1BBZwQvJQLhtkf6ZP2DmKn/BJVKOyZZ6Gag9Q8+3+Wk1fgrPBGXInVRMKCTvr+HSkk
GyG6l27TUmpmogQvciRDFdjiNYl/Bc5cLQHMZp3Jz1t/mlaN1cXNrQzDTOvITTerVfhDilaIghBu
PFAyB66b4RUV2/5p12al9AenvLgxOKOYlrxZGpT4SzpgqRVNVMLxgBpiiE2E0RMpqo151gTt23Ng
HvHWW2Mc2GLv+FVmOJ5i+zFHs1ygpq/uF/uMycRHAEtfyk1wNLJpFXNUGsqruUjwRTi0AJON78A+
WkOHzO4o6gWTKOs9rEfIzjSins+ejrf7ECaM8IwBa/eiQ1AsemkJ/fehVq0SQUBXUkZ85OvanSZx
AzILazQ80YVXyzNNRi/B0kdiMcOXwFTL7XaAku7YZHP1ZowOcrMbSrVZMI2JsDNQ2lfE2D/IRjeP
hK4ti1WzLmdiXkBzWHVGky53tF0UXh3puJC7jA2D0I7kKynLjmplmp8ZK7KKgO9pdxWRMqC8RoYP
jvypyV++P0x9wQP0/tCpv+j2BdlXnz8tmtjzEZkKfkTiYgD36/SK7jvakBmTRLd4lDD3JJt3tx+6
pw8o/kEtWPL2gZhsK6bQMyfd7+Wuj0HCUoJVuOnas+60R2sGG0MqwTFBVnX6QwGEDGbtwb2vJKnN
s/8KIUv8UKaKizn7ucfp7MDlSVICa47zVpsNlXIp4IVTqgIEQWEgUx/hZlQLTWDsxVzb8eDy4FQs
SpeEoBnLoroGdX4X+vMn6sSENaOpsEILryTevlzbPq1viQJiWErZP9G23VjhRoda/GC6XdFaVdYh
H317Ei1dwcIDgMesnxwCvCHfUDSnnWTkvYYzKwdOGm7IZ+mPNFlNWO6el/tc9TgU1Dkl0oODlP7k
YLBF/jB8ICEHhe64aNLIzApJQ+Xye65l1G/hVHRhXY/RQUyITSFcagAO4PbNBR7h9BLlqG3OzF0+
H9qQ4Uftx9BfijRWX2dt20zsbi9cd6Tk+QBwiMJGKi69p8aQ2Hc80LAjkF2tRBWBs2hW2QFQwv4S
6QHzGlM2z+jGJlA8tZI7LsA5ixIrGnBtUaqSLrpoIzCImDZDj3Sjow8Uz5GBiyi9xDkSkweHu55V
Uw16t73CTqyUQp35O4hzqV8LBa91aRqRJAeDWrC7XrsMJiV5kK483aK9xujbkw0dvKhZXwE5DrVS
EhrQSvV+lBZu0NozEhFcXSvE3pDmU8tAnHSqj4KsXxtOEGicVoBJ37mSdKTFBJLY7aVbH1by9ZIA
9WvYW8SvQrScHorl0Ax5wQDRTfP1mt7L9dr79CJfe/9gamW3tuxZRXRiTnaNRYPt4TapnjN48FrH
KMIBj7Xagsr3OGIMoFwiGh8oJeaXE2umJKpSi11wYYmsTwk8cEumEFZmW7FjRX7GsHBscSONn9jL
A4hZ/rNxkys1NpXyW7U6IhOcTiU/VimujCfdvA4YIcN2K11b7EvjuuLiJt0WXGFFGM262ZG2x2b0
VUG6BVfZVxg6dQUUsD+3HFW/lrnw4tkDH457w4PiW0bZjzv2wr7+QcaTmBX0dsCsFPIhqos74quj
NLiD3KHq7O6D5tUTybgnsWKXeezZpo+wqFTm5csU90/mlCiPYcNiOJQsCD3KB7xZYUFpt7axx7Ol
GOQbvaGLhWMyQZgK9x5c5xHcZxMb5JhnhWxd0IFD3adqqrlaRUhSi3HC57a9faAdTza9ywyhyEuf
XBgpTST8WwKe5i79N0CJqRFcT1s29CoMglrCC1LoccHqDa03NxY1kjg0+35Hg9JkwTlDUXgp1251
YSoAOWXI6RkuAfJT22P62XSgPeHhgEQ6XyNqGm89X8mxiz0JmXefrjjS3Jj1ouOE5SFZ6s0O3gzL
VGXydrqTTZNQ/iQFEQVw9P1PjyEtHXOlRdin8hI/cbzvxAtz9+x3MjZU6hko5ZMnvWrwmc/wHRsI
qSytQOIU9K1Gf/V/KYXf3vAtqwcAx1oT+cNhQDfpGB7eDADxESmCNIYMCtUDmXG5bd7OwXmOcL8R
+wvnwzGhDnjS1MH7kOXhMtlhDnm94kRfpyeTyi6bY32yEK/YoBBAKTipQjoLrseloZC39VIITaNY
d96vNVT3raDYgJsuWVmfYyyQervzkl+yycLqF8qnFXJhv73wCTYQcYgcqbxQY6LQsr8Gs3z2XGtE
cimhnuPOpPTFVkLjKEmsQu09yG7xnLSxA6BiyvWefX5SUtr0gX2WxDlmfhCSNVhibvqcrMczEluw
CyPTYfODa4dMue/uaJUKZYkrQAJ4Wr/xdzVg542XAzwYFCntbFjznqgsnWeqS8CpTy4u9gIQHwPR
ZNnd8JayRrBcWCTQpNq6zuDp87G4PHMxn+OhnMoZHcOQvUODERnDIuWAumGOrpI6InAjvqsHiwGG
DBzdm9wmkQ9nVP5LZy/TzboTbKmwTdNcs2vD9ptLjWcnBJgU7LDYvUXQA/zzxmKX788j2qoXIMQ3
79OTOjz4dEQvHKbKtOuhvGMZbdr+8JZPUPiSMHSOGgiSDdxUBF6VAkE4ISu6NT9M29CGXKdPWphB
CbksBYblEsNptmCOQWhWw4rIIb/ydYVhRoWQYKwEw8nHTl53gVKqU7vD0BPN8DOodTeHxVcN/Pbh
Hb0hIdGAUZrmgPfYXYN6TXYIbwI2Nm49MP4C/FmfurAxCV80Tkl1WAT3vU3aZLMugQaxhemHvgmh
bKpaWaCcx1nbX5ENVVyHwkmhtP4dRodEWMuETecZMRXPmm0odE8GxcIzPApE7Jhy0KB+VdqUUZR3
5hAUMN28mYliWNEojq07N5dcvR8etSIhG5yu44Zc9VF5qHf9hjc35J/aqbXqipGjmcTajF43WHt8
IZd4z8cUVDNvRpcPso+Wuz1UlKHWVmaMTI46bU21Z9vRl8o3tRSXswv/gSyMvkryqjlSmbnSiiFv
iHaPOD7v6FYQE15P0HpUcjFskYX44R/zMkP33Uq70xGVmckY54COKSj2pn8iN6Vtq2+3gN4p2M1P
7RHYVE426QjR1hKfW/5zDMx9Q0ZVdu3fryjZLBoLzK45/izS/lh9fDeIy+IWySCZdE9lduQ3B+B4
hXsywD2ZsmhobABlDHRO32fqmB6T9s3mhhYtx9pxOBF9QAGpGv014s0nErKTgnBlNKkNvBWwqrmh
Rtpp1WPy9oCeYkqccdrSTF3lGJiGHI2IoU7WHGg5VWKq+KUGLAkihz5pgKIn30mtRs79qZKlyFWz
qoC2p4tg56fRjjYdeJIicpPDEweXGe4dmvESLsuMmeXufHT1/3pgAAiGajgsQU3cSt+JBCjcnkWY
uC0X86MAP+j9TaVoRwhA7X4bjqp+JMklv7B6m3EkSAKuSH5cuPcg3R5zDMVIyCBh0Gs4rzvAi777
fILVMH72g+5rQ3euugUI8XpCpkkx2ALLxepy/LpXELP4fZR3tomalXr7E2kX/MfVc0bh1zTgi7rR
M3pqomoTfWskUO92E4rkkrcOQZU/CwDZ4yH+L5fa8aYLxdzHC5Vanw+tFyDrOodpcCWezcO0GEPG
47DVvRjDl+z7RVAybDQdvQUf4ceOzPizLDYWk6XEBz2ehiqc4HGpSU99YnqFrUBFl7Z+HhnWV5I5
mn1h1YqXQ7f8h7M2xz0oUjK8sRNDThVzIZ/JGUmDelluLlTJuRIAhge4a0i6AtGdUHIY6M2WeZXa
dtAtclhmPPcrgro7NWGemwYLyrgiCc8jzCXOe/XP/B+2WtikS/yRdxKih0fcxub0DYBRY4fy5Q1Z
k7htMsqQh3ocCJ1TZTdZsl2hk1KmjiHRXkxt5H2zqlOBUPf44gR249w3y7dTWuhl3jYRYVfyRfE5
BFt21BnzZtrO+V5Y2DuGGUFdwYCHdcCTzd728nGo26po6/8zyop3hM8gNs2sob8kTHyvICuXa0X7
j0yrcaRHsZFbZoq3mBCqf9244e4an49Vaaq4/zXl7X+dw5hJ3+agbB2NfZoqK5i8F9+cTE9w6cdf
hIX7MVm7hKVaPlELgcPajrcQjT4U3+KWe+zHqWLwda6habHN/jyt1/WXqoZ08xdXb8Ws9hcan1qz
Vb9l+gGG7hdpDPbhL1NlNRaZR+mH7f2QvIaQWjrPVxPg0NmQ78LOs89IYJNWJxlwDQWqarqudTue
eYYuU1R+VpNN+uqSfri9ncldPJ4gNgVTeHBGT5KExDFllYYdzk7pHVY8Dc1UouxMJaN9QKLE/FKQ
na2pKFxAloRjstYSE8mYDvkqgcqxbY+zC4ABJAv/BJZeX6C61dzhlZrGSFS1B2vIaCI2VQ0/eqew
0ZQ3VKmG7NhF4xRXMrPnE6zxrB5fHaRHjo2CmnlGN9Y8vyb0dfbYFELGr0rMuAy2WK8ispa21nV2
TGVswTYVM0w3Ss1Zz1KiWA7ymtHFsQSPMan3Nia52BSLS/LIEakmqmkF1J0BN0B2jbKuMID6gE6K
3NvBN6QCyh1AUW3uPUuf1GYnqyxxHq61brzaOE2vCwfvvkrtk43nopvfFS1cWFs+d1FXipJewk/S
pqVhFzD96Vs+T6gzupEw1qRUiBD2eF0vqAwyv8BnXZVKhIG3jNMGKv4WMOIdowKo/8iiFsIotDuO
FetKnyUpN3dbfmRpgMnJtNb1h9By16IPXyXzKU7QO9atjvRcFQOa5q1wvsD02ZhdUtHNvJ6nYmFO
/icBANyASlwlhMexHK3lnGXyqpNaQ2mTyD976Hcl19gaPR/QC0EsHsOKrs1VMDENVAS9wKIxPapo
Z9mW6aODZDa4gjLrTr1abzSJmABRCC0dnErT+7goSiRa9xMw7k4JOG2AaGJGTA/bYRM/kqERAhcm
FGb1Tavo6i5poJLYjTfo6HdyP1hotRX+W5x6Ed1d+wq1qJ/QPwtauW7rgMD26Gf58jdROvdwbac1
7rrE892nIjp1qNRqnxFaraNFxf6z3tHx3oftx5h67/2A6+MQLMKlg5DtpExzkzpGBGFGxie/e+V0
nvDbcGE9NrlxUZjNndgZaxzjfSdOpl1ZKzBr6chE/Q46PR/tsjCW5n+p1cfiuusRZPWWobEHNeAg
UamzhbljtViu7JjCGFHX0ZxBf2CbLHdqrxZzMAAeLXcybr/glnSeX83y2CKD6gQGNWA9oAvINMMJ
4Yc13IZnlsNSxOT9CY5qewzRzNy6qHgu/fDqerjOqr3oh0XpGcIWusLmtORA3snj3btRQMk7EFys
Pyuw97M7RIdMvZDApGm8brQMpc6+VAlZ8vSpLxCGCOYq/k7kyRaiY7FOdGP+J7DrLVWSsI26XQyx
opxptxRgx52G36Savjqng7q5uJ6nEYmNLxCi4kPfAc8iEXwkl0fovcGPOgnGZwr3vopsHcRC/fSm
fpbDJKkTnQIHgtrK/34ueNZILiy+1yIp+hrB0UVIqhLdNc0TnNhsQGyaS0ixoYmc+KYvwqNRk0HX
6Q3LG9sZzDJysypppYsvOwSlhEIB8xWbxY+uTRz+XoI/CmlZ9LNB6uYAIAJmXHHQiEut6pNR1SNn
iVHDt+xslNz5iTZmhujKcY96BykYOJVs/6af7RKVQIGrqCrguShasI+J/KVIsKWmQkDggl9dpU0I
wbh2Pu1hKmjKVbO5PLA4ziBZD1HF+4yYem4ztfjVqBqnPDf4g824C3QuTkd+mZnNTi7PqFFQm8Ev
+Ik6Qnedre4oxY4vq8eZ9RwKl5iBC/pyfTBJEudMj/eFemkFjSiDGBx4scgWgvANvkCgNyR3ymO6
6FfC/TlIH02NgxaE8071zJoZz50Ynx6qDeA597Amllxo8I8RfiYTq04b+KZEvQPV3s/6Oyvqf4Fa
mXgRThcpks60NfcPr/60NBPJkppnSEOrQ/XVgG0Iv0TARlbk6Xr99yraYkpUHGVsMkHsZ4bJXyBW
uYjSStaKz8lvFdZSYPaApBG+7vO+cZzI30IE53o8eV/LsHb/b4JDV7B/sGRpb0ZJg2ptqTnyZhO0
X2uthTrsesipb00maK/ZX0KqNGTGpdokUxS0zKDNGIVG6qkT7vuHdVR761D1JFvNz9lWbjwTD7r+
LjBrIH+Tm0zYJWVWvnmFyMw4L3xOGduny0k96s0ewDS0qtwqSojPvls1Rcgvo9LwH8lLGGCvZxrC
hkaMVe7p8VzhmMWFdUrKQXIHDPTNKglg0D2F84fN5UolF6dDoScO01U+5yJicEdDB/trs5I4nLXH
Ct5Rydh5F+093HbVOVtHjPhR5fqBQ90a4VokfqiBr0EYM1lEgO73uJ6rMzA2ZG+E5VU9rU3cpDVh
ax2Z5Dc+b107OOfjyH1fpQ8+kN+dGuCiJ8ykSlyy/BVE4dqxRcpy43bNO3yW0fXT9YPQhTdbg9q5
r44vGtA9QDo/gtcgdf1PxvaIAC7Uo8b27mPAiGEKj4yYyS+exWpU4TJnzZUOTLJEvbxQh9rUD/nu
yNwjaTsZEDxAYvLq3/3GScbLlP8WTRDc9YSYCKhUTBuTk+/T9hYTOywOdSWePydMmTyzrxL+3xHs
vU+b6FgKht4Ww1ZPgAqxpReec2WlXRQnUQMkx/ydeyBYfpYruHb7+h7/LP1gccmbTiACvqFIxJJf
iLmXwiAKvpFg4Ll9/VyloEK3HhV81XntXh8EBpxNIa6m/fuBipska3GHZO6AaQI555IClNbmZmKU
o1l9sULYY4LUf9eLVvBnvW0lt6tnC3XxvoQBZFYCDKcO1TpV7ZnMu6JAGjehoD7+ffbQ6IQWygVz
KjWX102bNn9tLnXCh+mRFuLd6Sn17RuKw0fbXxWw1x7p3l9O4S72o9AK9fqcviha0zXfsTu/9qBN
3nGQYRpIXnK21KO1GM8Tn0vMH2CS7m2RVErRMAtbzocHDNCfKRUmWD0EJ+xnb9ptSbs6s/vfTlJF
WiZKcrVcxxS+CnCGbVeY2kC9qhiMq1SZ+rpsUz3LlQ7ibd1R1HgjRAmiGcTCgtXRVC4aPac+Hfj9
vu4IIx3ihiqVSIJG0rMNBpPSejuRqCPOZ6g3X4KvTea6XqoGYUr5lsc78eetYAy9gWASzpl16jBM
iWk1hel5QeH8/GBxx31Dzi7U1Ijv0j9uD5/VkUxvI4Fk61vJW2PI2cci4h4Xub+zCGxpWPfJOIlH
iiDk8HDVhkD5dcoCDnL8If2oLc5S1c7bJN2u4bTN9mkARUcws++cVqyas2/bOZp5Yo5iwcGMe6vp
Ar1JYBxAiznhzknWQGCo7Lq1LptyxDt40lNNk1g5nebqIrmHt034Hkm/B5c9jClLXHPM+08Fzuj5
ZYjmT4/ymelut0SRB8kRiYCk1+YkPjVlE++kOFJ8i9jbVPZ2UqqUyhfc/MgzPzBSdu2mjZM7jkpH
tka0fTFFIviGRi1HIq0mRa+LRovRG2Ajc1tyExfR6WdDJ+AGGh8PIbUkYSSl2X4M8mMD/c42rH7/
KYFJaXlssGIArmNfWFwi/n1tV1Ys26fi/80QJ4DWX8M9cyTmSULYnHvNk3idfR/0sH6Ng5xE0B0v
W8clkIlJsbz971c1Gi/QccCXYQqqnvkZ04VX0Uc5Z2If5uEH9iggRjMiVl345FjzaRLxRi+3MiVr
w+wUeaGqhWH8fGd/+WlJKVHD13Hz/2LI4EbxNqUU2UYx6zzuJlGihjh71zO/oNkWmqAIrRuoWst7
mVXKyh/XJtLOxHFrYFJyDausPO7kiJ9wg4EGb+Jrch+8wrjQsDLISoVDoRqUtjePg8DBvKQy02BY
4CvFxioVFHLWlGcGrQbk/AQK4CWaE7yQOiCLfr9mYyzhd1VQkXvCCkFiMVcohshemSfVBnTTJRbP
ZxdgeXUhIT4vvy8+Pzk56e1XzL8/AMrgG2I+WN6TlCwav5gJVKXVWsj+ufW5ahXeNdSAVuuW0kwJ
5rITie8xgTjeUuhG3EhQQE2CxkzrZsfoyrwHX4PzIzQsftNcIZaQ0KeeU8Ha0YFL24V9lkKC0Bma
CDJcQEyt8/gNVZ5cja78DlCeqUgVaJ3JRNB872AVhCKnYDWEfnPzdp9vwtBM+brxd31IzoeIILMM
eTS/VcYzyEy63cwZQqGmC75z3DNataamJu1uVEjg7xbjb6LhbtiuUD8fgYCsxQvhGxsNSGaCFO8U
HPQAAGQfZqEeTjykibvAMt1cwIXVOukwlJg8AFFjiBkr6eQbueJKHTFHNb/Y/qSS8tQa45SS8kGK
d47T8v8n3A6D1BxEdAbiUxBkmmq5a8aWtR8RQIlm4f39hJASQEg3kax+U/XVGZ1O/qB8+t+JgVTV
CXawdh1gGN3G74d6VIqKVcA6Xvy6X80KMDoVo6gbCizhfAEsm8nXN9tz/QVZ9GVPgOlAaTyuzMu5
0NdA+Q1WmFb/hTKBF/uSSfW6+ddI/qOVFsMzUyVaSsWoyKr9JrIn/CxHFLPJaQF7CdeteiHXcrtb
P2QTMEfZlHzw1IM/DwBLtvVBzEXkuR9PoOUs/CYFRPIHjM6zRv9rJCwqTmx3oWLmkaLBxipXZp7N
S7SnfwYN6/IJjp9tM3aCY+h0rvF6OSRf+j0XvyOVpUjUsBfIqRO+Ee2Lx6XzEJ/PhQWi6A+bgzF/
8SPPvhg0Wqkg5jbuOEXHiTjWregO3ukMKOdH0BLjmttmvvpcDJyAFdFhc2urzUbNyc/B5nTa/AWc
3dSJPC6k1NwnLtrZGx5hUtY5F0DkOwB4ckHnZAPe86byL4oVXxYGMuVW1UVIlxd2LN1IrrGwqrTa
DgshH2u1M2Ta97tn7hrhIY2oU4mg2aVQl86KgYMoV+JfMKZFwEGpGtsCprZs8KTSvLsNQsPDG41f
Q39EUUZayT0sdvzp7A8O+XM7rgTz+zSKF6cFVPsn/gK1BavbE3DZHShDRKpX2RXQFPisjQKrezKe
eY9OFM3CEKz1N37mSelhLTnjUIQJCQckfZY5YKyLo76/tmJjAucMbH1u/MMPKLJE+Y2nv8a5vdxC
t5ElySehH7KESfYROghG4TTWleFkPP8yyRv6iGqMuGrUFKiHQ1li/E4jY1uy+jI54PbvKDHFgYnv
wVEIgQZ6o/O8JTczFMnc0IoOdc8OS7TTjHJdRCmqWsXaG/JSMXsSNOdoOThKkIp5r0bAnD0eDvo0
taWIVtY8mnlwOlMtBCOMNRHSX5Y38MWoO2mRV5BtSbfy3uX4dcVMOxmHfuRGhRDGK8FdTyevvzBj
CXA7gSh9QToCq53asddyOktJ1OckcM5iTebpHShoMDsQo/IMJewEAnx8r0VL4lZ59auXRVOaJKbc
0ti33LarJdI6ziS6m3qz8dA7GD1IanoFbdYz7z4a3pbRK6uI6rnwrD3LlVaUgSXm/IbRAa17WgCZ
d8E56kUdVL0bAXf459i8mekzmDZSUP36aHPs6dxdlGtsC76TkKtixX94LU5vcrG+htwr8ftGgDGp
A/F+cxJTOJqz5WRyV9uMx3vLtjReKptlAxkbKXDImeVHU92Wy/iwdakwinxNvE4o/N66GbP2FyIw
THEaJ0SVoFliIAaeU7zqf5q4IOWf9CH6qfBnu2FG0I6S+cbvgxuvVygtsABVijDSolKXtm6ucMI7
cacda4HwUR0r30yqUJ5YeVJw5FWmApm5eEpbCwIyHhXP0SLTzqXHSPPIiOzU/JX5ywtT5C/+nIJJ
wYgFvIr0L7zFyUs/uT7b3D9uYArMvjM6kPxplrjD2+9Fv9rNot8Jf/4x6H8nqx0jNod80zO4aIHm
G5+MrXHLNbAcHycrIvutPB5ddfjl3wnv3BD8bL1BkVN7sSmgLwsrGbKjvaBeKVTkhadgvpCkS9zM
rFWTAbflVe6i3GiO5mCHuNaymGnq06jI8ZAgMoCMtCKh2ZZKVBNM5JHQIODNsEwww0cpJcLEA7dJ
/j4FESVSfikFpqHpTaM6BqpunJ8dcFMr9m2K28Wr7QO091rHsRsFd5wG0aLflMxadCzLXpC3F8Jv
u3mKmPjdk2SxPx/EfL5iKdxH/4GCVBH/PHh5SqxGlUhh4+JvP5v1ECWxS9wDbEcHNEee7EYoVXYL
9lPgLZHWN2M9Dj6iEh3zfZg1VzMnVCd5+4vyqV3XCu1Bpjkfs9K5jM8n3CpVYQsdjKacnaLvxYy1
a4GssIr1vKfjFHJp7rp8Ovha4t0JD/9+qCX+QqYwCexY3EugEJLJAZ+5OjwsQETyeVgrEedh4/Lv
n/AQIa4VS80pOk1+hF34hgMNRd9xxVJ6jNeCBcu0wDax5/tV71H3fxM0wiAQIKxwn0HmbudLzz7e
3gyTcxBnlKT9rscljgFF8niRnWMKVCUhue0coQ+STbHMBkqEwolWjSRTcROwmwgS/qXxGRokqGK7
XuqYV1JpYsP0MH38IstS/Z9HXZQr7/MGkJg6PPURDVnau+IcSQUJp8DV+7W7Fo7ICkPMP6OBcRLd
IrdqeykbjIrJz9uCy1R6ZFb5zZ9p5HFnNnY1Waevs6doXCJDpED+kTLPiAyDXr1c1CFmOZKD0z2c
DImmsU+pkEL0OkBSlIANRn1NaYMPEabStXnE53XtznAlM/b4+Arx6bAJ6bIj9+gQQU9oCX/kbMdC
XB6T0Qogj9jKY8yf0pi8wR+7Da2zllW4IdzQr10UwSvdk0siadL2QrmdjluFI+daid29wTmLsxgf
VA9PCvKcPcJJBc/33VCZfnSnEJHDaUWIA4MY5Rcd7ctQx8rMEtZQ+fnEvzcwFtivPT0tVSChY+DN
2BaxL4j8eYWIN+ZjZzWinlMba+/kL+k6T6/lDFdwWLrzD1Q4eSxVy44exRp417pUSwsWxdXEWQu0
+NOmDjqzxbOGIQVX7wttIH8vOUI5nhDLg80DOxqL+go5G/OPuCQs8g7vuiWjPLfvyVkNLFXlauIP
RYtEo7gwtJe7c0OEU5HLBgoUVKYPp6kPdEec2dQvU2GxnAGi42gvxqaBUK50W/PHkVQ0qSQmevQx
R3IdLX5etu1VK7YXo2DBFk34JEDBVHRZXyz+RB6hxX6mGzoR7ZA9wdUwoHxlxkNtVL04uaANVGpX
UKfAfuYIMfRJTr8zI0qniXpFvO1DhiAJ237d3IJPSz/NtlshJHD/p80Hgu925HaMZT68leWHbFmS
JuH2aoOYTQgy25BXDyMCl+1+IPa0BX+Q+BEU1MvC/k95Q2t8MVzjPs45UGB3L+9F3qLdJhPVx/Ph
H5WxxRDx3AYiw4JZ+n4dGz4l516JCAhMNOlNTVACsFX1OpKXtYIUaw3g6y5MfXCasn+J8w4k8Ceg
mSQFluCnP2j7lvEhaMv4Pms/ivkFnJZ/SOwZuVKo1aQ3QTzlLB/H2nmWYUVYT6xxrRf+sXccIYw8
MqSTJ9cwLi1ynyHnAj1DNOxbRY0tOkf0Cwq+56iOjWE93EHeBqyLIqrqF4EJS3jfkp6E0w4KEg11
kLPXReJaze2i2jYpT9Q5jcRDUCKddvpq6gvfhPWtPK+DCI5IQhErTWoCBjBClhfGf8tjIOxzCir0
CXONcPreU/kSqSMCBfVsrOmw77CX1Z26Pm6zR2TKNOmz5rD+CBofRq7uHRRHzdvxcEoGTwBgZ9QX
XXkjar2xAEq+DkPgRAvliAzvLDgPxtO/QTo/1mmzssy/yOeFx3ryjMPGi6+8XtL8ojpuP81UW29a
TaPorcafWS3IIrbZrrAgHeOG9vflgQBsjsSz7t+S/puR6Y3eCmb2g5yn9vjNw6laIgn5c4+pD5cp
gapM9AQNlG/5+5+5BNtK4BdY/YUhikUsY8Ns9RgCy5ITeudXsw+JzGUdEIigvPKle0I8kHGz8t4h
Pbrn0SkLiFGPNWXFUAvkvRhA2InxP8py3CDQfGBSYTE3YqxA0ID1UB15pfiF/5HonjKvOp5JSI3r
U8l8rj30VljCVq3Q1KcYiVpH6jcEt/Mq3XS6E8IUV0QQWvBgv3wXMjQ3cEbRxv/+0ZQztOT75qdJ
IEGp/28Rue/s6wugGS5UGvL5UQX7EtgqGdOSKYsqHCpwOSHmMpCOpXwQOhrl/QGboV8G0Mp8MpRk
VLgn4gQRDzJ77gde8EHlY8/a3kgB+8JX8LFXTvgsyEkEB9n5Yn5xL56ia6pmmuYbX7OswOZNB2KG
0AMd1/WEIdNT24+hiyigJPRlK2gUr+mhrlhdugrnGRbVoMwQVwRiMopPCAVse+sXUuo49PubNsJe
9rpLdHCP9MYwsPtSWr0u26kDh6+DoiF1iZAFwF/t4AXgwTfBgaw9FjaasWTNOt9wCGOSzxemU3o4
yb3R1AFZYXR+TBMx60GIxRK3u1+/sUTqeol+FEV/EC4GsXPf6cZkQD7AUZLUgQjr3h2aISSSs3vN
QfjGh/+DOWaYJ9hP9flNItDKGugi4SWEtA/S+zhhej4+vh1VthOvBIf0L5yFdMNedxInYm5YJLpo
2x64MEseqbLvWCEZ/xMseSMB6j9TH8CWQdA7vrR99ig2G/NTtVXrL5xYRgEkEqsAIAZjcYBGoL2s
KIYYiD9jB62WzCldrfsNnE5X3KAXxS69YVrAL7HPqu/0qJzz8vc3b69NdIjQehAL+dcfdavwZBL4
IFyEB2lvWAbI19XWgruYI2AxurrgVwY8bz9JVTxtZ/t8D7JAshjIxT7GF5xnyQxBEGJM9bb3YdG/
2nnO0MYSWlAkQKb9ZmlfrwiCLYjn+/o02/MDzGhE+J+UsN8Gk6r/0eZUnlADOsPSaJAQGy+/D4Sq
T4enTlxVmyZW7Jw2TWu05y1EbNPvfhzgGYJuJhy51P+hQoDzl6Jzl0VRTn2H0Z1X4VGdHcUEkn0q
CNdX/O5AExWhJtMnM7tVABIq6ad2oflJ9ntNjAS0b+89xMDq3O6RI/GS7uLQKdDMGRfH3P5q4b8t
y5riODxpH5e/uLtB60LBkvf/wRxaqlyU+wax3ef1tBF6DPn9XenXx7u2rNhyN2HkM07NBYEWOr8k
/EfHUP3/niUZbTxs8dTVuX2vbVSyQ2T23HqdlDuK7iFNZjg0ml+JE31MKriUZCWg6sX6VGOSpn8p
eUQhrZ79itx1TIn/boslS2FQH0bOvmz+I7NoKTkoUEdHJ5XNvAnRFc6uf9gj3nLgRr2kx73LBgrU
oxS4WEklfQcmWd2omraDFF+855W+4RU8bsO0NpNSuFGZTTCo2fCBbZjfk2hYjXCyW082vURmCogl
rz1Qf8hvXsJ5UPzdLT1d6vwVz9jlvCRzz8jH525V9dqeE2/D5W906d+E9iiRH1hYsuNdSq1XCfZ3
B+dSbqtFwrGOeyqpzCcdN8t+fsAyI/7NlG0ENEZ3TrdxbirbEbXnvL/2na+bXjJceOkyqb69YuCA
MFJlXHnQojkmNOxOqaBGiNxrE9P1NS893tHnfDBllDVf5B3vFfGd0M1PfuQ8UxBuoHCWcbZUHNka
NT5dlvFuobPyWV38069WxGEBFjIMnr/aQySIPmth4Agp7H7lB+kIjn6OWLvS1JeiHRfPmyL/k3td
3BvzP5ovS2ZvuiBJwUGmApysFzB7HoaidlJm9AgwJKeBX6SOjK02K5CmVb0RFwh5/yf7o261RBS/
KrtG7jLgUvvEFMXewN+9zhPDvEHPuKz5CfoviO0vHJ5n8ORUzDQLavxUi7vTqP1+DU/X04iJ+Klc
pIDxx8LjAI02yL5f/mxwEnnEWdsDbLfSNQ/VCx5ZajmIAqoqkwPLNzGu0Ld1/ru748rYmMgCrcRJ
WcavZT1wkWAi3RZBEnC+Ff8kYV7sWJHF4waCSdJF7rVFj8VCuuijDbuYHMiIl/LD1ArBbmG/3pxk
2khZdMNcneusCA//nARZpQ/+132oqd5lq5ar+ix3iSwy+wANoagjKQ/2iSFdwcJ4m41Ls2X7Tgfh
/TvUHl7xedOoJEH1gD8fymkBX/2EAo1H9OSwQZppLfNaLh83HhtwslHPjTDR7z3uYWP8rtPW1bTp
uhuPafX7I3m60CsHqYvi7meiAAF+dvA+llO6/KNxoy68lVWZz9tRzAt6Q4RGvr9TYDF7IhN8yB06
TmiZOeTyCD28sY8mnc2lnhWnVhPfUMpI9gMGkyk6Y5I4oxzy/PixUAV/YsaJIVwd17fh6gOe+8js
vvPqs2MaxYd1ATJgKZ9GZbX5e84tYLD0CUsDjspOI7MSD9uxexnX2eZI2ljbGBMRhuFUvpl28aUJ
rTboAzU3Ig5GmtvOVcAarzcCupmnYhppk4/ELWxluKOH+gTyXzo2my441kLZM0CBvqtPnyr9h6AY
1Pla6TzPDHf3SCaLTA7tH9Kq13UYRcU5GtfZzVexyEo0hbB24nbUQubWTGTN4WMaD3dLI+jX795A
svAVlRShH9cQs3kXL11YMUMHZEfzAouHYNYMp8sZDiVYcN/dzcs87xIzn1FbisLGakA9jn4RMseR
5NlGpZ1K+ovM93xxfvfikS565+Gi0SyGAsAl5CYNNdFqiAMMJcOwt+qEtm3LMKD/IDw+HzCdX0I/
Y3lkFdlLM9d5ct1uUrOwMMk3pXw4Mb18Fn/10/+mT6gnDppBbIxMqfrhbQiDHX1f7dgzSWt/Eg97
RxuacfGHuElQRec0PI1AH/VoOIsDSGyfVKSlDMv05MtTub6Z/HgP6jml2yPZm/pw3ShkFsYzVHQQ
2dHkIvjL7XGU3LLSfd1wh6H7auDGPlLcBcacG/7OTZjQI0IvltrofVXy/roM82X/TMjm4VF/5s+j
dG2df/DXEZlv5DrklGpnkBGdJZcTQuvIzFTEF9hWObf+ZhbSW1Zi0j9alAD9+gBfQ+IBUHH+K4Ii
MRQRGJJSA3IK2uiuaNnt1AKMMx9Qp5Bu6dzVhyDvsIj6A1Rp0uUfh46JV7HOrE7UBabfcQ1/viT3
1wDSGHaBxdwj/ATfsL1O3914hfT416uaCPKxX7FhdF4LX6EnopPsGVzLyJKW8gzKxQcKovHv+nW4
/9HtOqcCDRXOa9fRStgAxHaauJLk0LNDXvpMfTCXOsbDBEyjGJMoox2VR/lrESCmD8Xih7BbvzEy
8Mrtc9j39YsKjq1K9P8pnHYIy81HS7Xt9q8ncBs/5BeZO04xdFeE4p4HNvmFaJrbzteZlGR6xzn8
3oWKBgiKsxv06DFaQLBDK9/J4UHaGxmDeBD/3ofK32FjP/LCK9G5MGoHLM0IvEbODR5WGZPFk/ms
xJWDYh2IoNOsqf29VxjK6wi17LuPFt6Jy1iE5fAsuWodB4jdtKlUBrbmAKur1fEwljcTPpBwuaGA
ZZy4ARZuG8IeS2zfi2dO+Z0klBaIvkkj9Eeybx2LrTCGIw+Ad3Bc/gCCUQHbMc8c6n29xuiEekdM
mxwIR4Ob0koszUBZSO+KLY3GtopNNkcH06uNR6BuUdXPaqDkMJTOw5u4AZl/8vEuCw4IbTXJwbbE
l5d0slgeEBY298DuYyjsJ2qhwLUbuhJTiaJKtna7jCk51MNz5fdg/LOnlMLdVYe5MGKTOk3nfNj/
3nz5SOl9+gME/vUrUnmkoWyXeQOuqKuxfjvVqY+vE+9GGpkwSxpmzZurM2bWIt8D8l2ffqpFiWQD
R0wAHj/1cYeysYieMPsvdbY33RMx8mZ8O/ss9qei34clOuBiJhkKbzWUKXvyBPJdTvg3V5DwyFz5
1n4LSN2PydSOkzy0WffcNco69+hDwy/HJsfvYg7MKub+yobhx2iFZlOVT2ZZTeWlyoYWsSg88t0Z
PDj/UvDldscH4/JGSV62FHJ5UaoJo5ZI2IV3L3gMMtlSbo+G1D1fga1V+1CDyhDPJ2St1EG+p+Mc
b6uWryMlCX2OQpNWRX1GGvHn6s797HCsZvAYP8ORsMvrhT5b3x4fL6o01KyK5BMI9exKbd/tOPvy
ic/Dq78yvl5vPZHry5v4GqgpNNdHWJ80XC/ft/TABhWedtKFJ7zfEBRor0L4BdjKYaRsuG4jaICd
jGrUbB/6nMgooh4xHp/asPcV7mcFh8fZ/IrF7+xkwo60iDJ4YpBN10jCzbhwxjx2w3HYRRx7Kbug
85pPKe9yQ4BVhMvyT5WqA/mrbbpHSW0ABHmREkoIbel0hok2Uys9zeMtL39TIhaaIRcCv1b71Kxn
6Cp2m/c3Gins7eEMYn93tY+ZxinykREOQ1VogPe2ed7w7dXfiBB4dHTmlaQdRFlODTJmB2TNl8lI
TbGvyDsHcYtJzhCHzd1MqyRO2/0nDlqtEf2DEB3HfeLBoL6Hqfxz/PYAx5p8yxnqOlUMeaEdVsCV
OyFHuBTSNQnZEoWrP6d8IH7k34dp5/226XfkLEgP8GM+VMVN7FYGELnoU1kg6vVpdIsVzF9MsT6/
zWJJi+jTpbSKTBSyuhzenQjhOu4+Fl5N3TF9sLWppI21Nxu8SqD/QVh2bESuKqRc4DTbkIk8I0S7
IImruCuvBZYM271VLZqikqBKk4KQuJuzLKJ947lH94mHh5T/APn7+joZZ5cnJeKC+xPcKr66X7Ek
RNxS16KtN4loYuh5E3vtpU1IB7fXYOYQ2xSNqg2zemN+IYBK9Y7M6w+/E1wuQ8hWrz4la3LNoICP
XCHQ/RZ/DkWU1eviOy75Dpq8EnInDM4lrP1BU7muEc3KeIqee9AvzYVInQq0lXjIw2elrg7o+1Nn
OxqYLWbn80b+5Aw5/C5YHBt+Y1flsKQSqro0Gp9FVoIReZkyRq0P3WRIZh5v+OtQrr90tYkZY5Y9
VBUjjFMh9v9mLzY2XN00/RSEDNIot9f25Z2MONuAPyEkUJfbFOhVJvyRKA9Gbp24fS7iSulvAtkv
JzK9e6mGrYOYcpEok9R5BD8UFTRxQ20xz/LlhktBagm225RZj2sYklVgxVhxX5VxWfeZSYjtmPdW
Bs6CLT97ER8b+QF2CefFASt+RmlzoA754kgUA0DZnK8yBk2My1pdgaKzIbTW4b9MgkmGW1qUf7K+
PEPEEpmbec+9K+/wmjxwOkqb1XbDZJ+r74z3TQzErsa091or2yszbtyer0llbZvb/Rc2odBHlBuN
KPQVqFXZdhUg76zgNNHvB3ovmJBq7MbFKsY4usqUHlILpC8JjzVDpHmLLHQ+mIs5ngdpcLVBqAxf
xn+dBAecMHCA8Z1Dsl9jtjP0g1GTzGAvTpdREUV+V+HbYronRU57cnv4Q3RYridBu4fayUOcDzX2
U09+hx7466w8FoH9zOF/KyoRNjfSKKaPq4jpL0O2LBMBUs2CVeX7zas4BuoWaZt0BNzyplRtXTRR
KHTizboMPCFRVOV3wo07O+PHloJBQXWBX1aOPsqpTMP8LJGkVGjYpwe0Bl4qENubbZeEzgQgkS6j
LRnn2Z4DRneqfP9HZ2kOQVz8qTx2Ib6js9uCWb0ItFpfgERtUEjY7JYhH95zOt5WgXBp6BvV+vyR
hixTuL58GxOAF8+CJLPAUePXPVyi/0tCto9gW7HBWuuRcCCMA3qD5Zq0jWKiU5i7F+POIYBzLM3L
0H68Cs8VvFOrWwEqEuEDVRX9dA202AKxQ3HiYu3g+AKZqcTDG8A5WCqMxj7WqPjslZtqPnxc3tlG
K20ZC1EF+2U+/R2OuvIxIQ8wli18oXJ/hERRERlTqfoJxK8oEOaAeXzYZZuLTwhvnxCd52UK4HHV
CVMgpZzyEr7aqLO2q7A5d4UFjI4AkLbV9IXDkhoUtgtbd7EyEwLXa29TpkR53FFNVVXKAPTmbh1Z
nJmlcXWEKwJnlYDDRMMz5hZZfFOxhcXk6bb7Kq3lhlqV8JTtqFAW3tSaf3A/FdLhRm/dTLA2Ppgq
M42eUyGQ7rFcZ0TIQw3zDWFHdqag1A59TI5jxfh5OGzPYjncfK0awGjdjYMCPHjOfDmGRYmHriWN
idTs18ivv56VQb2Zbw/lTBlIpZCgDHW7wPIgLOTmW9+P0JHZEF5SxF+pyMKu93n0j3Ue7GregvWE
1ILVMnGVAZF0HK4G2t6E3jfxq/2tpzJfTFCxFH4dfb+2LWWl0LfYb1M7GZzf6b5b82QZ8G4ev6rW
Q2UDp77Inu1gNaeS0U8Eoh39xHGa3rBLiQyTdUDdKsVFen3Lfc2Z37X+V3fyRYYzu8rlWXQrzj8m
4PR4LyvWt7IOSVN6fAW1urE4mbhLIN81b0SnUnBMSgPOx2cDcjQQWghMq4HDsC0KmBx4f+TWodJE
uuSu1OaoBv0GqXS8QFDev43XmLxIS01hEYup87seQqV6NNl0r0drYdtInqVW/+Of9Uyq2RQaCwlT
RI+lyorOsF1DZ4fiagWDk6AHB5yszFAIfw1GNwD0SOxpNrg04pShN0Yt1P7UYvjLRWPn2WIB/0Tm
psww4DdhD+GvbNeTPPUsuIAF92N1+tnY+qd0PshZxxfHxSgUn+swp/LFUUNLAGPMh5H/MCTYEmJl
SkSLodBzqKxRCfSpjHC15SHSdyAiYVGe8Z+M/L/GAat/EU9sOWAaW1dW5qhlvF+nZxQcneJDuG6f
C7mMUd88lJ6hiPh8u99rNwqEN/h/bS6RTAV2qj+UpvjeadM29awSLqSu+7BCkM9rwKxtqCEIs+ei
O+ax+gFRB3tu9MuNyKdOvSVovCb4+YDi+6NhhZ4R+BHGbyiRzhKjmbH5Sq0pB290aTY154e3/QNY
HOn1UtcGQ/Mzw8CmFNobkCh7iRTMCUMspcWTz3B94qnk7qFAXHoG8gWYJdj65Wbxn0Ywc8kvZM2L
6T6G5Jhut6s+2+0n6KlH/ar9Tgtw/jmrpqyOXZD06gIJSkRNqh/WXvq+dOX33Ykd4kWigy0VMjIb
jxICVCSTPxp0OZInoPobvfFvJK3eBVygrRGkpB8B4uy/6+fxLJIh09uzTG1N8kO216LU2Tdi1x3k
SxtOYHOGPbw8RzGUo9t2SgDXkG4WFFcdsePxGQoOK9FncOnpwovFZqKc0YEV/GQa7tCJYk/Lbrmp
x+APiIKz1n9WF6JF/LOTJBPRerZNYk1z8nkfCj55UKNhpgXmA02fkBt7nLgLwRZ2B4Oq57Huwt5Q
nWSakznlPdUSmY+l+BdcD8UB5KN0Ftyv0OK0KyfGBEoDZ4ltNGNlMcjCmrwzHPJjFHAQutYw/6PS
sidrkBP2CIO698jdOdm71MZrfIKqLd+Hjh5W/1axtAMaWXBDjSF/0dO2lMG1aluTQfevDlgHf6Q+
4oIJCuPcUed/L1HmjJzqvRZxAqsj9TNKWNsZiQZHa7d1TfkT5ej4LOt1fZfUailE/ABhDdQLAOzt
KQBstMnfOoNZfdDI4fKdQ+nlbnPkjZS7wEQcDEHv831Oj21S0dZNn4CtZaME3iiftIodYIXWpMem
D/+7aN2kEsirgHWc0bkoNWX7FttI+fPTmHRVFZ2j9IHdVP0vg2UFq2UPChCG0XTCAi+e4cM4gvbn
HB0X4B6FV/izChtrSneVUisDd0oqYUtj7RqeEc5/j8zEmeFGm205MlRo0A1bkB5Xja7yqOcAZAYC
Iuf7lnJ9zxLp9aI+Mp+2xfMfGNe5axJDT8AG/pXauBf8aUfZXkDuXvsNYC+E8gy4cLW2ac6h0IDp
USnR94rDjvzFvw3auBwy3pQldbZ2lnMUZaqgNgbdcwkGTvphcMW4+ZYAG60/eESyArZxOICo+avi
wizgvIVFCPGO0PamlISX5ByLtLyoieKrRi9Mevevnbbc2B0ZWa/jRJAkk9/zkBSihP0LuN927PMx
H5C80I/9Ff2i3pMu7diUif1ersJQjeAfFtHffpQfMM0pImSuX+sAcfCpckFah8ltIWcABcYoLsXa
S6JRaFlY4PCU0/UexgONEDc8X1BFbDiIMkLnTOcWS2E4vonUDwUoYKcXARDdEzrS+7Ofu5yTB2Wc
KfT9eEMUmNWPFFSLrJ2IQi1tkVx0cByXMvwj9TxoMmRaJykkl7Upz6fhlFN0rR2E1bq3dCu/3eaz
b63r3OFeShD3oMymQXUbS64joC5yENor15Mq70RoqBR7AFIZyDGPBnWmu9pxQU2xcE4XKgzPCevT
fhZaf7o/SDoLqqKBs7a7lMQz9+p+6mzytURwHZIZawL3bg4z5KhUhUk3UtMKsiKjGsNS7FlxVrKs
Jdu2FPsbiQN+1Xg2jOQMS1y/Cgcvg2yrHbYb5clxsUH82IOofrlpDzUzLEY69j3N16j7xQtdy7E4
Uy6jI6a7U+qRhLWGPGfu2wcDycP3GKsp3huo08lAy/lCgxUt6fICxtyIwq6MnCeQtukxiFhiS7Ba
QYb+tdEkATK/aTPrqxpLRAIad9Qcz7Tmml7pC4/ply0b87wFNFCUvOkdj1TLkUm5qX3tJOue3wC3
89rULRtktoiDUbaMUqLkMo5d9gtCu0OzLHEaM4tTKbi99cQ2IgV444K4f5NP8xjY6YeIMPx03ieJ
Wrv9YG56aklxkvyuZ1REHcA2ivWI7qe+bJYmJJsetPgOZPJ41+bvhfnxQ7rjkc+fSY77Ie6bpcLq
V0fpjBwhKkouzYGcxF5wpUoHCcVka+40yz4CrIpVuzBAPND1GPl2wAoIyheeSjHdi9LvjmvVC4Iv
w/o9yDPU1tpZtdIlNwGZKvnoHE44fpfbCQftzeGSPHm1GytG2kzx1FPuod5dnZBvYqaOBGTR7IhG
62LoGD8vUl3abJZQ2YGDH9dZpQf+sqiCpKZD/K1I9dbIv3JiGILNhgiXwHA7nH1W/U6qw6pvE2Q7
KudSCf+uClK3urd7ezAKD8x6ZBOCAr8tlDH7QmhYbrXH/9Sk6jpv/pDSEmURHmwWOoy5oWp3HPE8
zFxQf638Mynx+jFOgcKIWcIoHhEKAdU9Dq+8kaDCZxaM8mKd+hSzDWEwAF8QWRPONsOBInMof8/z
oIusttpiwxUtEFoePlUCokqdJGUhsZoyloZZeIEiN+drX686ZT5WU/mShMt/MxkThAgr7OjbtOTd
KjQYFaH+LDjd5m3fuCmGLyFaqpFHDa12c5pNe8kcX3VT54n466wDlDBb+uW7BeVTNExjMZXG7Bc4
wHnbnfC04qo1xdeitlxlF1ZmVcLswaVOOddGWEa3rtRrP1X5JRnPKO2+fhVjjgRHe7eS0rkrJpMK
PGQVph8m3jnAl1OjhPCLaPbXKsbgouOnEqyhG+geq69/jHSvLTzhrCqRkR0fjmttMwyGuL/2vMd3
9K6kwb4wjtz/1VAGnaHiNmhPmSSTWzK77xCVtsId7P5fF/pdNlOB4OuoiMYVCuvpBrnUxfNFFJM2
xQa6IQ+A6wr9Nb39lZhUEco5gEC1AL3+vXlqResuUDjE5IF1H7tDgmwaz9T6ziWK5Ztn0yOs7qT6
APD4/hva/F9bkVbjuFgwFB4WaZXxU0HX0tF9eH3xe7S7gdz6mdp/If3rUOlllDXeucKqFaDHqr4Q
LTwUYGkYmIu4nt3xydIdFfAtrclx354ByVCkecIJOnLHvasIzOcn8dmRrGlKKishsxn5gQaoZTek
kiu61mm1bmSOO3VZWI886bftPHqGMDuEdVUUF5fMRkT0867DTjJ+KdK9sL7p3cnYx8fmAdlwnDb1
w5u77FMRmT3S+xqNo+CumzOMfnkiFH1K9TYNlmpQN9U/xFe56+lgyRW55EeehLb+9lzIt4wIgGei
V8P7bC9VktwCrZ97mNYq+axOfbF4hCptxgRLOEMwICSfnNzGpLUI0ETDv8nUbyc8VLmwsgVW5gaK
epA2W5Lov7SJD/CwJlFT+T6YSYmuEq1nz97CRSX/r2eqoWZDKTnd5uEL6Fmo1Myc8eKgUyGNb6XP
7q6RqDKNALIGGsbd3HzJcLFYtrRjgmVFZbdglqqmvQYK5RQhO1kM7o9HM+VLA4Vp64c1vM6p/+qk
HxDJANFcy75uDXA6Gsv/wnHXlotfypiqt70ZYdYLF5k/7fIPB1nMqepKO5O4FmhH5hBGf16iCWA9
UbxvWP484+PqA2IqXCtV6qLOu16wkc8hOaql4GyA2CKzDzJYglAlHr+DAj3hV5d+AwWpTW9gUssX
/O9eY9B/y7kz2ZQdEGcxCUim3cMlJCg2J/dEUqprCkA2ffHqdi5Xn99gS+tKA+EW3+7FG8ooaU0k
T2LwaP2HXpc5APpLTPtmmuj4fpNV2XC95cx4U2hPSVDcS4ESyDi+af51kgAS8ecYUdAbZUXeGrmq
8iE2wulELtDzr77GYtwHxr6uBIw33fzTESJx1uht2TpeqLwP2h/EVcH2fNjrSCztZ9VXeTJgVenn
F4Q2XsRzFfhD8q/WeowvHXTIe5zyC1hHjaTs5Np7w4WC0FOa63cTHiznAzljWhgFQeNsDpdAs7Aj
JfbFGLfuTpfWviEx6R7a0D9XrggYGKJgP6SnOU9L6Bb4gU+rG4B+h6djLwXi8mvpmERwjNPgjhXs
WFqxFyFx4VtMdp4CxILUzNQz0Zbhn9GxPksxP+9C+35EphPQGn+fORFwWhWNsR5qLoS0vWOuhdnG
xcpoZ8sbgYPECRaHLJZR5V9HywXgvsg1sDv8FvxaoxD6fbPK/7iKgXyYuH07XfydWYVmEBPzMGOY
AvEvGDHnnJzeig4lvIkWC+Zk3zARCL9s+XG4chlJGTivOze5h5KBS6hpXwX0QgVZTg0i4ikv4tFg
crTqkAULG38arWd35POnGxsy5oN7GyQlgbtvXEFdjAC+eK9nzPgb5ibw8VigWkEp6VGPQFiucr6R
w9DenAsbn8bhsnnWSKDoOACG4+wGgAXt587SCD1+h5m+R/9gB4lm99ME3cq8mVFsHXBxD/Ys+0eK
WQXuWGbTW6+Q1LPPp4pXItLVRWROQzevRwX94gl1oSYkZjs+8Yf8cBP1LLQIrFFFAS0nswvnjaG+
PBQ7zh4iTv3dQxUzYjrQVQEv0oYwppjFMFLyCFOA+uT84gS0mcZCE1Nyw5gP5O/waH8Q3CVxzzYz
amr6Kbal2Toh5ptAv7OWtAGN1wXoc7rQAGF16PKM0+lKPYkiC4QljGu8WkzLdY/3q18NxVZy1ruz
TlV5ziWIF3TFNZTFcxcaoIKiR7u9NE+d2+Jyrv9QIEJ74kudM3mBoBRPrtci84lGKgolZnaq97Di
Hkd8LNsOPbQJN/zQpxxJSDjAAABQRdyvwC7MTcXoQTrM1iUcpy/bx1bZx3M/7DDTh7ZGMfnrf+Jx
OONRxkIBVhY5+cbNMPArktxSAUtNdhHJfaXoWZfwv9H94WhzES1POwlsEDnlGhiq5ebnITkXdDVn
dNwQtQdTTt8amA4YO11zAQmflHu4+BSZziXnEfpBPykroexkHbTEyt4r1giaZlle5MQmU43300Qt
GpD4PwR6TjNluNv1+UFB08cH7hgjesyX3tVlJwbUi3PEogJ/PysWfs9W+xKz32p2tnO76nRxaqly
1ShZhdPEJgdhs945eKDdHcrmKSC8fbf3Ke1F29OeeY+0FW+Q+Ix0bulmLqmadm7uBL+LEDBOc56k
VQziyiheXlpEwh2z5fkL8w00ij2n71CnDdgf/lWKEj6xBXNPtFHcgyxB3C6kZgHAA9gbz4GEDdQf
Nv3Z8I2OCJS6ZAH2NfCEpu23qWNaSm52ex1/D7F5L211jnuuXkBW+ZCHxaoXYdCMpoZ7EN5zElgE
8TZssj7Y6u8E/kbGcEkDuqlyCDPDzdAkVIJNsmXuTdbosTz/BjSZtFLhCu3XArFrd/1uNe+QlZi0
+MDoLmtc79VPA1LE/I/VGPxLFg8pCB9WJFqkCNnES15nJdB6ZS/cODkg25J7nWAsQfkiLtU4EkSY
2mm8rEXFoRV34mqZ8XJaginYsMhmU20CxsK4IybJFPP3vKI0+KHotUH5Yh99dealpU+LieVuhk0w
+s44gNueLCHP2tEuexk1KvaIC16C8hPyStmKHkbi2al9DwK1Jnoq7jch9U84flACqVLICTzWN5Ws
C1si/zOWofwTRQ+U7tZ+swDHXD4jfhj9LBJgbfxV3Tdgvqf5NCZwmif+EwN1uouWVKC0q+B5odZk
WlUx7WTewn+bU/Ydv7cZOdV5Gi+pDrNd9WvzyOomb3HdSGiICzuDttAUAOSjKDc7JOLa8qv0ihJq
ZX8NgGdrZ2rT5WqAo4WvZCcUWjuqyFZG8UyhNDYSLZUncX4FSWkYwzQMPVbotExq4DS4q8k+mIE9
TlUgXRLXnEagY6JKvqSQYJtoWvmZ6Gaw1jruP+XPos7SY0Fbo9GWWCWavB0mV9CmqxaYDnl/I42Q
xYOrYjgXqQLPuCTkZrur4Ew6lZGstOdN6TeiM31AXBZM07Esl9QB3r4FUWALuCHy9Cibs8+/wdD+
bgLEuIUO4MjYi28SbQw6OG71+nMJDLivmlAst/FYyWau0KXpKSUyX1+goJB+08vsfCW+q42swlfb
Fk8JyrZPqR/gKuGCvnGeHeCGPw91RJAOF8OBKCrQDOQ0kEBdDulKR7ZYKN2Vbn59TzdnLGYNMwSQ
B8EWP2BiVLoKvSCOYqFIYj11hHYP8B0xeqfHwwXLXs2OCVt2SvEjGGPxjECY7rvofKTmeXHwiyhs
Nfzaf33DXON4vPNTd8ZCzqXS4eFpQQNP+8Za2iQPtf+HoUDLV5NKeOWKoV3omi6cPmTAd5R0bmXk
mFgvAOqAIIv1jaddv7q25lVsDMl9Ri5JSQ5LPeiXLz2RXGX6D0h1ICvWeg52HC8VGGW0QaLHuov0
+tW92gDWVa+fRU1S+NeQfz9o6XntapJXQY5GcqmSJS7K82bPkHjTJhRq5ng1qBn9+hQQnTpCjFfc
kK4ukzBXPRtEnG+eq9pDyx5II6HrJeNoAV3b6qRIkzwoLtFo4C0RPuyWzw2j+trhSqxkbsDPIPPt
A9DPv6SLAX6HLjZKNqDsZivMNli9bw4M7HXudnXv9smmSzaG9stzzKxp0Ip4z9QacgJCIWZnynSk
HFSJVxfz7vU36GksGkc9qxypb7S0sYS0eft9QsOns/zUfEqdTA9YkuW+tRXClJiLIATDTIu9UiZu
c3TitQPA/7Jb/Vg+QjKHP/9fccKUV9C7JynkdAVXAMY4P/DihS93ivNSKtozcGt4Tu0kEtU5IcOo
YghOOZoZBNlSZT+oQ2arzMvaR5zi6V3skOAJGY6CvILdAXhYkjxmWizc1n+fvzKLUE33J2bilTOC
EO8jYlM4QSMEcZzOXBqeXwrAGK+xwTX4FSfBCSuAo8Bh3D2WKzxyTCbIQgwcvA7jZtujJwbvb5is
2e7wQdid1xxA1XCGvyTHLPjiv5LcNw2f7EkVOWl8Dc96/cKvP9IbipD9wgbpAWJxLYVMlZt56BtS
gJNZyZXnN/rPcdGj7MNJiBWP6r8SYknz8IbAgVC6xBgIM67qkJqE5YnWaf85ss/S2hBj2in6+1Fo
GuMtFHIBpJrXNHcXEYUOkDHQTupkCgVyEGr1DZudGCggu/QNpWirlXUeaRE4Rg//bC6IeXenLFoG
SLC8a0FH23RWJZo=
`protect end_protected
