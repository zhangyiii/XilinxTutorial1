`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20960)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAOTAApZ5P5hFPOW7R3HyZw9qgz7rbWscdzh2IReCRHnqRyGpinv9BHxp
0RKvsPaf8Nr9cs+tVk4pMfAQebpLNyPF2DKF+szcqd8jNuQ0BwD1uFwy1IFnuF/W4/LUAcGR+/yz
tblfWeaSdWWNWoDspkmWOnIb8uncPmtc3HNtcGdEeaLcCV5hOD3UakMxgPxVxH+G5zyNr2NiyzGh
Zkl+YmpzJmU6GmZV7j7dPExWDvbbpLjK4WXnXDhhxYgRU0H6fVbry42tU3/AKinlgvrmIFbpZAUW
XacEL9dbDEuhBjZRR8f02ET+cY+bXqcmv+b+T84PbxWFOGQx8obwhTOkKUpVloyIFsqYz4rEzSC9
4ZBdbkN/YFgyJBTxNqOcxOJ9qTJbCOZJ5IcpirtDLf1vB+Ad8Fldp7ukbBsGSUZqZ+vuQbr0NZ+m
rQhFmPbSGTG3mf91AuKMUBzrsCJSJohNBwMBHeTm3ekYq/N/3VLcfFVvmciZZDohm3Nkn1IKCftS
J6z0fItpN3OLW+2qRfDS0tC4FqoWMquYnQx7LaRtxxLX2jYfdhL7CBS+vQn3IaGLo65oZnh3k9TZ
Tip7vExS6wt0WJX325uM2egO/EimwS+spoyR6hbpuE1nhdzyj6WU2dv+uYxEwFRjIpzmhq/3n22E
9oFoFEeqQ8JDwqA1nOHAr8+SsWmO8MVwx/vFZqOqIBAt4ml0PaiziPqKTQvR/mQX43viLNNnWjk+
JLA2GL776QOZje2mC/8aunjF9pqzFOwPqQvsEvobF+fOh2tKfKHTDUvcqoJaicA469JYKfQRc3Zu
1IP4L4JZDCx26ayv76agBZ1D8jq7BFbS6NKrMt+somcwPTvQf2JtfcyiICYIrKMppJQArt3+Jgs8
424oQrBROBTKfbNcmE+l/SEOB5YcKt+e50F0t5G/zxCOr37WgYfnIKbCtFNRaSZ9rwHMNkcq7hRZ
GCkyOzhcIRXasrPjOnP1xEIqRCZchLjvgzljEd7NONUWcjB8nmSuizfy0mezuNWgE/NkR9sEYmDf
WVNPTAlQzXtuK9rr9iPt8MUNLgZZMW5ooTm7RoLksV5d1xg0NljSPoxXafNmqU4mh6l+y/0razqC
Ib+K6A2VvqiPTstsLzmJ3dvz6zGdhq3ssRkqp6PtIXPHc+iXoAnkwnzJRWaR58SxIWvQWXDuphUv
JvAZDW6BuYAYdxldecusEjv2t9Uwnl2SMhBti5AuJhgUKeL0jjosUzj4+E0ctJRuN/zzw3X0EwLg
90gev/OA2mCA+0JMVA34CYf7rp4mJ5+U58/1lCCSWfPSgF4mPt0Rh/bxa1ANkBMMLkMw4WSPRFRU
HruGM3QCXya+Hths2oSd9bxkWMt8tVVwKDMgNEsuB+CMmwkBrlfMhaMVq7cLFe+SBrGUjsRQbSJV
98Z+hzR7YMZ4eWZ8znf+NF91OFdIacf78ve4bmoC7VfhvJ2GahMWtJsVl/XDWZUI17wRscIRvarO
AipqdDq4yI67dA3mnG1BAnJKViME1yBIEin8lOXXCiFkNBbVpo14b2VNgDFqMf5ssFYI1l7qz12J
0aE/Fa4+/OFaLaSgmxUGG836JeiCjNNV/tacViHbvDM7ZIk1cuFEU1SSWDLB8CCZTHZqGpuP+TFX
lXz1jCMOQYW9lnTO5kRPlDO+fSSImE9jR/qYoWN2T8tgTT7MjmNSM10WxOYsZ2N91ejJGEe5AW53
8DD2SMfnOCKX8DLlSRbPLKNyarMZtJPxc7GmO5cW189HsF+ETf4FpkL6KlDe3+b4FJH8uTV6cCrf
wlSKRQVgDRumG6jFCXwD44i+SCAxj9HSxNqrIC/AniqUOAj5ZcNBstF4IaCt9JrFb2PBh3VNDvql
n96l7PgOp9LsvjoPvpxOcFPW/LfoF9brgHVISvG4OR4uyq274qqxB6jlLPYZd2XlxtYEwRRVmdxN
zOoCIqq68PVSUYlNMhlOar2IQNwJv8JMb/EMfL571AzV1GP3XBEatwa6tSMoZWri6dtu2xOzv1Na
601l+ufi5UUSyQ27D5mjWtURM5whfMEFbHRUtrCma8rCVjzrFc1OlvL7/7/srLGMDiE0wiOTEbtu
pcg9eKSBnekTXdHa8/bsNo1hnCNSy5SJYc2HCMsWDO7D5pqPxz/m4gKtyi1i8qV53mo2UyKTndQH
DoIyVFQ6cKkeAHjHsSuAooMDPLL/kPqSZRBwf7ReF4oWxGo6Ocwz5gMpOJ+Ay+7r5yLskQEAWm5p
QluVRl0eJyf2E+64kkEfKLz7wbKJFCFjqpz3JzTBP87dA1RR/x8eM5FNFF5CHjB+NUPY5Bq9mgq6
w8UnZ3WdTWFwn7FCzT18O+HZ1Fej50MRk78lMgNN1lfEIqORi73iALiJ5bJQOf7oWTzH4BcMUQew
d8nZGDhixDAmYJW5c2pbEq5r38bDAT9txJ/HAHqAFPTg6iItqlo14HE7ig5oh+f5svz98Lhev49K
9FjGp+87rhHFZlsEUMe02sXPkMf78Eontvao9ONqIkTaoF5nqfmg3pBp3K4ZpgN6D+6ZKFzPslKU
ZBS6DMukK0I0ErDB+TJpr4j5446kg8+itc4IHod6Cl1DsgvQp7PVlaZq37oSkqDVchaNlxsuGf8B
G+ixevCiY5MFYHUn4TLTbTqKkQOoSOKIDHuhN+angSBI/UCcXt3s8qgIjwVt9In84hK19c//4Shp
EaflOYZeQLVJni/XqKT00FlSpKr3R6TcT7V0a8IDS0Mzt7Jxjmy7rs8pyT0n7Y8FXiAfu5A4IG7c
wjX0tYp8PPqNpWHiWV6OKdxJLd8iOQ/jqhqiqsAHIVziIHVKc40bgN91jhf/Jwak7pUeThtOInSX
aeTiGIn1ELusGuFp48jzB6Z8b6QkUMWVYda2GHZXHIwJ1m7PMyzx/Fhrv73RuUHR6PdyPWiS/22W
u0ToqhUawKJiZssJJRW8GsfnaWnkgc3jirOorLTx9aj7FlhIKeJuL5seOxXAUoKV6RVZUUVkejUQ
HVJfGLRKHfB4coSRK9pafxQIwiSENU9f4fKVR1EwWVvCVH0MPc9HY3b55d7Lg3v2BNZ+n/TdJn/C
rUZRyhe3f+7IsBu+iy92KH+yV5my52glBhP0FB6kdLw4aK02V14OFac9yewyX7a9t44vhh8xgsSE
aPWiX0UdVkcn7Ca5AE0abwDta+YC4Z3SjttVd3TRZM1d8xijLEDVZ1OzlFjJI0T9kfvVHuovspbp
NQYHpptr8X4vtuFJ67FQjcf8c6OzHxJfbTOUw3AMFXDNb+nnegNYNF/G0FgzkMBLQJ1q6Q7XNWFD
tJmc6NLc2Cli9tVwEkXdKqjG6Hpd6eihULGdEehFsHUKQ3LNfxw/aAmX+LWhFRQdWBmL+iavo7Cz
KYSO37ZAhjBKn2+bhyjxsWoHHKgn+OQ8pBVPTSkSocNXRRgruQzdtcI9wk2x2lipgDd5qf8rKDXN
LmPQh386XoDBx3e9znOZdQwYV++1A4yrk1p/94/xE2bqkuMzqsc1VlsVUzh1Y49Rqjmd3y5CTSVI
aWuotzPe6IBiTjzvM6Q/gS5zxRruILn9HdfMsH76J04pnL0NRf668JvRu3xVS6RAVy1ZiPYF5067
tZC075loSBc+m3akJ5grO8Upy6atUS5asiWSDy8oMawakn0diH7Svqvel04o158SngaWZjma1C8n
T3wXqtsQu5so9mMxYyN6wUkUBpQf3iHlce7PDKhWdOkMbyDtlYlNAdfGiMZWX/Z5EERvWn2KGGjc
VE1lcYu1B03DkIpeKX3dpNwphyyiQjXjRNYLZNFx6mwBD7lMypFRerY8pEgKtu/s8th8mHkNZgyA
rOR/ZNzT9FyOE+MPcSSUUGQzVrg5twnpcGPgzsjL51nkIpawsKUi8G2EFUohA2DZorFn/eDAX7G8
ULxpReiKNMmfVwEM7IT7BxM2UYa7quqNNpOupM0lljUUV/qqQq2V5RHOEKEetSKlNEc8GkqnAdEf
m9w1tF/avtAimbcOBCJRgdeHIRu5x33IktP6NnVw7+jZP7iYK2pZomUjvpI/ZKDG+dYPeeD2eLKl
pgQbYs0XCePNlSf2xr5w73bGqhsUKrlYxXwaDm8pe+OnLXftUS7OXT2dL/MgX3Q6DcfdgzRaxnzY
cR7RsG5aXSx5kHsVENq2cF7y7cnEKJHAQVRRzKVf4ZtcqFtzupiDb9EkpEbESBSLVZrpiYWxeE54
R5u/ro5Dd+S/+OwYQQ+tTs6HVvwPoO1yRRcGHM4kJCvswyvY3IP6gDlch0jgCd8LvQIENGtXVa/M
XXDVhW9nl52qVhRWG6zIRhm4u6+g+XDEWCa9TpjzaxfxpiSUfAVnuQkSUV77OGabIAlBu9k2oyxc
zvrnmQ53M/jU/tmFi/32sWBUOeE0IGNaquY+yZWLoUm82XUt5vt3E9ahZ7g7gLqIg6OQLBgYc9J+
AaBLkqoF5+UrpAb1c5FUYauoWuXhHiSiN/Cie/KZduIngceUWHcL6/1ztKnAsfVlEcgR0dYKQv/t
OIxpltspRbvRHDDYksRhx8D8/mG1OVzq+z+2VmtyYnCLlY6jUN8VPScmI7DrOYb1ScdF3TKtq//1
WZi7zCUQx+YhvoEqwNTi3h8MnwtrAkLX+9bcPGnrdUvqtTuTmCjmbFpU1cOlU2auK9pXhsLmA8W+
tDW5yoPuPOfa4nFfFyIZ+kPEUTVmbS5sQN+JxICYVvb6tI/9php0+6eDJYq0ej9mRmss1fPEeJIf
qcttoz0xZMS+8sv/gQxtb+EqyiziPiq+1qcmg5CA/uTkeyE36578O3v3032KuILiJ3zSjvCp9vKC
fI/pI6YC9vmAGdRpoCKKomHEeZplM2EKgIYT7IrKKZ2rU5DyCqrXxovk1mGcktW5vvASquHF6Um/
pG26g5I7MRt0dioz0zMQAy05tU4Olz9zzqXvGu3Pemd7z5rKi5AJW0NPr5DwGMT3Gc6nQXHIdWvJ
KuhoY7C7veUedAvrFeSnw7Tbc0/zqSg2eos1t25iC3pETQdSi1qYsFddX1wkBQ/yBnH/KL/WMQZU
Xg0HlOVoISxCqlzMYabU8VDZOzSR0Wi+GmB3LmF8Ys61lMignfTsyPLtHei8/KbW0VtDgXXzpJCM
9ZyylZe/B5QTbKpzLyS7uAxgiG16JNJb55K5RFxBtt8U9hxKGx8mk4gg77yf9LPz5GO4EKqXT6Cj
MNxECNeqEcUevhIWEA0dNU+lh8t81Wsh3WC9+SMvMfOuduUkAtui/VEu+1FGRJ5qbc6h+M73JOKf
AxWJDwZel31/Ly+Go5JBCTsMTK5o7pL3ARGWn/qggCfBiu25cRuCQRRl+3PfLOSic00cVaUNIY6C
UbW3+tlOT9mvnKQgupI+JIosHzX2W3dQJIxIe8Rrm7FZsB5S0BvvZbCtmuI92VBnqodF8o9XyqBK
UAd2Q0tFZ4kA3u7QDKq9LyQgyfDi9a+xV8nJTBPqflpjv/CfIHLa+HGa2gFV6vZDv69qp21E8hyQ
xJdIwxLHpZzFxSD5tUXPlrIm0HRc4HJsrx1p69ts1kYosMCccr0pHofflAOwrjq1QCQqU+KqpL4e
Y7t6BsVF64/wpWJYRRZfj7zZZrWwJIDHoM8JdOwyYbphq2bYqR4Fr3Bp3aGvgg/NOrUOO1HNHXmZ
w7kks4nXwnJvH98ZIqYyom0d/MGBD6qiMTjjgkRBjbr4TBC9viGLSNig9MvD/C+gqsFV8G356J1r
1gLOpCOxuAo8mGPItgpea07fH7XCLA/wdH+KTHtffsCeuadfWSGytD4fJ4rMh5ioZtpgd9tj3urC
i+093Rk6EwtY+5M38Myjz7qjCG5UbjHKvCpZbb1UD/kcWODoaRdsJXk3AJpiuvUFfukHUce5p5qR
MJdDz5EpfUDdg2aTG4pg6cub4SX0ajyhv7pF4W2MJegvIcFtJrjmzusTvBIWJJ93lmRyWzf8en5/
TWUJ/+BfaiL9CZ/Yo+i4+P24HLH5L+2p3Vjt09y7t9vbL6SoL8zZC6RCgx68WwifnsduYbgOUhqM
eZnCbjqZJeFSlReD5z+BpnpK8ufzdc4ngwekJD8Q/UrgaDK0CpCnMsj1M2epn/k/OXFc8o30Aewi
o701ZZs+MfnFys7oOESTk4BKylaTD/9AGF+6gcU+gixmBjtF8nr4CPBmPn7CJ0seQb33wLxd5Pim
eLliq2ITvdDY9+Y9mR3Nj/6coaApKwjI+kaiJ4yvwpFnvVuXgD9d3vX/bSLcfbfxJZN8u6Gb3r60
0815w1VLakyoBJz3zC4v1TKhQZHn41xV/PhikmMvgM/YvkiuZgiYbPG2SE9913qKHmRLBRGGC+Vv
xutddAfdUwToxYdQQsvae5xIp3GasrzTOV2eBN534dv5ecIW6wBHK3ov9zmFpyMLIzaTQhSLP/kA
DiOy5wnBPpUrW5XUnDXUcu5tfqATtGSo5f4i6GkCFUq2k+qwmIALH3gJTI7vqkG7EhRWUprFZXhh
k5HSWWdoalbuzVnfP1R99nisRKSBnmYIT5CguetMIIdrq4FtxgZT0pWWzkJJl8rdW1QV6HZo1lWm
EkQFT4DVxGtc7sayJUpQv9yFbCO3amnlm5eY8OgCh1zAxNU0xZ5kXh7mWmPqOhbgxYkMcTx3QhlW
oAm/aCFkKV8go+sj8TTXhQ/UFs0db3guv4M4CPMI7rdDxn4yF93mjdPYlMUsGdWdnaYCxvFhgJaH
3E3HZbfBTA0vTDcksmysLwzNKqiWAW3rZpxySp3IZ+FpO8IYOnug/EpUt9HU5Sdc62qx7pbODQV+
Z4hJ0wkZlaLGaZ9Bp5FFSWHez0rxcih6GPngwCvSR7x445ynU7wkqjpe6cSh2sRiihtMZmCEZ8Hh
a6w0pI9gtwrEzn5UrA34wYEuZxWPDjDDTzLEmaii/BHLkSApMa9QjWHT6SF4Vq6yoXpjeO8Rvrk9
0JhLK+4g/7UPrKkoheRzCWIGgGtxZ96T5Z7Qp2cZ34jYKBcdf4lhMjsCEYkF5qs8PVYPEGj5QNIQ
F5+2IA2ts09t1mvszDIV11aGVStBu5rI0fd/lpYW0k2VvrBo2DVm+ekIy03ux6YpDeRdVUrfa9NC
qNFW9ODFqfZqPNUYfVkoSuUCzSrR82SS7LoV7oh2leBVAHDYKBfUOL6OMJfqmR2o7s+uPzCjx9Pr
si/XKreu4O34qftXjm62fyXeOmjXx9hy2PgQ0t8LTXN/eDDCYHeAuKurwm5cW2XN4ETiti3xkDc7
uSqyqnxtCoWHAc+CkpNplIqO9u2MONsAyDv8DQut+6hF1U27psmHfRla4gZEMK4334/Nc1h+nPjj
AaDu5BuE7KbV1iIOoxoIPxZei+GIbK/kfRXGF+v1bbYXJe5jHwgl6AOyKpSeLlO3TtPSgupGVJOC
gKmrNpJctnisFaLRrAot1Jwn/iYQsZ29E4QQqovsMwRzPhuHZ7aUf0YBcSX17vM3bUymZgmQs327
k/DphE7F1s/bEfrJdoxyMNTTTSIQ4h4F1pC91DBgEisORHWrwcXfY1RcNdemwB8U4putvokbnJ3P
zkcREqeYJPlvdty8VvARforEdX25+1jM6UboRSd8VjQCZU7Bvzzwl+ylud9DS7l5NvtsoX2oqLKU
1buPr9ivvxQsUhq2m5JnRIyhQ+Jf/lUsO3ZUY7m5KFe8VHORJcf6joNtyYLJ6WLooAKLAelRS7Bv
laZRg7NtvZbdriPe9wz4ax5C2peBWuFmS/eGR+MqltIlJFeBxO7l/9rDXZ0YWgKttWc2Xv8wqtfd
XCegwcEsBNGTFqusO0SiBBtQ1NOFtgnHXBHZPELQOsnm0/2wQJ5cfE5VuHkXVcRGgnNne4AqThi3
A3/7SU411fpIUHxFyoGy9qyPPwS0WbsRT47n9WGXmEPZPh9XHSpbsct76za66+PSBmhN8OexR/lC
qNWbicTvSNj9JNL6CGAgJ8SNT7M4p0qOxew//LDH4JBXOYXkdYCoFsYtYu583fX10PPBVo6Gh34r
TpNdKCGZY08ENuM3yeadkI2gvjjMygOmlzel40TNJnYAFucC+2vPBHDEF2RcbFXbn1Sv+u3kF0QU
CUD9k0G3C5fXg93PS0UfYQFkLRyFiIh6QBU541Lm/fSJb+PhBzhCtR02PMo69VWfl4PRYIPW+S7u
L9p0XeV112GiMmvuiql0/6GZCcnXeWaePKop0XzYusETmX4112mKvghnf0U0Kr+CJSJTqI/rz+XE
rdjdIKcymKGuy4l0kZOg3owpLXrZFKlkhBsHcXwJh74nAtqLLIGzKhc458Y7Hkr3ZrkfJAQvKkmy
qJQF/6Jjg7cVgbGPqyqrIyHIE71Oe8XaxvZCZ5koScPdbGiae4IlbQrqSCP/HJDUtkE5qY5zSh8G
5tauDa063kY7+N6OVq0pQjQyNvjePcGljeoZYXhKmcbo7bSNYHxUEQs0e/ngTDZfFdN0OIGP2+rB
uoY8VbLl3tUutvg7P4Mqu673O0k6blep6mMC+xBfYOX5QI9ER6mzrJJMybHaQnnIKucFcc/csXKP
2DF+whWvavncxjWYaejjkudGu9wn5DPyAE+KWuiry2xcWkNxF2PP595SP/SdkO9uwZDDkhGCRDi3
dF11p7FHYfJ7CXVBJhtTLxZnGVm64s6sJygwQxd04O6QguNKVedmaQNg3247jks65zA+Msd7Cz0J
C+Zk2xrhPGqCEnP8w0TxwbMSHXZFusfAol9riSmUFMxhw7eDdRiEttqrPoL/nL+QsrMG9X16uzIZ
UWFhmqQ8B4AsYDGIiKFpf97t/9FFjlIROTBvn/ZTKN5mWEVuIZIQb5EO6u9n9PenrTPRUEyfk0DS
olQ/iAON7gEW126jaz+h9xC4gvIop8TV0njsCJA1x0ysQllqjbvwLgjfyL4alvK3TmGSZ3WpeuWF
CMJqa3fQBffWpLHt5jgW0m7OmE6rnec3v/O3Kx/NF1SoDkPeL30Adw7rrgVzuc2TKJOD6oRkRKRk
wrx5VimWHuAIV8+AvKDADKycfrqg0L80CoXdPmqoXSM6rTne/I1ECTKZKru4DVm5TQ+JkdGy77j3
fT94R+YPjVOFvi1pxXp+p0xPzMp1lavVVwmlgcS60COXIu9dwDr8tdkl+qJwdCXEuC3lwt/g0ACF
arYsk/JoBrzfXcEovUWvTJTMI8gpvl7zEOzPLgE6Km8MCg2dB5Axxpl5ykiQZyzFlht0lsPvc50u
Jvn3VWqtDPvUIt++SM96PDLivt1pCw4smShrEBMQsf/xRhViNewrwubnETPDR4C/7wvd2/1RvJlj
SqkbKx2Aj0h+Nb7QRvTAHD7V4H7gcxsfo/uJST47Is0O0wwquVNDQffz4oeE2VFs3r6D9Jlak4Gc
KeETVDJVqeEnUowntn/lt28vkMlKrgmX4bvVx0iwA+ZOJwVRW39nH057lFHAnenJyu68KnZA66gL
HsFaml78afTQHzBKkuGp0roNTfivQR0RgmRcePQHdsDN/vWvQCNpRjEh9djYC4GeYR1UHjOBLDMx
kCo84xG174yOWgc834FaxMerWXB+cAjY8+JJVMn4HOkPasMIUesS+pdRxDgM1ayfK56NJO30sK1o
sb9AMGLSrIJAoGLFJssWDj45u/fNOQy6H8XwSCjgqTGIEVO1qwKUARULpglmooccEfdkK89P5aRi
0a/iy2zghhXs8Jl9CWJDrZpRoi1MD24UdeELYgMB+tQbUUZgM5lZYfIyyfXvOk6qGtp+j75kJc7l
2VBS3gtNpn6Xdm+QubhNXA0Y9W8bQUWqBO7ANlTxbG5EqY0FUNEf7VsnNIGpTJGjQLcZiCE5DCLe
cpW6nOvdztCiu1ZjL6utA+aHxigP5c/yAc1GOmS5STZQtvBGipQLOhh023GFQmKOES4bWfcao2nD
40sS6GLQ6Cp9JZgFUYXWHB15Dr5iSLUx/qsyhnSU33uestLB3VNPKSv7ra5RgucWCeCiF9J7ii3G
1A+86NqH51KzakMIsAUVlaoujTkye8/EqgUPc/gEK/lNiSEb/DwKp4gmupdcQmQb4gqXZeqVyeD5
i890UIVI8QsEHb9F+Rkbm/I1Hpjc0fphsAQES4IUrUCnuXsSBwd6AQFJbCLX79zopIdA6EQZsFDy
pu1c26+vYhxwaaItfESftGhYeb9z5WQ2NgCTAg67H9EabBqvmbMsnH43smXBdBJAhsVaaxwVBtoF
N/vaPMw0Pgt1T3b1Ujb8OdjO9SGdE/dgpcYsPpcAYRbxIyRBIogQWwJQbpUTnyGQo11wvTwmN3De
EXdgt85J0IEtyBGuYlKJGS08K7jplH0bXlXuDa+VptTu9iNfIewrA8IaFYjFYQ7Dr71GVdgnQ13C
PJfbKedbyH5MNPyBmR97V/5kjpjOAq4PokTu2Zg0x37/QHjYtqM21GvUT9aP4k8TrjuwY72j8nFZ
kKBh5XWX+ShEJXgt1t+zNFCa8wbPRXUMKPTOAt5RiZjzuzQYGWcMYPtg5NJov41iIZVZ4TvSpJSb
VUIEb+DgltzB543uOVSh0sMx3P5+OKKDMxxoFEpQiNkLHjyYZ9mzKZi0xJqtr5119uhwO7Cw+BGK
jeI0jaTxUXvKO9SHKKZzp6wcDzW+JBtkItTEGk4dcrByoh+zOeHyeyy3gRnnZzzxfMPPJCajUNSm
rQrzngbHNZ3iYiQRZj6dFnkQEiL/PlSm2tD914KAf1s0BuE+Lkq7Po78lU355XyO3H+eSH0KlvNM
dllMy54tKwal6DMsoRTNIE7uTtoNP1E575DfvBX301fFbygVgFvUUHgV3v2vA9ziLTF72WnfiNN1
rJDe5rlFmK8oWXImgWOunxdYLXyljph0yoOasBc3zXEjPS0mcNulmr5N+u4vEpGWnOrxQB1KNGyA
7I/Fo06SmuB+j2lhFwx/5OHlVy0xxorQ9EanSS8xIj8zJ6/2Tn5basblydJoPqHlECqUPP/e48Pr
y+wQOTYP7/robexrHQowLNUAhwkqZweKJBkWL7YXOtnTmQgry4NAKt5DkjmmiQ+Y3D6aATn8xcSE
xlwj0qpg85havBhDCglhUQrrMRdwnxbMXntOgp+eHOVdrP5fEbS21REFv87qn8dYataRQKTCKNdy
5OVMceMTAxDNCS2DM4r5lqELSqL9BadutFblmp281qKur6RB0pmU8XhnSxUxxAtSqmr6BsJps5Ae
cZP58oGKO+fT/J51O+B++fj9+A/ao5bcBQr/UaBo9nLYJ4HmNJredDUqAfQp+L+8YKSG2jD2DEUq
fJu9QeJFn5REVMEtygcKXcpOcJDn/rRKfxb/dI8tmV82IOvBy0EbedPPxIvaMVZn0a75Wmxzo73R
RKTmhEG5bTC4BsnoR4Im/Q5weK2OUylXCMxO4+XHqYhBnUodSWFxy6zSy2QS6Q0D50CWBxm1LbzZ
Rh3RnfjvTL48QuswfakOF0zQQJohUXL2gz6waWHaJyBzuuDz/PTs2htwuRBIm2zH6xHnKEiGZbVN
FPKqtYZcvGC7hQM/rxrpQV7ViRYmBmRFa5J5h2mYdVPhvotQ5LTtsD9Pny/6WpaI1VjFU9TUK7Pk
9tAsT7dPiusdprOGk54mXqOBTaOuns504ihe5/mbMOaMOz8YAGMLVU46pr9PVQuVWSYa4qONu9hg
zs3lbxzGCR6wA4QlntM2hxOZEIZporWFa0GgJM0tBNC1BFzDw2FOtWkh17kh5ebBUwEodrqFSeyB
4ObxEDsgihOLIkM+EomvQpjUAV2EJb47rWxYDVXZ1l/1xXERK+lw0XCDsYZ4RgfeqRIS/VkJuzEv
yzN8H3EN29QrPTplp7E3MbYMdGmp6Cyi+8cV/ExgkLr6164UvAEMqFAt+IoBl7YicI5PE2+y/G8y
zFY39QkxeZsvPRE9iKfPo3TX5iZU9NlxFsANZBrbXEmMIWmxJOVHhawafWGGjZLP36JvzqfW38Mz
A3gTqZS8DDhhXI7c/170I0Mj18sVwbOTmJMR/vVbk7mqu9qqZWzJ1AIe7Hj4S3XZG1TH8/wrjDQM
Wf6oRSYKVKQKprDYoaYltKvqpbwOHxsgpK8IqRQwnUTfKaZ+MMX8TOr1Lfzwk0TwJh6WC5ijKbqN
F+uU00ll3evuKKXxQW8glfy477+GQehv/x7t0z3jW1ZDFJ/Ms7S3SdzEiO7SOAEDHgPCahf/iaem
Su4I+HpZju0VRSXGYkLvoHxDa8bnqo2vWjBAzUopuu3HA9tWzz502wupQiLOlncIFUomprnBn8Hm
u27IyL+qJ3nmM1kiErs5FtzwzMBY0EzLkDlqMwOvgpjJ3woMIRntLB/DDoUmEZRK2eaeBvleup3O
xepL40o5BJuOa5z95UQIrcrYva6zx9niwS6G1xWQgNr6PRGEMO3ONBi6pUa3KBlMZwaB9aqC4uUB
KdvPwc1ShJKBzMClyeWndbbrC0PdFWG4uQHxV8wQowfXni3LI+T9RuJPz29UZ/jX+3N7YKPAFIYW
r49dB40Ht5LxShi6F3jkkaGg4msMc7k72X5LuXT76dmfz3R/3l0FUZGOjG0z3pBFr8IZpKda9CDA
VUzcCM9NNCvmfaWj+NTW3H9HNgf+T6OvgyBYRKL1s+zEkxl2xAaTLel5wY2aasTYqlyJtkBaggW/
gPNEjTHZTgzHSbnEBhvHngDEM7Fit5DRBGQ5Pkj63jdwuEIzJdRJhbKSp031IALMvaL1BAKIMw2H
2jYWIofSKLn4YxE6nk83P+oiMZCVXVMZUvrRf/ZrGi7YirYHh435aTnsBITYKWiBbg/kExX+ZaeE
04nJE5QNQEP+ta716qsXiGm5q6FOhPD28A/E/WAi4dIgnO2dSg6q+6NEyjEM5RkGaR1I0tkQaZ74
PVjCtjru5oDc3RwGBT2ITdgeUZAFhn/I6uVO7qSdUs525ZTs4QSIMBU4ebvZNQpYwW3V92dbCgQ/
T6/8qW1+2SCTgK1HmLZEArDFbdOHkogguwGZRCQcsPQ1cmwrCIn5J0irLIF/jzRJz4mdTrX6eJ9f
vmOER2HvKpyVl9jW3c4b1FbrXLJy5A9W0XolMdARHdqZ06vFKhJzd+CXk7vyib1HXIrZYDlvHn3y
YOUu8F5Hk1WWqUxecgYMqFTMEZIvT3Z2JdQQjTCLlR56JqqaLVvrb0DGNMYEYrcCDTAFbvq1sGWm
hA2KC9cC6KXJWTrlenwGyMDAlDvaIsV2C4ZuHVEuk6NnwL9BxaV3DKTusYfw6eznJqUg7lOKDvXI
U6KF+Dv8bBtzLlEmUyJiGnvPhLzQYjvvdTKmBuqpMteJ3LOzHIuqUwKniUd99MX/vT1fM0X9UgmS
1nQaQhfneiIZkuDNdg+7xUsHrQQXxWNJtwAyXOO+n+R+kRdey+6nqYYGGl+EnZaDFCYKc98TpvId
q/zzj3aZvwCcePP13216ITJqCfPfh1SA6JLRdoY+vjinscL0ab04U7sTd2g0rfeuTmA8NN9Ga2Sv
MC0tYUYDNyV/R9GeHP3VOCGNvQx9xWD1WMx1LuQvt+apbQXLOeqoOuz0+3XNSAlGhdJBsMelWM4V
bau3Ay2uTLxufQgawBIFfFy7oMnx55Ht/xpVJGzhxQhqINzAGy8+Q0ayZ3Pvf0dQzWDRsVICEnF1
aM+4UxtcrnmSJG4wKsyDBVdNHnfA3Jw/+e+pHZTqowBp8VM7iCTC7FZkuRCTdpL99+hgMpHGMpXH
0dvOtHt6xLURgxfrQi0hV6HFsv2xzgjCzOieyVKUoq6BoH9s16m71hry25Yd33mb6+tipvdllBRn
6GDHJmdJrTjq7nfTD9lEm4+qb9APMj3pHdYspkpWVYrc/r1TwRWA8e9Zjsf/8GC3bbvQHwXf/60u
FsEYz2RaWJNtmV281MKMk4sMkPSOKE7vhj6egP77hAp3iCN/QxpgpwlRqFXlE62Bz2dqkcmU634L
F2hYp/iO3ZNuLgz9HT+eX4ixUapuwb9p4cYTx/RwRUnUoEb0snZhC1bmfwd8t8bIz5g7j37smz8w
5MPqcjEktLOZnbpHXOlObh051Iw+ZTzLX9snO5t91UL1xkZYAz18lpO/kfQiys38OeQkytY9TtrR
W6MT4fFVVaz92hdkPlH7SXTb7NAfKbUKClbur0pJdtQRaTUMMXb7w9dX79b5C+hKQ7aZvNt6zzgI
WuIaB99oftDYrmwCxWIce5fghvglgvmzF4GozA3AW6Op28DJAJzNgld9dhtx1g5k+gQPocI5nd+q
8DbAgGQVVMk3oPawrM/L2NWB3Z63611ItIw1YVWndZukzk1MnwwC7p+kvLXjdwNwDQWO82t1c0tT
4NapBxRUsp3W9/Gt16xLgcdZsmub+3OSlXkgI3CswBa7qCVtoi4OsgiqzwvOUPeiYl/F8eut6Db3
VOdMgK7PONRBcz887bHVmkbeqwpd19jO9lV8EW12NRj4XO2XER4Tem1253QwuGWFsgEZeXUMHKAX
IwgO59XLzlToFjE9imt5rT2bkz1FkuNhKr6k8vwwka4QDjQKRIYvLFWnL4Upw+qztomImaqh5r6n
d4oS8ckkhsdPKTY6qKDaQqlJRRPvZzgHbG278RrfxbIXIbJuAZCgWL/xT1fTAG1Fvz5JUxI16UtH
WsgF60fqxnfLt05wQjXS0zSlBhD7VSveCkwlxXney9jfCKph2DcC7ycjX7wCa+pVtnfDvYKYXeMD
yw+Na0RFEjo6D2Hv63BKg+Bo4cB8Ml2ZXYpac30PZJE6LBg1AibLwCsoEl717oiM6nWeFVHtVonh
npaIT0yKQYe7Htav7GLkad4LF9IIUQbOqfTfHvmhba4r9scWThu4b7m/cYhQ9Z563YeTsiub4pLJ
XKfeoIfAdB2/3srZEdZ+Ivl8FyV73+UU1IVNqxQ4/FQIbB6+WHN27mw1PEO80aFtRLnnSAhAsrxp
nAHUR/wWA/fOs+jDTa8oiAczylv1kd0QjVDPKk8S+oLlW/T9A1iAzl3zKw102xu22rSIoCjlsKaE
GPBEQvt/CW9qjYsBTmgDWxzq3Ez1c9TUCrIJ6BJyhGQekWef2gar5PtkAoqvGbremutRh8q7Lk+t
RWumM0aT5P1qeTIsfNpP1yT4Gb7gJIaBBbml/PGYt6QR6clJx00VUpZ5bg3J7ohCOqjmVvtFkfrL
R1ia5ty2RiEbqUBZZyf1T7+TMYcPgqFCaEwAs7aSryVq79VwUnDmIZ2a3GuzTIVL19pQEUBypQEx
hKZC224Ca6w+51TquH27IHoFi0jRYnqCOerR1NHU7CBzriQacA/V2r395dP5zubs9NzGp/XIbNK2
yPkAqtb1uc4KecRR36C7xDZ5M8iza6Y7hs9aBbGoK/F3czDDSALHEvSfjU+S5m08OcjxzZVEMiqv
PL5cilWmOTFAv/Sjf32aCnRwBNrX8QW8PrEcwWwSVJ69GVRjE2yu5kg8MSTot5XnoNlaC7pQvT3C
/Bg1N1Y8EjJSXTD1JH2bwUjZA5Yf9cDIosZEBtNDBz9hcNjW6Rxd8aNmXtX9+s8KcLeJwFAtmeVh
pXyaaFS1LUzqW1sqmEMC3KAeXaPFtBeD61lELqlMt2BW3N7nSljLcGA7Xv17IsyAkd6YOHqAg1sT
f8wyQWg1ju6QCBxaAPlj0J1OEGEtS2tsK35auTHQIcmcW/4BOerTDAhS4RvY9v2zvjY45oS4q8DL
hMkZg+6whXoK7VFXH8IrS/6qKjkMnFHmh/baYHAQ+DSFy7uUnSJ4ElmVIZ4TsAFnlbfoyKSIm8VG
pLWBu1cFZTe7Tyy1mNAYj+stp38FLqshrfoKNzAoc7NvNbbwX+tO47hFYPQb8BF0tdv/E0LhpRGx
rZU6JFPjJ7lFJZPzgzTwgD0hOXSow4fbTiHY0lMSEGDa8gvu6VT5Z4R/dprsx7HCE8ZjGWy/apxI
G69LGwDwIYccAlKfRztgecokdF7t4YqR3zkx5dSrsCCC/J3yqdId10n1IM2NMVL5wFvwm1HFOdR/
HH2wyOqwwk+ZRdFQvLdZXnibZ8sf8dXcOesKBtksz4MKRpvWY7uCeKxySb39uLCFOjHuQa7cKYWz
J3GuQhUlFngvmFLLjRabe49r2hXD5KAQL6fTDguvEmmYtLmHzbDKJF/bvyL1uLhCUwCnJKbR/G3u
SmBf+G8YJa3V/vvrcHhNTf7q4oFgP0Fd2GXOTaZWiezZaC/vh/YhkyWE1MnFd2nZqHO87lYgOthI
TOmp48gE6L4E4GjFznG8iFkyANDw27ksN9BzhQM4+mUv1PfSyoRJF1ImTGnVi7rY7SZAOGuGXrNj
poB1e3P6HVeeMTVAHnSUTkDQlKUHUN8ASZPnN0Svu3hvJKa2vDz0k6cQ/5XmyGEaanE2G0C1ZzKb
axMlypaK5fcAMVVM+fq6jaUgANjy2+n4A7xV2zq/1J0TFBNxzTzaS+niI+Ry7AF7vpjgnta0hseG
EWTxjy7CZUXv5Ok4auNgXkAhz5hjkCgIbzwNil31fXjaJACg9emrXTfsBza1OTHkpsLXFfnPb2oB
vcoM5Q1ImKKCko4528gPONn3OuBjicHHKZHOjNPjCrEu9dEiUFCRTIbnj957RS8/BZM/09YOw3rh
SPBAb+UGWcvo0M22CTvu4Bw0DGt8POxuo/Z22+LGEge3ROUiQv/wfP4PJAglUlw2QuJRRIoivosr
MzojCOchf+38DIlf/QDeh5hHPC61vynA+AXBMZdw8Fv3zpAHJrSbBe2tXn4A7nVvrCkb6bGPQOKY
dA2TYcJXFjLMhZmi0N3KXsPm3xwxZdWeru35JOlq7n90YIU4UVAVBK2qSGjDDJEovD8sMNozK3tV
/8qiCO8LCbzPwQSqgeYlExVjYgjxZ/F2+Ze7Y/DOyu1mbHhSl0VMtj4lt8LxKk9eMgwTzlOfPRy6
4Juey4lpR6BSlgLpBYPGAGLNt+6ACq8Y66Cf3h7pn4DfaSKdGt4QiCptEnaAGQRBZ69sfNeiZ2Nk
R1kYSNIcZA5GQHHUFm1Nuwgw4pNL9EoQkToHxAY31K6O4v0HWrFiDSM/tpjq3wF4oPg82ogl7JmZ
4mB23ilCry+XIHypBo0LRwNP51EG92QXqtEW5BsQfdLOmm4qLPSTyqVX6ZYopyjJ4xKFYqJbFU6Z
cZ3Veeba1KYE9A6Td/JRaH8tomRzqhjYO5tF9sWMEhd8AXfQvL9PrAVHGqLQE76bkQAtoT82mlHV
HUWC9tByRNqTjmgF0ovmJMBi9eTrfdwy7I8deW9Nibu5jqIpXc7iGHuXGkGh9LYp3xMYJeaK18HD
LWNgeAcYd4m/WnTE+WjMK32Cz78PpI7y74QJjtBF/rTt5rQwRfVNhVfJCTnHV+FHnXFpm99m19/i
Bv5vfs1nk2Xl5/dcsd6H+XWyOKr7iDY8G3WO1tDDP/0IbZYkP8NANQEfBx5sNaubSP6WwZxs8w7B
iS6deSplynvso/R88DLfzaNSkZzNGLKwVQ0J9l6npnuqXwQFz1EsmY2X8aSTilOrdyN6ucGKRLkL
NW1HQ8E8H/FkNtfZdGngYQrrMJAdZQdZd07Rf3Phf+eii+zg9RBrx7pvgyYauxYKXxG+r2e3OY0G
ssd5AMsnKNDNvMpoReiIpY0TzWVk770+CGcC+bLkvW2LasFFF0vCdueBWdsKJKWLcepofQDud7TZ
hnHYz5q0bZX6tJOZuUsLA46Yiif0QXvLIs+qvVAySnIC+teCEaS01nIRtNFtgCPFV8Sll3KafxKd
7B2jaaokmA//C7xpJ3qj8iGnH9ng7moYEahzgehH/JeWGG96VguNMzAFg1YlOeHIx9eq+XcVSa1i
pkEBJlOq+lw1H0HuZ/ITru2IsYhgC14TARyQuq99UGhsBTNgGZ6AscGFwbUUDX28CsOU67Ym2G9+
XNE/8dODxfMYnUvoCndmf+PE2A3yB2DwZ2/luNvJrra5uvIh8T+wBhiktxhCtgMp+hK0ra7hhyCU
maY3gRFEzmfvvdJSfjNMvtpbV7dSaP25hPJ45tNa/MABzRLP471+xoIHDVhxSkNg3ITlm3o/WYi6
TWFt1mYjDGqk4/yiHeMpJHNIU0JWH5rwXjjvF13toV6EyOp5uAjIcd1WkFgQmc4Szp1UskltQPO7
7iVlkeQSgF82BYTULQcIQi5i4Yi1zcNQ4jQ28QsTQUIuqrSceNCWMjIZh+BT1a1ZXIRlkzv/2cKC
BFaWZhK0NhKJ/vIwHQiVTkVHE93yIk3MjDszIsL261LKptpEb+OndCnnTCPxvHEu5DG5VVycJnCv
kqUjM0P8Mr95RHSe4ipjKMnqs4tgWBkqphqyTSq4CcBynyGl5GGdEYZrIccfSsO+Nl3VjjU0UU7l
guhuS7PchEY0f+cTHPamr3JsyN4CcomnIFaAe+6RGJcI5SYv91wPViNVbcplgw1ZMRxPKJhM4eCD
oxcyZHYpxEbvCsqng/GubiPZcjrdLP0sZbjoTnOmW6lzlroQORaxoT3hlKN1IDfzF+JB/AMO/gCw
RC/RT4fr76jghGg/uA7W69kcDN7MmgTollXlTWQlhJ2LXKMLjKWogQtztsMPPGxfs53+qetUN16d
yz53mgwBn7B/TKlW5GOis+bUq/yDb3sDogRTPOG9Aix81clyDZvvN3M7at61nnIMTDYhoZjdtHVk
fQDkNj/NcjcMfiyq04Iycu2Bg5LS+FvsFUsJNjYa9MyfEPSDQSFgjF7+TIWQmxDnqgrlVC6x0Qiu
aue5WtL+G8ZGXNRjNsApqTOmGGK3fI+/IKJx9WEiPA5BksT/PhXDDOsedWeCyTR4qFclRZvNAzvt
7XZ9YYZiP3NZ4seYEWAn+AHILmGfPKa/mxbn+iSSBR6JrZuoLAgrvtlFzVGE/m5RUuDKRV3A4EtW
qG6gRsbA4biemcmx0qqfhOEJsOnGvVmb1y3DNJE0aqe0gCPf06LgTFIMF0Dh3QAaoRjUCJg/6ZUo
DtaFcfnFV8Zigcj3RQ77nfXnBQvYAJERrODnJfOKMAXL32IIETKvQYTXL4vo4k6KPg2sDLsdXSyT
U016WVtzZAsdno3YLXlHlz4Yq+bXOBqTlOyzB8qiYvsvlHJ16pmKS7RfrAlwPyOtU2mKSq3fnws2
wguzYex4NsMYZBLiBWerNHeVjJy9AXcrjLBd7zs2kbhRnduA0MWhN3boKrrFLTCPcINGxMA0JYHZ
mqkF4Mc+gF8svCFY1Z+aXuaUIFmpGkcYqhKTBcRAD6cyg26JwEDrs41Ly4lIhu8kQLB9X46zshg+
mFjYibO2iqorNK6j1ZDv25r1EN9cu7dConm/TNA/a0k+W94SAbYf3ocQbxfg5Y1pzdl7MsZT4awn
uagY9eCYuxNTxcgy/zph8OaRY5DIPkgvxSSy7uCsnf69F+btdcwbXFoQFxVOINBW5NWJhqjNMpvp
LAY4JPf7H+Ah/pnCfHmzPvk6CNQYCiBV4wZ0uVtxlFybm8a5NXvivrIwCSPTkIHMMZRTxfP9zhMv
p+YqyGmO70QAMQ8V7DR8UoW5eQyFKSA3gR1wD479PqLpAInNiKiK+prypGD/9t/hp2uCDl/9kaNg
tY8nXpNY+m2tbDDnxlQm9E7wKLmmrvKQ9UcJSt9wwO2DjH+B8x8bz/zimIvyT3E+s5v6lUAwD8Zw
ygX7YPxg2uidBI2t+gqTY/JRV/x1UA0wDX0e29MRL/rXViGDsLpd7uVrWD32FIqk0XCSBDmio6Lw
OaRHFuIijhTBlmSBur7Cw6Xn5i1buwaL4514NcAXo3OzeB8C8WcVoiNE2kRYWMr9KsONFleKYO2S
OvhtQnGWz4nP3mNWOVI1arHn0gecubPtkU/KR6uv1FkhMzlyXcMMDkOFTTvw9wPZr2ryjMSAX8Mv
baHVl02Z8x0yryCGOCC0iR/L02LAFhG7akq0p/ENXeZQnqhH3bBnI7pktdqhq2IAvTCpIa7/OjZM
++Nqsa5QocstbclfOw7UB7/QL6xh4gdRzJG2NeOA6KBvIoQEHpBNLZrQWgzRxj2AAUFoEAam2uZF
JCIi6xddxyjtgFpQWrrvQVS4A47zyu7cs2GvP1aC49rdTAq1EZJUuJie8+/uvrujW9QCjZp/Tiv+
7NOLC0X07GyiQUO3uxCIWnizVUje5MmICKibHNzJlxKb09o+AkOvDDyFDDa683e6Ns659CaQ32NM
H95rCyfs+9FNabBjC7Cr1Ejb7Nbp/oQoHUaNmqkKfeuSgX1l0vrZcENO8zyBGJEWM9slg2qKA2r3
3cj4PdRB8EWVYDytrTSF9to7ZZpnCPlmrjbUpybL8MR/GzMG9T/CFKvUsnpRb9ucMl6E3xSn9YGB
JqoAyK/7nMGzPtnyqVYbnMxI7PT7rtKeUvpp9NAGCFb2lYhSOc9oclNA2TdQ156PBod/vEizl4NR
RbtbB3JFXI8B8O/0e+yIo61w68uAMYVA0+6Qo2Ozf8jL0LZ+7f1tQeD/5Yyjd+sakC70aPKSty+k
yZgPYxDtoxaos8e0sUv2vi3bnhj9dj+eXe/BdFDtQ8LtuGMx47AOs9x8Al+3o7Cu0XB/mr3PNInE
047UqsT/FR5yLQAyDzx5qIUfKSzOb/mg6FrBBfsS9KV3/ZNoF/LHNlN2qXw5y82BzN7jwvWwiJ+g
hhxwhexWrSb87ALTlz1t/F/ZiT0ym1WrL8lRz5R/uAJW3y/s7z1fIsrKAW6RTpzSyBOTLnUWExDR
YrUZFx8Rz0ieIH1E/yK9RnXYNKseGwJWMdfZ2oAEfD1MCoN5cOxYzGCvDEFFUdLfAjupsNTIT7EM
jTEOpGDf9DpFR4NQVXenp2TL35FGWh3HpjCi5ng8GkcZ+Z13hrU1eN4eE7nF79NAQRlp8Q0EktAq
LNUMgCvXt9cKz3Z11MtF/0gKNAY8QaYKkIvbSVfAB36xGKq5qlTtIZYz6v37jR9dVVWQC8p7KRiy
HfD5Txnz2mOOTpjGPiVdouNMzrfp3T+n26OB/2urE2j28iJjhGdrejIUJkmlWCiLvRCVgcwTLPlD
MHlcr2EitM78KZVIiWNUuFW6CTDWfkowd7HEPEbPRBJ/mqyTu+ErTUZlLHyUrdDUQLM3bsu9qKt6
Y+JGepwHTOjPmOf2FJe7MWEYujVUtWpGSxiFytelbxIHX6Ri1eqQ7PC402YwC2PwH9AMIa6QIQDl
SUi+YtYZNPkEyRmOBglVO3gFS+wWOl3kL07gU1vNwRB+4E/e/peN/iK1hS2AgyMqctdwvhfWZKwJ
JGaKMAKlUbiI4XFJTfikebD2ylimnRBkaJHofiHoUzO+XJ2YFx1pVMLfGkJCQXnnsAzDmXFHCl1H
nGjXMqLEDCGhJLzlhGwzrEL6sGQtu2irSZPAH/+HxqeJ2/GnvR5eElkk7fvOeDVIKsLAee+eeYCa
IIx1cQEfUhY5WOOEvV+Pd0qRUnTL/qG+K3xoqqUr0ChhnA0lDyBmvchoLWhOq1SpCoY/zsPhg9O0
R6WKuROuN9U06Si563Ml8PivrtENKmt0r9UvD+17OGT4rPwLF3rIgCgliDmpaSWFnC05fDgzwVRb
AJ5/D2ZH6tQGSZXsulxXx4itWIrOxZxgO/O+MnZM1jsTDBeYqekQFVjETzshKWa1s4hlIU7VZYAS
pug9nbuMTnimJ9xlJ9n2GgGIprc2UYsC6venlBgwBydJfYCrAsaM63xzo/VbSaXswoVV1l8EqR3u
04EF0LS9t1rPozkCgTQy6pxqfZss6p0mDRRs2RiIPwHWeUKuXSupPxpu0E/KnrLniM9fldAteYJV
cUqe65KqOy4geIJ0JVAG0Kuk+EqQMcvMwBSqX8a+wHMV8lVzdFCf6nG0wYqIy81PpYEP3ZE/j4j2
zyBtpF1hoPKzrGhZIDo4acmTeQTSUetCH5BUQy282I9reZe4AwgWUfiIUboPhFre16quGGKwr67A
o+OwqO+puY6nvCn1SyEDaK5DVd3mf/joGCTp0bKgtSwbklYifBz5f53Z7CB/GIcTqN1SsDmDsdX2
BDU9X6QUQwaNQplT8/cfPHgH20fJMI4OIYzoSizRdvHbb4uG4RrZGnJwCr0jB1dWvlY4O86tRnFX
GHB/J1B7FrM36FxkE8Fxc5td2HLZu2ZuEuH9cojNFYDnO8x/p1FkbQT2GYdOlp+AYEspAyyQYobF
Biw/u+kOHUVn+3lpfbOdGAt+BrXQFHiEHBj3Bk2Y5+BaLERrhFH5RnNW9Apvpy3/cheGgJmIG+eg
2BRmGTF+3luhY9fsBJ1DumWZJyqhPfe4xrxsOrjy/X360Zp3IH/sXQFes41mQoecsb0zZiwGzSqb
cn0jWapRpe77wb9uUWVfJmkTTIcudPANe4JhenzwLdgnq1DC6BEAQe8jaosRwTLTVLephh35uGLY
zBdTd3/jMuhN5gL9BaMeqcYUadXW52EaC7L3EGaC59J/XGBKtl5O2OqNWk4YSXWz3NBoimzg0NUZ
42tcRdNHPFidwaz0GbJk8fzlRnWhFpVBJoB87xGidV3lHv0oFjTE24KDqE033e7Yz1H+Fh/B0FT7
VvsGhdBy3eUyiYrwC0PVgDIHVVJXdJxIQTW3l9vz04Ia4D9iQIeigDAAFAVyRO8FJKTviZLHkPqG
stuJvb8pE4mpHaq6oXlfXM3J8ka2NyOhH6PxoOI6wjY4xN1dfl5fd/VsroYt/ci0nOi9qCtZ0DCY
/KWcMZepT+YuneMAx1pgzhZHHJN8NjcUIvqEHwvF+Arb+9Pvc0Jp9gaVmlRreO46EU3ovTP0Lm1V
emid/tzUcU7MTbDUFHIzUD+WapC5ZVHwz6sXiRs1ydpe9pN87H8AaZ70aWiCBUqsIBFX7ZUwLerC
UonTkCanMuy0DlAFiQ2lYsYmQAR1EaOZASyS3qnJuEyBlzoGxlIGiMGuiGP0jywNOtwMRxWi2a0r
RwsCah5FY5m3yiMVLTbXFK8+O1Wjody2iWgTx486bL+fU+V7xk+u+etsnn6Z8q2T2CC1KZSmIwfn
SU2ezalo4Rw6bNxfEuj9LeWJ2S2vtsKpQZX8+PjPYlDKn3NXdQ0AGFfV/8tUdKy9Zydn93H86law
AWvJqwaLmluHE6vfZk4eiPLA/HodUu27E679+M+L02mq0Kob0J3k3eDcd1qf3tuJFNXY/sGI0vCp
ahjtxufcmmNu6Zx7AMnUjjyFFbJCxI71RPdkq0yEt379jDPibpSqqoE8naUxu0g4l7BWa0RqQDnN
fFJh/xg26WxhsEOhzWnSSk5VkTu/pukt3lxIgGbElkh98znxHnLKu3X8IXBE1n0FCfJN4NeYxrHV
dzzrJq6+XjeHauOgpjkl+9UEsUkixC8IAte/WMYk5pqWvCTBLb62/v12nDOHYmLzRN9BRUnqaS/P
NXVT+0Sk4mRN2Z57s9GuGDzelDDLUyM3XLaiuyppjPT76wa2+1+iN+BpyXdqaY6XsY3wGdzRABWO
URgMyzlO4xH72GwTgmgTjd3iJcdE/+JwGQQmwjj0yS/V42yIjt7pnW11i7fA4QrNIVI9mb7TWtz5
pqUAn3oXKsl/32tX+H9Cp6bY/YGl1/l9Upxr/x4LBZlTu2FRAisnoT6oKMNrxa8CyDvbO21s6LEh
6HEMuN7PVFJnc4ZRNdah+RYmxUsLCQE3XMIkc6gaAFsJek7jDN5Cj3RlRvsEAabI9L/ep20YrDJz
X7J9J/AuAIGJ5Xxe15np2L81BeAoro3qjXvw4PhlwY5NQLZ0u7gt9UXUh0lK+h4M+pe6pdWWQ87i
PYnX3/zFA2MjmyavWc148Jrhi5Gi44pw3O2eAYm4jtzqbGD0ieXhUoyECY4MxHuVck8F3l5occm1
FM35L/uymaoC/ZK0UMRsDVZjwtv1JSHVsdXfS8Pl7mV+nQJoEVoy1qt3v+LJGnx4Gxi1oDwaaZJB
Qe52RjUVEMOgbBL+wdEdU7N6w/GEcM5lDeNcqNIUVvBurU+WlOMMKwVdNV16tcTHgmpeD9KMfhTv
5mX+iZVJHLCxkR0OI+1JWt34fkWma4i6xpnPudbsPqxyAx2FfCbGrGkbp6mPRJv31ChAJ2MKJXkr
mem2r6q/KLQ+4iZ393JoGzT8S0Bvl0KAHNi+ykMu7zqeyCJdgt1rg4NSyEtwuJxYM4PcJCqrzYsY
JUEuf/IyzRenMuMBaM2oB96Ol6hBc6rw1MTY+8H5gZJslX8poaT9/EkKgKzcCCeGzoGycwzRUQjH
ZgYIjPdhEtpsoQqEIIebyfQx3Ml/d15LjbH8tCySHHWL8Lq9QRTuEDK/WYxxAG1cHFNxOuxy3kT4
WulOqHgwE0hK3NqrRCY67nuYDqVKQP77v+GWkSP3GbuEL3tA2UPNtdvmBXonTQtu1LbT8Qtian8h
WPtBgDQb3LWc0VO8Aq6bbNIENGWSBO52Bj/PikokLUmQZM8achR20+1mhASWHz2OajlUdSk9nfLK
EGGDDrBH1iVjBRY3Ed/YqfV6mqr5iv+Hmv3Ps43r+6cVUfM93HQVG/G7d0/+rYKIDccZWlsauRLj
UfSSeSZ9CvU5y7NZ6TesKBCdqNCc5VCymLJRaQucl+28d4yKtJqNCSZPzTMVV2fi68yQMvuD1pHZ
Zrzs/6z/Nc2h0okhcJUOgYyp6+BZS0GTG21zf4Puvkf47iBPwpDjh+QqtZqwEawMtJcMUIdFb2mT
k7V0DVIBU1DVxi5jFkWzf6bkYHYtxCjfWFzI6ArHwn7LpqCAMYPbr5/ekGqHPF8mkrWJ11pgXAO6
604dgnjmRJ/yymoRvK0J3/Svy3/scKGhfgz0+SA5pufH0dkGs1/kTlrbWTfrnE2Np7gqYtMfpOQ+
Llq6bj00XtfGDshutTvXjnCePSW1bGtxczHWxx51b57BUe+uR84vwssUrOKrmYkBucDgSCxFZlIb
1aG0iDHSzhfE0Xp3y5et6pMrnyrKP03mqrEnuRktFuyHNPPJfwwbfHojdpd7oRFhDWPZeE4V6ZT4
NGTUSSWgILcwzz2juhd/IyZpLXGHNlRjeenhmykER22li+0vY/PWdOpxEB7W7Dlyi22f8rjmoU0Q
mWXmHh46Cf1vDNfvt/QNuT8gvPiaoZ4r9fYrHoPwljlTiZYG0LimzoO6I0YDzJlZoBOJpb85R+KW
/emvjlYLZR8ROHp92BQbqQYDPX8OwKjEp3nlTQ06zDtljlRalfyR9TyaY0i6bnCcZ43o4DeHmE+x
Q3wPkO8lxL98XuZ+Jd9sm3Zc3094YRvRSze0fxYq4XuNbAjPFyd43QBDaW39hTi3ioJmajgIB+ew
iENtIT5JnNvmoYwZbmNvEQMJnYxcNGrou+KJ6732RQMfdDDMNS4gWySNDyOzxUHg0dUJtE0Mm5OK
4BWuOwE8NGJWd7xrPHyLaYLU4QHaoP5pv7Onky28XxCC3RuY+Qh4SMs/9lBxj+TQPYtq5g+B/+gQ
UmNA1chXQN07gufG4HmrMMWDsFb0LB+ATTaiy+KYzA9R/pCBm9at81tgr2Ek8AHvZjWt9vxIYZeJ
JQrz6G4BR+Ywr/irP5GTT4V6Yr+jnMqKn6C4DUGcMQ1ER+NJf+hlZ2TMTUVZ0w96pmp0hzYoRbsi
AlsoCzR/ZFGi5yZCu1jJcw5D6E9H6Ay6GVsOVIc1x7tUQs8dzcTpc545Fd7Rddzv5bX/tJxx5EQ3
A8n1sY4EcLaiKwafENn944a7KB7dzXzDFLrEgxILZOxn5VeaIWtnuRVutYkHm59OLdsapHIt2vdn
rbWG+anj+uFGH+kp+/nsrRmfFv1x7hTZO3hXsPjMS/c+6wRcFRiUg5PSYe7RIQD91sRK1QYmFlDL
H5k3i9eXXofUeUYcG545PvBHh4pSinfJMoTX33SEksyRYOf5A2/ITX+TeyWS6TMlchqXFKvq9CRa
FVgk83rbVHW87lf5/JPIrLVTk4WVkYXqjD0jW2lab/Xo7c+owyMZrazONbe2QdogqJTJbiPKaSER
m3dEUTR99AL6GQjjauqu0hPp7XUvqR53b2V6erGxEXFh4q/w0C+Mg70eRnSA15XbPumszIDfucKW
DGkXHHaDyH8RSzDvPqBmIGMOOa/Kef6EuPtofqmEceAWRUam710AVAYAvx6DoiJQ0jAwzajhWln+
SncVnjN1laItnZ/L66aB38aPJBwlhEgM+HMXHh2E40J29jF6CjaCjZe03vHPMS6cA2voUXa1UaHt
61/N63k+g853dHzjKxCDQ3YkOLCeNQcLvzjfaEoBPkxWWgvBLlqE23CEAF4Vp5EnKLq4pUD7JrnT
7Z2OS2TEJBDKoR4SYt80O+a+mRiXIjSgzGQkL42sge0KBDVqaXaLS5g+y2DKQEj8uwImh/bshPYn
KfFMqB8NeE5kSg0MvneGyOxRnXYV5mbk47zEKhfYMEHiJ9zUAdmxCtX7NBT5UyYfeq4hDkCrZRjC
pnaa2v4f8rW5rpJ9VdKcsRzQ8fs3iNXEo0l3sDIisu60baCUIvIuOoJ1uLPr0MSKJCIFAdAOXtqo
CI4JDcAYF73qxMaxbUXVM3M6tC6VkIWc+iMr7KZg37iFMpuSt/HKBY0tnlpHlnCwc4gIlsUpiq8b
Tb6u+LKiTycx/jmXOpI20Gk+pd2DGewdBgsjigIoER95Jwu9D3f8b6tBwsSZWVZizE1y0UmFGnrj
8j26M+n6lw4WOkN/imdx4DPUplDwc5/r3BkLo7QL07s+Df5ArYPLplSReHU1WY+SXotmqya2xoNN
U+YS0XdLIfKxspzJxUFS8JTaq9XrmkKvBYbGxM+2OXEW8Q1o/E5OHGphpqImIAPF+TqTt1FUjMqN
QEEqpdddq+NWp+aUx3TOTeQO64MR0FbzERJ8QJkda+Nf+LXrtbhluiv/Vc9tS9WAZPULiA1ibzmE
223LEOtN+AEpeUWD//sDtdJaH/FIT0C8BFgA8tJw+Wro3m6WR+etBrkV2yfOHSh6XvzBfiFmfbSB
jQzJYsbykyeWy3bTUxPAqKuljS8mnAZzzVXQ51Ue//zpq60jn4/9uWJdhkSK5Vy9WCXjaQt+Foou
8SO0Phhhwd1yVePk5D91WJ8bqm+tUotWHazhPD+/POf3KPBN0KMCHC1KMnu7J4uWE81gN9mogYSx
ny0aielRjZuUatw3dmqYj5ZjXhcqgH3I2/at+DOI+aTS1osY0YAjFslpi868D33X7XKMcA8tSD49
IG5fG7B5LJt09znw6fIMvcP+Vg2vVeHt75cLQMfVgYBhFlWDeVkPKqfVHD/9kn4tuN5EL61NrywH
8Q0ILkYrpkHjHItvhLa76G1NoUz0caZQ1rtQoE9AGxujkTKc2A/1fZ3yfeTVmleiEzssFTcoRFEc
Rfl242jKJiBn237HTXso3lIsE4B/IOIFZVpNSmc2MG1khp0sUYgYkVetbfQkbn/JjhUCOSfz7M0j
wDq2QFcxco5rS0ANIY2z5SYeDeVS5GQHXaKL80G+UdER90fJ4Gpp5oQ5bQvsce10L5soILJPAsRD
9//9r+Ed6G9nzAVRJQT4KmGfpdYYkgYa6/BHl986LmsYd0BuhozEFPYptP9BssyjZqxmikbiQWYh
QHSejp/39hFVSjstHqnHUttwdcdsHgyH59Ws98jkjg0y6DezXXjxziw9km3XFnFoV6mEaidYUIXb
lVAzqdJwer7aBj7XWyWq/ekGu+8dVKZUt1kSS3lngp3IolKMZ0sWfRPHGSxHsEUO5vgoVKCU90Eg
shaOhutqysWahImJoqQgLfK5aAzXc/3n+cpa+/657MrJDgSmkBw3RNomTMpRyZkH1XY35y60cHIs
YffMjPVbF/kDDyUQTjKjP2AyPVPdDcad9fazJxnlW86sLraFtKNmJsdgoGjJr6/dpocJNNvAoPbs
aZViETEANJkfp8MLljLkj6QNtCESACyoyGAhCQl8PiBXuls2A9PUy0c=
`protect end_protected
