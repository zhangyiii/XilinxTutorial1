`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22384)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aPkk/LZprZljgyNzZTGF6gcxBz
LkEl/7f+3dcASD/i/Kj5BrGQGPFMOaSER1KNI3/XJEw+A1hoa3l3Mk12tZ9RVZl4yR0gfjsXCzk6
pL/uQfackgxxFW0V1t8M4/p2TcbiXwKT5clPXgXR+iyTgUowldovcKaRmXf85kiU3Irr1UwQWvHu
R24W3Na/q7/o3j1kbFf44meZZLYabbnFToQe6cjJIUdSmO6hczK6AWx5CvKu0ertjRXiyzDfZCI4
RD9FojLlVWJD3w62utwVOMasyY738Qz1xn4mDtex6JXoGqkr7ghtiopFgo+3NXuw4ibM6p3OXfcM
qWvY3GWRUrMGX5yNDxyeoNNiDDNxfGdf5wftiyj26Q3AbfOIIutHtOBTCZLFcJsBSPJbR/Dv3ALp
XZBjJWYtFQ1bVaP1BDp5ZYoBYhkpgWnyD/NRw73On9vzK/EUoPAJ6HytDnGTqRqpdFXcHZT8Z25u
8YVu787E3bIqNgBfm6I5ipRNJ0Lkv8jD1PcN+X82ArH0cHK9Opj4zklLOd7isUMqTgnkClEoema3
f33UBWDq0/EX6gEMOnZAF5DhXPfCaqyhe7mCH+KQ2nxvSnbljGeRiGO07XTsFw+m3lG6x0kzxchr
r6xis/mNCmAp8t9eP9/cq7RIQMWmuDYZtMrUhk9L7GnZy9oVavqiukDOLk4nH3itOHY3YRd7DiRZ
869mTBMucPcC4oXhwnFtz/T7W8iZhvLc5atYlzopreflT3MLOcTZXRT7wqPUVQVk68SVB/buTqIn
Ifa3M0gl2Ow6KuV+4jaFxHCqWF8fI1LTe7MmZq+yqvKMb+Hgkh7Ebrs4nnBYsBOlODHjaq09k0yu
aw1iUVv6pZ3vnfkrn7fVXGEgXwvlM510sAIrxi6EbldpKBdxjlY5xjxK4C7H8sr7PP8O1euHml3K
DlgRU90otHRFaMpDKiuEZh3tir7629r8RpnFDFrp1yh4zqiZcD334vExxMpEdr6dyOXVOLrNM6yK
NjIJcKztxLmiAPcRDTuJLpCluxkd5fgsVoHaNnXobKqEzu3Zt9RkJeGvup8BkNaH0u3I5fxkjDz0
o7B2cz46e1DUxGxZN0+q7KeRbsTCB0HvN4sOp6m5X/BIdK3Q53EuEeI97FvWCDWNyjN5SUvf+TBb
vjlZgmhBa78CDij/5gaL1v2/h4CfMqQyYlGAxTkODWJ8a/4YctxQrEK2UAoK7T5FOGqtyE1BprXZ
XhF3gkGflztHD87UupOc7F3kvfXxOptO+qhisOaRJeA9qAzXyWATS9AR/9DEpq0Gc8UCSBnaEb6a
2bYTTqPpowzMH0PC/CwkGImUXiwL3x6gGhhEXvgjB70RFoOf3JU2bhCAYOKcCU/x+tj4+uQHEKNI
wNlISY+R82PPWyBYdW1BOOxyhddGt/xIapwlx2BhcHfoWhw3ebQM9Uf4MN6YM56F57mf/SZKcNyq
T++zHzPKivcQnPZXAgvlRxdegCFOR6Li8zFJnehxqsma4K346p5fL4Op/WB5hrIX7xDlUshZ2pjF
xvUPIe6S+l7XrRyjUJD70gxePUlMigpGeLu9oMH+6N60jSkrfIhr+ta12eRaCO6nFgRpUhw11qpt
lcJG2sRnY0F0Qa0IwBcD42HmnZMY98B6gFoqbzqK9d0uvfYemgOTeDBkk84JitzfAfnBRW1L6o5g
DpdRmpHKRT2TuGwlRQL86EfgOBfMXahcQTnpo5iG5wOvUWqGua2ANERPSC+rM09RyyHuwXUXRSlo
rHx7fu/FWfaRcn+kyoU0b+765yesZQd4b0q/sL/QeEMWM1l1Yq/k/DtexC2uIU/epqnMJbQ33g+j
SC8gbwt+9bxyxc8gTaHE+O+g8kv+LzlPxtv91PEYrpMML2FmlielEytKPKdhTIbR13XznZBoLg1Q
+Zb1dUH0gFCbLUre3dBZXvAJvj+Agpb1u+A3YSbRzMhrKLOWnTJG4KG3lDSDwJvcvWW3iCX9BdZx
3zITSEAaFc6gxaQxmMuGAlchGOHybZ9EacOBZB1VxHO9RstaEUf6PzSlSjcHYEL5rQIHovIKTfGg
05iVCiP4kT+YeiXVeXfjx1roq+RuI0DuB/YOT02KO7wh7G41u12968qR6DSJKiao4lLNnSIqlTYo
yJan2LXHXI7BdriApJkAbJl8ox7FsjkjmhjmQycOlC5qDwtrHreUu8qfdnYX3Dn4aJ1MG06wP/Ys
y1q+GB957s78WJGkwmgvDx6UDe3DwbDERAutBikmD4tSYoMi8zAgem0jnIAwrS9rBwEjLCNaKlEU
BL9sDAdYIDvlb61/1pyWpnbgaHUl0vE1rbmSevkvhSOVy0I1A3Aw2hydO8K2wMIvfva6beEX/e7o
YKA4iMzYrRIW+mrYPQJzKopkSjj50NFgEzmGKpXohsjYIlb8dVrse+eKZpINscMDT/5rIFSBc1YY
kGArYFZp7alxhc29MyoiUAmWoiIiVcAfnPG6zUwMbd8cmaCs5eqF1UJgrhDUX53sWc5ECxpbRWCF
m0ybe+kuBveH5h+8QlFR1huUADIpeMqbQ2PNqvwS46Vi0sjGaj8DtSb/xUaHu5zfTqBZeXmnowvW
M8YCxV0cGNOTf6mVgP8wxs7nKDCsTzzrRTEwcD6A1j5b7nEFrm3mccNieTPpG7LYZAiV4nGWHnPY
9ubW8dAC3QFxdn2jsB1cVNRoIsLF+81M1RqExobWCONkqMPD5tn9CKci9PW32FSX/EfBjFMJP277
0D1dF+XyoFZtO1RcZ2YePeaoNbIEXkjPG9ga6faKrycIeUNjc2J6Gr+GCZS7gWWMwynVJsxDL6wO
NtXWIrUcoaU4h0/J4feyrgptphCB7i/bVwTI6LgBT0Z948mwM4giFx9Rt78urjPeCCP+Xnen4qSk
Rlgvix4dA9HEcXb93W1vwW/qjhnxE4AzFoQqeTdFCrMQV3/vhfUfzSVPk6o9W/QFJxLFvhQNSh0N
/rWHYHqN9nLeafj9BcJoSaJGbIOn8joZJe+VM72Tfk0ss/WklvBd7r0DyNi0X98W6JD794nswVTF
P5rrJRB3Imo5PiwqIriFsJwy9ue+4mY/yP8m/u8bREkDkQ0Oz8LoFu7EHXICtx30pmgp4GBf9Zqi
aJdwXrc9Ztj16/HxOmZJhxn0EGkQ4ddxaUpi+kaSGyQcFISD1Rex/aftJ2TGOX72lrWNDfgD4vui
9nW7DLPc4G9rCqttrryCJ1m7oxiI8pI0gHP2BgOc5cASvnSZjpogFEXy+CwknDOHtXtpCHKhjAe4
6f1T0HmjvYThHBz7/pfo1AgRyCQ3Ds6FluV4NyMB5AREh/26fnOzlPrXSOweEFRMvAFROEN7fjZg
U20HufQ3Eb3icV6AainlZy3dbf8/9jyYNfFu00imJCeRCuzr4ETrFau3wqxXHjJhxpz7gPFVd5CC
d8Z0Lm03DnoU5jqSmnui2t3r2TNqbvc9+F0oasbpl7prgpM87iXSYuyYWnlhEs/UKvlJUKrbjI9J
qFACzEtSJ12bVAmQGNd+j/SczkPmfsSSWTdgHjF/brXKOQa0RR6T8Qt2JGmdyTBm6mh59lkPNLF3
OeiTJO+FRPv2fA0+sSmNwNGR31yGJoBCJhURrrdtv78ZZqfp5NyNj0JiYcFb+zTHc1VP6n60uKl5
EMpkWdMREU/CIEc9M6pk8MsVft91uKtE9+9iMSCrWUw957Ad9EX/Sg+uC4OajqsYY6AXWcGlWrvK
zkD4ON2R/oU5KyF1BbQJY9tHpai53qvmyBVGzVhif+L+DXRHqom3DMylAoamiwVoozMHTFsAq8pq
oanxexBDDw/qTU09qTz9oWda7EB4l7Suaz4LaziL3tl+jIJ3QAv5/DEH5xf/9z3uQppKFbkyb7YR
B/EJzD2w9gsvIIof/7XUyuUGLSqE+J59G/N7aCO5EedF1QE7LeztKmjZ5nAU4n00WFLwid68WYAo
N19wITBleomyF3mslVmFmhTHHQdj59kbE1zVP3K6GJy+qEGTb+mdvrDnRCSERumZPE2iSpg10L5U
KuBha1h96r9wKnSkkvtBQJK8l1FbM9TNpSCJ4sIGyCy4a/ty5j6mU6SWDpmqurSjbpIQSN0gg88w
eZyqoE5iW/PowFKwXILdHecNdKgIp/ctuyBBCQBsTOZ3UdISnkwwserzf/swW8PQ27QqihiTWz9R
1wVd/D3rY7E0wueMOYqSB7ztjYMJrZ3G6MCNatUowMzF3C58WEWoKdTWNv4oO2XjlXo3uDkb2n7A
tiwCz9TSnirja5ajd1ywqJql+86Bggf5xzjOkXbjQ8FUGYsM+sfADdaTJ7HRdiehruflSCKeFyJf
p2sDWqTlN+Tjsag+PbsfQ2k2IKtC3y8BwTxgI5Znse3SVyqyspz59Yz2aNR8wQfxbZk18g5R+8bG
J30bQTTlnupBYGjHLo/Yn0tchuEUhcbH7i+Lr2tKX3ALNKyF3Dhok2v5JVt69DIl//U2hID1X6Ad
kRINrVHna9sXTq+hzyNSt6EChaKkIE4ftnyp+0Lu/QdpxEfRYFNwXC0j+sth9uP61gkVFM92/FWA
2zpeZMcz639G2v1o2Q6etwgblvpAmlok/AYYOPAMhuS+5wP2927p9R4vdiZozpODnCDJ64nKhXvF
ZBMOXPb0lGzzUJPWq7s3YXj3r6+JChwP5Zi01Y1Hoih72IPm5JkIBJYLCPUzo6ufXZFLF8P0DOu6
gm6sgTUtrjiLLMZjqajcwdFcvp41G0Osgy66SKHyQJWNjMkDcx0pft6k6CriFZfDMVbBIw4n08RY
9/LHnXVeyYpj/VK2+KUQbuzb6evK74VIacLJYnl1IRA/PiYOXhfXnZIIZysf64sRLYqNHBuaficY
hx+GJzIHp34svPstwhMchNskp/UDEcm2ePdRcAKzj+L4wiYxkECuGXDr15kIdKF+elfJQX6oOc0C
48g0QISbDjd3ExGriEmyihQW+j1eQPn2B0UQyYva1eAK2G+hL3KF8x+89bquFp8dbFhaDxD0pZJa
ZtZHRMfqrksL+ZEcJNAmYQHICRWfG5/uuw+aCWoEJhiFtmhheY/KkhY0AzGJQ3Kw8wfDsj1w5or4
Cl4dFPCz0GEwsWno2eiCZR1i7Vu4TzebUng3ZIECAG9rCCYJB2f91To6UWg7anojNuoRnZLpAMOr
WN5O98TzwrYl2bKeyXVJni+ufgTXz+HmU2Fx2xoyb5hzc+/fmP7MXb5qUv7/aZfX/WuAh0j/QbyX
xxOAf55IiPZOEKppK/qMHUP48i2l8dsOxT84gjgUTVorGfLufzXr5LpFbqJmNRCCjCiVGrPjFXuY
lYZwmo5bQ0I/Tx2sqEKzX30sCmHDfXPeorHpnYOfz5KmyIE1ROt3laFAjjJ9Yt+6Hg96736KhcHP
KmiOmzfsfEeNZ2pq47AIwUdnAGBt+pv3gblReTKDb/bSen4QvcT1Izda7nnMSytUyJhMOkyg3/hg
c3tn8l0PdFhxs830hWH6lnsR9wIXYL2O4DOBK/H+Dnxjn+KrToRnIxzb6Xzx4ZjUSPU0XN55WYfF
282pRiPaz+EG8mZ7dXLg926cymWgO5ZTIv+mZSj98omy3BUGp+KwpldT5b82EJiqv0rcv/+t1Ypx
YRcil+dtLe7iFgtOPqhA23RVVASq5gqvfOIHm7+OEJBamQHXadEEC+GlbzdTb8uXLDqc3TLjMTEf
qAaBSAb8PSA0G7Rk2UOfvooRVQNTe0nptzfQQFp/QcjmXkMGZmOwI7t6U1U/LMpHgt94ILBvGX1H
UmhsFvD4qLUhtP0Du9CocpMDosX/3Mn3eqWnjknyhNTmzPEbBzYRoo3NP+0NYAb3310C6SL5OwBH
wcMJNC9AsKT/H3Em/KWF+DTjcQB9OIB7VuACt4RKnNlEorpwxlUCDVSvY5rW7/+xAunF6S5SE9OO
6exrlgo0bIjBjQ0f257Z6PNhg9lLIisxUjg8XLXm12aLlJihN9NMcLJW6C6YzN6kjU68gbWL/pPy
DOhgO88Du0or1wtcCQ4Exeb9p01JDs9kZ2nciDcZgrVhyOnDMCezFdErGCG+R6lMCGtpMoP7TUgq
i2upRQUjjp12hK1/Y/i4/w6043sLfiTDIpsVdc6ojx34y10P6eO0leN57SAUbTyCVUAG6ITcXa1r
NS50UBEhzEGdkw94dRZssdHXGwBC4qemYI+MiWfvvFc5/aAFRp+HQWw8+tFo7P8PdZ3cRbH0QyMN
NobEbQN3uPAt3BYV8gS2gb5Bsm/WrS+bazepNLN2hl7AIJuoobXM5ekw04gaHsDpjL7aUJNg4mSo
tC0fjQIq++zbL+KEe70ynid0OUulsYoz/XZnYozBA0t1csAaWw6y+HtM44JK8xlrYEHVpgvRp1Qc
JupkKf/Suk1V35lDxS5EvrD/FAoGgBvwlzjQtOBUPK1mYKsdBozjkdEdBNJKxHYesf2Mche2fdu7
YviIIrz4tqSg68nwtacyD/UUO2FvNYlwoltY8kzcgU1sDuz57VFjEY1n+FKBF110u05taHY7Mb/v
REkEXvBI8GyeTOS8rJs9x2sDoZnrnV9mp662SyXyB4PlJiD9bnG6VVJLspe6F6tylv2OKs+jVhAV
60P7/svnhn5ig8AYZ8h9+pQ/7IHWEqTdIEPlw6cPe4Id22SyaUYIC5TTTkkizOFcN5pQnc2+kUvS
HkJ4lRmZxaVRy4HJTkuwWCfcMlEvNeTtWGQTx+fX/3aLAhRSO0vY1irq5gqZHrciO+sYQYrgs/7K
+mlVyG0o7o19eF/QeIHV43IKse4MSxsb85quQlLafiW/8vODH2KTWq0d10CLqDMLXK1ODPhQ9LPv
+1iHKEUkjlQhnrXM1u8KkB+FvvwtRFwFuZ5nSXe9bqMcMfw5XOREX+DjvNOsHp+x/3ErYjuJogp4
cSNQ9CuLsodDnxhb3kokF2Q2TCj5WnAC8IpwDULmAWM2TxuV/pcIqEbSZkY5YTn0dNIrtdbUUsyo
OWs/fitDmDZUBxQJhVnSjLvHF749gPrYTPWtcPc8wXfUyN40tE561HOHWAxoQD0FZ0KsHHEDV0TI
jzoGDgtOpJ+tiUxjSpg6wg4JqJWAtmBjt7/RCc1PhfCGdls4deQEq62wCTykPb963UOTL028VC2i
nN9rwTxMJwQWOunJGAkpqnFsr4kl+LtmfDVGL3SHMZhcZFZvh+JF2TpoeW684XuFSFQlHDgXtv3a
Fc/l5D/MwCOAyvXSM8HsLkKYGpfQHRyLZ+WZ6H4NTjIu50u8Bm8ytmzP3xzfKstM/GS5GK07Tnz5
nwxWM8YEMR6pH1RFQ8QGzhowI3hxkdAZ02vURLWUV4jwxcSr9KFt8WYk/CZD1jJJfJ6Z0LdygGu2
KxsYGsUpQCCQggShZN/z2FIDjbyInaRBFvajkgvgZMHTMj/xaLwCzF+t4wzyVmDobi8sbGwpET2D
j0CIvUU54ilk86Cyf12yWXP5NqUNhO8+hWklEyi1pudg4+dqf9ezu1ctotnbDwF3v/URPE/WxghD
c2LyZXQEyNewjuDN4uVDNBzRTs06e2GgdQRoRvpbEOklkavU7A7k1KAg5asXraXh8LuyF2LNg6II
32Ao4FE3ksrCuQtUz14/rLWnjIYb+ruEakRWSiQXNxSvtTpi5Me9wcwhmguB3Inwq6Dpmri6EmXi
nLn2tTywfyso+MwdgramO4RQRDeUxdZbDpBCalRH+6SZuze1oB/76aCN+G4k7/h9+/xowLkdVaG2
uXj0/LnmzQgIB7LrxYvSHGFB+HVnc+1+Q6P3QmBIMP/JyOM/malWwlHyx6ZzDIGgkaXuC+yCh2sy
yemQzgsxvN3Z+sIrmgg0nov5cYa+DjuFMmke6A0UktQ+MfjDjHzB7jG0/r4MuPogqOovh9HgK7dx
Ij3ylXbgy8+OB3rRtaEw/eHqi/E8n0fv3diaWaxoLFYTX5e43UHJ0erCkxQGJRX8MI18CCG7ez2r
4uHAITpSW7xmOaYAlZSkUDRA+JQE1Y8Qfia+wY6Tp6jF7s1BJBtUK9UAVydrv1wfCBy4ocB1KLLl
c9oTlCMrq4r6cQoEStTsr0Cvm/aToTMhqsDrWIPnWIoBB4HmHEBptWtDtktcW3v9xtnNv94mENJh
IY/lIhhCziKIh7ll7UfqOl37RhkJ5Z4fiQDrQHE+drMfk0oe70a1FGxGq0P0lLlk5cdmf7yWj7nK
pDcYV3yrmvmNZ59DiyBXkmgV2jgcRQhe4jVbaMiQ25rZcB3aIf7Zj56fpKsXm2y0l/wAIT+zqScK
K207/y6SwrZcWjTcprfKQWAL+Hw7GCCGoEQ5SumcmxD3tLqMsgI6QAURZVCu76wdVfi7ZDYbXgAw
7pHOl5lL7IKYlXM65wwy72WcKlbRjOj6orbneeiYRYq8m6+I3rssK2SK5KGCh1NazdcJ0JwuseBW
2nxS6Ex98JmQMrkwGusNdnRssY7NetGsj4GgGZ8G23vC1r2PtpJxsyPsvXCSAixebO2jLdmKOUQL
ngtlIR9vWdl3oYiYK0Wxe/A4iafXI4d0VVUBSTSN714PArqGoWIRwb2Xu7AFUFdBWIZhlKk53ZAk
q8BEU662kDVjhDljrKKzTMA7Qbjhr78FqSUfi8kQu+LeMxFGqGY8uFMTtvv3ZUkwmVNwFBqx0+cf
59yM3qO/mHaXN/VnmFA6g1yBlcTIRMhyxYElao69gGb31IdEXzLRLJQ7+2bd8XKPEfK0IfoiZT9l
mlq76SOLazy9heMKcqP8ict0M2yfVwkRVvGMgAkuTib3G1Eqn2lr+a5mwT02ZklBFJZLpJVJSMo3
9DAUAEJjaGxVJA0AEw7Kz0IINTerKlky9aXYD/kekzttCcoHP3YqvYNkEKOd/hVmCY3h+uT4xF4E
Q18RoqTLbMiMBHHQ43h+EzYm6nZnYq8lr9xWGlnYSRWVmUKx2APhRNrZQ//di37g09NI+q49SOuf
8EZLl4pXhCCVbz93yIDsPw236oXKK15liJC1ibP0LjX3c4ksQGNZhQINr0yn2pXSxvndqQoU2LQ2
xubYc3sdgMRDLo1/39nFBgExj1NWZPuOJlTJQXvGKV9+8QG31xEExkmgj4AukQjgBKSGDmrAKhff
djLLPAkeKrrTf4C24XnqPRK0RWgJ5CeCrMI9mxo+fhtB2yQg3O9dbruvqlnotRlmDGGc/E8KcsmO
2fj9ew4alZ3ZQVS6Ht5cd6GscWuHF2sZVTDS7iJiRWvqbCavCVEvjR4h/QQd0iJcrSjKAOkLrIpH
fBgg52AzoeibGcVBhlctLJHW4vGaHcDrsFdHJ+v8JfE/aDsL9iSz6zhVvsLCB4U+/6FiL9Gl4c9y
uDKGVTW1MI1iubp7oSR5YbC0i/NTRIcu/fELhy2t/35eo8q7OmPoyajI0bw//I83x7XsF7BWCd43
s07VpEy5Vouzwi+HMrBMUWiGoH5jvrVAd6T3+/nqRVPZAujB+EaJml8g+QXSLFy4umENpFYHYCbP
DiUyoopDNlaJIi0HIrsmHhHMyemixZP53qyaZ3cFIqAOm4on1OvGFwnzZNa1t3ePuqjlrgtGLQf/
+bBzpymVRdPU7uXrkxiPhXjLIl5//EB1khVZVCwibCIKj2akpffbC5dQrd5EJT0iRMkvvQys50sL
ClazdhD7C97JHqeyor7VgsJLKOSfALLq8WLNsxdCohUbHQUtfjynNqCLEGbit1bEg8jL5RPRCHjX
6a1mO/cr9ec7LtTajnFqr8hAVN6aAvRDyYqEdxzecxTqiybh52YrQrwWm26bConlGPeAQKgVe9U7
mF6uNHb55CDKKDnub6GO/sIynBsqIGEj+Ha3YhLos5ytAqv/wFUc0aWrGexWne9b1gTwn4stMDAV
BpnAKBLtEMCiTnmx2nqE3Ci2UcI9ypm9+uAjevizFTub4CnvaOZQWGFEr1d2MPC3zpj8iKTaVV0/
TVemXWGh3172FNPAbksH3o9ZXAjkNDFAcjAX+vPPOXdRddYLgpQ5WDN+FluA5tQt7MCyugN6iEbe
TK7wpNwcagwObmrrzy+qywnur8ExXSAEklSWiAey8/KpB8O+WA7Qh3kAXalVTOy28KOHlIc/BvJ1
dpq/FLNAuHBgut3VIaIajWtD8x2z2oxtzG2mLsbiZ9hLFbcL9dI18hRGK3I7z6Q6RlxIXfvIxvIQ
ly2jR9oCH1QlyeVIiyyMUN1DBdQOIYaq4o+YCcs5kxeuHpC+RZyMmGQeqZg4oA88gosw7J8orYJZ
voN4J+PuSnOv3A8lLaSNZ1ML5CeP7KVv0RGqQSpX9Qp+olxsumg58Sj9jN21S24h1NJp9NCykrS4
ykqFGmEAOIqh3N3kCLuBOg/fmaovHL37pt+hrUb3fPQqj0VHfHLeC6aCBZSOdK1SWwcLT4iAvEtP
8xF6nMxYG5HQutiSpKikg32wd19+r70aU4pMGofZF8+O1xzMvCbm8bIaxjUXUIOdWnDmSjORoGEK
aqrmzCSqLnK1swhtpvx0+bxmRkTS4EaQKPg7VKk9CGWVTED9nXnV9G3Q65F+JfTHj83/3quhTrsh
HJTvDB6ccVSuLPMPErR0Gze45KTK9KuC/YZRt0LIBEVc/q6D/aAKDshxcuI+en6OwW6s7NgumgsB
6nwny62SJvP9PtKVZk+1FWWlYmv5Ef8LpC2aeLSWBg5idJYgINBGJ5CEQLkiW3ErueTrqV1K20wu
WGvRIff1xPK6QKj5L3DhBwYX8Uq5l27oh1lWxxYYlKtQggrK9tNI5XKDO/X6w2XZ7o/uKBKoojF6
JAc13PcZqEOxR4/AE9KspYrOekUV9l1Qv5CTvbEcVlPMIKdvgnclJ392G4UZDfIJ4pv/oEjO5Wch
NSjU1yqZIdESVB0NedJA5OzvDb5w3+arZW/zjfm6oksFcV2Po5U4r9PxdPukQD1C0fevOPuWSkZJ
VzQdv7B09jxr+PWtFNodRGvVeWk6q1zLDminroM9jDHfYTSGQBFjLO7euZ/Y20PJ4NaWb+ewoZcg
J7VJFd/H9e8L+xxD2+kxvitOI2IzLOCUO6QHZ10fgfeMJPbiHza3HbhNJhzWjqoYhW/KoVEJUa8/
qLJ5KmrtCvWuY3VEjwonM7zNoiAo3QmqrC7MKFe8c5M5u1rSF2WFaUvLGRny9fluurYRUfDnJDMY
No/dXstWGy+LjDk4SWP6RKPfgTCYL1r2OOmZlXeiUVthp6f3aV4KiqWzVydMAOu9M/NGjVJZaXmX
AsKDcgnCErDbrqn8ASV6A4mwFw3Jd4wrUSRw2F5QfCMeooE6aiHM8TmvrTYdTNLpfV4Op4K2ZIzs
n9h4l9k9xCHaeobgfGlYIWGV/IM+5twIsT3yBObYoBuCiZ39w5xACrQTUGhDm/9FC4yKz/8A482Y
1SXASXcgM/qOUrt0a2/0n5+KOdxKbxG3YabySqDpgeMnN7BljWyA3EbxBbT/pVJdH/DA7PvHewq2
sIE87APNLxTzLYyh1qcs5v2IpO3DlYOtcDvg5KIUxc3Y2Kxz1IwJn/fJxeeBZpXLROo8pIYdfQ+K
Kqj8NPp8aKfjgrG7oa8+oFruH3/2AA1vcofDb2zXfvsDbf/j3/cRkbliNFwAHWW3rerPTAh7LuTj
n9812DpWz0FYFt16ej1bcc4MnfmGB2nZtZDpcU9bzPrSi0TKilQuwg9SZtQqpYG/Yq3mBOJTkUMn
qM/I9in/RDxVc0JdXjBOFG2UTk7vLQfvKbacCAFSmlBzUgf08xR+e5IXxBsOgg/cYY7xEVj1/LaO
92tnWb0O1lr4Kml3fRxgxXrxzed8xbvWKUO5Fq5kuR1NMHc1qvg8ARCIYky5VDFr1RdkhF/Kd56k
PTSVgfoFtcaVzwMUMROYRy9+hZgb33JS6r5gQVT63kb44LfsiAgt+QAdTJ58bZKop/SuLce0K2Xx
HolYM8YbHNsVyp6DtmZUbNR9YoLQomv8FFrfWcI72TnMfF+4C8xG4MdhxwzftUyUyMIVC1hErQQw
N2zAfLFqYnvMdjd+9oeB0Jn95snvYsWBOTpwgLsZf//ckpHCKYEQX6xQR7kuHIbI6ZxRXBhwaLH+
ZpTMGIajaIDEqqQ7cOWtaGo5clsp5ORoaC5iC53TrXANIq0ZGCYGYQ0qfwSeesxvTi3UtlU9q9eU
dRecPDGlA2+DIsDr/aOHLNoq82R6XJ1qK5yExnYEo8GdYUkvCkjsTl6TFWU3DfloNPjYWcXVyW7n
bbfJ9eoakryhhR6xHZ7hZil3Z4dzPrLlnk9hbOUh7Q78xhSUyVJ00K8n5ErQrbE84JVWoK43uO+e
x57c2H4WE2gx5I98zG5lBEIyW23EhckQi8JQigRPUljI09JaXlIc4zc8FCG9mvHxmb7vI5qn+xCd
pOprNACgsKdMokUOR8C842tT5xLO5YC8ewv2zOxCQsZA5RF5ogrkBBWMIShrwFhzCUH/zPt1Kgxe
QGl+g+XVL+6DiFd4b7AcdxtghAP24Kktx/X0KJeH+YhwPodBAXRqJ0aeUj6pKaPauFBp2CBcAt/t
wRGuXlk0fc5SAhW+vAwz+QvrBqT7YC/6tIwfc/X0g0iKBQfcfdYAi9kAVAvoRIn4O6wTvo7863xN
VJC5zxYMNsXm7Kdklb2SsnHpjlzQK+jgewH/AeBCeYtOz+/inwzgO09g/dK/Ek8e67JUtLWC5wku
VGofjKSYqk8FdIl5BzMrfYAyYSnZwzraFxXkzQFyLJO/j5O3Nv4BhqLBUQawafJgJSi32Ts1jG5M
zu+GoX+4qAQ3fQMbevNDB/Lvw2/dAjCFFjR0sUPnJi65aysL6yHXhY2Gyd2D+ib74ISEAB+5UvD0
WTACfbhMIQFrqHHQbY/LOti0bKUGmvBlWWkPqjbyk5xsUlNABpKxVoVQyqV77Lqp9LfpL8RB8c1M
+qB6praqcxJ+ugw+U9KYhwUK7VocJZnC5QNHszkhsj8pH3+qn278LxUb9zVXP0haaJhxKwNOAdMT
MuzT+09klgsH2QeUpvdjJQzl/M7urAcAsizM5aThk3rwjluuYvTeRUmey3skLjyzPOytiy/tFtPb
Kmj4cM9Jon10VQ55MUB4k/rvLKvhP3Yh0+dTLzsxL6hp13IPD+rqgtA8yLnm0OpzKwA07wVvk8uI
uAQMukohDM1LuJDlYoXfNfDmskZ1WimHHbdFDY2cruPxpKQMJ7Z98gfAUFMvyUW/aMvGv0VeUj3J
Dxmy7kYShVvgvNqbG8R/LFPrTaTCPr0OtLoKZ3ZbePhl6Bgf6OwQ9xk1NIYB1uiy4acKlsKoqgdG
6jMdB/SGMO8MqQtwKKmQ29zBYaWWPvlhhZGzH61bZSSNjs8JriuCS8QyTKl8I0yYrwlPUC4Cc/j4
Cpj/DnBJrVSSeWj2zAdShG1pnWctiR5YtFO4ftpsbSUlwDjy1vvj14xziReziIwPZidE/q7p0EDO
e/rj14EowHsVJoSw6WcYfPMxVBQuHPhscjgHOPGi3JfchhTNy+nQgfoSTJv+iC0a4mJawLPIOfTD
IuRi/1p8BNcjWyENvyn+Ge+o0Af26n8gvJp5dfroVFxQm2Wl+XDKX9DuGck5X8GxhBK6y7hc9RgF
i+y8TVge2EjD8z7vNY6elNojVGllWl4V5n/7qAvtlN91hUFtRnOIdmqLI2jtYvc2FCb7Zan59/pd
iOmU03ZYkEB4y1muchiWKqTS3bP1YhXcmSdXvhl1Ll+L7o2BZsVV3U9XgK0JIv5XQV9gmr2AeOJL
gwI5OZJuh6rjvfk56phmVpYeNVZNtapNu8q7osqSjrRV8H32uSDrA9Su5Jpk4S6GokoaGk1wTeJY
ug1DvZBo/9k8i3cNUjKGb3Y1ZdGM4tM9i4zKhA7KgaKxN8DhlKySmuuaO4P1uyDXReMCLxhloHsD
QVgkMBYQ8/3QlR0y39JINet9BUGaSLnlD3aiBPofSqNVUbHdpWNeUpvh3ZQfq8s3XZt2oUBZ/1Zr
CW/jSl96t5uTWek6lp774XntFsE0Lsi0PpvpNSlsIukW8JWf6/M6rrIE4bgie68OpZS5lwL1evXI
JRFYC41HA+1TsKZJMf+yQHqyO1zjjQ7rXfk7efr8Q9yd6x02KvUP504Ic2KvzmJohPgIhqdodUSV
JwLvVij77FgvhANpCdFKv5AbEvWeQFrLHGxzS4GyUhhjARv0dQ4D3Zi82dTmE2xCfoYhx15aooV9
+PtcdK+Bs7A9YQLWNnNww8wxaOAXKMOApUnLCYO94UEB/wItbspfnSulkoIGa5E5Oq/k0lLM1DhT
87uwKyYil+omEPkgsEKppDgCM9hChKrG88IvR4wEgai0IA63DjrAvR+RvD3eo3f4rUJOTX2iAV1t
M4gQyaQccSnW8DmKvGzuOuDcVEntUDSoJna1ON2//hVAtWUHzau/WGbXjAxgTOfmnz5Zl7kUWzcb
AAprv3ZCaY+DOttFQfTUQDorWz0Hx+Qi5NW30/cpgrlvhJoeY5VbeA66UwFjsFTw1MqxHurq2g4/
eAyv9J1oqteW7jUOyooGihv6G08LxiNZ9YwZBv0xovT0ym4TnGNFItGrwV2pKGxvcG8OQSu8B/aS
qgIfYzu114olWm7JX6ksyj/Loc4KMsmeCGJm7lsSCO1QJT7Spit9cNWNCgDdN6lluVMcLy2lA9Vu
2Ag4n0vxgMZkLQ7BUb5DtO4H2JRh1kzttR6Muox6Cm4NMHl/5ORGvRoM595vaggNg8URIspUuRbX
LGti0v2P0gsED51b96t4ZROJfvBw+xsZ8IaljP7bL6ZFzRnCRAvHxz4d+0Jn3mpXHJF1oIV5Nz16
649X5CdY27RhLMpf18YrEjeD2W/u3j3zFX3mljDAbAl76i/q+7hKCkgQyAsNgsR6rEyfV+fE+c/7
VSvo/q3CgUE/3/TARlRhWkICjVX7457TaNqYhMZCuWVVm9PdIiTUzSNipthHpQBL5rLKMMFOZJBW
COlogm28FT8GDqr0oIGF9B5O1mf+r+6Q3ZOBovPW36gJSZzX4jr+7zR6n6MsKyKK+QECCKDfcLVB
gw1jfD6sN4Ku0aJmtrn+Za3oucSBkYn1ydpinAULMyVv/TOJ70TOopVPPND9+p7MyUF72AxYqvXv
/+AE8pKhVsdN19LopSz/hCmUPnOpQzzcOMe1jLEoOs/dp70DqrFconmRewOYrraylHeBKSmyVhk4
5D5q/vO/MwnJNExqtPB7MHvplACAihpoI862/GXGpQjzABmirqyZHLfgaDk73lVLudaz2Y6wzegQ
lLgVchJDIDOJGeO0peyhAFFhn+IEypYWaHnIgKw7MXZfTeH8yYutLGfdJMFlyVu00ZgtalXAlSx+
M7M8ZTJ1o+C3KY3avLFcMEahGofl2gTvoX7+H5fpI+k5QqQrInxjgsvm63c4GFOaZhjOXUQb8BmV
SQR6s+9huwc+0xMbgT44P7CUiws8+1NzgctCBBGVZ8ubMtRllX/pQGfI9TJrLtnYNMvFqDVgB5mh
Mkr8CpFXaBLJjp7RNTxl+ZhipgRMkMGs/Y/D0+3EKCOAB7O63Tljggxt7L1Flg+fCL7fZfKiC78I
4oM6c2JgxQ3xJJs5B99aTZVGm9Bp+yMoHd4MpifOzU8hb4i/QUgQCyFWOnc+ymobpbZ8E7Xy0iVY
J2kEHiIC7FAsx/yF75eKF4PUOZtA2yRQSuoeQC0IOW6NjCpp0clIlrG5vRKMiplSH0CNm2QbSvVG
AP0oCmVXq40FPlXlKTe3LhXOA8tMSPe/2hXEgqtpSkP1Zkw4+VKdPbJfogods/nqof8vmh49Se8l
2uTK+16r+GUtwSmhudr1GX4P4HKpfPmQSdzX7OsZGXz+UK5ghYJYXq97YLtMWX0ZzRJXudJBOXTy
U3rZRtySRGbb2b+qHVQcKUtxcqdNMjzaWEUsr/zYftWOMA3RMT/zagjX9omFSVoURMTlosQnxcwe
OuQ+0irixS45zB3ONSGtligj1VR+tusIOPtWkuvxuQw6g1QHeSamMi6ji8F9NG5cnf1GXqeZe7Hc
a9gjmy68HZYlmW3zf/dgZ7RAuX3ouVM1kxPf6lqW55inUzcZ85aFC0YhwGVbXrm7x35GUXBfv8J/
VyJswxMXKzyJEABlMQskB+V0li2K9O0lAZOgx6I5a29nmconXaczzMA86MKUZT2On02hStjMi3gh
DM4ASZ8JX6TRzeZKI0RWeUEIatFAZoRzU6nEuedgwrdc9qNqffFTELP/qmTsZKvXjw+BA9TTAbIG
91j7gIeVOsAE7vqpGN/aOu5CuQAQp3fickIvRRvjY4J6sSRXp8gA/4wKD8+lAxCO3adLKi5Zgeb3
chREBsh3IV+ckuSgWvui+F21ob2CBroRPVJVwIkbDCYNyigIshcq+a8XHOcllrCE2crV2CtXCfb/
aO+s/mNwx+waD6OXoqQRFq9/mOt7GiN4RjyIei8HG7rPuVfFNj5PU76E9tUuge/o0Tet1pQLYp8t
9T9Xd53H+wefP3Kr3Yr3TGSNd1daDOx3X4zaIKFiukK0p5cdbUMbz6ARe/rp++Jua4n+cpArX55e
Z06KOGbvanFnsNl4YJBDSJyZiwqB/Znfc7g2f97Q2nXTIePAgaw5K+SmeDyXez2krD7vfzA0Juti
nDyHhLIzag2nV8R5Nre2fNR3+687lyoXCRtFLEN+jq/JbDWGa/bVsdJLKjTEc7hCf5+cBQr+nyF0
LQSUePjm63SsH0tGmRw7nsuWplMqGJ252/IPsapb+Nt4422f/eqq7J7Ei6RHA+uiq+OGoyUJLJti
86ebAv/GgPBgF2lT6Sq5emQnCHxc1yUA2ZBg8fXA3Z5vfHQI4rQHz35T9Q2ah93mSV1DrEY8AV51
f99wOASB+PMh+xXhh5SEe3jVc3bOjZsv1CnR3pmBTL+susaf3Tu4YtSHZcq619WrxnSty3YSJi7I
dCNMMPofA5snFRQ6nx3aF1yQZeBgYQ0awDjJCD1Ofs3gQIzg1Y16g1k6Pws0A8xYqtwioaPyxVVw
wDnJkXRwsDdk7cpd3qzkVz8y678cz2t6horjUUh/6aNppY2+uWz5Y6VEf53acm5Em5xifkC781h+
cQ0A+G5nTJfIR3uIykc6S1KzAMIcQOY3j1Og+VpG9HgbQ0rbCHvJqWYLtCUJrzZTbxL4ezGAZoTD
p7BCgeTe0ulwtEduUP5R4yJm++X4PRirPIUUkhEmZ/qkYZbDXBdBJJl8EGpgizMvJyZTlhw6RmrH
ZH0I3OV3Oygn0cX4dwNuFTFAcimwbK4xeLImKn6WILEA+e8aXgsErlgAD/8ddpG9omYLG8KWO79s
rU/RTNtqcB7jSwPQNfxJy91hV8OPz8lks2fQU4Zkzz12wm7JFpbmcN6zwAspf35AvUQo4G2CPnUG
/gJo5xhB4gKAkkSPtHCDENfm8vx0rG5+HamOsYK3Z4gujyRyxlRnTwhPb5q5Ju5/TlPg5TXgZ1pQ
nSYbQk5AfELVxmMubISvk3rnAIGFHDC80jrWOOdvPEpNKF1PoZ78+PQ59m+fsqG3O5tH5Z8a3rb+
iah6xyaNqc8cQZBDGqWfx24iolyoeLL50zcv30vagY6SrZt8IpA8SaFL+66RjPDXrIRWRmXCE7/f
K6LrMfY8NH+JwcT4HjG5RSj1m88sIAiXpu18phLadJ7AEhEZeGpjzObYomE6YdGjoz+2RyrKIKJV
fOVisibiJRywABYEoyauHHQwSiBN71vmdqMz5/9kpv7P977CyyRScaSoG5hflBUmx/7/crqnTuL2
4+TVZw3UDVGucEfeFaSp2B8VZjETaIG8KZ8Yw0CotPsayEpuqFcbkGfrhaZKiNGzYA8bkTw8Tr6n
Az3BqDqeP2SK5Z5ZizoBn0auQOmFNxHajqoVFlh7VFOX3v5dulGFE6oHoq1DAO6Rpx0U5hU912e3
nxfwyikRvGWZcajn5MVULdwB/s01U4RJ8Bfk0dyWKJYjOpXNPmw9t2JZ546f3O9V6WJ91M76Xlx2
Nw+gA8lwWmDehbMr2xD6y/XpcZqwjhHz0K0freqdksqzP2Rf/H9BLU0fO4G0z3MM7VjEbDceRkC1
SO6RxHqT4jIKEjInetRo88eLGmDRh88FvaUq76DLkPW3MPeop0jdaCRPGLEQfyrNK5EOjCdvrUEf
Feqz8BDkAX7WCToSeMSQmH584J8b4ttaw0PQDhLMxXPmnEN1JEYqerU0vDJUxTDJK+fgovhk/fXU
Tywu8rpFoRJFYTkDUCVUAfQruPuToFH3j97oFqYNJojbSNUyFY1O3mhyfWE/ejEwlZnNicevIun2
wRD5pQLKMkF92xZgeC4bFc1VRQ+Hk2oEHCoKX9FM7vH/c3Vi6lul8dVNDIEa+GZDQxquWgewW/kK
s77TMisuBUqhJmd/egf6R5QlyoR2kx1xzm5mPHD7noo4VdtgueTDIGLcL9ofp+DZqD6wuOpj2X0I
L9/uKBeQvSFO5WU099a40APsEVp3h8nubupiRKsxlUurYfqy/IG/V0wKo+Opw+XVAUGMkn5VcJ8G
itqLeYZj+GPLnE+dJ/0watKHD2WV1bHxd0ZCrKcR7r8sSRjbFgPdvWc4QuI+WvELXhkcQiYyabkr
jsH3MHAbXfyO81NEVtST0I484JWAPprpMeWN6yCLRMCyzNONJKbOXlk1NOlRhtnp8gPm2ltUoWNe
boaSwnPWZNA1kvL1kA8Lhmcew4aa2qjZqv69rmvvmr9Ba+SK5k4dozLEVMbB10lr9WxBcvK7Ubxv
ciuXXhrLhiEOkFPEinMMJGQuby7JsPosSWHlqtr0MukqlWRZdIp6hHDKIdBKufpUCP2OIMwzo48k
KtRhWlkuAd7X6Q6ued7JM1GKh2p13AsS4ou9NqlIEUFLfzecXW4RXOxpoNsiMiJeNjhK/RvogcdY
qxvtlw3V02S89vzbrgpv8d++7+w4G8fna7uT92KmhaWDlLcwAvc98Csxgy5tGObg2O+vuOiCTTL1
M9H2N0rj1Tf8A2bCqKaJTNpo7D0EGwIvMIYjVJ5vVRUMxohRdLh4oiI0FYYA3hkjD1Vvgm0Fy71h
BwslzilVMsgMy3VYXrWGerb69IRdGD2UeiIGHJw/OjtkMNOBL7SNjib2/wfPmO30KtzYfhySRtJ4
B8mimHByHNsPz07FCJytZq5UCN5EYzgP7vKu9mSvuDn+vD2jLUfKrwnz/pLdG6oOsc+xKgovKGxF
/mFZpc6toHVwFKusE4m6+Ce9J744DfjsEUngGiGv+tA2JPKqRF1n4yXh16wdB6EJxq4zB1xT+vX1
5v3DeemtF+lMdigW9rpVRueGxKggLowPA55exDQj7g8gkZ/+Ff+iBLRGeQcpPSzc+0kjtKIXh0o+
uJEW3/joRlCzjxZb/ZnLtBtvOUOyUCCV89Eo0cbMzkrUyYnCpq0ZN9x9cYfkSq6zIt7qiHmdEyT1
3CLed1MQKYbXjhiDkof+3zczEP6Qx3AsTTMeLDno1dZ7Ua4xBV8GBUCXPUW4uICFiiRjHJ+uouli
UkKRbs7fZmtL5o01mSzy2+4VEqdvou3UxcRqsRd9rJ71uNduzHmnN7nX0QVE+qoqkbbc7xhbjrps
OSJDJueAIYbRhWbc39IFHHg4EU5lpWFMmaSCHEfCB/8iTv5qZ1pHqdLdr9oq+TcqO6ZwyYTwPdj3
fNo9D1VdBHGwzxUY+qnfQVkaaW81WZV6dWl0ImIRyGjdAUSnlE9vps3c7GzbRRRRyOH8lpcYyqV3
m+frno1JnSh3tIUmxjF+p1aLHaHHdDvVr5+bhkbPnP8Y9aF3ZVjlGokCnLBWuc8k0eWqS9u1/6zy
kWKzsEceVJ1msw/b7ZiAJycW9oyT3AbEUe3L/XmoEqZkW6RofIn/Is1HJbTFxVh5Yg6sdkLvUGX5
0yvvCRekIUC6BOqa9DlJaHxMfLF7Qh/Zb7wX/Gg3lvBNyavKM/VESM0XpjpGlMlIvxxUpCtdKuj3
GuAhLh/OOPO3Btdo8kqf15uP6V3laxsXq7ZPHaFLjPAVs7jhbTlYYvM7DFUrxywmDVUYYvjAFF0S
CfYz4tMu77dH8qv3uq/S+HFPa7l7Jp2Mi/6EnMr4tzb/X8YHJlWKYrRhdGLIjPnrGNsR5xRhXh2Q
ZjWpghrBcIpCIExc+B/b/wjMwvhUaW2VmRknNqsAzyUczbWmobGj+SFmpljeMtfRyy8PDI6qVQ8T
ct2t/wtmhnI8imcYHwvrYDMOtUxpu/G3tmRbGXotiel8c+1XbCd34faRVjV6C1H0uC96VJ0RvV0R
BzQ4z/dqJgHNu7EQf2upW8EPi+k9WbCka8G+WEefrR8LqLWd8DPY1x3IYdNJg9kBfnBxicQnBZL3
jmF9IwTDMByaNnL/A6YTOvXL5ylg1U0hdvOCx7vBmdsb+SmLbZ15hw7WfPhzeN0ieXUROnpTTlAL
pT568FPeKGEJYqGRi/+5+xJZB2uGF/YV00L4ifRjzEHI0lhIxsqDJQUpWBP30CoYr9H+Ey5DB+K5
s9zPpbvny8odddV3pd8JJRL4jVCXCcilZU/irDCdSPHtmE4c+Ovm8RIG05LNDGKxKzxx2YJGs9DA
qB806Z+9cR2b/TDBdsriIMujOywI6W3vUU5Vz3yzKric901FLu/6deBtMA/UCu2fwEUwpb8gQs4W
4a/gYDsF0ckupu8OYe0iSrfC+5NfA99v2PqdI0j5T7BbsqYUjK7QKBSdfJdayg2Qg7LenlfB8HGF
AHa4Rqw2k9qmEAabbLQFdcTNYepIdY1R7qIOVl4QIG0yjAI8GZ0FUoBPQWkaFu21NRqBFDIoKwDx
a02LnwFEF4coXsagD+8+FAMISu51nEM2lIz4TLb7tcJNeCZUkoeaITLapEbLBp+tjKhAfG731u1G
VRy4FMuxuIjRZROl1gWR40Uec9yQGu/EfgfgXf/MPE0y8eZkYuuMsq1iS9EYFt1Kg+3Jyylw/G9h
MyzjXgpejRU8xdJPnCXYFplSF3yfUuFDJjgvymHCwvvKbOeVCX/rMEKwJQwFbHs6aHV9nksak7PB
syLzMpAwz0YsWuVmgBz5hZlsxG44samAamBWg21M7baF8N5iIXERm+ftdQlPpQ1E67Jp1Bqg8FsH
owdu1gtr/8Gfg5K60A3l3T2qah7NuGjLv1PgB7B9dSLWo6gJAb43VJ6ukODZIAfHj5gjO7/B08OE
ZzNlUWHzjgWOh5GIBiv4oqRZEUUFoYnLg8V2Wn3vEhMd6afO2YJ7VEv82dIT8XxatA9aatAS7w6z
sR5MmjmASppxJPbTTOt4Ynf3wyB6BieJYtTaXJNa9p0qcshCFY5NgalhYj2kQ6ZmPAxid1ERP3s+
b9vlL4w58YYzVQBTA8+Rjksmoro3CiD0z4yA24YanuHr+kGPXI0drVPunPIDl+byChuj+eYz71MW
Xnr+yImqUWdVphkY/naR5bFbh0Lxo5f0gVnV9IaKva9DwUquRyb+S/Hp6flPpW5x0Q+RnEaBZRVc
/ZpgkSOxSY2M7E3mGq4+1i6fFr4ZClUiP6jv5za0IQfF1aVtL5c5rN6VtyeV18wGVl2fGzqxwixy
HDgzQKcz/0IfiT7H+pTE2BQJPiGj/gTQW4oVPs5euou2C1UU4VHKDSSBB1aIKCtK5LOZtPBMH7E3
nRb8OZ9oN0sw+UkdVjtT8nc8vNSFyEmHvvt70AKSSSwoX+vvFew7tHb0Qu+XKWKNdULr7ibGwfhL
fGbHz3hF4dspp4Owsoq1vUNdg5RJNpHIQyDVhDkSmKy1qqLheC5S1fUYLUbG7dUCRcZI6ULQ0WsO
r3psRXCTwQDMtGT6vDpMHi6yBEpLVM0me8NVeKsppwh2f5OvMuXH0U8qxKAV9vM22TLKnTFhTCCE
+ojQcUDc+E6CsbRR8AoYqrZP+ok0ejSM1ZQNdKkGdiCeVYEP7Pd3zeKVLaNRMbFwJxTWuFOMNfLy
mS00nmnXI9XWnItasw6rl+Q8OjHrtNyV1K2Xg6tXRbwMMeH/Xp6OFR3j6IcuGuxOS6sbC+7NjkIw
49HvMq0Sht89vbPqQRNY9g/NlqG3CtHna2bq6PqWeXA8fTecNNkAZxruTMdcN10lhHBYKNtdumB4
ulrEm5FbrmilO+SxVmkcloZrP8e3t6cqq1w0I1k4ycQZtdVfPXr5xKV0dddY14kBoZ5AP5KtmLQE
Y4TFPkCPR1Gk5RrTkzcMvR6GV7ugNN4MZXKOuFpiAltNVGgpVA2WPe8Deg8PSZ/IoUYBkMgtyYuI
8/JIm1de4G2Qo6AetYdgkPI/UF/TGgsJlk1Dp0wSvoqY2eK307zDAq4fk+hb/HLkWYkbC0p9jYkX
Rq2P4gD5e6hi4d98aoB6xEZAh4aGawsOzgEKaKsY3Ot5Z2JILRIz80Zc7T9aXF66E5egF6+K6YGu
xwDp+J6Y+RnI+0vPGegMYYEsPznlQJCeuZeJ9UPrpE/NS20/32byw3ag0N7oIymlYEuQ8LERYX+u
Q8ztGLwF8G2xZcJkzClDrTVfJ7frAi/+u4RDDpmFx+0qZrHqoar1ymxxcBz/HdrxuS5Vf9zcIcTq
iuObA36N2ZWMlDwgd/64+9GkAk6kW4RGFcvoTapqzauHRNIoS6vo1eQAm6ORgEhd9HsS95yR/x9N
Uypx/wLsEXE5FxskPcBUV0Dv6HtZ5KBeQWeFgVgSzl0kkxjhhEM2B7Wz9ryVPmd/0X8ngLwNRzzd
Q69knpbupq+CLpZ9LawBOaMaAfuDNnhNjIO38DPmLuRIebD714JPYK00e/PtNwMZCZZLh4H8BG2f
iUgt+6W7XFOp/xxsSh2+WlFtzCiPR+yEvuRp+VBCb68XKQSDQVxvKhuXlpXHIL6RGdodLYC4Nwbj
FQ0JP/fbBzkqT5YTBH0vJ9h7/6ETBZFaBRB1qaRXswatLwB6zXlqhNaCAqMQdnbmrIPvjQ8+4jCB
irhZY0BanhW6fQinsnXZNsqHyeIWVIzNVixJOZ3rwGEzwchIjrCH7cOdG4ttMhIzV4yd4xvuD2mF
of/XfRsDwD3blH+AJSgvvhKCuKLWSsPrPhYtUIP+VxcxDtmto5yvKB0/zxTrnnI/lgc5MUDGiJ6H
TUiGE82E75QWoQxwRtglqGZKiWooOWUmMYnDObD9aDx/NmPfX0lu+seu+dicK2O7MeVRHkvE7Qb/
Hwfkm/dOLGaV7k94vZnT6ncUIlIaUvS/7TlE/nnG2ZnTX2PrLLNjjJJmiXAJPXJGmLi/H3NG1q5J
To8kIezfvrjSloBXgXEcYN3y3YKD9vfBKMdMICuQGGR7O2lyjPD5RhgOu0Ap2aKA/o+fEQn7YIcG
Kf4OVvZjkOgEICud2+P9kRXWzQbZSDagu2GJp97Jox9GtssecrhLaKskLOym7WgDUCs8w46kesgj
bvSe/LFXjxMYoIBHof+gFtAq86usBH4WbcTwDU+yRMZm02DJBrrbWpRUYCZalahPLDTFIlooNrNN
zuuysrUA3yRK3uBizFIdeHrLwVFOIjojhllkmpW0v8v6gr4mabvbA1nWZq3Q7IT5wSdx1XAaY34i
ZBlclVHD+UTzKS388iewbbfta3Fx+GIfUGUBusX9lRfz3blI+zSGYXBzwLvvoZ0z8EkrTJTxE6Ek
cPsb5ju/i2IPLw0TGwcy+LdGzs/+h9Qhmp1B1C1zhDyE2d+b294JoxR3dddgRalmePUPJ9xVFKm0
mxYUbkNEMA2AZojZTeaBo/JkI9dsPTUy7QJlblCZnz/WdeU5L+0aTWEN8VDRXdMoHGswcCPVcf9m
TREMR8Xr3p5Tk7kWHKu/qajzsiBZT9gwSbnBbGkJWd9GJT9pMAwuW5xkvDInmPP0sd9wLfD/LLi5
vc+KSDz0lF+9/66N8uRQDlGVWeXQ65u1xmL4VJOGXuzhyO9gchsDsy18BPXotKy+1xZbJEQgxjlT
Sz2iDDS3MOZ8x8kk7sf+hjZfTQ396kRYj+4hrDM72t53pLj8JHAgGZaKQbYzacWps4ge2fm3DWIo
6EqfiSK8earuSxrAJrVMfCffMCW+zXkIb16IAdmeCc55j9LWoOMJGQ9z+xnuIYji76OTOLolYDn7
DnUVMGoqPLGhOHabStS/n4UGJa+jchIEQxaQsbUFeircqbmtWxjCi9uVsG2IWfZv7asouPvmu4wm
8vQ0jN0Z97MuN2G4AQA0Rwqn7rP0BkHpHeYiQXx6pXXMRf9kr97w5h5BTqZiZctIikMCu6flP2RP
cO5l0zYekWRZ/YrEQFhN++1x98AF7uCS7vMdqcqqOKApeXUHpw/e4lOO49RpDsWZ9kflUvocpd+a
4XXIjoF0pDKV/3V1oGihb/np51D5j4yXVc76wLSU5JKriYo8AEcLnD0hTfaeOfz4lg6bllWdHHae
R3Ao4NmVhcw26nTf6mphSEs7biEbLAfxkJwoLEUS92AXmIaOIXXE73jpgbfazzSeWx6+vvDLhyU8
ETDSJTy1m+f6DRc0CUNdvaCAUqAeWQpHqC3L5h0VO/eG1n/FHSnbU3ONyp9T7EV6FmlTe6aDK5Qq
eULz98YPUZcV4pLgbTVMN6BDR9TqOX1TplUoy59+Tm9JWRRo7cG4KVtcdbX3yu4CZaT84ngIqsky
W0uMqmwkX+nswrh0t4obpMHQu0yfGghhsACofxCqiRcIY6sKeDCz18nNrhysV24KJfu8WolW9Fxp
nOCIFK5oHIWOXq+Yd7oyQzvbF6Xxc2d2GxaEhCDdvYpVJ582JZh7oktJ7MFsUOLqT2Df/QHpF2Vs
xzib1D8sRU7kPCgKBlGQKUXy+461nYTzHvbjEfH0JsjQKCau+btkxZ0j2YKj2vEQomQ1aXXhHvH/
wdG6m5PWvUQVLCxLbc8nIZ0R7LTHlGANIBI2Dto4MUbGIWZ0xvf6isWcUcdIdP9NFSvGSrETPdb5
WS8lNzGWJ0EvcdxktDaxd2Az6ssSJNJEzXPHJ+HaMwOT9YBknW/3l1Hkj0AMBeaQ+rY5Dj5+Nopo
0wEcEL0Z0aSQdQ5jn6veXAKYbTGTX1iyRReVTXjZimzDaX8iPTPxUGiLX5zkJm1Onn3OL11fFL5T
Up6IJiBJuu6yegKxyAt/bYvS2pGA7tufx9m95Riic+R7wigA4gqwjVcHO3eZv6zvfkxqidFAvU5l
OUOiv0guf/NcRMgxbgow94/Xpow12JD2vsbyqdzjtXsf30N522FvEx7t3q6ci3e4FJi0cBsk99FX
aqL3QrpJpJdDB2bQ+ddMjjJ22OiwSmKe6RNH7hYb30ieDmswO6gml33c8vrCRMxV3h3za4rVs7Do
4VLDOLOzNyAvnOii/s1SapTgGMh65D5a2hg7usq7RdsCZUtAW8Ac+iOX7QNZx4ti02Iphc4IUgnx
QcbnDBUdhuIP/4MU01CnpxSTy7YoBx1lartfjHFmfnq3g9A9Ixo1Zh81TC20TA0kriENK5nN/5y+
8RsdIkCrtJ66nzrhHEovTxPYhfJxPEvdQSNPy4UdAJD81c7a/jU4br+bnLQl2MVKrpoTWJJGAZz+
LA65ZDVObO3u0Vd62YtrKQPU37g6JdMKpb1TXKKQhq3AcclYtHcN1HXMdLnzkI+gZZXGeMKOlHH9
5jgo233J8CUkwchbeucm0kAt1WuM3Fab0jk52doBP/ICeVk4rTLmk2u09lbuI0V/sQXr8kJ2jB9Q
/4hMAB4QtH8qQ+FSdCQ36YbJhbgrRJ94rXzrs8h1GHw+UIlv6QEd/TmTJxIU1RHZGB2oglhEqjvs
GqeWcW2688tcTE+NrbIOf8jiJv+bQfz2a/yrkGT7eyF4y8DLKEF8Qt4lc6WoFz4lM9or+8REyuEy
Gmdg9fnTZsun7V2ofPzBpOhlOEYwNucEEsqCdgoiibH0yFUFWJB/Bc1ptlJ3qaWPDUMwy7MiX+wg
tXRfpUxE2XJ3noDmrjfqP/fsXMoaG7iKQrFQ82lQDB4ZNZRoBahTUOq2MZVF9pjuV96X34M6eO/h
E/1FK+W3yFnqh+J9n/jz8QhQGX53RRd6fELpyqBpAVXFfIbEEwyaKD3CA7TvZlAB1SD/STmVwCYi
hdHFXcn3mPC0nKrOm+XsKqBM7ISyGpROdIfXL7eiqSl2lCguLZxNfOX2Mid43vonIBN6Zc/dXAZ/
Xsw1XtY2y858sB2Z8U1f1RzVxMuX0k42aGTV+0w7w5Fh95HqsuAs/FHP3rkX7+BcjMH5Kw+Vx+db
z2GtvK0ieBBBZrhNULN91u/1PdkaUx7Kjc+DEKJ1EqtCQ6igkprg8bqQUJtONJfjd1HYQ5zYVqkb
utXvC6iCOp8jQ+Y0Tof4oM57GzJZqNXYzscF0Nrbi5NZ3BiZfEISaKU1leDTQ97BNDkqbMpkFRAx
W9T1CJV8cyV89eTrrRW9M+Nl/p6Kf5lGI24dsSUcxcH10RnaILAL9thvf0jlmdkT7YZKnS2Nj/hg
Fxkr6kZCqC3YGW2v/rVKU612XncI44L+zwuy9pOge06NaRXp3GNOt9eX/FpoGIeM5BwA3op2Q1LJ
HM1PKxdQGUxqm/DlPhKSy0tmOzd9gIpiB3XtJ5TXR5CPs5YOIv6ySV4WzgLgf2n5L8Tu3eV+MVxl
S9BZNtwTAgk2CoA6oeVSyijq9QI5GqXOHODOtxwg1OCufzrR1iNoqGmrIRGG2CHdbRAC+kbrwYQC
Pzhy1uYKvKnQFXzkS4h6fhYDfKEY3ApMRP5zK3R37TwhjVt9ZCr4IBsjGn9wzXUlcDJSVibm7PkK
fnKeSj5daDOJ/Cvz3IG33HAgd2nWW29gaMHIXcb98haiC0u3+cB7451VeGyc0D/EGK1hUATauT9X
aZALPAJWsjxJFHAU4sXrM2qzMK5Xir32xzhBjz9KIHyv9bANtLEwY4g2r381JEjNh1abdDt7ku43
xZaG/HOsv3DmwMlxGIam7CI/H8q3OBRmD9BoVkrO7+RuxrPbO12W6qLg4mfZG7K0RUcxAMD95uvl
TtL60Et7YfiMk3eQpH+JKAC2W1sgrmHwsH42z7qlPRwwPywuaC9yGRWN76iBBC8k/P4FaDNqORQF
tvAOFYABl930L33LIwcpT5tlwHEmcQG8yNJ/WD7I2ttPv/W1pExzQISRVnfDAhvEhcAYOUyT1+AZ
P1WHwzCwgvFEivL0kGz+ri0/6VAHjrtbZqvj1wJnOINhKsWWcCKeM2jSl+NlhKXiZ+DMTYYLcFhB
nGfWTP49D7ACdc5fmWVx2Bjtj2mC6X27yQdxO6qJSpbzx2Aq6uMw7MyZp0FMUNazJaVmw7ywR4KB
5O/vqr9M+GsYnOcAFTjkwoyAZ1s3Ge7fQ/XIN8pu/9Sb01KGAFDSIMGq+7ZsHUqoXDmdK6l7lwLL
KbC0dlAMTp/kXtLNvJDrh3AUBsfRi8pkn6Zr8TddCPk65xyKuKi+1oPfmGH4kflW31r7sAb0yNZc
fFsjNCA1u8+i1GlO22D8vglzi797rybB4VxVV+FS9lvZhajDbsbdsbxjVG4jd7S/JU7wxNxhzam4
h6A7MCL6DHMqGJ/2KTB2qyT//ZYCvIioFk9QlKlSfCur/KLC/6S60kcb+YLRWbi8CSWmF3xWiZkR
ppSjo5kQLAkabQc9hNDH1RvT+LDRYufTETD3MAMabI1V2my3qe2h0zzbQ7ZXwAGhEoP6QB/9mkpH
O1jYcu7MjDyFKnfj939w9dPBPjTgWrKnEtbh56aWqbb9jC82XPT99A8bWep8Mz9j44GV92vMpdZ1
aKRs755QaX+pdwO8LMQBC+E9UfR97KfXfI64bLfenkTwO/7QUaDp7op77eLZ3d91i5oT5l2TkLTg
9CcV2dOnufZ7EHu5jGDeEn4Veay/5uaYmRTne8CMfMChbvULk/5ZA6SgHaqSE4J/hL+FjBtqqBwb
Z3sEBLVpiTysBHoTpRr74NznxoEj7TJ2IU9e58Y1ovVhFciXfir6PZ8Nj59eT1xJPtjkUHxNQEzs
nxUmAFXiNeGHjhIly0divjsMbX+rVI6i/J7f/TcuWPubZuAMFOQv44YUyY6W065lo5R5XyOLaNAM
RPitX3sNzq/T/oA/o5TKh8DzD7sn4FPzlqBqrhphPjpHTHRXFEynEIY5ntgSQmPg8Q84ym2zBRRA
8gC1bPmiVNbY4H21s9AcSdy5IfSXcqQMemBtv5pMneYEl0DFv4FsXUS6qddxzDa8OPL/BtdtIAsH
uho2KN7VGSxwtMZETHPHfntw2kQl3DMKwPtzJ6xMT+7c5wHAUgdCe0pjwA54k0pv968sPgR4cJHi
w9MrCCJE9wmgPFLwavekJmkOJ7LXxgJnpe8W3mfrxcnk1tb9e5npNbX459RoqXSv6xgdgT00rJ2p
MZmS1kc1WbsYEpRKfI2xGExsQBcFRRiZG/fTcvMRLWhZ5YO9HCG/W1X5/taK9mw3VlcaYYZ3Y1IN
cGXy16aNTycCCGusr6bQwv01qsHd2GOdl+1siD/IQddHPGmC6quOoowEBwAk7rAcb9b/GrflrJU5
2a/kA93rZQnbcZNYS2pKfHPFXyVfVCVL7bM2NdYoZBGc47oJtyBmVyxgqgK4z1cRS0J9mkDbt/kU
psQhhw7pVY8XMiLn9GkI5cchaf7S9CWOqaBydsWSWk6mw2/73dW+J8D7EfcrV+3N1Cyug07dnQ2C
L8UAfX5JYvrsdHLcALzaq+vVxihn8t92vp/1US0H1i0ap3PIKu5n81IPZoDXUgcT3OjqWqT5D2Q3
L5Ug9PA+o2w70MRfVDhnKqrdZVMQN+Z15pQUNkL3nshXvu0pwtQV1REsq7Q0Ne+o6kgLN4gE0UDx
FfTK1pJVK1k/KIEh30MQTqorTXdp9sGt460+w9Y6avyzFeaS/LOYODW8fjNemduUDJjBYX82fqIu
p+/ZPt6pmp8wFz05TvASBq0M7R/1H5vuX/EOmbcYPzgQWCU9aYHgkplz6Clwh290nR8B9ipx3AKc
06savP8Hjkt2++CNE7mUL/uhKs2wiPuo46OmTRLYtKCrxoF2+xRB1jlTX5qa4o14jEDdCcym3oHT
e6v5fF+iFfBmwMFMadVGHUBlqFTUt0FI3I+tL99dhL4hV1RoTRdSX+c2RRN69fi6VL8ngTp1LI38
fyw3hDJPrEXDJ3Pz+ULyH09Zgvh5GByIA5GazSGdo9SK/Ws3uOcEz5hAZ25LWDR3ioUqlpgCyD1o
S3e/RYUgvBhlf9LweIsT7pjCVG4zJAJTEY8FkhDyamqQzx4MiJ5uLKHLGF54jNpkcFVViCtdYuca
1D+WsyWBIbw9/R0fdQuCyY7HqwFORgakUkSR2i10ETuG0FjL8aGFReS4Oj1b+DcpXaThMPfNNfxW
oSvLdg5KJ2TUUKbQCoq/e4HlIssJqR70fJ2bL18YkQbMC9YR2TauNT8RLAICeXiH3gmxO4Nrjwph
k6AsifUn2t7U3FiPHWuPG+2YFtkk1GWMuh95PemoFZvfYgCp6bBvqfI2UGlRKAAAViSwSANt5hHm
4Y2VBdOuhmLWfcU59C3bdiAfvlWcaNkM4SO5kjOOiRhTbZ42RChY6KrqQOx8aOv0rUcyn2M0stKK
I+ibFp7jbiB1Dk9Hfs6ZKVFGY9A4yxWr9dIlOvJC4BcTXNM88fWTUGOOnmi03g2eeTH0Tb83IqBG
K7XFQarkU+mPj90sLmZiSzr0GTtM1ildMYhuCc7rEZ1xB2qLWgsNWg==
`protect end_protected
