`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cI66OANCJw8fIIQbdpCG1eUZiUrVUYlTNQ823416CUh5RU0Z0lUSscJg0VdsbyeOG0GIlqnKKDcJ
g+441OyZKQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UgqPJ9i9WiJwgzx9hA1QFTAyJQbYygHQhueZLDtbtfbgNYIe9Vf6qQf08t96mKA1gKActJ7BeV+K
6uNMiJfx/3aUXCSX1zJ6wf3n++OQDmqvxVVq3gnHpb+740+sx3yxZnt+NIQn5YfqgmEXSODHM65H
T6IlCQG0Rk76FUmssyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JffVUoJGoNenA9JkXMLk3KS8XcomfWAzcMGUl6pS4bKWUvYmY13D3pemGWR5ICLizj6/IEASX4qM
MrcOHNOZ78VNNGbrwydnmhep2T8HUJ/34A8F6RlIg3EPqaoJseDBIuA+1YYmvMYUPXWmDmWnG1uq
4OVHNHuSMmViCS9G0XZMw9OZMd079W0WWlGjxgCIsCbTxgr5NySjw/l7QR6gLw2PWlOAIibLSL/6
FYbf9Pq748eBFOa73RMaFJULQdNMNcUKu7XbHElWwAbBAEQETSA5PY/T0Ovuh5VWjxfKceXk9gE2
s16k5nL5jvgzFecQSuS2lSlURIB4qY5hje3ZOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6n3r5uCHMurGEnMpYNf4UX/MkeElsrXqvd4MQdfthvZDOuXHZxcs4tSf3laM+WPFVbsOKpN2K9r
vOlcg4pO3R/XBxH8buk6fx/j1Txb83yD004eikrbAzhD/XMeJoB+vwnOXVjryL4Tq7ewJGiuFj3j
3aajz5Netn79SPqpagQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ux6EQpdIiEpdxg0F62ecUw7+0Os42ovKYC5a4J5nt6L0NXwWYNruQn6thnH20HG3CkZMjYPVsVdV
6fsAhKiqralBKaBG/Ej9eLWDO0kqJYBDBHDr1KxCmmsfP7tgcSeensV8aAfsf43ITwJDMIO8VHys
LbnRxuW/uncBTBd8BpuuF6FOlCwImGuVwEh0SYaZjLlAA/zvuQGePlYAraOXp22pKz1CICW9YEbL
RHIga+6SQ98q3/eoFGq1j3ZXVJuLYcvW94K/kJlph+VD6UU5Kix62jbW5vyq5E8KMpqmJr9NNRFn
j81j5XKXBOZlfp+VVqMs7Hlviysaj593wan5HQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62832)
`protect data_block
td5QFuuLITbKOtkE3oI0mLzB/U3OEn5lA8+gSvm4NzDgr1xoKZ6KXCYimdZuYcgLb1Oo/1ycim8W
PFfdiPDalf8RhWG8Bm3Uye1fGmokMIeViJJFpudOlf2QwkH2Q9nSjhByWCvm5V/7FzruOcyzJZl8
uis+1q6Ca3nhUQR21H8IcHbv6Xy9XdyKOtDQhDkDGI8SOYvdtcIlVOvSvgg1PlHx6usdcjRT0U4H
P6/B+j6sbCmxYTaRSW+MrSFDCMABIOsqlOFl9PQ33XhNbwlnmHhR7+TVp+HznqI+LmuIQWc3StMC
FLXQkrxIvNX7mEKE/W9synmWVxp9FuRQ6tuVNg8KGhglhiwD7f7G+wTaFD3D4g8wczI7YzhR00Ln
P6G+1KyxxbKgHZ1w9X8twlSaNz3HwkPr3JM0Bnm+Lek41ACBllrIwOT5Qk0wqluVuwqkmNl5frv5
QAFQZMqozkW3gqe7zePnRIDY1hQAMnhKvsb7f9TsmZPXLSkEEONCx0QeISsPedMzb6/Bv1gUkRpX
iQssrnGxFh1qkivZCpbAac30BahF/epvmW271oRt9Tfn2PS8ZqqTARrTZPmsWZUWOMq8EQt2B1uR
OBnn89cPyi8ETcHQHey28GSUgueKAYN1DIibITf1aKTvmjTLLGpTVnB3QpLju5LsKfqL9l+lWrLp
KPDYQFePZXOxj0WQjtOnDLSIm4ylALZEyP4ue0y1PyQ2QgnI9fFDRnZt2Zj2f6NGPp6Z/FWOGZlN
br7qLVaM0AUHYlo8/hSZda6b2Zu9tlrGRQ9aNoIVsrIJURG1+wVSNPd+dxwxxDssTNzRsbBz9fra
+i0f6rporVY3QHrFYs+LV4aXES0g3kbFQSiCLtn4R9QHdUP/t0wwyvAReiJNq7nn5tL3i5SeA2wS
Y2ZpaejPRmwWmkt2ZaoJEYrFBWdIwg/rHt5pLKo/Ab9O/GRUWWbLIwcBidb2hcq3AnWfuvB6SAgy
p5bZWOBXby17vlXoFLCVaoTGBQioOOrdj1pMzdTyn5r5gqM1tpRiaDArucIbqyYRlCqIpNRYNfzU
BdacoKcagOCiBigk3b6BvTBg2IzoxA3No9H59UYVPFmwEJ+LAukbboCQ2R8jWa9qKyS7ctIaoDOJ
yINMXAYM3iuCZclxxvDWIR4E4AP08+7nUDhqHqKGzdu9BGCzCbgBEIQIijX1z5M9M9noPOZoC96z
Lzo+44UIKtVVZs89mVkKPmT7XtjTTVlhSgOswDcucWqEomOWzeGkH06TXH9gXPA8UAEX/qUj7WKA
Oc28TBLg0vYPYwbxoF2lzyB262B1S5S4sEv3XkRG/0ayStYM+TbyPHj3s8vaDtVJLprj57EvsPg9
YPqOgZ7tg/Q67ak55jUjm5ASIo98CwvHqr2iofzEaXDmh9VQKYic34iVrez8qpPtL6h3A7MxMaDQ
y+WKr4ta19uZTbygOkudMqwrEuGefvWiEEyTQNFrmZ09jssLOoBKt63Kbs3C8vxT/dwS2dR2XlNL
H9X+aOrFV3CvULcAURWdogiu3UatBSwqeFYDy7lrrUHzit5pejohjPyeLn3+2eWtddWwEGYrOEmC
irdPn10IxFTCpeQs/RqbnRmwOKql1L29fDKMcH9F4KrLfRlSy8kHKdzxe/nEsFHwRDHo5eAB8RRq
NUQwtA5kxqHyxTu5rvya0UbifC6hO0TeKfUjUIRy3cf0FtA9RweH+1N6X0eut2Pi8dJDZKVk/m+l
ze4MJawmu/p9GPQv+8h+Niz5FAP1NRbA5xY85y2dPLEKVhH8v7XZxMhy2jb8yvWZ0oykxmWVnQRM
5qGcQ2BiuRjR7SVO166SLZJCMHiUuz+Ria3Xqm63Vp16dLYKlMiiE2raDDldHvswNduLNckEHsci
rKDa7Pidvxt+Kaemvjo4XQ+NFaDCgeJf/9X2s7oLfc/2MO/MZ7t4wEZkEm5wIrJdsraq5RPIfNBe
0yyp2ArHaGTeTPrjKYf9hwHaKvldff5Xyp4QNr1qhF+Qk74uIMO90vmEq34ljKw8i5R32WyNR32b
iFXm43CCB+Ufar4laZH0Y906LGrubiu5ZcT0RxR7Pxrh+xqNHRkxhaZ412UiCH9sdVdhR2KHbZib
NyOnydBfOANLLlkEBER8tdU2+Z/BfVE/yDJUO7GxAEI0FO6wGi2oYypH8BINrg1Z7OhI1Cz4CH32
Goh/mCG4hmeMpRGZaIUpdO3HtqWC4U36TzX9iGD7JQCVG18FzeiIah8noK94pXUn7lTlUoFYQc7X
pFqPg4qvwM3+By5UleOiuzQIOrNg3droe6wTFOpW4VnAr8Ufil/kDZ5kCbpsB5YFN8JL5vbNLzm3
WRsK4QawkpYYQLyC2pgKTXoOmnRlsp3JE8qcqhEkrCXHIQ6LiLsbtwQihuiFqP9tHlXsvl4Lk2Oc
72tIJxcf8Qh3UxHEdipKfhwbGVWbhLhw3amt6zdsKrya9/JbwtpHO+km0FZlmkd5t9wf/DGvKEwg
ymtTVPko3KkhEzlkdD2SBXa6gY1GRfYdt4yYs5hfLdE9WnBQIDnCFLHKMEJJF/Ys2VfG9J0OPtLK
J1p/e+O7wYAJYNhYwdHVjCrvKIyuzODRPJ0Ovv33lvSdONTxTi2P7xPVd8/9TsDYy1wieXHF7gen
u9CFzC4hppPDPFV9IMe3wusj8+FlHeqH7H7Al3oMQOF1Mlj5ziNhl7v7jkfRxl+t7rVPrTEbeKvX
aoaW8RBVeK6BVtZyZpzMu4bPSpc1Ssnf39MHXW8NnND/n8q21KTjfvOIVxCaofJqyWCyUUkNAJif
YxUb8d7+Gl4+PrpFv72aNis4qkjBrULrvUskm17sg3KfFbsILTcfgGbVsJjx70SkEhYvUAM7UOje
17wlEmamuJp7M3rWhlI0+B3xTv7LuAeQK72vBxtJcOwUzg4dcRsi2u235Nob2trP/1O2Okf2Cwp3
UPIutHzpg1vVoZ7K3aihsge9EP0muFH6MmQuAbdi0Fu5Or3bKd8b1OKgAWtQyk5VKHTLlnSNq4hJ
0g3z2QDqc36fa1tuDuHxw0+HweZcE8poK1DmoKYjL9sTwOF8hMwyA8+8tKiFfH+55O3wi4IApd48
8Xq1Q9KDKgJyXj4bs9hpQXtfQQsVTU+nyL4lbdxQ1U4fQAgXByaVHZpymxeAjyfkUI8ijOkCcnHg
wodvIBebfXXsVttzF6BiOL9q1Tm2iIhL1ZQcQz3tRvRpchQJL0RY23Y0le+bWYcfofqO3p6sGyeg
3O2Cr/ZHyIKlr27GvPxt+Co8RGMwsqqgUgOyQw1bRg3VSuma4HyH6FiJZObd5+q27FB63uGmx0ev
R7JBd6OwKY9I6P5SPGBLNIgY/wblnDoOsEX4LGFFZEBTtDquth+s7BLRtKM9A/AxvgRQBj7eZmlY
hilCP0b2s7rtGBXpvCiWxu1dTwpk15ykTvu3oAvpCnOBCdtpJWO7zpi3+c/xKqeb/5vLb7yfLLNB
cpdwHrZa1XXvgFreYKMD5bPdBQWh3NfZnVMWxZw9nzg0W7Qj/P7EPkjuOgjKRnCBXVgDTFPjOh0l
qWXYQYzej8in+jKjifmkw6qnVykzIdctDgjk8hhpg12tCpviIO2MiXEvC6icbiGplinGHPFAjA7g
S7OLulJiNV9OPurI9mADIi4wF9ei2xllt/4WVhDKIQK4UJGxYXwZVEfykQ3wJpPL4WIBinEJOLv7
SezwLdOZu3XAVy89tNiW6+1SxdoDiR/kppSl3fnfQXXDGfjHZ+285FqP4maLkcTZGHGRofYKVojp
HxbfE8deey7HBGZpNLRDl9al74h++dQ2csBZ2LB3JVwbhbXEnICZueooHF1THciN4HEyefkBGBx7
d07ful/S6XjRF04BaSiYC7BWG8F5ZPWGdAXLpRVIbNLx+la2CD5UVHrX7u6ZR78HuJZVP16WLkvL
Goplqrn6I85xC87hToEE/SrvSacK0f8mkFchoBVArvYkI/2XyVhXp79540ihi6hGY5SNWtUv6sfC
Dy4C1vDS2e302wsfbVenhcJsJ9cicRs1NGRZ0O+m22a6Jws1B6lb663wBt1nIa0SFFeMXWeLtF84
VmCfa3cGZQvgnQShedI4O8KDte1lYRQWRQ7mwPoKMS9SeYuOg3Ga7jWX68eGHvju1QgXZR5Fd9qt
0Z8PhHCwmOPX6URHwOyyEHtk0WSl3+XkU+RwWlOhJEjaLVyWKrgHT4ypAyeILoZZ6Tk4ut6gFLTz
t2Qwmpe+977nNLv1kCqTcdE425Tuj1iCtrzj7eH85euTx1k1dymOVdrkkTlOU4zj1IA83jPoYMd4
GvI2MswW9HjOaMtXZ6TN4XUBd924h3MNARTIPASehHNhRla+zkRiLYs5kH7r2P+6Ad7sr0Ts0qiL
3l2GalW6Wf9wUPP9fatqApJzBWCiQhoDSpV4zbH8gl+PgrruFdXiUxuQ2sIhpH6lMHSftgPxvZWi
NOeUbCo8wXWU77RIPrvRHU934B2n0IhSaGAICu0a4hwlowuy48x8KT7qHRaI+PbQrAJS4Z/R1o+Q
uKorfBNwFLTtnkQBVDV33+l6sznolPDrmO6pIT1pw85TCUlgGO8otzW33E3WBt890sbpDIRrIC+z
dzw7po0DOxEiSgCkvEoWdTzhp4GSEJkBQWOUxs/e/fPpwX1bDaDQyUhiH9jrH14/4kkZ6UXdiisW
iLpBgeVG7D3OqhnWiCtJKHS9qtbqeoK5ALNYyWVlvV9UlNp/FZOCt4P9bsDrm6Mel+gcfgGkoUVR
l+0JWlkBPnwJ7izB6usEEbb6uzDIS+fDam83V4Kw5+XPOAHGeDVEVHFWuRMkrODjbs45sEnRL5zW
NtSWRqdd90aLN85anhQok6KTqkmJhT9u5xgrttcHXHqr+6jUViztjr5f6K6LqfUBWtGQx4UwXGKO
yWvE2NshO+10hC0DgW/3I8wgNnpH4iLmpzBLKRwpkvxcfBscEd0nti652wQkGNDyIggHYzvV6rcO
HyGTpOatDWxro7bYSYwsRSrppc0LSM3Il6dg/H+DS/+/7ftMjhKUGoCUydI+hiPJPoBwpjOxIdU7
wlElgdKSHRo+nwV1WLGBTFCW/5szGzyC3nqPTk1BU0Nfn+DQ4cjk+T2opUBpizS8F1c2jPSEgm57
MUi56E5t1x8EP6B8rFb7AaAheK3DP8Dka5Qa76mmHRfWTk09r0QbqTY87xgpLgFLrpOuM43AaXU7
zASdQ1zLJUX5a+gfNwO4cB8dESileHe7m4M2eFjzbpPNAAoZSCqUixTTdYy+o2e8yLKLZpqdFWEf
RWGlvXNZdaK3zHzoT8j6QAKlKrnwPIjPNDkGyIcgTSsjxpCzHebKbLnZPmNVtqExLXAVoNDRRxtt
QflJ5ikZT+8Yy7cn4xgRgkrLhG7Ui/GJ1SRLRxV7NnI8sPi8rimLH3JOQ7Lp6MjC4veunmaZDEFa
WpfbI/WuVNOj2xnr6/yM21HJEK6wDzUGynlzyVJaCFupo9KiT5ckx4OZS+qOElbd+YL9eS4Dyokn
DAvHbOzlgt4SVIUx/TvWOuXz06arfLW2YEruvhz+P/GP0dAy8BHzLAHqEkOTBD+6iTvpQ1SzIqEl
WsNd0N4KqFSh33ANFove5zT9qWWpYeAKYY4Nir+lsOXIpx7lGW9Ff+j6OZviiUTv3IXKDlPZ2SYS
OJACIpfoy71AEd5ZkTrbYYsNi3rkFR1D5TDRJy/iXH7YX+xoN+jdTUGx0OoMM6wlGWFf+j/B1iiE
VxgLJCPloxqSFqVNE3WNfOujodYlWt7BimEv1MvIvhd3VGU6MwKn5PzrcDV5GDJQAf2fsq/w+xsm
J/7kLeDcRBpBzBKiz1nu9aRQTfErSqMd17Y31raSG+k8sE+ZBp23uy8QXMr+1ZN74ejvz53gRSKJ
WfNfiauKhc09r3l4MWs+m2eJjpwAqiPIJMHaHKwBWwMjLu/lb5Me47FqFVYKMtpgfwz+TO7JBx6C
XRRvlTn6etsCE8gxC4562CUTch1om4ZmbXxg1AZLZOitfSaQ2Lq2MMk4Og5OPel6fVmVYVXhVJTH
uf2qF58NnWNweieZQqiTRyh0RwbxlLw25HZluv93CluieviGzExkpjjcl/aD3aP9M+fKKp7pLbBg
IGGV5NzrQXMVtxoo/+Eh3MzQFGH80Jif5MskFYVrnlwFaimqvUEccsrXv0pEwaxInxUkq4aslSCD
W2M77pZV/Bn4i7gQdu+910u7wgivxTeY0RCbpx6/nVnzwFWEc7YpZcEguD75kIEWNP1lq/tDXceV
4PJQZdEFO+iS196NIcMrApWRy0fanedvMzEXRwZNHqs8XYZAeBY3hRL60kLt6ixJzRS0CGxP+1gE
QyXwdK+uqUMtlVrqB/yQ8/yecOecVQpQKfvgnsur0TsZmCJstzYfwdoTe89elw8xGTrf4WPQMS4L
8GrPIgU6Zqr/1IbRMQq6gH6LU9MAttOWj9ATWbO+eTKWLixC6x4A9lrJzz4q1EjaOqkRnZ8b5MqY
+fxIkXqyH9ka8kjJMLE0M9lGguwASNAonZN4J19+5QSpho3w65Bf4IvOnqidUBpR8eMkfHBv46Qk
jJS+t35GZ7Okx7bitrM9Bq0reCGtBcCeA4+WK4WalzmFPgvhFm3UfR7c78XFxDvJNfot2eeuZRRb
wHbS1dnQIJSWiwSXhznmtk5/+lz9d2fp9Vjn4mhx9fcXAzmfjqh5jIUSzcveY7d+aXJOIDMaEMqK
z8m6sy6cxIHatkI0Jl/6axd2/LhkPIBMqjWyeTwMKaG4XoahyjmAgrdATt5v9P0Gb1opkFpN1VVp
pjgYNM9Wx7z4xhZ4lWVwi10KQvqGtnyeWVvQOmFmvyfnp6AHk5PkIn4vAtbY9Zv4xRNZ7KlTSdfk
LX8KqrGk07/XuNiDPmNbxJWwSKA4cOz8SYfgJTeUXnfSHovHutX4mlkspsrtuk5VHpvWe1dFE/Jm
84UWfyoBxKT3SOXCP9taA2g+BJ/tbyYpL6X99eDW0OZP4jOl72Pj0/QcRN5/rgygeMnPEmm187/2
TDV+/McgOUJxEsRhkKkMAEFsuvOHBPFkUpi6A0OxwO7SLwlhql9qEA0p2f0qReot+2RYv1mDFQl7
FMGmJGSBWNUiBkQVSLgJrnRhX1iX9FmdQjGIYOilGi/4cgYib4SjVA1LpJpIvCz/ut2fSDLtm+kW
eVe+otvFC5jbJfWVJRq87tdqY5sE/yTbfPZQxbD08pqvDG7D0qS//q0UrclWD/Lpk8HMt/aMjNQa
01DZ0aYbY82jJ4hlCOwmPn+xc1YHte2kUHVZJ3SWiZPQBObz8tFYYr2A/LkXpggxYwAsgsxOqTxL
7H4YMxlxUYlDnVgcOFss10nLIyqNgHY4mX7wI2MBBslp1jTo/De7ecY0Qa5VbI4HsdGfopMM1bt3
1V6qovArIGe9eoATaBcqttmdAvrJAfyxQHXdlMjKGWipCdzb2Jb460j1ezAdxh6LKrfr9orz2DhB
2QKVb8T9eLBs1gC22orCxiugJUACZQO+bH+urTPWEJhO6vb6e/W+8C7Du6LMv7QWUxhx+zIF1K6R
lu8sl5FDwf0Tr+WuaPO5utOT95NkVO28SxvaWk8KDslNH7HYDDxlVW8PNE5rzg4fKaQ5ej7U5qh+
zzlEESZpXHpkzLw9+7YHtZ//mHz936O70WpgziqN440K7hHLe0Gz8DxS4bzrTTkmhhiNFL7fA2Vi
n9hx+f43Il8oasVNhgkhJt3hpeI+2ALSVIJHTbzn9lUzCppBdUF8onw+fVYCVs7IasVQKhh2y526
24ST0sJHVhdQCX1/bcA4G6Yz1RaZ62+i0Gn5Wva8TBHZiQs5NUs2kDWmm0jGayq4XTkeit5cSSYE
ulFJgNApzp75RhwvxQhzyJbdi00wicZt5slNyGBjMMJkSOScrbyaEuIb7fIXLxlUQGlnPpRC/d/Z
FX/z+o/frFGWQjYgE9XieroIm5YqauAsIwFrfmLMvKhTpl+4EBI/D+3fMXwo8AlVnTg3PA+DBSSf
M1MTGFfA8WAE2RSBWTFwsfmwI4vVn2B4K9nEcm3bgWIAKHP5oUijrJp2kn7XJziA2xGbfirWeys5
cHUGvOoEW2s5rKXiAw0dyg7y56yhSffZr6s6Ozp3iYjtyCjz5AUAtzUj1AGQjO9eeV2DraFGN+XS
pbXnMeMUqqYbzvEXSI4qwJPoJP/Q/WSzjj8/iZcdMhY1WiVdEgceLxkuoJZi7vjduBZkvrm/ufCQ
hK7n1ivgUdWBbG9hfbpTajawIRRR0N0KJln+pW11/8UABMIQ6hiZjKLiPbZIfU6Fid7FznzJgz5s
031jnGtUj4O+nKNrOjFRMZaIDM8UV2kiMV4G36GYGqmjyFQkfWYnNdgE7P6FEFRWQmmL+WvgGG4t
V/aOW6vE+vMg1xfuvXLRXX/5jecIS2Y4SjUw9DSOtlWaJf/CwoH+5U84bTb4JD+h8SuyxCogzK9J
vyghZpYhF0Im/olxdRdfO7wpv131eYG8zOASLhh2I9YKLKttOU9W0aEhCJAv20ZdBuzP/D42QID8
+mSUmYELX1WvFG5McpXdffju1tvjJ8CoQ3klLt+tq2lqRYrFoIWph1pqu31T5YY1G7aL13FTMo38
23vh5DaEiLFlxbMerPR1xg+5VvaT7AgDxqXEiuN/+QM9KAj7Cy4exJlcnEjK7RsmNiFqnrq3EYgA
NRBLSCI5sKfb1GqI4G+8aiWcayUiAFMCLhjbCtsIeSRhL5m6FGKMaQFAeodd+Q36/EPgFkaO/Wsx
YDAXew6ml5J5smi2mqaTSpB7AOolkdP6j8pl8MIA56g0DTuzWuIzU0Ke9jBLhfrIiG2E66oKR8F4
U59O2ZnLfR7VBEJBgjtstaZKtVxm8qE7T26YkDeEQnWwywh8Vp4ahR9L4/xy2IsK403JKwL5e9rK
AvTzjRICb67/tj5fOjbkZLyVhYjWPR+MUsATLofrdH/qqlX9iJh8LBlALSqBYDtk0WqPUZbpw9Xq
nPpPYIfNqyD1BEF40U1fnqJPnv+oqNziK+eAVrsi6Mc7MMmP7QrBhlAGnEWiH1u/s8yh+TNNrRbN
Dpdc4zHe/JgimmzyiK/JMQI1xbQ+FeehB11api248GtE00wzNtr1iOYlsnZG2KG9IUpgreX85o78
STARQ7hl6dCqWqHiA6hwMuQvMG8WvZo4unUa6VSLKcWwIPdab8NtDCt0Fl0GehErbJn2lEuQtSnU
hdwGEBmPeGgXQhL3hglwOc0/HNecbaZNvmfczfhPSCSoWfnvv3aRYQwkdG84F0CpP3+qWwAa8QWK
U/Ik+59uS1UMhsE1OEMP+r2fFLXlUZQDFgplarHXzgKc4NCc+QapcBDa6HDSPpANqa0WSuRMBnYm
2fDmO/mLltkoJrJiGWeu7z067TU08wogtq+m9ov671FwlWGksVhwlD8EMgwjLQd9TOnwHfCwYuuR
Q9ef4dEmrK1qsz44cXplx1Q0bMzlYz7bqMT+U8SZjQBnk1qVQwWviTlUdSBxiKsONxt41Qc51fur
Bh8lRY1N7U3GUVJhg0ZOPzizqWzhAfOr9dfsg5NRx4llFjE4qAsvAuRUrsuGyQmY1UKVXpQh96Kq
LvLKWetzOYeOzkfz56k8xKfEdyIx0mMKQq55ZGwFLlPJAqDpEWGUITay2nX0IXcRcT50wC92/2k1
AhZnpAuYAgZkZnrmTdx99EoPrjOnCjzN8LVjQH/yiQv5I1cW4Z2Y4Hm+dXTGO8y1UxkRSej3dBkH
n12X2NJXtvQVyItYf/xOGgTZF+WlY3wAcXe8Qt46uQ/8+QaORTdNNoYmiF0OOYqg/lqsG8GtzbG3
gotpjcULjUTREcwFojYfqX/SaKUjNDU4vMsOs5tLHCMYebr+V3Ak5Bs3CNmKlfX0sJbZswUPTfRS
AsInabJGTuMH/9kqSObqk+jlxpRUEyRa/i6b6dlKtMeVLaL0GSNtv0DCPiAZPzHZLbqMQlDhp7gd
dRfLHOK6fEX8WNn9P6GCmr+bHalXX4OBC8Yxq9SrmXAhkOUc8cSwmhXZJ6TAgVo/yKScq1U1opyL
Ccs25Au1LK/Q0xv+iBjr2iyd3UOPuZLtH0ri8rnQDeOqe4uH9t3LXIPQYYuBO38jE9/UVG9BVwTn
1B/vS2oqgd8Uu2DCuGeEOEtAJ0+rnzFiBtANoBciKSsF8B0g/iqv/MPf9PGBPJ7AquPIUBklE5Mz
vM60UvaPMcE2U4jlxQgxmaQVG+L5vwpI+SHQI3/PB8QsDbZpkUmWca8R4SvHnDDCqzuxWJWRHtNA
Qg7fE6tMbuvLaiBa3+JJnWdfr0UsRTK7QfInDPGAQh56Sb4ET9ZEE1diZkiDeK7qxYkLV1V3OMPd
XMHRLeY9Gd2Eak3TEcks3sF3wankdnMoOBJSyIYZfTByQV3gNTw69EsR6ICHoK2gQrkHV9qs2k0D
O0FRTxi3eU29a4ZAKgPu9oJtmn6bZpqAy3D5bGq8RxO3ZEwG/4hpmsOeZmQvKSI68dPmju61PY0v
yMOwBTYP/PajHU5ngfpgIYq2uKFcnWqvI/KH0yfmTOEJF9ZJIDQqM36+ENj8AbLw+kKhV5nOS7G8
UgV8u9Adw6UpWwc5Snl6FxyR606zpfZGdOUxZUX3I3P4L9nL7NMG2AnGo7WcwdbH/QYFV0HJ8oqh
mpqezpNGUN+9ANVNC7hzuMZK79xm/MJahsLcnsA7aFk3AeuJFP2wzAyJuNd0p8wOLtPcxO5L6f/l
mLh0I7ycwSzMeWYDlvCkYJRL2PLPB7xn9Dwbt9LN3leVKEmhk6V+pxf1bqMvFmkGwkuaDN/gtKQd
vTKoWt1d4lat0GX11tSlZRK1KmaLdzPOrF51E60QXXPPHSYVy280+z7+zwXdn9G9VULQhsu1V00/
TXcT8y3BJ39jDHyUJbZEIyHhL4FdcrxZ+E/aLjvaaRH7B+DEqBHachTI2D7Z+7Tf17THZtDT3afR
TK3WoAFzyNsdR87WMZQykrO5n27FlPJLrFO6WjoW3k6QPe18lAfeEfh+bUHZ5YFpTJ/QBBllXtwF
+L1cirU0U7TgoUtqMbfxi6RD2CslxGX6Hm+GWLkBOzlwVt14S/ln3nESPfqu2uksC3fMg5G06Agu
xbadBRvnsYxVgcTWeSZ603EQ8jv5xIx/HHiUc7ewZbI4umBjaimgy550wFXz3z2VJ07KDyU6l7Mj
X8q7u35DdX3zLz3XxZRg1d01hijZMzXk740Fum5eZZR8pi4ngK5NaPpQ3/T0TgboCTSgdXmD48nO
FhItMlzrov9pcCwXyQtq9lpapp0/C58yo3EkBXM3RmNooiN9F1xlplOxNHFA9ZNlmLY8AvKw3E4C
tAmcbVzwKXyKFEhlhmr1hJk7e+3YWhsnQWQ1KcO3ZfdzYo+BGepgPMOcajgJH5aKDNM3siXkj2ds
aAlHtX4xeeCBiKHlSagGo/wF8Z5RexcbPZHyE9+ZhPZoDRl+7Hw1ZOqaUP2bmuYTxEmKn/23STuw
IU+w+NSGSlbZSdbKbqJ1ihTJWF1KprmKVj3SjQE1GL4kgh9TcqvsdNnmpN0sOV2pTNsPKbJ4zpUI
tsh8wWulGHqzj681i+4bcIey7QnzbLWMtgl2xl6ScA6V7TotlfCwC69lgYj1AMSIKzHpXSFv9fNO
X76HZP+54Loiwm2rdYyOC7jw5Tr3htekMjV1kaiddjn44gofGD4+5Iq9mRC6fsXv4W9ctvBp36Ng
btcfzRIcCUr/Gg+QGkKp7udh8R6z3XHrac97tSXEPkzmQCLFHr+gRgy9OhxtrkTkEDCRU+1Z+YOF
KfhGqtVTzso+DkqwlsFwgoe+/THxhSiCbHRZcWPy8CCOtW389hfGKWY+a88TWM3fHI2hV31ShtH+
a6VyprchpjgSX6sY/P0I5U57rAyBiJMIHGC6iurdKuWLC4f8O8Xlefe7mqqSkPiSvFkr1XAQuJaS
CEhwCOSWR7NqYHB81lCrv4Lb3ep1sB61OiTFkIfxCJtYwwjBUjDCP6FkaT93dy2RXor9GIbYHHA0
ikTjF2EDVwHSXOdI/i1KV+AZKGyaWmnYN+Kj/TNY+HG0JUguIRtdfLEoxKjeePrkjugV5q6n03Ws
wbpGvqXnRgJQeVgRbkbqaof7HJIYphICWZT3qRs/XNzDc0CeBMdQsaec+dFLSLGc/sV0KHChmVaZ
dq7phcrpw/hCZl4+ruum3HKpWPUT0BQeTRJq16b/DJHaK8icLy1aICfCMwluMli4TxtzoZEiphRv
MNiXQjLZRvR5IEaYq7yvVh02ltqnZfIjnFn6K7A1CJFXzU39DCx1FLYVg0+hnPWnSZp8QxclMArM
P4DC+xobdA5hANbVTj6xxzlT9N6RdS9bmLtWPK1MYAlbLlbUjOVMkK1s7aL/PmmSZ980peGmHk26
3McAcWWURj0VBPNHFlrVYc0C+VPuYxzfDFXIHOUrG+ij4jlaDlHih/yzq8ODEnBpJOeXIyaBeASv
v0b+BsqqM34v7gPsNARUv7OMl2ORANHi4KqCD3YqYM/ClbjPEy39mbsZYnz6ynJ5EY3hvVtMEU48
hq9B79zlAfJ/PSI+ve2Ewr97fM+YiD4p/SPjmVgFunPNjybklP6mLbgTXGw7e/5VJG3vFhn/bTCA
NkaAZ5Tnj60X4upJsCn9CaAJGi+MxETE1Jd00Vd5Q1x2waY6McMLNmOazuodeVXImuDRW+gnlHOS
xMxUPNSDDTl2HtYtK1lID+Z6LiR7t6r3WUlwJWHr2zmNEVDEwV8pxj06JH8a2K4uxWmHYqUDCsOR
2F7SSnjjAHm3oqpSo39wkHZ/b85OkNyXkHtBDT/lZ3SDOugboP7cAJUz+lNioRd3slap5WWNeqFN
9+ilhFPG8EClN8+R3Np1VEsZooOB3a2Y/P4W+zqmWGcqD1lqJN7UVG0Yc8Niz84Ra/FRiD8RGcaz
uPjaZt0aA4/mEAYPJZ2K5WXP8h7mTpFwGexC229/yGzl+7I6DExPv+xnbkyZVwixkDim0HjhQI5T
2f5nVcwGvXD9o2Is3CWLc8isGmIUMqRKTAfOdyl7MimosPp2f+sfBrElYYKwu5IIVFTQRo76TIN3
MPyaK7uzxjeKuTHg0rmT9KZcpf3yZQsUDJLnbBtUSIKwpTs0/wYQxpIcSXRY0HazpCTbUYLlzdrD
T4qhtzFD/U5ELQeLsRM6Wg7g8HGCHzqqOtyd/C9TPLIVn3rvPaodKLPNPQnwWH+Y36Tu+d1S1VRY
Hz+AUmJjcd79AByG/y74Q34IERObl9umhdRmx8qe2ElofZdVp+oI5WAheVjP0JtV2fxxcSFmJ1Md
MNACTfCfHHj4AldQfSjqV9yeTt9bhSa8CBK8ejh7sPdCC/X0DoLmi7bDNO2WPoCvOmlrUdKFw9vI
gtjm0Ln7GL1RioYmqCAKeD8mlJ4OE0BXBMg179Uk+jZKZc1v9/qcpULQhLV3UDeEePSuD5zmHawF
p85qLfXUwmi63Z5V6KvH5RqVWBtOiMTJE6AAsT3f8Ec2CaamfPcVr1+O1Bq4mcBJJi10j8AzcT83
23Pl6Qdw3YZfBxuRTzh8eJJZNmdlFBfDkY641yHXB/+gmTgRCPHtEQ+GKMg5IZIvuBuaoHZDVT73
lHEqLipkk8DizBmhQ445TRDGB7Bpx/S2DzwVKciBleytPRInf1BYwmD27ds1F0QXE9UXpDZ13cBW
2YA2NUnNrsvwGFadhFsxtjKTe97eXIyMvbTF5NPuRMguRv4HbQRNgKS7MKVqYDoS/B93lirOQbIZ
5y3PgJtbobWBcl9dM4YV/l4Xp46Gzp9RzqXj6TKra3EqKqeajvmNWsXeGiqKGBjeJBv3Q2ofcYVF
/jdiVH5fZrlCey/A82gSnv/1MrKmhXwXtgbQihALhZRrcREU26vQpDAz9DRoOntLvN2PNVZqm25q
7us+ZNAUAiRN3tkEhBsohcHjO6RAKT70CV1qTJluSTYKjUJeOqxd84ERUw7xvHzfnyFAHSx3oFMj
um+NYirQBUvyJHBXWwOjPNH693CjHevhJ//2Yz7hTAKStO2rLUSO9emdSjlnuduIKiOo4eezu9mQ
/DaALrm/uy7v7g6yIaUqqyqFgah9RzggGx2CaRF2Ct2V6b188MejpZFjSBzIARzZn4hh+LR4k5o0
k3KIdoiUtB+MgBSYqYgYNdjmh/EnSGVKotABTU1s2NhfeKhzG/aUm2zRSLXBds306MEDX0KTAaaK
fYhGGRvC4Y9tXfzrPZVcT5jo09KZ2wfP+VZ0D5YtYHfKGyZyKsak7zGhc/MsdsrEP4FhoxgB669I
hxX+JctCM5eMxy7Fgela/BHoIz5mkGoNxl/P0hjazXsEbxuSQUbTA4ISUNWG+UTT6FKo01++u6z+
DFJJRMalPwV+VVA+8oSpYETKVwS+Z6DNSV14UN6xEQzxzOgt3OeI0OISyHw5FPOXoC+VMcD3V4f7
3aW2IfrbFKq45XCf6swBFnGDAuDT0rAyHzRcjAvKhzri9UVfN0xRVH+OF4D4aWlnJ98C6V86wci0
l6be2Uy1ZwDFl6/8w9pmJz9T9hbVlcOjh73CJk6bGAf1TacnTR8Gcqs8RS/J7QiBcXDZOsIWZ9se
J02iwbtLzvWAxUAu2+2ksbF3h6ffGcxrk64e7ErqbOGWuTVuzFsKg6IW3shbTBHdNcFCr7oHZtuR
Zp2XDWcl5KzShzuBsFX70U1NWBlJUDfgA1VX20F7BRTkEhBok6rUBeUN3fA2foJ/3ikmccVQwkPl
5DQSyfKCVjtOZkUWctA+HF1y0g69sfK1tiFHko1pS73ATqQM0l2I4430/+KukolkgaOtjg9BoEJv
S4y/B8J/BAXiBugw1DfE4/2ZXHoAE0j/gHUzV1WxEjEPf0WEk1lhUemRx7rvltRzWBK7vY1x7w36
qrf3gSvQvtRUbqJmfFLBnXGHE7DdyKUBhF4QgutvsfOh73eKBD1p8vHDgG7qYqHLCxmg+9fFaLZI
jHbKW6JxbS0J4ER5HMdwzAuGZzFWUfh7UALWGCvnW6RLrX+3EyIdMqN2th80v8j4aoHa0b46GWO1
wrpqUmRxI0zD2Sc7rdxSAxaku/6fCt3RnVy4ZclY3KvX/CDCQIpnQhlxWPGx5uh/MzzdwQINmLBm
xXX3o+BGrRsly8EtlcShEvVkAZFVNJ+kWoq7Y7PDtXHwj2+VCRj1b8x107ghRSRD44i7RsKoIdph
kVAqrr2Tu89nNhYQAaO71AH7EqUsiDS4B+dR+i14oisqFO/w4uj/e5qj0ESHbeSyV5JmIfnpNnKt
QyJrv/GCtw2o4vCzgfRF3GTKUjReigSy+SPo4XV0r6AkZRpOyxrU2YNSjS6jVfPh8hLaxuOArPnM
4TMF89BtNXO2N+Ni3MggCFfZ+F69h5REygHxyZ3nbVWa9gytDjb5HseXt31AmUsgcWXmd57EWx0E
nipGQR2kcMbyuQ2XhlMTeGUsUz+TwGPXHbC4ITgW/0Fnn+N+2HHUiVo+v917OkC7rQnxofPS4qXx
6NdfEV/QOM/qggg1Jeu53euNKzUqR/Z1uiW/jn681eu2PPbBIycLEKn5fQ/TPCmjUUlkpoj2r4si
EMFLhiIKKzxPhwMVG7MoKelyRSsFu5Ou8edwndpzNzL9v4sAQ3AvbCFvwml/rN/3mq1sMPYAzhM6
73+kihqM6aFBAEjYwvGmE9fmafaZpv8UjCo9pBxmQgbjhIgL0G1wyUMGRUb4hG3Yhllz1N7gK1jI
owSGoui+1JwltKDmvBC/ffyuRaZoG74Z9SmGrj08WjLO1haRUKwPV/0MIyhB7d8VtqjhSM60VTHc
GcRFPlaoWoAfmXgtzbp6KEq23NDyvwjNrs3RrEYDHMVpKcwwSEItzGBdg7w/Q9eySPEayN6MRTYk
EhcAOn1LErraitTxNnJwgjHyzcsi8bpgJI3A6EBPjlAp+VS1E/vybfEsMwg+PbBFEGc6GGoAt8Qc
51zfHrZoRc0q2EAgY46B6sIKkXFVo8PozipetyDHNEYS8jTxetE9yf1oN4gX3f44Ccnrz71M2QPe
i2CB9PY67bOT1Ta/zxxsYiV+dCZ5NCDWNQ9pVcvQNYdIvPnEPVDOAK0X4Bz11xzLwczbkGrh9Ot1
JDT8PZe7aMZDA6qDyzZUkNU687MDMBcK4HDK5v2fjV0rJgmrn8iwqrCVrGNO/1AjyE/CkOirOZcY
I8rFFa6g96watntpO/A49q5m2St2CJbK90WuY0yVVydWyVB69JzFamFQPx1dDlwuvi8bVbaHpnv1
Z2NuLUvaNpsR45XV8xWhWKvR2GV6kPpp6Q/WKeCvGHQkpXEc9NoFW4RRFV1Jd56pomluDeil5L2+
1sxKeYYlaltUL2oLsfX36eBjdlXPOtqljvAsyza4D+65tUWVrawafmd5Y66TRaeH2KBWrNbpIh7o
qItWiMq0ez7hzMzRkNSnFqaiUEd/BbZYEAwYfab5JHAqBefhYYU3skiPMTEUKa+DOyJuooXq4zbr
1eSTTysTYLeI6vwV3YQd9BSuZZSpN7bzezm1QdhzMT5JkX2KsBn3QH0dpu4ORnQJOa24Zt4uFzl7
kHu6HQIKB+3CM/9wyniwmbfSVzbei7366E3hB0hFOtGP2/HlhOV5EFlpiRYUPPkRS3L8JR1YFQmA
Im56gJ3VCoonuNt6i9dqPQJ4qCjr/Qxt3SIUg1wGO4PTAzf36ewOJ05T/bAScP6h3X+ta6LkdUgv
BiCDYk3SRtDPdMZTZuch1W/GkVG5704LxThxtW5WBLYJF1iJ8ik456v12EVcHCX+Adbn/jL58dkd
bhX/BjDuUT4IeFbVz/VPxAporwHygYbVUbFtf1uoBRgXHhfmBJmmxh41aBxlV17QXqF17E1I8F+P
50MzeeKhORkRmQenjTft+ODXTC0Ujn/ICMP96tnwfoMR7t8YHx7kO4xBvECzLkKSrp53W6OyFNGo
3GOHSwFJqv/qCbIrZ/5fTHXrSGNpxMzT2m/t0JubyMyZfNAeavme617AG7ZnVaxM7TR3h496Y1p1
laA7hx4hEHcrJ7f3D66sZVgs7c6YAOQC3yOQQVKeNjzxs0+3KKL1RbfGXspmUl5zgmQWzd09GupR
EH6H36hEMsnn4WlTMAym6kqRK149qlES+oZGYub3xQQh2ESl9w2BTUezrg6wyXtid0CXI/IL+e4Z
hqBlkdCKmld3ff1wXxmn9LDlUnEjVX7I93RE1+MGOPFGw9x4doy6Q+pSD6LkRmsHsSN+BZ4qIYdm
obALNNxKmKInGDw6Ejupom3oD14xAyCAgqhPSsNEx4HrLxuf+ZifqnqgIYMrToR5a8woqKOqacN1
Fk+nQhnCjsvZnn4U2T4dH4XJiNG5Dw92+Jn2IQujv1X+O2qPP5/cNsagqKX1T28UEQMSQ4ZtBdNF
H3VBtCcfezxFDtFxEPezxeUTq1B8zqFkd4Ls9Jcq7PQ1nPPAA72nNFo/D4mBnAMoqXs+yqXAYtnS
kqcPCPhwtF4brdJvg8AMn6aXdaw/DgT/7e7+YC9GwyDDoK6yiR3n8kZZib7jvdXzafv/e82llzf/
dPaRpaZSwNwgG9H4b7HlrkrRykQpKGdBoRxysWVjbQRJ8/sDZLdzwKYv+6aQfM1eI4iwS4TgDoqz
LKIoIFg4yU7EMgihEU+Gx2te6Q8i6uGHvoxckxL2MemJ0rKv6ioy2841Efu0g5k5yfiIaUEg0/d8
XoIbxDX53nKAnkm5kqgsXBxGaDsuhx0Bta3UDmvFN27EojbWfcQSLLOk2howE5X7XBfnG5T1Xea9
FKcLR8QJQgwiFemzCDhYn/5ElKIxklnICF4HjF3M40o+dozy8qbHV3eAIjM38Us/E13eKJrgznYL
xYl0zkrUdHeZBWKwE3u7sgkSzRajYDyGcRK51heNQMqy1sd8YpK6v7VaaU7nYomc+WCh/OCYn2Xl
A619F1cTw35R0zhK/YRIM/OqKk0HzG80uWWviE2yHkPZzIIV+W+ve256h0/9GxSq+nFmRmPs97bM
1sCfDKvh8fmsgmnxV26ZuC0TZMleVU3laqd+mEIZ/++qODmHz6ohQ/qHbU6f72CEP0ranwCdv3/2
nUAYsFrga52mlC4/k17cDDpubYsCE2XZWHZueK8IDGUzYvlTwVdx9GyY2+XAHbEyPzMfjtaC0lGZ
OB6kiAXnNWHepwSI32+cm+ORImqbVVVfloUtKsggIh3lnOtpAeZ5vtHQbOz0IRT46EZHLjC8l5n/
MhwYcd7/DOc8Y+lLf2X4S3yFVsnYUSzsFuM9K6E505uDxihHK304JiLuF9qDlngFgmxpqflwUO7v
oqRq7EaMfudda3zdGNDaP720M9mFzntglky3B4eJiqAz2TO9x/QgLB1hRy61YmUfDxTGWw3JzJ5i
5dDkN9Q9S94YnRlkyGHBv8ZOwJJosu50LeODIg8bTmDrIuH5yQUwrtyQ37nngOmYikUl1vGnJATx
AbyR8hDSbn+Il3N3Nx8ZcSeiMswCKPY2rXJMrThpihyxMFx0eCm/LifP32canASu0P2I5aWywqlk
/rG6QaoKAdo0tTb/RhP6/Oesr6d6ATsvxeDs+++R961Vzuf2eEO97/oiZMOl6bEs9GcVDhSONOBE
ci8MrLDd7Mq87UjeCUWuTw9nX9sbhdnbYyIXgTSaRDl2X8U2BqwbsmlaYkTnGxK33FUHWn5IimDc
9hVOVVF8LBaL3yMXwHdtXbmALy7leddd9LJAWqn8CTEjtyj/yzmRqSwbl+IBtX6aUhLG7TnhWjRp
JISWRZZkO7dqFOHCuwsWLLqh/xue0bLz0xJ4ORrNyZCl1J0254h6cZkDB5o/gAhvGf1gNAu81+wb
Heztu5nLw9tY+LV9KNk8AapCw/1+2BHFeYPHckRcyQrVRKpO8DmpJRg2HMTKA3brDIrru6LBBJjS
oIvNt8OyLtx25V5cbbYZnzrRa0HCLX+4i0x95r62+76fxSAdv+Pn5+M8IKkYjU7wUNQ6LV7gF9cg
zM5LktAbdtFk1L8yl+Ws8auBxOTYWJqk2iasaeokcYJufaw+rV7c8U3EeAw/hDoNx3ch31eOcblI
htzLZgPaGNJz6Kjp8fcoUlbjzyZnUejb/PRW1oY01B0Tz3Aqlfo3+ZZi+XVl4LstcpiFeocKPxa/
xl9WH0E984e6tF90e/Vodq8fWY+6AVdijykz7/Uwt4wY26KWfURKjgaZMJnpjIja0x6rP7YzIy5F
ZGTclniUdyA20YONXeekGP/z10t6KHZDu1XRLo3ebOYr1tkC5z/kedwbnYEW8yVwCNZ1nOD2aoJf
C412gaBJd1P5RTPSLwbls4rwFysMhQ/QUH4LDfquvXOfJ3BoiBdktxWcs2QlPmvD9PQRx9Z63iSi
nmUnNjdOboec2PfOtAxVL3bOxSZ3sMKKsDR0YJwPQgvu03sLUEJbBTByt55VH2EFX4k+6IqR4heE
/1zkrsyi275K+3TB8xVZoRjnXYHFSxt3ai5JGb3MFDiPGgODP63gzva4BjP++b1yO2yt1kGxbRE2
E2mYNplJeknEIZEkpZiz6M6aT7hfBaATq+XYzjbnk+9sACpvAPIAWELCL2ChCJf3Kn4MHFf8V3lt
bGD3MEq2w2mOxax1byKR9uefYJ5dDfTeB+rl8KOC3cXAmHuoKqx7Dbt4WNhLp51rj+Ac2I8vQFZx
cLYj5C/Zuj7Sfiwle1P/nFD4g41RvL0Hr+l2AJt1L+LKDeWOPQGjTkTIWTLO8ZL2u6hJ7jgFqW8X
Zbftfrl+t+Z6UHedYNTpJIFTuVmkdRJTX4sL+UI3SIUP0W7qoPcElavznf1GA74h5enmfEYMMXBM
e82zAv4my4pjRSnjZnlJz48M9Ih22mp3gDMtvLAaYXXHXkZsOYXOeD941CwtHZAO+MEcK0ANflb7
Bp08vmro5HyxShab+49BfGkOKNG8FwBVYr5pUqQCkYozVJ5MbcXy8eEZbv/KiNP0tihhXslxBJkq
3SAfMNXqXXEPAY5ozrGO+cIV02d0JRfBM5Bdb10AlMIM9mak9464o2FH/9XMGJJ5OonbGre4cPrw
tGjVULwgCPaffqfN/w/bfBLWxMDpgRp2yIVDNvXpFa576iU+zUDVqG8hWnduDO4xPjfiKhbOI78j
TDbtoH0pLT/G03ki/5m9bzkO/DrEnqVhEXt8KKvyJF0bdvL0+efcSBGffVNvC7jhNGUKWii9+Cdh
ybxIJqd0HIA2aiSEQTQSK60BL4u2trCpLCxn25aMtpVrN5qf1dgqJRY/JlhPHyzfdegLjdG4DTdw
55BvJynmKfyKQqQJ7fguCWSa2BDU3t2xC5TQk73Ly+2WSatJIJpzmlm/0gl5BPoHoFfdryb95yzc
S8SxKZHajHgDkDDNfLScf2G8YG0s8NpSnhCzWmbqxEqT5RMX+K6nKFK3W5XmEhJZxCSGxNaS2CQN
ZjDlqOqmB5oLW2i0ZuEoJEyqRmLH0hFPxQ2SiLnopSxbAjujBTq9FUk6sl/OfQxz/OoF+rVvyidJ
xGnVEJ978+rhukT5MEQjHG7kr6o7RJ/URFPFcJvYTAC9Bk0Y3XgCG+I0qop63OB3Mm83MDQSHhqk
T5KvQK7l5Yz0JCrtjkkEi1UA4LzlefO+ohm8B6sH06zm7kop2z6woUHcXWe1ZPYHCPxMq2OwA5ZX
XZkNXj59S+Ua67RZVWsJ53U14guhbXy+16Fe/3nOq/GEJIiz7L3G6w1jtimqwOOy4AsHiUpKuUwM
mrL//dXx5vAy/I9zP+znTtHwORz+YSy8R2HxeLjU94qF2jI8zQIgLXKnqcHy92s10xa0btCipxnv
xJNozUAKwMw/YaC7La/DUUAawiAjGJgyUpwQHrfvKvAeEzaMp20CdCeUtM8dL3ysxxK5mc14TSAx
p/7rqvK6JCFxi2EYK+oCEYzvVV7wIoXPVbReJuDhNzQTJNulq448XIUj077e8rW6ti9LBPZSdzAJ
HGvDK+Fm66Bxn3GQOZSzeNMlL9pvRswZOlEZj7qJAiM4edHLBG77gCpDHzgs9r6HSPDoIjSiJd7q
bYS+zRC/mirffTf3DINAyR50ck/QtsHR6YMQWmCundbB3tUCU8nqTCjGFt2sgbaGphqZYLdciUc5
a1wmT/x5ILhdFNLcxzD22dyAFCaRuULJurmf+EevxAB62bPHTBtey7iX1l17i3Y2dMrHqxOVEsvq
i5Kr7iYR7NYluAo6FCQglWupyhc/wrgq6yzK7xRGg3i2MXqB+yLUWl54QO/fOAhzB7O/vqcSOYsL
9PY3QtERA59HPjQSX+d47aC8X/1REsoNhnLLXUaw1QqdaUlv2Vl3wnhVBa9cicBIHzaVsi9OkQg9
2z+hikFc2PHmEyafmVEv1PRulrhMP7cAVwhXxCOxbjG2CDo1FcxMBGahV4F4FYYeX/DAclHOftlb
X8B9Cu+6gpl/Et/h7tkH1YV0f0eqiKaU4kkQsX4fETauol32pSLrX4z2TcPmRV5wqCkw/GhVnjoW
VaIThAAJ+PlOXZgyQx7sJ+XJKKp6pxEr+FimfeLVdcRDoppHzrcP3XcmzjVWd4LbaxDmwuQJzIt4
q6jkSqKEp/nX8V9+P2Y1ov4cKLqI+kk/2LziM0fOlVZMs3AykCFSlaO20CPzyfwnnPzQCLhJltWK
kTjRgevi5Czie4OXXQnetNY4b00FZ1Aswt2VmSlX+/xfwa65Iz1lpvqqyedaKFaXzWaVWbgtH2yh
H1kZSLfmLXT5uFzK2Sb8Q4j2XA7+1iKRbMLeT1nfMg1J2eHbXWu6atE9EDJ8cHp7bdK0McypNJZh
MLna6ZcSowWAkDUgX929TuOMMqGT2xF8IcWpWq/7MkUsQWzgcbDj0GEep9jBH1kBKqo4mNEp+zLF
NVjQTXl3S/A94r1n8J69ubqhTxiWMdQXIoJ+mJN5YCQbK6JlYwb2OGHBgilJqYK3PURTcvQo6E8l
rl2550N1Ku6Xy6EBL+dsEJd5o0nB8BttHUJXc7a5DEYQTK2ub796/SR0uXAMcwW/ZhsSPf1gfm9F
vPknNf4Omj181LVGXeOwD/6+56W2qaWp0zykSzoclKdvYx1XaM8ZrZvMazWrAk1NujrejGvZO3IW
HjQAE8320bht4TMiWbLJbilZjNsrzlPZarmG9WnEtSA/WWzcdNx3GSZf2zhmExW7cowSVnsL5SDs
dDSpIMRSg+AzKmWpTjb8s8J9RfA3uOWzO2ztNLCS8do8R79bJRtLP+ya4eLmb1cG4RTvg/LMJYJO
apFznAqQm6b/0lJxibrcvLkxOE4czOtSmoC6uSTNJB3JpDKAgGSqaIbszDcX+mwHhqpwbjmsV7Ew
FKzYXSFN6PGztOYkFZeOGzXhklwdPUsDLn7v0nz12A84qG8eiQ8jAsJPWzq5dWAOlEMtPZdDKRfS
1AgoYWfi/Xak/FE0bNn+aDZOjerHUfOOwR+uVetjnP63NXfHmYN9EU3BHp/XkZ0Zr44bZXw3cUOC
nV5r/lKkLjTLKTQvNVecdL7RKSALdmTIa3tYF5DGeKs3gqwHQdkJbuBeoDyGj5ERebyHvnr/UFTc
RQkUlb7JAB0QDmIt/6m6+44dfljkCPmbRm5n3dSrKehKwcX+GYyNiM4JudF6PmG3nM9V4pk18dz+
ZsHH1RsIpd/5G5Tqonz4nNC5m8VF18M339bfq8EWi+Z9CIg06bYfLP3Pm/p0ksf3xqAbcX4weNQB
6WAXqB2p5vWmLwhfajICGGzzuqhyXi05SrHsSxvP4ai2pg8Ob81I9KzbTi966YhuOY+tihBuAlxF
8z3bgWJGZrcHIzwtERsgtyErViSMD3HCJQJjodsu+JqiTIHjBL37Vq2CrKDcorEcvhNpzLjKOJZR
q3Vojy5xMwBw6S345m+A8VBxxuij4TK0MsfHs2QaDaoDyiW8n91N7HIsUimslybsSl95W5aeMipN
5UbHs98mkftxZ9faU9ZtX2pWgb+UpZvIG56KGaK9SezGP79Q+OVOBoLWxDU/4+ikZwFgQqJ8P8/0
Phzak5HDTuSoJ4VHiGR42K5SHr6xY5olUqnGCRCevNwcmQmHwW/7zWqgzFepwmgkD2ZjyWV4s13w
sg9PvWy3p6XnKJgn5k8ft3QSbWgCtWJeRRid8NdlScw9FTqGkeNIj7NYjbg3+OkfdZxYSQQeFlYs
JkV5VfkK9TVH2Dq2jlOvj0UEP6tv/IGiPYK0exfR4a728OD6h5NGGuo8Q7gDLCeuSEK8OtAxVY0Z
ceME8PvBacrPciiOo8dN5Hq0ebqSmA1LFtPxvYsWe2CRYa+XOqo/+Jdh0C/uCxLphdQzctdf5++o
/OIaXi/THAfRcnI5t2OnV111nhPT5bnxxNzaos6WVH5/WQELVdW2OlJPyU0qcuupURRTRN2bH32n
QFsUBPWZxhlYlB7iCnob8JwS9TjNk6bQw7kLNM2F9AdOwtfIcgMYSokzRjS+H71SaGPwnChkzfaG
QVBmjHv+Tp4l+vy1690Nr+/hVaeW9IsFT9udIl/heyVcA1qFUOcbS7ivtUthTq8tFt8gLeKrTkad
wkGPrk6anOIhyFdMATkx5Gcha/O34IF89eZeV64ZIwrRYeR9jkwgEdJPrVjDrOoNJQ6hd3djNBzx
Img3nGAIXUUQ4hD8XwMtFFS0ZWV0snldOxIXKQ8+CAb9qjqjIR6JZ5MbGEcGp0A0b9o1DmrcrrYx
w4sMTWH4KEMXYFcwe7iBcVnd/YKZjEnlE9ID3gccSbRPoFnM65YTJlQpBW07MPqgEn7WIOjR+i/r
5yOTMv9o4dxrPxQdwzHy7grLqi5jWuAmiNySA/f6lOqJzz6JpA3uYYRWbuX1iFCDCS+FUnCno8Vs
dy9h2wpTzHdESgVkljY2J7qRuO5vq1oss13IHry+2Xvc+Qzdpy5SMpJ7+qmOxrPm6amYeWaip5Fr
q2GnTzIFvW7rWKcLKbwF54TC4dfBhn2YOpqhey23isTrg5cniwol2h0cJayKnU5qWvfzfCoLKtag
jsm94A9WBjcxk4UbsY3ME+pIiSeAShzu9SStTcidaUctaL8E22C0iLqZI1G2tlroLfKApSDT3qSd
ekx3e7accBFIv53jr8pzWGAN/MNT6METV7XlLaIGcjf/H8CNjSbr9O7LDUZErnrSVD0WbEQbLiNc
wJ9jiqrrLlPA+C7XvBs07SE2LgmXX5HQj1jR9eWikMcRjMSYLEMcObzsKbyWGFcYFLFqPb9Xp+U2
keeBbjOqtPFs1EFMwoFBNDwyDnpV9pGMTpAyPQOA7GMw+fEsO92KpbRvXZlYRaELwW1XZQ0zmG9G
TQGc3I5PJKfIkxn2MV4gXT2DS7Pf13tfHrZeGAH19huzo4dp1usRCqQUN0pO4DlDdyapOhwwU7LY
6VOfoQBL6oXLh6kVo9Itgm0zLEVh0fZ87AUSWif1qVJSrVHCDUuls3mZeGhiP3ClisYpaXPbGhW8
l17lIEAWvTD7fpI+jmzXl/5zDS/GuSDHdBmkbI3g0F3Fuyjm9lnTy68Yrd91JoUUV8N9BtNAy3vP
E4rfqm0Xfu07RHpPvn+ws+yrPwRF+3eX18qbc1JKjP3oQ/+9/N44/eKBipxss5eRe/z0ROzIEYzC
ZXcg4g7FlJDP4MgK6kA77nAUNGGTrt7AWhHimGz/Rqo7rBY7/svhzs/JmOS6TjRn9LTipVMOYKC1
3MkHh5EAK9V/AgLMEg+h0mvMftZHpyfile3o41qVmhJNsRwk49BvJn6nMmbovMHzTyMR7rR/gr9V
LpVOVinp9Z2whQsuB2uU1/3fwnBi6YeU+NM/AuAnqMlSDrBZ3PP6ir7oJVExz/InJDeDLhGFqOBd
qrKZJWc1W5NfqKiuWdh/r4l+8qim86tNVD9/whwEGpF+IFO/5VCzcknA4uK6WOz/R1adGzr289td
O1KfDeOGj+Ibtdr8Tdpe1tv9qTxBnVkRgbPxlXYBjB2a838vjWxPWBUT8/UZdKqU3YYY68d0miPJ
Kiv+WNXfnauDIcD6c2TH5UI2yuMPZfvV1x4j+hVloLPhorzUGVx3dzm9E8YRgXOia9ihBP28NtuS
IOT2uM3IfSmelhCFEKnlL33X2si/Blnnqu+8ACUuzazXVe5maPY2jz8+IFrsQ90dpvy4dUDHSmId
YtD28dDjRBXRpxXzuv8lNZAQdr0dtdM2OBokBz+hiF0TEiOyr3TFjjBXWrX4UIWUc9QtqQ6Igf55
x2LrfnpzYiZwjTSVg/VWPnYNSLfDFFF0rfmbQoqAS3B5dPnBZ8uHJOVFO5XfSGw95CCEoAHcjOTI
FQjfUDp967tH7V+tbkhfS4XYaXm9zEEqYBCtB6e5xtYFHY24xCmaV5E56GWJmnMlv3U5p/Ti+ndh
VC6NRfuO0VwvkyQ02FSxdFwXIVLeZzjEbfeb4Xom+igHZ3Nt7f5WYY3PEAf4o8TTXjfnclT6nlhF
Nx/rBVjCrVnsgsDjKpiPl8el1L/AoOu+yMg7SkjheeWrrWiJYTJro/iEDLBlMs5nk3O8MXnquBHb
uiXILLzRZsCmuNZK/0oLFnW7xSlBk8vlRPs21agHP+VboRGnkZGJ/3QBkfBJf/5ipTozCcqFSubd
IUJ+FuSpKZGq6B1/j/rTMam9RUXzxKdpSIh9jOuBD46TUJe+/FFVzH9Gof1RBLmaw1xuMp8iOFvk
4WIMTvMp77rdyrV70ohXi3zOqHHsqWhgTKVpKxJwHuKk5JMwYYKOeBvV6vt5aeKDokwb1g6d/QlD
Jo3ypUUWqgXN4P6LV3MQHQfOQGj8HNSmpyCrRoLv1DGdCl+jHe3lgrTiv54GxGc45Ax2rbv0lZ40
WfPGq0otMLUnBatQliVahHqrd9OZCfk/wuwtoP4w+NBMxtIYlWdkOSSyfmWJU8oJ4sCMK2HBY1Sh
zeoHBA6hsBBg/UbG8hqjp5a2M/cvmANTJqHvbZ1gch0sTxY8PJ4c9ZCICjolQSykGbOYZCqPm8vZ
DPnxF1yY1XkLQ/CwDUH1le4NAEp8Mq2IEAoOv+2ZFx07PX2tsWGE+c3sPMUXwnHPLlQEUmUBpzV3
z0M0iMt+xMjLcCwp5DQX3+wgRaJ5ZXf3vBbXsW4FUUu8NxpcSjvU/r+vVNjX5dDSmBQOQgfBBC32
1Nc1/wXPuXr/uq1ueVRECuJ8OlcqQBQqXmNM0I/UoCaj2v2RGrbZsxScQ6X2WY9D/79Iyxcj9H/+
SyKesot7H4GA8YKO66SkxKqCoZJSnLJzleVjtc76+buwCNSC41E1OWMkG9Fd2d3KHDKwiHt+8qWM
TlSF5L/GJL3k9m5Vdu14AQMU3icfdc0RqEcF6OLADWStucMDs4ex53TLVUVgZcBtSU1E3nWcup32
O+I6Y9gTKJRs8X1zU627xhdU0sx58/QdDgOdjefDvRXqPZy+RCIobIBXB/drTIDyMVTfrjgDA2jo
ej/cDqc501x+62lro3jUujmR2hz10GJJ5D0oZHlJuawYcIZJJP0G8CeKkvpAAMYZiwW09yrgybIM
kk8IO5+PixYyI/tFi9/mqteJ6CIrfiT0W/zYU5JHtnH3OErD+lngcqFlnKgDS5C0kswVdn3DM8c8
f+HQvDHjv44c6vR1L7Kc/EOKiJYibhgV1owhsIyjLJCG4vJPChFQfFvTFJd1ekrGh8iRvjCRUcsr
bV6ROxESk57MIxkiTol9xvuS1gpE+SjVt5wOs3AcsqJDZJLtWK7rCz2FIvaPGDFA7rJ8m88MtqRa
ouIyoe1sRLHiZ78PCXpAcU4hgBUNG9aX4K6ZlLRNfdCh/vvAC7FSWmhBatoTv9eIvyxJ4uA6MOC2
upP2I7hbxS6KTKL9f7bQeNCVOuWjtW49v5QU0infy+VWVEo8vDWqB48H+Tn77fTaTkNdOcTbAf/9
CWfb1L8sUurmDSCkUhRm+t7g/3b6jx2Et1Lni5m6FGAtbKZYO3VFMQv5abfVDovYuUFzVyV6VHdN
Djm5hMIua0+pwgIdrHvSiBLUEQ5w40Q0BWg7sJmVtIEIHb1cfu6V5JuGoqGOPVz1PtroZ2h14pWc
qxC0iHv0k5lDjGuAZh7lxSKFvnQ11EVJdu1hBQqKAKjH14BbT38EilIKq1huhafBJCa7IINiu+uq
FJ7h+ZxwoFt3zT7i7kwxXof8O98yprN3NlxwbDlek4OP3+CBDEzbIht/Bi1ehnxpOekMlfUzVTqS
VgTKK1TM7yGXk/msyobRv1dJ+bqDFhNr1pY0WfWnohpyoOXvh4TFYX1yJG0yxEgxId2seqDxP5Rn
A91BfZbvk+20RIdrfr1hLmqxR70PKg448Du7g9gcWzKHPzpi5ouKMkUhvBXZhJZjuo3sRoUQMafl
xmR1tYkpkMZh4DyWja9gyofsJYsLi8z6G6dGGIZerfSHolYcqHFe7RgHRhm5alMulBiykEZ2WXbn
hUGR8ysrDi9R+cXCiIgX4Yaj4LdmneqhHq/mLqWf/75MpfXzcM0251u743j9hNzgalHb8X19qgyu
7KVS8bt929qkyAn1SzT92/JQNm8pjG2A5g0gjZiW6Eji721w+D/M7ou8jTRuj/dwffJQltQR6yEW
otHIJYFVHONZQe9YLXJOKhE0zLP3oXiDOB82hIB/XDLrF+O7yC3tx2f03anEQsM6noR8LmWTNhae
OJg5S3+KF+p0R8wVMhPVpP1dD22JVjpbnlAyjpxGlaNCen/r32jAik6FPg1Njn4UfWMfJmJ0OtkP
LKnD9rlcXxFYow8dUuMoRtwF5QyxE8DdfQZ3G1eQv8CdAecGjeNDPFK7XaPaGjJ1in4pXdFowwkA
96z4ewNIlIV6Wun/01opMnQ1LzVaZyqVQIUAU2aR4F69A8f1PZ8GPLSHqj0TtfgOi50F9fU8ETXF
3Ie4jXOm3oTZE0xtxDELIMumu6DMd6YLsp6FRxEKVeyv3/Vq6or5SoZg2Vf2IHL+yc6m1+uiWckV
Hk85XgaKtmI3pxyJQWBA9vlfhAM5yi6S/EVxEd1eM5TdBHDK5HjaLaYMCSOurnBpMCVjZzfy15uR
He9EPI0QGMYieSjr2JWq9iNRnwK6YV0OfnVJfR0nQHhnoLGkhb/0d4p3236uE51urJeqmILxKIpm
vv48Q3vX97O+UBd+nFiSIXvhPL7Yodcgpx+QHa5MWdb/95AyfoQY6RWsK1o8ZuxvnqRSl26xxTxU
9uoNva9GiT4/e3q0AvBc8J8tbT5OT0R5vyhSsQ0s5IwvGxyoAny9rd5dfgRq+FLFBIEmoJqL6ONK
YbQodzbSNketPzI79jTT5YQUkc8Z1L/9MAVJxx2lfhcMY2kaRYxApQ38pwWRs5AID/M54yj9Wyqp
hKUR6MhyY3djWbt9xTmbGqIkLWDjr+4s5hErnITfbk2xucq4bks99XZ5T9DoOF7e222CCgXVasW4
hIuf10ofucaTT2Bg01PeRRpWF3eoiw/FKWR1VDu/WdxmI5GqKC6wbO5jyMjG/Cg+GF3DSuazzH4e
NhBPoWd444i+l1j8EECmyjgJrjUf7teoKZ9U1HFDM840EL9olFpaEW0wbZgZW67WfA1u3MwNAlyh
jWEPVCGrYIXYR6ONle0lQynGhz4xE2ObKz5jXrE7J/OPMnX+wIWbjq3HgWAsBg5bz9iHIOHKlkcR
FmidGkyZUMkW58LXv2Id8ikY7YGC4si4v4dWJ/mYf0us6zTX0VEcEUCjrwc4U9E4D6o9DkCsq2yA
lyFOmH5HyAQmyGLBH4+1+f85xMZ1/cGFuO/nQv8baNdQZW9wf9TTC/MkTif+FaGz2C2KQL/gBrjN
SHtF47HITecT9LxGp/1wB5CK8Fy2w7hfQRJlKF6ZiOGyVH8xeOPP2Rq/qMEhrq0eBfcNo0LdJ31x
ZG14xvkYOuDUNoZJ597y6wnIAu5kMrg9dV9rflwa6B9NXLGUkyOv0HuOO9m3IhAQuMbvUJ3kbEt1
yTpyRkjzQgArCjz1fWMM6qfHxRb5gLZXhoDjoXSkberHEDCutY1UUew2PCIMaIPjSkzfXLAXeabv
hxckRRi9Nfu61rxqQj/ZvtPzB82lQA2PrWZMODu1e+svlVcCGejG/Xyr8qP9SuVPoY9RqxGN86+C
5Q4RkJE7TxJdTWmq95a13Gc7To6XCDlArjbsAoDnTMhVloJT+FhDw5QbcxYT+rZEW4Ux0zhTuBBj
Nm9c5Qu3oKwtcMfZaSaHwlgKFQQZB14GkJ8t+qngoIuM1Dg5BZebyf/RuEXnmQibkoQCpoZp9Dr9
hpAhOgAyxWgJdRWxrCglURumINLd28VxgKb1vjp9TLzReuOGxuOyQc4o/Z7sw9s6eNHe54ctnG8x
/Qzr90TJUZPUcCiTVhbJPW092WtHWA9gYIC5SJfy9N3wIyGUPeryemKguZdvyRr4r6a8K7jmsgbm
Pw0uVsWnWt+G73fl8KqslEEOOwHniC0MqmJqI4F+oWVGBpjS10AGgLA7OxVUf02yD13hDQEse+vP
AF2WXX3sZobafXlCKa7Nre23UEP1sfI0RmeggJeb7nRm9yMh4u1u3pum+cvaP4dzNnFBnpVKi9cq
QYtWMty5J9Soraz9VT4skrA2MGRaY28PSkUW2h5ZR0HNkYlLvkBOOjoF7S8xq4zjbJr/K6r5Tnxc
yrNWqR702nY603LGelHNzckwH3BYboqNwrzub3IacJ+5wvBV1LrZ+CVT1Kwv7X/1gnsHJUitDFfM
GXu/GSwYPahw/tGm3LObnuWfambqaSLNK+Jo6m6smBQYGKDJjIU92dBPaM6FF9htxfSxzaqE6xme
y9GO/kAkFdaEdRmRuwr6SzwsqOAYb71h785Zc46hZNZK9YKtpb63DW5FMhr/2+SHQRHYqcdnf9Le
rWbsTRZYQRoY5ke/PveJjMmt99XQJjuVE3uvGv0IoRw451OBgTb/uoTMBQEUomotf9vb34Z3PUWk
Cf+pBM9KcfSGbe+FKxdDDNBIRL/zilnJvarIA2LmzseKv6JMJ7Jwn/FhOyQ0pgSjEa1+DNdJCh5W
C7OBrJHEWDH6wKqCOo+MtG9DRmUCCUv4s2rqzHuP9+MG76hgL8NfvzBcdT0P1P+al8DqVlTlijrU
M+AtGoJ91t745NcOJ4JAW3lf+2p8CTMlmwaFnOyga5VDSrApV2oUS6m3WOpJ/g3CfwWF5Z4Zm+jk
gVSJimZvKCcDdv/cqYo9OVrdW1epXmQvNSJGo/v0BO1q4keXbQ6mYZQPn1O1Nk7MjgaDVzBzf5xC
jzHQfozFv7gYK0zRKiqkE3rcaaydCmGNakQqAxMc7f2B0lEjrSEGadY3ydIhdsf8FLlu0vnmVSb3
Lldg4CPMNdttTSc0TXDaDNoM05fJyMGEIY96puwi5HE55wkc+ZgnNtHXdZBZftf8OLhNaL5hanb4
hvSH7JxvdhhCrn/JUr1XP1AbJIIe5jjH5Jf526q5PC/GSx5iUzXn99vWNjNnIsrkwpb943kKw+VB
z3TLcFCyIwvZ5AwogzR9E28ch2407BZ9KyWV5yO//GNDxDJVp+wU4/0p2H9MKwcIpuY+FEew+6o1
yHuOCdioxTxxP9Lh2El8X7ntrMjw2a35JNVchTdx6goIf/cCXx4HuvRkouoSTUZa1xlkZnKB99IE
DBUExYVh54mRI+lZTLnKWPyAtWSIhx7Ip5W3JJswepRRyB2hLwXGBlK2wvtuDZ+0csNCYq5zr8CZ
2+/7/CAJMZwhdag4Lm880rB7Gq+nAZd9VSUQ/TNVJ2bJa8H7g9uNJjYcRTXHM5w9arc4uqpiWaf5
nQdWYxZzJ9ZyjMdQzFTcDf+PROxuKyHmEPPfLb1Ni0FWhyoD11MFA3yts3mZe+FjUH9sKB7zQ+pK
eNPL3FcE17J+dnx7e1B1nlT53qYeIPT8NGMH2xfEw1lWZkacqzclv0vdv2b8AzQFzMxbePFiA/aQ
AOZqh8vwOl7/JRrsXxLiuKfPKSeuMAskf3jHwMt/ZG1OKT7GlK2UbiVjG2hWZGLRyW0uhYh43cK9
tcTNshqTDmC0edRP09TRL00RBsXDgZNayayMRqJluUKwM9vtqSEa04K6UlbBgcEi6iT0i+drrvJK
CT88LhNHi81zf41njG5BkjMfcFutyH9HnSk5pjW6VZIHqpQvXp2y1flyOF/H9LHflzqfA5FtwQkU
idYgQBZWrl3knEYlsZRRJExO0JMB4oyzjgCgUw7hLK5FaWEfL56QQgxUJw8GSSX6ZBweLIkKY/Y2
NOzfZDWthRdXH/R8PTzVDWm07HBqGU8/e1oIZszwWRNjocU3TjvZXIpGAKysP3t9IidPyfEKi63/
sxUTtLzlTz0AyrxPKhQetO1re7eZdmZXd8ShmROPm5xhrO9YmGGSNw5HMaj2QUiLoA5b1Xwor8VA
DVazna25/4L69jGoM02IMq/bZyZPsGhaM7JZAsm9sYYj4yTLmeIb46TIokJ7QErgRnlZD6jwNZXY
PzElev9F1RRXe1GuSz1z8okgXNpqjhhz+14NMPrawPbi5bRWBVoKYaCKQnBNVg5Nj7yhKHa0pb5J
VSwMh+TkCthfP1yLPip9zsHUYip3hBHzRI/702kb9p++2zb+09CMpUi2NT/jhxeJq1ELC5H53cqp
5tOFTq2bohnTwnqHh04C178l45fDU6H0XvAP4gaA8jxmNb8o7eTCb+j72dukUf0f93RD+EGDb3V+
fCjD79JQ18I2w68P0MP9q+wSRK971Js3xspKt/YLBWrgHhdHkP0hsSk+o6FwV/r+vbePK7+5Ylyd
HSWebqpx3Kh4EHo1HvmSns7K1ZJlCVqs1ps7s4J6dIDrNCHyMwQxXVOuzBDF9ODriU2HVrlNy7mh
soLyEi+Al7ZQSRFtClD8Gjl2NA9KPwawits/sHBxr0AbFpb6581+dj1kKgB7dtl2uvxYF1RPIktu
OH/YpGBeL8n5WWRli4Xkg+7cXQ2UPk+GJo7DSCc3krNriadKXzptEOhEm1LQbtug/q9rPej2E99u
tVANrSVWm+CY5fI9l71d4J4e0PU1i/r+8OhqtijlUbc+HjKnI/bNCLKgo1X7YN3fX7Lvl73XPQz4
sGGCC/V4PBonvZqyTsfmr0IFGXXwr1mq7slxu2uYRWbMMxta7f9Sxz39rHUDvKjXmy7amsvcNKLP
uqt/SR/OX1IhWmt+rf2guHMe0wC97u3iasFlZJBQaFf/LOZ4+ZtQ57fWPZu0FSudhgv6QmbTc53t
ryQeLfWuMZN7QKcyZJr9admDrEjVrWKfBi5UzB4FnJwE0871pVls0wvI+FSBKf4Sj+J0ZJ6Pead1
Yw+fb525zao29z4YT/AfMlO3jfr+zbiL9ahuM6GSMR7+khEMNVqYXQicR0pS6VkVoGPRU6kBFoRa
c08PACtEXsJ+jzJ/mDI9IalYT3dnVXVM6yxGl48hoeOjK+f0qHcsammCVcnU4IvSpeanL8/KB8i2
GBZWqhc8w8ofl++zW2gLFxAM7ZoCVtbRSq7t5Vmlg3i2DmIFL7P2016/kCGfQcpWPnJLQRPSC0Fg
PInZfoDJlW4No8Y/yUzjV5ZX3pa8+38OxhFpZ1A2s8WpNPUoAGcosWad41hl0ThuxPlf06g3wof2
30key2tUpNpPa1UA8KqSxjtaLG7eK1k2JSINbdlUAlIsd22upLegUHY1I7U4/3kxpOdUKXgL7Jg3
dga5p/xFNE7Nfhg9ZRPj7kKuXLr5DGxsTuFGjDOGC3g1Pk41Lm94U77fcMWS+26mCpajpKBguQ8Q
aN1/qTD4Xrjr2bWoJXvbtgRbmaS0hl/S+3iiF/tlMrpaewcRl8nrxCC30VqALZYXASlOXuytYlgs
CJlw2zR4UPPz+uQ63DulFezjJlTolYkz1Duryaxk2xwJZq9tFJRTzTenu00uc+5QETRKjCAdoETH
jbpRCJ+0DGUoUSbIp2MAohxE/aFcaThkDWc5hp0s+v2WHT7TdRTDG22FRyGOIcOlQcp+/kf23haE
uh+5jy7E1AKmbCsmfPO9+gchuvaoqYtWRdeh9Gl/ipAJ/XQxHRXH3nWc0uKIU+x6BMmVQoeCwMju
pIGegalhVaNmWAXhWxLMpfIQt86wlgLFb4lqlNxuF3c+yB3eZefyezsOnlqmX+oCocrUc4RXms5A
oYHb6CzNPnd203dHQa/wTbsC8hrs0TwZi14hpf56d3I7TI1YyfWekyn40ONTB2ch1I6TVU3iocrR
CX/ia1sPHZG0QSw5JGsP9x1dw9Fyo23PDlhXTVgGtppq/X3C37e8lRexHfQOSnPl26/u+5opF9gD
OEc0Q0HjMbKQetpTjcxXsMb5TPDxW6v2p7BNMXe/T9S1lHySMKbEoZX3AUURO7s21e52pFky+0sh
dCHvC0eQTldAV2s45Cn9vNEMfQV671LCg/6MSl1wDI6BHsADeawCtcqqs5K92rPEALY0sIS++Vvz
tezp9OhHOpAYO1hdCUJzZesmIxrR57G9e9ERFkMVBEZqubvfla22FfCwtSV5j4n2YIz/upY1/oQD
xM6v5vspUcP4+EO2x284+2PE6gmhEFkXToaZSkaYduZtEvPCZvWocIgs9PBIo746pFk2pZXkvrKb
lA72xTgJHq/p+wYyYc1M4LX2NjgM3VHgcpfUqgtW9WIt3bCH9nBNpholu/388toz6oXUESqetaPT
LbvPEt356bIatUYOozpBodmP3OXqyRuw1Y/mOJmGIDm3EY/8+NQUroIcKpkIXehNy4CR4bSSLFCZ
9P3huu9mgZvK5eCFiAOsHFYotKqJ3yaX7MiEcM/Enn97RVvi3C4mpCCRKYaiWWnjnb3ZocAlAQ/w
PF3kdbDZC3EUrWK+NKIcBqUqgQ1TjIdM/TwVOvJa6SugBL4iNqtP3lfy737Bzf8Kgr0uaa1NmIlt
CEbGxyUm4C8+xIFeDS6rpwzynngeHKfjr17vJI6hV7KMFARHHHyF97ZzB4gGA+GkmJ714/oYwJiv
QT57DhGNGFvoqKxjP+eywnv0ggHSU4RILBcFc5Em5fTixAVTf2JxO4v7miPeMGlGrpsaCbFM2H/S
eQOUwM1tVXjRprzY0SzIga3LnFxi+P4Rh7kcnbp0XN+Gsw8HsqisxfayhrVge7aVPtoZ4OYTcRov
2fX406ewrrQmWf4UhWrzPVTui4whaI4Soy2IsNu7C/Qp+JpX4bVwjeN+qJD0uh2CBeUc3KJlp2cJ
+iDBMoIUiC5oX1TimufcFiydpcCgqr15i6MVjXLyBvqUy5SlMaheVeNPocIgTqV5LJDfHGLGBQYw
bqXkEcSkF1UPIeQcuEZeN+EhA6/EobV3EQknIk7eOTru+GwXNr/H+/dLj64CSmpuR/Je2F/phEcW
BsFs+xI/ZjgYCs6zrcb7CvW9KOApqIPYTE2JPF73dNrwQYBG5VqsVvTA6lVZSh0b/OVdoZ3OSvZK
eHXL4ZdYAyEeof2Por3JYCKigDJ19eyRnWHeyZ3QSG62P8t7HZ/BVqXgBKr+H1JmXNxtCVF5MH5B
+sLLwGYVcF0zxZqQ6c4jwUdEF9kdR33jx6AVz4P6k0ARzGZW8T5NHPhhPMNFFfom1veaUcGIILR/
nnEpat8hhFuH0sxKJ0BDZCXyn4e7s8bwBMtzpqo+ToR4VXbvhU7ZrKGkxPTAZI3UXC/L8okUvhi9
bufIQJPNFSFvM4lNib0Pq54awdqdzvNC3Yfzu7uP/p6/r37MpEK19+WafTEenQ7hdo+GeGoonm0r
tPI3EZ9jOsLU8mhG4G/zjW/jsF57yCeeJiVni683ChxDBnCYMyDh5/z5EUOpOSbToXK8VPn7etG7
t9rdTgTbdLR0WB19Ddo7nGd3NDeYNvXgWtIFb2g4JgV3ajdsRXNl7IJlTAGmyNtn55pD9WjdyiFK
yvoeuWR5l1bB8QL9XbE8DCsq1h/WG4O0TF9kBqxhtT/lkJxKTmnWA5DJWNS7MDNtBnBilNOjcfsF
nEbroX0a+XzPgNcbj/tpqZeq2IF3bykq0QlSGGlOeaW9vLGyLWlX9zMituseb9jJTm084QoKQoXY
tk1ruLqgTfomFjYCm65Jqx6GgvUqgnFOygc/qaPO2/Mg/uaVb/p9Fy2vEggzDLECE3mdfT/NF51k
18GJ/nzk2izHWwPTGP7BX5OnQ0nNfSKqyW9mepEg/fRLiwJ9NVShxTsDARe5c6jK9R5vi7zfWsLT
tKTslJ0vRsibvWoOIWJoR5OyCxmFebyYaRD589TfDTt/u1MejNEXCDwcrE9wNkmfLXJiawtCizUk
/2Vy+GS9mFK/MD0FBEH0ART33FDh2F9BtBNnBWhdVFFfAdICtXNLeM1gfdia+0V6nZXbYlmiA0/8
gbrdDmssNWUNC6pPUnz9FpgVooS0vGR1RPZTXVx0seELanj/O1YILje8xXiZOjYQEXVZml9fCgnT
w6GMDqpVOOlyIOtTuNIf8Uc1o06uuTspKVkDN1l2mRnLnH58isKW2fyTKWMZ61oYiUsJfCaD2VS7
lzH6dNcKw7PZZIJJVf5pcJKrnymAOl2UwppRoGJKDK0t1Thj3t0k5Ekb29xXk0ycPQYLxggPm9iD
f7nC77t02TdbLfnH9MDsywzt6dLP0EM58P3aLKxSqTlaebNAdbSgs094ijHYRF0SMcGea6c3KoNx
u9pOoFxSL2VZJTt9ygAysXygzsfpjupC+GGPGZEqmfMhz0ZoZubwIiIeqDBHjxW3LbglKTVQPTG1
uwRZLC4h+SvGzX3VfHo9hFiYWVPUhYJwFUM3ce/HOUZqLbK94XVh8QbleQSImZ8OwJ9v6Mp3l5TP
7+Ek3RLHdyLm/OJjOcWPMNm9JZs4J30gh7V2ZlQ14QGoBR/tESpZGIACZzQljWByv547BZUVp+z5
x1wao/54mvBKMug1BQNb2lGAKqEjUcU8OuWOvcd2DbQrSM5bPIEl/vKbOUrFrfms41HbZfUM7MTS
B0UFZ+n8rJOVkRXtKYyp5Ypv41kkiedf110BGfsqFB9EsPq8bDe9BOEolp3Uo4CMFHRUaaLzuEQf
PcFwdKpAvVoZOd64PuSULz/ajeIjtr0RC8kXAxF8zqHTo+0IDp6POKHaH6NZWYHQTi6BkkH+sLRb
daIVB39WqGMbsASp5hYLDOf0j9QH5oFEeDr8anjSQRGOBZTW23HNyYN/AEQJtYLElNR+8fp5hyIO
TkMq66YOoS1zSuhS8ITXvW6q1mAKklnMqH7t+yHgU1Y1rgvcL2F73ksTAShkwZ+7jbUNUqiBcZbe
0Qvb5ujw5D4cPaBwh0z9AalF1gvALlNV8kHrBWbrVl0aQN0BsDygZnhIV3ZjAUB7Rlii19QTwBGq
kliEgrdGDXvI1jBZfLhjXlfUmkmiJnMfhjwCWIoCMGW3udolYyV8PKpvFUvaQLnbw+le1H5CUT+z
fuMkdq3gD8gOABpSrDD/w/hISiP0YeOmj8MQnM6iM/Cc7pkL6vY9C1snIjJ4ydU9CYWUyaxClDaP
mOCqTIOieZUehVHJVMnmSrO45qiwUCNxv1vLsfhX5EIWR5Y7xubEWy1NzIqBr7Xg5nBiQa5pVI/h
b4BPjLOCJXlkp21QW4/KCI+xk4G10EPsuGGU10jC/AKza50C/nsu+bEcE2/sNX67A8dDy91vLf+t
B9ie4K/tooobxlMliojBzbzXX7c5Nmunl4s5/8I6UE3beS9yQM4SvbqjHPr23C8NqiAX9mmR+kX0
OoKHG/q7czGbSUL8VDe+fLhTQed1fAQzOtp7AwtSFGfir1ciY9NBqg2w6pvo3awUC2lHwinANw93
kKWJHgg/LTSESlQEbKjVTHNdWSDLS+OFebKh99jpJPc4o7urZIQml9VAhxjcEZ1jMkA5C80GQqdr
z2eP3DTuOfCUNIpevp2wkrPzkgpnBch53iKsArILN4HBlacM+jHQyq7e2APrFaLiQ9aygg9px/Qb
VWQkdxdM5mse4OlHd+l1IMp3EYcw6AV9CFHaxaAZ5R8VNtflUavM5qEmoGJ9a9mkhqbdCL75FPwm
8osKukY3w0piUu9Ge76yOsYb2M2f9Zi0JRa4pOeMmjlLsaOu4BtyHq4tRCSiY+KvIQXiiO71HX8J
Wy9lozotjZlzYLj34gd48EnRG7mmLMDW5Q6hLp40eCE6wryGoRfSdNR20aHOCEf12cAiOfzLsgig
sfjj3GwhU4SXKtmwP/h/4IHhkxLATr7NifWFo89a77IO+sHMtSl621ddPcBaWJrord7CJRBumlCb
oTALxrStF4GVpUAgiu7ue+sr5w03VzKB7hCw4Xkc1GchpL6QSQXJoZ7d4e1iw8WTYUnsmRCA9vIL
QtxRWiP4HkmWb5h3GubIbGFg6zRUObhOoyaQlxINExBL2GL7lY+JGsS6inz+GsRGTQVjrFCTrjG1
3Se+cbnAZ84oWxaHEqr5G6zuyBiZkdA2x8RjypuRtdtDbjL+N1bMj7lhcPGXiRVcvy1pF5wMUe49
gLzUxiTmgQwxM6tMieAUn0J3yNc/unXYYANgrum2+uWOF7av2WxAdPpt1JAnBthsyVA7n2DNo9l6
6hQk0mddPd8vo/HsmYWbtaWrKhvx6rVVbAUfu9YzWojs7Qx+tdRQIQlIhJ6NW0YCpJ6dO9JKyc1t
V00ZGofMz5IDt+WbpWgPdX9im5XSRUADqFSyk7hG3icJ1WhP6zgCcB/JWp+Gv/VfM8ojeREqPATS
m3NV2ojU5UagE6B1boioVoV5YKA55fqs1cz8jYHh8dzjnW8kp4d/u+omwj1hcAVWA6xHlcjsbIR9
X4d1v+TB6Evckfw1/8h+uIu5YrRldOVdfEtsFik94B+Kx+hqfCMHho9T5A+7Zzj9arOXeMd9l5Jr
7gviYH7NdbqPaoK/pTu0Q25ZjavWvGL3UAApW3JZPKWeqwRajZ6Es9RzhoE9jDkWkaVbLa4TDIVY
HdpQHUB8E6ZVF3LtHWliZVxVcMaBxR9xwyOsaDcbW4vohfNrs+8zRt0zr/PB/hwRNdjtpHhwn0Lo
C5GyYN0I8DCo6OK2zMEfG2U676Bepqenx0edB6snAlSGku6CyR/XpT6o7fBkHW+JdJ8XuwX48QKb
8leCWCZtkdL/R9mZzLSusWKT6PEBXot9iAC+5VIujPNP1ylUja2eF97GgctBhXfHR0VlEv8kgBbG
aw8dXcsgiyy8u3JGUov3HIYsP5XS6c38S7BiLK1VH9YijJjuzh4c7BvEc9ijT7i+vAboDqvwxAp4
1zts6bs2IX5bAgae8Vf7gJ4Py0gK1E1hCwr0ux3aQcszaPg9UyJ5ttMBgf8IYZZz1bwkF2SJb+Nw
n5MiHiUEZ90Rzgj6BRCMvPomnEUU/lTNy2S1xw6NkAiu3huEfpg8+akKrLrdbGN4Mwx9H7cFZtRo
Dn1d77CbzGu/ohmhLMuJCDkFrNvLqceBUFnKBl6Q7BM3UT7L1OJM2XLWWspUv160Z49IkYqHMIjK
A9NST/ue1dj7wOH9HX87LWSo3n4sGM/nD+kVlyjOGtgQjiHpEsF2qOtt5xbtTNUo6jJy6XxlPspu
wk4beiI6AFvKdjwou6QEJwc+r50DUtv8gHuaeGB5QgMB9q4hzymhIXnqkeY9FGzigbzzLld5uYn1
oRU82RqQsQezMyp8Gt6stzQPHcplA62B3C022P7UsKGA5zRU8jqA0qTwOK55ipDFoSzbf9F6BRZW
FRUyZL4LRhnTTiGC2pgurHsL8IxtglaXpRHLen7ZzbW5oLOUcogRCAf2Uizg0OHOIQKY2js40KVO
VlInhc3sU+hSHQHVhoecmTHtQRk2Eo2hPPdJGeXK2w3gwnRxHWveP4ghbjNMzStJWcTIrnW7K6yb
TstMjnftEYHFL6kPBAmZyKK9YOtqB/7Lqgr9JAbV7DEav3P/nYwsHFd3z6pir2xxJqlnOsQ4RODB
sBnOpvLtmnTCWG2I+NG6zqoQy9T6zMwU0+C5I7Cu32UBNUwy/oTasRC04hj62FU2G9DkI7+GQ1dV
EJk/K0JeefW5kfrndNIS01GdeDKZY8vAdG5GGHfVlU2sqHqz0PUajIwA6xP/14qepohrlLXweRHV
lgW8tUIRyRLqBwEk8byPdQgkazMtPKq7tbIAV8nkfXNIYe8EuXWbWF0jrWnDgH0xMrl5qfBs4TRb
S3s+TrK0Z5GT5zvT4jmUb94CEXZvzU3kE+hZo5V6jUNXBYvfIJrBiqhIrfV9MFooSugNrj388BF2
9sNZEReJFfJXVBSyE6TtYj2wDz3rtAWNdbDmUc5Al9X7fopZ7eYL8J+kVSHUAGEWnRcnRrO+MQlQ
LLdvF1dyFBoXvjendp86RG/MiSSugr7OtmXKzr2z/NwTSwYqVAdYgLS+KY/bxBjqPmWMTqJHTi0h
V1/jfqoth7RQXXwNQDaBcF/dhgdEb/sWnoE59N/Rx0VR2EKNAx+7tPVSzm3Rk1uqO71mVBvpVpz7
w3j8QFbmmHVMctMPsMYifnqUJbSbQRXUj3C/SylbPULB2u3H+qwib+3sw0QRX1TOsfENEp8IToAm
5nbprHKnWk7lpHUXAzQrVbADFL/pTK8zK39UnLDXJc7Kb4MG0avU5RdODOhR/UQ1rB3e/U3H3/9B
7dubasRJDfHOvfM4fP+8+Bq7s1rLnwxvbDNuI9uLQ7cpnZOTcosWsQEaQdk2Y2n/jh7cjlZ92byG
kpk0fjqwa8P3ocIVHhQXJD/TNOYV2eMe/a5StBxFVYaz+OnXveTydAzNPkZKeRDRV0bjb8v1RWzF
k18wv+YrkbOrzI93sdA8vwm81ZKDT06M1vsT41pENp0Ouxpjc5E27G79pv7CXLZAOAL419/iug/N
fs09qoaU7S5acJOMQx2V52iOwfRQApWFVmK2Ag6dj+QPdF8TB03w9vdtSTDdA/u9NaOAZGp7x8kW
YyV00p69euK1e3XMdoMS5qLYImDp0GWMSju5jJdFGBsSlXVvUEtukmXCw/RPEeVEGbDZl17o6FLb
xHHPfSY6tBnf/48eSCHD+a7RguYwZtxgmn+Ipfoep1bK9BHq72yay/ZSh1Wepk5L9goB33zY0T7B
015l81WZNQLpe3tjAe+vyv6lt81oDgOWvherK4Xn6GmrniXQZi50zy4D8OtgDz/xVMjxmA94vcc7
6bnKz1jgksB4Tg+RWejFYUGtrhd65Na3pabaLM/Z93PfzJDAEWUNhKqWZDeMwtU55nqWWyBYjppT
G5oLSO6bayQZqnA3qwe8pNv58ozSGVt8eWKNVflRfcCzs/PzUa4mHyGyUyPZ0JzLSMKCffZN3Ez/
EVXH95A30SQfHleRoYQGd8W2C9Vlf5r7egIeXv/Qy2KXDU1vikg3M8V9UQ9fx8gLdRhKBsSJNJS3
YxfGSKlhTtAID9DT3kQouLgVde4TZ9y3ZySvNeooT1rsDmBfOO0BR8ZKaIDAnmUKM4VyzKN86hDD
YWFSURv3HwpzG2OgXZBQ3yLZo4Xh7cTTeYEj6XWf/iH2+O0uFhRgZLzWoHD09gPAYgrCKcUbV4CZ
jyfjuV6/Owu5alaLwrcTR3SLH1KcDoexy8T2rPL3fDIGUOvJfYvdtngC/Nr9ufqJBlZgU5IWvmm8
Q7XrTq6auKM/92OfYd8O4fRkPwL53g2sSlKTUMB6b+BqW0jb51fpGOerME3ZLIhkEXQggy9M6k5Y
7d3yNq9Jud710vDB8zJaiSTb8jUdFaCcQgEf7p1RCtToQfp9w07AW+xFNwjtRVxV7wB8vrxoK1FF
oMbUXU7/TLKYykJ8JRXVk/xrf+G3r/OwjEu0vLXWd03kFGH+UpJjl3LIoOP8UHoZs5Ew3liEWFuR
R/tOrKHVYp3QxcUJoSW0XxOSEza8Xr24SziW5C1tWohkVQc8WenRLy5YWft4gUsM0WjSUQ78rQJb
Swyj8So8F0tCgMMbDsLIDUu3BXQ9HeEreYJYVG6jPJRqWjVR5Apgr2CT6aI+YJJ399chzDVdoo+/
Sc/0JECNnEgpGgiSZn+0FBolT7Ayh95Bytv1i6OsCssQTDMdGLN6SdNAEEo67LiHNjh6gmUVcMU6
A6VWjNRs4USehnNxDuEV3xlMlO3V3BfW57LOj6+tFvIqI+SZ1pECykOfNL/LnNE2f2jF0/nQJYND
HSprxdi0wd8lmVWrrqCrW0F0b4htkfYI/aLFcCyVlrSU85MHJEvYwS+JYl6txXv4vi7OnAMz36FV
R5bym1dh9wfFw1UvhcX6dtdoGhDUMwL1nipMJ1RpepCdW7tE8tbtOVDDRX9QLanMowY6vrVqP2ZW
CPtJshNLq9H2msH90EVgPE7VDU1boKVZGwrfyUSCE0GSTT7v71CmOZgArkajpjl2svFwUS0MH1FD
FTxex7LXE1TNlr/qN4tvcqsh6GL/V4VZukcBcvrauMbQfJ+VmmbO55M0rZQmFw9kD8zWKaRZr7ES
Uz22xbDhDlI0R64Mkmb3PcpA4sIxTSIh9Nz5uJDupGGJBUxqw/oK/9Q+qzDkWn/1nCF80k8YPPJF
gB+PfaWzYM03Q+8RfCXYcTlqUNZaZptD3xe8XX4GuSDwguestsCK6DeQ4jM6tBOc7QrEcnRL4OZI
ttP8eJOw5JR46uLBEorvUsbh/zguVlGYBlqUrSeiHOwfBFv7cnPxAOO0viFeRZTrqCOFstkXSTix
mindMeu3yTZSo8WKu1zCRDU6OEe0D+gzUUbOcuY8cbeexyjH2e/DcNHejuzUb16IUfIybRm8EbJ3
+afXyYe3E9gzLAw+hsomC895ttgzNv6hz5hI+b+EQAMc4b4mQxZPdKeLcpKrY/1ZdRxUKNSbIJzV
+8rSLZo/pNawkbFFnMw3r1w7TArDneALvqFaCverFteKxgfCAVrHUkYju57gXDogqFw2BffkajdP
3y2K1rQisG/qjgYXSGJOQ16scfFTVkdy+OqPJq0yMlQ7AeRcqB6zkjNR1RnU6aLpF/pbIcFLjJlW
i0p8Lr228t9Y8o7iEZcbfUwHi9Hb86X9lIle7MKlbHRJcpXU7/HRYi4cYD84l6scui0h9iDUl9lp
cqChA3jRESxCSbkaJfXyHrQlbdKEGKOWK2ZmfHXRa58hdaPmWSr5dIr/1xUwzyHLtyIsUpZxDPhX
pBSdpypyelItNNbb6LOrDa8BfQja1SS4d3Zo2DZcSII0IPJEdmZvHotQtGrCqJeL4VZEAFMdZlSD
g0z+8qrpD0fMAAbH6gNdAbtyQojECuCPMq74KcVJh1I1mKRAsdb1hrLOaf/nq9zwotF3aPwbOXRa
fXEXTCluFLQLBeYktrSIRw+Qc5QXwk0Y3tOuxAddEoE4nRkDaZUZNspZTX8dxMxzZM7ISSrdzbrk
NQwzgCmv9K8ZNjhJrf5ih9CfmMXeWaRUdUWKoErggdMJ3mdCaGHEMuwSvlDUuwfNSH6cJiRZKa2J
PHwWQmW61qOSMMNcO4NZ296dX18o4OIHWv6+/VvtFBdUSC4dZ9WhJh6Nu5hRexdRKd7CU0/bzQmV
rt4Dkm2p5Oy33R/uFSTuHrMZsIbQveLgvObyXoa5IaQDdw2hJa91ppW+p7bjpPYh/oRBh6v0D9Nq
FBjLMmM8u85UfekEMtklGXCd4ENeTFrTKljjWhKoM5TcZwCflkf562CBK+te/EUeln4XAjB/0JQc
eYDn/eKsdE+yieiIQXeonoSoq2r8jgvuZWc8T38cqgW0MnXzPoSTqbBQs6sORwnuVrQ4xCuCY6lX
eUeH/c41xgeEFMLyNWyKfDip4pt5dhWl6pgKRJXtozT3qSqFbqzcNYJCmlLq2FDZErOb622KJ/hy
Y70cswmDWqICV4Oo8eENp2/9Gkca3e0BceNPUd8K0IjXEIK4k08O1WZZrRnt+FXIqzXor2z+MBkK
83/FjuekpZGY8AytE6damDUhZf/0n/B78nDUBzDy/yAf3MI9ctDxu0TXU3C6D3fMMQC6V0Ah6wjD
i3zssABPlVX73XK/VKqRZ8shIuASDUkQGApz8VoUGYyXqDOa5spH0CM7t4sG/3CpPJB1X8YlX2dC
Rz40/tzUo0nRCOsIAJLFkBvqAVGh6VfMByAAktH3Ar/uMPxJmvls1qs2YHFRnNPKFhdAfpDJO4Uy
JWGzUEflSSorVxnaWoK+L5Hg/TOVw2JNoCh7KZI5ttuNmmeCW+6r7KckKjPCl5EzMp2XbJdFmUWu
d84YwCkaxROeFwFDLQ4TGIeyXC5hc1C12rEHeCP86zP8eDDaRXNVf3ZeO69OC1CQTn23m25f9JFQ
J5+wSPWrQzsrHJdlttytG3Ky1l1ih2g7SdEk3sHp1IGaSIhZkdTBIyP5XT8YexoMsUcEuquevFeN
a4vdZ93PY2JuNUcomDNC+z3z43c3zzzKHwJOEavrmjCbCG1Zft60qWp6qPDA8x/vGrk7bG4uzd7X
Tcqz97nmndMTqHZcDTdrU4vb6v4JCU4PfxYUUCa1I1RUIuIoln6so3dEs1f/BQjg4SL8fJ/+26wd
9WTHm0BTTAMBUqCilyOxE0FYpWakf6ZLyCt6av0jBJ8+ORHlT77sKFTOAGcXkrMrv0597xvbdKI5
SPb8sBpUHLGgxIKaqKwjdnfqjZhEod8ReEAKW/4cbtNojQGpx0IjWx9fOJQLZGEesXOvSC5pPSgW
w5kZGDCWdOYtnkYUHdlRtAEjAqXNTlUmBT0qK04t4gLktwD024tmkzzuR8lvpTb4qTerpV+fddmz
PUvp3qkajgDXLhRNtb2vIofmKaRg+UKQ3Gf5bdISFAZ2YaeeU93v/ImAGorm75ALcf367/aRjO/j
pyXajjLskqY2HcQ//M8Xfg6XhzIJzHDyTs5El5wsQTAAych1VMS/dxNCuIXcHPzxxYQx81/ENWVK
6vvKU0AdRDQbZS+vZF4M/022BbGHlzaYvYwjk2wDJBz4kw0+y2kr17dT/fNWrBRFV1oFMc660a7f
ztMrFP6+kO42aSs9cQsXy7FnBwkK8CUOzUA/uBgmemF/VotVB7Songr5LUG1t3a+ZG18WWy7w0QW
p5QKqvir2xpe9QulpZvMOSpswf8H2X6UvdnUgP9MKBEL+WkVNmwByf3tssUqY1mlj/1N2LembGf3
h1VP8KaPUczZT83KZSQNA4JiVNzs/vKjBsQMrrg15LLvUKKWk6hnOQRdOYdWpfBrZAseJNIUb65Q
A/ZIWC/mjzS3HRytmPyElNybY6Fv6ApzYDWjUFH3H56gRDsa4HFwrx3nSeRQ6LM8FPXbgzXg1vC4
vWe7oBktmTcy66LpUh4mKeMCG569STjaKRACs45h/V32yw2AFPHd3X3fre2bT45/l+v4kttbvAwX
ctHt50UTfG33TL4ViI4tbtazfLBBYc87Xth9OHoKJb5scEyasROpSLTMhZbXyXzAlgfWxuiWO5p4
KCisUYukn/pZOWTEeyFPMdu8gz/N8r31leUn45X09D589az8CmxcfJFKnH/3JYQe5vu/ZUHithD6
3JPmjxAgZ3TiYKnUUxkZGs8rIQFwI+DE2z6ofsosORJYCE0pyxY+DpOgFpEqohOr1c/WWmpjAHh+
i/hOIuozDTe0KXh65wgMMsPRmErAlz37I3dzSv3bYxcSpl2jKTsSFiG4WywyTF5IwW9qNggjHvcl
VCrP2cibXhXu5Kkyo0SuAJ7fPyQpayKXOIiIFrY1yWJwqXl5P84gMQXl1eZCF2ax/ExnT+qnqNiD
BIAcqpzQA1e4L6IBHlDJnLVl0Unm8EhSKpEMDOvwbfm5jpz1JlecNRc1xf32UdjTz0rk3noyxSUn
b/O6IBfigw1B7G5jki5ERPvZ7DdV75K7MaRDrFdFxVOX0D+r7Qf/N2RX6xyoAel/bIAzcu8nLmE7
bRkW/4kpu2EhZWa+NFQvN4M6Vf9z8MEmQr5krTXHFkQDz1vfDGdHqGum0kcGggzyayP1n4IX/rqP
Ep+CEO4fhkPqii01YzQvMp3i9KkonpHDxI34cjppAh1U/Q/m0lkrh6fo4LhyWlprrNVFeCtWFQPb
HcruuHC9PAcSRxl5emQVm6aR/6UemdKDpvAt2umfVdwLPLJQj9WlLtRFF56mrjdN9xSd9433fuuq
QcFnOBs77lJxq4AhvJQlT8LGS4ZgFSOpfPJFXmkZ3HFB+tRWdWN5ucWGMPhk3qe8pfTAmNW4QVZ4
0OK4cm+cmDCoCnsbRue0fMcuZvELUqTL7S4Uch06za9khdSHxWQ80s5i6rV9yWzEnlEiy4O9NnY0
RiO7AN3WaWPVJ6e2n6UIT6vt0Ld80xUpqzz5kI3nBB2XE74PzNP/c0uGTHKDn8w9T9JVjwTQu8LG
Ee3cpUoOsO/kjQ8EId7hmrd0jxosVB+E2z95WnzegKRbbjSCFHUyTQRYsw5MoRgnVLB/KYDHV74k
P9a+YhiNEYP+BKOlPRYwGGWu0uBaY/rNhq8LD4CKYtLF0WzfOuXZXh1roYZRzBjpdkXxvTwU9Fd0
hGE0778K/adULeBX1fK/TB8X4wNntatGAX32hslo9kDzkmDfC7UVqM0/SWxUxJwQ3dgUM7tI7jeq
sghxCPq+tqMiIRAYE5vg1z6yNegezxDDMSe5MK85es3FJheUV4fRNRAk2wKGK6liQ46TOU5yTInM
FGV8BD4JofZIw/LOM2r8IGawRETuYs+BBppy39MbPsPgvaAsTiDSJL+m8FOBifjYXzBCgYOsRGud
jNixfGfvIPwkCoB+673xaBBQgbE4KQr+rPjKNVUWsMyRtiv+jmEQVMFaygAuDQLKbl9ulcWDAWjK
CH8kFTJt1CHxxvfbPl/FruE7sHNsdWvIQeblVnSEkJyFVVGfRuFojHgaiLFwSbuhTjyLcumqxSeg
W/zPdJZx1buDQqSIIeG0YSiQxIEgZ6XH51C1Y1YVQKxWnff+sQfNDa1Mt8CY081Vowotd8/A0yWk
Pwx0n9E/J/M2TnnzHfmpFLsYfa6jJkfG+XShNHEOi4q3lTKIqcSgoDhhPm6zSC9LfzXVwS9iMyiV
QTJCNbXFYYAZDxj6MvlG8wzIawTclJKYzfBH2mH1wHFVoQWtSlvGPj58GbBugL6euEgXS07ClzAn
JtLDdWNuPI12iJ0cdDNVt7eMZLcwpNdl12hT5aIfz0BR9XzA7OeGl5javEefP7zeHXg0M85jOsCY
RKMNVlQLmpWzvYcfj2zwqhycfZeFO40wDoBl5A0SbgZZja6aZ6H96rYQdolxbD0JjTTdfBPjy8qq
/vYm3UJYv2lj2PC3BKhQZ1Rm1jhsPdyiJZ8uoK8l5tW0c7/mHTwRU2yGdPWXTC4l9Z4Eo5WDYvRW
uuKbsWWHg3hFClglcOSJNwTRgr/19EuVLAkxEPxo3y5lyFFnA4dvruH2/iO66I+do/eb2D30Cea2
+fxhbD+0zvkTqWv8T13c4mjirLMktbP5T1kI/uzhoMi+CXuQOyVG1hmmKI1JV+dr1568PFvO1Mpb
pRPZSjVEXGAtDH12TW/PIVMBFWie3Mu4dOeggmRXDwuU/2EHIQToT5HgW1tDUHKWnF/6fuqZPY7G
nxBjw5lB9hg2xWUNUa/2tyty5dlnmuDH90JV+LDioPhVI61D1K8sP7wMYYUguEKdAT5g/Y7oV9H4
s1FWRnfskGvfHmjg2l5Oon5+7HfvzXSH8b4m9QOtL0YFv71W+9wlSReLYGMHOp8sYsFQdL5uPhFp
BDlcZCRuwuUgim7vp8ByFgosR0eu3Bg1nqwvDEUp8icYucQYGh1ca2/lh+a7sN+GCqJ67VrzX0Uw
dFnY0872XslS9tWBqa4IgkoJowNbGb/e+7eq4BXZxrO9tu3iQ3RX9CGd9tiqwma0hZEt2WsIBy82
FsuKQyAcJfLPk8g+gHb7JFjlky0xIbvl+M7BdJpfufmE0sQsB1ScH9XtnAge+k3uyTNrT8NxwEF8
7ITKe6L6jmZNwVqdJdWMCiGNxxQTUlc6c4eLAkupTlEqn7w8G45SGG/4ynLRbzTDQ1BWR9BLaj2z
9vECahGDiZoaKO4r7/FRTG2pkHIk0/4yXJI0kZ3Xxs8W+FmKqomr7EmiuNNgkMUTbClv3bk0nl5G
6z0+9ir1pCq/3KrX3VuKoEfPGhU02gq0HhBHBRU8eN8m2r9CVUphFLXP1aEZZsDCLqznvQqGPTQ9
XdjXbHcLEwWdX5HHK0QSGQYzjdo6kO26nOEsPoSfiLMRTZj/XXFVg4Ri/zrd5B1stud+aQNGEE++
GAxsUOuchwOH/kM9hREnTFZ0OpASyKJygiY/5uNgX6M1uD4/TcodlgKjXQkW6HkCu0eiDTqXlQjW
I+laAjY6exinXbwgqsv2oi9Rd9A/uB09JmBXyMRWQZFT5JjNe8SPgUgrZiOj2RdmVqV438ahCqdp
XjEaWOv427TyleQ1LzDFSxpTSwu90bMiInhj3LNqy+6JVjAHBJwDzpAK3MEGr952UV717RCv57BG
xPhVmuRQ/pptGvD5BE/sDafgMElTLWD54dCjrbw39XxTUfUcgPK916vveq6SauehMUmd3WSqSnF4
MYhRHNNZICZWD8QLpe2XubuRAMSPV07crG+wpJsBU21n3JuIXCuLhiL5m6fKlCsGak+a9pE3upIw
Zw2/Kf6yNoiPpLWCRozgOWg/i4uulQDQQktdBBUxhpBhJd3A0uSO/w0gpNgpL9A1IB1R5SiNf2Et
Pzy9ci1TsyYcNLA/0CljEYiuJzSuUUSaMHOH9ROzHb2ZUQJ55Y0hfODaOw9TAAhvveuCF5NmetFc
tFYkkayNvzUcHMVA2F3fPKnCMk7zLVuizRtX/47dP7cVF0vUmLSbIDGPqaKK0EJtK4QPlNuxvOQw
A7IZfdyMwg+k4FRSvUflVjewJ+osCUj158ZcqJwl1//EynEVX0qEixpfA6hwhpTkdUmJxV3riYGK
MDEX9z8J9dteaj9GSzIUQnC9+Y9mfilGjag5ccvKEhwBoGMAjponHw2NSEoPGbmHYsnAldBF1D79
JfJ0KWgimR52ketNFP1rPdxnQu35ekFU3NyhM6UFlE+4Wxzku8BR36xgyChSZMC8uLeUpSa0EXW8
48+E+wVdaOnr7YIt3Vgz/TI+xk0XXpKIfyjFxfsyNScUoPCEkqMAFhR9WXicWiMUBJa32uR5Uzqs
kqrHGZqSrWZv2wn9MTzl6Rb5LwRicRReUIxqlg2VACLhR4SORTEvOfLwflgQHnKPwy87e/tlIJGi
NTdakqh62Oh45xRBeqJ/9/1YVbx9JLNE5U0QiRPb4BT+/90Qk6nTIbLw0C2r6KftDv6ZXG6FlurN
DmkVE1Gg58SYTNoia/KmBfZUNZgc8xmQCQE+lOrDBcBSAaZCQ5iSIQDOJflT5GPX9Qq4bkeq3pSY
VtI3BVI241X/jTKM1iFIKCCZqeN1qXbOGsZBKC6270vdcmsnQ9CflXA/OKlX888p+xP9ouUIMqhN
tUuW1jt3ifhmhyFs2ZuUHDIo0MKt+Z+0/FRlwTXrOhMaElZPjLAGolX0KshBvTxm4friuvEi2gBk
avehB1SSUUfcCHHbhGaIFFAQWydJWrrvA65NDjmdV+3eHHtP7NGAgcTqZ9xMl3SIaHZAO8huZ+Ni
il6uQpVS2lxOkJcMBuwl5PhdUjZsDbD74Kqw9TP4upCNj2v68ga7YEU+qOfPqvG0PLfXteyqMa/N
SZ03XOTRiVBqEFIz/QCPKF/fBFRPHJV47wNA3apdWNreybAoRHj6i2bLjFyPIv9U/L9zmGPi0pZZ
SWSFe4toMKVmV4GZYBzFpCauiqnTHjg8R6T1z0rDNVkRAiymd5VGFODPe6DC30KkMrBA5PuLfF8a
RPNVz8x+nTkij5+uVGqSDnFYIvV/Kmbz6r/QB+LFvcWjLE3I7hHrdylxGaAUQzY+IdBSq/3P/EhL
++0y885oiqpel3GYy7d6fn6qGNoaYT3olx3aMX/aGJA8UkDzE/7/lqtSNLu07Byip1+1SW1mwhru
vKvp/liY5iNvY9BnkWBazJNptTJCNnKXxFe9KxbFrGwvHzaY0pfJRVdbqQ6dLVELanz9VsjyKPZP
xCCTtztvM4gj2rIm0qU1x12Z9pjt5sk5kv4Q/qZu8aYqCxX5I1cO3RP1+C8ZqskNHdyygTxzJHrP
uWKoJcokxXlT98m7SDTfIEcpYNQ39tjvzWdSOcug/PYwweBxBlVf+Y+qugoH08vO7iFZk+XsZh/D
KgHIaie5pJE2SUOfWS4yXYGxUwa+BvrcXq5fU207R8qiQm+SFm86HDXbH4RKJc75c38BpyY5pEKL
eamXOqsIs/rG7Pa4toRefEbk71gp/KFuQsK8quNl81zKG1rwc1QalYgigpfaolhZpWBFRG6hHtti
avgdu5REK1mTRoQpnlCX+C0Gp2s/DS+FO+EptGAqGxjFRVm/RRLYNqMcCSTMfVMZWHN9oI69KbZy
TnaILoejSP5ZaZkZdLWdlLPSA3KrfraF8AXCFYdMOgNbscH3v1dcvZ/TZlXc2tBxFxF3lhnTaoCl
g3siQ9/ILr3SlPNGV/t/E8vIidRivvscAoMvWzEx+lFeY2DET/VR/j9AOwVuLftvkciHU1stkIBQ
HKeE24REgA7MZyc/u+1Tx4LYoQIzDH1dcyTV+FD2ivPbL6zFPBVGRo28NGmh5VOTn+zsBgnCBO56
xAX/RVc3XZQh2WQxG3wAq+R/KBVgREiOT1kV8sCbJt6wCIZDHonCI0pR4ksnZ7ksffgClBCswCRc
dP1BJAgqkaXfAgGXW5yRYEsAzyAh9OmgJoO+90B/g5y+tYJSsERU4dhdLpJolz1kbGo/O3QSP5qI
YhQGaEMIOY/1yD8wRr0MZrVMUC8KbWxIoQ9Axfo4C84QWowJEUq/JoT/cEOdVO09qMDL/dFRS7d+
l02tyjJVfkN2RtNv9fSpdUzxXI8fzWgF8hN9xEmPpj/5iKpdl+4sYYBkmk0MP2c4RFjbEV1kCY8M
kEzZvNETdFPyD/K7xV/nudRvKblcpNue54wCGA02MxPo6/qE9fWUE6bxlJSxnZJ7ijW0Y/J/lB56
jgnBb0HsfyBo0XRTNtFLjuiRg3634qsZzkQTe0if2g1qNAHmoFtHq7WNEqjC5xgE9obyJsGf/Cdg
bxjoMGUSPPQLxobWNc1BM8a0djaEii8Qfd4A9We3frtjdj1KrX8Q/EN7EvyUeHu9u3i07Ud/kqxp
2pVgYun0n1Ye3qfWx7i9L7nUmtPduRADwV2sbqwvNZBQPmgKA+AAxFhfZvTencxMP/dgy+9AXzH8
QIytAdS2AIA2+yDq5H83+YOA9E/l6KcomxSQlLFmRGngOv1LCiPX58z0j0om0Nzw8S2CWL3orUSH
OyDpdQRRBcAD8iTwOpOwna2D+VpD6lo7I0QMp2laXG5Lo73iRYHElwmDM69R86N/kOTnju3FhNkV
PtsnJUBTvRIAbkEOw0zBV0GvvznSnkcHOQcm9T5cocBu5m+Q0OlpWseXq2ImEbA4Th41CZEf7lHg
MKv44ZX2xYzBCiMtqbtd7nr5Ua1Q2AjL4ol/QvWoeeLgiaDakclKZNh998T3ilfRH9+77Pg9nHM+
aU5wJ8wnMHNK+jS64aSYKIRl6+B2W2X7dRBoNGMRX2WAojMIESR3Vhqnqu3473zGK2OQDtLtrylD
bug4p5/pnRk1AqKNjR3e/ekkESGWeeCefcAS7h1Mh7V6+Nj0wWCJHMwhb86z2L99nyIPUfeqfieS
vMdGnB9DEAvU36rWOX63Aga7OCXUc8TqaR3cBOrUvP7HEtIx2PWpPnE3ENLo57ku0xxSuDEe4H2u
S1znD9EoBO67HQKqta9H+dOHDvJSyhHyyP6kGv60TQ4QM2026HJN4AK43Gl5AInyhsD9KS1vx+Kj
0xdPP4bNcormfZnqJeuEgjL7ngn4RdMs9jiOQeozwMmZmQNjzIcQNereBgMMEy1560S4cX6atdFX
iZN2ux68EvxyJ7Dx3xyyT9HecXfVYEBFFJUkm5VEo0UDYUyN3xHQGqOlKxXr+dQbFboG0TpB4V/t
eK2sx109iRvK3vggIYbang/jv+AoZ0O3OwpnbQMIRIHUuvn8fMEKARKshHB7SeNNIpRuXwcM071U
HdlhsKF5Vcg6IPsNAWcmBH/s4NwmQW1zjWfSx6atvx0uhy/niGjoqDaUeibArjulfghMG2STPvoJ
6sX3OFK8Pl65iuSM9Tw1QzCUp6NGQezlOaDFzMWlXsXYyqpLRjBMTZV9YeiWJ2iZSKIhZ/HYjQsi
dE4Jt2Lo49B5XwNQFTKm003GuKKa5HOkIToLaX4tKEBBE3ZWc6Fxqv8gWX9ZIPjOSq8hiXyNpLX+
t2wK14QzpfS+1xxcshGwQjGa831OJPjKg0UcKDbWBkafEl9FlWsFUsE75va9IkpFIaWm1ezpkDNT
XfCfTNdixUnVWrwO5rgWK0VqgEQxDwfrx/GtUPD1ZrdasNzWCrMiX9FMVel8TZV/P66bkDhEl/Pt
asCHYUALLNBc53kwG21Rut41tYm/agybEexFe1NxS/hURLVX6W/aac5OJlecQjstEu57DtL73R9l
HAItg3Ab0E/yefRaMx5ALJnc7oYVaVKFhGsIBp1w/0lq3bh2wIfOvGPwjbuQY0LZfCR5LiV6byix
ba7zA7rV8NpggmfGCP7ZY0Xcp4RJ5wDBsQHYJHTuDdubHDDoEBY6cULtKgRlsV5JNGE/PPNYvHtY
FUxWE3HZEdO+ZYIuSfz1944+k3b6nL03FIuezpDi4oIKoZi+I/hv5j3nnUrIyD2wKylvFYqnI91m
gY+K1j2xEm94R/9pNVatAXkOvNSo0/+5TvmMiLn6XxN+1OmoXZkN7mHHDH2g5qSAq6QX9Jf/oJAK
wyBl+aFWmTlcjl9/T0QQhniIoP5HoqzPdsTpcrszNCbuo8/kZDjgtrh5911P5NzNfDs9vDZoPF/+
yBrhO76EyEO6WrWNzGNHzHLoY28QzCQzGTo0xls7gi8HFaFhMBi7cxfzbHoS78r54IyExP7LtCAS
qiN3CDTlZ46vfHHSK1mzqydFt/J20ZqpoTBfP8qD6KhSEVokZ7xCWf6Adj/9iFszTbtqcCeGNrxF
PrFpuV1WbjU4XzHp9A7vXQuwty2XZ5/wRfTwZmM13FQKwtosQBi1eEGQKpXc8XB0+kX2TD+hOiYT
fPDqaSZ3R+/r65t+04jM5z3vnHuqWU8SqWyG57u+gilcLaktt02OuvtDQzqa5mjRMTjrVqv4y97F
/Q9WdmJ4ftbI+y+tXQqkZffchpP74aO1sxQh+m727fyslgrkLBKb2NZ2rKEY1snwzm6rsVqKF47m
qHLTIl8wpDmzM0kgHRG5y/VXVJ8WbIluJhy+I9u52aDoTmHkrPa3ilNjWfz4Rbo3ArJbV+WML9rc
Ba5ZoY8f8qJ0Mr3epyxj7aSlGpA8UNDJ5hHQ03NQRroJiE7rWm1Ll+UJl7zvwGZi5dLW0LVWdJiD
dqLAvsOQ57TCbdA6tn9dSSlwm5KKtg915ZJp9VZgU5J8TAZai0rZ3U1pl8Lv6DLTXreK5K6/X02c
rD8UnJn3W3gfdGWWr5H66iQIlRX62XSFFEE7gBrYfuLz0p+vkOcc8hn8Xx6SO+aJkfKuP+tnt5QT
+SB9WvNQRy8Fp4hTGFmAsOV7obyiMbzYMH2Mm/32379cNRsFI1lf2Zq5EX26yPV43AAE/iXDvv8u
9191qwKoGhfED5xtR83VdXPOfjRdGF/S6j8jjmcHvuMKRk+bzDmaab0qZR0lSUAs4DeUDPIVPaOc
bf840TfTmx9/5TSOsh8CpNZTC4rcQSGUb4zaDXCxnWreg3YX8rUS+WE1tsnOybNtHwSGCj5aKcoB
YHas27TDocGi/XIPfQ0QKB8syJBVj+giXV277NgmqXTHcXLoO+eEKh4tgPqLWD/+OANLmI29o5aa
ulg/9h9yYB15LmIjh8WQcs8cNNCxWbcg0CHbzSea9Uo5HT0EyqRedEJp6dRqITCshQQ/8QEIYCFM
uwdCKPOG8NxO4IoYCA9ReQqQQNd7WDb1qfyuP2MRFxcRt2PTmT75hYYqsJZUGXuiMEhXa6sDblhK
f12GH/I+wVBTM2qs+ymLx/Y3C7aGIQk1ULf1mUBsAjApT5G34zd2d9FW1CfTTvNpso/izGKVSKOq
1fObtcluMhuMgaAixF7wQiTMBRKwtG7ukb0KSkIA/VNa+As/CSzE2m4ntmyxkhI/8rUH8RWoYhJa
/i7KoJfMeDbjBsdSq/87xYVJzBX5/xlveKO3MV4BFT253QBi2GCsCFtEhODybGBoCprTtxHfhxSP
brmqLF4V8h0CwCkIFgCu8nZatPBvMi4fGja/FPKJ+ZGkZ8O6Qhen74znJPvhwWQyQd2obNxm+CsL
PqbEQiRcjJmwDHYWr/3rUlR3uppSXp8GQ1FN0vEHhVHpa8XQL6NMUH2Fspfny1HNRcnGwgNiGm16
jwd3ciP/xCKNDkbTN/kK2AKnwsrdGzvgVnrJuDgVEokMvH7pbu02MyFWRohT8rpYydECWiLK0url
YWJaI536Hd7dCH8yF8JWoWqx47Mv5x8F3e9Ig/lBn3ZeaTjUrZ/ed2+OYQdvXhcSNEFVK4Uo/3TW
Ggx+HnAmKsEdmt0NNcF/Kg8kvcYYz/k8niR6S85Co8xSVewh6ks2wCDGmdQ0ssaoJqRNM3Ku7B0F
ngjV3uvUkAxXwd1YdIvdKfMPl5xLdmAfqQKyyg2MmBvPjDZMfynUpXq8SvJr67ZbECPe3EBGTxXZ
nxQIgKW4f/YArat9MsV4TbrBh3mfzI6xh3dZivXb/Xd3luLlXoq6GS+4vnQ+lev5fuL9UCawSzfX
2aOqIXU9MiX8Roh/bKbVSMnK2dO851LUcZEd57NbVvtOzEea9pdDTHJoGwAlIgEvgwNm2q8MYei7
hYW/Vg0iChb08wye6OIafbevwV5GcA4lNWIzYAsZZzw7RVrmwiB4BTZuhz/IjgUMs6h4vXYU8rI+
73MOQWJcMM4t2Dufu3d2dUY8mvlF6asv1Tq+IXzUMS0PE4KbtexEY+4j4o5SCtzqzDsWsK2oQRsm
+nleImhhEAsjm6EyvGooOF52ouGCX/OVUAmnjETLjzxkXHuf2Oo+xvWJqUz28ytE2kzV5fyKC6S6
A6llIwbxSMJC3Oq7nOKMUsiyxisI7JIxY+l8AA3fAVVJJC7/+TSsaSIbehOdrdZRDrVcUCp90v2z
mHnKMAh37Gl3FyIkhlGuUHKYH4/Ou7fvwqb4bmai6ijINg+xGAuGfc97QjVDCDcGu0ftOsC8L3Ax
PtM9jap2G4qCfPN2KjH4VEYbRPlnmqW/Ab086a6pAhj2a8kCKum18hKHzQNiJfsPPF18xwld8+jw
lDV48jaYfqaAnuqS7BSX+66gCEvfYo4+kVcjhUP+vDEV8jPdR7hoKIR/+wkzCpSWaKndKasAMuBH
HWXZ6qxP8aLLYzoFhUs+XrPmcJ/xT7auufgInIeHdVWFCQyaK/ngKXAGaEefanJzflIzikOUHG5b
/0Fh6jjdMLpJ4wno1yYm0x4LSoMIvUgLkupCal73Nnx0LSFcW+vFU3gLVBHlC6FRfJopJNyThmcw
UB1q64r1dWGbNveKJmkPtOd/JUCiHBIJC+856O9+mxFV3hYXcT9vn71AJ8fG4KASrVo6gqmCFd0/
8ipnS++Tg9GgP0P2ZMYGbZ8/qlaLw97j+gnY559sWm9f+ui0+JoDtqWU1lXAZ7Ua5DX5nU7lFnDd
YkSLgSkbi+C7w4kebtRh5VT6Bt4r2K1TZ2GCxOhaof8DINIFOEgap5TwW/ak4z4IiCdJ4AMfHCNz
YwUXxQ6waV5P9+QL+0OIbfhh/7CC0xf/CXyJ+jM21QenKXK0Xv5KNe62naQ+PVjcOk2B0qUY7t/+
6baoQmAx7ajpk7XPrm3wEUg4Zmkp1Bk8w4UjBNwvxBjHM2Rgk8qGDANNtKIzvUyidXpdmoLofPh0
NeIflzY5kQxTNpegBitJAfnn2bl7hc5H8BOfOQO1dzedxnTjcO6q7opIW2NqIaVDhm0O6QdWjHEY
v7sqkvruXONklFBmHPDePPKwz0UxNEbmDasseP1vZSdEmPBf4zHohNGyxxzEombTDd5poFYtcBrl
tnvF5ss7Cd0F9eXrozOKAXIpteKse9JJcGFnwt30+e/2+NaMi/PZTV1343ZHJwpYtSPhJK7wyUG+
teVMx9RwIiRCBFtohISz1HxgJw9wStJiJ/fbWApHLrZeA53ktO7BfWLqRFRHtyT/g2a4iaIWxmBF
Vo5m204799pnGtVotug/F/pUFv5tVJXWG9d6ldB+mViVTfd4qA/A4Z+JBI85LVoIw0Opvr3X4459
x6r7dJs4McsT+qt0Q2oI9/UDJ5A0PJ8GSJ2SALjkV+wycmrcDVIjXq9N8fB8mKuUZGbxUndUTsS8
5yJ5fTmKd3znKrDokLQgAJFHdvaepxP1B2jh90PAueWlwmVPDqXME1TxKO9nGIhukg6lsmTlTk1q
9SdYCny1FJj7WS/qeGhThQa6ffWm2eOaZoOxzxmVo2RrlvXUVTS5s/AsCEiRsK8kIXxwNx6mc9Qz
Qwi2iqj2LjJTNZH8qJV3FNFqEixjTCiB1YwlM9UTqf2LUP8m4w1TJkoCoa4WvOSCtUjU4UBA8z1k
8A8exzow+D+PV5hy6nGv5EQPtH/iM5TLXRAS6F1ODkgVnCqBpTzOTCVfU4U7luQWgls8gY25UfXn
aHU6K48UXCkfAcQvT1ca8ubv/MlR1CDdlrgFUW7/hmneQXA3yLc3oJl51yZ96lwlQaTbCnNKn9mk
1P3v5iQ2i07AlzXI1014QaBd/0Odee3r8He07KGPIoEQSofDEaVs3xfsI2bgAIXueHhWybeA5hWs
MavSGC0pGY2cpnPTEQnKEOWuuUM5S57UrHmx1sJjquhxBlVbxXO0bYBhISHQJ1a3gK66Hsf5lDYo
Ng5h2/H8S9tPqdjsdNyY9z0S9pnqDyNtMRKpNvmLJuvMKe7vSKfa3XVM+qF4IaxdP5GTzw1AiUo1
qseq+2H4rEcg0mOOxYTWDsTQe2G2l5Muzui4NhDKB8ftBRr+92jYXehqXcl6JHtBba51RD9xeal+
TwnCJlsPJR85WMqiDyJ3pakSuF2BLT6aPUD8XHYDSo5m1s3o4nbsgC45k6p+ES0gwQhhifoI4XTP
lQT4wgNDyL0lKLTR++y/SEnzBkgajkQmjQtDPQ8iL6XdalFiM5/uOKpBBPSVq7rXJ+sefoyGXjaQ
mM1uUzVsSnS1WTKORYYKazOTrjgDrQGqaSJn+69RgE537esPBvrQPwoqv8YXQqOUv0mwNOCMleEP
3SVbxc6uD+doh3FJ5Pyn9HkmncdTG83lxm4gyR8gRw8JfCpPUQ3HA7QuRqUG8G6kWPXkGuNeKB8F
9n2IOVfIQiOWdUzP6YmWemDyWI3BkfOKaOAwF4MurgQLYnEFaoUYTVzlSXS27vmbyv1hSg4pq2i/
OyFfcSChrNE4Ol+wRqX3MAOs7UZ+v1KLXY8zJ2gu1kMIr+wFo6iGXdxlvOfpgCcHMq4zmm/P+Hfv
nk22ziVr643dThiZQzAB1Jy2E1j6YA2qs+4LtiUswsHtY9NPECeEftfuhnJJm/160dJ3gFIHKWNw
9teC4+hpnSmvOG+rI11iIyRqnvVyBEpoaw7u4AaRFXfdUXlFEnLTBKTMUA1WZSTy6IcQNpbS+t3V
mCf0SLyVbM00/XQE027574IlDP5XhjeVvMlq093TgV5oEgYjZwINGcZtYTxun4z4yKpxz18WPEkP
y05+OWHBfscj579YFPsB15Q5VnlecCCtZ0v3SMrf9aQALvjmtZv49PJJoG4jZsenLMWTJYkEt3Y/
lA8FoG6jeNlbi7YVyMu0aSTb9uGGvtO1i4ZctXIWBbuhnS8wqWMKCxyjntUD7bdXQ41vM4t8qzXI
mzIrmpfJU76aiPsNfKgJlXSq5gCePy+uX8N12Zuiok1007vVMOjQo+ANL25vjo7LBmVs8+j0sdAN
6MeqpP61AKMwW8/td5MQRBESXojQ7cT26+66BZp7fMBpxoKQAW00qtdSas9QdqWKssnDz8rXRE0w
ItyVgFev1BmWyeaKvVaq7Lwjr2zf3i+fubi4qDfa/vKmVl3KVCqyv/8JBPvyo6+sI+kHR9prj6lx
M9/MON6xUGQeRi6qU3vnrc3RBs5HRTUvoncOU3EX7Lnd9rHPX+0yDol3+SxGW4jQZ6hUS7pektqU
ynIZB4DSv9uD3hCRqZUmxX3I+yiTyNLoelm9xxE0a+zvrL3umoOx7w6wnmE75n1eCi1nPAxEvxsc
jiuzvHcjANGpUteINceBcGaSflPU5nZm/6jA60G9qd21etk74WyRTPHb7kLNsEdVlVD2VdegWT9r
UX4AfzYBt/odTP4pdJjsV9l7CpAcbBlytO4BNmzaJZMgKQvA+NfYMA00U/1InrprUxYsLLvvHmmx
bDym9oridZiM/kMXccTyPI4WaokbznSsGMh7MhwVyNkyI4GgaEQX2I1uuf6tWzOng0+RB1RB0FBb
MJtdKdmCIAqw5ht4bjU6v2heUfjEnzvmKEnXPZNtovjYA6i3tUbRQVy+y2rAW7x2y6HpGAb3/Y7g
eYo+Ruc9TRP+Fvm37ZWQpvfnYDaEoXEkFxdi6Ren4/Q6jYT/HzzOlRBE9IA1KDv5LN0ZnNx2sguM
h2K8vR1T5MvhKBYAniTQd/e/j7gGI0+9A2acpvQWKoe10+5EvFgT5cd7Ht1SCMdXFwgjZmFWls3Y
IoymieXqUAibq9K+rPFi7zbvpqHsozrjO8BLNYsEptcRGoU4rSnHjyBsNfvea5UR9Uc3TvqyolLX
cyWXaOPvhP9k8WESZ/5Da0aZW+dQGOieh6php0t/7Jhi3TulyjKQShSoFGv3ymPjnxV0wgidjcE/
jbBhi6HZgXzyGO9whQHJSYOo0tU00CYkv+jo8UxV2DfGxh4XbVICp3sU+rYddtt4V65uFBihCXnV
MBjlZzob8czJDbtAGxxjrqx6PDZ5JYYDMbhFn5zPX1VZu0Nv469fA1LTTKUSs8aTg0pOxzgAh8rq
O50lyYCia+1wqxRC+MvlZpzPrss7tiTJ+kXPde5uUBSU46VSWi2KefT0xC3jbpcDqwc402MwGwEY
g9MhzrTcZUj2/quyJWmKqMRKXfByQTnb4gAR6cTjuFmXlD5gv/lGEfZM0hKEIK7vlHO37sJfQ+1/
dpG7m+FkpCY2a6rfU6P+TOS3pAXpbDi3tPatXcvbDxo3b5ImwhfZoOlEnyHOHgYqgCpXQScTrnre
Xphi8fMI3zu1bvylFgj75stMJHTfXM6uIAi7vvu8LSuWqpBZd0yHugCQBn7tsrWkZ0RDxMwYLuEQ
eRm1VbyIPlGRVDrPE02oD+6BtbyLKhMYHzhLIMrVIvuD1Kz2rkFHUqWt+chbHvsFyJkAFDW2/Kf/
+Lh4ZiISpO1OIHntn83Via888/u9rq5lRdIanK+DLqnowBagYszX0qOchghLB9r+kq1XE8yGc33C
OACQoSdKYkbMyjBoft5RamV9M5sgrZxPhXRUKeMeq3o+iI/puQN1Sbe5UoxOjE9KViZlFqVr0IMj
ZmaPubw4N/kN3cgKjw/ehv9tmO8Gf6rl5sCdfPktnF4uxncSjO1n2TEhNbL9Ph2N5cuZok0LoOL4
GqNGiGZYzexKM8Bo3fIVq9L52stzQFr/JUuCv7TPCksJt07akNAx8du9bUy3j5ScXRsPOazMjlwU
1mX8jjJyC1MdFOH+BH6MWZvz8UVOSjOBuxjoOn5FKkAWhpL2Csz/qfAt8G/uwTVCp20sJLHP0rDv
rzbudfvCGAik2rKhACNaOp/1nYGFFHgYLicr2esYE5QhO/ZNP8S5sXr8F1bv5BaX9dx5vUEjSqBi
4sUNergGRx8Huvm424Bo0FZ5z0aUTdqZoBmSgXmZtWcRLaJej+O5HJrLICU34q7kwXIzXIBRfv13
476sGI59txMQhxwg50hYrqv4IqCTBFOv734Xd4Aafm2pD0Vks48vb7X0qf5fNLC1g3U7ViOICqH/
yI48evB7iquzcryQBZsQjS0yLK12rlERi51GVxGfqx4lD592T04E6/dTA9Hhpk85b5/TV4J4IR4E
eYw7ky4S47TNL8QxilA/vgPRonzsqdj06+HFKurAIZYnef2v1M27QXj1fTOLuUaTis+zMRrDwI9N
tfxT8kb6mnT63JsUm3y5ibpyRsBaZx6+wClDTClN9Ma9Uczy1+Vifb/DP1m0C2KzMBoQHe1Bsx5b
ledVLph7KegJjQfdyECqKkCdyHQxBBirAKAR4h79zFrHJQOg04C3gWH1ZYb9LVmIdA651A4h6NVo
BkHQfYkcSwtvxvk1RXUbLr2kkTp7vFListxoUcxBzw9T82vqRDwRts4DhDgDZBUEIN7Cu46nJGNF
AtCL9vXME5Zn/taJsVAdR1x3mQVxnOwxD5BarlVMcy5pXaKQQTv2JHeHYPjjBTiwla748FEgiEyQ
K9X3NPck9hQTcCeoBgYDWqEB7ECBGCUFMWk9Ux6W7pqF+lQ6H9LLFJKGVN+17PQj7ZngICYsZvLC
0eq0a4EU1ZDghDTnGfm13JUQSMJ1hEn8TjzoR88N0+SwvdhQSstnQGie0dD8ikGmFi1fdaf3OyDZ
QJkKT/+Z7nHn1VpPrCnA5J/21nyL2jSHoNEq8gFzea0wY8jbKqAn0iualMPRYYtV5LR18gnsPn0c
nz1Yhm2oqFfEbdQre8yDadUpzl/eFZS1e2XDG4R+TtjwnTu6z+3ZazEXtzpeC2D6SdLf+GDBiYjY
Nm0n5YJkq5DlUW7ioL6//NtGtFRSECrZyo+Pxchd+eLwXs2Zog0VQGpD8yE87VvsNy4mQXjzkwaN
/3Ri4o3x+eCW9JT0ZRoopq6KBogrW+WfO6vJwjG4G6cGbJIrZA+6VmzNxyobR6EtLQZZ4sfyAZ3i
JWdzzlvMnB/GBFIMELNFwiYEKj06XAfh5JaosC6VtzI9TtXowQDIhmd/2NXRNcknTNNAGn1wpmpI
mIlmlof1W+siuF2qz1hewf9FAbqPM3X9b+dQZRF/kwHxuvrXzCKJyInOw8IjKmcNtoHa+orGUhT5
wwWpOBG3C3S+Rx6V55E2uXWstpoecmWflYE/tJOHCstHqQ08TQBAgCAh/xzJ4Tunkhgm7VN8yQJV
VhzHJz6+P73Ke4maD179kN3FkIE2W77Lpb4a4jycdU+vX7OiwuBG58aTrEKOdSzg8lRiwSrHuH1/
mKaWPEW4CuU0V5Ji9mQfyutt0HvLIEzYxc/GlFWaSKpLBr5B3Ub9nYEoo6RfYsIAL2igmXSaJP6Z
1QSuicD9HDHIogxDCdJLG1RFprBtViaXAn60mvqDQfykEYsteYjLN0UXvOUVXTeqZ7a/K4PKYu11
/aIwlendOzVd/vdvaj2pL4PCki0iq1eoSdgiPKGANMDPraS4UvxFobJLk6qPw2aSyxI0owZpOTVS
164GUcTNDSY830jQDg3rIEPBAk54saWASmDucYzRGXlPQX09Q/tU+0Z01dKdxHzC7hGU6A4tidNX
im01IjZnIdTmHacIFCZQyMlRcqsEFLe5P99T5inOGGNNeFZM8JqhyEvtm3l1aDUK1WVkq9+epf2W
RpMAnA6NL1rv/XuuKc7Kx94py1PwHWo7U3QOHm3DZtnFl47txMvkn3eymxfXfy6IHpdmJCH2ZgNL
n97XOg9SivLN2E8L3S/U54ZkXy8hoCLsTbepzoNj1PxnRiSTPWIvm2PwvKYZ6xsUUGkTqwrSbSBm
bsFG64OLyKsMRWj6JyC/W+UMvJaSivqwAHamSfbZ1c2CE8ytgAA1KH9/nhNfom9NV0AgWNErMmlA
8FJkMIC5oO1fJxEBrYUV43qLbIVTlBqC8HO93FwvbEhutRFDHSErqX4Ky4pByCElemMlaaASCEgD
zUqeZdGbvMzZCwX22vyZIGxQnT6WmmZNVR2DVDjpZrlx5LQIrsqAR74t6lXOTBT0ksEMirmSL7Sv
7kVgUQgV/jjMZJBOAjWWoeKe36Lsxl9PavWl+nGZy2jlL7+MFxrrqRJyOr3psX8d3mva0VAHXIyX
9U9Zu4t8pDDesD8q6uHO9A4ojbAnDqNoQy2CY8vblBBMeqGe3jsyopLhHqNZ3fkBHqfKxIDx51PS
iS4CWc91O9WggCSSct4kTgr1eU56gVTNsGfE0ebou6lCgWK+1IK/T0jwrvvwMoEoyeL80QMelH7o
8DKurnyliMpzSzXdzkyBUwOJuHHa9J1aeoN/lmNVxWeZbOm8KMtvJr4viDd9PHvK9+2+fA535xW+
1h1edLvnEG63F7V5Elp4joP7fxbtWddFz8pR7emjf3gPDG4AI4XX87Z5Fz9uQEN+SZEj2plevEcG
aFW2gWzfLGr/gRWPEFV0q9czi6+2je72au+fD68gVdcom1/0wUy8eNe1ws9GdWv+5bp/HZxJ9JoS
FEix6fVu8s9Ogr5x+FRvSX1dWKVysAg5egiupmh4NZFWp6ut7VW+XE8vWTq7hSs+HTdWjn3WDdB8
bdVlvH2xVSQD6t+0/GqcN9bR3D1yhcDfT9wboTS04wCa7K3/7v5JmnvuLW4230tc2D/6u8T0Ynju
jNScaMQyNn+4sDhHA3NQdluhTJTk3U80iVina6QGxs6JwSkeV2Gcy8WD7mUEeYR9tW8QtLoqeOSS
uR2gBBHzAEbWxCUKtBmU6ZT3d3o3AAJajT0nIu2r6XHfKygVOos2v+4UeLYgDPR2VZOTpGEasMkb
PshpGfR3RqATAfXAg+QS8vhegDrbR6GvyDBHmAhkjD64zpjHIDFJRIXG23eM0Nh2hfnnbUEHwn2H
C3XuNwzH6DudBT5FL5F5tEo4Fq215tYke0XDasIGzmlrNEGRTssNX6GEwYPYmT6QzU6LKowhyHae
zn3NHu5acTBE0Tip+vnTq68sXktZSwHDHtkHQx4zSUrilXqG0N11kzAz0ky4GpcgUiSXjXQE363C
hXgOdkxIU/nuIohRVFsgYLOVSLrWZE3OGLJXk5k7qUV0owtDuvj2u0Bnt4pgl4KeV9lc4QxXZaW1
qRnC7IP05uuSt4U/bEiEKSQaTaqNRPUnfPx5uxQ9jYWDms6ioG7Vb6iR47NZgbTuMHjp2C4ztwh8
4d+Ja51ZnJp+56umiYGyHi1N1DojbAJq5qXEtamPhngRdiprVRJnMhi0pN+Y6BOIvrxIxuJzKw9R
55sNMZDd8recH3SJ7jEA1HhASSfu/9Y2X4fsDuyWq6JMd0GdqA5slsnHd8abkPToQvN9/xi7cn+1
M5fuxTth6t0eVSbWjfCEZ9imPB5VuWQq+6mSz5mrsAp1kmEZMWAdFZZyoUFfn1tHYE02rr8vtJuU
UzwQWJNK5SKstU2W6bkrb3yL9D2YXmltBupRfOwG+MnNzNi1xMtPoQDG/ka2URHX1cS/Q2sgz1nm
GF6yAf8eGEvp0kbmycnumDMGR8thf9O/EekWa/EowEscA1kM6UBqODVZo6m8Nr0PYT73XrEU35x1
A4u4qxg4wl6U1ZrCXwn9J0fl9YLi/0ESJ5QGnqDjE4cOQ48vE9UbBxVUqlo0M86I3hrzPMwlR+Ps
qSxqnvX/iEITVaM6LRP/sbTjQXLxnn1u04DQSjDd9VkMwQSc5c0iQwRFIqoxk8QzsdwO73pzhEvz
L70vSIKFakusMQqT1ZoKwDBbfFPQz/JOONaMr9sOUDa9mIMHz4vLGA55UzRPzKBwQu26c/2C08Vm
ZDdPFXfyyBgF6VMulm3HYEVtKQAwaW5epKXOYSuuPLsRoOzvpbDKdzERqgKNVF561c+w4priEsBg
j0B4KkHb7Gwc2Y3mjLj5PITGQsbYPUI7P3wFChUHaJb9AccealQDc7n1k6Wl3/EfMMg3BBfw0lo7
mzWJT7U78vad100U/fqM4DMsy+EpOhLoLoex2vz59oft5qIHWsbnXdjKfPx/pcGnfk8qixOZoTL2
474ntzKjsz0DLgJQLPTv998SUqC4r8tYE/j8NKUDscqO21r9XptRqa6JZZxqU9CMUiRuJpq6t7VY
HEx/Lw3vkeiWNCkOEl04u8Pe8eK4bnJUrZpnSAbL87aFiYl0GlilZOke9INqWQFwlWQY17Df1kG1
5/EeC/wNUIPG6Q2avWzpTpOqYhv0aSnU5WNd7Y20YoUW+SEhgyWt2QFNf2u5zOj9M3HfaM1JZY5l
uHmpPs6EV9Bn3KVZs0ODjrD0y7xvpPM/NaCn1HYtKU46HoJtq3TVS+krVlwgzxg9rPPRI7Ug+5f0
0YQzeOFOkG/SithFmk5HSd1iGW7NQPaAuSOdFEQHGGFnkBmSgr2mU/00p65HoYhRXSSXT3skNBHt
cvzDUw4MaAeSSBvqXfqlAslhEHoMO3ghM4oxhbuTs02Ax41Zkdp83C6vKR+URw10u1b6e7BBh8iP
eGocfvnO0UzFzN26Q+53bqL6k7Cwas0dRKkvmwlMh+GC9Fg+TjGjCwQhAoQAlgoV4wW+tJOm46lL
UIKpfWsGSYC/qwC2rMeYDpla073h7pjbAh/iYvBK2wp3Uof/ewy9vtSQ7OfI4lr8DsY/cprhJMlb
QmV0jbxo3iYg5iokvGOtQaD3u/3+xVu9aL2CsYBr6w4oqUwij9qHbPLKZkjdOVDpV/Hv/izeIDoT
VxbT24vNi98UL/oyGRpfuzkx4Y6Px1u3LMjGzcPcP4j8av2mENwqsEW3mApXZnWECGWAlsvciJNw
mlMCrrRy+e0dQU3flcjxYFTZGadB6HnEiT1HbbD2aXhZIeEJsSA/m+OetyRzXYXyOe1WIPBBRwCM
uHXBM8k7XsiLe1JKaKsDAICQHeb4F9wP+V7Fr5RzmjprxFDeulV4F3xVVFU4GKQ/Pm8RsunacLBG
u+rEwqQnLNe4G5gBqdciHNLf0mlTDfAw0kqYbQ+p0HUcNAgoIguOX9NQpLy+NRdDo95eBV7T0qcG
pya7EXlE/rytDlhw5ZoY23YJntqwLI3Py/viaNL1nBbgp1sOUCR16e6vtz9tllC0rSqbN1KqGkRJ
hvBjtRcW6gcTqqnWf9M8jE8Gjpjx6DzJNGM95/HjCE17xJ4OrGl8xk/eSiHsyX6h+0UT5bAiuZ+Z
WgfDh1o081Wpg2qNPf/iefO0r0pcXq3oM0SWrXy+KVRgDNii1YfCJWIOHhI5tvwWTGMAYKew8kz7
vKe544i0piabqblPG+gK5hDpbCGvDXKMXd2gyLiF46UCmrm0LPGrXrJKkBHOitjL7VpVma2cvDKs
412X2FCYw6oY2eTo5lOzXiMbzV+vZDmbW6DC6nO9i2epUkH+lFGEpht5KQfJ2XD1SyU2BoxdYjkf
f41d2voqe/5tw0qEiXx8iMtHOnoijPCJBQ0PVfqzrBs5NTK7zeLO5O38TrY5Ja2clAEHfw76gU5s
sSe9QmtoSBb/QhX7xxBVgongirMPrGMiMHn/JSTnkQDgw7lQbB6XAjdCex1dHX0dxQLCJA3EuHF1
uy5tdyMuq3gwlS6uH6Rc6l9IS0UaKjz+HxXOeZjZ4Nmd3ZYxp+hxepusc3fJ1aK7GtJ7cAmQb3kK
xol/xLfiVe3PJBeylwVUFvRkekcuSW2588Wvp88vbjoNyWSlxwgGIUAsnFvuop4sLpfpX59ZBgNf
HDRyF+HqlIDA0EeeqyFKZ/BL6cfsQdIXtXLTq7etApNwD/bzFsHNAiEEetbnMQ1Oqi1UkpPOGVbP
ngQhCsZLgZaVAZnpuu2W/TSSWqgsTz+9gc5xyYTRrbM14p6zpu8AlbaPsfx0E39+j28i1q5apdO1
t+8outIeWSceKlWaJkXVEopV+8n8EFYiqpTiHtfJO/e/U8XCmHfKkabWRh6Hd4EG67iNyO8f6+uH
64ZPemo8IE5tjiRXxSXpDSYJjK+aNKomVusWPZYYmimHzlUVrZ9o7qPeDlIotE2XbZNxltPQGSRw
IQSHzxy6vtLDwUp0zJsApJ3KLoDzRpte8LYVKH8uwLXEsEi5jhrR3Ircz0HHJgjOPg9bJrhGgJEX
4b181ij4hAp1mpmHyZmVnrP0s0sk/Je7US1qZ0XQElphlG+xaJqEzikjFR96Pxf1QJsAxdIW67Ht
FjIgERLK0qOC+ERDTpvHK9VUeZ1fmIFNMJTGsOCOxiyEmyLB9eRDOYfnluLTTQ60hziVEAOTMUZx
mvhk1wwyWK+TCKYJK5kukQJ25mbQAIOgaKrJEZOaBemWawcj5mgTEy/QCOjbAjlqMendMEprZUst
SdK/qKEaq5eXX1vPGxeX6osNK9OPAPv8XlsvZumCp3t7itWYy1PcjIHV5ReG2pBRsj/FC9NBKjwm
9vrfB0zUr9G9H2vL9vh7GgrkxHo23yJe1rfSd61eTu/uIoS1qQl+AsOJPXhaBUGgPZIfpW+x+kNv
6PCFQGEPi63PGdqitdsTipO2ZV7tOesmsXqPrJeTV4AG8ei8h7KsXEAMHSiZV/RESs3Iv6ZnxQ3A
xSAEVCmbpcMCSVZXa9BsL+bi6BsmzZ3E+5kPo35Di7WGktsFv9JcZFPgRXTHZJEjMgjTMZtczz6g
p5lEHCbj1gbLZ32lu36Xvf6aDsze2NRsrR8lypQgghms7S1sNLfrFwIuzYsP69ayoI9aF+E8/kuV
Ly5sDVbhT0UVDvWSJ0YyG9G9U1vPsK3u/REpX+av9D/v8MWI7E92G9S2/W3smwurTzlKYaujCuMq
G8H5QMyjdfoy9h8vN5U5RicqoRn3Oug1X+jkNMcY9+nYDzs/H4L3+GJ0pYrmWCYCUaqFcVo00zRr
jkdz2vhCOQLT5NtKRk+l7LuMX7Q+A2XZnNWSDMYldPeTWliDfjIrUiVA+iC2AzJuIkCgAJwavKoW
g0/YYVHBbJ1N5kut9NCtXArpo68pdviUA6JAB8T8jgqp51KNatvgrIrJF1g0kC2tXWeBZv2whfAM
MRlEMOOL2Z072fsV970TEbIXUUxNKpvzytHZiMiBeBN3QN1K9q7odToG0GgSbVMuOwZZi/SQrZ8D
yprotWl9ttL3xF4kefqgtDr9npmqYG4aTz2Xun7gzVQsCXuhSCAmuswmek/+eW7lfJetkbx48/wv
I6SiQ73xaODG4A0TaQScqHbQpg1S0XKphsOILzn3/Sc/lto0gEoobl4FdcoTc/hx9xXAamBUUW6R
JLWB2K25rHYwY0OIfeHau7jYZ+Y01/sXFu+HK2jwhp9B0uV9cKFDQZTXHoXlUHkh6ppPHiM1IajV
92VSSr1CSPyZYNRFGu0jX2Q5UXcSBniEdbmRkhUPEAqJ5474xAYBmpEDHSTvioESE1PPZRJBULgi
a5+gwEiC6w24pgEzQw5/LQ1LL29R/abcY2uVhLXV8lIgaMGPsIdiwqVJ5lNsP7x2b7jzpJX1iU5i
0sKPgLgwZq9MABKjPO5yEjBAIeqrv3v4AJJ8rIU/bY8wTaVGidJo40JEuMt0LSdJVc276W+9o2ON
FlvCOIuCPI8UZTkTYx47P1iP/aL6uisyhvFU8L8WEkfgD+As2At23QFFa7NJhSm7ptmr4GQpzQTs
cHyPm4kiQNwjcm4b5QFvBnNE4sj2KSCctYMOBSKSOJ+gKKPRo5IgHR+lq8piJs88Wt65+EWYmatf
Xf0y0JpD7dM3zuxX7UxWiVzUctH5ZcT6fAgje8iN9j5gBSDjqmjgQQyvT8rHtht3hd1p4lnV1rHv
Wv17Y9K23VFOTAWRHaAnqt2pZgoGxkbkcxchalAg6oAj3AOS6zIg5mRb7cjQ4lqs7FY6p3Dv8Zfp
V5H+VyAVjPT8gn3eoNaLTPzZl+55RA0CdvYcHh7rViMXHvC/OeqtUmEywVBErpYShwEYe1FfQTFP
uGNf1DPOTLY3istzjq8FtottL+4uhlrFEJhYvlSgrcI2r0y7levej2yls0azkfFY4iZUHQms+pH4
zzuRi6Q/4xVNubOs4+ay4/DF2t6/9DMnNK48/MjrJ3FRVfiEnlq6zt+u0TVmBUJwWta0XvUesPIj
N74eTBuKH7/+3Ic5J0YJXbXC0SWmAbgFj+nYZmIwpahC/cmvagpOobeV33Tn339HHE3bwEPNaZW2
f2vWIivOXfA+sE9bMpiNYKtFoJq0rpQedClkQvAAuaPEsiMhQa0pYeS8Y0BBzDan0asJRfrO2S5c
QC6DEKq4uw3aJUuL+MXgj5MqUSeg/TxzcJz/HWglLVjbZMZjTIHAo4FZ1Bar5gYu90zNDOOJ7Bhq
wcOg5DLL7QJOKQNiYPhzPlehDoRndEGI6KQWAKhHPCXjjs4dJJn2oxQH4fhPA1ELO29uKdnOlkAF
ZvkuVvjtezrdhHFLg3J2ZGhyTIZIya/b51e07jcEMm5A3tJ65EAFJbmYf6Ht81QllJaR0uTXCaC8
GmT1cfiSwzi8+VLZ2aG934iw8ltTp1hsiPgNMpZr1TADbTbcmnW2LQiP++vNXsW03S2IWHezvbfn
8aFBP3UNxKikfg3Wirgm0fT0omELJs/X4nKRU3wwh+bPlSBV8lEcvF9ruhW8XDoXb3/ol10vUwSP
k6WngtbLMy0VxicrduIQD9N+AEu3b/nerxkKdyqgg7Ofifdca8pZHorEl8jubGPkO6A2cy2fjuTF
wbxmanu6+GwaRvoKTFtbhbvQXQOOlp1wHue6Ymbvy4UsnPRFQQcO9WyHg9qTzwdB8nAjdO8QGNXe
gTvF2/TuZ9mrP4c4SGgYxm811AyVIqgWxOGK8yveLyUIyMf5YOluKMaebdZiCjj5MG+tLzRrGcbq
NmMinVuQTZcrKHIDgeOoMhWhSFZl+8uCl9Lnk+QN1hibjtZ7v3HLz6cE7F3XZEfkuZMRK1JiAhII
6QGF/NT2z6bXp9FRblV/zrnDziKJ7hYCsIMcjB5tNlVSiT6ENT1C5HtYOSPmmJZfIXY7b5rzaOhV
UIIcVtDfrMpalPhtN2rDyRhyKIsg0MRRXgVB0COXJTbF++0IuM9W5rDCJQorRDLZXz+unxJ6EA5v
Xp7wSEzjesmldeU4LbWkxS4gLC9S93UW6dmkKJADePaGrLI4gI5rX+iclD2+H7qlE9I4uFAOZyWb
LG24F/iP9OsnlH0p9avz+TX/8v1LByQ0DxOtPEh0aAQdsaN3CW8OkmgW8x8yR7q5LjHSmGBb3xSV
3peK78739SUkwG10hNiV7zyqI1F7A7bt1HHwmXs0QvYBU2UxPTFkQNEzMGA9bMezKX6eiKMUwn7S
igGaGw+aE4J6XLFEfvuyKvdRsxEcWC5q+ZFqdHMBfFweLYG5E/o7vITgHM0Uom8XnA5V1KrhT6eI
DmNQlFAfZcDHDPCej3cprB6iJNF1aFr6KtxD5Et+ivJDGT0+xO4qf/U5xzRqiGNIYu3FMhmR813l
8tUxLruS+aA22RDlkwrzdSUDkwLsgO510zMeG6Dy3z83TYNbVMW7UImdA4wijDSAtM+MLk2ESbb6
bfMdzx0KXV9Em3dOSi7VqMtofRe6FZVa8udFVdI20xKz4jUSQSNbSx/iisJWZj4qSYTpiRMM1yc+
5OJ6HpJyxqzNjwUEjUmGoLjXK9GR+yTGgw5PII5Ch9lN+UWjdh6NynDP/O0W7eBPX9Qly77fkVgs
mkGBsRCWWHwdpWQarQK4U8tWODw9ivnrWtFOEnVbmvxRyd3+Zh8NgWg9kQc/JfcMKUheh+bEW0rf
19A6i3i0Sh3LjYGvD/l+IwMNXONleZc+Bvo7bQduab5iuEA4ReYMlXTAWeyQLBBw2K3JqUhLfrEd
fyJSC7vGXbQW5KpXMOmH+IlV1WZwHkkSMrcqN+0VveJ0rnXz2/Acl03IxtZvcSmHvTyCoMn0YK7P
OtVPMmcgY1Zu2xZqUIqMFrcMp/lo6R+yQpPRscWa7Iuz+DxF95MNWy0c3XYP8+33rv9d+a4gUVI4
/tJKe777XA2oYMB853yoJpgk5GOJ+rNW7ONhR6lunYlpnvPtykLyGWaKS1aE4x8WAJoRc5jdUszl
5uLFjp7kyHOTLYzP4pcf5Jrj2rqJXNmvViiGqtrnXMzIOuDHfBQ5e/8tSlKyYDL2P3nmvgK4FcOa
id53y8U/UoZpPd9uHsPu+SOhiNOCSp083nqukuzsttaDXVfO7Vyw7jn48Zxw3ts9ZqPQlyamsMZp
jBQXJqQWXR0tBE2LBqSua0Y5+OsyDmAyy6jT/zx5/HFvUh7qysd0wsjUhBmZS9bbaYqC4fLWzruz
U9Cr17guZudxHYMA2fyOTZYC56XVL5SfHEFWaTF8McbpSJypWDu5kEAIzXpqdiW1qEObJ12rbavS
qq8nIv0x2w56ND18Tw6C1qztptqCUWNUeEXIT/jmIIgP2xyZcXVr1oD3Nsg1oXXwUCS1e+quENfu
zdTQV2q+fJPz7HycBAS7u+cSwAOkCgsbBAmvXwKXvOCZvf5hXb7aGUk1qpS2dImlsyMADgc22Rki
HVs/qP5fqx684yXrJXKduvyzp9ULK4rzlvKOEKwF6Tl9xdxhb+FMuOURgDa+EuO9ky/a1DTdzz8/
NMjknqKB/qWtzSwnbgCb5URpjOyXFFJtf6UEaX2g8SF4nVDl99iGziULLTZnb/xwvuEEjBtapEhR
mHSszxPgA6p9YQPYi7s2J2ae7sC9Y+U8lJPjt2lnF0+SNw5cogC8lcQmekQa8kH2J3krx411/Yl/
+rHCmmawgMxt6ChMgKjiN5JoynEOvNj/jjovG6RjQt1X4clhleL2Jn7CA2AWjqLMGy8rLF3dkhRj
vegto4XzUn81j1c3LWwofNtWb82jAqX4/vYxz+GwdDg7DmeYcE0QpMc4vOAMzGQq269QM73rc1Oi
4CBELnWPyH/xxBAiS81OzwbYYUGXZLCDVafgjvOhXsHNoWREPkti6jw854tjd7OFFmtOzwe2ws+m
c9kd1T+ToYp7oL+b34SaGOjewfNz/8tmx3sxFNr0iIaBr5EXUCEB5Xr37TtEOp/a/Iz5GudNiU9u
+X7odIV2cJiJVA1WMNm4pCnM8jULDoGVIa2j96bEpbNfNO7CNxiumunvfMRynwrUGQ7BiLbBn3vb
0Ue1vm5Dqq40BLsL6Bgdno6Ho2HD0Brxn3rmepnvCenxLzFVfR5a8cn8jDq10GAw0ZF+jdHN8uV7
UrjU0EFWMRuL4YtXIZnkiWAJ6A/sqLa4ElEoAfyYVrAn/FVC4cDx59urml0+Ky/T1ZaIWsSiXcBq
w4gaUOnQ+kNJTh6UgrlIIrkC9oGKRtBLCYNLbVKezWXDPdAcTkyWM7aX6Y+j48glPkxcl3KvgMQ3
+LSe+jsA6u+1xa2C0SUneucYoTlA6FaG1wpqpq2zNmrUn0N1EJyMaFiINov4NUj8Vdji5qp1hQ8c
8BPn+t4o8DZPo10uuJ6J2j/1Rp01DnTxBqVoHSFBob4MTSjM5FVEdHrRMEAal0+CNxI6S/m7PqiB
/pIjOTwLmG3bhSGsN+njpo2KgbkBOJ7JBSPPxl3d3dnyWDoihyR/KUPxMxo7c4eMmdijs4K/DjWn
sIPABP1KfKW1/DOoztEGHm4fiKSh0o40YRYnPTODxuQwsnKJDzRbd6rsMHTVMaQAT3FRcdsVA/D7
Z6+wfV5Rz+9dmO8Sh9M+IPjLvugXiFrFRGQVPpJ+HfcXNduc8hikd/RyxjJgTYMHJhk1Qc9jmqYS
gltYaU3p2plUofG9UX/vrD2kD8fbcS90CvlPeoaNYpgH4wnfKspDJHs+NyAwJKPXb5j15NYY+rzo
l8oev9ldM0vD1aHGvMnMRxomXr5Bd4zSe8e5SN+FuDhIyoSzNzdRkiIbw8qugopja4qur+nyeYj3
mbDIk0wvGKI2w0ahrAUQ5wsn+CZXM5qDAAtvUUWzpVWls6387nc8RV3cX6RPB4PIUiOtzuLVGZ1d
VmSBjTKls2xrmdKuiBJWiQfxpyL+hO9v78MoPRxkJRaJMmY9yGa3ZTgX5K54Ml3vOx/4X9zaI1pO
ozl612KY3LnSQwdDBl3Vrndhbcm9SXzN8FLvMV4/v4bIps8CCM0ep3/JaKvnfHJbvqGaRwESYzX0
+ta4KfHBgAbS6RKC+Mq6iON1V1IIl5OzRIGwf7wgffNB6OWx0uFsU88trBInJom8snTcX4U0FWi3
2E1yIRKmeoxFAvuM9Qpylm9inX0IRqHdn0wgQ84zwHVKkwI+fVWwA0UwFzT9a574QHtOcj7BPrqU
6FMxtsPtTm07jxLRwgk3uJFeq00B4hjRuhNtEYqFNwBNXI7bDwkxh6bbmxjtNL0emoITuKtAz3cQ
LX7X4s36Yoc5aIKeyqHzUzm+PNQUIXCGEbxb3hIOrnWPMOtgg5lDhLtnt+E4+u0fRY83C2OnGO66
ykLS0oYplm/X6jL13EPXlN/dkL38uCBZBIQrF8BKSXYOB9VrBZkoNPqWMuVNOFmkWMc+FA82Ts5z
P6Ot6nr3Y3uwYv63Ten+fhcGTMPJQGIQLYe5CCqz4u3TaIV1EQ9vLvkVHvMpFU4bbAl99HwV2rb7
h4fwW2MBirxv8aZRr5MLjQPGNYxFPoXxE24lumJyvFw1XCxKMcW73L6sU3kGzfwymEEw73bHlMjq
F/7dpeW0/Tt/WmIYTfa+y4OchBqTnXRacUd8b0TcKJqCh61mQ0yHonQJMk4Sun4Mx7zspfMQCRGx
ArC+WIfwnme0j+uV7WxZ8rVEAYQ5wL49xd48Y8jmmBTeSPZ8jCKkdzwOoPon6lYHj+rq/LfV3AKK
HxvkJkdJQZNV3N1GloxBBa6cNOFpcSu2gkqbDQu2Llyn8Co9O+Yvk0rYbP8FWEZSf3fIa5WoJwhX
ihye5P8VSocNtL+I9dnsBfA/QEDVThWiAZ2MI55I7vLR7QVfoFRn0JiHDxnq+YHzDsIB8mK6nOZE
vudCbvmmspHDYC00pq8wR+5CyXnkiFJDglVxQIXhmOqeK7+X4kdnt43tp7MPhgZTGcxiFQ4GLCcO
mDAM+D188B9apuJXdyTCmnbEP7O/4S6t2mLVnlB51Df6A/V2eoDzFhiO/ZrY4wY1Uy7DJS68UNwq
EU4T8aD9i9Kk3HLCr2mHRUOoHg1w3qVGRumdOzyFzAFrfSIn9nYIFZ7q4Ab6+XV9bjOwvrI0MFEt
BJUHt65amGg/NohpyVjerhWxowXI8lM0uAj77Ldwm1/JJV76NJpZBINSDQAG4EsYHlsKcLKuR5Ft
V2k+zattVmgQOLJCgProZthXUw6s9oEOZyWgpEiuUSTR9JSUxoEniKX1Z9U8LvdK+QcJhTYHkjYJ
Uq240ygcrVnktVIt0ypUhZ2Zu2Qa64yv1sshuWgFwX11k0KrtMFZTGN0wIQ9UB/9GMSs4OnapR9j
cD8KoK2+bofGQRbHqrgZkg7p8yrNuP0sLq4ZqDKe9I97VclSntxswo5tUucnZppakMnGJ2r1oYdQ
BHm6S5cMA94Zg0f2VyaEL9Q6xYQHC++THmXeilwUKDGDrzSocc6NRmSvqzw6+0dceUGzAPZ7MkVk
ZdztX/oBmhhtJyi4LoUyVrbhaNmoGZDOMlFNRmZms4HeLWRlwp66WlfU8bzB/EHoAOlWwSmCM0DF
zpk2F6NL4IW+recSIY1e/ebI4kwmyNvWNb+qeg1K9gLxAOh6+e9n7oK4uNAqoCkRQSSBVNdnIcMj
UH5PK1jrybYBe8yoW+8mtBk650RYNF3pz1IwsbiV14zQMsGsxZtyY70PRQQqeM3mUsmgsMFKPo/j
Rk3nQW3miZRv98jeazAXXBABVo3HtOYDI//1UClcf570dGTyslP5E/mkab1a+c8V1AFaRuYWnd/o
xIa/FYyj3D3y0GVEaCupMIltLOHagQEs76jVA3/YZH9R9w4SffDZgKspgxcGgWSY3EImta7B8kLA
8H5YRULJnETg0JHddLtyD4Y6+tHS1x31eU+whuQbGVXyZYSIBurIo9y28hlwmb0QbFej0RYHLUwb
X1rHi6wGVf2VVwIejuHeU3mjFIHJnfVc7AcKvdkcBCUUkhqYjWacg0z9sPu9loxYBRLnKXTRC40S
KoSTk69LpbRPuTz27JrfZvhnHQXbcpejFmOkpwfiGnugbhdWlOkwPjbtOuM/fXccgjYyV8Kz4oIG
JrwfvS8geyjyeogqduilbbuii+mDmMO/e1qV4ajtB3nckyb8hOqsuriZkC/U1sKUHe+UXRnjvCAJ
XNc7d03xzh6Jy2SkKyqbxmJJiQSNDHolKnAC4mQxO2CuzJfwQjZs80JQEeix5xihjjqTo4+TRMQ6
LrEmRrMoWl3/6rjZzvGRZeqD3nyZrLzixByQwgl2GA9pNDbkqSXBRQoTIJTnsTrITpg3VlB46eug
jzQXRP5rFNi7/B3GJ0q9M6Cq33kR2EZE09nweI5VCRBHGyG8RjG2kyvwb+gv081yKFc/SZtkiIRz
o8JGQhcNz2tgdVwr4QZWqOC1vRpBZ1/LZo3AvKD3GyxhtSiE1ERV7aodWsQWzX8agEhHg/F7Up7x
/ZGrU/HlIRU6tvTTRDOxRRSi/ag0CYZ6MvVMWZ8ribjTLvOjrCA96+AybDXvCI3okgPhKpvXk/rj
j5UlUazb0YVoIU/xXz7qLoh2Hv6cFafYLHJ48gy/FZO5fPM7/X+5f9DhqruP0sSyIlb1zQCaQqMe
qLt3cQrDoermKnSlax5RaKs417aayt0SxqklrdKvZX7X+SqXXpFWGiI3/p37QgjheY1k8eGbn1Wh
l0u0Au/mb7qOyjp1NwKtuu4xJVe3VQPJsSrIsVkMC9BYnhuPnIsk4XQGv17WjNg7ZIqtdTOfa6Xc
TbAgxwjrgHRZwutjqN2Ojx4Zng1sNgzr2S0VQ6WVwDf3I6f1FvG3N77ReVMlwab5DdRFV8S6bXuL
1IDZUoudEQ/482bdu2HbILp555ywkpalHNGt3G741GV0NZJTssnn29haDoRnpxB8dEdCABjYodr+
+EQXDnzVXiWrNJDprQ+c/5tSIorTBqQZ5HpQuQ45fSdoajaZhKX//hVD1U48lTPiIde3xYY2lEjb
3iNq7FtDRNKvDQF+LiTKQL7Onz2g/81fjvrJoIjqYVEGVh1M95+wdzYwJkqOKe+++BNPQL0MVL7g
nS774FZi+52WgGUC0RV+QMBtSlnd/mHVxZNoxIG+BDqxLfmfIl7cjHhWz34FVZ/CkSih1/1WDle8
4da6t+WacHKuBFJOvITxH4vCRcsHgXDvXCJECpQUFavlrtaB0Jhm4QGpdRLiviw6itQ6golql2go
NTCWGd7xReMZnSAkvX5KbyzsfIc7JiVM6EmmKeXbxeJRhRgT//Wr/zTTlhH275iZ7u82t8Kidjn7
4I6lkOHRQAiX/nq65gkKJeV8jRZ38x82CsGtdL/+TFTn/v6b4rwoLteOdrnRcBbUPhyoii9jEBn5
i1eEVT7BuRto2VkBsPgP4v0kFQxJWT4XS02sY62ag4lV5CgE/5wYFYGD52sYazF8yfegDcbVEbRy
+++3yCy79k9PDyL1WSm1NgSkOhxwCjvWC+g569hMOPDG0IvyXKVYTHcaABj+9XZpT/eJ/1Y91ANP
a0l773vEVFY804B1CSPhJx/qHTHm4uxWEEReQ+pxipaGL4M1RBIPGeyCdpiMePXCO9ftixoT3oQ/
THeF9acVCYGhDlvZilU3NgcqrSrS4nJ/mlEztQUkTEu7zcozcubr2TO0VXcRvox7CYcBjSSNkb9E
uF8EQd1xb14oEyPnKwdAX6uBnWjfg+lEF+CHCqavsUp6+amAnNYqcNZcYFeoKF+i2sVJvPRl8YLB
vrqywVCmfxE0DQMF9EKR2P+PsSTwuGKHyENfRkTzq+MHolnCL3ClHZJW6J9dasQ0TEq2hyXLqMMT
bdbbGeRbKjuTFFhjYg+ZqWJbD2Byn0MLj+qTmJbQ9EabFDZZ09DexOAvjiumX1KNsSrXgokONA2g
CbkhFXPUTxajQ4lZeht77hMjDdhGNW5GEZnatQEEk8y+Jwg5lUwc4aHV7chfzVtlwWToUqNE0SdH
IqqcmTfmDGjJ08MR3RDTOiZeLBAf10oDlNZFxoAwRYzKQmrxPleUzMsxR3+I42ealCmKuBLK/0SV
DtQZWO55h/R+az3dpgsMk3rLgKln0M3Mdmw3kpU6FxF/UeyBOC3+JGL15xwFUv0rec2p2280po7U
DCCEaXW5oBi112Gd4JdjYFahly/d+GOV6oKhKoHHJyRStMO5pH7l/gdxHNb5SQYfuD5V3QT3fTtK
7N21s9WYnVO0wGie9RpN9wg8wLMjHCABCi/td7PAb85qXjyLRbEgBTSSMdDK8xpqSLGKQ/kGTgkf
ODZff7s7FuZ2K3W4vpe3B0+I+iTD7xdaAyx8p9vKMW9Ujjdlypsdzuoo4k/jvs9X7oqYDBXSvgfb
42ftcrtNd6+2DMaffdl5ftxPXaQ3E8DO2/+vIUXT8HKeS0hXVwV7Qi1vA83i703gqUJ5R7+KzFO/
66bXKIUuq4xA4HQRBFb0B8IWj4zjmaZb3p/751G7m9HIEnlwxU46x85EmWmxa0WaeKnWP95EEGH0
KDKjoEzmVeJ41Fl/58Jj6z6/5/X0V7na1aC76sVl3WDSq9qiok5r71UJ63s4cornT/ULJrSeif9R
mw3+rJI4QDYHSL+7W/SbUupQNxOV0xL8pCUcX/JnXMbqPDXxlfJcSWB1lTvdCR3txoH9j58ngonu
VUsNCCWu9pL5IrygryE7zHWkc7EZ8GITC/N6wsIB/QF8sEOKp97/wVzp8Md9DHq1/bUifhdcbB7k
Ugk4AchdfUc6uazJ5kO/VpUfaAZaDS08qZ/AviCvDFJ7mNyuwzV38tSFDSLWylaCqcUrBOZrRiPM
XBqEHvyM9tGWpRm3UaR7jEewOi9ZB8UaXRa99oXETTKYvaFrRRQxQtWY7W+0ZBU6sKQPOTY9CWq9
H0KR6trRyRHF+UrN418OotNa24w9X5EmXbB+TM9Rj3l/17qL2aOqrY+rIY6+1ouihd6+lJj63Qbn
mN59afgFuaUh/uHSh1JJ7MYDJWLjvUBnNfzfARBu6bLWCwtVhYLFFFKIVozdb4A3h1qY4ZiIP8Vc
kW/EFWfqdpUbKVqJix/PqKAeoPvtOu2nR7GmXlL/BWEDMbc4Ne9JQwz604wRga1mcYA1GtaPSKz7
gSxHcrnPZxO60+1B7g4cwFqyhOeClH/u79RU8PlLmhR2mhnZB7CYtxRxZ/hNyDT0uNU1cabFmde1
tvR0aNNNXVt9KUCjmz6PauFu/lkzu0ppABWP5V0v1OYsL8OWh68ctaDeJiut54oPG/Qawq0JdKEI
riuFPeYCU6dgiE1ms0i0BLCXr8wI9l6FIHfSxnzNjfi+YP7Lp5E2SaQ2mYQM+a220E0EJR+RhPpd
tPcJOYvIq95oQWv4lB/lJf7UztZdQPKGVzo12+fGr+2g9hLsfrW/sWImbRztuWDXsK4hc4lA8wg3
OYfXlhur6a6QZHzwgnhO2ULZR5qRWX59Dxw9OK2Ev0n5/OVckIEOnKKOsoT/+b3OHtL7mZxalmYn
IokB+pp00MKFO3HivJ2AH6rr9X09IqMUiYPCaFZsemDGd1KNqLz57IKWIrxmIdvk5X5sRtSHMLB+
cA9i4RWD4v74/CYFQtemSOee1z8P4NrUO0YdeWvny0aUrE2HBN5lTnu0rc8GXPlb7kXXYdr275nl
O95AJCwrmAG/E8RRe/NM1P2eZHFTJyBp93XCc3Zvwkh+s3dqRooqeI0Yfl9u4udr/69zZFD3pxy5
/+hoGcMkU/bqw+R0wFElQI7zcBqgEDtGvuPpe/JNaYgrCJhao0T9EExT2IQA8YiarXsRQ47Za/sZ
2ZLLwC6uzp4n1AK4bFN9/smZbGRFmjTfNK1vRuamAeqtUkqOSQZOSoWQTeyeaG771+LRfFDaenfW
4R2GTgQ35zLKkbPmsKnwPYkQCYBSNuB3G00QCxDkfXNkp9fmJI8v04UE/nUerCarEXBGTiXaoam1
gAaH+JvknAG0eIDHTVnLO9pXpB+IMy0GuXatAAve+VWw9YEp5IH1j4Er9IayjqnjUmqjXEsPQHm6
T3VuwGJWOk+6Ay0tWv79LpGLgOBPSRUNBS2A05CAjkcuLNHd/s/CNyaKSP1s2eQwJkiupyvaIyEO
FFYrHsZoS/Mur/jSwvZcIv84ahbk1/+ww4/3pvd9CseTk8dWUs+BbmaZivQnhHtsTL2YRxmXHALU
Ps6VjGZJRmGohEox2i4hKH2Xil9P/rrAGNz9fQCD2p9ZZZ1szSM3nXMbF00et5nDXTbtRo9dC9yx
JdMMq7AfANQsa58v5nByppNpjbpfgoUGiKZQnv+7WacxCEoRJPtdBX9+NqQFLlFMAIjY9ONApyCp
Cp2qQ1jy71t60mvLV5F5QwTCnpOgcEap+t8lsyrOI3Z7Ex6ltjdoWRkPcFiiz5ej+6BKT55rI41R
CXQMQi6kcvoJ/PiamyWdo1tu+PDbS5iq5vEwHuW5+o8OTOn+fmruTUVYLE366qKtjv6vrWiwbZcV
QXYhlUofmjwWm7O5lzPqSh6pJRcdISFOr7jnm2xeswjNiaebpzRuNyh58nGBI+IjqCQBI0eE0XpA
S0c+04J9vAlus6Z00ZpqWYsrsjjYhCqyeNSoNsYVX/Gcj6u7bGohrGfdQdyoqspTbxpoUrs/SM7I
wzXi4+ocTZodCIcgdwxRpdMKgGU+58wDDZ7J5Uwxd0TLNxhzGAuHgYbiMMfOXX/dgZZBpupF8mvW
Uz529H7o+/KFsPu1e1H2qeoeIFt0MLC5yHIuKbNsHpjy+woUIL+9cvljQY0VPlJGQQi3z8LIJ1KD
WvK6QGizQZLm3KpsDoW8Y4LEiz+0FwaH2tG/pF3LuQJYklRB6BnxeTd0DZ7mtNiwhbhx8bt2eNLp
qLI/VJE788xmBbnfdQjldwJky3sRd71yCcO+wncPL8gZA6l70ZlrufonRmaZLWYfZ/XGpmCDZHHX
dj9IxUDos5adcj6Co8jPsFfqkiKCjT2iCW2srlIAI+0cljV/6auxZ47XxsKV7Fc0l68lC88jmumj
OkPGBxaveTrv8VODl3J+PO4k/FhWVlL1ykY6OrN/NyFwXKc9mUVg1zfXoCoZPp+v9BVt6Oh+Y+5H
kO2DIVHIVdZ7PNTAineiX/sMe60cs2DLi8TG5NZcV7sS8xBNDMk6TUpwZE9lcCvwRKWMeRq+WqtC
HXsdcmESPJDrD4roY0TBlzomBAcQeGwd7CwP2EFUdAPhpnrkTfZdrWv5qE7/IQQLikZMpbCArXAp
MzT68ubhh3HCMoYlwin3qC7hQsBPmYdCj74cu896L5uB4NSUSrnWZLWeeoGyILbjVNDBQJPAPyzq
sTmxhjV6tefiUcEWivJroElLy7egfCxYelY2mvAkJwCb4MZiRRhZVdpHhtdQrx9vBlVjdpL3YGW8
yOOEDwfYLWEwIBgFQPj9PaLwgAjg7CQxO7avbESqS6M4a0jERVzbdUuspnThchYklt9eLdBB8O8L
7cpRmjcpNR9PADVLTVfIDdWGJq99Ns/GpA2kiVDJupG7mjTeBQ4y3pbiq48QheK9AuMflgCsJUXK
UNI3M0nJOVywDdnkGYSMjj8iIGeJXValwH+S/LUqXoRnYIe3Su+oJwMXRlAQ6tDMf2GbQwEgaZD6
Bqb9pS3LTteoeeJ3t8Kuu0W9UOf6cPovXwM+qt0ndhoJMnBv672wTIEOmDJU5QprDQqwOjMJH1Zz
C2zFAd+2hyvbK/KUQ5jwGLinppLW/S/6jJuch+JJjRLoCmTsLtJsHkCVtLarS9o/5CeDIdACwOX6
u3lZDAeMqdatuXmTMoNx1OF+tF/VtIg59QAxIY62KQm70+MarSR9KZljnREjAShL10F0mJ7R+van
x1+Au+YVRkpM/LG270k6iOTA9JuSHn3Mz8i3fXNC860W6pMDiMGf8mFAkGlwfGHtKl2xbtNhG/we
ZlmwDYLE2ycfY4iGWARfFiSBGzl2q31Sq3wmadB4HI+BGET3NQ9Ph6TtiOgBH0IRc89PB4MN6uFq
lAQj3W6Dyv+3+U4Tf2WJyIjZHg7cI5gKCOP6p0rvXnikHyq7PJefPJpsJR8ITsUEt7otOilzG9iw
BoZDIOxwnkpiMrRL3oE0nhKQbRV+cpboeMCGutrSVdX0QNYhsfHR2WoC5Ok/Ha0rx83KNLySt/sz
KecYL9IL0LTwsAffp9hY2djw7OcAnw60ZQEQXNZ8vizHoF/+G8808gmX6vLSnQx/7H9nGWIdg5Ko
xjCqdAbW1IDxTTPBtKDrB2ghIQFdRVXGOrSyb06FmI0hcP/B3cFDgJisay9K+o7pm8OsOGGnO2Qo
C8Sss+fBPodjAGBU4ObQUaxVW4dtYnmrzGUQrk5PAqTojhz73WBKSgizSVEncLLViKQxRk7BBD6a
4h1+BayDwosvs9ml81YAhW9WQsLkbCBDwA5xPMuzJOZj0LsZ4adEeHf8wToQlD77sblwcJ2rrvP3
XEJOV3OvUmaitdTaz3TY1pAD2htiwXclKSqKL9GtSNpILtswxxURxjXo5GdNNyq2yi0ojn2Yamix
3VY+NwPdBdPJsPQVkK5P+Z06j7dzd2oicuy067oZC1PFVw0Lqj53j4VeDAv7tl2kLytKZkIVnzBI
bg9xMcLC1x7QnlJDE+gPK/F88fiZsoHJ2E1VukSWqzmt4DRE7n7kTlIYIBIbysmqHLFyB9gzK2lq
pWENu5CDCeMJr1f6ommslhXf5zkla8EqWbegFcxGBQ4bs916klgJPnielqgsveIC8CQBNTQoK68D
xJAL1BOjMFj/eNGbtBQ1oz8DMICgGGMlpLDc4LJlzjwKPgs7EdDo88MJPPP92B+dhOv9Xer1B4fm
A/FTxSLKCD38KWvTIZbtBq/XwOS74b1SFu/mMrx2QfgLFC/sax2/j89IBSSFIKBkGopFBMrBq8Nx
HMt+upgvqxttQ+OUwHG9nJ4Ev6WdW5YiuOx3Lz5gLuQU+0gWST6R2Q9sFwN3am8ws0PFeEkXWXEg
vOxkSAYThPIDTESVRb6GbLyT26aEHlyQwQyicqYYK+dgKyLmRpmvhIIUwnvS0NTd0Xs9Zb37LwUN
746HOyLdxvONacoIucHvmg5Hdd72BYPMaWGsrz5f23Z/3lABOYC+HOTF/2uVS1RcmFpEK0fLB5jB
Om0qxkK6/ixEzpNdc9FjzKTBxBBhZ6b5f5noAdeoyksOysKt7T+YTJWkb864VmvdEiObblPg54E7
scFMz6fRibSw0rsFbGTkP9+rAQMls5fwFxvtA6cLhfOX12k5peYsZqhvym7SxedgucSihoC+vh48
WIwTUnTxf/RWsF9/HPxI+/CJhO8eYd222p65v1fChMDXC6/wv1lWDOBi8sBKeA+VWbIyCtAW6xzG
dTdue3uMBfHbwzGX9hZwDgGzj98JJXhiPZEluHNBUoWxrc8tcBQ7nbNyG2WBbFxEuPNaXqJDgLcu
/oXdufCRHcy50SmnO6t23/SZWjguQgygSKcsyFs2FETcznaLukZWuirPYLu7EKet6app759cSMtU
JpXy9zr6Xuiu3yhb1P6I/0tqTBCQYYZN1Mq3mMajhbiaa9wmREFdZAITzA2LjZQnZ3Zk4S4bHTZW
G//FYk1O+XLI9KnFpeTzx6YYlMrVV0I5gNoP7YCPaCg5DMJ0rmzx/Kg1rDEsNXS1+hWUt8UYfEan
IWQoCEj+3WxitkGGpbwQCYesfB60IRAhLsWSlVU0YTDLm+cjAUzLEhcy5SAc6kxbFccT4cSC2elk
wFE1tHDqm7haWGx1e7rCxDB/J527ejcGUsQFtA4JOaptsVFIyNVM5cXn1tniuY/Iz1r4hK7KOQbf
yH0Uf1hZtb7dcIlpq/3T1mCLqYkJXP8OIvAoCTQMlKVwM7eXVuXDTnPvsfawOXENyBCxOMW2SAlY
Wb4HjydcPR/ScvjH/UTOytRzEkKUCa+fOefo6Q7xdEUoGlT1mXaBQjuY3IQJqmDo2CTYZ+PDiHzs
q83zJuhD6KlCs27nyYv6TWbfbQU0oi1UnuEORA/h37jZ/OOZW+i6pdmeoAqjWlPbFwvecvN5nQ6H
jOE7/bJeefM5ik8QuOEN198pzfHOw2cQMdyNfberymMhfqWqoVodbrYgDLmy6ubooT89NNFLw0L8
McKy67G36bt4b78Jvr9FzzsmXLpJ6uyALtl0KyCg27gZWSsrWzYMuCr2PWIfoUTmgV0ErcGqtu/8
GBVmD6C39MmQ9D1c6HsbjKICTsTTBVPNOBpUHvxiZ+NGsMBZZm+oIm48o/yE4wh9TSNygwLmhQuZ
0TbonAJ4+YSc1mLgeqvu94J4MAo35B8LN7ey9A6GtpSO7IFL/9FaCs7Kv8qhsVJPmuIhTiXKruAy
PbUPxrVLNCa78YF87chpqtG9WP+VP6SvhqpuUTx5JqL2wx3DL2tWSJrSIhdAUgWgCKezdbIIR9pJ
T8eruWXWYIS5SVfPmB7unPPcgLuOU763aLAMAtavF3P5YOmsFOjky/YQHvmGtJH4Ua6+Tos7twmO
hOGFbmTsYrrz1RgRh1ir6dngGRDDKzV/JmKka2U+Xr62H5epw+px7xwxlo7l/Zqry5lE35By2y8D
GxcXHBFHnhJFNldLeO0xAf5DJjeBko09Uv8Ra9fEysYoA4DKQjqgsVv39xiGANOoZxFdTPVfLcTb
fwc17HsJ2d65wjxucJU27w1QeR/87pf+UtOOn7HviS5c26AIUEOaKFru5nPSN1Hl8HpbYArARepP
+AqU4gTmJiz2GZlznoudIAxzm67q4kNUjgqTIQyf+FQrrjkMR7lZNfRuyLhZlr1S4eoE9Z8vrPcU
1z1keqBQ+ida41dZEQw4nNlQw2E5+EhiiCaHpIFFP2PphUrRYZ2pfXHdPLRR7mtHj+GN1LmJzNwc
+x2x4FTzGvmBpUB6zlS8KyjY3u/tFYju9ysCQtsbBS35hnCk9uO/KlUndDW8xcRQCGgFr1RMVmsU
hz8JQ+4VvbttKL0X8IYyxNvB1J1W4ZoEcvbfKp/0+Qiv1YhogJTS4y0z/FA72cCM/lXsOvgFMs4t
RssJZn5GGQKbZuZRl2GUmMIK27Eq3ao1BGkKtjHHGGM5pbBPbsplzRKDwss5NgdUUmj+Job7FyCY
j6XHkwDmoFMLBK1mfrmOVUNibPnxdynNq01o+EeNBxolGcemL2aY/7khI0tVcRUh3Pn6U5AenM15
eAA4d88KnCr7TyAThnWisCrcMiRQ8DVWNjYbJya5BvvPD41LqMq5HMzTb64nvCI4CgJnamFAl6IE
kqTW6wGiGn8x+Khpwim0cJsuxfXmjvrHbl7T0c8sPE+YuMwAyCLgIfak07DXrD98qbIYHLUU+Ddq
A8ZbWrKXU8Bd7vYVjiIHYNdn9kgp928XWQ3mzS5LPVB0kKQR3DYpZsrJ4XbdhBs7MjCHE7exPTAw
zI/71+q3fSQHUf08JMVkG1Pwy/KUnDcnZqdd16Uh1cViwf+RoRgub7KvQky6tUFAlrc8z6tHtPfO
UQ9c5LALlTNlc6IlqomSuRz9nNJGgPdHnp/RUOg/2OkO9lwnMPhgF9FjKOQYv7z9E6JafPohJbv2
Tvi27H6BMUNMW47haVV0neq0pHJx1Nowey8e4h6CQxXkmL71elkKYVgzGdXi7QHSg9puX490NDr5
AnXNF/PrL9jXHp90T7C0En7wNiyyOD8XlMhB5EPma8PcGwGM8OD3598+rsG+AtCjZp9BfVMfNLV7
Y2UipvVCtCdiKs+hGB7bMa1mDf7CDEPOCxQUim3qT8cRx9ZrVrFzxFak4lLd1YeRASn0qPkvHgyw
CA9upeixvrEHvlBvbpIqe3jpaZbCryP1Clp1+eJ1sXmZt9wHxYZ+zVeex2Mr5B4hAN+us/d1cWPg
5wK0ajskPRSguUEaNUbcFP7x9frTL7794JqtbypiBtpXl1xq+ZmPVOURAHqfD5P4Ny0GcKs+enTW
z/wV7+cwPntwpBLkEqxMz6GbmAjSmikexeni8aFpmWRUKTXC+eR6k/+OsO5XybOkxugYU1gZAcI8
6AhnrVH0ktfBOfrGSjQ+yPI2Y+Sy5mLLIe7oOhWLh3FNsjJj46Nf1w0kfiTGNXFRyaOvqbTC7OkN
9K1+kTtKcOFaeWsLBiYKCMMtugFfQW1AfLaaR5o1Esdwj0WxeVzWJ6XGkt43YmQoNWR/veuWN19I
s6QQ79HMIcw2riieu4Eys4mhzwUb0T+5gsaFS+zim1fi7QnPjBEcuPzFA6MznWu1g5i0LuynhRbo
7QauycyqwNIaRE1DU7fzerhzgHa07DMC02B5nOqyqzTdVPeMLnA5A6jI4z5lUkaqY7vo3C8JoVyf
UtfhT7DFkL0PsNvXOfpv1kyHREHRoGvFM2VbRQcOyb6aEQyGfYi091ZqxEtEWEcwf+/NZa4YIpwt
dE8ccyn5G0z+HTP0/Y/diEu9eSFdkYP4cl7aUgBPy0D0vJSDNLHAnivrCIA8KlTjD8NQ4aiY9YqX
FmC7EjScoifz2pUve+8zU1Uv47lZ6NHEfRO1uYVZGUxgmAy/TkVT3Z9eTMVLFwyGOgY0vSluAGaX
ZhHgwyh1rNEA1jQ6n4y26+JMn+XnP3AC9gt/5iLl9lTWdYls9x94QTsz+jKpJ0KaeXnwBmuCmDUY
cvS+eP/KQ1vWjNdOaJmgXKf0
`protect end_protected
