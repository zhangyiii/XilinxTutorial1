`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18624)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbkV3TO4Ee1mp364NJ3ApJ1FbWY3IB
02vUs3YLSDgyj9eZXMh4yaqzcKbXOgmmjbKlHV7VT/2nPr/n176PYqHpH5WOQgLDKVcRyUPmFCqo
Vp5sbvSZ4QuceQ/e7X+XUNUhZ3OzLPWnDOniYwtTagc1ZwJD8OccWAo3ob42xNhq100XFAgav2Ka
svIGe+t+WsRZO6eL54E2sqqxIySewOzEWm4PIe6ICW+nLDZcICddalIcZYbYiIdS0JehmWwv0UkN
pcwtSRq+STrfBz+r5SXKYg04zc/jFKH+OW5ygtJTcL8OId1LA0QdeAXzErkGkr9IOv6Bw5jNMoGK
JlA+ymZaWWvovxinBl/9jQgvA66eg65RGHI9LRwviz5JkSXnKONyzUrcjyIBfCLJphHKm5JQTbI4
tcMGEhbZrc47kOjgRSJQP5BgF5kqX8PKp9UsHSRK4zoyuX/ub2GWl1JvwYgM41vqPrC/jpRTNCeR
+VcjSwiGjfJNAVhMIW9M4adVOtE9dRmR7p87BJ15OSKpVd1c7u+JYoglZUU2ZnX5P/GXRWtEXlPI
AjC0inBf/ZaoYZkrNcSZcN4tNUFeWOr0GnCO0Rqt5tWC9Msv3OddQqkQMw3JA3nh6MClaDl6qwBj
4OjCrNXvVda5yxN9JMcZbI065QJmBAnOK4uEn/hOEsmMrEhPUTMp1LoZS2vEIVnGx9DWai9FlOzq
+P8nxC3RrvsEVlJNeTxCWPyy0TyRNTPa++CG9JxN+Ip0pPjNvW7+STSuyVvMrHitGfZQWHAckmDL
PfL1GYce1beBjeNu+3lJA2LXhbjunBh2qBJOxt2cUc8ohMrWZBkU2uHQwfWB3Qxls5m46ZhvvTe/
UydVb+IDSoyQG5ee83eogsetEQyu8qn6tV502Ao1UAbEAUoNFSJr7fFG/XaVE01te4ApTcWsmXlI
vwHaX8YvAOwvuvn59u8CpMFTtkZJDMexdqa1Hz9k9rl68h3joZUlSLh8yld1zqPWOml/pNbvOdFc
ww9C4j0rQkyM1VyM0Y3GJlg0QiZlHLn3PP+F4JAVJO5OMsM/ItvkQQHKdyVZU5p7Kfvlz6Q6ohGY
zqKqbepyVfxAHUD3cIcebCS44fxY71Zc0U3lC+9GSCtbB7E28faXP8SS+VU8g5HM0wWROgMaZwjE
6domSD+zcCzv746BsLucCVyPd6/kefIdBMnwx+5BC9dmRXwefqfSgukwKZoMYC/lYrF+t+xxkptA
Tw2dN6sFgsd4d4a53t6DW8/dCaJ8TcxWm3MAvBTmUTypQbcxSEEOi3dCS40Znj1ZB57+diR5+Y8m
9qDtAg7goCCLHYOAMCeVSHSm3YgstsA+I4J2TVQXMfZQrEOCP+inMxowiFsboQzUJvMdpoSJTWJr
l4RgEKCSC2XOqbb0pH64LqxsX/c6dHB/rQ222D8wWty0ZRKxRyZOr6ACEE4ogNKhdM7D7fbSgIqZ
l/EaWwRrM0C0xpwpTf//RWwzv5k42bUqvVRwvGDGFT1CjHOp8xGlgi/XXVNYlRJiVypZ9IcZLfAI
Efvyxg8sHvssxp+F1zqclXQ5HLrmGadR5frfdyfiQNzP89gG08vAP1Ax3PNximO5yldUz9F75CqW
jO0AdsiMDAqB3e3NJBd7g/gQ6aem30yMp/ef3LUQ3Q+LS0jzVjpeObI8qzr0+vaydnTPy5DweKyj
+/NT4pZHVM5rqghTl1PEY5xDPxHhcUxkErCRfDvN/AshxsCOVXw9/9fGyY8h5Eu+iYzGECRfjSMW
YMkBnrzpeAULq2/ibh/p1FoNfKqYTZ+mm4Uka/lfyQwklMJpPx+1SZaa4macAa55OZ5Tu0SigwKN
XOmb18fzS+3HRmLlcg0ZA2wo+amqUWRGf0bTmNrw38qXkvBlHqUkWkX/LGGE7tEaGeVsK+H6dJH3
1fax4ku6DAJ2tjI1bRRPHksUhzsyvV6Yz6Ppd5fwwv8VuuGvKuRVZBA3sQSFidGge2hwpA5nQl/z
Jbv2sGIwyYfRCkul6KJFFkRSpFC3XSt7ISYeD/d1hZn1ITRQ5JljkDketXhQjrPTCpSHksgM8Nbt
fJUJpqViwbzAijZ9cNXpr2OftB5j+sz5G7VPAphhzNbv3XRsG+A+pm8xk5SGExaN7fzGsBH3gHRK
UNiwUzLGRCFzgVXsEXRXsuFNyoCdUAoMtdC2nAgvgNSxON13aH2eRbUz+q68degSrlM2JNHL7H/3
sacuyGQvSpYlVvP9FKHFYQ03EYzeb1+IrYQ6bUkNI8rwAW/tD+GfuJm6ZEl6aNvtQ7lZj0x/ofAE
Kzh5q3A7hXsYOYLHsw4hoPTnrD2Tl4QmBQO260xyDdWyaicoH+fsFjj4dTe36rAUcb/6Nx+tJwK6
pNXjNA7pRma+Whx35Zw1PkmELPVId0f53Q+7pr5HhmfiVETGHJKVGUMHg0QktO71UjVeTSx5WAtZ
uJbGe15kHgdQ2GWFZPd4bSQYBlF69VBUYVRQf1WMxpuxy9lWHzFB0TYhq15GeB4y2P990XqtNyub
tGxvHCRIBsbHKHA6Hv2935yyPU0/HxEIiJclajqhwdBZuKutGSv873m0otwHboFDA9jPxIsQCahy
hC9+oDFkWfM3GqE/bFsUmGfkpN49fHXHZ+PWFYGe14/5kY8XQEdOFu4sCgM4BDcVCw55QVmVqBwF
eHMCk2uxm5NRhCmmSzlQVdXaNR98SJU+w1PEa4yHq0d068+LeohjRrgSPA7cwsKK2t0wfG8wOYxV
3Em8h2yMZuUZjYE4eKS7eycWN0SobbC7ABWZawaa4X/OtOpuAi0uvsh5Sk7qQ6wcsj7gFLPeZ+nH
2Bd/AWuWfMbBuhvOgXTkq4v8GEjSVS5xNQZCPpIMVVI/2tbJg9QKmxwEqYccScqpmMoaeZeKEUQh
Yr7TZoNb5Xb8c31wEuqt5N4Tq1VVvVStrDdlC3ObNVbgTUFeCJimvtb32dZyXJb1MFvFrnpvTpdw
O9Di5NHrMImJ7LiJKvp9zvcPSsCSqdMVWkaSc4WaonzYJZZbs9nJMVRAcMpTb5qsw3vN9hWTzgm0
LzV+SHn/lYAvKNTYGBU5ZA38V3Nob8Nf7BTcK224Q/pFDeccA2XLhABt1Lr4QHF2PlhU3/BFXLLF
eefqeh3ziSWbka2VYj16Q5g1yjQUjjGQ98fTxuE4n0SKIK3QO8uwfkCBjrtnv1mbn6Ah3HwGB1o4
sPstI7Triz7jej1ap6jpIuqT4eFL5rfa3BJHk15CNxu5XPVQ8s7x8uX29F8IWh1IV/15sEc/tGb9
OkEzOECVKO66xt4jNOPz3g+JLSzro5cyMIc12dXG1o44j8lNNTbEOXFOs8c0N4W5vyYlgcU4+XgG
Ppx3rxPeoHDfhaFRtsGzJqIQKVTVmqIC6EpuTT4nVfg0W76LqyFtlqPcw+iFlZAJ8NdOci/cKhpH
Gf7Q2uP8WhX82hD2pMvLInzSkTUshK4pi44F5DWe0MtYec/KiJ7VDyoFPgGhF7b1GXFkWOy6mZXb
iyOuwUr4RKi6DWN8u/nq3AxZyc+CyLBZc/19ILFqZzonFUE/jA9AxYAUjwHKQQMas80gq0IgC7vB
jGHrKunZlg7h2cL9UN2SdIt+VRhYgUn499pe+n0tc2PfnWpLZX8dUpG8zVkv2HScuiwwKkuShoJ1
P4452mSVDvPC+wNG0EL9ESFqVG2rr9i8J1lCrf93LRhOEsvkhpT1M16qxC+jhgjRs+AJPIWZU9Rj
GndGzVzCyaj9k9GslV++9QnMBOEILqu2XLHgs0yeEnkg6Y6hljxLpyG3Y2Jvp3MtqItTEeLq9qB7
vGlDjRTxz0txgM07MYYrfBR6Mm0Vzo8m6vNDfDEVm+hbRIJvoIHa6YSvsILKpc066TX6/nhR6mrV
rQtRQ8t38FWDqugAtBXnvrdy7rsRoKKAewIO9Bbvfpa6xqw5/18DY4w8hWVIsxdTfILzTSSLHVfe
UCZa3tvVHzPEuT5I7g1xkNy68mhOHLbuMZjVBlS+rW64mzWbyRP/qv5KJU/CkzRPYUgNpsc2VQQ7
yzdjslDrWoy8A6uKOUKXfmXca6YdcPoZ7FgnILx3bNp6/84qFaQSfOUWkW8y1y2I2EbmbIdujneD
7sV2RucNCHkzQ1u5Iu1qH562xAe+CRVPxnqsYrQl5VEAKd/60ew1/9G2IuBn+dWYcl6rfgq5pP4N
eGgkwsrZkE15qKuOJ0fERw10wZPYllgAlLGZ5t3H3CpH/J4e1plUwpy+798iGvVa8cuVi+GnhImV
ivhVrDH6wrfYAhdXRa/KaQcOZ7WionzBz8bilpSnLGxpIyK3++LdOTNqPIgTZqupdj0pIjtySqGp
aANWWx2mfMcgKLZ9rrVb/QAbHX0mQuAsznLhoM8uqrmSWkVwMubdPEQO3mbhVVMWiyC3SSDH/kr8
uSKyJeiSkAFnbN5LkjFFxDvM4TZIl0lUgPFkZ+Er+BQcJzhG38QVe0z+Z4XD0y57dn4tWHGGg4ub
B9WptEGQiveJFFk9s7oEX7WF2MbRSEU9DLWXDi718/iAWXXEnk1Mz+WcrSXHinSWmqszwzmSoT+R
Mjkm3TeWO4uN6D+FhT1b9RzIvEQuE2TmifV6CJyKHJWF3U9hLyrYSSJOgz+3lP+1EtrGwbJQMwe/
5XE/IDC8TRkuw2IhivIp0rvD7+2BtHUQ3ukr/o0UiPTEyxo2mQXqAjteYdsH7l1hnOf6Lg5kGR/e
WeKMTkL/58ogP3+Z9luqbHh4Oad++GENxXQd41xBwsvMXvJjkAzUhJ0U8Tnt0BU4VU+o/gXndxNp
6Zv1NIhhVuCOr3iDf47odx7rnl7wMIZtGZ8+fk9J/3Gruz4Ms+xAv8bZrMV2FmldI9qgaGpUTMi7
BRvv9XLn0HfFuPzmUKQGrxgEPMMdDruNuGzWmcie/imbLQ4LFBfiglUTTgtqZEp/KoXRhlqBmWse
+fJ+0jRWtu4VDVrye0z/LonG7EstVzBYiFmzxZzSARUXuI7zyvIaPojT5xBnj9ia8g4nsUs7jPmm
38ads8+R1PR34LPYHF+h6jsCU8hsecwLId7Z6ZxDP39dP9ywkhjPCxCJbgB8+8B4N/GYprYtl6Uv
FiqS46bUZqgwECV2WB2CiG9ZFy7aEEbFJ2TiDf9FMu4NE7dXGU81PqDyOJwzQfbXmRI+g3qJF4qC
qH3NX5NN70n1QRyO5hpIfXJYjcCTTfWp993/p+C1jMo5Mvhb9qqjpL4PZgX+aWk/LPk716+0OpxG
BItJLm5V2xqqebz5JNHfJweEv9WPlcPZQXLZb6ZPq0JdjNF4aO+TFWX5ZIrd2yxqCnGp1moNsr+S
mtuSlI8ozV5XJ7QXZQrEEG5rK5sMcz6xYCLL1D+N9/ObHF9iLq1layhU68qHKUvaoJwHN1LWvyP8
KxoEcyZEbppDaYuYMUXuvpijeO22bNVtNSLWkewcEKB0Srz3Hdx7K6CtS392gjjB/NmvYlm8BdFT
ogD4EH2mbQhQ3B12s0BeZB4B3fz7H0381cQGxPwOwAB5qJs+608dJ9TU/dFT+ONAQ8rxXBNTdx5W
UKkrPyQnooWAkLuawUHlgrTDkEfJOy7rkVVjzksV5Yav3HpLI+vpwqnheGSs4X4C3TW8tLvHrPJr
jjk1T3hEqXMANYLsFrgO1FklsiMcJXO/yyJkC5GkDWkiAAWWb5vm7qBlICvuD4CNkfLuIma19Wmk
LYZShhb0RIRU18JQibuvPBjcch2bpv7UN7LwR2atllQLXjwfvpDjUqWFKvWnfAnrCoK0LPwVFxbd
UqgPdU7rA5DHZXpflzQ2idHnHoXlU9YnLTya/7H6ogUHA6Tc+BY6RqdIx0p9LmcAfEu1+UFt2VD4
l3TFmJeMmO4AtknWd7aSiDagmEsNEZmVLv2yyztJzPHr2OLe4j+KK2CfEGb9Q+gzecsoCsTslMiv
Gk4zSBIczhLdm1VMCMa/623mT/QRTzj253RhcJoWOj7azatInpu8hl3YXfVHql2MtDYEJ98oWPmQ
6E/AbFCPobaenw5GbI5Z9bCGcLLIsvKUzdzHFWOsMFTV5myGa9Tusa9b8c0cAKve80lsjTTsXIgV
Z78EZZNqnD/DcJ/0uD2ZsTtXwPhOiUtmNkuxu8Kztl8eEramUn+pn6J98cd1ebhQpnkT3dM9iDYv
pkMadzwGgdMFDjXfGrPtGo0DqhHVIZJkWqg4RgunIYeCRaDXzbEHwNHHXo5eIJ9jIDNxSMCUYU2B
VJXYGTceZXq1XbQ40myQdERtXC76sJWckpvlWY5j9BUCG2z2YZoSXGwcGmJAyk3EvNVATr2Fagbs
HNGgIki3ZEPfrrhK0imdZIZsfPn95CyiLudoBZKee3T7YWNqvgf0qk0TolgqHwQm1YDPRHSjOKso
UCxzmaA2fLXl8j34Vr6NzQucWEFe4TAAP3d+lqfK6QQ4yR4jRdHHGwOGr5SP5zNZJ24649y2ETU2
6OK6uuGP4C/f6ywLH8nR/TOwE+xsgBweuRhHL10KRMKhjXFfxAxZJC6/aBG/mdO5ACfAAmr9K/Qb
i89vWHQpmBgG3wbeYZmcB5si+YeE7ikuRXsrjC/stN+6gwLzEwhqRjVIcRsdRpX6TOxSmO29tIX4
1LSK7EFYbHD6QZHXwQON2BVkVPn6qi7skbEjGDAx2teGu6W1owDjMEofBRQ4W+UaWlUvlWPGzTtg
LYWFvOag2Byy+tyaj2/hmthbjANvB40qSCzoqt1FutchHchQRnoBWZx78jd4WtAc8mxJZ49gS29v
34bfr5sEHwy474FE+nnHH1dU70rUNyoDMYfUH4onBxV7ytFA8wRC2L3EKzoLJRe7sTWg8FbAxfE3
igruigac8REZhBALBBHblIpbFUNwL/57+N2qiUxlwsTVOZZF3hleI5Ya333sZ8P3AYsKsiLuGeNJ
dD8+Tax7qmWtYPH/RQjLYD6WpudCKvG8QfjeuhYcOm4VwdzpJxtusg/1VeU+a79kqIivTGqQ4FlA
EBVFeOKeyDouT9xxXG2qXlyZ38ug03TYrSps0rmI4+ggb6+KrXfmhRjR8GfiBzKSA49dodm9QpwA
G4JKa8BBA/Et/s6zuDiy0rtPYAqB5Nf4eTlTJyDPEUhXi6Z0NnjvuvWw8ICnpH+GpRhxJep+tJ7D
2olRtfVLOFFH16xoWEZXX4gb7lf56+Ezx7ty5QiJqh9/GiTwLMxbvEmd5eDsGTdqU109J3Rlk1t4
fOBQ1imhLprGlMkl0aewiywHb2bAxpvU7XqWUh6hnhqe5JqMEbSIOSdLHAzBJaKTtF0dHw8/7h5P
teSc/yISjmG3uwLg1HOaaJ0NQ6yYbB+TcOFqtqD28TXKJXwCvCLwrZ02iEaKoFITCT61Q8Ha020R
WK+n/Y1l2FF1Pao1ICtNPo4pcumPCj8uEi1gfI5YTVbzLwxCRzIG+Osde30RYET/obykmOjuoc3I
Ip3dDHZ2lNE3/Ot3E/JYHnTEMgOO/whyUwIGYiu4MVz8b7S2Y+DIalisBWDsqgVHwml7u8eMmZL8
Ih+2GQTm92hhFEzjn6Vyw6254fNpg01v0BnJWMlfPJVHgpTvOXRiVicbR2t1FnyfqFg+xyfQL+Fz
kQjBqy1HvL1wx/KVBxiOHGH3IghVU3BqJtTAjq3mTX7uxVgY5da3fg53sildoZ2MKBNzNuUEBU52
9evDGmPi9aJuILmbbuw10ifEAW81CZd7RgjKs27o6hswbYrWGKs4xl87q6HD26sjxm8/EhLQZKeB
sLbA4bfzbCTu+EEjn4kQBhVxhG3lIOClKHT9sCnk1cWJL77VpDI0n7LQrWRQ88iXDlgGCKO9OsK5
p4GJEbe0NsoEsWB73ZjMzCDY2/SUsjFRkbay37ZOrAHwq142c2C4ZvXBT5aEZSVHa1kGx1wklC0B
ng4pkk6JnvS7M5hu4YkuPftB+KS3iz8nJhCfXVhr8QsNAA7i1lKukRzLXaIHx7goBaXQ/UVarSA9
IrU1cJda3W6uBvN6lRvbsEGSi1TgXYA2ak2d6IOCovKd6ooJcfjuaqCOZa1tN6awJGU27uQY2gW2
Xy26N6gwoLFdN9LRfCMzCsJqQmJfFVt09V7Dss7JK9CponY+zLEJMOkHwO8hpTkVeb4TZS8wPTOf
CBeJFBdhKcVKp6WOvuSBWcRAQ6ySUZThtuXzQihAPn0f2xJ9gOe800tyH+n7MwLhXz/Mo2UO1EWj
k939uwl+o/TONqLQtK5us6ZH2x4KXtN+lpdsI2XUzDL934Vk5B4fLAjY52AIj9vJjnGYl6RwvsdD
YGsurbWh6dzdkm7cnrihqyQLNvogIWej8KI1mmt1Nnc9XpRPKcGtyn4ybDuHjeDEORtDWPR69q5h
Am51eRtauZzq1wA17aegYQo7Pi6P3P8vj1hkAWsxtDOtZyo5KHL897lktxu4lE52/RSWLS71KdEm
05FGZFYwgSrXnIwHl2tYPwYYUuR5fOzZjjdcUwZdxFnbf08rqmvu/ezt9W3DStK1gK0sxcjFNYNu
e/gg5H8cpErhlUr4sWrEACk+A5QcWn1xlgn48J6OSekUi03DieEkfFKgUv7e8Zb0UQGN5DOhh8TZ
aviV8ZkjDS6geUeEO2fQWx1uA6UWcAOXq4fGoIdjQlSRqN+MJz1L2L+3Z/gJzujjiuCE53oxXmEG
BGfRffVYxZ42+TWZIW4s5qBSdYDjxNMkqy/ttzwTBeJUjq7jeSaXS12va09Mx/QI+mudhZFKNIb9
er9P8uE2WMFxTetzwOx91Cm6Lm7l+IzJaTO2NHvRxMaxWIwyWoZkMUjFxgs8NCR0bBcw883xmVUv
lwGncLN2M2B9PF5T/Mvg8CDIE3qKxyqAlakQ3HSB8inDF13isG+C6HbP3MwxOc6yHfObQK6pdX/q
okXqHXXWmPqbjrDV1qQ6wcUcBbVwqcHlEvR6/Jck08so6Bx5bJlZHTqgkJT0PMsw4l89mJ9LNoou
TBvrmukcADUGGG0T+kd/U6C2zZ6dQODEaE7M+JNRuimVIauuHsaubEww8R32M3X1NC2qd9rRed5O
M3U08VahFwarEhrEISNDK8J95e7R2OGdEz8tpbIl6+88ctu7t0aos4JQhXUUVt2xB9O6YoJQUg9Y
eXH3hkocX/Vll+UOG/fqhZ9tkjMsl/meJuXiUFGHILQb5uSs4w2ESVFe4ZVs/mbEdUy6/H2UPIbg
miCUsQJoCLpFbdTnAVyrjSs3iQU8tqicX6D3rDvgixuBnSyUpDwh63LlfKrBNVgF6INYmyV7WHvx
7jmEzRnAnzKW9Vj3SOHjCBPtStIuwZx/Swjs/80S2n0dUopwjrxUSytv6AlgOSqQWR+W6zh8PhJ6
Ib4af4v3J/ZgY3nv4pdT4tNylp2FbS5xcB//dwVyD0R5zAcxGNQ9AjcN0sfl7IJ8N7edLLeQS4i4
eIpYSlGal0+H9w4KwCcKFHgyzZA7Df6ZyupKT+aUHSk4BuyjI/XvwjOmDw7JeG/Ac9drhkXbehQM
kf0MJtvbIntB/Oesrv/QduezXtWS0b09MPQbccEe772kODXQsYRMNMJy7Mi7sDlzvOCz8z1/MGhl
LzArLz4D9y+IANwfjPDSzemth3LjEHaiuOUJU0EaOrcEXXRZANWpRzJyKd6jqKEJsksQE185LWzg
4WaP+3s5lmyo2M9vkxa+xsHXuyHTcd0c3yxrUhvkPZeA2CpM+dqUXqVRnM5yKbMVkBdFl0zAJV4t
LOpOhtc0i8lz9Z2fYtEqsF7VlHLvPGHqHRaRCNgGQuF6DbfHzEUSEq0Sb15qObWXvu0dKQsBQrbK
2GkvCRTRw+xnihWtXd8U2YA1eYt+rQDNym3x70Dpqi+Qo7Q5sDYale7o8Za/00m3d/LWM8im5k9m
m3OhyLjx3gPwe6jUmDqhcDOhJrspvIxh/jeLp5EEQrchNv6DCuu5ao6gg81REF/Dh4d8TBo0FrNC
N/PjNaH953QKdAl5jWhnMfmHxY8G74kQgIG33LsphCLGAucIGrFRwr3YNBRNNa9/p+l5SGnNbdzh
ssdSQQNP2xbO6uX9w2VCKzIx5iBufA5iG10siv3knonGa8LoYvEfCRAgQjmhTJa0J2Ks26Fa6pAZ
dTfrxa+D7PiFvETtqTNZR5LNDg1plfkWVjGkQpyjHZlgM4mc6JZfcAWhU1lGwLIb1SPMGnOrBxvH
PNqQ4j54Eb2m0ueXp0iT0wW/rWaduPNwwKpXARvUIUkW70n2J05m/FLOHdWRc0x2mUK3d0EGZUx2
nBFiNavvkVIj/91ZGOdzive+THPa4Vyjgnxj6E/PxlnNy1pZjE7iUKMC01qOXBWcxzsqFnz1orj3
cZ2taSAW5V/7WRvHqtYX1YcmaPewtGZSLFmQrowGna7Hq3pKjeX5mK/vjFYwPV4z6W8YppQ83gRr
sWTQY1bjxmOzDtGCnpaR+M5dUG4Kh3da143KULQonX7nb3bsbe/qm7jZ+3xRm/PoV2ezL6z/Rjq5
25BGUn7HRmHEgpcd0B1zsa8OSYxaEXWKYjcqLp/Ba6NQYR1GwIJFe0kibTkhIQqwO9pvl8sTtY0Y
jlvnUvJa3aD7ynJAhLPaf2qiif2oj7ZDAre2hH3UG9t91/TLLbb/DsitZ8azdOUa1kThmzMips11
FMuJCDflxgxdqryjMEgAUFrcOJSzfUp3K8eibyQfA/Zu4V1gkqGqK0+gzW3EmPElX9qipy6xpxo/
lymw2Xtqg1EOwHt+/OLsqEzjEA14B+fZLNiIjDJw2ebWN9qDEJ7tr1RKi3nTr1MhaITvIYkRAjy0
L5JieMFbyY1+ACm6lVIBKY1euLv5IIAtdwD4p1qlctN1A3wGD6r5Q3RicB/K7WrxcLUUmTlnt9aj
Ec1ImK07ULxjX9zDkKD+LsVav3Tc/1oYKEVQxIdeK6iQNUNNvSvQGHNcmKIv16YXS5V4xbqRe8R1
t666oK4UJHLNxTaqryFEuSP476tPQ0gUcFrDZUHCeIpAWOPiz54oS4kvW4RiuLaTIpbWC+MKxGE7
ZJEn1U/j66SkqeEVsKDBI5uj53Kv+Ga32j+1W/OLs+goIufff+HCK7cmbWofbNZYl3sDCxDia3g6
8qhb0kwE8YsWTlx3bAUMXEdNVHwDwmVQvXfyao9aHpgTSO3pqQrIjxIU8Cc1dtGaUGuJ0TLh+te/
Z9kohzBNSP6z/MEg9+0eKnJg7paI4kBvhLG+FQuCzR8MdU3kLcZDDCDLoPKl24Sip+N59oXbVBwr
+aexVvW2f1fEAJ3Ac2NrsZXNGu3PwszMjca9bKf8riw4cHxn1+dRqxrAgvrU3E/JVzrz13Qw3Yfw
uetWOvdOYed0s3Itlk5ve/Wsacc9m+R6GzXKJ1ZvngVSOxgEGv/SKa8UHj7WyFv4pRzkPvlAMHfn
A/f6m+EZeUbQdWBvyUcrkFWH/iobpJP7c5ZlbTj5d5UOolXGxaEZGvLy94PZMmLKeDI4JHs6ieuO
10pdlaCLTNbs0MBPcvCxns06IOTOsHRjPSgbK6Dm3ByP/sW002QnHHcU+ribUI8ARsQsXt2dusTz
+1UGhldMJJRg9qXnsQZrlgZLRuke0GVyh1s3gKAZiVFuC/ZQve7cilE8hm1Po6/w1pEpHk7vboX6
fHpr1Ra22IV+UIMinGlT7uXoEBy8KCPf7VO2N7/swkgnOnG9M8pG40G7PZp0lJt4RswEKGZ4Fo88
3gfcZaP1KGWR0JCcBKST49n28VvAvGLz2GfJGlmeYEBGCuzJE12M8NHdhxNL10HwT7uMzbaIMB6i
l7/qNyhT30ryMCQ4jwJIrCRDAW9udXIvdMCFQCn+/NTz4s3eDhyopuhkAjm+6P1IT1z0l1huLXcL
4gJLQyZr32UeKIdRlF7KSWoYViZqJ99vqbEck/NWGmiM1U4eFGt1w5F1ZX4oHlG2laZ1EeoS8amQ
P6/lCnr9x+P5AQTwpdMTGK83jRpT3d/BfG+HqCoQVcY3gup/NyeLmOwi5/4srD/GCt2r7xSPoMWN
X8PWALx+BqqnrCMTpb5GXkS3lBVTsEzp4xLAeUS53ggfjqw/Pt4oN9bqiNy2mBitQLNdkU87UHV1
oDGUrXJVIeVYXl/uhlQCjVLPLBuXXk8TW8r8fE60Nc641QhngM63k2XI9O1eiQiBXLEYPnnbuppu
H2TRggG6LBJ0cgC1ANHHyNt1xcoFWxK5uNxohCgMZkCjSYLVjZFqnhrlUwoSpMzT4WXJDor7fnh6
FZmAMnbzKVvQQzxMNf6gnZKxGJL3JBFUsCNdsFjtt8s8YyR2nuEcxA107E5Cx23sXLM5QE1r+GLg
uOrCs1zkpiygvXYi4kjNPEnXp5QW7G/I4rWMGrjD3y6whJr2TdAb+GhB8Zlsm6ROHylGXHvtId99
MyPujRGCRCg93ncEAOTDmF2fHACdPmfhTEmaEiBmvGHvvVLczaspypVzt9iDexbik678zDVudNXn
6QZHuqoPM/1oqa0XO6MuUKQ6yw9qC/BCs+Vl7p1Jwachtozp8A21+mVppY2wcbVIrBedpCpbhoDE
3d6R/vLZXzz9uGVOJeE3tGjarO/rXOJThy7ZrsVRWI7xaO3451Bq0Ej4EQlQ/nrUH9SOX5T7tfbw
iN2Qa9BciUbjp3CkOWA46Ohl3pOKflxcxE26gdorwyVdDel/PAFewx7BpHoHQSDZxoFJWOLwPcLw
MfjkVs3JLNv93PTrslhMZklK7mwvTXdEhUxBUvqZ+cbWFqq6UDNH7o7tnGS8Vi+JEWlTySCRVNtp
OFBIzCUxUPcYYIshTzL5Fo1BKDQJCYKQw73GROfyXBa8iXwofQ4NCKKIrYkll6e5QLGrF4qqK9X+
2xbjPy8BvA893OnM7gWREkbocShctQCG21Lx64ib1QE+NxagqDHlCFvP+oerhcmEDni9OJTsRVIc
6Vy947lnvMeM46m0dIJOpl0Tas8AU62DmxgAmZqO1vHJ0dmORYvlJvImt1zitL9uc+2R2UXu4Gv6
WNTh2VPhMS6ihrjNMaAPDmdRJAclx6qWKDDvXSsyCSLow/wnHaJb/EVzh8jhxFKoX4oASw4l/Flc
QHL8DPaFRfqX4KXs9thTToNH3brxo9cKBLNqG7tWDGBRKplrJLAvsKZlE2tdcO0rvKAhrzqNDoJ/
tAVFuSR3+sj9c/TZitfrgNmVGpRUr9C2sYqRP+JDPvGo088io9+/A5WB6/PTDeCihOyhdn0kiMBr
AVv8PkTnIu+clLxq4fjttZq0AlZcVAS1oGKZThHq4+mv6X5KW7JMy8UZ/5lvnPhC8wLZkCrsjyag
lSyitBpzk0Se6WLDtcXUXfsq0NBbzVNLyUGD0Oej/GsYjNyOZPwCthhSVqo45Q9+wfxX43E37MGO
2MzUEGW7lOtN+yBxGb5LWDnCpY4pXL9ByTT3XqVgpmmxawhUTAqwWJ6lQsDREhER+fAZv/XBYUQN
upf//aTrWK9hhttNPKPQuuW1kVE9lAsSFxAZicRuXErvy67P8pAjJ3ssVvtI52k46g5qe0Duz9Kd
2/5l9kofFGFQv05wb7fDMqey7tpeNC5cXS2e3R8apWb+veNldz6Co/mzLs6bbPnvrUmjnOIv67lw
BdvJxQNF4wfc50DWRUMnb0OWcefbWK8rdmowoLaGbTfVyeP0o10mIxpKnB2BURlP31b0y4EZXQ0V
4vlbVhk/PLmdEVXhNowJblURQTh+QHFE56izJoFdbsGAa7hGdqHKaf+kX6gF/Pfa7/wJnNqOio4M
7DnKRwg3aolzandrPCA6ijvzvTH1jj9hR6wFBtaNbzFGovnZLcIh1+x85d1HH6VziG5V0Ourd3Wl
XCKOUj9lClOoA5MkAmqNneiJ6B+p5nA+aSOsU4JX3Y6cpnuoJr3VAqSJ2Lb7x0Tf6RkJ78wOG4x8
bCRHBDLor1jooKV8PgeM/qEPc+UtDxCuJWdL6uDb9hWn1T5FMlr1LQ2mmhbmoHH4nlrBo9jYXpE+
Kuo/ZeEKv3eTQa6dhXM1AmPFwqZ2QFgpeB8hC7cK0vj7n8DBAQKtIOHREpXE9ugPJEsFd9g4UgIg
VLLxjbmtbde3R/4orAwTYQcl39mJfayDMsV7R6l/BqSBdjdCSQegLajvWTJkjpjnCOktpfyMEUzG
7xdjWn3j8C6dbCqfr0PLnoEbg/keHnM50KQCblxI+DSXrzAObMdxLYwKRH2b2QKHf6IAy+PTmClc
UO9zAXNdiwSRzJvGcusx8bSGSjm8iOCvyzqjSBkg221og8pfLrFzseFd6XL9GGw3m/dY05vpJMeb
CCFv7+CowX1QagrC7RE0s244oCdyP3d4tgEPIGtTQPGBOBAxgPGKeuELAIDV/GJ+0vksAUU4kLv9
H5OgrXO7omBytQujHxPMsIeInczNdzDfUoqRw8y7wNEgExTNXBaGjlatQyysD1OgvqJumre9fjD1
gc3kpHAIPzvafMB5FzxoJFtErE3ciqDSakqfA9ruEa9I4a5VUO6UuluA8JXyWqZjRyb5CmFRgLki
hzap5H+ZN49IBk1+Izu3Zl7vJBRgTDob48LkpU0AP+W5Y3BqLkkePRuP76//T4RD8ngRITLgCal/
lLiAJ1/4sV3gzWjL5mPWkn9DR7mKKky7mkRsk5Qvl4UOytgOS54TlXccEMowaLw4EvTeCIib0rdN
XhliOqMWgq00acr6crRo+mxqx8TAi7zAiVg8jQjbQFobhHMbkom819dNd6XjXPPknnvszKccRSvZ
AEL1ZeHR5BwuuaSJw2okO2dvQ5gFxwbNXpb8ltPgJnfNJFcpMMNtXasS/2ZVIvcj5vOObhb+USiq
heD2U0BLlSuDz60zjA0pHnB3h8PLSU3E27d4wwyCZVrMG6mNpBygOyoyKqoYZ/GOgvAREp29J65a
OvpLOpMCzxnPIJkeBIDjQZgrbccYYh1GgKkgBEf6Of13TCTa3mp9B8QVclJOuePurTRAcV6EwLIN
fOl50UVU8HuwF4wsCvXJfqdJIyudMn/+yMW1BPdQRkdKQMiOezWgr9N6XNLT2VmPNFy0e7geYShp
3wR5sM8v/gmRm/QBOCVwU5ypAlyYD1p4w1E4NjZXQsT3Z1TajOKsDzZ7EYyJDK9LT/AHUYTu6+XL
JO0fOD0hrH6d7vxNgBqPPreAdvMypTzrT68H88UuRlHR/TX+n9MmN1W3j3XZzxavhCU79yA+lTXK
aElAKxeUriYAEahEagpoCe6tMhyQBe266Y4cORjRz1UuVIvsFKZNGfAleZ0CSzA6iA8MCdPb0d36
8XPy4mddmkMvhCio6Ampj+TW0HPrciqx2iQxWREDREWDMo/CUXas1CwmDUn6XpZ2EZMm7XZAzIXf
84kHh5jk4AFYS2W0yByacKZASM20/obPSL79zjHdAbDwgysAjJNgTUkmILaXvMJRnSJ7ODi6iQAr
c3YAF1XML6Cshwu6f/uQEa0Fv+5AelEYZQ7tcBP3retG99rSHLU8FLn/7LjfxOKrLI2o2NCwi/O5
iQgZax3M7H/LT93IvA6UIYiTZLSggSdGJYwoPZ/gscaju69A+eT7ZWf5EDkmpx0q/Rkt+WCuSFcn
1CIkdm6PkVqaJ3WsYvuY2z46GFvMGEpAeI1oA12Xtm8CVP3MOtnAUenx/pMxb5qalH8OH88H4PuJ
sNd9lt+UN6L6nt8kpZOP5Ccpa8dZohENOdFuLxsIu17PssIJOZ2WtO94EUpJUdjoRtT6qb8D/7zI
BmT4TJUqqhnTCVRZR+gl5ULVOJ1DekGbOx7YwNLQpro1+CYIM+NY8pc/QHKYPpjxwT1vkj2W3fav
tokOHJDu9wkfzye1fJbYQQvzapz4+cgWt3IwKpOTpdLpngJDgco/2wNsEujDDk/1GsVSelFrE1yO
Peh2+DscCekeEuQr2FhkUNmyRApwBoSb17b3V1FVwRHfSC/1eSrjtARsqy9JgivU0Zog3fuGqOj/
J7cMGRuEMKX2KCVEhROA7F/WDQSW5nmwzTsrvfwWWRN04kfXG0I3daQNsLX6tMA9oFEGgtzBHz9S
9m7rnN82jla9oTPYyfnwTG8LqtHpVYgYW2kl8aF9RV5yns2LEPbPhuOR6Zcyzo23itii5fIUK+z/
MvluN4EBXmqwZDjtgyUaSxXUE7lz2+dWMnEV3hyhJbnJjpigsZ+dXjTwNqrbXFgI8PVJoa0nl7/+
wRb7wDTu6AeznbdKYjRhhabSWZaSfe5zOF6wd39s/75xneUdwtmvvooA7RrFP5xfyXsZ3YwMtujG
VFG5fEaQxIs3uQTmomgmUqsw96jpP6SWtC/jHUpyFYXupXKNkc4cmxLk/PR3L/SBmdJ0PyYYhx6+
kTZFUwxIBzykUwyc5YFnPFsG+EE5tmyfKHDFqWlanwRBHVjwjnPwIEhrKxsXtHGrELWVfQIugPsZ
mONg6aMiJ/4Sx9aBij2yJnow7YMHqAiJmlQ5f/l8CONzNVlJqyS6UWEVMdce84R+0inGfdX9CBBV
POUVkGshRwXh9S3lyicu1asapHdJDtFpoO9dWzyKUy4TONMSmRti/z5d2HCzhcLM+Vdidgn0XW3h
5phd6qDozECY1OkB9lElgmLxV24YHzJ7nt0/OLSgkbCDDW9r/S1+uZZblbFFTxbesGGX5aHD76rT
PwjifG+6Ab2tiVhpAfjrmqZ1acf6LHpgpXkRaV880bzF/xhVU4JVIWugvjWoLnXQNoembTS1ZjlI
b3QsoZxW59mhSfN2bnbOeF5ubGeE2lyICSnkOWHvMGolCYfUaatpikZcCsRPSPpE2qZId9EGpnp7
YQ8Sikv07zYxc6nKhemFcThc3Q/WVdxAt1G3uU8Z/Ej3QJqfT/BLwc8UQmN4uftrSB8u/04pui/u
7GT4E+HtkB9yqKx9jv9X+rBHQiuUAHXCCY0bKn0IV8hqorLM8RB/rkl8muXfMamlOoSsQTmvQx1u
2OK3SQB7njFrUNt4iLptIxUsYncENu2Kv/n5pZbahxQQfYQ12JbsUcQfqkfvCITz/vWf6AKDUlCg
7b+WusCob92FDSQGF3OjYs4YQCTyYLuIkxSkvDw38eEU5wQenvvDNt4xak8Sn6xhvkWgiNpe5+VI
udfEIfEmJABOnywQ2fGSspJFu2ZcCE9u3RzShmcmAY4ZXdGBhlhagY3RYmpAvxGh0ivjFVBIE2dw
KFnob01SCoHjvKNs6hkidRJq8sE3KxFUxlUAN4LfI55zHotrMGyN5qhVZyYEa3f59dLUIX1+im8M
IKGv0WOkYEvNeAbFOXp7ic6DO1zm5jWP6HIbG+IeXszR7yH1cq/fNHIHGlaQ/GzaXjQcw8PGN+es
XyBtB+jQjSZh5bjeCW16DvTQZZdKRF5rH72ppBXoPKlt5sQbtIhIQYgENS3V3oLgvyCIqwe5G68t
+VR4G+Evhyd0qZ6MZS1bRZzwqJKZx3Fxqqb0crdNwZjKI2ANXqmLNyDyYz1lrzs7ZgjxavaoXdry
z9B0D1HyaoC1wV8mn+dgZWuKwU+2izId75kFR7+z/tk1VvGtMFvHSQ1YfUfHK7t/NIK/5BLxt2e6
pVAmfcsV1dyoOvm4d2lz0YXTUNf/VsQZQ8FaWPZryLXKYl1XFUPAX4JyhwVTPqZYNEIuMZsAErCX
hliz/+ppUXR+2rcFBY644rfXQDbWDk8vokXcPipyop6RlDVAJZOaaw0PBvGTsgmivDEAIHAqf2ww
nvog7poR5yX/6yqy7FCI1+/DYv3xLq1WA5hMXs+BJVLbiJ0B47qAv2K8POROSKMgV8rCPykHBOEE
LXeqicrC5SHRBCOeote8idmm5WCVe2zEE/d0QpANVLXXsEza5tSrgprHWMtqOHQB2zcKXZVZg7Cc
oqED0FBorDNifxvo8V4B913xknz1BNbN475Jnu6CtcxWl1pLZu4caqdwXXlkhJ7lLRg8A5cPckHH
FeaPzdOw1kpucXtS4Yd6KKHfyaV/jt0CCliTp7PHjmjI7z8hS5aYttmu4COfICIZLSU1u3kvS8LV
5sO7/oIz1YpgyppXvwaZVncdPgI+rtHzcGxVf4XiCV11wachh8cWfJTKWEbS1JHpzXEY/Acot5oL
cV9B4Q0YnSmFVbDe9gRHehHyoG4VCQp+S4pE1RguX4y5frIZDYu64Y0oPwbO2pwUkFLwdrEULwKG
sI5wKK7QdJbVrctfj2xt8ijORlBoxp85NlONDzX3P0gOMiEuhkuEfMs6tlJVvyCVgTInc1EUeelT
pkXMWvEyseGCYwPIfuJOPQaCvROfmkQZ2IUhl31zyxG+Xs2Z/tE9ta5x0KJMV6DBDeicigXNcFr5
MMj+iCI5sXLHJB4hk/rMXBNMHxqaOad8WD21USPiIKgpdpjjaZ7UeI5zvFMypXZFHLA5ug8GeabZ
PhAiurQ7Yn/dDj2wcVpoTOfSkVEB16RMQKPG5E3MqssotyNBke8G24aLJnGkgPWnwEbMbD8ZCbXy
yPLfMTaVcB3UO0c1FwbNaAMXJnzoIqk6uWBPbKonI0lkaAMDX0tV+v9DxZONWxjSZas0HToHmxrt
JvAsZqv79y5u1WB007fC8n1qTMDL6rQZ5tXc3IpcHeLsvlBLtJYUr0TKtwRnE6gzi1+L3PnADg/r
3LVcPtzMprsPeZB4oNV5yALFO2yP0h7MhfKdeScssGbCf7ghFd79pGRGEyDCmOs5lSIvYm11fxNy
aFR6sVC+9CM2O8sWR3D8BtWg4T7X0DWTF1ICMQHy0PUaUao+O+WuPgUHyzFjewwvFLHuPvz7rfdl
3s2kHcbBNFXlLcJgXDxX9exIP+mmh1Td15gGNyLzQuBn5LVVsSJ+Rfk2AP3QoktsxSHoflHnMUZy
FRloMidYoknyCiK4f9QQlATJOEjMKWKmt7myURQ6T4nwTFuUdDjQI/bpUvwgMc7DBuLvTSAHCrqA
KJQD6XdjhK3XgGD98xEunfMpGt/oIibu0tmWhRj+bDZ5+P4fxyZ6zoXjCf9WOGsIRxvyZmpt5/rr
0Lcq+gsiVT54gjrBsupFD+mMt5ZiddGFH/lknRIZ1uS/qDy1EA0YGBRyp4ET3tOhVDMZbmGU3scW
rb857lnQqdtThoPlWdD22fTMf+wBFF8AX5HYJVwNDOdIZEZ3+BToeC8u52hX47G3z2CVXreIy7z2
0/2DyJUbkkEwfYI3UQM1c091466S+GcRffhSOA/fQJk8gksKYhfLtRRyOdRwYEwqbC9PTZrxh8aU
9zyLL5vlTc7U0pZSCUdYX2dQkKYfRHCGkB7ODSpo3r+qYp8sQj85QseDvrTiQObe9Mq53+Bfc1cc
amXb25G7e3Ytv+X7+8w8FumIo/m0y8DqbR+3osoK++IljLlpnieOfpP7gh5rN8ne4oJnNaWlS9AG
9HUPupU3us43ttIrvyZPkpn8jC+8PYMNMdecfpZxjcUORGltr3Bu7O7se2qMn7IWeT0zdH3yoCZ3
LBWk8G3DKUYDB2OoWDgfqq2SPPoFlkkxWnt5UITfpYKeduhJYPnHrCSAfHItk345nKr6EefZyN3C
sGnbO1h4DNUqcVr16atgQd+iu1xqGAZ5tG6xgqPpyXMhb5Wb4LD8JbUG7o03bGZmdtxY5VKHwqCA
Yz3UD51xoEWqX4kyteJoB239DrCjrL4NxubNHO4uyJGVHou+HrJysAZvdR5l9ddFxtDyGDN5Cs2j
CELiIExNcpCwpozZNQJRiJcJcet2FAiY2iiNBY34OLi7DUIdNwGqYj0fWm1JXa5D6Osb+/EeCKHH
q3EoZXWOGMnVKrze7encA5g1PyE/dUXwhexWBR1fEZplbfQYtzNEyY3oN0JTbHxS9Kxk5/E6gRKV
0mosdquksb4bqNEEVO4fnwKlWX7fZs+MiRGF8Qsx+LZTuqeKdcD7yl8EL6zhpMSE7fY/azNCs9mG
XKidG4qaoeVL8W92PZePgY3FUSvlSB5dPsr52rdOs8zaA99CGd6NaVwPmkg+aoFRmPhyHAy5xqJO
l4eVcLHJpP0YHuc0qrvhO5k+MpmIpRYl+U788u9SrWCi+roFh2ys9snbUzPNOzeKWRpU8uSTTqY4
3cy6BTMxEz7kla5nWlIZMvcswmGDueKuQzxeY+ZMp0VdlCH5py0dFtarw/FExGESHpjf0HZvTA2n
w+z7RJXvxH+n4KjX/Jes8rfHJ8MQ3ZENP8A3+BwmQNQJHsId2hBZ3Y8loN0PORlWoLSx3+rJukAZ
sPnXeyeVcBNCQUwA57mdFc2/2MQOtqTKemYVENcdsy9V1acBg/IJEwdG6mLWxuljUm4woytf9THq
/DLVDKWquRXJwGZfoiCk0kOCzAILKWgwPtnJ4He5yirpu//EvPlrDBrcJOiP4D47kSDRJh1Qn5+j
AcWSNKqhuPttWrbmVkTs5XsrCpwdOg3WIHfEtxWLR3BzJNiI2BK8wkXmpbCYvlfaXqkGXL2dGyN+
lJb/NczH1B2wxzKOdp/sa2UIj8FTfbne+t0mz6y16DMbC5oKxP1yw9AAoh/G4K5OpbaE06n0x0UV
Vex470sDCbzW1hyIM7eyJfVN6Y/Wc7h3pnXADIeUWdVJTptXLiG9l6QVE7sV2ODCuJZpFR8OYDse
QtZ0my0pIzc88DQYKnmEwIbAQQVkpwFaUH8IM9/udC8wEpgYcq2StY0EllzciE1kU7SzdzMl50Tf
jGibocQVsrGDKAqG5sKuk0WlSMxCbH7a0teH7vEhcwrm47lB/Tl0tjJnoG9jFlleqCjsqo0YHNUx
gND+kUwuIUynGqAmbYxSB7/Bw8W6TuvuzyiRoBgeM5cvSFN7OB9heZO5w5lRk44YUT17EoKPAewK
tZrtZIh0OLYeDTvJQwpor8bYcsolAT9/Z78LDF5+keEBQqA5dnSjsyt7SIYzd5GflYojfC591GA1
Fi5sRDezbxF2FDkeFqbGOArn9nLHLuAzs88Fj5IQJj2Pe+P3OpM7jo5M1TBEz/6fnr+NW+cIaHmq
nvXamkWKFnbRqFhOV5CPg/hSqBMOW6L5oCh6i6fcKF/KdShmSViUvcfyawGYDCG0gjYlymga7o3i
1Zf0DiFt2SmZDxoh6Dof3rpI7Uldiajo1IT990illSe7UrzduZCKqDDnICTSlumOKhXPer8yvs3U
fLUscHh8PDPhH+8vbJrzuROmTE+of3cMDruz3XARVeV6WNAQtFCRLe41LT5CT0cQEc8ZP93JXQ0M
cfnYBCRhicbMZf3alHowS/d5GyGM4nWUOqS1UgKWGvVFG78bAJ8KQCeubeiO9SQDODasABEe8yyJ
hctbL4QufxwAZTlnD5zojWZmLobxRo+jsAkWEASLmXJCrF6f8mbb/wyKXhHG0jKYZaj2WKo7Fe0j
1Q6DeR/ZR2pIWlFLFHu9NHoWi33AN+gKWb6PLwcj+7HWeZfgd1bhaQiJ
`protect end_protected
