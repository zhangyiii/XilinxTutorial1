`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
d5VJXu82JfSwswDjhvbEU9He9tQ5/1Rw+4/2nB84LUuT0wfekcnbAADJNd0/JtXdeaCUlOw7Zwks
Bp1VvQeB3w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T1a12gH9+o/WCd/uq6lAozrIbwFwnflilDyEA/rZKRAxvRmKOSqBXtjVpxVSoEgX9El2BLPK+36k
Vd8y/iFx5HcwlteYeuYuGTvgQerRA9ycH4Qwt9s5DC83MaSGod9ecMMI8PPrmdJ+hCOX8sXwEsN9
IHAKBa7h08XDRsgW0os=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZE3CBd8eugZohbo93EvXvQkUxCnosHfYT2eG0uuvFgW4E1aUdxFin2hcHpeAodvxBTyPhYz4Lsqw
3nsUxnz9hTb8Lhj5XnlqKx2mVFP8Z35n8lJk21C09QHBGoSukklDPI8dbQUv/KxN+k1qsLBHfCBA
FWz2UAwKlgCaoOPe87s5MUwwDM1/P/D4+XgEQCRDz/7JDN7p8ZFVtltMEx51xjJOCvfGoEeTzG2k
908lkYgt+B4pvwsuFOHwC28xicC9lqwuIR+OiqTI+hvqIl3tijnK9dhEHXmlIo9PqdVp3p9K5niF
C0wKwI1gK4zk+Z+Qv31AV2g5KDXjXxSpUgHlpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1K/c2Exmx3hO4tktdfNX/hsUCqBDw6bH/vDRPja11f/SX2mhefMgy+yYp/XXIVeJlyTPI7AwLQ+m
jPsm9qUsxInkPzY00BDkxz+XjPmDvPZhWK1LaTfp3S2KuDInJ2AYP1AwgClVQtpRFpipBFYqQeNS
QrfV5V8iPYsCh6rtCZ0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z2R2Fz5uoP9gCKKJ4H8ByaZdL0II83JUVbmmEiqboGhJOssYqqghHZS4Xla1DO6PE/W7lUbFZBMN
taobe7WZ5vLL3z9KT5znQ5u/8vqZfQZBnNTCM9ij+NRl3PRmkUPrtcd6xURukGspBspXFvJDNTq6
HoC8rJF2dAK3E2hXtQ2qzFXYx2JspRBZw2ARE4ENjzYZSYK5AhF3nV89pEvyjDlChnkSNr7Ec2sz
zSK49rQXLtbokqxvvzCHRCEs+NoMqKlklN93OyjJFAIzYffS6GiGtNeycU755Cv+/fAQynybNWn5
4vdHnb+JcudvHzAJFK7/azTzKOJrOSm9uJYTZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9024)
`protect data_block
mvi3i3MBI7n8zvuunOT1BL4eDGhQlMnzDOzVrYI8XHOS3ZoKFTTDP4UmKkCCDyXvukS63/BOGJv3
NoJdfMFYhDx7pjz50AatTRm5dOIAKktHZJVnSGt5h4GNaEO2RZrMb78Xxh3U1zVrxlZ3qI2EnHdF
J6WRO15EzLY/6cuKO5Kv8UeekAl/ckD2I4ewipiajYWKZO3uf8k/Rh1mOKwYOfnYldGTejGDolVs
dAkFAfrWoFa5NH/hK0UfaK5r+ImOHpNiKgNwhCpYZss4JIw5iG8FkGHdaqxmX1rlDFXe39WkxKir
MY17LQX/R7LlQuKgCjJ5JAvcFinc3JBA2T1QO+ZPuEX4zKiev65FhCWHKtJ0J0MuTk3n3krtYxe2
CKPBduPyVAzhHDUgxleRzfcBeWIjPpAEe2EvJQ4P6LNI0DIhHXTGJa/lZPGuuWVzfoEkR/iDX3+O
piInkMC0XtYsn6PhdXjH55FW5JFDIdxhUKDtIAzUsnFIbjm2VOLWjDSU3iaMP1lNTdvFPbTcZsFv
ZgBt8D6HikPuCjSviuh6qnTqYY67dza7FvYlUL2uhm3UhQL15HtLASQPuOleyqsG1Vw5Zw2MfuuH
k2+FG/JAAte/n2gQt6vQOuOVZDy/RKZrxKtw0PHl4JMi8T4K1te5cvpsOz7JtzzNMhtx4IGqYNxk
YUnAobChi5jsFN+NBalH2ImOiiEH5RxYkGqVwderIUKArCAdnLBb5qjU1TSR5KA/4qIZRPHCfKvD
UPF7cSAYNEN5Vl6ts4N6KLVKYjrOPzyPkHLtxT6uQ6jg+vg40K7q+teNSAeiy58/QY4P3Ed8aoSg
U9FQx3/VHFxinuM3/VlITTFUf1VgKTzv/N3f4sZFC14mEwjGMExpnVCBVoJw02MpPJw0/687N4yB
u7pNOhO50hSjk4EBbukK6U/9tUfKMR85QooRcc24c7CrRy7mb76yppiwctYsGzw2/G6EuSsmj4jm
hKL+UMuMJOxSI6xPUs6hVmHZ+DlVVxRumpWET3z43gDf9Ct70tKTyGSg/RFBTNnqZdz+QXZTxueE
Esli/TTIwqYDUwiTr8yzyNY8SDyb9h6N586UdOZeIdrn7MLl472QFIr/hMN9BSDdUVtSDS6i/P+n
oksL+L7Hc/uHElKdJyeo1wkVytMYCBKItRAafq/sGXO66uTKI97nt5veGYX6HfsvT/XM2YgBxaR1
XVeIJyPCV0aQJDoHappsUWTod0DGJc4Ub2ag1nONSHG8tMhBljhsDCiKVBcwX3DL9qxuFoYrKu8q
db9wjT404veLJQ3PlmS/ema2HNiy6lzu4il6bIVyqiO+Nu9sbg6q1NI2NQzuDUjLuIQT/xk3lTBH
q3XnUhbr4pr+zce2vyDQDihPge06av+o2GY84jKNI0+k63NCVyEPoUyndTatZ/z+kT8yRUACFNhx
CVPYdiSj0EKYTISE92ZPcdo1WcXozGwxVv769DQrxHyaCmOy7695CRvgcYJR9uvQrB49ZukAPa+c
qnPgvVp+aOCmoYTzTuULLcjbHPBIITMC0rk3Pq1Xhm7aIlEPOOIHHyJfXaj1SazlBEAi22WSbhb3
sKO5FJFAoDjYUshGnTKtknl1Uae9QTH8m+ngabhoyDY+be4TWlmgPC+/V5bK0EdxlslQTObqyq4C
VZdj1HJ0UK+b/KSla8moZKmX1FMemSzywzKlE/UOttJNN5l/PiwGGIzHtsv3NFwYP3cPIOdubgSV
HEMN29IQEzmIZ+buZ1+Vmuv/t8x+pqASJ6TUkF1BkdRQnEakaK8XPQIcIbDdirEePWYRVLcSOmSU
P0OxDiVjgNfrEzpGbFYxUrni5dfT0uXAy2YBBdJNA6KnwB8+mW+/RnZ13TbhH1MfvSH9SJ+tyXyc
/Ve/YanF8RY8E6O+S/J5pPjcWYgULsmgk7hwKY/p4wf8gbQ1m9GW/xMQgP5OpHeKeNsuh52JikIx
MTUz767XX375cLc/HJW0aCC7GG8wX2MF5BWvq7EGfvSHs7Am++bBQBv3PRHHjBpPJhE831GqaNJx
GyLdRm48z38OATCqlz10hCQjHrLfkNSfbmBkj5f0A1T//IqFbS8hVhv25d98P7MlejvCEh5Y8yty
XOS8ebsgnazp5+mj2FPCObW1wO+qLaosUwhghxoIdqA6NzMhc92cw9GVhYR/sPl8UaMSpwvLQdTY
JoxQV5SBt2S+PWyas71YXgshteDIF49/5Wjaz5G2Q1w7nmddSFSQPYz031svtNDBHHmX7wUR58io
JFql4MWPWd8vn7MKh2lcmhyM5T61AftaGwLzTWu+7+bdTxhTnhvPICpRiA+scgWKQPwTHZWypidx
9O8ulu0C39oeyT/mSz9e0YAjUX5YALgGV8IaTmOYZy4h9pifOqHlDDSZET31Jc+G9R3pO9YXMwRn
gXdumgq5BtaVEzzKDiWzkB+0yJgAe37PsqW+78Aj6RIVFIARy3HozwJEU/Nxpv0Z4MJN8i3v75f6
7J1+BehR9eALgCeWcwwQPYANQ+biY2Dpu8b0en8nBSyMyhmiroute4wr71v/PrVCvbZXCQvFmOmY
v7aZi2/7/F/XmpOLgAFnmDXok3gQF3ldnK+tMIIuuixmx3fBYCfTMEMCfGBdjFZ25mg+DsCcTCyk
rjl8ANalJjJIF0Bj6pN6GDe+PPRAFWT/Ngk+EDUuvVPtL262FTeUxBBIG3LDVaiMngYFqZGRH32k
z5Hbh74d8N5A14lBnNSkb2NbXmimVZ/WDBKMuRDtORL3Fbxr2VxxExtXFu05wcvxBI2UV5HjuZ1p
SfWFV+JI2S0LtVeAv5hYWDS0RRBPaCC09NOfeFGRQFzx7wGbDptxxrrWbE1GCiQGRlCKlQJQOHO3
SXEJMz3yRgmSdoJuZOQTBeDPSWPfUj0nY+ysajPWrsSoYyTjSeNcE51gyWEJihHOZtpONQOTyzeI
/c8C+1WZTtLKuHc6kgGsa7WJrnT8ebOQdx0zO3NHGp1w3WH1qnd5N/wQRKBZ/x5Vucr07wQ9/KHs
17oct2KrYA610vvR59f/amctURWMb3MLIHdTJ4CFLeN/sdvFsgurJuXic5kevcCWkSFoeJ8TefX0
8FVANYLHIJkPoJFfsufI56v30UL8sJU8xq8Mtm+2WmM58/yFaTSK20vdprAEc7wRl+8UcJalPW00
lLbLiVy9NjjXq4Juo1r39pjl8VNOwcYm+ozWsp73fWOkCh5J8GxmJsq3gYDkdpEVZ8hJpubavABh
ytFqQ6Ll34yZOtWiWb82Sc8rOfpN6ODfMWkzif/wLyB6m2SlPCZDx643UGW73u4Ga0XwZk+DNuq3
vr0P9ZDgheJi/38UfCMQUSx50wQYCmCWPnZQDEnJUasm0aFLzDvRHbGqk4gErW8D4cIp6oDr0qRo
B+wM6DSU/OIgW4NGzDkLm2scSx5bSqBjQaxcZaeRmNo72Ot/xWjMNhASkZ1bTyXkZaPjCDemVOq5
dHAWM00+KMvjl9A8v2Uos61ixEOrI33McqMr7JD8UxSa1R7+2wawH6ErwW4JFFHy7RBXFKYIjr93
RkD1NHjN6/tVJWn2DeioWuBw0MHwPJnEWHLZt1fOe1pC49uaKHU5bP1BopWtAu6e4UzCTTYp7cqF
aHhb7cDs1eBlABPd/KkUhEL6qM72i7qYwKSUDKTn+XN9KqMcrbu9hAMCLxlJDxtSf9pNEAlYaI5e
g+vMYx+A+m+HUVhlTp6PwrLQI33DhNvALTUNBweheNHAyMGD3Ak8lh12du4VlN+TA1dTRCcFQA6o
MB0vl+7RFXo7CQMnV9fvwGnlvE0sIdch9ue66o2gyboGanEmedrfUnjKyuIdpYa1J3tZsfR/+qeR
5BqlkCu+Qy/pUmT8d0Wy3s1MpmT1j8DGPhMgzj5+vOs2JgpfVnRp56yoqSVAO5t0IZAvcMcGK6QL
NMNMQSeKqIWjUhkiUBulSYsZ62hQRkLpGYwhO3EsLmktd9BzkMv0v3xOgxQxSznopfatIQ1brpXv
yStvtpuL8aVaWhCqBrQmCJRp1LiS2LLmCyPmNcsFZ6XDkLn9qsu1wkFWUHLxPvc4lz0KznNJS1xN
FTuz2jjjAZ3D2DtWmzwy6YBCG5FB25qg3bAP9PbTMsKbJrIxE4D4ImcU6MOKv7p7WK2K9aUOexN5
mF2bpSsc7w2AR1AGP3aMzmp0IQuQqtq3IDlRZlcrH7BOa94iOxLBsRwSponU6bEPu8fmkqOPj2Ld
bkXtTstakjFYoJt4atOG5NPjt1auUPT2QZ+8aNd61EBNAP4R41fniH2LqQQnE+koarjP0xL8iq4B
HgdwQAE9tplRB4lbKd1DliXgY50KUBfVx8fB7sJs/MkBAuPeQ4W4eILRQGnRmfRCkqrgExB9V/LS
CYkug9sbh2VH+KESUQxWtqiwSal2nAtMzHeZg9xOh1sWt8ULPqQStFmhylTzkBT0MW3DXxB+BMXA
ARAOzLchP8lREXgN9Sa4y0JsStYQ98B453+wl3seTMBQjNICHmiIyeJW5tZ0yc+IpSKQE+T42D+E
CGHkQYJdAEcsKSFsYfkQu+1cBX6VdwZOXpwQRMBIoAtl1z9uf58ZXONdZff9TIhDbEefZRuhS5Kl
j/q5C6ECRhk2m/ouD9E02lGof7vk+1q/cwjYQ91RBd91xlCiNRDaNs4ZuLVVjiDiy+sTbQO8SA2W
Day0XeoZ9VUvrynutRQ/KfHBTQJONVFGvE3dPIRGCv6Elk8djIuIphJKqbx8HNaLaGlcTYcYE9t8
Zdcp8oKAkysvmAL4Gr2XtG2iOBArMAcv7zRKj++20bK5hEampTIJ4FqfnzjhQBy5sDgkaXv3fvNM
fi7cPBC+VUabxmoryV8jc4A12rYqSDswrJV2sVPoO4rYGKBRwDJfnbpbmClyDztjf4kE+q4M9UWs
QwHFHbOEZHYKwl/Goc0T5QyqVrdNfIl01UJai40n4KFVAoH0vjM+gC+FpSelVa0rQUyX76ZKuJC4
GV++LwRtvUCxyXODPI1tbq786k+A0X6eAV98t0xP/vwPLEWaMXYsKc/0u69k4giJnui2zphl08oi
y7w2kXCkNHXACLUPODW8Lix8lXINSNDrzfs4uBeSY6+y81Kh0bD8QT1CNDLY5LJkqMmAnSwoiKgY
VpIdn1qHCqMKvubCFrcUqJp3TE7QPoOaGcxF3yr4CiKkJkcG0u8V1QA17eaRapzMW6AHGDf2H6kK
u1na2madrHMJ8CrEewwzxpDGaVJfuqlcgsTO4buUvbTDPlSVCAlzg/MwKsfdGk24UWP3M5oMPv6s
hx7tZOutH4+UwY5SfDRwq5+WrsWFOpXlIsrvhyylAnw/nDGHXV3LQoO1juh3bcggqx7lzm0tN12H
RZMQKYBhomxknrGib8jUSp0bqzV3TuTXx/i5hebWNrOr472j0DjVHBxwvunG2U/qRzpwCTWxdE6m
SSmeHbk4V8+DcuZsQy2M99N5zbsQ5c1Bkg6AWbf+4b2plK2xjtWLiEvSFL46T+RnsCjeA9EHmHDD
mBqx9kwas14wC5eGaVU1F2uTZsw2rmjmoapDVdXSaYs4LGxRFH/OKrK3Z74VWtjqauDPfllKhStu
VtwLZluEDVOaKJudNKbwTkRPDAdUsI95wsFzMXHKLMA3qfwTc68wf+VfvT3gy3NKhW9ennOQFuLB
nl3MAlu4oEZXn19mf28Cnrdpy44ytTlcrRqdFICKgeCxb3wpTHf1iqASlKS+/F9CBajjeZfXm47f
qFn4WhJL2s3aKGobVvhEeopTUInzcdYZi1OS5QGtXA4PNGBXHwnmX8Plq/0QuVQKJ8HBjbA/RMQc
8lyccYOlCsdgwJTbmCFgcHHsbB5NM6xXyzLnFSIa5GD4KTVt2gkEPP7P986d6boMkwsc0myOgKvd
EniviPxyYQtFnR9qEAPN1vAI3cwSoC2z7+JKZ/rrxa5++ApZXcogKxCycsDaU8iMS5XLiDxuc6hE
25UopqnNLDAh+rMgqSGdxXBwTGZ0xq71zr+pq3UKJ21bxfwlG+FqMy+k5nlb3+mVcbbdMPfOkvaD
mPf2O6LjdGbjl+Ybv0ldd69FUZFzUGEvOsMyQ6EM9j0PSJO+EdinudcBEhDvWADFcrDvZ9M22i5F
VyKPcDKQ4Tz1Y6UFuxSuKFaCoYj50GIaygyes+nrvsA6uxqCw3rfD08DQQbt1SAr5TyJaZQatS8J
bUjruSPUdP8BLqYkhSEp5f2/xCCQyX2vzVOVbAo6IBETsH8Lv0DleiT8r44XmgYRrPR0FHfozk3g
YjFud3mOcDMS5yyUVEaWLkJSoUrpsGWzUgfwgitdqIx6fASf5o0HnW+7Jx8bMSQ18Ul7yo/ssvfa
eodGT5oHXKG8VdLIlpgg3YPczcqFcsUpzDQbv3HA57xwUCtBBkrZYawZ+D1VAE7rzNIJzW1xWrl+
OhRHImcJFH7fsEf2O6XvpMBhhDeoBgWKRqIB9fTcpdclSh7z6quvqyd6s1WjM6vyl/0gklc0jCcs
R4lGaZrnyyF9K6UpIs3y7Vh66zIzrvTDMW9Bd/hgp9oDgxdzyGOpHMChI6UuBiHjX3rkHUYqyUI0
Uyx0xgT9ESw85N0msui4H0p5qNg50f2AXBI0LyDBwwvfYiKVLeWsWX6HStPXAJAndp6LvMWJqgsz
uumd2wGMfjKbjs2TdNGtzyiSdMiP1UyaD8q8A3brg82gcqSG6xz0O2JxB+8EVPNxBCTjeF2JUNgQ
FwTmqGXxTyHqCVQRYr/eS63Zs/kLOD/7e809yIamMQ4f2vPPXvaGoow8bypH4lYL5XwMk9ckEUXx
VpkLvbbSeGetciuPgBKWCRqo4of/CaGkSEssbqYnbSko2K5mA+keQQ62exR/gvt3Gc64OOcqe7ZY
nxxtSganJYv9v6/3YMnByagW/DWAWovbkASaUCxNTUb/c2uw+dEOkgfgxZQ2AurAKE+1T0VrUvzW
DyZgbtQQDGSROr5wNnF5eWksqkVRQUEBYHcbkOG8DkoIEHiLOBfSqX5vZNStTEdUaR9BHYQzqZxM
9jkk70jsWqtBhJbhRFa14oVs/1GdDotYG918PpTAXOxnn7SnHOF0fEoCbrX44SZ+XDpTa/HJ5CJF
CUYUvSAMLewadiZfhC2Ewl/orpJNfYERSTN26zSslIB4Dat+Yp51/5VPvjov9h59UVsOlvX1ewOC
ZZWAYLJjjjShu3dKFUoLjqckK6PNHtaXM/N42TRQQ3J1Rypwzc3ABVapl5IMwcmLC+gE9qX+Swhx
o7FoaAQ3oUB6CGv90NdUBqN4BjDRAcLZefG1x4JpfLcSvHcq38OsGQLw+vkBgJiD0l/vVYCW9StF
KDcbjxqT80/IG0MLX0QrA6kBv2CV5isrnyAzYhZ0DEZXR+mUzo/q3vGdcRhIpwCeNeGaJ/P74GFE
M1GlGd4QYCsq+cJpJC705xqzuFimijbogVriSPJfBV0pS1KyS1KcGYqZB/kkLylZG0scoWbUrKcw
W20w9ADfFkXFc6sO8Vvb15mIBNa8Cu0I04uwBpxafSi5Yd4B88TG1LNSCbianD+0XCmDyMShZH62
/H+0/fecs+xFkBv40aa3TlmByZhODemefT+aUcuSV1bMwysKWIgN8lspLcGKNgMTQ/ASe7mgBpmh
Xw/746NA9BzaIx2iOXLtP3d0eFyMWZfiJSFbdOtgObY1hAn6GhzowHa5XPK7jLA/NHZD5lOKOzsn
gWPKVzrwlsvh4uVpFbXXNq6v0NsKgB28YI2BCSe+Ulb57pvRE1edzTEMfT1lCIdBOfpAuvOSo+Ya
4zEwx4QrWbsB8Ny+lm59gMWbbunQHuZMBqkWhGTql6WG3356yS6nJysZaxhJsz3zkS30Flu7yp86
bO+/M0360GDO1XS2EukvoIjJlS9WARRRkQzqUdUop86imTyfEscH2ntOnAAjRYM7RukrSzdnuGw9
NQWvkG6/0NKrfVA1p5DV4IgSxJsUdrySu0em/UwOYIZoPOMq2mG4jTjlMk3uEVEY5CP3sSsnwpiY
1I01m113JJdPraE6/RzPCuHnxcT1w2CWlfRKuExZGrRTAxhAMJnfYMilip1AIV8060y7wX2W037M
ynZNccqKHKyA7IUMqT0HTgECL7LMToZc1PT06h011paZGPTJC2O2oLDbDA4dJnyTmwE/gLg3gm8W
/k3fJhSfxE8BWUAOuACnCCtflV4qPl83RPYV67DHCanAJ0yBmNCJnwe50oQSgLcr6fUtQfYqX7i3
FKSZqE0G1C7V1VBEjTHvjIZOkHYN42q2aUX9QmxfT7QqyvR1s9llgAlX2OJNiNjE43pc7YSVF/HE
fXCy3mlSmOeKgyQ5mxXuhfGTfnKu58Hfdgqj5c9AR0FJPOKSjwEid/Cxx4reVTC+LyTGtuNWeF3N
vQngC8r/sjUORpT4zycJlBM34OlwLXlYJslFgtuFWNk87PElkg1sDhnbUBhcdPmpg+nc0XeRHjj0
MrL47fvzajowK2hIoSKqaJl5wbQibkoY+WLB+goN7US4Rai8gzC7ct8+sg9seeRfGA4lcWPp22+A
2P4eqSjAPsRHkUTg3VPx9XPF8hO24ZodZqHnfRt3tJtoEpAm6LzT8EphmBC4BmDFdgY876d2lVN4
uEJOxoy1nWZsFBFIxPCtdR6IekKeK30q0So9ucziXfZ6cStxMIfudxyZEMdf5e81ZDAyyyxX7HLp
catElUW09woSFvRKziTl9hEXA51v6imgKZf85QyoRQwRcLv6cQv0Ctkfgfi2e2C21h3Qz8bwjNo2
JGg6U1OdwxO3NJS5f4hThWr5blohZu3p+DQo5shuGivo6QzA1z+CclxamTZ5DqbecAkaD/91fxEH
/Ta3QvZvLUIR2H1WjvT29i82B7TdO2U6FPaFTXoc1wAiVauOESxynWBcvuVh0onpAYRXiaKwton6
lUmBrqm032VPG1e/J4x5mHWgpsDU9OUolKnKkBo0b4sLSYTfUcE9tDyRzuWS7Cnb79Ltyq/lEVIU
Bhc7cHYzM41rF51mH7mQIK8Qr2bDrOIcmQLJOPwMKvOT/rTALjfXg2dhIoTrDPy4E9a5N9bNj2ON
NsdGrBfo1uy2QIHeoeIwHSehphuAnGdcFiXmZnhMU55XoFnz4JgwX8sAfLIziTS0nevKKiU2W6iG
2MOk5jev5sVi/jsqOrQABaJAougA3IrdrEoF/t0S6xwG0/dnZFmbrLOLHAd7Dewx56nJpi5uKvLv
SQ+X4GI5SowWCVoqFJBaUZBGMbHMa2fDQ1QrGNAq31iUs+anbPtYKuFOZs6KZBkvJz15t9rcCa+Y
vm3LsW5MMJIV7z/YUDgIOdsrmIpZE8+cF64rGrfObeNseg83J5qIVfin1jm2lgJrRsoOGTLo4MO5
meC0veRzhizKK05aOpzFdviGFNo8ErKkp3dK3y3I1URsbzDuXrp4IZ2D4fGLI6JuFqxkDalfauty
v6vLtCCXw7suXy65f5A48jXbKZAa5/lnSjBQkan89cufBI/yGMFb2lcFmLDaq/kqwq8CvMGa7dhx
ey+iBOvDlOm+nQg7nJrCFfg5CXzOKG9H6fywivuIxemuk5k8nRYLq9J45z74+s51r1FQ27trzjEk
Urb08kieag13eJLusAXjgIh8/T6GfSkQvPfvwxboYYh2X2YB4nkQ2M3KqXZBNfB59YhmwqtXe/VR
0372YBE2bR9eCSLuKem6RM8103NcTHDZg6M/l/FIpTyGg3dmAzQwGa7EhLmsxf9jMfmuoqg7mnJd
eyru3TYuQ5xYJ6JhlbSLNRKq6LxAfx0/jxpcspPpkXhOy4ysBW79uMv4a6t6S1GizF4gobIxBjbU
KUzwvrdSuSX6DFwyk5LGjvqtrrGlyu0SEbHe1kaY1GGm9A/TJkk0xsTFpFe+lB+VG6APz3heXGV0
H9j7vd7yPVPFRZJkSayfnAzHTx68jXLvsCRV4GY4Qw+8L3aYz4T4jRKnWuBn7z7sUvcw18CssGQb
vu4nTENEdVlEA4QVpEnvD+rK/TH6v8VAG45aQNs8ChNch12IyKAm4DVwRnmfibgsm+r9y+EbxULu
KZ4dFwzI9uGtLK4Oj1ARCMzJJ25ymvw7euPoteEhzVp5Sm42o8xGbi0Xv+am2GtjAGpXlWOLobbP
YzSDMvg6S/UdFNYRK+5guE+f4yW2tYMXYROEbNTN/c8F3uTMpXdSO0TLhMssLFxPUsyR40sr8vat
RV8aKzmd0jCbPRSJxgxvbPO5l9Ld+rWLDwd60L3w8rHav5xQmUo4hxq8zOeqQLAW3LLZsCzA45lE
dlWv53LL1nubtAQADqya0jLaDiR7AAb8kTI+ZrlMqnnafAb/PnmFmzI/JtpFv3RW1e8dNoRdWtkj
sSDMw8Hw1fXTPjVdt+i4tEMn7IlEVQwQ49DiOYnJRZKhnhCwf1wp1gzLURu95afBvnZ+u7Ey8eL1
crWNcM17PUvWXwPDUh4s0D3tD38aJ92EHNNcW2mHhEyjPfDYtqg/H07lC+ojaANnPPNJTYznzThY
u2biye+aHh07ZHG8EPFq/EfFbmYZ7Oo8d2R2BbouzPADxD4sYLVekSyLHpxSn4ikEWPu/xJ4hbSv
iqe0yEwAVIkGAox8yvjPYTSID/jNJRt1eJdqN9wipsO6Q0UIrUCrXnG4fl7mqjeJTCY9+Hp4BALS
jDD7UYCcnBKXCC40qcI+jDEFL3uvrxJ7SmueC+LBHstCDYebxipqjJHcvHzwZJTogXWaK8pxs91Z
MCSt4rmmt4ADdlfDL49zZu8Al0tiQ+Fv/6oeF8x91uUgbO4h8bo5mpeB3ogCPrT3IKaRGolWIdS1
20VHBEbf2BaAZJoFimRnKfIivS/6qJyqtWlPe2qe0clAw6pGGUQpzijfOfqBeJTCYBm/fejjmEwj
YqF+Pf/rG7wXbv7oHWVuN6R/84skX4SJ35JRoBwV3fxAjSzgu0nUxqVqWY/eCPRm3VUvmnF/fM9F
agVw7jE3O88NziGsmoHL7Ob6pNOFurLoBnxsvqNQ9U5NNhp4FFTsV1eL1g3T7o48Zk/GIVT5auaq
KSmNC0nU1OPx0INDntsqw2HnTBanwu+BAYx796gPm/RyVn9cpyjcjqQWTZEow+ZWBivx9jkyoiw4
+cCq7XHGusOIjIBXuODSnUBpl4yMbaFB9jrWNIZXxoL9JRrZOGaEOSFISyNlPHGQN6jO05G8Yy60
LuNHcuAzukh0EYCjspKv4OGVwC9HN6Sx4m86SxeauYpRXhPK6wFk5udwpeIJCn2LUZDLIGhUczkD
6CN3280pTR0Wxe3b7MmjDfEnaT54FG/0zhfAm57LSqUe5FrqnC9UnZWQyMza73iTj8y0lcRqB3x0
YBWrcmeBcdGYM1Ox4K3jZr5Yif/fvGCgExwHxwiZosEeRhKuVK+YfxJZ/TVl7X1XXEDsUU0FXZ+k
UoJwZQzR2NATYeyXTEaQ23sbB6pJi26wTo/hV+wLmrkGeUCrEhIfPbyV6MY9SorssxL70MFrtDEm
1nre5K80WAkiUUhPegjBRZyE1vBeZN70ZRYO1SJ76zX8k1Bkb0pLf2WcOFOf6B5+JBZkZCl6jlc5
C8JfNBRypK1kQhym3QIvuLt/+tNQ6ci9WOAj5DmKPXzTriLBmszdavZzpIdWx1zD+ROpBYTe2gpS
ysMlWxjkP3+JPicoYNOGIVZKBqhthUbSRINidpB9uCpjA0oBS0C+a3Mbpq84uuOQb+BjrtakztDn
N5nJ85wuCKW0TNisqmZnyVzSVHJ0aakD2EYgHH0R1UdFUiYyBQ1Bin5mSZQDCk0hMcFgpoTPNiFx
D+7co6UPMDAJu3YV6M28CMyRf5CGDjVaYk/TIeF012dtRCURfp3nFBaCalxS69kNMQuxrQPLznVt
ev8sQb77Vzpv4jjY8kgzaAACtkXhoTvJiePWWjIDPxobN4FjDXl8/r7tCbY6XuGoM64h8c93Hng+
f9aTcLuGh1j7jp1DSwYNel+m
`protect end_protected
