`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cI66OANCJw8fIIQbdpCG1eUZiUrVUYlTNQ823416CUh5RU0Z0lUSscJg0VdsbyeOG0GIlqnKKDcJ
g+441OyZKQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UgqPJ9i9WiJwgzx9hA1QFTAyJQbYygHQhueZLDtbtfbgNYIe9Vf6qQf08t96mKA1gKActJ7BeV+K
6uNMiJfx/3aUXCSX1zJ6wf3n++OQDmqvxVVq3gnHpb+740+sx3yxZnt+NIQn5YfqgmEXSODHM65H
T6IlCQG0Rk76FUmssyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JffVUoJGoNenA9JkXMLk3KS8XcomfWAzcMGUl6pS4bKWUvYmY13D3pemGWR5ICLizj6/IEASX4qM
MrcOHNOZ78VNNGbrwydnmhep2T8HUJ/34A8F6RlIg3EPqaoJseDBIuA+1YYmvMYUPXWmDmWnG1uq
4OVHNHuSMmViCS9G0XZMw9OZMd079W0WWlGjxgCIsCbTxgr5NySjw/l7QR6gLw2PWlOAIibLSL/6
FYbf9Pq748eBFOa73RMaFJULQdNMNcUKu7XbHElWwAbBAEQETSA5PY/T0Ovuh5VWjxfKceXk9gE2
s16k5nL5jvgzFecQSuS2lSlURIB4qY5hje3ZOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6n3r5uCHMurGEnMpYNf4UX/MkeElsrXqvd4MQdfthvZDOuXHZxcs4tSf3laM+WPFVbsOKpN2K9r
vOlcg4pO3R/XBxH8buk6fx/j1Txb83yD004eikrbAzhD/XMeJoB+vwnOXVjryL4Tq7ewJGiuFj3j
3aajz5Netn79SPqpagQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ux6EQpdIiEpdxg0F62ecUw7+0Os42ovKYC5a4J5nt6L0NXwWYNruQn6thnH20HG3CkZMjYPVsVdV
6fsAhKiqralBKaBG/Ej9eLWDO0kqJYBDBHDr1KxCmmsfP7tgcSeensV8aAfsf43ITwJDMIO8VHys
LbnRxuW/uncBTBd8BpuuF6FOlCwImGuVwEh0SYaZjLlAA/zvuQGePlYAraOXp22pKz1CICW9YEbL
RHIga+6SQ98q3/eoFGq1j3ZXVJuLYcvW94K/kJlph+VD6UU5Kix62jbW5vyq5E8KMpqmJr9NNRFn
j81j5XKXBOZlfp+VVqMs7Hlviysaj593wan5HQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33184)
`protect data_block
td5QFuuLITbKOtkE3oI0mGg81uxEpl4OzFN3dx3S1ftkr1FB28AsEjJ1JzlMER3jugQ0XxNHpZ6B
MQSg9LCC2ub5LNwlhvbYEAYYqCK6ZgIfuBIOXcuFFCv38YT5eHX9DfFv82XjsC1Pwn/wMP5pa3ai
+CgroYRHrtDe2OQ7DDSoKthMBOUrZtCQsLcpjdBklVQoHle42cJze+4ZXpPCwHRIDOHSWwcXVFVH
Z5PDJyhiEo88YeY4Vx4a8GJAYjI09qomGasMdNkk2A+JVS/7GhyNak3wJFnlJX/k7LPenVoItKUB
s/5iWiCmE11UdejaLz6uyAocKBkWSlogCXoG02RiM8BXhoIKKtYL0aVBK9H7qEdvnC4pabrGQ+a3
5Nhk8hoUU1OO9XnwNjdkvce+wDiRqOL4aZyURFDtGCZs/7AT48+cEB8w6abDh34mrLMunExIHThR
Amdt/L3h6MmmaaIWX9eT3rZSgNtGcoANmzaiQFhk137m3Ud0LRhrsKAjhVhjqVGlGxAE91sl6Gt9
H/oWsIEiVPyNJCgsW4RKtgvBMqmVYOz+BVynh6oYqM5W5KavTyacVPPPbMPKKs7+fRXbewFttQsQ
HI+4k/h2+YPsjPBBWqZ2vasUvbQQUxi0X2VAJXOD1vzt1QlGlu+bimTMCg5G7VbIGEf29U1jJiCi
EISw7JKofVo5rF5DkqJ4lnBD/kgf1Cr4FXXhyESZnxOFJbTx1MO/Ehw5WciqmYpXyonkvDtjAGRp
1SydFfM1SQ1XfJCqNH1YS8CubrZkqLL9q61j6se5RlmpJ3Pg4SVbla+YfHoE44hG1wiQoHrVsEdu
pu8s1/+Tpn02rREVGHIBEVONy5LHF7yYthb8c/IriHUl3BNJldwAxL7VHftj5YUeukd53JRf/fNC
cxlDbs3P21VsBOoV9swE5QAUHo+lmh3udcf1FC0fSa+5o0qnJ//NGjbwGZ/TyFSNd+VS7OGW6s4a
acgs7aP09EZN6UheMm1ORfAe9LYVs213E0bP48bUaYI0a6IbMPtye2boiqa747e9o8HJroll3JJU
dc/fQCO2AjTRTXeI53RtrUn2+m6IByy61c80CXo1kyVfS3wmwKUzkr8N0xZETubxmEe3OpviEbPu
cGbknIaS37eexJlSFJZnIhm4ffxiN7yQKXk1iORo+XiNRHHKLbUPojK4BNGfCKx8LW+ZyzxAMEJg
Hy2s/4G3OO5QdV7dLlGxav8i/9m+0ENQLM6AKkUliGNvmS/js6EAOa8kI7iVRY7/9aR8iDbhFZD9
DhIbRCO5MoxqDe2Y72PIA/lYDSzjoXnw7GnD/tgnkQc9Rt2wkm6+fzaCzCGJ7P2mZ6fqjDLVsfdu
xJW/l0LUvPANtnKWs2wJTC4ya/kXWN2yj57cP1hVS8V6glgInIUvogJkRfogL6ozw+SzezMMpLte
Z7Q3kYJLCm79jBYCWjVY3hDgO34lM4SlLSrIMs38r3n7G9NEliIaD2T3zJMuHjQ7ewKIYviZp+eG
wymJFAc+/6OBu0OnGwub4YGHFAD4IY3Lppg+9Hld4CaEM0yKe/fLFd1c/Lf9YUObfsXkCHl+KyvZ
+kwpJ9c1Xm2yoMp1qLx3bowbHuB0jE5H3f5pfE1yz0YoxeBJAlcUm9p2goSsnGDYxBstyR0kagFA
TiCiwX+SYstArHj4SySJlUi83ygq/8rgfH8YZ7LTan5PxA9xebrq7l3H2JWxUPyGRCW+qnh3Gb7U
KXyjjPvuDBY0TvKam9PRwSGBSgvtNb0bYbknlkvniE5wSwajW9QR7Ynfl1uy0UhzJYzOgQnfR1+v
vO9xGAJywLS4bvZZNTFnDUitNfOyQ6FGZ1sb73rTdMno52ljLKMsBXlV07jbBVeilGAua3jhA1+h
zEq341VauDCCw//rd2roL45WJ2FQVr58B41UeCapzItv4c/QGoNW+c4iQpzYRXVhDpOGCtnjjJH0
GIYw3nr3+XyY6j1FvIQeT7dAmv8Fj+KvhZ+jfNy/9ZHJ2qIP7TCt4CAtf3Wn9PoGJqDEc1dKVMPj
xi8ECBUcxkAKQGvNEgjuPRFcVlHr3lsOBY81e2K6H8CFkjP+wjA+FJyl/yCmayp8UBFWn/7s/uAj
DEUnRxjCMC+BoS4AuXAXJiybWn9NDV6+ikO4/Z4U1/T1/p3VVBy0mwXi3Du2dUVat0pm0x72GoqY
nH4y5Zocy+uzI+2tkB+GUKvCy4OYBZvi+zH6VZiGgy0tzAehskpFbpn7Kw0YOS9dwQCsRxWGVKqQ
O4A5Wog/2DlTXctdZa1Dw3qCLAtftNr642+RXgqkPutiZxQvqQGKZxhXGGtMlCTeIxRISBi/JH8w
dIiZb9q0r2xZgCzqkDFEb5nDivtDEIzU7P0L5RsDmznRVPfYo+bj6axI11EnIyOri6rOTI7EtnD+
/6UZ/cKXAVE8w7HZ3pD/ILej/3v6PRzHWJDI7aI8F9LQQ6ERi5zXySH/2+bFfOXrW1KQNH9HjpZA
cr5xDrT/ttiEEcc+1oS4xJW7bnngQfDHqwuhIjIlaRrWcjz58SCD87g8avTkIoOtvQpVHRJrqHwV
WOjfYzTPZZRup8HUJzzGuACqjvhTegg78ik/sus/iWN7Io7cIfPMniDNc6lKSKdQpnnzivsC3DX1
+QH8g/KSzAlxQhn0hFQf9omnR/Bp0JkikRioqJW/SKBHGm4MeIoe3j2hYOGSLdB7pBpBdP8zmJqW
b0Q2SgSsOxS0A5wmvB7kiNR3BDNzOZq5Bq92APKc+fm5TPyUomEOen+vEtRSoiahIxMqSaSAz9Lq
3KeUaoOX+tleaME9FoPYU7r9DLFTZzMEx7BYsQxFFI1RQI9iHORN3s9j66DzRp858759XcEjV5yw
3i7jk9uFbtseOv2aG3Xn7mgNBC8cZtxljkrR9LcZzmNLwu7w1tI1CYoZ4tQ+EmYB2Lq5EYLeDcif
6GFLUxB4swhTPWBkOhDnEODxQADKq8HZE34B/sGtwd5nbfPzocFBeCHu1LQYVbsjjOnZZn8HO3Bl
23Pad7xHijSo14uZj2rPR/DHvwV8pGLqd3ioUPQ0+jqC4O73bu43d4R051mWnhLECo1i/+nRzFRa
vyloybNnfhNhXU3HGtJuNOd+7btYgusAeGnwoULdD5eRn8ot+HW/BY9jdSM6+chFzT0PqL+QVTtS
vSk22vjJLBTeiF97EA8gnGtLSDKqhAPxACRjToy4LkkGxQvWj+PnMP/rggEZKG51VDOvpTlA8UnD
83sHDzSEAb5urFIMuL1jTlHJBIKl9sd1kNzKI2gKiFz7Kl86HGHiu/vHLBbr8iBJk9QPFRc9XrBU
kFi7e4NARYwNYcw+jSnoxVXZ02UOwF4+VJY5DuUmJ67ulj2gkpcYpLSIV0cRRj+Db3hk8CNPA2Ce
smLLLVreh8gVnsT/llQlaDViIOlKeYEWEUD1+V3IBnO+RzMFsR5sj/ibeT58kk1rosr9l3cdMLD9
az8GEqWNm8Tyci33uEKTwnjenYtu5Cei0X7SkXmNi3SXQSZvQ7u3IcZ7l8qZvPMl56ZDJlPgZVov
7tzkZsgHvk5nSltmFICN+DlExAq0GNA7E89d9hRFbw9bqKh9SPllAKAwpoy2R6pnIhsN9mqyL6td
DSAO26VclKrtGvFATWxCpOGLV0KZbcsojOfaXT/gen5BbKW6KU90QLipiTj5C/K1la4OLUTmp4Kd
rY7mcXo+9duqwYQS6RWOenLqvukZTCcujzVi2pyMOu2UM/COYQWLoAsknBM5fZPMwKlqKhnDCEQC
Fr6Of66PjVHNOrmd2sBI8ppg6kxn46PP9ohn8vDdyg2pnh71f7cd79Ng9PedBPqn16LpD2Ax7Tgt
PCoXNSOqCDJ+PAiszw36YGO2xcMkdXrzoXmI0TSEjQ0v7EjNGOWsT4Z3oMSgV91tj2Ovg1EV/4uB
WqQdP1FvWcXCrTzpKKx6uApGaIOoV16GCmfNcSquzH6/NfL/s3CqSdf8NT10IqI+C0UyVHLbf8y1
s7S7OzCLvPUDVG6cIiAONxTkORu/Oh7xcsToS31/o7M0zf8ux8QB6q33J5bNBlX8xhfIUmgG9riD
NCx/QrlRkbBt/tMiYZ9wfrlqpWEule0ZpONcHL5bTn0sr0e7+wT8RUTBgK8IB014RR+mJCMSkKFp
QSR60zh7/j+iyqnomKYqjy9UrmqDLTggCslN8CqsGI/BvxcqiTXqR+CDs4BzpHekX/lzn8TEatdY
BuawWt3vDR/80/QtyQfuZNn2479i5ETjZNJGhgl4asj/pxcW5SxaGkeoTToQaPBUasLVb/cCSloE
YXliHvZE+2/6O/G1KqyBkGdf0U7WjwUFv2XaKLNzw9l9YicPM5l71HaxegtEgW7zEnD8vxTdvj/z
dLUGb5K6+ilD8bbWwBVqJXXUTISCY6bW0dt0nUtpkF/8hTlDyzPE6ryWaGIH4c+LUjk99TXpsjzu
shWJxyGJSlgOhPwtRyQBKZBhJQemBi6nW2wkw6RhzelQZJIurx8/pLncLgLz9LpLpYsfv7l6dOOj
NDqOK72Hen5SpbAr1W7zftEXJFXxxT8yd1dr4XCvJnBb182SBHEXXW8HAUUfAIEraD5WGAf15psP
2VlRvBdQlWdOFDQtfhpQXQZsf96u7wmH+FUeL7bRHI+Sdfsx6X71OjvBb5MONIG+JTVKannqoyXh
R/Hz7+xxYpwZk5Y4awquDsDew1ys6HIa3gX4kSft6wB8IYcL8azdAVHsYXHeSOSCQXWmSwfoiBSu
DvztY703Q2F4ONQ08cf0DTtcVjcKqfCHOHLpFopSEWi4/2usqRHSMJ50H09UI8bOsGh4fLJexjmM
WiabZBfa8vSwM1b+NJMUzz6aqZlB7RPD1hGilWGRd05kdMz0oztK2veDgsiL2DzroUMyg3VFs36e
S0pkqe2+O1mdFRvsOG7jQiatMoe6v4r7x3TK9YivAjUsjrDyzaL3IvJFFNVNdYMFPI0GyCsZ80fV
/1NcGBrFfd/czv54hiz9g27A+ksIEPI9lSvx7gq/XD05HN1ydOmcmNesFNytJ5kLVuBl3LrpGXKV
gLOxFVM5ONl43Sms4dht0l0XP9ZizSboXRtIfpRq2ZRYKsyJO2c2C3OfYUlxI5xgm7Ezt2q9LULw
vn+ptDEfwtG5Yn2sHbzpRiCehSxBGBJcMqIEnOisyO21EvdpE05No6j84Pc7Rhss6gm54QZsrWKp
4kN3NpQN3huD/Z9TLItJ+GAxF6ziGlOM5o5Cz6I4v8TvTDD26JDzR6yU4ZR2EO2QK/JmNGOXnVXf
pZqDWC4p257v/+pbJWQONvtHViQIXp8IGmDvVR6oHBwSTor2+o0+2mLCpEJQ0ENsNGXUI3wfSwpy
BBPYsduDdnANHWCGqdjWJzttoI3QbvHOpYqSuxbEzM7Iso7M+UHbWUsy+Kjv8vDnqpUhCx+kJQ7p
YVzDI0n6Us9s4IZRgwif/nsg4lSJTynQOk9/xqb8UDy5yWhhBPVSwagqMSuLYd6SxV+/jBHRxXQV
Pfmi1gFrs6DS6dhNG9SqmA4mY+bp4hj2NU9eu915n44Zfas8uoVexeYj1ghJxwVP8JMBoowtXaAU
v8ZaaC2cKButhGKcGNwnfG+w4Gqp17VsP77rqW44D2HnkIKZ/ILw1B9BFvIiY7t/XWjcaVEtvMwG
On5fwOf1qZpJTWw5W8wkUJeQHPOGQjFTFaIgmm5jrLTwQK3LstN4DGOe3yJMDDrciQXC2WDo9RjP
2kPkgc0gSNgEvoFEPXcBXAnS+KRYc+09GkjR8NdN/1VZdm+kIiV/W0X2ouU4ftJgjgIeOlmy52qg
jKlKXbvGqDh6mZLEj51FEhOfrEXab4NLld+DiV9PFLMzHfWpqEc2MhmnpHELyBNz+nvbPw5YJrfw
GX1OWJ9BgLwCItz8A3BAT2UppIQ2HBUz+9ukiNs7WGqqu8hDmehcoTqw12VYCXGeen1KD/kq7Dmd
AH0prwKy2ur4X+dznZ6bq+1VO+LvfnEs+ytqRGx1rbazrR0JC5HOvqY4To1OHGEqEmpP9DgJG3Jz
0HPM/tD1wu3WcLlFVFB2Dg75IOtXEqqSJl9rhpVnZOP7q2Oi7d9nPjV8WpzlQyK06Nf12EKudFAP
XGHCqbdKQZKOE+EUCK3KfP+EymLILtAwtIY6xKgs+wjJTMEsa8D8oVub++Rc97SvbajhIp9lw0Qu
eJjLGL63cilktRyDvhDZ/Y7+C26Sb1NNW/Mq33knVjTK2E6MCkzLUQHhxcnGPOnBD5T7BGpBIUUn
5lqiI7ntPSnCph8F61Ysgi2v7QRhuJWhio95G22AanAkbrx7TWIxSRNp1CdpIJ3Q7mj3NpEYgtzF
uRgafM02c9iXuHWe5B+S5U0J0U8CfnQQgqgLEXFGcOTOvcEl7tintgYEzzowXQWeRbl1cSEXLDgU
9fsG0A6ehWGkNLYLgmzecXQqQ0L/D1E9zrSw17dX6xWHo2vN3rlTRUokWFkdPxPwvwIMwlkF3JKn
0VowTHObqlOIPPzcIuKy70HEy5REkf6AgBS2rKGmS57s6rkO55K5BFQ2Unl7ACNOQeqPV2cZFn1C
4Jp1ICYvq2+zEsUrJitKq1RC1l93HnSvqjQualxPzvLbcsAHh7f0PR96T97CUUOB4fRAScHHWVa/
ubN6zhQEX8ksHFGw1MwWVnisTYK7UNZbkgTckrsUR9Nbrqj5B8dt8mKae5TZEjqmu7PsfukH9kEF
E0mJfg4Ii8GBFT2AEnL0iq8gD9Jdv86MrH3YrNxw+JOoeon+4fjg5I3iI3NdpE4KKZK4srTKn/ZQ
e6Zlrm90ItM1kjHcmiey6NCBpAourWrjYBk2+vOrIjMP9p1EkN77HCA+Hel5I8dpCGNfpU+hJf7y
J6CHLmcuwLAE+DCWCg24jMY7rADjFlpMlCdLvIk7y1WGeIYU1j+IQB8VHCDRJKmNLOuQ5gyhMZcT
TcQEK3G02k5j6wd4CVQIuI2FMiWwAeJY1JvNOnH9+qiPYEbsNpyExYYvTCtAV/bqZ7BeCnOrebJJ
TiV8NCy4d2HqtC5kJVwSWjof1x9f6du+ftKg6aA3D5ysKhCg5NQCEYXGIQpTLv/VKuomvXbxZZVE
cEwSfSPLhhxz5pus2cRpPN0ObNA3ZdFjlUvezjiS2NLiYq25azylUfU/Uh0MVu9nG6KNU14oMIGz
GkEsZ5FkM/WbgKocv9rLOa4uUA5X3lahY91iMKJXtsQOUuE+RabOTckb3jJ5ELEbL4xXUipjk+QB
oHl/bozkSHVru+mA6roqPSFOGxwxNslIiMqYJxrkiNTUTqu5X3nof/nu6abnQ3qXKNf/thh1ahan
+tIxL2muRQi9ZSg7UIgZE/5ED184sHP9UvVeqmH31Uy9l6hOQTIIJL2Vut/UAGWbqJLjpo14Y72A
hqerIqzAZs/ljLJ6Gwmix21ZbuzWpMANy6SjO9GP6LPTgRM3raYdHAzNWpG/Rm6zad8mSzUym1EU
ZeG+RIFuHUUJqp6Elbh+cVzt/YMZfGvfzRDY864zawmNHcuZsSqiInzmsMyMXPSgyQFfmncym6Zn
GA8ohGz5aNnhtvC1HIqCvxAF5hahy+sBAqEnpMDtyh4Yqkn9qyMXZHsAWAtVGbjt1eT9TTmAlyjc
IQP56Zq3hTy6+fIh07E1DqeoIgq2fuMr7Q11DxhoKuL8zcbi+krfyk1OO9n3yNE3b7QeiRBMIEFX
3wm1tObsthma4V0kSKBUBoC7eCuIbxY8LLqFkvjJ5TdbSNg+oLocGpDxDGKROrENn4JvKivnyPcM
6ovjVtQPzQSqoo05QacodK/qCBaGNloEQVeSqsXbsnU4+PrbGeO+jb5/argHc21zUOC9O06ClBjJ
X0qxntlYfeefY1odWfv608+j2GnaVNWtFYQpzWV3fw0/dFjBM+DisehytxrMdun8wKcYknYV4QAC
++O8ChT9vyDKPGWilUgn8HG5W62gYjbLYMW6qryjL2/oUQQUkres0CSvMWlPbi2e6KMaF08wPBqX
QKyJ7ZqlRjCP975d3V6iUoxL1jTyFsaHdRcWq3lDDOlMjex5wHszMaqPdQeadFzBB0oCfKMEz5bZ
PxssxsuKr2mIYyL61Is5pHC5EzLAF3oIrx9RJdtURlb/fuhtL4XFLTtGLlxNaaCc3GQj2WVWp+6I
NO82j/WCOw5HY99cFprSF4czUJ5PjoIDqbM7Yverxdi9Nkmv7LP8422fwPueQ2aC8gptzzaib94+
yVzaoi9f//3GLSuV5fdYYqCUXJkXHwE/qdZe0FifS7faiB5Ia+JpR4rI1evIxaq+rdh1mvupddpP
qOYXOjCNivML6gk2H/sTdEo7wkNIb+EbIBXGyIsbe0/WNhcsh4Bd+eoHwCa4CoIcxkWL4AMENCZa
Rw6sLTmUMjfP1zgSKMbJkSruD/KTJxwfx4wBt6FesX/v2ZKpi8ae6BS1uyr0uUP2SFtpS8f+l+nM
Q03T6t6uu9BTVnBOxzW5I9tp6PIpDn2iXGcR/J/0INoPwCzA3b4Teunym5Hb6cSvG6q/1sxmAI9t
zquYAFbprRhYx5SzKjVfhinTv83h+6DaMYZlXoB3/Bzql3CzAB4LmSFaW/E45lrhk5yiJI0LsEB7
fi/SRQItno6rs9bbEF644CZXJ34TKleMQ2TjiXL4SOL1PecQbm8XaTDHkMjLNLHNGxwDOU/aiZ3X
nG3dP12BO0xpD0eNdO5PdZRAk8kxEWiIhG/ac6qJ5e+juuUblL4f0cZxrcof07Wb/jRxI7ya/kNQ
WDprf1Jj7XkeyomyM333DG/4eNsOztOrhlcF9Tl4weBsDV490GsFX3THnpVnWlilhfMRywza1jnx
Y0z9N6GrH8b6D3orc90GvwRDAJH7srvhEVcdJPGGoPOd1OoTm1fd9g6F4DXBgOknR+xMPMTdAQE4
b4r7u8dafJZ5V4Om0IC5eW2VZ0WRqEy4N5QdWW8JmRWcPuA26VxE00mOVnLylEfeTc3KD0XC1KSu
F5Im8vVOhyuSh3bchJ1d+pOqUKzoORHgI7cXCM72sg+RIEOs2M6KHr5vcu2NKXWDEuLk+ozd1W7Z
4IsUu82UuAkZaOUb7cA/N+AZiOjstnvM8d6z/w7vyNKpqPlfQRM4n41VSolUgoUW93hF5tGA5obR
X+14U/OKuvFUukHR1caRr9OKiNa6AW2f6zp54VJbof53/Ato2NyX2HwEZqaajpemCK9qHnJupBun
yZXpBaMctEdyJrrAUukPPVVu47/GpFxBv1safl4taR7HH3jhSXwftce05TrpRFcMNL06zRgyaoMU
g4uOpgg7g1xddxpSZBI29M4xwmi9NQeZKIaZVHstGZZP02z3mgSM11lzzlZRPb4eCH4azniQUkuG
Vp4I6jgAqZYfISVFSNqMBXCjoGghQ61LsB8thRrPBScIjDP2lAKDjk7Qf9MqEhFGMZI2LPZN6QJ7
4botb2sa6wDrvgli6hP44aWPrReVKacY9swtI2ONPWYQk43o3V6GAyLQ4/dc9qWbQ/R47Zzm7xsY
y/0Hx95MAa/gzsGd14EmQNU3wI8/qZtmMBhf6PPnHuFjX4EuaJjn/1zaJLM937tQPv49C0lcs9xD
5y2Hq1ymuoSpTWXLcDrQbR0Ao30qup9xSIUqo4FKWp7UhrDdTPvlQ++R1bZXUtby49KaX0mqnNQy
DKobDRjWPxjWbtcxzCnkjIhSlJk1CaGhsYCTKJaPkHgku6kNRR1G8YtcVgDuR0/9Nkc2zdlL3ivP
qVVvA1gdbl12YkUW101cKXdqXL/pXv22Ug0YMMJoIzRoGkgCvHAcqjKtCXfWRYTIEGcgaEj/r0es
u9NZaOiY8H3JMi/c/HZKVPnBbGMCGRkQrUOECoNqWR0gfRSLs7Ltrfm//HoOLAnuSge5QlUNkmUv
H/gqdBskx1pcw8LMExfWdcGHM97GcqIW0Gj/TZugjSJo5dADHhZVynkNigGNnJcW/S6r8/1m0EA0
9hE/erx3mS2Y+m+anL7xEr7aBEBb9FKorSIz/s9Mv8xv5YBEYBKNWwFZvTmY83X9YPQDJMmdleur
VyCJn9zt+YdPTDwtvYdCNHuBhAulX4Ai10Wwsh9WOkLWSnp6iQ37lZLJ661erxi/H4N6Lo8L1sJW
nwW4+Q8QGkIshjZssSGa8H+CKiuXReZNn6ebluowIfsrfIMftAfw//reGxvllBxNMIWS4PWX37wU
9hRKC6p6qEmRJwNSFr4pke6lG7ZhxkU/CqtjQT83UA0Ey4Yq4PBYqRlBhoJRc7/EomJh0BG1p+IS
l4R0xWrrOJ2TKeRU6hRwJg+XB6ty+qFwzNrmDtrkuiHVG3UC3p7LQf8qedsYAFiOQhDf+v38MhH4
VoMXoVJw+tImRMcG2pSVeUzN7FuqKjOWBqHPuWZ1/VpeUZ/a1eEzIC24hqAof+Zr8K2qKlY+4X/r
O8X4MKfd6DFcoHvFURkiYkx9JmDNwrlkfayoPXXYobw5rgwk9V6FM/QJD/8QxaNwOvpuklzM/cTm
WUZ3OSJjl9JU7r0jeqbGtGehGpSiJ+5NKzX8VA8gHVXiJfdqPtvkdiEkpBodqZOVh73DEWuHJ3O7
yKQmrULYRwD7gKAXmNqmUAPVMf1tZNYhjLNU07+oI8ha50JagjI5I6GIctLF2yTPqgA9ycsSJeCe
aHVJd/Dk+tVgTeuAGUZhi4HAVPJ5spAfuboglTmvlxs0aa4yNlBmHndkzVTuolrt81yqzV3qYKyu
oiSUt93tcC2WOXXqL878BZ982OxdFfXHzo9TZgHGRc1oOoIM/bUGvbxXO+YCmyuV8IVodftBwpp/
QPfKeliOoSMiyZ7Xd9G98e8xPlun6GaGyLjAc790jSX9V3IfIXD0lRqJQBb3e4j6Fl7dw5zK1ZOO
iaI8kZ5RSozTbhrHRkHzYhVGVKLFZ8jbM8hvayD8850t+OxFiLVMwXKJbq97ytVtRVbavlF2uTsN
9Gcva6rgX033biE4BFAhNottS11XsM65rBoShdw0loRaiFj0CFhY8yexKRS/0CumMfTEzB0RcH0y
E8jSLZMgJ32ypFHyeaO37JgowgFNj41ifGihGAeENzXNkvfzlKefXTUf3q2jMECARkb5TtOOZxmf
SV0gRof5HyI4S0uOYKG8ZGIfOtD9X5i6bu611H13tFBjgmy/JWU3oK/il1wPHRYz1uKNAxAaulle
pe0kz2PWRufJwSV1oQ97ViSG1K38o6NvJWkKd0V38Rhd9wrU94wr/Jqcaw4D011FcNhlP70sUy0s
h4MIaJ4svO3eJWrouzvsmtZLeT8N/PqBVecenoVqhXZoySWW1SBrlBE9UCCVaw1BH27Yq2+xIjFl
B1yGI25dJBPQlkee+hLsUiJ5NYL47F7iwPFnEIMJloqm4CTXx8q9PIbm6BpJUOFZLELfhfGhWisZ
fpzQx9sqCn1/lSle6gHLxVzoGBGv+GB/nvz9liSUwbEBhAnelpO1FHxtAp2J8Hu7ADDdgAnyIU06
/qXMt9bRxdDa8zxjDIUhXy1UtDLfw4eDuDRY2fF4lBXoJvpFmPGeORN4AiuggZ1tWw6bW9la6uc8
ubrU19d6vW+l7W42fLqaYitpH1xdYfq/Qjbwf+T+JjKh0RYClBFIRQRhK/kO48kyP8IlEx1pSg6k
Qw1TF8zEgUvv0Ic2XPmibqCkUHviS6tgwYADjUf+A/zPYZo//66YQbny/5a1cMeMorEGgffUtvSO
dawZPrII0adWYh+4C6UGURIP10wHguwiuihKcRz1K0h5yjDcfumeOKdnppb17AkMZIkXI/+KlQA7
yukgjnf+5Eg7IqzouYKIKfK3i3fCy5WDAaAjLn3OvtMnCYGOWNIqxCaJx2vzff4vL0rt5dKcYMWT
JQSHDx81by9Q0fzVa+ib638jeXLnP4vBGwxUBU8D1rHJd76M06hQ1hFO7oKRJoHAmcDN0QxZ5h3v
/90s/G9uS3CsejVMMg56YSw+rqTgX5oDa/+CyhSU3vhtjHWO8kvgv5XKfxqVfkKck1tz1lsiEZTd
Cv/wVPy8ziny0vtnL5Q7NEqRrnmlK54tXxxXguBLRxCvkUlNx2cykBCl/4tjFEl8WqptX2iLSRF+
oCjVpUPjbjDTHWB+h1j/RlLbPS5VcQ6gVnXTluuVkpJ1Z/zuGJtS8Tife3Uo/nrVQrr8gWu+GyeQ
97GYslaajr5AxpZKOm6BN2nMunRzUR+/Lrf17OO1TcjJgGIdvanVMlVo6QgTByx3BJGJWQssnU6I
KGsX2BST5avBDO0MaXdhlkhwPTSlU0LG3aFLaEKGW9gI6LCS/kHu4wYs2UyzOSl8sklWM5tVPhlJ
vgpAEbnuH6v+pOtBUGGkiIWEjV6x1YVt5L5FiLtimQXv0mVBeoHoH8mHq5Psam40czqfAM4/zCxi
JQVC+GDlD+UF/sFS4KIxrBTPQauz6bsUuiiUzDylcwzNF7B6+traB4UG7CBthTcf0b+HgjuzBKHQ
Alin4/Iy8OEm/mAvc4enAQQYZ8eiUhiSbEi1uEr99wsJUPQsqOO4puhDwAlIHgZjCtOUsF/q1AsH
av/TE87Fb/Wn5/iWU2DsYm3WN0wwhNldjdw/SEsboAlzP6pF/l0a0Ls47Dm099i5uE00imj3Xj64
MpAnB383C7DfqxulxOPVypJ+r6gtHpGMb28QIz2jcV7axtFOMnZfnql7T2z2Nc/m4+YYeJuHOHij
L0jrKSFOpuwIIusphlPQjPFLoqEs9gWZhKdhgw34gbBcguj19DZ3IPXm5qyQKxxLwxhTsG/Hssd7
NJz2Plx7wXlXyCGy0Q/JYfC+jC+9R/wjA1Wn6BFSG7qu+PEKZfW2B0YAGdEFH4G8WAIkKwZSR43R
aQ44rJO+qP6m8LR9oBxkLjuYOYzRsg81W9oI/iJtYVEg4q8r6bdWDskHhpZcvgmaHfexoggGNqKE
VwgVv5Zn2eU00ARyOa3bhtfJIsS1tifAwyXVrNqJz1wSf7MoQtRLnNYvw1xWKShb8ItcSxz/vjcl
OSv+R+M0YL6RQxDVcKau3R0Od48JGFPlbNMTuoY9w0phLDeQfb9WF15vdmJM5+4LafJnC6Kp7rTf
WlVZ0uXUwk4rNczn/6x2s2dNpdYS3RwsOLItejUmZrQ6oOUeyKnCvrTzTRDLO1wjWoEj6uSPQ0rj
izZ/Fec3U/UfHcCSSyb98rutYPlg30HgB7yRy/rwM1MzEREA2NHGdmKfJJrEN4SqB4O9krIIH0K8
3CkG5GArIcC5sn/FxzjvdA76iXonDIYrUKvSjSR9kcnPFqJlrRCKzAZsC51FCkIRobT2+7Tgaer3
04zEPHPYEFLf4mTUS2GAPBPb/ADU1GEedDcDuZ7CRK6Os/ySJRIo35h5s1jac1gIwkXMQV3Ig5FK
jSLZimK94lc3LkGvy5Z80EqvNYlMmpSizVc2VW4ovYpEaQz688c/mTqcZlwjMVF8a9Fi/5K+olQz
wl0nMegJWTvYPbu9JVLmIlx6OhgYFEYtb1fGtqbPhcsFX9nUn8KaQ7DoTX7lb2F/uUVXMmz31xPM
OIUc9xhf3PJuOlySuLPrXMsFcQxfYF0cbx/Px0Lw+M/4tGQQdSNbs0OXousO6I8DvGAhqLIk0F6i
FyXg5pY6Rf14aHswWs4lk3ZG7dKCb+fN1pP3yCWDNXPNCaNrWcmolxKm7pM8hv36dLxMBvnsPPw5
0p6XvxrO6wTO6RHJLh7qhLD8Y1FytV4oqI+Mo4k/sy8yhuT9BoR1r82UG9FBKRIwEHCL5mDGhDUk
tP+GQq/lfrY4KIJkAu2B7oJfrS5Sjq+nXiwrRBbO+rHzeAPpqm5N/nyQjuvz0GoGQv3jpg7tf4bz
3wkJSw1x7URtaskFKTF0HAVPi8X1xrFenDWIanhdeBKJdWTouoIr2nPrb87Ce/4uqN0w/w1uUXhe
yUluTnJDUl7UnQVnWGSvb0Sz27vCl6h2Qj4wzcR9rGuS0U2ldQgQEy64CVNSTyoalVmd8XCwcJRY
tf8Gla56UhmHaBHkdvjvE4NAlwrBHT6XXPyIxOnmJBhxx+9ucE32iqNLiSbFFQqA6zKSyRQUZ1ph
doG5Xu83fU0kWnrfolc6Qf6Znx9eLSukgLvvz5fjU5waMysQFWHh0Cb7dHnXkj5Bb1vKeEJ9Lx4T
F4e7wPxGNiMrn5KWejBYfwn2RV1qoTIIKeW2x9n/kASqAfkUhlkNdAtPedw8RRj5BvRUbKoNhPWG
5bYXlWJ/aKnaVaFOpKbX+uW0ncLVrA57dWFGeguMMeCo6UuhCoSmt5MRggnqplsQSUsEIbIj7LWO
De1rB3F9+25LFLycyYFyKlmA5NDXK5iUJ4jkbINDwMHFqtGsptUPrDRHVvTyWKnq3Ny1aUPkZWYk
ILiJhq7up+ppfPjRwB/uGtJasI9YUWlk84FjMVmL1KIrRlieh7hu29+kcf7NTRRWUuDhPC68eLho
+VFPNFP5XIgUTYiQzgQhYGvkUhTdT9QMYh02growtvXHWDodnTdoQ7zC55yKLAko2oKD3b5dw8NA
cElLdwqwL1GF/oWcwZgZtM4+iu3DxX/n42oJQ6uz4VkNcKCkG8Hj2xpNyOuOvUKydLaoKvLPZ6gN
2TMNr/o5r+a8YiIggbk6vJPtQ8K7M7Pwq/wMfyQgx0YP2KPcy1hCCrp90wRRcdOTe00T233pyBjD
MELcLk6atIPVoH/Db+puo5agsvuCPyT/lhqktgcD0hyx1U/wa74VvtkvdCKmrAISn1REuH0GPjup
oAjEdgBmvf6005d0QelvfzXXBICyZ+i/n4tTcH5oB+hf6do+L4MguzQ6SumVkcjMJugJg2ZKM+sn
VxVwg7PqTk7o1EQg06E/hsYmqOCGojV8nPuNX629yFkRqU3azSbjUFCVyRlIc/BQZ1TOWSd2jQTI
In5V4GsGxBKm7bsyXcWacisWyQzI6Kn8alAigjdclR1/YIuBV9+/znDhQwQIga8xekunosA0p9bk
bN719Ali4oICuIIaEZU4E43e0IK+fgrIbTsIzGFiaQ5w255QeJv1h2W9HNq0Gex8OstRogKMSh4w
I4aTSB5cQ5/IRAsD6XIoxcLDTbzeYJhsYKhnrXZBl0Gu7mjTH3sQOpgBBD0LBI3/OjveMgN9LSvu
gyxd3sHNkZ3O56NGYcCIszraf/WHOysIXll/+an6wcYeJX9NMXAhT6kRD6Gcxeqig30WFs1EcsC2
LLeIjnv4j+SEuUX6fSlTzWO6TPvB36evI/LN0SnJYEa7NZh9C40iWQ7lz+roZ3pm22Pk8e+4fKLw
dXft7VQ0MKhlveFvU/smUsNDKzTRri3R8Oisx5doAhVjTr0py5GhR+GBvRgYTUtWub6VebJMZjkV
p0+DtYU5WRYVGjuryJZDJ9K6A3fozcMSy6hCb+s1MiPhIkZfWPcxz/XW9O6zi+8DjfP2tAhhmgJw
atADC4o/O4GWwTNqh3yxn1jkb7+6sbBSCPIZ2mKbOyH9NuOwwhWgpIyEuFiMrBdt2W/F1nSKaqIa
wWYtlMpuI18BjnDOc2ybXAaDYIICZgFPBEbPRlSPIS8YeB+BiTTXvAh3NM5ulu2ihQ9++/SluQR+
yzFfJ9a+RgVib+jpbtA5oWJmEWyyIenf0rmzWgfBGJBjbywGQNVNQEgTSrDwEvmIkht1oUbHQWH9
3U6d1dUgaa+HWX3KcW9Lv041bHa6m/wCJqBwSeVhM1D5n6rgCPoDyziiJMGOHoLPDO4SQICTjNpy
koQ07bYB7DX/8sbamNPSwUMhy0hAWat7QI9Mvm9pqhYiCKs7mW3T1ckwzZh2doaa6SNWHWr3FC49
HjTcjUN7B6NTuStAS1Wv+q7/vz7HYkGYgX5jEZ2UrYQ2ES1ry1oXYmNNXwZSZRbI9hPGDKeKf6hg
XZdVuCScOSqMEThnSWRMbHYN155teaywlg4Y9dwRcK1nvStklgrFq8G3nDZ45M61yQrle/FzZhpQ
guYp8Gf/cEMYvVp0r/ZMsff+iU1OVsLMfR4gkxNOyqbHfCklFGlCfNY6AObOIs16Q78NmdyhKSi0
jMiXsfBzdHXpKLTbip6uUB4uwmW1zuymLKNsowtjlnDtpaiQ/y8UWjUaW7QprndY7ttZG0k+O9D9
cWtG4DZmrmEyJlU4TyDzbo87sTIrDktGNWJOichPnxMhXyrlB1cWFZQNQsywEd6jjy3gPxpU9B2F
vyGUHh495XT5EFVyHOtqDvHvKfmkjACifOluI1WLk4KW/NdMa7LQ5q7uN4jLwEQozIoUK2yM+Tdk
Bj9LafHChz1HGVfAi229U4UpXhQiyulxhbllaF6UD8k6dWSQc9KNvGLrdVot2joyXj/I7d/tx2R5
aWbEI6X6UB4yJGo3EXVeKhDEj3Ztek93RdGzDTeUO/VT8CudwtniS8FMwayOeqJFqrle/SlhERQH
OPib9L8batiCCZEDsm0il+J8PdaEH5oVZQS+qxFuRLeye7B8h3v+iunbNKii1NbKfhkm3m2HGY42
fntmjB92YtgaOQ8dmxD0hv0SRXh1t+0dfdZl54uLmIzHgojqbEFTycbUky5jTg5nSq6Vp4TNMvip
UzSlTiT+oLbnFrHIjEGFHr9+iMiRuhFSsWLd/75VJ/wnM+GLHOzrHV4GdaCHQUVBOjc7W6PUGJQS
6ctY7eim6nOMZo2azDWEVw2Tc1khzo64SYwFF5/zw0QqtdTO4KhWrGQu7IH2jYzx/r4x9dq+pda8
vTJmZfHUfvKLv1NDVvLqYnLkHQGJdHjGGhtBrloP0Qk/yozzmUK/6RTdj1u8oBvtJT2l3YxJ/5SP
tnUy8v3IZCWfj3v+uT0RrsJhtEoll+1j2BLM+RuKA3mqb6pHeI92Ti9mR6TYejiaMBnU4RJUzAZ/
IVMezQugr/vXwcuyaO8sgAT3795yqq/Ac/3r5+Jn8kKy9Sb2kCteo5Bo1JgF236SqFcuLSyhQggz
QlWARa27ZNuvna5gIt75Gm9ISBTKKqXZyk3P7d80bratJDPO8eSI4TNXlZMDBNv21+HaPShyyjvG
pG7bgv4tE5WadzJLhOsj6GehbMSS49TRXbfYeqbZJwIGOeVuZ9BDCS2BVQVJZm5IGKE+IDVRxRJu
pLO4f8Drl396rRJBwC6p8/tIVrzIUqJRAh145EOXzZ8ZJPH6MNbe7pBCaZkNSr441N6/lmL64eZf
bCg9ycvRjh9hYMDhaf3usxZRNwUgyzJinD7cthxEk7qU6wL/WAxIU6PCvPdrWsqY/cxiRyMx8q3F
3J3Bz5KC5QZv67OKwPpif8X1eAjvZR0N7C5GjOm35J/DSizEDeN8K409pp8P/gt93+urcKF7mMSg
QvYri8GOF15/Ofg+j88C9cnG3vnqm5MsoS1qHNVlHwlVReL2i2j1jfQtp4oDGx8ZKmQeUy0XhxMU
PYA6DJ9jTiJPsUKJkR/BLD7VnSaY0Ym9TfbylY+0z7Lerfmo0wQWkOuIAxYtlQZykx3y9KPPpL3T
D5lQkmE2J6LPER2QsS4xYzsqi5oWSt6vv++1pCCeNJgqXWI/UGqHQH9q6L3/iS2zj3ebNu3rfgEU
xi3HaoVAKZ/dpuz/ss4gGEZftg5UiNWD5f8E1NuLwFHZ27cNeduvUoXa/GJQpoxif+OQ0C6VRpxq
cZkbZ4510mDpWISbhQe5ZIBJRTC1LR/j9Fb2D7bjYgzqEqW9edXdYHQNXj5jKSMdPKcnEhPLoGTt
vW1AioRVs3sM0fTP0oAZkZdowbNkvw3e+czG1Iufn670R1x6H83BIK1j9AMRLctkn4Ej3uHyg6op
QemN/KNh1hU624b+I1+ijQroGN5uy0uNSpp9t8SmKOmTu5d+Adw5IMSWdSQvLo2FCRSNyjnpUFAo
gLGO2zoSLCQzOc6ZMdPxY9z8gung6u1I/mRZnuroH6VfQIZ6hcYf0atNs3HXd2QsLc0yd52KWV1C
lOpzirXqlOUkCgnz4WBEt0Q6yk5YQmRbjk/L0jTMFexzRuvOd791V4zjGVR7Fqs1GM7boKv2z7eZ
C5P5g8XvdC7OoIFK22C2VnU0rAk+6C0eTTP3UHivrxs16b77k2T4el8zsb6vCPVw51X3L1wfxNBM
Thwxtvmm/z4h2WWf7YR5oQIXXdeIOoPYr729mfcD6vT3M7VfVJT4LdAO6WB5uKk+gxczZ/D0ouaj
+qHGIHS4HAYZqHdng5sa7461zpgjGQDgpP6rHZRefHrZZKjwHIVu8ZiBdPGTgqO75Ote1fT3Nvud
LbZ6A8RaCgUupqk+D824oNY9FpHkMMrHK2zMEszKPef9S5jaTQccn7yRaMaZ4etqf0ooxpyJO7vi
CrYjgcTV6Y3YD48piHp9ea4af4+GiL37D/xq5uNI9IqxFdy+G0xrosoWxJE2Q6CcqJLomIkUnIIB
Ird3nZefR0qL0vuHZPy+gdzHhxJKjJMf8nZYvitmCIu/mJB8Ok05VHuoBVNfaEpOEKUuE7JSjwqj
ys6+etCQsnSTSD02+yUvtkMW8Mm2Qsj46tqd6Sm0ljPjm3OgofWF6gnrbA57369WekB/exWhOV1X
HLNxkPC3kE0S8eRhyjC85/0TrhwgKWBLGc25elL/YThCqbBAKJurJyO6chznHSBCkLgaMZHr66uo
N4N6MW4X5fGUVStfEFU7GoWcVnoitHZhLTfys+EOSFr4Gp2XEnIyV9q1Xdkk+sylKxC/iW1Vd+ha
iq7z5A1tTCGrPeSCI/Lnyvvan5xjFr4yjJl878LJbZLGWmYUX8Tl3SGUfh7YmnUU0jAvyZ4u60z5
DKPLr61b1t7eQ3DvA5zPg88Q1GxmaXz/E8sY4PaALoxwz9vLlguioNQZ0YZdRzF9UIlo95uhCcWL
L1N+ZdQoR1VfdoxM85ygB4n7m9bKZoOEKF8ZBGn0pRhgScL3UlDyqGPOokAuWEHpJY+jfjki5T4c
5W2Tr8rj5B4agTPXPYz23F0C7NyZzID9wECYMzbIu4TQk9znZs6ca4nI/pUUQq5O5YipJ586Ad+p
TekdtZzYq87IlK36+ql/7zYady415KDr8ZDZQQ6xD4YWmWhe7m7QpgkRnyd9hCThqV9USE9UE5GF
uIkt05RqOAST4vR1D0QbofgmXBZ2b1P0bSBKGN/6iwemu2tJQ7s3YlQtjOfkjKgqjlIjc1abLliA
+iQxMOJGi02CLN3cinWL2k4pZERBuuYBcsGwRm/3LNnszbDqr4laS7ikB3wQ5Yqx0v3EiPZEQAC7
iXcNRs79WMM5rglnUdUp39hb0qeaN5SD7CyNcQ+E81QRQKVfIsfoMDN15e5sf38+Y8dB93f0O+5C
6fl8Wo2BRsKO7sFHkTIbYkC3u6SkdfNxXgyBVbrkVHgyAzqt8LgFlGEs/d52L9wfdHonAR16U5AN
XAsE6P4C1zWoFF6kRKLAkJ7VOKdtbUwy4eAPPUVpbKl92YCFpBjlBPDUQMS9E4qwJ56Im/+f6KkB
eAAeAW8B0jQMSSP5xIbQokJdiNyXCnAT5g0THpDYMBObWx8Y9qjQP3OFLLnvQv2KaX/clKIITr7p
95JIoBEI1rIcdSSEHVT8YQfGhxSnNbv105Ha9wdP8nxRrE5Ww9XOsh2LlPSVrWNqWOHYAQf6tADt
s5DGwTwVIlU5k8RAGkgVolc9uBpLszKxTC7wnZ1AIunnbux5VM29ck/pZcdPiYTMvoNRSpZwamCN
pv7NdmPzOfYmt/l4ka2DHbRQMl05BLZpeR4tlKbO454N4NmToHGBob4qbj3R5lGBeO67SHJmaTJw
mghyAHsj+l+WZpM1gdRWEXwcryN9FPgZmFzSOqWlkf2LA7YGkv9KDlllME4/JAWG7HdYRJKTJrCs
C/2lXS6g/YSUGS4qTFvE+7XG4k/yg8S8Vf34d8rz2wgMc105Uxfr/Z7XyUtud3gOmrydGMKX7YS9
9vtIU1Y1CBPsaTTZ24if/kuT8EWlBUFyM6zJlHCCRTyFbocCT5aqPyNavW8VL7Cc4MD4TZvMrxcu
hUnVKkO/mgQygtR5Fv0POBdp4hzDlbdcgm3YGytNBfoVDGvD0lW0o3LoBjGG393RYROXwtIIliPO
oQ56FWfqJ4/nLXu7d6I/fE8f1sMFiV9+XRJNAUHB1JP7A6tgr9wZ5QOthZcMG3l+IsTAamKY4TL0
0guZ3iWuYPlpeyibbJqt11Qob2UO9PRNzuDEoI+JzpS8Je0kz+GSd0i1rDrhKbeaX/X3uW+pnNRh
Ccg1/BKffPJcC00wq135lsHveGhuCxB3EV+AOy7Le6q/ZDcyRwRzfjO3icTWwkk9G7aMLDhernuZ
Be18jUMQsUyYR+78/qAulncz5lIjlpCimBpVOFBfDIRVtSmzpzFXceRdorA5fNPTRAjeKpl5Q/jc
JGZFWgP5H5jcY8zwu54g9B0KhR6LcKor+SO4dusHT2RiKGz9Llc+9inJ9unkLh0cb7dsY8WJwb6a
PDCFvcjlc+OQVHJmYXaN/qWb3uCvrl0c7ms7NgQMLdEP3jo87h93Q0uBb/qy4e/Rlbh2A5hkzbay
rZjEh+bZWOC1PhwWZ9d6ny73gID5Kfiv5xfxc5AHajZB3cnyHjMF+fCzZAAgC+IuZdlg+CdPoZRE
uEHEPjpA1McpoNCRfyOFXSAPW5x+eRPtoBbc/7+IokZ6+qVwImATtjoQyJHIe0FMwNy+HkaS74sj
T/zP9euTQPWtbGRgnGD5DYyr2kkkaMYHK24MmxyT5KHunSMRB8UFYWQsgZp8ibIr46kbKcL+N0vl
DrfepyQMXpT/v1DCGhx6iJX9l/tXfYREJEjJzv2nO2FfEeXNxPyP0ofIgGgs41H0Nbdoqtqc+SwU
h3WxwSFRiaNubfsQAwSHSRc+/FM3KE2CQHxsh+hUdcOrFVwH8ZmSoGp9PsAc7vNX+C7VlgUoVu6O
INqRrsY9VlEbFQZcBLEPqsIEpmspmAhilpa6dX8uBG7TnV+q8W+6OOoiAVMrNdp0IV9y9GJDtm64
TikUK6BHvwfsNCorgwWdDOuizCa9gG1Gh6IPAUJ+DBP7onxH2qFprPJL0AdWkaUVTf7VA40AyJyU
BQTWQ5D/CXBBUOMlMg37WJpk7u7k8y+aeejONI4JgAtlpC6M91BnF0DP+68h1gPEW+ZwEj8zUZPV
I8kEddi8YmiRFNJlm1Qhs78v2rX9pFMR/gLD1tJJ3RhNnV0bqWt9ocevDk7XrpDPQQZZXQX/fcYf
3ujA/CbgN1oWftFBe8nCq2aYXM8nR6AiLRpQmB7RMzAaqDY+z0dYOVr/jQCJAX9B//AMEo7b2Zxg
aBAbn5CzqNLemT/IUQFC4X1YNNja1/57TCfChDKKdyvV71Ig1xmAQWXCv2WgXPFDmDUf+io7OYq8
1//ShPAz3a614QSyO/dCj5vn0tTkFfD8cVGoe9ajx5k+r3677SD5wtmAcr4LA/8Ni9qp8ju88gYT
n/VwmilBPJHrZH01Hblrng8tztTTiA12h5LcGPmICs9lLCbWYtMAqZEktwf3BetK8E5Wn4B0bD1G
dJC3Jeg77cy6rPmCu36dlHh1BFMrDTeZGGc3nY0YQaHbEW0uk1BXlNQiQgxlGhQQ0t+07z4+B5ZS
U4JxyRpVsv1g/tBCSWtRArSFFqaFhqtr1ru6Syr2iElYTwdX5bFgb+WN7eeDvcTEvwp2nnd+OxcT
ue/kOiVPHQ2VnuFO1Q4glxthXuOYDOsWMr2PgHfNq/4G0I2UpED3prwvoMyepgosjVsBVTHwYSyc
qRfbpdtkesU8NXCp1pcQLOZpo1tJFy57DiwSBTC/sFmmvQPpzNKcoJKG0h8gF7oAtCAiK5qL4LPg
cYFAoDdPiW0EqfN42sHKhoe19LN2PA73Ko2u0hA0ftgOfhBjMh0mO+26tNLVmQB1Q7WudZtQhFxQ
9BqTmyBNRBSmO+Y6z7iG34R0eN0C0LwmM0x3i/7etGh0GOxqRFbAVh+unV2+a5GpPj8TnkUZqYNp
t6OSN5uusegd/UZOElr4OwWC/XlLAm0IJHgNmCdM6IDuXPqywbDyU1qhoeG8/7hTDMCjElfL9IaG
Sgkp41LnA+HZXk1+SBWnJD6VKdLLD2Z3HaY6GQbBkPbdvsz3/lcdjHwF3vx4Mj53J56TWjBS1OzN
w18Dqnno+2XqvTIfeAdKIwaBZxBevYVkhvsTh9M0aTCOqGu6tA4EwfK543PY2XzvLl3EPUzXu00G
JS2E7C8oSOWqLaq4ocWqK+3Eds2I3kU9HUype3E+UXLv2v0jfnAQy/7pR4UdZDd6JDkShOBlQZA9
HxRnPpGsXRGDJZLelJyt6cUJT9ljzfOHdNLHvv4ibUe2+R2HW+HJBuGBq5JCrxXNe8r8fi/xtPHG
xK9/bnfoh8tC4cY1eL8ZXUX2jMdaB4c8Q7o9BrFmJ41paOObQaeNbAGitTDChKA8N5BFmj6Hb0nr
vW3ThKPcwZ11JujnravkxBKttnQJ/tPqcVpQphMsr1eAKzfdieMLKg+lM9Yf3cew/3laAkKW4XrL
yCF9Iw+fuy3KV9oiPbMG99e+GfIIfRGT3/IDPa3gfYhfseURutcWZ8X370p1Fd+NbLEk0IMAMnft
37qL3k04og4+nav3F4wb1lY9xPdCIpttHpiyPsQDLdtgRTdKAA8lQhekGERjp5QIhZPnLGJ5ucBU
i8Ymv6kF8BOXks5NwsEV6gGPxeZ5mvP2cqjQYGIj+J3G5cbTP6DYmgc2DqZDdNIJkOaHkO41LKxS
K6ELI4ySbAgtcNam6gULrcIqAnO8DRVqSRLa7y6xG2ZyZ++K+lMLp71J6fDKxNayN7lNEHEtF3EA
qLy79ulRgoDe8E2m4mKSZwz4Pmbix1dU8pwtpMWeOf+fjCIdzVmBLMls7tNreh54XUpoRbxBYaso
rgOzrQzpxubURJ7tjIkykubPX8yuH7TPh9cfnsBkZ1S3Es5YnSSvzYOlhorErntpAIbqy9Be45HJ
XSXx7l7BXmLEselrZgpq8qUWEee1p23qeQFjaDz7HyMFsuTH1Xd0fd1EqSC8O9iNRmtbvwHMDlat
8ae7MyHiDs4t5G+MlHf0NirS6z+1Ko5AxCtBPd4TbOwqtwYMUQZViXaiWBoNW8WfAQG0ZKBet9O1
f8QvUjf3WVg0pQYiO8K5X8eEi1ousiMPqdfTPY5JmmhqVyeK4mDrXBosizJKORl0MRFTC7MoQ/Yl
Jn5rFcRk/06vdnt200Zq2DIIUkgESYRv+mEWBbd1PE9McM8jnohl07cui2Strs2qkPQpntezR7AU
EvtQRR07Iv4ZHhofoOQmKwRYAc4fs9OugwXQG7oq0CuBhaIWicIJb52aPWva5KgEpDXHsX5xxnsk
Bo6J8scd4hNuKqMhueaonAOPLEdEqED4+MUHJgBU3oRxGpL79DICgGoTvFazhRs3V+NgA7teSKwo
sg/9qqSwG9EZB4jgCr0lBGnkAm0m9KONCqwX+qNtY26Xak0Tmfwc+JspPUwhkkPYGtMbFZjjYxWr
fpVmMTvW9+0omJjwz8NI3TmpR04hXHOFHgQcz/HhXk/FypU/tvKr6qV7mvpar1NmoByeClvVobL/
1SiSUXot3nUV1gVE9NNqL3kKnr92TwkzrQ2YT8Hzgt2mIATN6PPJqIPYE6es0XpEs0/38BLT+5YC
08MYolWMnxVIdfny+PiB6hoetZFzDsXmsobwsNf6NQ2NbmMziM6MHpSOqk/BznnGFuK57gksXdTU
aWk4vks1pNURK2tesIW1KzgvxV6GcFH2gUGbt0YXMzYF2qnB6IC5QfOfIh/JowZwDp0iegpK//uD
fkefZfJl/3u/+4LWzcyJMJVkWnca3LqmvCBMnkWyygGapYFsEICLqDW41+n2TIIT1uWlpCvtkVIt
po5gl07PnuPMMoCL6ixglsZYmhrmgBf/ipri43Nb8Cevz8Q5GFk5onkmS2ZibJk1gfq1TnJ0Oa7J
S8Ra2+YPOWMlNw5p7f8DI4lgo/MbIvEVWO3QkXyX7waFkcrkZDNrdhQ3zJI5nj9JKiPBsylWVUbP
VfkQ0c2vcRgYknVuzFIFMxtmghe6buYwUswMsaFSIJCU5dfYq9gHBhlPnfxkU9ZsXyXvVPDFHh4N
ze0b5XhssYexi2f7Eix8J0IcRLNE3N1CwA8rjtBi1iD4ew7h4HPlzk3x4fgMHtga+7glOYtyZqsb
WSHJolIcMtf872AEH94/KpYnMBGbKkrwqb3uGaovyz12fDu4IsEx7q7jmDuKyR/5W0ZDLYOoJdlX
an0wo5/MzdAXBJcCfUUc4BXo2LCSqOYXwd0gLJJxHvXqWRZaLRIVLl8NrfTEOc9P0wPncTDmFfB3
CIGtRWrvctFYbbxmTgf1jpR2h1F4PO1/MMiSy0IW/qC3k7A9oC7RccFKmpyq1pRkGH1831YpinJx
3IlDMumJpmq/B32AlzBLNSr6HjSUS+RqnO56DcGnNOoJmnFXQ6madpH2AcCbh1OvproUhrZgUiZF
hc7t2Dlnd+V/JHvDx1Fzbu77poOLWjPA8osdaoNWpLu/50oMhToM5nsPd9AvDyMVv+7GQLxs2JPQ
A+GMGlwhDmKJv4teBCSK7IM7fa3veEmlztqhQhpQRGfJ7juj4NbQqmbRj57fEnE7Fz1eCz6+Ww3c
pzecgT3EqsyrtkRw5iLh7JE6OGR7wF2v63PVx+HvPA/V04GCUuohCS23kl+a2GCoOm2GwrhPnAds
KZrwmIjpEtkjMT2Fmq2tAMFruQIZwhN3hDaFob3Sq8OSxKLb09yor6nU0a7KflfHdqD5sRhAhEt4
bGed6+fPcPf1rryhANAmjk/sGa0Mwz/G+FCgnTGPb2dRliAki84WI64EZ/vUayu3fCsogLs2PwAd
nQwl4BV4qxv7i/HPQ7UReWCJs7YkfFMrL7qvusky82qj9+LtYgQxYm8sOht9jop2PrPO+x7rAMWx
tNQe2bmh/T5dAWxdElMbdJyfDjUo2T3A9M+rrs4AStfRAq7928w5BDvHOEJsNOGqRNhswZoes2OO
v6EcHF0Up8ol9pH4GsMYuXXgA0MKlFjuiuR3tYZkfqOUBJ4f8DpKm4jeodThgiwBdPXss4KuygCB
2Z/oNFPEuUlaPz5LDFZVor45YmEhgU9AhBT/e2F3vECWmjx/0UvOiaNJGhHrEheB6gEcE/y9NfIj
/dfkXv5uEmGDI4G0ShkMJKmzLAkFB48sQgF5R2LAF5OGbXShOvDXfeU+BYv/sCi6KZQuDOFkm3S4
dDvhdy8vpStkSEXBjtWUgz7VF0oNPG3jnx02mviAr7ArnJtAI2TUUi6xNHcDbV7BXliXPUjmZPq+
LJiJey/X7eejsSQm+wgxTmOiORJViZ7urku1Hyokq3dz5YRgKNHZVB+jMFdWqcWnNleTilCMVciZ
ctoyWmhuD/W2CBG7gMKzgji6bJ4uF5PHkKGX/CKriUnyvgDA0HB73Zmi1scgAKEoOXw+yPpvjPGf
Em4kCUZJFzsEYck5LB7hpSyU047GWqLEKM+N38OHa5IGFW0kFMCxiRFE7Tli6BjAiv9VPE4xxNWs
lHmAymOGp3dXI9bsggJaFbk/5cP1bVN40dbaKZN74hr5B9i9GmTN9ip3bNSDMMSSDaYwGv8QeLC5
akwz5JsIWsPNbOHUWzXgqt65wflRf5MtRN18URCOGwl3ZYa6oa99JiHLU2T0AOdhCjQDS74cFSdf
tbvUCwAj/vBm9UIjn3fESdmNC5gQ4sd3kiEccqdoFdtnBQ3zJL4v1w7CwYid0EHeJyaO9nz0ffNo
r51jmwo4PaJAuMPHZ9dpdc0mY/CaJyDCVTepBEyGzz6wKYoNRzduhJBSkSnJCRlat0eWa1mwCkrD
R1qGRECwdOno4fFyUcv1MGF6OpNSMah6wEh6fUit84uEvZ6FmWmhi/bWO+JZTxOoNvRNaKphXLIG
ER7UQMFpxF5k3g4WIng/BzwWgE8nCXyTHe6/FV7EfmDpfFP2w5m/30BTNrRzrc7TSjbWH2adu05C
YcubPWPn1QrWCuoANRiSLvKOE7ECMR6/SK6UWwqOUEVOoF54jZT/EKimwrT/nJl4npGsf9V/zSPP
Vs77ZymOEszgrlu70m7vWw+pY+SdDuaskZtnhAFB/yRDi8O7Y+8B0IDaRr5cpLmo21k/jL/zG1QB
alJ5ZrabLiVyQNxYrs0+Pdz4MFtwOjYiNJiMhEtg2I/Zjr7pH69SobI7qMsTsinK+fKD4sJqiFum
dB4sJvpB1JQlsBudGp153RtRp+kO36Xrcf035/HvXbXPrmdhEPEF9HZVqgyJ5SqFYNVT9tJGSJCb
q1fvNNY4lIQ3ShLfM2rVbbg2JVMaKGedHdSYs6KVKuY1lmOrsUoPHZ42DBOt0hdiy5oCUiWn7U4Y
Cy2pjkAL5VNCCcppdiZyqatRAFCl3br/C3bndzZDzEATcDJfLZG1zYVNQPnfLed2v+Kv5uOoMEM4
PDpUtmA9Ud0CZUO39pKxf2js7/d4lwtxMozvJMBZFMWkfswrp25lycLf5053YHtjRMJ4ZjYCkfdW
vND5JkwBNSeOZXMbm2UfQz0OxpcILGHBfGAB2AlFOfDEMcc6bdbX4OM3K1Xa/C2KS8t7binNK91L
2kRCAuI6EKR4/SkZ9ClwPtFcPJV63UAWDVCMbq9Hu7f5Ak4Qds2wnTYuUauXPBwsau9tkiA1Lx1q
UTYr5W6t3lnOSyEG0SOrhoSJxlTFC0RvA0sDYhstgQzP6ZDXxp9LrUh55UB2vIwHzmL5D1/CCvhi
JOjEO5o+qtCZ0y63VMJn6rjGv5CmdpHjHClIIjGzV2SRV11/BwBmkfvnu80dZnhwp3uZ77RpmzPH
BFPLXvVkyMrfHfIsp7UpOfTzw8hmD/4FOHP+mSA9e3vFn/uTlM0M6GIvIQDgrG+E2XNNFt+v4OYq
Z8YetkH3aZ1ttctNzNyFOpjdCt5bbaXRxIC1VWXdyAKmFx7rPxvTZOfI6l4iNrEKYMco4y4ctQFJ
Ts0ceqUNJcRaMVpQDMdY5auxkVatfqLpGFKs7cRFqfYszmk48iIa5ssK1VlXKsSRxX0PwGpc4x/5
wz+YB1yYi1HpR5KkRrFAik/GBkQZ2rc6w6kNlnABZO7hwKXJFPhpQlcH9CvpQze8qlerb/Ypn/xv
MZ05oFPg/FB9ot13F7fz5WXE41AXRrQm/O3NkeoYqm0AcB6xTt9YimakzPsJ/4RHfxHNkLZGFssm
A5G9d3cD0+OYIuj5Hs4KsShwWoWJ9mf8iiwmiou/9M0aUSeKla40+H3/mbenvgd7I2WbIYFbIraK
CimpbICjv2j/P6g1ovrvOjP8HIglrL0Mrf3jeIwgQN0GKQd+uZdFPrsFZJkCsA5/j/Qy9GEr6iuO
w849Ufb99ETqtWm0DEarW4ddl339MfTon8yvJ8v4dvCQwDVLY1KFtPsUEmylA0bxNG0/DojJ/t8z
cLxUEW8tkpnkBX0yTPRjLF0zWYdlHvB2+RjvPsVz6IoQcue1itqDt7mz7UJEjDqYMc1kG1m2gWH9
+E79feeSiNssJ3dlEsHTr27FZtXoKHP3SU6MQvW9fmKb+A6zwpn8Y2k+93MfCos3IvRhshdAIKRc
qx96SXPHAjrUUJRkox+0RsSD+c9rfLScpeLXSJOhnzLW+wdRETYUozuau0RiGegjCOYgM7PHORbW
sSwiJBWRNDZyWzdgy7OjU48f5KLXUW3w5bDt6+yjZd4cqmEwmRmRsZIiSLHAR9LpOAsMrNOoyas4
Hxbt92z3CTM+9KBnPtlWFW9xUQVkYXe6eTqVzI4mA6VKaRgUQD/5fatNWTrEEXmaUXi4lG96/zVF
+AfyfV0rGZEphDDfj+0MhEMWoKwFTv5aQSkVGzfmnjcIFhS5B6ly+f9m2qktCn6vTryZyEtBNvE9
YPL8bIx90sE5Lb90agyVZpvPXkKUpHpuKZzgGunw7wmLsqrpu1Kd4AR9KnviVHutgy7O093S0+eF
aASzToY6RsK1LrCBhxMy50kD0Ep6gjKRvnWtB7l6KGVRSkkMf/lC7fUeuyda9u5jYXIK7n98LdrY
EaxFJaDf2RxazL8wPqOviLIMb5psbEB0RICvnm2SA/e/biizKes8WVQ5VqDlG1m+9GT4CQ+ZsCEQ
3hV1F2aGAAvCojIvEChTzMpM5v+zDDpKjHDizClB0tqGjUiSyGnWpxmjcAzI3QMfsslNsP5Otl02
vOBDJOKh+uC3BaPB8GuirVQgskcdElStvqR8CW3ALJUMmGkmhOqCWDINLGxmDLNU+74HPga6YQtE
W8o0yyanj+g+/j3vh2eg4IWgz+G1c/8fble060WKlH37cZiSqNTTVfOI+0sQGhQoSlALWMqVaxir
Ue9ZZuXsh//PNghWdH1Nj8NRVLq7ONg7pxnPf+DpC0Q5rRpClMD1Gpf6hfwFvim0NAVoQcJZ99w2
KlRd5Cr3D87JxfOjvOwUZKqrRRHZdUcHGG2JfKclSac3vG4sVJvrMzpnhH3OtMLvfCoUnXbfSo8A
6XGilPomDm+yse2x9ecUanwjECR/PFGiMNXtOzmkFPtv1gRFiJGcXaRis02Yls7XiCXRsdeI0zFO
NZkglkNIS6SPPsA017OrBvEsZQhdpDYvn9mHcFpsBXBTLbyaFM08RzaokVJJT6KMNSPWU9LGSBsJ
g6NZTZ7bDRJ+8wuR99C6bAHDtduj5YoOr4pztww9ycXjtrQjZS2XuQPsaQDTZGr6lJZbtgahYwwR
bKjCi7qfKyX2W9Y7X1GkU/0kpCqAQMGm0lpHlMChY3zT14ccM2tO61KhbZR5PJpWy+A9wO8AxDIL
1qsGemc6yfyl+azMmo1d3fCgf4B/vuKEe/ZaZ47HhGjqEI05Z9FfGopYzaL/guktZmxdriE3cKx2
uAkSA5HXFtqC8haL2ik8USp4U9osXK+jaWMicid5sNxdEW3y065z9gUL/qLyaIsSusP1xXZ02Wfd
J9xggAALNQtSDoKTy588E2KJzMNIPAa29CuWpLsB0kKHNhfQZ2CcIYzU1WCX5sgvW0DsDHCcTg2Y
yHZDmv3e4D8ZTFR0H6cRpjWV/508H+h1gp25aTBASpAUWH19g+lqtZLtarftL6eWdoO35mEZGCsI
rpBVWfBfhFYeuGAutyRHoUGkHQ977bDQiUT1b25jqOfAUSYqPk5CUx9qTwIUiMrs7k+G87ijOYSB
0MS/1FzKpyUphIOVm02GtNC2ES0yprwws8j4buwdDOzvhA+ocFQhN9dLRUVppX58lDNPqZET2nB2
qBldiLxwmTNaxleApBuVjYPojGouAuc52oBQMS/7IG+oCac2iNDbezFi4bHp9Gmkq6FNBgjFSTle
U//khBAjB7939+r8JDg7HkbbLZmNhaJT2zaMdT5D1XHB90G5yolDvR6R2eL94K+QruCqa8Sd81sI
P1b9DDQozQEqX3BsPA/2q5k2HEOXB5Y9fK6y1pariTCeSz9U7Z9h8ZKxm+q1/pPO9VXEPgwar03g
Q4vzg192uEElGUF03OVFaW+VLfBPqzQrNp3EmsODcnIL/hpSaJ9GJo3aF/u6TDMond/0BtFcIO+3
o4FoVioV1JZS9G7BqylATc29MMrkb7IQzcNlFug1w+N8itEmNxnlQKzuSPlaNrUxj51EszdmmZQ2
N5LNoaN6gePb4/XpyzNv7kYZ/kBf4vpHpq+FnRbpTkayeBVXLtYxRaVLbuTDJ4Ze0PrDgew4L+6u
P3QY0PY6EC1ge7hCTV1BAWVyz4xK2S9DXLKI22XPjszBiHlY5q3nmmh27mjlrhGrGwQ41ieFjt61
WQyMROwSEdFXVSoY/UcQyGv3wZzt8/Jgcs3cJMwBjizUo7xjUZIOcgH3rs2SiEPoqQZMqG9AfE+I
4TTTnvQ9WalORalJcpKpkVTtj8HFA+Led1HJs5HCHvnHKqL+aO+I2YALcukvNlBRppNzfO2Wkg7o
PLt1jk8VH4Dc/9rRtVGh18TPuE2uIB9S8tKmtpUe0r6qmolS/YVlHMfKNdIT5AtocGG4IGmRrKJj
IrKsZUatpUpGULKhJngmmcI1DU4AXwF4v0b8PAns11ah2+rVN6tRxOTTjojL99CwFFFpUs2MrEB/
CfZZSugPNI9gEL70sX+AlCzFHA0Ybbhc5aO4s8aUS6VeevifDf+qu8kBNPZKro76xKfTLpzYcos0
5AyBQFnHO8VDgtmpXwzqQSKvDlouBnIa03nsd/iHlS+saozAQ7Wn7RCDify4xMavu74aYzme+REI
5qDY6LnoUE5woINiBEjeqccIdKLjj3J4yvSXkJSLuQKJLaqPFdGhG4ODOm+3kHnNq2aDMmZRwkdG
7m31LGDsYPlw3fQ0ol3pkGPgw1xJZmVkFbtnZeJLbHXAUXYDB0E/ksWz/Z84rOIn5f6fnfzsJF98
BNkaAbSVU0n55paYB70c3MF4IBLGVw72hcgqFH359lMH9ir1qVv0/R1F2B+RRgAectGqGF4A1LjS
1V0L68rkzQK0BXGyl1hEvbvVPiXRlcKFYwA3cdq1ofcuJg7Oti6rzqCrW8ZQ+JETZqd59gbT6GL/
oNRtwCoQS+LDV8Fz9jac864trlZjaGkFwt9eAFkuv+N7Vqv2bYt7yh6fQ6NEwIu4GLAGBjU7ECL1
9cn7IdXmYFMyFHF5WbIxCc8L9fMQ7LVDjleFpvM6KhYCkG/6Q8u3HVDlp0bNwKr7ryIFbU2eRgPE
Akpj82Woy6TIhx91JpGmkhI6jv5RZhaAzGH8dLHpueMlQIZGvx/FcuR6Eq/sODCGFLPP30NGJAwY
dCWfZ5xJrDm0gbqLbuf9v2VcwVdrRfxByN7lOEYbvyGtHQgwdO6L5ZcTYjLitZ+/X+m2kFvqDqqJ
ca5N1tqiN1QxNuntRp4zoTZh95FfBlG09frvHKJXyu3POKj2Kp/bB2dipMiUFP8kfXv3vVod6gJq
oRn/4yKVHSpNFgc3wmo/SFsIJ6+ggXT7oTZKrE/neNQKiGNPdKbbEs3uVgfbxnTmrZptR3TtrrMx
z1Myf+1CmTjm7XuFsQpcAAUfFQudh6wPUcFlq/2S94IfdcMJNXqW4iIF1lZVxdRxTdkowo7kNyGa
vJuKloqIfSE0yP0tDgUGaiLuQMnDQUJw5QjyfNwahiD3vFeV2bRqLVMj+EMnLr/myWA7x+z9rOp0
pT+A1R7Z1QqNVEGMnj9L0xhWy7Egxw1CBkuf9agnsdWs1je40hbMgg4+RGaGZ1wjvKpz6SH/+fMz
qL3bbBEQcvXK468UZ2TZ377IgmMx2SLEdYgwFmvNxg/I3rK6Fh5XP1WZS75fq3YqiNlZo7xrhzv2
TcSIUF987JY8jcg1YysfCo99zQiChZGrEDh5N1xs1+QA+hqmrKFisP1VcImWwhSy3w/RGDv6HOWe
/V4qZiC+iFuTvRG4JIYPKsy4kvOUAST+en54w3hATWJUCQuQj/a6ifc8szjLjp+bojyFYXHAxAgZ
phjwkB//tawi5If7q/Dj1L58GgD8NPZRIDE2zjpCWKOs5kYO0neldkXGmAwu1Pody03fzwjnxRTo
stU0RnA1XsgP5v+NQimJN/BOZyRhkmefK84pEfAJBFmR8sIh51WJ0N43sgAnI8Kai9nSy/7JNdf9
QS8BDWZk3MRf3dkU2yIWu1GiMNFyIR666dCxgq+vjUrwn6TU2LgI5q3Ny02k0I1VT+FQAUzOubAa
9GqeDQwo9t4bW93h6TE5XbBfzmagC8RzV1E5jO6vNWL2v2RQgZSQYRLy10eddBhnR4qARWSQDAwo
GBgwXg8nxDVZKNSlcpSypmzs5XLf+dR9HhB1iGCulvfam4dIG2XCw1e/4u3KQH4EFKrTTofl8VEX
v3h06Ani6H/amNfJwZddAu82Duap2WV1TLN9ab6olRS4fuhfFQwbJMoMDWNGYafLMYN2p+4W6Vay
G1yk3nUD1YG8N6r6yygXn61+3r1+LECAb95BS7msYE9Dx0Y2pwnrS6xFQVMKhHUzHyA900xaB8t1
UIO4SizByZf7GzeafZGNqDSVN3lpmPsz42TxoA0G5CJ9TP/IuhWtrLrPUJD9KEN0996SmPSvbEBg
tiEdVS/sIXE1Vw7azNTXEitupyn9ANgzdR9nDPSssBZ/r5PWTpuTX6O7k+DIhUknTv3fUO/k8yCw
6xpauixUJMAAFDj8HU1xu64eU36YNVkDG4r2kGNCCW0NxlEcLaUcNCBUpPwCBTkdQoshjtaHYdu9
KgwGA/3xprDgePATCbi+yvNxuLhnTzVFGlxl7krTdBnUvOGvYk5Fv6xSVQ7bP01PLUQVFXDVCVQk
K3v/e3xzdIyGCBMmePVlv/mwkKXUrDISTFkjibrL1FbaDwI0ermnqR7JuJZxtJbJ5KDUw1jRdHFw
Ff2Rt8yuYik/RS9X9Qev94g53px3mm2eeBwuJTa7Lb0b9Ige70o3vFwSepVT5bvxoNcOiyRvHc7a
wcSBUnvvYPboqgB1io/Q94s3EDIWoehy61QbEIWwusJAkxGv3ZUHC/Y0vPpIrHxFI8XdtSHMoDJm
FyGq7c8zCyTqQwlfjV1juLdXMBClcgJtAypskuekFZx7slDUFwW4xrlxBSVt58Ls887x3an7jRhj
k9LslgQn2l6yqCW2vb/hvE93GEYNL/OYAqvdS4KZLIjzzNFMBJNBFIs9epcKZtqyfavkyUomuKPg
Jz0khSq0jAkFLM+jn0AmbHNcwvn1F0RKf2KZoNM40+KeLRACyQDnW+LVwAeHqpvW/AfhB0eUkfJ5
Btk92LP4+z+2FDqJ47q+pE6S4V4CFge9tE1yOEYt+fmGpS6hYmcfNzJeaZdkhsq5rij5nx4LFlJY
LN1FlcNLQp1BR3gsB0sHFbBnRBIDP5405O89nRrwcUGO/1Nxwv1EGJSEFfDJaCAwdZvDMR8ckrP7
O1ssuX3WmTr0QrUk3bLXqanCfvHV5MeHYezG+c1VBOZyD++EypqY9dVkiieAPDFxy/yJ/FHHBLni
VnwKXwAWw4aj5bxYtlBrf7GWzpa2b5COQWaDkutoRxJ8+HrMS6uOEM1GQ4TkM0gYdEXZwT0DFWYX
B/SjBADmO82Me657sRrdUFBTQv0MqqFUVvaSFDsBAtmSBv0JsJlGWY9tV1ZkMfSDn+1HUS6/qLBy
7cDZEf/Me+1MU+3ebI4FNnxNPqPqDt/xWCIMIICZP0VNg7QthoV/zgMBe6cp7jLhMaAkcfuOf7PT
JU52Y2HGzKH3DSsTjs9FjzEhZI/ixlHZTFZ0gkP363UqJhFnFu6qEQYqvA6DTqMjdPD+1844YgSf
pV8zV1szlxR7sIQqjxWMRWGiMtdNTWhAXyDpAmXZL5e8E1gaRz2nXfgKnaFIqU+sW0gS37A5Uqfz
b1ib+hOrLtvg2m6803WvTERIo0wuUTXQExVfE33PeMYM3Athmv7ySsntcImZqJ18ObBIN53AGDFn
NZiIeYnlEvm59/gkFP8A+57S2aqEW127HibRQ3NST2FMXc9+FujKLF6KLjagh7b6KbD+naKOX49i
QxJ8a8c/mnUirvoIwTUalETysXm9Zc5KOhjtICDS+nDiwm7gwGz94x8ApLft83CfqDZk4yxhGN+R
oMV2SJ0hyQy3VDkUsKGhP7CQQsq3NDKMKt3N1+B4Sd2zbjDzFoFnqDYg5u8wBKCqvJRKiY9Vaxu1
DNHldeZsBlBPRKDcc9Q8evEzce57MXhmRQvIj+CPtv3LcxKcmzBnaAAprKcz5gHZ9zesxHWy9P3q
LZmbRqb+nHaVUr3DzUHTRk5NO+XlxetnjTGw6c5yn2ZGdJZVnGoJHufl/5XuunvReyAVPSrxGyBs
6MakgJX/6s7CIFrdF5SKilgbm876aTKVEwKAH2eSZO5VYtBTR+I5BA5ih+yO98tI7KZtX/kogORQ
mDMmwYuJJKI/MRD0j+Q5DgkXrkMlqMO7KwNX/TM9ai2zTbP+UA3HzIRMxw3ZWdZychAApL6SGo7L
SeIOVY+OQfl5nyht0Jgxbnc6CZplFxfxeYxro4Kmr19+4QuJkMhe1cwRUxthhmVhX+V+yELPj+cc
F2Ceg8QbqbGbcmd/LGm0OBGF51eKoOUKhOnb1jystFrb+EpwM3iH1ZJNhq+ePSBl60CcVGXAQz6K
bHVWMLCzH8H5FcHMjvtT6mPu6uO44G6sPOqMO3HRwSrzBWgl7Ee4/F4ooEwct9dkFtCO9PDqvTDo
8PM/iMQcko44+MFgwXQlDoJP2/WwEuYWcndYp1o+D3shexvmwnGo2zSt4TU7gCaCww7nNRiGOwNd
5Xi3EIXMdwazFJpcdWGalATof0jQ7KbX/TF8s0QDmD1q8qXtq0M8k9sR7PFhFxvOBkAbWKEQvzmi
7H+021q6KE5O/pdSSQpQTwHeh5/WmF49YhYeHOWkXuuw6fiqq4gnLWTMcw/cuhc56qZ/JGsLF9Nd
I0BuYejejXhKqC/H1Tvk/IWRV49pW3ijHbGHQWJxT9end8GIPi2H4EogyVyRHuARY2cMkUFS1k/7
zjq3ado48yyAdh1z7PKbM9jrrY9tUT/n4ZeVV4kGqVxZ+ZfffD5brfdMcHBbgtbMybU+e8cqTIFg
agp0/G03jKS7yDBmR+8gHy04edoKY4+3sxyHaSP8rn61KcpPWR1li+UrtVX9umeo9pcVpBs2R/Na
1fmpoRxVFU3xP1I2iwjvRvxKYnFAs+5pllUAGTIcGi0M88P/GCyShlf5fKxzXZhzdRZ54InIk9GT
8jFRd7LdVuFq2ObRLhEdkqytGkMLdebdlmSz8VKabh90aBEAEemvKb1IMfJ8T9agTK9sfeHsLvb2
6qICfYADubC50ngooVAhbz7cbsZ4WwosWD9CjwSLFuXqe98RKghENcdM21w4pW6Vb3J9UKV4Dmxr
rTtCIXwpO4UmbuWJ94dr4+2zr8KEzw7NrU30TE7AgWq4D7O3nDfbiMn2Q28L9VosAZm/X2L29ct+
/ecDgJR+jndxuRzANYLTL+Oym8YGHhh7petmCrGYvUtRQP6IDPVopKXY+XuDEU7v0156v79pruaT
MfPWgxfK6a1rEqEB6useC0+jW6/dbHpDzANCvF9Cbe4/kTn+kp6trVLhDNfWcfOasIXN2ZtmnMFZ
847KqUxsF2BfHCwLKn4CLX5Q8Zu5WAbLJFygj7c6npxaj552EdlG3ExiQBAE1rIVBEEevmrArDTF
zCuNbHRT8M5/GSVqJA6GXnjDnhmTzOxxnlGFdlOVmqhaJQWnHoDQ/PJsfkfOJCYr4AQjFtltKIo3
lksxDBOUrbkS1E+UcJKFw7mEcXJ/dKMtoa0vyNFcrEigMzay39mpPU+NNnDvqp7QjACpFKxF8Qu6
wKH4Jtbpt8pf4cdi2b6H+B15STTz8aYnjP/PY8JyF5R2Wh4igEi5UeuzO7hug2Mk3pszmmnrX3Qh
+b1xq97wbCOowV12HjSnti6ZotHOhKxpZS1g0MOj2ToB0+EH9YMBMQ5vOL8wn5Z0vj0dDpVuEry1
91S/y+C2lbhxkT1irKnncOVrEJrTmCZ8YKrHQQ9/I+VSQ7Cnf5j1d1oZQNhs6IEX0moaz8hTl4ug
E4cTdXuRrhw3+H4ro/3VBtYrAEyISV6oQgOPBJs7kgDGdFrJq1jpzh1icEkGIfszBgl29P8T46lo
0l/16/unlRLc2hSFnXeTilstqwxYGKCfvJEerawQV4GDyzA9mPZVEf8NJfTYS6gffMXTYuRsKBSr
50ZXkdbGuYehfA4h0kIg4v2Z9nr74OrZiedr/umaYIneeGhFvyO+En2Db7UuvQO4kDYHOgQmfrgS
i1g/JvtFaoGjk5ZmjgRKmKc/3cLxZWhdQNcchzxyxVGzDVMZGpLgzDh3SZVGvvQVE9HGiiMlXUmN
ljHzGXCsJ4zQcNz+5YcLuKbSVhXcsRJ28ZpwCTrzANJBbHleIAkJxlf7Ej+4EEX2R1NuaWezQiSH
Bk5zkMc3BwDu1EITEmXu5wpTALnTaGbA+d3hPx/rz29biXWoKdNbeOwYBofgyHUisRop9CFQPR52
MowrHw9hC+ecd5ew8hTieXrY0FrQvpaDkTfDqKNkmieXVb3+gsaP9zlATAEWWTvrjacLo1j5J4XY
DY5VPiOjksFiaM5cKnuvZrl2T6V4fonr1hCoxv9wtoCbozGYzYcoxebo2gqqy+ndEE+kZDBm+x0U
7bSjv6rK/qY1HTbDrV4OUFnSpvTRUI1M02B8C6aCoiF3qt07adawWNmMS6biD1MS3a/s9Btuf8eB
+/0rdrlY5IU9KYRD38PEMlJNq1+/v7CKQ2AZMItTkClf57IoN5nrfYQcNFkvGea3sdt8zekH0IeD
NG5mQIHvPQJW09rEdi9+fT/LbdkFd+XT/HsrWFFXgQyVlbY1BSTWzyq8j1Xji9X0ScdwLF5dkNXj
yVWSvWq5RnRwlrqJ0isZkjX5glEwef3BRrw7SijYtnJySpUN5TWrGUi9nPwNWrX33DhlcH2rtt9O
g6Y4d5Hn8Njc8q+5UwGhgjQnlsMzNKIaZTi9ig7ZOkGIZtrqAGie2JC6YV8a6BcVT39OhxLRSg+1
QwqjbFM9fA4XcD877TfOjp01CrXJkxrcwFH5j3NonNc4pE1ZaRBSI0RJIZ5gkebH3/oDKEBxlx3n
1463VW2+rdvTPnVOowSCorg2yM7wDHS8n8sbXvjswb57GLn9qQWzsBYSdJ+yezLfBbKLNWMJ4FgZ
mlOjWiWL5ic8mCW1mfEra8KPN/v3scVAVDovzqgObFKN8k00zHrAp/BpAmKFl2ekhe4XAELDWhKW
+BnW43WMOHNcs/gy9NTj1kMu/+hKC/Q6gzNhuANsPRn48YKpWu5/RWrQSOEeOQFrOx8ui0C8Nvgn
hi+mcIHMVEeYFo3AbsaiBGEiTGclyhw0oEZIWMi6mO2v0IKSCwB8AO+WMl+RsSatE3aIRP9MUBxi
338vcJezDXB7IqXk4MrDbkR5Zl5vTJriWOMXvZrM9gzanduUUEHsteTSZ1ZNra5Ofm+1asJ9V6M8
lf0TA9v8yyb6KWjFpfWsP5bed0Q1QIk9n/nATQIQV2+u2mH54qmUhz9UHSSNvXVDv+T4oxdAPq0T
lpIYtliyVsXcNAWC5Z4L4dt7jBzVUm4Ok2WO8nzUAdOfO0SjQCclGrGOdRa4NB5O6QOQKfyQlgpj
/1f10RzS+xTKB4EPVmhWMXBnQZTgEMBl5f/fIuLk4N5rYw3ShLYoj9Tp0P4RFr08ACtiL6eIZUu+
YEXBz1nLa30MrY+9QiDtKTDUy/87IxTutIHQZw8tX5IGIp5XDoqIeuWdweZcLVWa+akTcDfA08qB
EzSEiujrCt5dDcr/BKWRgB+pZ7opldu7ePhgHJnV2ZFyRqZWjz+kLHQXwD8f6NK3xxJ7oRgm5m5H
3fmSMhHqsLr6Bch8syS0kEKZl1dJQa3DgUg8tiPzDXl53z1Qra+fah65+8mL3J376mPQyrBoJZVM
BtesVKRHy8/D+z2j4Rem9dcNq2oTxkV1i9QpUu0M4c1U0PZk12qNpxJR/1/lkMHgjEAgFW//AkaZ
9K18V7LswgoYRJxCeNKkxtfubjRWWlmU/u00I0BoUZtFi2+auZMHYSdvvja0HC6cIZpRQXnyPF7I
I4M8eRvqq0ld4JM9B39CujTy8z1VlD2S/hM7O/ogzXHytax3iEo4Ja0L/Cd6goHyu8rYCrUjWd6j
XfUWO7Q7wW3ehkA4g/YYrNELizfsuue2rFsdG/o+dk8TZdCHsQe2zORABgE4zCOvH2OVNUpF+YZR
rW/XftaR7IlLbvfEb2AhYHDD0jPqNGgdyUkIPiowTWXSOI/bGEOUe4vE8CwzpW5LkDQ9NIn9lhrp
rf7knhG2aevAWxHsb8GyxjiXcn2euWj0/18/i7krf3c/nlR5xW6GUi+mxvUbbabNHP3z4Yq5TiS7
ehue7SgEiuxrJawqwB+CUZy9OPkSsIo8rFbQ4oLQ2UtCCM3PMG+h8ujyQfrvGqQTtwpiOIwcSCNG
lRdTJDbcYcU7XMpX7Tta0sD1LBOfesMC5xIavBdSJQqdOB8jOm7fDy+ObyD5QNxl6x6nWCh62Ixg
Jrb+LdgOs/JeYf2hl+xSlxsIbFPaP9vso1plda1Q0FGmxzaCixcGNle0pW/hCIC2B7xr1dcEQ/z4
Si/7CvFxVUUsjiW5/6Tcbyxe3OzivCsDWgjmTRd1fELwkTCRtISDtxjqIPzanR+XJE1ipANkuZ0Y
jA2+Y9hB9jDZk9iMV61IxE0Xt7ys36IVispn8jRcVoq/ZuIHPhdWq3G065YB9Io/Z4QFavgSkOXK
gVn7+q4/RyHJwR9j02JAf+8OTyIgpp0pmtBudRBIdsi4PZqUE26kVHufYVpvM32hjYCF19O0cRfb
K5N1hydjLIYa4BbNhZ6UilR1FKfuQxCD3cagXtN3iBcQsbrfJiZ0HzNMX1GpaWZmvJApIs7efR0P
SL/SfT5hSpV4kky1j3voTOd3RNeA3RmXf0ThikbWGhuCa72a6B8xWRLA3dzLe9iWHrRgtbK5q3Mz
dbFX3qVb1j4OzgeflPLL0eE8L7SkrIclDtUfNAZbN2uCdYHE+5W5K3EwzRojH+kp7OpM/NMnP9/x
Af3fQWc3JIh9UN1/2sutF4JelKyUlcGU+e3/D8vQvwl6XCMTZZHx0EshX5ShiLWs9Z1luBg/K16E
sxHBPXfOuzKYrG9SFtlqSDYCK775XPWyD3C/e2YLD3gtIJW/jmIzSACmJQXkzge6qj678EN6RNcz
Pvq//yg7Vn+p4/CpV3sIKvVWu8cFkZd0jp5ORZnYw94AvzHn47+MoVvEU8xcBt7OsnAmXmT22qZw
K0mIhl7PlnXoCB5sogZ9Nvzm57htSFfP6HNeTGeCaF3iaKUHIJybPzk1dgeF6qKHd6xXXfcB3NWu
dDFwVk88pS7DgH3JqXZsxNu1pQjYRL5MbBIe5uPyk00f29s65ETNO7AlGRmwaFu72a7g+NDkW1jC
fDD+HABFvMFbXu/alLbI5DhVoXt8wwd+/blLc5/MnYDzpQHu0K5FcglG3hsGGqaPDuotN57H+wpQ
ltz5Wknc9jGGlToaFutgH/AWZZG/cFmm+u0+8ZMQivYGma2dWER0iXEgu9f99d8jaL11fipQg8lR
1PjUDBFxyC6zDP01JqRL5Ct2gw5fY0Djp0rKm7bH9z8nzI0Zl/5NYElG58WE4Gg5utTUpfe/IXr6
M6R5QttaOAg0vrFsCbv+VcJWpnCI2n10AByT+EQZy24Gu//mXPBtet/Dyb8wT7iqLY/NleIA4pji
uZ16OOgdm+ZlbmLx9/ukI3qe3Px7XVxWEJ4+Bp8w8I7aNkAYSVWEAq8HXRgIYlPv6t8fE0LMbzmI
vNCYFzG6H+HKJvGkeTL0hlAhX8kV8ziZlgCjcWD6f28DwTOIZ5hGJYY+nDJCNZ89L6gqFR/X0k3H
zUXJUbN5onCP2+JdNy3x1obsYo5Iv2zi1K5Rg6soYrtIFoinyoil1LgNtEH3kOIrltAAHNp7kSOA
PKT/JlG20/BXWxAlMV1mxIEFAsozjTUxvrVpG/9bFxmJ0pD1zc+k78L+p1/gkFHGI/5IYo7PObSq
8ib0uRuRPz7vLTNagzJfS8jRI3PHdLiCaYg7V2A6sowUf2FB6TPE8+pbjM+llPylpKXr3Oekboeq
Kurf3PJX1RGRuJ0LhikXurNF1D+aHnBn7Xo8HIs2RFGTXjNws58qQkc1NqhkH9v7RwYaPo+ZrmMr
HDmFO/Keu43HhjtNSSHEiiNlDwajhLZiwVWJcp8fHHXUYtC9+nUHfgbRxbqtOJ5lZBNFICZDPPQs
juXG1vCVv6l4+BxRYs55+2vd5RIfPSGUQ4W2XvB6sz+owwm69ZTJFqTptfbarTK/3yfk3EGSWNgv
CYahxKfkRN7yhoCWqtOK9xCTwT04jJhs/ad58S3jyotK0EzJ1IpiuybWHHI6PQ4gKY3sFiAl6SLM
eXehdoB5Y5fpUsMo498lakc4GrNPSB+tkHmAf/GQ1y0+PDayNmluRlYKzmpfBsNsox2qoC+CXm/d
D60xYDqPiBKBblZRLW4gkb3g4ZzFpH7OwesOsBp6bpOl/Wipf3wLsh/+d8qHIOjdrOs4EnTwKHLP
FW2dkc8JONIwoFYN3sklfohXnc5VHN4JH4MyeL+96dV8492Bz3CSAbpnj/sOpLA3/ef/8QAv4Ysl
jysMUKeYgpf0LOXXXw6II+/2jEJdb3UsOHzI1VBB3R6dAwwQHSBUf9nMnZIjrA7ErKYsSjA58RSE
komk8moacykEMMu44R/QBpDNwQ6yrQxkwGuxvnnPIoKUJvAl+XESOX+fGhJ1tpXtZkUVZEILzxbc
y9q7vRtgU1aobIhMTIPjjpciMWGUkHZmAWZZ0qWIsS2qFXTCrGKwUroK6cQ05OISTiN/7NiGEa0M
jbocqKnaL7e10zW8UPwrJHdZsNPutDYCxmQqjHaPTapH96/XojHh6a0K83hvoxJ5m/Ma94gwHlhM
53ejD09Ipukcfrd0UdQf7Y+rr3FDMAa5R/TVHSibcTESL592ABOJ9xHuvn9wHcPo3mKUduLE/jHh
oxqoDk+bkxCcQQiMbVjdfQ7s4Hv8m348d6Z9iFfUQ7YijgWCQ0Pb+34DqA8QfeH6mNHITN4oI4pF
xMvFPte1oQObzxUXFo86GhJJR2lbf1rca0pc4fOhoROmN7cVI46xOdq4+yTL2swlgiYR9pY/cBfY
vSiCqvUIfb2P8krURsIcqXr6e3/MJJfFcVhbk5IedHw8xqjGbY8O7g2EEEAdB5dllaJ34aA2Y0dG
C7mMhZ9WzzUzYZRjBiB2utmnzTx+DrGmmKfsd6KROPYuhzCzxT3HG6lpcR3BEyYY4iHgupCT0q+k
xmqpVUNwESjRVUy85xeY++eAQT+AuZ+uGJHUmMco+/eSCP2ZvAsmbPnSRukDTpIpJh/1e+k+bAvT
yrsYXuJArMd6xliRpc1y6CdJD/HyaFL7gmn2hrdWoCI77prISDzfz9Eg2mZkvBzvoe1zzxs8jj2E
p8CeSP29QJPdX2rb7GDET/Lrrp43n1er3iFStL/N9RR96mh51CPvw0t3f+0TncJVXK39XlERPdoZ
AdJ07ST9CF7UQZbu2bj4hg4P1jugoQPt82DewRWByi/tB4uJHA0L2iHUVXqVOUq+AhcWuIOx0R5C
Qbw/LspnEa0VORn7uPPKH4agCKG7ZleOv3FjNSiwdaknmBPmJJQgpJkvezvdTArWR/skfISU63vc
cWnfnRclG/hXleOvuQUIHB5lC+3hQTm9JA6eE8MkQUEjTlwjC4EkiWt6nk8JO744mJPgAqu5GSsw
PW1IBwETxo0Tw6PysWm858hjeiOa3ohmAFEJAmYG+9wjTY2fkrQerkYIQuO/a3NcG1MGjkqM/raw
6gOJTHfWIbY7F0/tRl/At29mtLiyQhcr6+v/lQnPEYjujc96PUqMa2r45prTShp4fJZkm6yOQ9q2
E/UiE1p2Nc9JShV+gPoWVhOW6S/PPD624Gcr1P0NyNisLuVvl+X4oHGePMdlEoVsnHc1702quKjR
fXlhgGex8zX2EJKTJdttRGzD3LOMDss+OwMuz7EBYVUb8wzrH9LQXzOD8JEby59oadwrAv/Tbxx/
uni5UCLqF0c++nwl0w9J5P6vArIJkfspQOkFamYQiuVOWq2T2aWRfBEHCIbmWokwyrZ2wOO+FDRP
VvV0OVaxvG+4tm0OGUHyIFqEgzmCmMqD5WUtreYr53HAlewXoLxsz/6a/xA2RklcxnhYP85MYB7D
93iDFm/Fdv0lobicVc82ZCofdgx7d+pi+B6iYLo+ZHfSjE4cKXfRBBA2P7BH1U1d3f2zDmW6GSCD
/5a75ZNZAoMQiyPpM+R4KHEno4CB0O3KxIyNHR3fgQdkYGhvBKazGXYF9TqWDgVcOAfN+tkAnXmw
1w3B9fc87c2NFIqrcOkbHIRp2ih6PXNAwATBzOoFcK2Q0Z2Uyy/DoOTTzE5oEDZVtUreLl8Fu8ac
jDNt2rKYkLZ79kULOM9BODIdHIDHfMDz9HiF1RxCJp7K75/EQK9rA725vozHO9PJ41MrfiVnvU6P
k9/nd0zxe3jeKqDz+cYyFhaf6OyWGw6YejapaBq/4UkRyBmJpjKEaagmCzIpPEZEzlyyAKSN4CD9
8Jr1ZyRl6jDK5gSTbbdF+kAvLRKJRIOFIeuplbm2CsleiRpF2kKWODgkYe0SlsRCCH805YTucGfy
/VX4DefdEdO0vsUTpKKGlNmUElnDhHDzfpNzrTdbOaGc3GRMgNCwPNOR2lq4z5oQSbpKpPMRswfw
qHDDxsOYLx3qvQWs0yjuWYStEnlEv58yiQ/FNryg69SWgFdx1CEwrTFWSJo54+1plGtiwVK+2c7G
04uygpe73qkqn5x78iQHespdq2gSi9b+Q6wP5bJUQwT7LmFGc/82h0TwVxpnK4lELsWHWT1Xg//P
8Tz/sAMfWnhwAxDz+ULOe3cl8EdAsIj3GYdPGcO5X1eZiel70aeJVH/KMcmRgdpa/V9nN2xaEHaw
PJDaRRYADUaW2CYm4l32Ki5kVNxe/msmrJl0sXS+XjiV669B1l5bsSJJkQTFX1FHzLK9eLIIWhkw
AvzS7o1gQQOdey6lii3cSXO17gHzaYGtV4mPJXBrVy0XbDxuc/DlMP1YEW8lD/9sDFWLzbe97RM6
a6n8XhVVrdXStDa/g3EH7Wfn2zX9wlci0Eq/4R6QCy7QRBNNUPjKJUhFLn33pRQsTw9Fd061q8si
xSaqvc2XogtRAY4704Uz5j1mhsMYvdKpZETM4kRqrtSV1CcvJsIuBvLmsxTV1e3g/C0ypwUXE/Mx
vsgkKO83//1IeQLYUxHfQNuKMZq7iYXoGlcso4oGxZBNQZGk9SnIzqHJ/BfnPEdQQAlo6q2cP4fQ
sbESHIkKXmQ+Vy7KrSmzZGXbIGmCNtudvgESsxie610B56WE70GLdR59Pg6mo4BW88lc2gb+t3yC
u4mG7CncfL7QK/6M+R7eZcKPJu+0owRaj9YgygO+3jr7QDe5it4IweXYzsE9PkQznTXBryXJoKeY
xPZwd1LohQI6lu5ax+b1s1PjeF+0Mkv+uOP7rT+VpmjjBPEn8ahuQkdYhATafJ2wyJi6t0ro6F7V
OT6rmkAUvwHdfSeHGejz9lW8RzkDI7fz8cyJKiFZMdO+S1GYHC/ktOpLDe/p1weicpuVhUQJn94d
R9cP0tCbBF4Q9uFAUchnyZaazhksOGeDtH1BTq4dTyoTMpYoCnoUs1PXLtaGmUKgJay0y5DFoGst
ZdHVbtx6cWpBdA9XaPSOoNSsWV55gJW0MpE8KBpCetT4gonUcZLVkmfuJeq4SqQWQ3vdbMm2gjgn
TPqz7IDatPX6EzzXXFftgq62QYJWZWRUk7akuhmEWCfUhGIDSRzx8+qVgnlZFcV+zqPgMdwmVg8L
KHv8sD2aT1nmb4ELXdB413qSpnRlIgsAnsPlPjrEZjrcosEZR8K4qLDWFgZPvUWr2eveb8SWw+t/
5DSIfz5Pn3GcfG23+pt6ooS+/INJyvbAkVvXWMOE/m/u9Q3FyknIHIJLUBw9v7VC9pRaDBpLgKPg
OSdhA9QuALOz3kRYUSMdVLDw/CxX7KC+8aEnay9BzBA5IaBrpq0CjnFb/pwMDupQ4hZC5yY6a/KV
1S/mGHPOac1CJMfZ2UZtZ8xGxAaQCaChbb9ygSIV2luINAwZS4KWqHgj1Zx10NIJ0tfSFhVEBrVS
3/wEQwbMaxu0IUXXDI+hR9hTIOTRxEA16dgkmP6vQyHKzaThXUa4kvCVzeZX3QFNl0mYRCZUkcE8
keoIuloOAOnMBDyM78eDqmbmieQYMbm3HAU2hyaRAVnW11+OUyEtjYoXLVXr2eG8DhWCu2uwZuma
hRuXd6pwjZdzkzeTIcZMdwTI6RIkKuGJH7dJr9yoYZrFAW5bh6pmo0mCqu5ApBV+7r8OInGlEqqp
UBpUfVZzTPtofCdufT25xtYn4xR7gzeeZ1jBVWh14ThrpQ+/cXz0dfo9TsTLJgWFRePpbskclfzA
lPtaRqePmmFJuPvryE5hCKzz343Os7xwaNciW0sc1DilhudvWdm9byqwMHkD22lpN8AkeeAzYnDe
zsqYi9V4o/OEYg==
`protect end_protected
