`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4160)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosb+EqZ1v3SQM5cugroTK0Ogv/nKwWu
IP3dGkUeW4FH+9YU+CCo0CN+uO6kZ4slP0LVtqG+59ekLqaba1VneiaBEjGRt1Gz97p/C1ncB81D
lvqjp/OeO71QSqf2Zhay4ZYl2tiy+Ew1f0ZkW47vQINNdKO/M0B4+2Kd2b2OwA5iNh4jb38Q8o3K
fFSQL5clNodY1kdOeu5Xj6KBtyhTrCkKd8EBaxyft3gKcQzAMEwlBsXsIqRMR7e7wmoo90CZ1T2V
h/FjVRslDCwsPLBcuR82KHAoQDhJYZoiZ85DE+wRg7oUU1MOGuX7o9lCVR9a3KTbYEW0MJAwz/IT
HiIqZrXLhn/zk4E2PFU2jeo28hX/mfHLvV3yPngxpwTjFFcb5j7ewghdvNnXVaA2CQGL+Mwbcfkc
PRLG4i/97b5lzMFbwJBFhM+U9z/fc15JjYngRZlx1i/xRFdiE0b1YvF8A2m7TFOO53hA7NH7d8Y8
84KmhPDpZt3nlTF86OzE+MjKa4ELyMGzsMJoijx6GgEDcYx2s6eIYxz576nb1al7IgMQGfAhJ83h
HX4zNrP7AOObnR/OZtx3yfT/0uJM+FDc5O272E6pXlrVoF/5L/KtZv3fqgxiYHtck+qMyXFE15eD
tQ6PEU6TSAUSOAy/0ktFByyCyKzA6rPf+IZpCgEpCTdp0qrrTWUghIaFgZMpHZJQeIGZV+klnO/r
9Li5iQWPsrVPnGs4I1R0rxS/WJz73vHpPkq7IhXA/Z8Lh1qjpoQRDVRhe2F6mJTOC7wF0yPpFPZy
Jt976g79m3BthOiBVRKFd/jmw7emcIZWWUufkeHGBrXLyXY/8XNhGa6fb9xhr8aaAT6qSwqsQ2Za
Zva38aBGRJfYt014TtTGhhN63kHvF+g5S9PbTlVH1J7dNUW2PZk4imYUCw43HxrgjCfSu9rkR/TL
YyLCg+oy/0HYLgWWr/Ek0Eabx5Lrn3YkO2QiLHiLBN+H/A33+bPIEwjJxutZXk+IY55A4vBLV/b3
FMtPoat1bcLkkz6A9G/1frD8krUyEQmCarJrL4bbHtOk07QyvWovIOArvyWlXt6f/bTGJb09DkiR
BfLQXfLcbnN5sZhyv6RcGFDqY8D6RkZEvZa57nZE0aTAI7spDwNsqUflPRoRePWZvQl4SeaCzL3H
ZacAvJ2+Of2nBTnGh0zbMeBNOdqJAsjVKYKB3qWIo9POk2BU18h1Q2s1K1jkiNBUe+CqfdokJVCj
WeLewZwAfO+kSehp6a3XjopisBkLDVfz5/6J4KI+3AX6z1gmXW0xTtL5IJhNkqQGFAPoIrQE9qs3
HCj7uqtzlkRcUELEumdmUEuVUcZN/wh4Z99eOanqZjv8y15ORVg4jP2+c2W7jELeyd5fBQXAeG/v
zsJ0+ke+eK2IIrJDL8bW5sfqj8hi0lXiOMJnz7+LXa1GozsF9yclxbVhBYgcsAz8OSKZ2737f9uf
462gEFM/v2c09SHIMjwi2oJ5jrMWBgpncsNW/YOaCWKv6VJM42RKEu0AZr7ukdjhRcrqYNMn43KR
7zL+80GMCxShJAId98bXGok3KkW2E9QxMwo1+fQl+6r2m4XMrr/B2p3aMjjSQM7F1VWZIc0R1Gqa
tSIln6lfHhVUaP01E8PhhaxY9vxfWY8LCGGxDdYKLTAJ9hbB6qG+glUgy7/oOJGKzxMbOL+Ejgh9
sLFXp7ZOZdNHRmrWpBgNphP221E81MPLXTZPlxa8AlpfRa9Mq45Xzp/HZcsSBkoXB7suphjPhoE0
p6dy084PYzVA4xNxjQqQCvabYd7JyWjOPGhCV7b1uMpq3f44QUnEU1jF+IObKxJ3t3juT/5+BXq9
Tm/K/bPSax3leY6PWv6IPCphbUIHmmp8jdrPctVHcHj4xsixNh8aIqaI7XB8cXKZBqleA2eh7csI
8Wm+JRu//4b3dSzHkaAOhU7wAb0tnqykGDwy7plpYR7AArh4VCQ481GRYWBcMp+ftP6glz2As2jZ
IjfS3BuHX2Rxk9LmG1D9+omypCOhzPiawZXaKCMu+OvesXqK/o/tMWCWeHc+HSoB3DNsqYTxkcXz
iWNGCytSdgsfXZWJL4r882C3hkQKem5QM3fgANznHKOJATTRL1xXJI3sQB7zGimZFZp6HR70a+I=
`protect end_protected
