`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62128)
`protect data_block
wrovcHZ5qwQL2M/nAAAAADoh3SP1zS4qUaggEsoaVmcLHFGzIcxpK4nQenRiP0GMvlBnq99bgbCC
sN8rrCZhixpmpHpJH8E0i3oa986B+D1QHg/brz06le3d7ff3/oIcxg68jUdO+aFyWeVbTNWDmLUZ
sIMH3VdGyTN+z9qrDhAoC9AXR9M9aWbgpi9C/XKAaW/ov4jlE0lOouxHOne8hHB6Db71Ax7NtSYy
RunB5cDBtUENvgvLsqx611T1QAwm+RvJCWO28ij308S5uKOfWNC4l6JSUKf2N9dLAh0BfRxKrfUq
sxvJSFfpCuN8rn50lq3R92CTxhU6qIal9u+vG/GLk00jMPBnXOBXiJeaR2K7Ph4RVz0kdwKeQ1Pe
QPhoXygEFPD2mHC/1Ao2f4sBIVLO2CPhBKkOPQQIcU1uWeEZn40f/AxY0Lyf61Lccwuq2QOlxZkt
0Y3jRfoaTW2McaQVuaV2J7vSnYvyQjfnicu2cynKDfBg9bXZk6XoRJugYAcq03ZsKtZlZ2KsnGhK
aw2tuMmecF/Bdyr2gJ01NzAmIjCXmkzrtaSH6TX9l2tJmkC4PmJDj/vJZjdOOOr7vLm4aGt3ATwY
PBjw54l21CW7tOBgy1vwQhMScZHQ20Y+hPvHiHAfF8tBArta7g2whGuXApKy0aPlFnOrquxcDnqd
PZkU66gxIq5qi+3lw0w7afQ+U8RTYBdYkf4JpTJMVz7beg47Ox7C1zhHxwDTe2iJTjF7rmmNG6qB
YDoR1+MASxmuEbIySz1/4pFJw8RzQOdFGqXjm+63+xpr7zSHhJ3uLOrwWzb1tPubF/e3NEeinvW9
qN0p+7YoYbOr241jZ5zV9x+aXhnUkfro42J7EqYdkMo8fsbvhazuAtJi+yt0rDdwLbaR2oghsXGX
hbOWue1I8g4Tk46m6UcB7CDL979oKsFKO0Eed4UUcpwxj36LKqWoMuyyy6PKpYqkIQZ8HTh8Vj4W
GgwTqVzu/nDjrjkC0px3wDj3cjRGlU0KSvxmQ1MtndiVVkodWx4aLxkl/gdKW+aGjac4W9HI+6H0
Gc/dJUixMDwLKeoorx++ZFgdXHCOEeNdq0D0N2yXEs+DyhjdplpGIi4YZgs6/r9sDY+nsbNJnbzE
2P372/eYXWRG8/ljVGhMbKlp0aToB6Iw/ljuf+4kjxQ8bZk1gpO6Z74jd/rbVasHux3JJC6C4B3m
lofDmSkYHBvlr+9M+07tMrrUJyeIrR3JowY+/nY9aVhFGNbjSUxWORIgDGKSQlVuYlEREQUqJnnB
fn09gJTLi+HHeHwqb/USE42G9AVA0MeusuG6fzSWsCe7GAHmIj0dW8MGVxLR1Zb9w2EyRu3mnSZT
pz074apu7Xb0JPP38W2MJrBWSxZSR2IqdqjnmdP5zclsPJ2U539kSD+YJ5tTbnhe9C3js6pxtQ1B
PQGDycN9ui6cL4ixDwdWQHPuawU1Y9nONirSpvng+H8qZTqIosm4I/9fBc0mZRr+DvBE8sAk+rbI
pplwbT/t5iGp0SIYCj6CZhvCTA67T/gLHbFutR9ycz2a2lWOJhTX78x50w8+qudeYLgAEKloBZVd
JJbT2LjOCJOV14JgQe8ba1xxOA+4KTSXyGWUrJVKmeTUIPTGkLrqbDHvARq/Tp34F9gc7I07Iu0i
4p+kzpWzJxnkW3i6uHjsX/He/RLfroddqdg35ASG1+uTVf2/sushfMofbfjnw/8OQEvj5vj5kJgq
PDo7XoAVLarz4SFjiN9vzCuq9rlxCgKv2h3sYjNkbGXu7XAph5jska0JJ0OOtD+pA+08pDe2sq7C
PCCEjnWLDZK2Tg/cn+Hbw+OhclZRUi4GDrKNO5c5vcohHXHlZ5omRkhsYSNhykcXp5AI9p4VDbcq
GGoEBf3cK4aYrlxybRnzLZ+pEgtt+Y3Kvs1YqjO/NADDdWsiF4RpZ73TNUnHlvf8Ndd50oR2bVQJ
C/qNTP4YTDGtvZLETScxtyqbHa4R99SS1gjY7bWMB7s/3iGRpvq5ScHFCN5u957lZKph5XVhd6Nr
H1PSzL4rwPKu7A0hxLqWui3gr7wTJktAHsGBLU4IHyFXRQorAcw/Yz7Fwyd9H7uBFYLIV6J1thq1
e8nLlm2ADEtBlRtgF9K/hG5nlD34pOi5ZUbX/ZTJo/kTuoIr9ZYP6akMzQUXxfVLfijfddC93Dsd
u6SYzG4b+NDPgq8X+R1leCEaTpawGW49XKBJcUdYI2AelHF3S9ugNvD/ZorotqHCy+SQ+uCcIaE0
cAPOQJxI+BR75Pt+x+mZsEKTxADAVVJyyqdRY02nqf+lEnCfWv7wLGCODcsTycT5U3kROpeq06Io
RC4cgcZZN0/Y3OtGz6VGKOe+brG4v1rHnZwaYuwyffhdzsn+BRtIREOlM+QLlx2G175IlWW/6s1T
xuItTBEhhjLlPImEJv2KNXkqebQwq78KAuYyXajZSaFXJ2PgoQOBLJANhCDR7kUUivmZHfxZB48p
fqfZ2apZfvsV3vjvxzTP2j0S71N2kPy0fEaBGly98VLL2vVK4oaoojKv0X8RAHU5f0lHzoN++pgz
BKKZocGUzgJYr9qVEeyDzcF3kbpUjZH9JWX7Y3lG1Y3VFHHcX62FCd8jgFthMzABIdWQyG7RIf2n
tl7oCSqVg0Y7V5XxSmHyeOh++zRPts8RkkYyhJiESwQxr5zf7FFPtYIEzpyExLoUOaG/mg7rU5hj
dZSld+k/n2nd+E8O2McBV23wUa2e/Faa654t0ixVU4I0gW+YM1KGtaOzRMK+qpeisFxBaB0U4pWd
edzjfmfvkZZDspUTTuNzxEt3mC2xbyuYnk459XFEnayC1zGQIsRVH840qGhppVoXZmWIaibH4aqU
Qzp0P9zkZ9UB/wgu6aE3w9VnTbU8j1+y5y/k/S1moSpXajAyoEawrPX6VsTQmUPYce69GWYCoir5
UG3LxUOQhq/Nm3G+MaZqhaJkt7q9nCocKf/SvhO/lTBAWw4Tv70hYo/P9j98SeZveH6db8c6vMOp
hiMbQ+FabPlV7uFfn6eITOEN8u86LryHIVVG0uqGrXe7D+66wJHuAroshtbAgQpEfr1z2eF91qQb
MLpuNzx16csLWU3cUj+y5T9I92TMJ0Lb59H7fZ2XKzJWPSK96GOSxli+mRlnC1WX2RKwLRJ56Fli
niFAiUM/ooiowQNuYEnjxmP8GbKcYvUMNz1SVAwXRUpvbS3+FJhJV/xfavEDzBvZRtvezadEHyBo
STj9Dzld4gy4BRPPsy91iXBNC74bz8J2H1QWtONYXvjmyH/gB4Ftn9dD1u+egDMkexipZq21mdK3
HDkvdpJLELRyHiw4rtY/wpIOsK6cOlAeSqHmgXCKTOtdp9H4xwWnknRH3eVLnsyg5Q1hYKq/2TvF
9nNNLSmI9yiuBKMPYFNzK0hlAKsFDVrTLx/PaosHLpwv4BNZ/1LORzSSlKUSiWHuUaBPcAduz7rp
ue35MusHN+rGAubNU3clmVD4S5Js4feeOHADX7lszwL9T0jAh8dVuzcOuriAqOyLmyGfTTQFDbF8
w9K7E/8RvOxX8HseZDmfVmxiQw+S6APVOVniimUvckFIAUTsLVYmhZDvmC40AXmVxTBFg2hWFoUU
rWymoPM3zu2lrR7OeHXEacbJHiVmsyG41yeiglBTqZ2EhVOsoxUSMjuZP2K0EqlzzHUIwBHNRnPv
RG9JeO+j+m9v/LUt0QNDRapH2bzBuMc8bO5Yipnz6t7lT4um3wbWflVTwuHvZa8HyZMHpiAGhHJX
ax6F3Go3DY2waaoDhAWtQ+jUOgOteh4CN6+pl0WkSK0zmvWUbhFp9zLlXQ+tlmHcoTfrtRvcwb2f
QDEuApYHT2bfSUVvbwcmRHFG5LNpkWcryqFHSL0nCK53ngSkxHQzylkXDeBNKyjDXs+a4kgSHJsU
jlcNNxPniMWqA3PwEdKO6b9fK6n3nMsYLb1ipML8i6XDBYQc3NLFzDQHygthqjOheCgAy7/dOXwA
HqRgiSFQUv6t9mWr6UYrGyL8fKtAmFmzDbuwnfYB2EyNxgoxlK8pny3gHERpYwLLov5c8b9osrqv
oK1x5Xoaf2wfVkBW2UwUL98qvIL0Yhg3Vk1K15yAgxtPBErw+mxvNAD3xfOQJSoQ3YtbCo3dFq6q
gK0DL9QjjYS0sJDpvJYGRHbHr0QyAfMx5AKLAb5IIuyzyrOJ0169jlQmC9Dvxbi9w6buTy1bEJhh
Q6md+TL96q4pj5UPbYHNTX0BdbnK3bcEOStEcFkvlEcEFeOlfqEd1WVss1iYE3hindCyut9RJlFP
VjmHEpT9xql1GtYRvO7C6rDSV1MB4F/OElKgGneqLicDloYPnqRIpX4AIKM2vvwFa2CTqQo57Fmz
jao0pNAIZJEkPgPd025i9NFi/VryIvbVmQRCTVO6a+Ah8152R1BCuZbBL1Ul55gcnCwLRODPe3qu
Dus83FvmRyhPqtuxgxX3cqTVLBSmysi/ZMexdFwtWiwytBnl0o27IG0LCDteH92+ylDwj1bY4jYC
4S7BL6d/BcuZwyb8/ZiUHpB/wK5520b5az0NZ2iLhWFsrDl4AjB0p8MqmcwYXz5FDPMiGFvFzXXN
W2vctjyyksiGWoBDk8jlj4xq/5DF2VDHUBH3Rtx+G8Ar/SZQZLFhaNQX7BFTiWduxfn//BoRPCFJ
26UGPd0m2JWkKwUL7IuhHiyzfPXxsFvoLKZ5jSXHxfWSajhbsQlhyASMK5+CozbMROsMNTDJhgZG
ts6NU5IAxEYVOsOUHEtVZtOkONXNDvMpDJTFNu6rVvoGTvd+OJh7r597ELRx/yaAfS1IB3smA44V
9sasdPNmQwxfTfbwcV9VbBLFsaRMsSyMOCwLeU3sSbUJB/0tSY2M1ttlyZhf9Cr1CvVkCQ3qif1b
14zeFhuOWiS8+TYMQ/d6GE4/vfrvPZmh/4SyNXPnOI+YuHzTOShdyAQNyi+r54QHozvMEebC1Sv4
IlTTsK0hUK2MhbXM2in/PRUJ3l97faoC5vytxp3j9sKU7kpgHkBOg/5Fw3ZEiKfdV/XUnI77Czsv
gP9Wiu/6GwJyjcbk58C2nknqWlMgLBRrydLPUZwQqvmMnzO1ZlkAdk+gjrC/E6rswhk/MC8ggSp+
aGPREbmfX0ipTXkkArui6lO4Vg0DoVyKG/1R//3TxtiIbM7MSr+LJxvvIsgsjnrg5lIV3kqu5hB4
6Mna7Bo9LbX+Lh2IAdxylXvEvmNXBizxe9iJAOc5RcHeJaFvp76Gtv8Zdwir440HiAN42FtPyHHE
5cxaaVLSCW5VrMNuZHbJa5ewQyzv12Xc2btFJ/YJUCWOUs8umKwFMzkzjma6UcBqGug4EShh15TG
B+jzeQjZp0F5NLmQzETRUV5SygPiLjSwYNrvn+AQXINJVS4OabVovo+51S7KdL4b76sLWi5/O0ur
KW/Hd4h+FWSL92owT9JsSXFNBBNmluD67oHCF5z2nvZEvTLKuonOuvwgiNik+j7bquBNmjAS+MRQ
hylLYqsgnNZ5aSl+05DH/GkVIENjieHQRbAr1s/BuGkWwGtH6y6YcbPltxIqB/FvK7dHOg4igxmY
V19rgSH5XxPozSi1NtS79lc+vaEHDQWRtOA21Yu2X4xp2XsiAgag06W8v2RifAy5aKPJX1fwmkg+
myu+Wdr1JL0spSRlxDL6iBKFzxkevVNMcKT8SpOR9b+57SJAFBQDfYzXzev8YaYFx82ql3Oo0PKv
gYZuvkC7kV+tAyzBD2Su5ff6r9JZfJUR77+qU9Xl9SijtYnFEd/DPz4UEE7XCkm0C+ShcvEhYp0p
Tjh1nBLuAgTZ222+ngwsBiamYDZaiHZXYND1gzB+iP1nqXtZblAAUP+03/HPSrmYul+utRI5SFcX
pPqQA5v9kRKCG0CApM4oz6L8iCEy2P/9O1EGHSZR95jZ6V9nsQgRLK563DXF1dJ4lse0zkbi/1dD
CwSk/7ZrpZJPqR9dnrjSbhqyNTLpbrY79kKT19iO/VkophNlfQ68Khw724qNE/BWOJuuKajy4KG7
o0k7GXzF9FOvYA4buAMZNl3LDQqvEim1y94FOKeHgNTJ+6m9Bxm1Y8hoVGji2Zu0CVSjevift0Ms
bLANzOqxzGKTE9+i2P6FXhfTmSGBWFQvT/MRuu7oqQywx38xOw2JjVKe15UAbc7p1gw5KO/hjRHe
xhHHa7OBILARPN1vARJvPsnfdZfB1cx6r/UIDPUWchLyPmqKLXeq9v3ZoOej6Jqx2ndyYHPLrIlx
liZjh8srSo3uzHqPMirAn0QguUF854hbUPdliH6D8PFVS2OAKNgkp7bEPEijTj98uhaouv4xRyay
inhBo30aeiw+AZYGRl5/Z7Ie2fu6/1agzXnh2dv+VMhFpUsoEBTPvU4SyjHzeSxiINjnHXtGKLiz
pKZoVXFf8KMiSp91UTOoJttOVGr7jlFZa/JfVpMzVCHjdQyD8TegS7kZrCbHgy/rWCKPoWSJidmM
0SHcAsGoVjDV2eDb1CNqEfjViDGuuByb3zLEh3yPTTvTEbksIe/mF2P5RsHEP5iqzKmX2nWSdRrx
fYxPrh4yeWsE/oJzv0vFvDPGlzqmIhFN0FwBWnkFZD4MRYT/mB7Hv5M9c7yTKvZx9PLmUuPRnbLW
OshB50KbKXK06OHCqnvPpYXd4HMYuvJpPK8W+mLrjZgOpMkUVmfoh6JGhuPd7gSjtN7lT924UaSI
Xu+dbVk2MC3xlnzG9AnIQV4yuVqltp1y98/m9JpBt0EfPZhKlfLIuGHECwx9ye6X8LctaEL8yZ/b
d+fwui8dsu14gscobZ73ciJ1ALmZMWOu5W4yGT9aTG+xeyeCsbgn14rfkx8YhlW/jdfygixH+tCK
l0Zcz8L6/c9ZLdpgWL53aPsgudfEAdZka8uDR4dQPxxfVmLYhS5IOuR4MkGCYxfKgy5HIP0TPiPc
GPepQa3/3mz/uPiyNmRWRaYqBteFYhidz+eOgH9ATPYrhlG6QeEbxEsuXZjRNsSDStho3wy+CJPL
74xLEOt5qIP7hGxZ5w3Wa4O6N98UbGFUaYUWN8u6g1/QlssSIu9FLl4R37RO/5/BQDXHgpKvHohp
OuF24rMuFPzCGxYw5D1R4iSiCqXj1uJj9DC0LbI2zb6bPZndm9p/0fujttcaDCxAzlBZsCN+SsKY
xyd6Beurw5rOjaDV7EXQ+SGUxkvYcojDmm2GlmtSF4UhugVTvfSqJmAqtZFz3xMztqnZ8jIwNjMH
x+EstAAGfqT0wGCN3fjoi620YYlwiJ3G3+yXWFsiuJoDsnQDhkE4XBQNnpLQtOLLT0IOKpAizY9P
xa6wkkrih914WfR5j0kGo62zy34Wr+K6aMp+29qvCvv+VQothv4K1K/c2qW8fxX5Hg7TFZp4NDZa
UIke41cmqxedtikT9b8CBP7Ayedi+i2GaXQc5mzYBhO5pm99DQnKTiLNO0FZPxrvVX7VBnRsEZ/n
E7CaB46wa90QygF8qSH+w6nJ/KZFhuRgXozj0YEcbmWqc6cYnALepaTVfaWhjBMvDO9zM6QVOqVo
gcVzm8I0owpN4c9A3N/iaBSaO83FPohl2pSX+6bWPS0H/DQcFv36fJgdx/mXM0nfXx8qD7kUokit
Fvj7CIeYFDuhppnc1rp8MqNikzfLcfCmNabo8Pf+WL1YYURYRwMf2b3GXjE+JordGOQ8YAv9nrgy
2YSsafu7utCBEEPlmK6aD8DPGfdt+dxC0jgmkzKxPj4YA7AtV1QqR+PCN1dPRUylN3302Nth4yBX
0i67wWeH3GXpTRSEfWKpuI0zY9zP5c1mFaH/G+7liUw9yQDb8j9vV5b5gPUiXq6lzpS8JARhDRGz
M1fZWlHBwDmJFqmAk8wDOfdhTo6OZdcpKMbUYB6AQ3ZLA0hY/zJg695a6PlRGuVvtwMRd2YbICQl
UHnafvhoVM/kC0fx7SyeIl+dHCtezBqRiAkN6LOkKkayy2Gqy7+kY7IgamL/NKS//OIyfXzfgU4f
e8C1p+hwTQlltD/gtByny/mODUesJH4bJMve1uedPPs8zwyKEty4K6aYLdedABJNHHlnKSj+bsNL
/JfzNc1Gnce0a1ghshNKz0hwyJEGnEX4Xn6JtjEuSVLqL0l77YcA9eh7edHpQky76cwEZJNGwv0M
xkIMCmHC2mA/QPaSjYx05WuSOWfRVpr5SdUyLn8WGFGnhaub2loQn7nEkX1R1RSkqGO68gOMBOzs
d/69EFvUki5bA+ShJMl/wWxpYPbXJshH8Sxa/NLKdztlanpn43fpEyzWoHmI5ue122ltpHuwYa9W
/dqJGB5CVeAcCXxOUuWoPoAN5FHMWTdyA3HMTUNpWqzcZGELf6nB2YXAkXLQuom3vX3F8v16CPZG
H8K0xF+Wh0dr9hNaStAnxlVqM01Isx/9rVucCTCKpd+iC9L3lsWscNX43QhoYT/t4ILX1+Kf2vIK
MaedXEYWemMw9tOtT6ni0a2iUrb7Sv/120SPuT0KS/HlzemSk491a3gD8b55ua+szX2Lujz5dvgM
rhdi9+ijeBFZ12ox1KEQWFv2QU1/AvSpA14mNVKrv4thvGJxKKfjYoazM3apXMOooVeeaxeLPB8Q
X1yEubE4TfufM51vXsiKClDR8mOr1P5NM5ndLNkNJEDo1ppTYzkxQCRohAGuhEJmsNY1IC0677K0
pJVH+B6lFQmIVisOdA1dvM/5JvjYvZ1GSbxsCDsVikWMjBbb+B0cXwSXkpAe0q8WzXPUbvbxOAuJ
ADBV5+3/s/HSDcjeKWf93PJwfB66tqI8lGGH1pyAhrTNTirhWmq93mSFywM3+FNglKoGMyo43L5u
YEZxdap6XTcn1VsRlbzWDEnPh+f96aBwNwdG6/LBMQnoE83rIxqTX6N6syXeNDbdofk2xZn5UZia
+6i/CgCfF3WNAc32jNbKFEHnliriGio3SX1Jq6/AvGEXqSXvzaKJ1Wx5BmR3weC+tUMFlMGeo+xK
R4TjsYzPe6R1dMTPl3cM9tQJHn0IZHS0xOxTZrDEYN1kfRy4cROHntAXq/+UXYTTrHtq0B6NjBH5
E+i1AqdnnUQA9IsGfHLcF4Q/CvHT/rGMHle1v5OOBBlV9y87DJFUkaZr8HFyUEaO1XkKyZ46+bJj
aWge4wG4D8oJtUwjJ9sgxYkuXeLKa+v1I1F6RgKKJbaBSpOtKLODsWqIxkJOC8GgDKLnz1yiRnnU
SPnUMxAl8duI88paV0uFEQd4veeVKdsyMu1vgn9IXjxA+e7wxin3wo0v5TvJkLLlkzNKaCmw/LNW
PVynpeBTYf3dIyvr6aKMEyslUuNsqAAoQF5yGHJ0Zs4sxk1IYODOt/xQmsgwZgxSIgFbMFBndwkX
lYDN4SnKZ1kXtl8yICdNObLHHj+xXrTz84GjSUTxOUPKukb6f7SbRXSxETD2EpW3HwmFOaI4qad8
xZgR8PvZ51RNXTA+QQmawbrDwdSstBrpSLOIn6kMyhdxWbnsfNx1xqUfxGqWhLAbaIB7j7wwpIeh
q9uc2/WVS1ylBYnxHdahgXdmT/bjrpg4pOT8i1yQqJl1Zp67ZHbeDnZPw/0e6YAQmSyS0oBY0kmZ
fdwGBtLbLoVRyRl+Dfi78bOqxxh5fFJJN2jLuvYchmL5+CT9Qinf48fxrHsUFLKVHeokrTYsDycI
loZGyndV92YSbkmxV59JrIe4dempd+W7vBIsPt5RO2kztd8oYdvKOkS1bsPC/m4sDcgnbsPtLi++
yJeqG1Gphy84B5t+2u63qtzxt8NgtoH25GKQ14TpjZbLK3+ZopHxYN+JefY7+tlnUVljVnMG4293
iPDTnt6Di7Go8LIcd7XNuZOtDJ6XccSW7qk6WxglXUX89ldUE0j/Lg8WQKxjbrhpicJZwm2l4gcf
xAlkRfe6L5pCSRk9sIvP+r4d47B8gBzbgtFDlaOF4KnxHjZX7bXyUO4oujRLYNEvbud42UDvkHoE
IyJ+YL58fKQOuePtcWE2EnSk94L4+dHwPZCPOYvNxPokxscdO1t3RX6AyNXlyquktQL2WGzLGnh7
FLbw1/CZAzNtZbK4hyDa/axL6w9pwLsiV1Lu84P3oRCKTiXg5zCCgg9wF27EZbfvtlcW07cS0hkR
dwTozxDjULE3irPeQh/LW+9hsPl7RG32x5lxgk8J008DHohmebyQkGGINeFxAjCmJzls8AX9ImL7
N5KWf29an6tC3AoX+ihlZjZXBNpvXXft9r0gWiq+eFAfoiaXUIbdjfkclYVG0lRbToI//utAUjFh
hbMO5ElnGt18zJfpoLdISEJW3enoJes1gPWGDMwfC19hW8YL6HEqp9vbNTIPPVOjVadou1Qe7kjt
fNzAd9FNK3ct9e4RN8VOKEPm1yi/QcXa5yplDQ1UIQLIAA8/iFh5kiSpqbydCdRiFqn66yVI6Oto
vamaZBoZtpN4ve6873AOFAjaEoDsKiGH7Pw1tANPsYAOflfhcZEF1moct1nrlgK7oQjyrCM3qlr/
REqp7IpPV+BzeD7NCci3ao1XfnMtEeCPiPJmNNPG2gNd6V5w+aCzY2WqJItOIKqDTLlLQHM9EjSW
ANC1hwEYMvFwZczEbdSxVBK9PxLIWZGDXrXhi2PO40tZNpFvZqN2W/v+a/veyJg0I/RZnn6lmeMs
KbN9e8ZDiOInsBfRWkdU4i2dXsmpzzY+Bqn8C2UAw32aeoE/nCku3Eys/JxJEx8QsLz73R+4a1YM
GXCCZcmcH2+kmd9jC2HX7XVZEnk7htU2id75vFfhbriHHgjKnvmMy82XKYATKeg0Qn2p2R+nXkyv
jCzuxoCgXV4aGhiVmq54hss7k/IQc2F0CA9MQGm7mXX2SriUND7uP5pPl+U6dcuLS++qMb+jNXY3
AUk+gm5wzqNdm17Z2S0tmEollzNKVKBbztGVMZMViONs39bKtahPTcelvmhtkxsnAW5+w6x7T+fR
aNVaesnOoozutXfBWZqZz9s0mXBqtFVYJfIeKk5/WPpPpnJV/cjyQMJHeItlapNb+Ld5l5vX0+h9
ZljjUYyETx8eZ6TDKtfrHTLMNCvtO+eSND1sY7LbAaXSEG6n1YkZMoen5LNkLYnXPY7i8V20Zp2f
k43T44IKr048ZnXenVLe/wpgW/sx8//ePw0Rt8ZUo8GZ4Kg6j/OAGbyiKo2Z4v23FCKxJuFYNJEg
G6cCTAam+OTjXjjz828RkeKwjGXoz1VqGrl5RCDOKDByyP8CJOErxKXpKm6lPsmUlbpIJPU8LcZD
mBXnubTvqp7CLCgUF8E71Cf6u7Qw8CeN7TFVIx01Dg6cbeKQlYAaZqKh9RrmlG4BpwYmaJj+TdAu
uewFaAMxNxgSGuin/TH7HawDH+PHNm5uy8YmtzoJSYQ2H9mwMUg+XoD5Kx2IwKmhMKuSiHQvbQlv
MLUIoin8A9JWsn0OhnQ0gtUP/y2AelsFhs6Cl8/dMNn/Sy0nvq/XjeGDiKosFQXxXoYRqyJ1cMzx
yClvFvRKZWzDYbncpDBswiuC5LI35/j3T+QAjRGwyDGMvK1CUykh8yS9I80eP+zqIEfv4imzwfR8
4E4tx6d1F3yLE5bF5glDW+emHXnDjyLvFEuIUgAvjahi7Drj+IxOMFOkCpchA4LbNCIqjYsUk711
kLVxqRYvaXUfeC0LUIcjI3kWPcWFHUceL7mySNiJwy4B1sPN4NhC8NOWHez/OGszqqHi9TWUpTiE
pwuBa5sLEPFgDQFrq6XIU1x323UPcxjAEzcgc/YD8UW/jE13ZONOeymt0w73Q6Tk98noThRD/Y9T
WBIn0LbD8LWmqTAmxfMSh9X31AMLC36rntQm4wY3wpNq8eBKVDOwIp1jDY5brbO3PRsxxPaoBMxo
LUTuAx86YxWHSZr+ks/vvRbJb4Mbdx6EI3TrvU14X0hUDU9+M3zN33DUiOP+rqUpn39n1YrLo84A
xTSBlvZ3ixKLwY2Qu58c1p4zPNM4vC9dxpsxcAlRUNIYI4CsTZM2f3MUYyoFA0uc04wGgIByquLN
uj7zGVC9igHDVh3RgWF7yux/BeHf570AstM+W6CMdaBe2mLtDpY4Pwy9aqd6aAOunRSlRybbx47r
13CD8HVquiDsX1VUPHXkWNLjHgz7OTeEWyHltieboLwptgeVmdj7SMov05CERYzAgyu40Latb/8l
1Yhsa9RquAidSH7ZGkswu3WUXvO4wXoH2mwpiaCT9t/H01elDc3GkUbWKLaRFjdTPMgrkgQyUTm4
5f16gUFM27DEG4+Rvc75GyCMrO07tizWspz7anh5g8hRFAdoAx/RMm45pw2K42IfWnEdH5DkSSfH
5B7UpmPnVZC3tEEBlZcatSPHSTj/GTVltaNh7wD6xIKOke06CA+siiX5wgf7HZK8jUkpNfiO6PEK
NntgtaUHgmhtUgIp34nrw0y0a5TzxTnSD8KDBd2gqYP0t3FaoxTKeCBnJVniqmgOfmJw4nhiprXh
pPLYx+Ji/f3uNTn/R1X53mYR28vwJJxVLfA70b72uvRh2jgGf7O5L7EKB/RMG71VyjUcgu16Al5i
ngKL95FRl8WTfhwe/O1hmcaV8H+4UCNdmO9fX18a/vPkYUvRcfgzi6UWDBjtz/RdoNmQJCzepBUf
Om1reHVPiU1lEn8GZavFpbZ+Fj3jotZuuPj+VNHbzrOaOvcpn8EtB99iDUciRphVhmpl0HoqhEPz
6vADxSb3nNTPeolkIrx+K0sKWd0ffudayTqS9eyTALK09nec9eVvxxAHdv9TGRsfoNXU2FtydnoE
1B+xLiBjr86UjgM8CgKu9HCvqwlhfkDJQysxbZBaqu8hUakSWvS+EvvevJ6E1wc99GDjIu2FfnVZ
5eLXu6vVmbLi+a5MgoDpKKZDERSOCWwkyzNuQp3QtTj17KOBiit2X8xtn6DDMViCooxjJgyeckWW
g3LIWLg6iBj+bL3S0dItU5Fspm7EdoCA38bGAxkSvwugCFCXJIoX+7PQ4GDeaCktljLnY1TjQKXe
z9y4bXpQVbeTy1jvSLNkyZMcu4audh7ZnjguyYSFvX9jJF8C3QeLierlDtJO6M+9zaY49L7nTnnT
2USZl1zAIIGkMsn1lChFIW9BDhNVj/N2HiXZKsWQcE04+v/iacI5B1aRxE19+UCNNyACNFFYZ8t9
N2QLyi0ALTQ0BeT3/Uo+vi0YVZshX5qeEppb5eS5YfaLnykcSXG/ooAm9dg+9ZRyIJK9mduo44Nz
XWEvkEh/e3O8L0Bm5r2tUIcaKnMHS9PHeJO9ZZJeEEYOpIJFCG857r4raT1IhzSyqfRcBK1kLPjz
tNiWAXiEmtq6i5ub46altKUYAZ0b4g+bNTOsdgyC93wDemK50kRKgHJugWgksGybYcybK6cxZ8zA
RRAh+D4+i3OejeG7izgsbS2fR8DpousSWT6LpGpcoTU1L1eHo7E3WPQ3Ti0IzmZJPAGuB/9eYqZb
aAzg7yyXbwjisoGxgQ4IHgzFX00iOITRgKf1in61aN12r7JxFllW0Td/BHJOBrSjz26FaOqjdlVe
8U6xa88ICpJlNHrMcy75TsoMdjXnQDDClDj6/qVnBKraa8WsVDP3h08ip6XeuZu8iZ7fhPz/8hsJ
W9TGII0GSmuIK5rEwh75kx5tkK5TaWVyph+HMqp2ctFp0XU/I4957sgKSwfATuSrMGmcqhbuwKK9
UMeGbOHPYfUs3ChU0y8lTOUJldiBKitkHwFd2j598vzzeJGTyz55TW7LVsMRk8npyscpXvM3cXVl
BkbWWoLbf6+diNEIdrkXbZcm0UmmyVcd+DF15gIwoBERp04V6l1rZLakvdFf8Z5QOHj71V440Zn/
y4MwvQX6QYYsfMX3BzZGhCNLtuX6Zb3qgynnxg4+amnRHWsfeWgwvDtEqdxPXWNJQ704amAzrwRZ
W2fGDX0Li+jSiUUHH+rH9pJ25Sapi6rS3kYqnpzJNiqKS1iHcjLmESzZ+vK0H5NdakZIqXiv3iDN
UC0BNT04Gz2XaT+W7SgPe5PAkFtDYDf/J58HAcIXRKQ8CA5L2BjiQCYvJAJLd0tS4K/nWHfgOjnc
d80xzMhu/EUietQ8ggctDImSHGryUOqEldfQM5XJoxwhtIGFlAJ87nQjACO26J7ArLbPnwowIg1Z
lN5k45d13NAXkTJdRPGwLUUenl+XQzjNKPugayTxrJ3KynubbeBb+xuf1oqrqzPYbnAKhzbBZOQ1
KPb6kq4Jx1YTzKGf0Zj3j7lJL2GmEVCC5ezOD2W3iXcRGBhrNe03soT8f91rpZcYURbDnxxHNk6g
cYDGCBVyoyhvxqygvpbA+65b7a8ypvPsy4UVjmyyqZKv/1N89L6rZnNYk3ECINqEBjRD6AWcyXWa
dUN8URK29NW27RzTZCWrnbBEV+Av6SHoUPxGS5UnbEe9u/7mjy/fmr/cvgCV9jHC1upd0u/0B1fQ
rhCQyECIunBsttT91qMaJZWNLgtOgG3BrtrDufbimTU+G5HXXk9PsVf4GaSE7l98i/Cx761B2wOD
Gkf+5bM62P4IMp4pPHi3y7ti1S/lPx8phAxE6/tvDSSbuQFQWYOQ83uytlUveM3GOQf6cTqwInvK
96hmXWn1ssc9Y3/B5bvtXgPP/jgRMQjxMcDg9O4IyluFpe4+Ouhgx0ZXsaViZbRBtvnYTwxOjI+M
zOdtI3MA9oLtyjaeIjAbnE/qJgiKkNAjtrjrf0uJeqgZB+Cm43tWuIO39JXR/RBYS3zWxStybJ89
yWK6jRjUCB/wL4Nj0RVVpdLf0SKgwcnVCkJqL6DJXWFfkbO2kEh+UZAOQPz8DIWto/iUOpJYq+wq
Djtg9fmPSUgtQo1g9N6OvuVSEgoqJUC9l44rkRXmf6uajOgZe/GDDrNpORePZMZ8+4uPxXsFVeQy
e4/y+yX17w0J3yYYPBzWAm83nitM0MJqazVOx1O/2Pg27e1/2qcol2w/zDrZgmgzSSoeK9KDF64R
KQ+B9ZnyJQrAOSDQ3QJCqZGg9Pk1KAoqSya4tKzMiOdoK6/hrOCwC+HxIwvBno/J6S2jZLllLnaH
0Rpaa/gqMwNI81dYhAeOw3Qrmeuyb9m7Yyh/exmgSlmt41saKU27LKDI80dh9oWDWIDgGDaMu9HW
GMqHuXXknDXpL0K6JIMLwLNoKAKuq/1mpbAW1ByxTPu5dqXTuugMAH7at7gmrhTRr3f0XwHtOqvf
tnIs4u2So3NVhYY9QdfjAEFGQa9Pletqd9N/RStbPvjWglAyhoDA/g+X4/WfyZq/Mz/OKWS0x8lI
RnrnENV30PHJK1FVlC3GeMlkizrjJTjAHszskCbejF2QGsqPRetCeZ47n3XSqjkd5mXMic33nb98
FK24Ghr8sVwUP5HvWwgyMB5B5CqhP72Qh+ZIgR7ul3TUSQbNzgzWZlBB67seDoU9L2smXQCaqofD
z2bke0E6m8c3qftLP/VeEdZMMChCLfxzBSMBjmV9U6Sru6+F69n2Xr671GfZMIm1Slc/S0XO83Kv
syRYooR/bHQ2E8EOnHTW36akubec+Oc/u0HxGrCFbC4NyQJKoiZN4zyfHL6Lt/9jLwIoxQjFtdtz
jbH6a+vBX8NVC+B0rdNF8yt7BzBIvRt3zbXaKnfNUNTrdNnkMoOR6uPZ0zglhRz8WH3LMCq7x6Uk
CvEqwvPKs+E6zGN4TUfNWhxvCozm7f2NKXyiltIBoIocmtzsxF+O0JK01A9Fr/sZ39dSlYHgJkZY
KImcKpm3IPamR8kHP2mnPxBb+Lk/H1mGZW8L25hoSWCpGJVUvUkSPVyptsllDo2xRE9YrQ5IRvlo
l4Giq2XQUNbTSmq4vp8F7BECaw+pBENxF2az2jxOOu3ZRlJfvtgD2Gzh6WJG/PAKe/A9DG55Q0Qv
pmD8FmVqQagyIguHaqiWoVzvS9T2gSvcLS4wB7WjrV0FNRDrd65VcYRjb4cge6SivKu86GmVLoed
jzy0WOqAoHjt7iw4/Rph8Ijqj9j7eKgIPID1TDIrQAo0gruLvMXUlbhgJpCUkavz+gcminmEJPIC
ioGyA6aZqCp4kouYU/sGr+3D0EN0z6VYNuk16eBEAQfF/numDk1FU4vSFgAlrNads1EKxBHe6Bhp
t1RKKeWG1XCdZHLwXFDVds2LD8z3RK/TYCSmewtMb1Lmr9y/O5lHV6Y0I+WIZk5GxuSSbzA7JA+7
CFxXnouDKSQM8k4cy/6vX9xAlcBHXTLEb3YR51cj1CDw38Fn43/pEQvXQyuELOPvvKWyHZE4ySju
0l1YIgPhrFkzdbVEjWGCc0Ci/HcW8MhjTrTNifGZYjVz/lJRfbfBqoGFZYgWj0+smYX36knVvXgp
wHyJHk65tvl6zYOWhPExWqcJsziIkGLBTNb8H5sswZIT+p87P6wmYouS3ve3PDZOBuOFAniLyrs6
oS2tp9Z/PUohC4EGy9fPRHjjAfL5uQ94r4rIqlqa7fJaEwipfaex9P+dh3VtSO0r/1SgOq3cTmjy
0T6D5nZQ/c+7AOlGhfnivFGSNSHJaTSYAA/IWjJOcqYsPrtm5ED3VKld0iTTVDmnTnbYmM/3lCIe
Jo9BPCq/kOVPOLwYWRSQ7YWc0fjRqN3asfNSMkqHri6HwPF8z6qKGDbT81hBgpAokCyeFJEOXkca
rozImhVy+eAkgh/DGU5IFZfNiDaSnKwMWqgKIO9rJUE+tgG3zXBosH7678bDLNnBsX1C4Km8AQ1w
3ThNZV3flgu731rfwr21Jj6mFNa/i+RZNU+zH6NPnBFc1C9TzUM3gDzp6Jg26PZkMTW+W+Opux/8
BUHdRk2sKmWgWIxqLMGIpkcbnl3iMoJphnhAASyEdsAKuEwugqcILHzqJKS1Nu6u1gdwMTI3zXBp
16gqJ6g0nIXchvGzmIDIoWgjgHBOXdu0RC+UI9YX3JfAJEMh1XCAw5HS44sX81nWDUKxuzkVHdzc
Rtuuzl6WGNnP3VcdFLYuqyPJK+mWe+0Y7lkoS5+t9F4U/TQquwwfWomOEACeshELSFAwwv46cQCo
2S4tJGC/HNQVx38UvecQXn2ELC1HNoeJQjZ8mrlYjwA/3eHnSnijkiwf8axhxKPJLcIdeiORd8hd
LUD5j2tBKlrDWJ0fRnvT0wIfFUB1H+bYVkZkqEEoyNPSvysSaEnuTiUBV2G/89AtNUCSgJTiOpn2
+s4c3bpOanWtBmUdNCigmCfKuv4P2B2zNgENvP1/14r//loomfy/FWvzQ0dVeGAQEXExrwDa5BGy
awfUilM/OPmpV5Lx43lzguF6/ukyzxJp/kIKyV3EySlh4vtYIx6w/e1mAUa4Xou6HgddAz1qvt9E
5NwhRot/As1UUsdciMm+v2Ayulsv5wSpAeSqvjMBkuw6SUfpiAknLl7KL2hsGSMKGkF3Qj1Jtsne
EvliedB/jjM9P8h+iKvh2sNZrzk6X/uLas6qOkHFbrAhhPRk9tOEP2YrE0PsjKCJyxc/IY7zWhDj
W7bJhto1G7U9dAZsrov4xaWqPhZuzZt4jTHDGgWDuBD4q9/BrPXNoVRzGgz7fp2xfM+Vv6/41soE
9SaHBll/Xz7VpTidL5NkQp6IBqyQg6tuONbMU7iCqB+rJaIU07q9FhJr25sm4h7PFFI6NI9vVJcS
lngxbuJ/qqdYzmPBy2N7YOdZp2+6uNAta7cR0JqynwJg2E24/mP/XWnFYuk1rFQ4bSkMUVnYU3fr
661Y84rdM9pPMsTY92+uFVURZSOgX0OhyS0NrmfBh4YQEVrsmDfvyb4OEJqTWAO3Yxm0mdrWFQ5f
MgeKf/xRTmoABBzppe6CG3HV65+V2+L5TU1cDWkkk8R+z1oJglqjsN3OmQgSlFwJqsMefrPb7FLo
mzwe3iPSB3UqglT1g24W2GJtY5dsLFft2LWT+y13/pNajss6Vld3yesDcW1jP6UiqyRfVA4Ybmzk
Re1Xoi8k0PCCMcAY0IEm2BsCbWdkwDGpAzNAKVGnaDkKYxmi0q8BpQ59oYON3DcnFTrCrXXfVORN
QLXyipPPRHvrSIi0co/OBPcocNzayh55ObSglOEvMiQNKNW4NBVjNM3vvHpbFsz/c7U9bonFgQTi
f62Pdu2oYmQ/+fEZzoHqm4fAhDKrMUFDOv4VIdxnLhpBND6ErjpjXynZNClQud2INsk2fFEzi0iZ
RfOxhyYRqzxIzIdM+FHzW4Pi5P18skJMcMk/9KxihT0M7nompAHAGzOjZL986wVq3xLU41t0lN6K
o59GL933tPXsesQvgVAk/fQJl4yIZr68wnJcSkfLOLEJu3n6i82QNpg0tDqSwDLOLK0+AIYCrABp
4WBdenLXS+eLyaRwlZKu39W2wbis2oM8rtBDcXt6lW/PVn81WdCXKZ3zboByLyd9oaPnfb/kEgtr
TvmU8aFBPhuFaN7DF+o9bgIbhMBbUEpzI+foiM5r8x2zpbeTwGqjyytIzWZLpWmseq5+an+gPhCg
Iy1J6GFQGRAHRczvB7qVPLtPo7MRb6SCt1xQgOd99rTlvlZrfHibl32/9rIlKWWH1QLPXdqr0Oh8
MgFjNbhm57V1EZufegwYBhNZLJSVYrvw+iGqaNsOIrLYvf+T5ZrHXVDVFdagUQE+U7Le6T7OotUp
MFvVU0djESAtimRGsoWAS9VKYG93AM6Vb3JAs7cKerhwFeEAKlarVe23LHGFoy6/30JgJ9zg6fc4
wAmczDqV7RxjU2vqjxulrqNsf3LlZF1vN0q0G+onR9GgqzgUsj3XgedwScdaheaDjOMO9hl3vJyY
mRRpTMNQ96kmQaLu4aNAAvfrSyQhNHD3PZr1rmnwxwl1EeBMYi5LEfNYO2mOo7TdoBep1OomY+74
E7OpI4zWWWaLtksKw9wXhj+Yfq0VtGNtg98TUgPQSLffaOAlOm1K1B98Pol+b7w/8vibwBKFAXO8
5JA029IdjGXZxkyALuf0bzsCN4jAEs8GjPX7ISD70SLK/5WyP11UPHAcYWLCc7BDqVQ7N5eAr43A
Iq6A3+o5CElXL6hgwIPWyGWgJur7I9sC8iZERITBrBE++pHoqCH3ZTJNOD2pGg5eAKd8ry2pLjUn
SxigLz/k8hQP9F+lV7exaQI7KdMUTAbbne9S0qEWL7cBEx+6fcUKCa0UEMMEPJjEUY+TpjINES/b
yquDWYJrOZptQMGmJ9SM7aaWhg71H5P694DK5th3doI+FdVOmOTTx1H4jef79FqzFXJJW7fu+JDU
2MkC/HUBH6lvSdAvhjgfX5PtZ4pxn9UEOlXfe9znuaJFeEWxFm5oWmrlWNGaJvVkja8BTKQpbBBm
n9fZfZ7G9DN0JGYwJ6Q9nWHedJohoCGoxmEkrLjQJWgmRqz/bYLPxb/a2jK+PTzfj7zfZwiGIvmz
p3kqnS7n1XHjvjJD/vZXcIEUkFYdPmvVSXbYD78tDl/kWv/kKyNc8DU5D54s5/tCTKhFZggGbzg+
mJr8tgb6xW+1ATheKV+EEfZZrtIVxVIh29xWaC3ooGwpLk3LW5Bqiz91RE97k39IcdAaocnBGm/z
8rSEmL3oz/hHCG7mgN4UrR/5yGtOIrQcO7TKmbsSnCKL5+PEdU6MYSMm+8ZZUo6lPx2dnDpCWlGU
W5NLABfNkVN/49qX+jOPbrAiXTNTRtT2xN+QvskTh4yaBg/gJQo22fcBbYodr0lO+hYt5JDLS8tU
1ERYSnZCSaUXna9j+MRx7DJmg6AkflWA+W9GEPCgnWQu43GXoOkG2szhf9cKkQo+rw2axyG1+Z8l
ITZDQaIlV/ovuRZmXqmHwbepfncXIpS0+YpbLS8X7Ookt0Sk8vhRNwEWzpFzLT/FoUWLxmVnV/7i
zI06at/8DH7LvSbqpfc0I1EKInf5BbOuY4pPq+E8kKpY0jvg2MQt94RR8QSxCb6yGrG9Um3SfCIe
vw8dlgZwq/b6C20YMKmXpJNYMi8XeVCl99DHe6JDq2e0vlWTcP5nlr+U4xXMIRmb6MMp54Ws1kVc
qZozRO/oJoEMq6JPDsT/uhVYT2A2v8iZ0icsM2r+prf2Jdroz0Om2s9Nfs9ao6LthEtoaAL5FxGS
5v4980go5YUZukZLiK8VSbctUXohfbnHinTFLyEnfbcetf6ar6DM1VJgFeA3Qwq87/GIi3ZynCH4
A+sWyAbWvffX/iNx2CUS55o2OxocadLKhoILO+rJcQf9AgQUIxKPNVqiSjCRyMiQhvzKgzM94OTv
ElEC51Vs5mcerSkN2msY49bHXUpKodOXEIb72V9/Rzv4waTuEwFhjqU4llZdsUX6VNcI8tsBwX0s
mGAZjLigdnNWdtq1SA1IrRlia/AZM8ARqIL185Ftl9lb/v7cSBWfiPtEAfDfTpID3PhArL/8XyQM
M3UcylyewoUlMF3LxnNAoHc8ONogbiJrIYQgwxRPAC5xIriZ9twVTFurdKw6iYkNWTeqWUMgisS0
hroVsfX7nDVI5V/92GjeNVoVNy6vKdfxNtwvHZs5BVHm0rrZ9UEharQtTW+jqGh6k0uYSnP5Twiv
D3s5dPZAyRv3R+cFbkbAVBHQMnTWViifYAgAvdX9ioCAjQZnG1Vfsu/uHElLlW+TTuI8dMe6gcj5
VwcKvf6ZllrLfrV6Nq+IZvLP7LO9ujSs2wqKAbDLkFQk2E9+KlCOWZxXZB/N1gfKaJD0KepQ3Pbm
xoWSkgTciJLhGSHJ8UubwRGui8CwEHYxqnkIDUr17Ac9lPZHD3SWQ2/iJUwpyc5PCPpkq4a0UWhq
dKYY5BaMGFKS7zs5bKU3AxqRUXV8DhjSw8aRWNwQjiPa47g7mUXtkaWef7t6P/s78bnZMHU0xGMX
5WSbY68HuT5LZ9C1iXcPnxLecWODo1YbF/SChAQKEqjUSO0VXSU3P+f0D3viLIWLmMA+BGz3IEmV
nE9s66oBfQk2xt21FASh6xU+ub7uCuFNFCNyr2u2055rzcUcokHuajd0uZY+S8CHwTpg5pMi7psX
a6h0dQS14RbBtXflfFIdqUqrOEyKrowoMMCW1IIOWLYUQS3E854BT/R3nb5QnSidD0IspT7D4pzE
2b6XW9B6AqwXiPcEdRwYUAsvUC1Dovl9yzxYmTZUa9U/3GCFeYELjWIxGJoGNU3SOzGFak9FHvyr
Lxygv3Lk2LpJqwXdpKysGj8wByq2axcS/hEvPm2FP12c1dle1QmSa7ZQq0eY7GJxHHg11VdvLonU
e967Q0CHBEIUw1hxphV8qC0Xj0gYjDoFluaUcNWJqdbRA+6SjN6brgKsqTyDlk1cjkLdv4Joov6v
rc5S3zIbg4w6AqthuwFWu4xPac98myyIle6aND9iQG4WkphR/+NuSNn4vUL3YvgPluOBhgtapVsb
7DHQKKeLJBa1QxJjoaO9DnGs3yNYxzXGq/oVZ8giwWjOg3LoUAtW+IuAc3wYDbxoxYrPva/5wruR
7Zf17iOFFOivnl4My7jz07q2m9ADHtfRq+A9wqkuIPsSl1pJ0SzicGDUQ8t29u26Ii7kLmXhGAXB
QbA4RHPWFRHjrig/HedV+c4vn1qZ6zfJzBNKf0HiYalKOJH86aM93s/KtHTVI6TU8EWHo1DORWqx
YcfUhjPZ6RGnLa0kDXyys39n5UNOMVIcaj++SNJ7h8cgyRHMjxduSRqcJjr+b23oql9jgXa337+R
Y84VoUSMmgNshFu4Xq8K+d0TDmoa7j9kTzp75K2O+R5lMCei5UD9i39ycs9lPRPQQSqNhgQSc+sE
wgrfE5+aoXnH6eWvpENrgfaUAUeQmDPSwl6z0Y7okgL4iCkJF6MhdvBGjpuU+dNVwvPaGaExWhB4
Er3CF5QHIUd5kS+SVSM7TrR8o+1eoS8n/t+wbpRvIZbhizIOOMgBAsXXIsSziCTn29x4vDmdFiwt
xgQzM5TJCfNqccgISgYEdORlwuA3bGsgQsoWGqgc/a5WXceRa/FJw8diQGTULz3NhwhxaI6skHMf
Y94mRn36yzS7k7Vq7Z8MkeBoabwRBfm15zZexosq3pBqTJTUUWolnPA3gz7cR7ggZFPYORSmS8Zs
FpDf2bK7f+l7xeD/pdMkgbwP6bloDjMg+2mckbU5RjHGrYQeB37vN2XD9Sm19A5E35YMFCO+kHdG
IFOcEpi/84eUdD2y/8DrprH2xUOHX7C1QoGFDG2V9DRlRxgAzMfWrN760Bwko4s5PtxKcRg9RxFG
5qtTPnipZk4UsMi+ff+uNPdvKUOxJVcoGV1s/3v2zOrC3861/LnUsOT8CO6cX+mD8Fdq3wIvA7in
ltgnZ9y/3hDxoP/VqsI4i8O6Wjk2z7PFrkU5/TfwYpCP3FXHNvp5v7kTPtpct+ULkJ5v0Nvz+Pl5
yu/R3VUtBTTU2gZApsA4v1UfLFmLgbTZi8upJTL1Xl8pp84+OEMRS3noz0LcQH4KtN7Th/0YJdFx
LNHhNz0XSO6OdQ+DVQiQKN+bbp+40s2EumWFXJNs2KmpbyWf2TEi0ma5wU5j0deAqJ8GN4pOFRYv
4mhAE/opRmdUbS/0PoSQwGaUjPEbEGiHHdWhP6yfMegAKGN75zcRHn3Rz2/Vxm2BOCrU3hSqSH2y
2hGPNKdaMX4OzGK2Bbnljcih4balNQNW4dwFs/tphiwWOjcs7byWljTG8tUdviYRzyvCh1C8/cOU
1ARTxoQEgpUZ8RbwMlN3uLo5b7GbB+QPm5kPHbVHdwDRTLNiDyXSf2lclBasjTfKqszOarG9uiB1
p7nFOPphgwtf3ERl8GUPTLWh8e39ovVR8Itx2/Yz3XpZZdhAYhZH4PZdHDa3ISoZgiGRVpMeS2ty
LPwSfkTY0ZsgrNDMN+JZLCIDz9JM43ljkOKa+Ezf5GpaFD60wOKy60rC1GFihLaSAk8em4TwYLJA
dzaJjt+20EzCLcLa+fI9WMyBEDw39YF0e5zZBqurqXGQ2XAV4HBHOTHGQAThrnEG9PtdKk4YidMZ
qzfS6vdXAFd8QBRBI2mvnyg9pJILoTy0PuM+5+KPmp5f0wq1980t60Nay/cKgRx+ai6aBRsG1oRW
uYeUqHBSunsDtax1yz3VCmQsf4dxqL23sg1iGdcwaPEXifYmcAvc9sGgXXYxT0wFtj+d5KPeww7T
qnSsWd0l9VM+1UvuRCR/uzisHByEOA5XA5JlxU5xAZF+INfitNYBlNsNkyrhFkXqo8mRSEcZg1+W
DhWkd7/TPdk49QHHWi1OEw+iRwa0MnUF8nJolqzp5iqlDE98n9SowZ7hLwhF23XjfxWD9INWQ/Mw
6wyxuZ4OSEKtY/sd8jScZUgUKVZeIEqV4fypIAe0LhIwKHjCkjJSp4Mix6m3lPjFprKBv8CxZ9xf
DlSHyqtMgpGTEt1xEydlJbHXzmYSU2arV4Z8F9phde929ULrsSuOjTKYm98CqxhD0+Chvtx1sQ0M
i4gmnC54+3kD2dkv4n3RcKCBARTfW4H+ATzKKmV2RXQ5OXYB6yaLBftR7E1y1dsv97X6ovUJaJyb
eBc2vTC62086G3U0PDvcDCixSj4MKAbkVKSedduOY+MAWq+mDz1PxPJdDdUAOWT1MS+dHiNkmBmM
TZkEr80oN4fMaOFYTXBVgFRDqIg6Aa+r87SPSXCpHkPBtZyLI3NhY4HschyeSALqXjIfj7PWlM/u
nMAisNm9KB/YdKtNYcN+qsGYEj0CdRgvFG8UIONLaAwXXSzKxbyNeuJGuNj0my+cKzUKrCPqaCiq
Z580jkUkpKEb8xhx6nn6XCS9rMq6SM5BkuCVgMhNpIBkTfM1IuDXJk1OWXxCkzni9r22d92B2GqA
QI7JjviqNuYFJNIC8MwNthGHH/6YE2Oo7Z3ADz+0vkAtqXW04WhD5iKMQ/1c3GqRidjDlijRt7jq
A1IR8Wn+OBl5DgRYvxU/Py+RFVMJMH2wMzh+IJPkiG9RvWLcxRySn2r2006V9E+eenRzqIesiPzX
E+VSHvJkru/oDx7SVKDhkJCtqh1R2X1ug3ZfNK2qa3EdowwrRhqK7XDEbK3RluF+tbhT/C8ktTrs
kXMl01DYaq9MiNr/uBDGs3V+Ba/UiHxlTlvS0Q+FdLxKcdIW+zZaIW4p44Wc6estC0UUJvREbJkF
XNMnj3zUNIA2Zdo/tQTOHkCwu+MB/03HXtU1t2XicYRldwHyIQyxk91qQVWltklDJjOz9EsXCLtX
IELIT/FCpB0yMBehKeytlypVuO3unrFFyOP6TNZdTvUL1DDcPXmJFWh9kCuJ3+mK5UKuJQFBWtWQ
yUFkRRPWLL9B6fnoAIUb6ibNr05R04zOarHRV6Lfb7fl18hh9SttUHZtehd7qzWgJxDHmM0XNWsr
RjKX4p4nojxsM0exsCHI35YHdK6x62sHh/s97c2kpbpFmz5ryivcVgm8OnKZ8cnXQOXd58IrlBBS
XgGeQ090MB1dS0kBrdVNcINRAG/4Tj7/2p8LcNbmzDGe58pvHVaElaW4qhZ8kW+hVY6FkvYo2IJ6
H+TiF+vMb9r1Q0wnCSs1f1wAmioKoToRv2Ywb6d8zYd52UBtlWfuFC26T++NR9RVQcBk8F8rn6sP
G4A0A6t8TB4bX9hi66vu8WK12plqkQnoLZtu15SF356styQvNgNMPu/JkvZSMKxGXEkBOafm0c3p
hL9aSSrJNqK/VYcesV7tQjTuuOLh4ddoU3Re3gpol3oy46+A10tUX2SEzHJNeoU1jy02UWXBEN9J
6XW6+/CoMuD+aJTkpxZoHW3K6FwaR88GKihBkPUZY4klDQ7g7ft2W02/7J15F2p+HV8XgI6OPqdv
lxTecv7dVyzgutj2J/cO7NkYiiqZDBAfz/V8UQi6GvGT4jSKCP1Z7+yhEMI00dNkVciTb5kIuK7e
uhUBkT0B2g70ECGAJFXrPQfGqVAFz3CqQKA55BUYUDgKKt1qI6kaAy9z9boOOH9CdnPnjRDkr6Q0
Uf5pIxwn7RKMvFyaeXeGt766KLTQDkuoDiYS+AMANCytS8vfFFrObNpPZS5IhjcCuTaW3vFgtjcE
vIDi0I+Y9r5ICuQBL1entIiSAC5ctduR3RaTQxj5GFgNhJ42ZaMsZ8p/Jj8WF+Ibj0D2BPBf9tEb
xQW7QeeVsbQWY92SxAog2FHUMN2z8JWAPKCF2k+Nky01+ShR+NnhkiusSFjBfh0FNbEC8fkKJfh2
RDwjQ/N+kWHySP4qC+DepoerR0Rf7JeV5Wu2/WJgNtplvTFlARa/Z1oDcn7KVVjxhmW5tCh1wgCn
+3ehCix5gw3bBYD1MZsmiEVkB3dLr1hp39VebeNAfv3zhOln8onkS6O7R21TlneJ0CniLFGhamUX
kAmVJOOk4RK8IBW+7mKWPdv9zE0LIy3OdCug5IhyxW3CKvKVqaYssVhByxaMPLownhICWPK0i172
NJbfwRsoFOLI9hU7uQ2zoh9iqnEZqW+IG7VdkRCWQhMu57Z9RkcI3Ppqv85rjkZa81DpxfmqB2QZ
NBxFD9/V0YPmG3d5UBv2OgeamLrZaKZxrWWAKhHbWfxMyXa+uPGYOw2Iwl5wKVuqk1D1nskrM3U7
wF+I8gqIMyvFamg3xkMBvG52e9lmXL5fLF49dEzUHTEb3gQvhXRCkuS+b2fyabmWDlSkVr/THnBV
KN5OOTpMorqaXL3NdXJKYf+8lb1VvDSd4tNuauMHvtvs7wJ53quBFxWecg8gE7Ey8FUNHSj84ZE0
fCLJN7D8SMy9OfMp2WIlRdC98nEHovJOWUgl0UovPk2BzrfzbBzOWcHHW3sT7gCnlmCzhskLEmIF
SllcGbQMQn8lv4v54MOs+NEgkvBH7nqYixT0q/wZnokfhk/SmtX2aN6F5oshEASQWILFRb5bIf0l
uSLoJ2mk5k/6UJC4Q2ue9xSao+xzwL4zu1ShfjdagAM1yxipTHnVCqtXRsqEa3plRlyytS9y7elI
DvFKCgUWlxZw1ftUfFJGi+d8IDVf6mmZPfZXgrspzW8x4XX07FuOUvdTmTGPsghhWIbjbwAIn2H9
g9mHoEUfXCVdcof3RZ7wnjhbzx0sRMYBGZLxhypsTK9BaT/q0ZvtYHN8BGgxneQC0VzBhhimsRxF
3THGuvYytocfvoeAfHDsUdFNMpS2s0IN8EVe7QS73uYF+uL9jvMhuaNSrtn5CWRSClXGiMOLN9I/
Yoi/VEJRzVtoVlJhPgj6TDXTsyhJDqbYX3jAmaLxJB8sHw6yJc5VaEQGgFs7GcGH/CeNT2pxVX/X
/g7MU2BsW3UhwOKRyJLqv7xEX53zcIWiii0Rd6HeM4Mf2K+LRzeCQJAyKqXgJEJ2rdosUih85haR
/AY93slxRpSVy0pn8gg0LmMfe0nm7sz4Vi8cSxtAdQmgYKLBjtlBS3X865bYc4eZsL5yk5K9zv6+
pKg/lamJmzRpHN7HNaPnJv5U3WiW5MOZUB9G+BdcVLX5AdK93dXBeKMbg2q+ag6Rw20vLUv0gRZO
D4IBP9Fm2dxMbFNtZr4o4npp8ZVjnqkeRli9kZfO0Qmgv0MSJlCbcgHJ2D+0EIvwIGeIY8xZeiAm
WGruzpicwmFMgdJ3r89tU4L2J354Ncme2JpKxuGMX+JeHr6tSwIP3Ql/e9goUuvEX1QXLzXn08Iu
0S0GP8xurxQYHlTxv0fbl62U7U7cxSi6nIWI1hEcYSzXuNA6Otf4KFaOe0iF3gjN0BBJbZYR071l
XjUU1fFLBTVWx/hXrGCZfgkcKwgurDoNiRSP/diEwC6Li6uXLLEKfV1Mg4msRWMaYG6c4YtrqFba
kEbM0NntvhoEdaq1fxzyiW8fFbSvipRqQJrMbCEQT+TZTIe7oEAsDYpBlPlCBHMAHPZMWcRw5AAy
YdCoMuAeasG+MOv/Z4zN1Me1tivUJZ6csYG+InbPr4v0jsdr+GJkuxK1uurO7AuNnqhI0cmo3Hk7
jgcTfC9cb+A9ROEuUxawpfv+PaY+A6ejKvT1NxLAKx8zSYBwZJC4tdDttBqSdUbNrnArlRqR8xdU
tWSTxq+DCxIfGoG2MpIoLdUXjuuEbeN0yKKRZQ6faeu/zZSqN2+EHZ01o/JTkiocWpxQd+4IpuyE
RNzEJrtbsIXUr7egTo8Rg1A+EbhDBRcDAC+t3+iDDAesSeE5SgX5Wz0qVn+9IAxT0MjPt2zbgjVQ
TMcL9zSQJsezL9Uum18TlzAi35FzVX/GKC0ASwa2awtbzZIPmW6ATitI4pyfX1/gawdf0YrLclrX
mBPtRRNn2hwYpD1a1tMu1r/tOXhOZPrrOU7iKpQa18vHalCQVhKkaJ0u1iQrdn2wAz07Ftco7Cpm
84obl7mIhMBM//fJps8l/I5AvPmEsCzYz1Y+pZDNkGlRFpCOqoQzHWRPdB2q8mernlHCW1aIfE3G
y96L7czYQBJtebLlHH0GxVXbbKseTky5yPD5AjiIZCJhqzGdRjqK9th64Dfyod8Zbf8cmB9nH2uh
cULdx9X9t6mbtLrS7A56Rb22hUP8STKOcvqY3F7H46ahPKpN893nTbvHkpecloubmScSJXklipdk
2jnWkiXvJzTc6rMOpbe+oRVSB7U88mbmtGhTwBQibzoDV/0/SntNViZFwepEgGEBGOuGzg/efGSk
+tPsmTkx2KEUKGlgXn7ENVdDexw1S3VtsWSVf3oqz1yqewdCF0PywcOhf2Z/A3TohlyrDfg1p87P
6ay/5jfTUczSjV5bv//IS+yAmZkCF82Zz98tulGHFHVzBdRQerTvCZVvvsJb8c79m4ONxTnjKEXy
dbZFLbaXX7tQ1f8CKSmKcyDUQiI8sld4C+z0Esiovptgr6VrLm6SznC0Vba2odCY09W1mAEuOCJi
w2rSBUG8jVMTVLX0eb+jkx5kP5lfW+wpy71OzfsgkW0cGxIeTiBhmnUmVOE7C8qwVdrqjzlNYjCw
+FooBfi2/PkQnVJB8RlOy8xj6bPU0BfNxqu72Xx1FkzN1fRrq9Mm2y7PbvJt9/XSMUihBUBbwkCG
9aZD1/Jw6WkNMfRUSPqr/b+XaRzjLcM86JMCE+rlleeWhf7cMTjO66bLLe8lTqtiGQKyFuO1emKX
ARyw/oEC1/jfOfGVskZYitThnUvWz1Cf8zCav8Alx/gg1+TVIIJK6YflsNUkgtTyY74FjFqBHz/U
OBZBErh27147+b+oSNZRX7sNXInGlTBurRLie1HSOvzxVHbGZ1ZBXmUdoeaQIvarxo0QdB5VOa9w
Cx4ENskK5S1KJS8Ux5VVDyhUa2QIMJ9TFVhBvBb7xIriOBZ8TgWSqM1bi+8RVdx+YcHZDWW1OjJd
IAf4OTtwtXeAgFjV+6YQ1fow9WLaNOJDEkbgx83GwFljzB7kvZboG+Mq5K+lgiXfMFa426oLzN+J
9NHai3TcKyamZVKON7V18tPc4Q/B93RIlC/4QzZNl35uCKYW99+RO3+Zl0/G6AHrkYNUyqhG+4AZ
yULQ9eK+Ho2Qo2AD5RBzfr/bzJmYK32zVsSoJrWXig8ctfk8c3eLEAXJZWQVjh57fDe/3zgBIipn
6PZX5KioDPKK49AnPlqddqqwX91yNuWj1XkIk0sZH83WHuJsXhGxT8eHHcvbcSfWR7mQ9m2z5RN1
KYV46xzs7I2pi/A4fsm1OTZqjEliuNvLVsdE/4N3LEF9xgW9HdGx46ics3XYSMAeCxbE4ztN5XQA
PFktyWy9whjGqA+TJy+NLbi9l0D28oHsUnAvtaLND1GHSN7az2wfyuWZ2iUDJcyeZ1gq4/7CUHQt
nnVdr22yTIx1DRrrztLojjptzmCCKHXqslAJGBl6Y0zRqcU3SLDEU4Na/LzaBcfumInEiOwBsKGz
B/dFbXG4szdNt7U2isR4/aTyVsgahCOfV36T/NCwq5H1EAxYRkYiiCD8daNz50U9Y3WutWDVbI1a
Kezyf50Ap36vYa88oYCKeEnmI4Qew7WSGmr+LTZbjftDSKIJuKiwMf1kzicYQIo2qa+KqeJww7An
etLLSYyhUGSbNxQgdGBdJNc62R1gN/by6I1jRwNTnMLH5rIr6kw4ZGa8XvtTTJL0fh0+wvkDkAr0
L2SM+MCWSjp01hi711lvO8Kx9opFu0uGRATB0Mia6FoGhWz/CUH2xZYOjTGPQ2WqDjdffK6O6EW2
aU8+gSVTVmoZxBjrLOCWRnaZ6aw4Vx6P2gvkNvrU3AZg2u5X9TIDfxYfbAyKvlMfFfuSeH0k/BAR
JVIepOlzcDQY46+ccAt3zsi/3ZKJkfP9LVxXnQ3w4g/JeUH1AxM+fqf9c/G99YBXhu31YFaVps5H
P63uSqYMeubDVGlt4/V5I5PeOSVfo9oKuoHWr2PDMO3kYuE4SCI7iwOkz8Tw8YB++j4fcvnbEfMV
xm66ZMhaQjl+DxEKdyJZablWL3VVN5me22iFKnn2S/Fmfw2dKBfCGI3P7/RyRBLDW/5Ti3v0kIA+
fvd6c7ULCPOBD2G20+LPayIjmaydcKkXXIfDa2WNMH3dKIuGalt9gIEslsFvCkRxnrIdxXzbUZe5
OwnwhuDoGKnxOCC7RuXeHTyVq0ST0Mzn2KD1FgygxtoPPZ5dulqffvNJ/uvDnQXwwZJmgVVqdNsq
+zDotMYCjpA5HEpKbflPFSkihvoEaiuZErZgkmrOVAf7N4pK4PXxaYJ5jOpSs0symOLKDtlSzZ+Q
b6nOy9acD+lG8+UyRN3I64nNz+GSR2FocOrfmTGThHNbeXVxiWUHRCsjb6A+gJlmidk5PYgtgYW/
Sk8GBnX07VN1jZE3VR9aF14q6j+3ritNgCmIHIoC9mRzmoZ9PihZJBYH5nt8RFbugQmgxWWuWZ5j
EfG5sk3El7/tZHDkHip2Vu+u5LY87OUcSM6TkM9Bb4QsrdfJdL1as5bMV471+OOC4DL0+f2zdOcj
+Kl4XJU4L2XUiGdu+FuGRd48q+zoW8Kxo51UKlotFZMVjEFBoKXXmafYHsCmjdihlDO2sJO3fjyu
GtGvEQFqjmKIyaxZcwi767Ioj3VtYkikfA2Ker7OmXPxk3uAvy82Cvxd3e7jXXOh8iF387z6tU1+
3a/EbQ1+93A9pky+hkPygLr8ikqK50mQ2jZj1b24LcwGZQPPJ6wHxBc7r0SpPtiodjuFefNjlZgn
LzXoZsNADp7WQiymUZB+HLwUz/dKhjuZGfZ5Mp6zhEJ7uudyRRE/KnHPjdNj6kQPNDJI9qPF9s1K
EqIfwfFTQTWQ5tFDBYDCIJa9KtupXHv1GR6zFQgYsClSRogdfV30bntb+m8bGEWEbIrdhDRsCjWK
Hc7Wwqm4RzdjQ7wQYY0fBljbFvevOh7zhUOHbjJ9iojeziMR+O4xY5IepVcj02QtTg4RgdUqsmUw
zrusIKe8b4HaVM+NJ/mvJBnXIQsjBJV64aSWRq1HS0He6Z/D7309oz8qHNjVMmQUlM5MBxgSTyT9
ZCsjBqR/ZweqRhajQlQ7O8M5lyhahllnYQ7uOnxWH3HHb4fG+RQeQSzMsWPtGKAQV3i2Zb4W+qmv
4BnOuF5IEMsYCGW22G71ScZwzLSk58qeU0xIJwPUzXVJ/rHEV6zGatWskWhzld5sijGSQQlLEqq1
iJHL+aTxY5ILMOwAw+kXto7jtLy9/phM8pKsZ2o83WzAqeoYvjf1sE+ewQx0lXrXYiU6CSI4OL5Q
3nm0xfjO/iaXjzGOSvT7ZhQmue3WQYt69AHUJt5TZU6fhhjIth/ho9uehsd/JmlUTVo/izBTm8Tf
NMtgMGVzCgrKse0ofSA14uXWIsIqae7sf7bKcjG/TJB/jt+rT+mSP5TkJT3AoU0qAT3u5tPv2OEY
BUlnv41tl/DdMfV4VyaWTENdTbWedaqycKvu410a3y27D7gca/kHNOilRdhIPduR/NeNt40e/U00
hB6UYYp83sCqn08ReK/tHzMbwiKMMKHXsTIjRLomb6jZU+AdwRiY6+SiDo0Xk6dTmLio1FHzC/cg
gDYfhQQNGW66szk80OnDH/VR9m5D9ngDmIjW/VVO8GtTDD3kytxxhXx+FQBU3S8oOalSkTZXEQyR
C0vpIXq6SzqiiimfBdKRx9DoZjDH3gNw7z1WXBp9KgYUiGqJ75asTTt/RXdb/9tiG3p82PHdDzq3
/qgW9jgBw6u96HX/pXoHju+GkmiksrgtoGAFIJVSxkNcpXkpqlxqR3s6J2GTt+7etC8zhzviPboT
g8nt7R9nElNoctTna4ZF1VVNeBvCJP5ypk9Zq+pfGHyhvgBc9D+YGPnY6dWNIA4uNsyZ74abitSw
ZBGFhND59tK6MyidtehiASKfxASEsXOWQ2mAHWcjCkMBHcKQy2KQAIT8CJrWAkAL2yWg5IGKwEQV
TvWHM8Pr/vSC58GwxdNu03uSNq7SNZPMYiObzymokOb/PHb9clumKY2UWmCn+TMckDmPg+l7FPU+
k1N536R1pUYMIFUewiNMSJpHuDc+cjCV13sD+bk4Y7SCPVcKFRhwjLHaXDq/u8XRYnjkuoqbH/Ag
j2FhqaaEADruBTc5U12oMvCrsDh+RyOMaPY3raLe6g/BZVZ91zqkBH4qJAsSxDcxcrAEWnibSYvY
Z6udvpKdy1GYfnLxJXk/1m60fKodOepdhgBX/QmGeI6K3sm1BpviNymUcpj6Hi2QmbsNcBiqZkkB
H+ahTwm9cpr49Xw/12XlsHXCSzgca8ErIAiUCz9jX0G9E8ahVyAZyMPbYL3QwqEv7TdpodRt2SxY
E6JeTHu1Ch/yWt/iYw1OZQtYgTRHHG39tiNqBnCYStK/yJJU7uPQidagfpCa/oPwB+C+LgAIlDRa
IPJ8OwYvJVYAN3z5Wpr8GSAcEr+xxwNns9tni+evLzrPBxypQd6vFKcLvxA2vsXBiF3jSDg4FM/b
zsmb/OiaAHwS5WMy6/STN6JSbVV3I8TRkCfflmCf8aOXlCoyTl2azBgRcKqPZlAdt3b8bNx+kxYm
31dmwEgcrjJvu4UwfJJUC77xWWGd9ZcWBPBW9xJ07TocPnEIDyuTRphkLYd0CFCo/ZPyFYCfNY1p
XBBk5I69G6WFFzY6k0tNNkwH080OKahtL5RIYbAkuVpWSj4ftV2JrzWndrtSuWU1Lgi6UsNMyYFh
ZUv88j/Zp5EaHz4RM46RPyjIs37wA2GGntto5z6Tlf1vIJaRUTSOtq2+5iEPew7iEiGul1CFiI5q
qzY0ou2i1Wg7uWPF7j7fb18bfo01VOuWAdwU+pf+zdUzoDNmaSEOsPGQKwC9Wl1x8zEflk1pfygL
07lH8oidsr4u1EEu2zCZYJPk4FM3wcACLGtjHUjwkEb4V4xIEttv64D1vdaDl3VgiRGcUrygnwpE
zl98WHtc34f+frlUshBgGUXEqUD+Qjk62Jbqfz3n2THO/IAAmHpzq1Qd013VkTAI/tXRb8/zDz4y
t0fnUlrS4W2r9CNxvHnsoQ8KJclJb5mEEncmlNZkWQFJgKvRmPM3oJanRUznlyz8O+kbOa4RKvDK
5/LvGbSDOkXDo5a8D6NhU9Q1u5FJLAJa6Lc7weZDKRzyA2UFWpB0JA63dzuJxE0EgogslR3dSl9V
VtEHT1wqTGCJ8NmHeK6EyOT71A9KuU1ONRoY92RjfJC7WMhgtMcB3tVRAdgCjmYxfoVvaAfw8Q+T
meT6fXwxzGSMX++OPGYZzN/mFkheAlpi0gQ613IfNNWpcnL2RMDpLZAw++yxCFGMkE4CiQCNlxRQ
nragp6kC0+duJUfAdGuxedONfbHCSxuw7Ci0zky4gEnZcf2g/hZ9b4sNpUpIyYj2rxsd50d0WHoC
5tdW95dssjBLYiru2EJJXuyvuJBLc07DvHFcMEnB4w2nrl9Hzms18X6oP8E4Glmhy7yEn5bnWV/o
ys/1m1GnJ7EUxUMymbvlDTNv5eoPiu7ZlYBs7+TABzzxOvsMpK9P/aCadQdRTZBpSQYUrKYQIjNj
mr3c/8TBmRwCWYK6r/fvlWUpbF7SRo1GWzmfD3Fkdzd8jF3/wHFcXy4iudLwO0E2UG1R8doOeW/1
TsKgEo53cXqEwdDDwLS+4pGcy7gX8Vv2J6R9kZV4EJ4vhTI0LaTpnhJPpioM7d/0TOPTEc8Aw8cO
JUPcLEuj+RlrmmTQqMpP2H2rdC/nJ45fNncqneXodkHRkEafhCnt4wwuiQxtt9b8fhmjOJJmTOrz
D7qDyWto3X+f25F2SbPD6/xVPTbO7ZK+MOSNxqnu47kr4BtkLf17gW1Jh4cFOrCj64LpLZyTDjHF
KSqzPtwo9r8tXhYWLq2i+Ttuj4lvKKB5rEkhf6hYP+cfMUI8k9UeY9sx4AKnL51OnOGPPhxPuDA9
OPH5e9gfm5e3LxBg24HXv7At0vMCJA0FTMXBSgzQynSImtf4sEl/PABXD7gN3YJB1xd0dQFynaPn
IqBszWUXgFCZuLUBgZz/jU03X3uc12fJxh2Vad1X71ufAC2T1J63SVWMCyxxmUhzJqiZmXiwkIi5
ZdguhTTNIakB3dWoG61y5NFnaej+r5ys4bEfO25PigE+RSx5PmpvBNqf7c8Mw7gGyOowc8jMClCm
mSvUse6uvLE/Z/ubV0PeWl/uJj6Rxa4tI0S2EfNWdyP/B9BAVI8tGQyhFK+WbaipqloxfKkxvw7g
FQcJblLOUHaGXCzxifAyqP1sJgUnmZcPtfFyUQuXsJytZ62CxU1LYT2O8C9T26fyUoB3MPEWLlrb
Moq0X9hNcqyslEYgZKT93uv/C9ZQtMiRfu85Fm47pICUIZlkjVCD/lftUxNGgi0ZXTrVOYmGzym5
BjfdtIRXZpyjLEe15wShfrPZZln4GuUtAbrc3yRhViGnlIKKUwcejOltpFw4jXnZj+o505gGmpli
FGR8WXmsTYN/5HGfPJGKRp8Cz++D+QMMVjU2iWfLo6H8vRH4T4Cb6vAuyvrK7kSbbcLVCnrynBwZ
ToFSc74Vbbr9VLis+e6bgY0PoZyc4eL+23oTb+0O+qGfcWFMq9KGGStU2tn9R1OpYwkbcYOA3WMZ
/BK+opZev/IXTz74rF8MbedG4fX/ZGR5ZtDAD+7CExGzGUMjwx3VftSq4IlbTTH2bGrUy4cZYjIe
BimguoTdPRgFfyCCxM7nyU+yNf8zUXVmkUgOpRwk7yauMHvDBXIbHZJiXdYKxEcebc0pbwg3spF5
N2mt0K0x/GKMW2na82r1w7J1EUUqg6B9RZVpGAhsU7of01jeNjHs/olUfjvBj4TLe3JjRi2tIDuP
NZxD3VH9SHAno/aJFdUP18flVapN4ncLT1fFgRrnVTX/ay04Z1ANsKfVDgwhDRZ1z25o+JJnH9E2
xBq5lztCthNpx9O0u+J/EsvsGOs0V6u56Tqbb9Vh+YYC60CgOAAV/RpCUd4HX+5X0QjjkvbmbJlR
gPEDuK8o8LpRvwkicXaksEwZJZEzKlodaKx9xbHVwWf7UHI1lqVtI+vqLACB86668iIjfm8mpub7
dTqp4ml8g9GaF1ZR0g8bP5N32sqXWYIAL2hwcm0nO89mRoVOiOan0gN8fgIexc4YhR8wBusAbZgi
nNkwaU/G0r3PzbeNwVa0Ow/Cy2k9Mniv2dLwM5SsgXO/BSTR/QcXq5Gx4Ed9Mq3UxjYTbjhnef/9
jz36xB18LauImg4h8/HmIKV9pTvqui77pDNA56gI75CDsgV6PsMUtBbdJrHn+G7ynDVqKzkKT6Nq
kvB9x8/qsC6htf4zIkMv2sc4DV5+em82Y1UgHDNRU4JNxYc0i/4ekQ01CBg4zZ/0I+7X36L4PQam
lRBdWswweIAkiZtnSnnvCQTiFDc+bnrLGRidGYS9g8ZO8L2hE9IJvD8pnQxwzoMevW/B73qBFpHc
gWZQiz8JvAlcMnVPKL4Kf3/5abhW4zomezu5MvJqqMkZIDDLRKaLg39rMYqjjRVVixAWcyqo/h6h
EuuYgWzEPHCEK8RANxP1P2Ik6m9+Iga50mnrBPXEDzyZMAFX37y19R/n8ukxzzt2F/jS9qMJPEAJ
j6ky27ltk0IE9A/T3jIeSIC6ggz3PMQXlJprn7YPd2i6B975S//j/rL3n0+4JcIjvj/Txftn94/n
zPwxv99OPxoWzJqLm+xs6Q45/STfVL4HCEUK3EXjMq12Zyk+sEgdJt/EhH5xkQpMh5dABPmYDf8W
vrYYk/qolpNaiiRXyibW0kFioD8gPWyzxDxmWMcS2MLE2sc5lBEaerL+4A7O+gGfdwlFzwLrdZ1z
76kGe2yzk9m3I0Q9yKcLuCGRQ7Fl5wGvLM4sT0h7nQlah61L9ePqhXITiRa2lDgeX6kmq5dS9O9e
VB/ql9UKKTbG92/LRgJ1Ch/vFcJvNE8NvP7avqa+JkYsmy+0LhjgM9QFE15g1K45L1bl4L/aItBH
pUPYCRgTFFHGEbOeS88w1VpCVpGNYUNQ8dXxfEX8pvBVWujqwWp9s+2UcvjuHqftx59idR8ZChKx
d/jiSkCLfXadwxXmBWOynAM9+gwHiQLbQosoc672Jyu8jfVaDogvH71zw34hhMY5vYNFBWYpC5z8
5Qr93v/bhqnGYWIDFZsNul5/ko+jTo+3bbz/AMRcf0yaDTQGmqpzfBgqs+dF+TXt4NEXQiVl770I
eSNhvPZx5ZVjphjQrIJxagcNpKieKSzJbDIbMwCETNf7As+kUmp/UHJPJyMG1IeBGpEuoQcQfgBZ
+XXeRrZt55r1DlfUSVRF76Q3ERGTXnVXuzm/MMOh54uGk9O4q86+G22vIWYBDPLmuF/VYzDtlaJj
AKZkRtWvwkNOv/OI+kgLWKvu9laJE9sOvVNmK0YmkavQb56J7EeUP8xMUgdz9+tAUrhnQknk4B3k
gQCiEBSnFAtTuyBymCRoc7AVzWc5S8I3YRGoOuj4T5++sBclSWDYykeu/5Jo72SO/MctOE4ZhyP1
xrxSeh2ShhdsigM6UMJcZfD0+6+hWiPRj2T+pLaIvm2o1Cj03z1o/6YGLO/ASxy6pUBo1wDilzwC
Mn8XZdqGsgmO0cHNJGGo+z+A6h7Q1EQiYA8UKYz+jQy5zfQ0z6d9k8m8i7fU+3bj9zc7pdjIhhmh
B8ERckkwWYGOfnJDvWWSmnJJPRqU27mtyOeJTuHC9crhK3W+bIHR/IdOoZYaO18yNxoj7PXqZYBq
ZLRSFIOI1uTqBGwjLkPdIiogDXaWVZH/zjb2xkXYWP/QEd3N5sxErZ6kLVDL+nW34mplsaCDWyC9
tgE6pr2MMXxuMuWK8bCfleW9tXcNEuWOkVhQAzzSr0h48jhvzL+zoFVsrwa9U2I5AozTQqd2TiJh
PAo+IvDtHGE6Uva9fh0Y7PMPlFdMMg5oFc9kzVxbKVhMzUlDaiEPZZV71T26hdfrkvTjhXPeo6yC
FHpuGA4JYcU0CU4lC+BF6/sdjQYIXlZ6+kdtzTSoBvwHdRC96Y14KqeOPqmObcxE67K9/llOAQu1
dBkr4eg7uMnQ14XTmUvvjh7O9t5wBYRkwKmq6sKxXV2fDkQ2mPcQuu3AmFmemBjcIYVxEfbcAFRD
didm6eF84Xz42DOQmTudf4YIHSAovPKBYGdtKz7tHEwDmoQvlFX9d/X4gaO0IOHHA3yIsI67OXLi
RENVdoEQm8e/+iM1LuT2oMXqSEq8AgPJ4zBXHEvPAP6TuNBXcpIflG+NMhska2A0fdNUIqfRGYRC
lquh8/1b9ydiQnvULaAnlnPFGksajlYq3I6dVL/ooHwpsxhPl1cDiOiCe3bX6/HSXPTm2ui6llDB
bECmgF2xNQUzhhcN7dBIVZuj9/F9Y9Ruj/yY2lqPo8KSqKdkhatJ+rCxBnwyRow0bvNy9UjcQtAm
aWO5pvbVS5yioAsxKmnJpvORcavsP4rDYfBgfmI19EsfhO7wOZ62B24NbnUFUNRrurxjjaa5ovlq
zOMOTBYNZK/Gl0HzRhM2Tulv/oDqlW+k6wCp7GpVfW0/zX2zeHMjEf7NpP+qnSwKvjjFM9Rexolu
GGp3K/KKHdfuvpSsdHhNNhJa8n+Pu+3V6Km83mtKt+hVxydFTMgqPU4azNeTBy05DVHpQ7wP5xeX
u4h1zJxfReqVyi2gQYydf/zpvQjTMc4G+EKC8iBvyOW/cbFcgv8DNw3PgZAYKGjacLGmNmCGwXM8
zzVDTg0TbQT7u1bk9Yvgq3Wr2ua0+l6utTPTv832/+LE+aOScz8GRjxSxI2mnX75v8C/B1sNKHN4
La+f+XzmEbcWf3FHOspZ/BDT+eCDdicSMsI+UiHnYYxO5HYcxiyUXqgSXGaKEmjQS5udgnClVM3f
AOo9SgHYLCxkg1Wq7qECWzR5SFUFi8pYrHTVayqySjRtYV+RMDXIlesVN5f5x5/IPtfguQI3xiXU
KP6zGP6OB34GMyevmyrrHpy5n3AjI3ZY6XtgqnTczm+pk6LQmZdjZGnnhH8cLhjvHMvpbso0+qB0
HTM0wYCQwtQGz4lplb/pm21BAGFkuPxE4wQ1c7RdH4VyuE0iYrsM3095MjckcoT61akJ8L6cKjDk
cMml4FzrlSWuvSZ3kk/WoHtRMbgAITjhzZkdzwonHEUvZIEA9Ak6n2L1MoBIkbdIsvNNQ3GtoUvC
yPY1gPsBR/CwyARvmKbLZvxIwiZe+qVkTwOGjOq5SjJGT1HljA/Px4onUJOzw/gks1EE4DlM61aW
2xQgJy6/Y3pwtA4ySzPhwE5CX13xEh2DXZNftRiedgHTJNXmZNXL1O8ayL74H0VqpDX3iAuaLoRY
LQJfCRswAUqC3+oZZRhEioo0u67GB1FVjJvM5Hmmb8H79ANvKu2nK+2pLtF2jPSnQ77484G5spP3
bZU0IQCIKVJZQhugv40Zbym6Fx6E/hYnBNIMQWkgDoVldp7WuYw/A99K8LtMX0ZQ8RZqx3QmtrpO
xFlq3LvO0ePKUQgc8PS32nGcrINTu51lvqAeEQPoUkzyO57hku2ARQD50lLkThXiUd7M+vWDtGR2
dSHd0n84r1q5PwkWvV4HcQkQV8acWgYLcfNX/DKqPm2JhgUZAQCE6CN23fQVPcF8tR/f8eo9QVky
xeoDY5QPYKgchiMxJEofCDXHmDmXgs+IQ+8oNI3z6dtdpCeezj9sfaRuhteWVXds7OZ3O0rATmHz
DvFilaZTYP8vv5PXBDzgMIz4gLL2bY8ZbZBuD8Q/eyfJnRvG32+vLbRwsbX4+fTJwpacyq/X0xMH
0b5dKEm30xxVUB5taV/lMoCgH7fE22C1kLRKCO27I/MQXOxBpOdSlixS++yhlXylPLJ/axTGJ8aH
t3kG/HUn1r6Q74exlraGng/ORFP0VJ42byqcwH65fO81gGV/iBPUcdSMTVooUyvm+ADJLWpCYTlH
RxGN0klXdN1HJJC7VlL6fB4kTPXSZeA2Dy7uYktOk+csUQWgKn+1YPbpql1Ad9VggzLD5MmQZL39
aQlJtrgCSL72Qs/LrUs8mvzHoiR3I0E465JEjI9LrMAxX6o18Je1A2l+Hm2GLIzYIRAcOcBB+3er
6ULBOK7kmNf6uMtxcJtat84E1i8VApZ3qnM16sbx1eJrYVpKS8trY2qKUz0qcT3MLtSc+oaru1PA
PYLB/4mbqPmCs6OYSteG4kbjID8mfUVaPyrxtUdj6cL1rlntqS1LOmEjhZI4hBZfUImI9el+Y0I5
/vvr8g6jQrIJZD6tIUUMm7locaz9Uub2jWiE0CzOFzsuqR00PQpXZJAoNqa0vaFdoKQyAW3MdqWz
ZmIeO7n1DWlxgKUXYVgd6NWH+TBU8sL+Q4jOG/H94O3cLeT1vtQaOMw65DCLbyxrLwtcdUc25wxw
qN0L/DL+NrBJfMBXFSiROOHVWft/w3J6WmJbb+Zmo4iXSPqNk3e6VK6kjzfDvsn1HHySF0qsYuaD
1FwMaO4gxflCp6QWqMOdooujJxpoagmqYtBT/0C1/4+EtD28JllUTBX0p0Fxzb08wMPIshLBeHy6
vg9t9O0286upzlz9Y5bGkkG7rqs3NwGZkeQjG/AxVG+xFs0jBSB1EZ/QRKTn5r5vdldZpH+ndIXj
bzc+E7L7c9qBWkiYkpaYzwcsOsdnCnR7xfU/7BDrMqDha5uMxY+jcu6GDVM5vut3CuIu3V603olx
j5KmKx1/Nkomw6ivwolpJohnHfWs+O/LupfgxiRmbMEGMaDqZ28Sti3kTJnUJZ944mWHC1I6DToe
SkmQri8TvdvOwKAh7Q5iye0ZIY/cSSWuq1wjnvZARYBMYZ3WmZrlHaTEKsBpamZRq89EkoixaVMo
kTZTrme9UARKcQ3Ous980YbXxEd+zIiDJJysL1rhUjzjrBkqQEYMXlG5bf9y5Unc5HCc5C3P8y7B
h9MVmv7HTOxTRhrEvsKxtoHy/3Pt/qjdmEwqsy8yoae/b8MBZNWhbpCgYEwKwSKvkhRXd+2EZNOs
3W1vmII3IJlodl/PKH+R9wqBUe5w4fcActL/C3C5FwnhoH6C3ICJNM3wbrnS3LETRnmquv+na5rH
lJj1NAb4hGSsf2z3VXDUGdvtvctctcGyudHCiyhhfl5R7TnRfxD6oeX3BvgWrnf6VWEs3xof21XN
t5d5QMIiNQkL61B0OPgRUrJTPnMNANfRIDAo+2eNFPU5mFhHBZ9WBRk59pRu4F+IiEIpyZSXu7rV
bOHOz0mamavjWimUtHkYS6yojNTno2+Ew/JlmTf00X3pcYGbg/nCpR6ChHHcx2jHMnuNfXMd33Xd
OTuV90uzDMa8Y2za1p5rEtSYK600jwvMOFVfWNnFYRP3buBBqYmDEuyEPu4+3v/Axm9IaBwJu8mF
Q3rWAmQ0xUiFxGqDCPB9dkA2eIXEnKNNLwNur1ap9DtkKzFYFgPs8Ajo6LyjLHMl++WjEWeTG7C5
gbF3haLfUAoLAerXSxv6EYTdr2A4MmpYRgpxHnAqJWJLVyB0uTGoTDdX7dQbMNjMxX8cFgfoMz/9
Zrf/MsFVHsAMjJd7HeX3TVis4I0KoWPKZ0znGZ0jQNI7KDzKa+3JFuPJFbMimEWAbVKG/hdd7sdJ
ddD4iOA+y+D6OBnUE6kRA3z2LBijLiiNyXKUJKYg+taZaFUI8MEqDcQgLLxvlo8OlReAm81Uojk8
+PkblwlkSCHKD3NcIvsk42We+9DQMvKvxRCSuQYYY7Uk4CBg9syRjEABXBk6FFVUQj6zupCu0QJ/
KOfpPXEJjRJZcgvst+M59brDV4z7nWzrZ30IEG1dhrMV4L0+91XC6BMXKJXTvPzxbSeyfr4GGk/2
QhYY10FX6vR2APaUjlUmfkzWMCvuRUfMRBFI0wF5ZGAo3ihq5yoqNSiYDMRW/P17LQjMjuL80K3H
EUjeq3VyraTL772sfyt5c2WVbrVf9PR14fycFkyHZrej4OP74cgX2BxvO4uTVoERH1gRKRHuFYcq
dso0DnVAe7eH0BmzLR8cyxY6IREQIGDtvjscBuz3idbl2Cw/d201kg6gAWl9nAaDPWNnUa+tnOfo
kZGvY5ZoXvEj5tsQvuxPtjTyuQlVNUhRvKTHxpaKpxPta9hSeVItOb1uEngKyHAy8c1hS3MU7yC2
GAC9g4ZTa9X623CYCxOfBye6IyGVfc6xS3TKpI6wfuDEocNTnXbK39aYPv4mk78fk9Fp4vMmS6A6
UwZUA0E00DeF5UsRrSBjPkq02AEN77juoSK1ObAee6Wml9ROG4/9rX1KVL9WylLj49r0jU5hYCIl
JcX1JKmrgRmRguRAdVgExcjyXAVzII9PwfgUsqZ5wPTxUuNdK4jQb1yfPSJ2ATeDBFuFuCTsDLVw
DpNBxOlLd3yGhZoPX8lt8QjIicsQ14GffLqkrfkBUngE1W6H8+tmC2RHre77nvF1WBtQU1k+xI7K
5Hc+iXzKlV0OcHF/Nl0En+s992gEn++u9KmA11OmpfxP4emP7dHZPwvcChGMU4q377PYCAsgpsKI
z91FTRo/LMQTvdGdW4F/u+g8CGDFv4kGt6p/xJjvgQbwK3CA73kSeGytXZTEbj42GeHe50TCE8nc
XOhnpcVQ98oxwya4LfDhjPe+dVczRY1wTtlJ/y7LBmj7e8N7PTQ34Fs29u2Fp+EqWgtCFaIY0h7W
GKT1zUc86tu3LvBMv2JCqPzNDdJAZzcvmm6Dp5NZgh5dSzMuW80aLvS/Fa2n+SLNlxM7yb04E80i
5TOhPi5LaoUDsVhZ51DC8xWQXkW2/W8TlNHLsizMyvqGBJLnZ6yt10ZJo+rp3PDIQt2WJ4l7Iz2Y
IPuyqPbBt6LY1937+xyHtLrlU4tlYnknNH1e0qFXhrlsIaEXf0mMgg5NKDK/mo1xxsSm6E3cGx2e
VF9u9VM8mFUWoevtCUZl2Zo1cjFTHjf/TqAyQcDhdfHVM7nZeQB9yvzyXXzh7zYKeDorKcbstPo/
DJ0dXWNfttVYlliNhz24f3TWw0KCIy7JgSNXpVqnkN+mA49BspqvPZDRpegaloQMEMK6O2coHmZ6
Qyzge453rscXmRsEqDBOim36qOnCRqQUOBcEdPSiKDhSOJ7Ul8YmMPSW+WEcD/LrGH5m+tulLsRb
pDlPe4a1BmUBIX5eR1GXQqTiuukkSVGdEMIl5FXRsZ6+p0JmptTO+DO2n5ZSFhDixU7iGkgQbckE
Zzapbb70ugntrfONg5FjQ8DBi/S4Qt2Y5gdv40UaoHa0Sc4ODOzG6BIQgRPPPVawrAkrjEQ0YveU
NkdTkTjLP+KcMNNWCwLtl9abBKS46xd6hc7e/gqJgz6qMRbgbM7keYRB9nvJ9sEqDU8ejbpsYa9D
V3lmUsCDhbogjJHYbNfCDopbohVNP0TSC0Isx52uERNY4ld/AfL1XOG95YlcK7AaV4i2WTnM6XBx
9w3SZMVq/tIK3SZNjtwbeH8Bs4T1LuGQP8SEsdErUYe44qLrLRZgjdNHK2mbX9lTDlSu0cSbQn2S
Tuk3s8YaitIo2VEuFMyQux2llDPSKVg34OqwqYRBeHoztfkDofMGpMn8eRSNiFP6wjXckD+l6z9S
aqzP8lzsEAZkNXSJ4JfdFaDRmx8SZbCJTDqpnjfjZ5seUILxJN6m2XWSh0QFT8YHeheI2YOewVXi
MEBVBegx/cejONRwvV9KKUOBqMR8QSIP0ezhSuti6ryHHndasAyD1yd2DI05bUKJu7F4EXdwQ+3N
Idq02K3awzWpxb9DTclQJLOeol1gfuVNvfJE6A+FmonFUZ0ZqpR6Od7qXh2soQIWiPOC1ANdhI2w
ySSwc6P91Q15x6dGxAHlx9MRo8bg8J/2awt3x1PEvNlaPGBdnnNWdADhykmiw7RUNWhKAE1Sfz7O
aLh8Xz2fvAVTsjaVB5Ufs6ksATMMmFsTkh3WMQUrs8WjMGtSi5SVwVFUMGIgQRAUbupC5j7iyHgQ
pwUjNjdKH7mYp/98Vqo3T01lhOJ6DBkADpTRxXl5IoWAzv4LrzZQ+xgG15GLDKs1YXlkQjONeYJs
7zfGLQgvwrzdWMw8i4bdQn2uo1E+7p58NncbVDC5wz0RNLNe4oA4/cvfkcEiCKgOOqxODiDAHnp3
q/7t9/QNcPS1HGIvQjbp5Fwp758SC50fVQKpLu60tMT+sn5doQVw0zmkSzdVFHqaxbs6tVsaGvhZ
zRC1AnGf33QB/ZNsUmjpDjIzWC2Ze7E3O/jP7mEpe7gy0XLf+jGZ8prgKvQZs987hM9h9P/TJiXC
wisW7k3lQVO0m/OwLKR2RwFfeb7qdYmlcP66zTo43u5PH7QzZqpES59uTMK5R9Mr32V01fuINtFL
By77AuQtuUbzAJchOWzu9KiNn6aSIIFDQ+loO6L3s+27a+QsWfLD+Q5LLB9AsFVLtREcl5LDfceh
Eafus7TqXxs1JlQBVOOHkcFYMbimzkyphBghZcnBQvm5LjlWH1XMXAAi27ZmyFupwTr6J7vdEo7Z
uEXeqmyEKuJAa6XZwFbGAswHh8AU93fytLQ/AvEKKS6aMHjUyZ2btshbp0muZxznGlJLsQecUrea
MfYYOF3ntVGJt6kLyZwm+a2aUmlw5yX03Q8QygbJCmhccYig/mu1A6LVWlr+8rNangjlVD5aT/zE
yckd5gabqh3tZSXTHSvrogTqV7quuRYwMJHKFcTh5UQxGkbqXLjFSvPL9H0VWGRT2ZMwLMWpiF4d
IRBnqiJM0Cp5PDGg667qNNhgi1eGS8uh3yGFwsWJqMQT6PouCsCDtGXYeSdO7E/lElk/ShmLgRoW
Wj178WYcYirfv50mZmmI5i4smOrViKRH99D33fzL8U0wxiVsfdwvPljKrMbuxMjhnXKDGAzCBRlF
YOalJEvZpK8f4NfVCUTA64/oujk5kixT01NEKH0ftj8Np4EIgQiqAOEM+3PWyjGSJ1uzTjuUHCCk
vuEL0mcYyrICUtpalBg93HYeOigjpejGwfSPwx99vdEHCRi++SRwe/yLwlR02BYNXIOQg1thXyeC
h+joeQqrFTwzBhD/dPQUZWnylzuJsLneu7a00M+DxBtTlaPQU6ewdmSfT2cXNck+JG5RjbZyXPpD
DeTTmemVQZvJkgmXNyyhoiKJ5a6IHE9qm20S8E8tUgtdDaF+dU7++URh/Cbf3NfgZF1IeigY5fDc
dpV3UUwZC2bzMtmTvLl5PpCWHJJGSRvQWxFEzQ2QqV4DZ90ZFlAQaHGvOX8eoUK6zL/w3WZyucw4
PbFi65vVIp2xR+Gmj//JQwaYs9D7ZJzRiwbkzRaGkr9ZtNkl15sJffX5rApbvK1TEv8dg6ZjvAeu
NivA4IwUJoIpawabPf9d6xSGbJ/h/gIZyYIKWiuXVYVzucgTzzXHjZ1zrRkFYcvfTY+y8sEm9BY9
hfOQzXqrEX2KriF6AkIugWWEjXPjPGGy6ieScXLqYBeZRwto2Hlp3SVNneDOMd1X8JNZiVJTxX2q
XckkVybesp61S7B3V+5u/AX8bYt4nYBHHkJScBiWX7CYowryQ3+Prk0w6is8h11LDxtZ/hnE0zF+
BiKApI1+upuy3BrlqjSkxKDxTdJcyLM7ykzVFAyLqAKUcZxH6IfUH6u5MgK82z94HGaeCravh6YM
IZkhJ1arcoGDwjcZtS4SQGgRG1lbmm+MF/sIYN8P7dnrpn8jXTpmMtHCAoykDkjG+G7sQXjfFFZm
s8PquNye8MSlsvq3IsQMYJS5KWtyDoispFIaCwyXnGMqWfQQQNcHz9Ri2+cTatIkwzVRqSA89Tym
TUv5byKUrSyAGDq/a/MZd40G3JVDcpWVN08cVKkOXeghNrUOk4svTTG2Tu05Zn8R0Ap7OF9tcqS/
DquJQNUaWcVYVO0eIFZZ3OkyhLKTUUT0O+xL27NG/8ct4lxZckoCxdJFHsXbRyP5xqB1bxXwfEj8
+bghoFG/uT4cUVp/LGQMoDtsUHnzb8lOCgqChgSJwQW1d8TdLF+F/VrU9/5wTrw8qoT86Ouahzhn
x7H9FapEJd2qySGDvvF2oUVwV1BxxdB5GZ0WTT/FBiAP6tWbcebD7q8+v2Pt548prGW9B+oCqMVB
2FddsDliBHZQ+3yPGIsAJj/lXr1qu6NPuB+2msbM62UDosIqHbXWue/GcVzE880dIrrfc9GxDKWe
g4nrIrKCtxLgTU6WrV0z84o2MJViTQB8GpqLeWqSJE/GbQ0nHYeVhCpwjd+OwEanoeqv91d4P0Gb
8m9f0GGZIcqNpa6FCwYxCP70PlIpisPsBXA2CfRqxduuOgzaoCmSRN2IHhPbwvaJPkTS8eD0Czuu
/HDARljXBumTuEcKRW2WLpKXeLuDK7HlJKGAsptoT0HXizIjD0+a9Xk688SVyABErWi4FbM1OIX1
Zp8dkCGRSmmAzaIOZ/9VrW6N+TNXV2QLV9GBNAkWvHwI180KWyIoyrEYaXN8R7piWcfwYvbrvxSh
Ia3MbESI6DjxCvt7PYj/flCcRsnxNXrctGZN6SchH2iUJGqv4/EOJjLJy4YlfZCjABKO1SmbLeKl
7AtIE+At9PmJkco+XvqLyzOVXMinzcC5kVZWyqmp/BUJJ9QBYIEHRWfIBIZEcIjgd8FWKOvM2GvX
MO/7kE0BaSX4mjidTx3Nz72/MNzA4XC5XfO7AZHPxFsxMjUQ2b5flrTb/40aOmXODIap6fGuxO+A
uQbOZulkBEjpI2iUWWSu2WXoFTZ0xEAZNegiEd4zjj/CUIj8rRGNMSfTbtVC0wQkNFtL3NXjmeTR
ZmTlgmKh+c+6BedTFmPZhJ3Gd0pTQm9oDJtVPUsBJfc0nrqK8NERz5IldwCrBXiJJWoj05RzNgAM
PBEwXEhu8RSC30S/UW/lN/0FpweWBpsed87umERJwGuODoiIsIxfgB6vka91sxA9igKcO2P56ndj
+4HRDWx4cDyOo6KeK5d8qcG9adE0mMYbYM6iMtOtyhzxZZLs1MwXBUc9Kk9GfbybyifppSrI05k3
d2yIHBIRq/ti9lyvVwQC6GqlUWmMgqoDPL3lPkS+3NHq8LVJl6jHvTCNG9msmK6aP3t65IqnajfL
iYnU71zH3HrfcsKFQD6si4myjMi8i0/Bls8cpX6VIkoFgBzpfxKoCcYiQRTvqolzawwV0nHIE6CO
ZApnxEBBSH+IYcrZ3LR7hKEco5qjGPVQyzQBkrarVw533AzNrgw19IUXQIEfqHsuOxoTiwGlR/xI
pe9mr+3e2e3E8DPIjNwCC+EHk9zqk7myqJGD4D7fOG7pKcHOFv8bp1MHx0gOlRXO3c2BfwZLvJD6
wiRPUKozx8e3S3gl2q38Zdg9kE149QD4Vwn60sS5XUhR5LwWLu2Tq/vM+u3ONIaanPvIX13gnCWA
3ZJieUnVsQFpp8PoDQdoSYxo9IzDpLZi1Lz34QCXo5Jdrxw+pa0h8mZy2yArTqPbOzxrfvOjUsQb
B0Eedn70gygxRQYrmmG1tDpRrL1zhJtMO/iErpEitfi089kuDBFwAG4nJnUlNhP3oogtR675dvjw
aPANhFTTBpMskFNSDeCXT7GjI7sa3jY4hIxJk9FLSEOjB36aeIJrpB8ZL4i7Agmxnp+rr2pX9GSZ
epZ0968IHgoQ+vJM95YcGwEVKhzkgcTfh6DUr4SeLl9BP6riZtfWgUBoA2ZS4+NaZ/4uaWkHeIbe
llm0d0po0yF/j8TB6oNUAhAoU4KwyUJnroqTbkMzywfRtv6vFgQGzKEBMBq5jFrbk7Ww6sTC/FGg
NuQI4f9vjzQ6ZxeG3/j9y3APXKgFIO3J3G810bBfyZr23pjszXjBkSx5NitaNoG4xRIrxZLkDPPy
hTz2GHk9Xd6A1ZSutxeTzmPvSHrU1lQYOpPqQjr0cBp9mtfZN3wLswHDduxQtnz942VNCxP3EdRx
FwDP/7N/DeUgX3dGQuRXvX3IOujUkLZmNFiU3HUVyfsuBwSvO8xm7OmukOc8ZZF1p+L1Ck+kAobi
xkm84MKNepenPUH2es9gIegPPnig6XmieScAklVy0GD6g77Z06OP+RNmFkCKkbrV8b9ElIlHq/Zw
5kShakChq6Jdujp2ixqOk1kbCqjjUdysFE0wgRhGNkIDw5DSCaNmDk2NNPKSpF8YoMPYuwlYJJ9J
KBhccuFvP3Fvka7jOkFMzbidfR43WgZYxg/M0dayX+I35yzAb7cHnomlW1+RNB0B0LW1uiArD23H
9arTJxBZKTvVOGNTTjd0oWAvTG9fT48gfkmKH5DPn/sITAW2tZvqMqCrjEtPeuK3zFPLcqmxbJbl
+sTBayMm3oFiodp4Jj7A2/v32przDRM010O+u2jSzcV6tWDIKJS3hYrSd+r51xbnfVXZw/8KsWGb
VdOBfdo+Cjzl66xJ8e32/Y5fxRcbgZv/3bDNH7k5EMxMPhdMLssrkPGW6SlKKVAJJXpNuT66Kiix
ot1XYUozY/B/nBlEZ3uusTxIuYPPimt0DnmwvOZofUHfYCFvTqKPXuYKqg6gbkJwe+SPGF+BZwIb
6eTePEJGEjGE9RHr72LLZqBiGP1OGrnFoRxgpBan8OoKkXpf5btxAKUIowPwu1vjB8bRPiGpdX9a
y4UvcbL/ANKAMk7nelexdz+gNQtwWOXuLxY7oXRmylwwBgZAiDfGvsDtahaSB/PnCQR2GmlIl8fm
dPbnCGUdnwUDkHYhwZKTCXIzVt/wZ7X4T6dayGkn7YT8NFy9Loix4EDDuCYDOuPVt4jSQKubst2v
PVE7U/UFWjCFaLhhkVw5aNyxfo4TRMeMiEacoPPHtolpZdY93nEIdHN9eeKwk9Sd8cEn96g442tC
GcWBSlCoZtFkcP/globA4T1P7/JyPZFP2+vgst002ZSLkKFL5K2Aavq4Lrcj6YrIQG2Yx6Knk40D
U2RJfdNVNCYT1cN+HLpV2Frs+5wm/qw4lze7SKZYWNXmBvJkacI3j/W/sJFaCyGHysJy1VeUzpqo
SYZYOy0pX/1TWe4ixkbruYJcqcamAvvEtKfG7/myBmD9dBX4kpP3u88YO2iLNoi9VfNxpFVdIS4k
I9nP+HWQUz/VWaJaaZo6NoZo2/Ou8I8zDzGuOXI0Ii/AWSRcZkJ65havXc/oLIwLUrN4baNuDGf1
659yY9SiSRkh+/P0k5VrNkzyfapoXG/X4N+GmrXClUvN5BOsOnY3i5E+IAT6n7OElW+E5PX5dVo6
qygqBFjMSN1hbwIT4L4QD8KTi77OOxmRn8UWryhHgILNwB6BzHgQxXpGRgB++R3VCBD41DzKxMbt
Ly/j5A3SRn1XvzfbdSvE4kYPCG3+XGlgdvRgZRTookGabIRd6jN9p6FIJ8nGzG/vKJPxuXqpxvXV
+7RJwRdFKtq5Nwwla4L+UotHDP5yI770ArzOSY8vhXhy+QXHxfopv65JaPfWz2Gr6bqo/AvjTckV
EIy/3WwkFUfi1SiOSeCT07bLNYlAxvcuog8GwvQYW6p0Ofbr6IeWIvm+u/GXzX1q3FvAe5ibqX/M
Qd8O41FLAqXTBaxbYdoZRjynMu/eoeuMEKD9E77l8cD2M5XqsE/f7ossHvpCxYVbg3VvMtwpGdHb
/cRpFlBIpm4kn1ZFC+XnpBpo2Iufl8QtNnAjTzVRR1X6MzAJ1JIv66z6P4+enTMVCJt8i1n2lX1a
kipvOsQCqhekZ5SRCd+JRm8VTjF4j+5u9JtvgZNAiiFvwvBrPe39ShWPtTtE7wmCxmf64a2Lf6nB
Vausg39f5te87ngcEXsTjZyilGdr8WoLf3TWFnmJrcE5YDvD7nxPWCdtRJkeP/2mmvQU4d86Athr
oy3+3umq+jxZO+3fKZb2pU0ZNOvbjaPQA42UB5QwA7lD7X5Qb7j1uQubaXy2L8UgSAlARTUBY7tv
exsUTUH+AyYrEfOW3xl0ElbgjlaT2dYDe06ivgLbcFiCtEeu43JWqbwpY3s2f21U0M0I0m3vTxYC
lhtVEbR1o/Ighy4h18EH448X1ofC7CGUAggSVin/T5QNGUkaHyi8YK2DTHauN+YW4+kBdzZ78Ilv
p6Hx0lb2RYq5N7T9TyjY1B8cWjMue3Ob0R2KHCDTEpUfNK3amulE5DeTYQJnIdcm+Cj6Hnzqxa68
jxOVsUVsNLS7zy8ZOmoja9F2jH2ShHomq6KIn0NIUbKrLHEWR77eytRrWX6YT7OxGwHL7IlONj36
ENbYRU1tkyyT54IE4HWlhKGksimRu5IBmg5nr6cLh1ku7oy3c+lXha82ydKDumIqdr1Hct2NfJK4
yloIM0WS34vl70S3aYV8HcTj/2N2o8cviHoGB5GYFgRk6j9k9p6vSk2ITIV7rWi2/7xnhueCzWVt
+2jRxkWWjMV2YUtdqA7Xb/gM0c8vQTOvosJvnqFpity0BE8H3i1xXGlhFDClCdegChg6kM1HhLBC
J5HwFqRGaySm/i7fPwBw6fy/KSYIZvxrMp1uTAuV+oVMgzx/lGq+ejO0JEkF4BAJVzTCGdVu7scV
zaNIG5bXMECySV7dFGfkG6Tm1edlvTVu2OgqFtUDKrE5Rk8jsYoj4GB680q2LTh8YnnHioMzsaaC
d4kean0h1cdFhfRdY8cAy8algxvOC3/PP+fPQSCIX2pCiG3bRIaU0UZRzqjSrEcE8WxNMyKrcOIU
41Cq7iMduNmh0886cp3GHzNrtcoRcf/1zt8Zd8R9Uhn3Dc2CJlslpTRQIzDqZnmhE4ZzZKPT3nu6
xPWEfLH3IZQL0E0mSQmTnnUyKLz/gALWQnka7rbnWVStAfw4R5AnYBlQJvv1EWrHWsuZFQW7yfSv
vKcHD7JiID3xFE8sxoOgw00Cl7Q+ZQ3wTE/qiHc+I14ODDaMYAk8T8RsUPscFm/G4Yzmo2QuN2rM
ab5nogHtb2sdR0opzZnah7XbrbgZ+QqSwRyt6xlQFH0uddcRFLCdZHNgDKbV113Jxz4E1tLuMODi
oEfapgSEvhk33VxoDkSmBwts8Oqpt7l/fd3e2U2hLMVNHCxgcJfYH2ljRZNBWITyYrJlLGxixm2u
H4y7m0Dgtctd38MRX9O4a12bbYB81brJyvFC/kOiiy52QsWYYCnwTvpq3ZfC/d920IL/ju3z1EtH
uTqnXPtZPfQI+L1K8IC6zcmbswNoyIE5dGtOxO5temUVs5C9pgkEbbJEkF9L+Kfl8D99UgZ6hTVD
+gja0AY5mDP3J7ZFvqDS4M7UciR1TbsNeNGAlyd18jPkVzQBCWGKLHPydQU/sgRztui6kNu25gMz
bplfjU4GpuFjCiS+ShAejzCigVVCyuMwYDi928I2Gr328EJJHPKhneXR0OeSNOvHHY/0jPH6vw0o
kUXw47YU76RU0BtmESwHXreMfvfojcJoWthvaQ7ZETPMOLQPfG5LPMwFkZ1iHRjFUeqV6YShniOk
1NKrhZCOxLYol1azufXldoF+G/1NBmeSrSDdurCeYFNU33ZsvDsOJRKx3ZBXqTX0+tTtkQjGQ0gG
w9jFiR+SORL7HStckFVtw4pHQDFxXcgbpbSup6rrdLQvHJSxN9/HC+WgNdFHpw/Ts0HUalDmgaGc
/4GtSAFPtbF8MrOreyG4OJc7hj4KUrMG9TcmQfV1iR3yL6HYaMNWa0XQCKlD392fZus1lInp1XBD
7CbdWFWTDPwLS6WG7vmhKQwHEM3Aw0Goygl7ZtIxuifDXDleMBxr9QZiyrz5cmMhG0WfegOH1SD+
EAdVNISsz7g5RyTZ6LJWEd0oSdpwlbLavRzOHtJH0AIt5kv3GubAH+aYpmlErYSwws2+qqYy1KiF
h4sEbtTPDA16jtsEuqhvvhaZvjgnryFknlY9yDaeUgNMI4MBPLgh2cXFgtxKuvF2NZcom75Ott4W
8nKNpWqLfSyk2YQEIcJ1v0eZTEJYH0XWdtzIewRQZvGrFrFwiId4KHBuHmtaXzUr30CRpP4kl6SI
UVp4v5gmsPmawNFfLtp1CZxLkEoOG8Xf3qmPOTa1oxG+N8ImMP3SwbFiTN/cPK6dxctkjekQ3nvl
Tg3elgyXxtB/yOxLj7kf9Q54ewz5VHt8hB4dmPFxHCN7nHh1c2kVJuoTL2Z7nwJHN3Kv0YVZhVcU
0zlGk9ZWnhd7TWRQqAP1XvK+fQ1NdURlfrKxxmOnwWkOoAChiukcloOZOsT03EkHCH1lv1hv0/ut
FUsdzsI0ar2zzfWmltbiJOIYOhGARBXKz7OBxqRlxe8MspxdmWX3hxOugXkUItYTZKQhqgRK0RzZ
umqGBP0HYX+1iQy1CdWF9BI6uE/i566u6+NS1/BXYmwUSiC9KCLNUJCAKxeLEx5hnP5wEdOvLray
GrmjPv4SwnTfOoJY9rM/oIVu9ALSh9dDRcGYuCTCNyodboxLeA01VEru2wllesrnc2layyAXN1fG
Rj2jH15bIvykwx8krLVCgxFBB7sZOwlzAmMyxGMLOQosyF+CttYIcEOzGIddtVE/617x/VgM1Hh2
hUeH0jCjCxVgeQ0b7X7f7WAP2rXRJmEqbyN2famjYCW/Gd/O0P+y7vHo6MsrHFynoDwzPoVzhnid
Yn4kx6Rp4F9/ueIsfvrMhWO6cpczUn08x2QKUNAvcqj2JowiaPoOO27/JEuvLDLUrWnpovcUp++D
WlpsoSKpZor1Yw01myrhEN+h4IVnfsRiMOveySpcL/zs9q2KdV8LAkwhnUx7rszRdz7jHApID3Tv
UEgRDYrkWEnC2fSh7SFRgr9YdUbUbiCl6kRQKZOdcN57RQoFgeyMc7tN7adkLJ9mkHr/YfwKx7Mb
W6GOl84OxgXyepWKpN+92MR/uRfmU0T85t1QjnetoMgaOoyw+prJDajXM0E0Vr7E+5O+NE63+UYL
HTrpWptzTx7qehoZOZSDol+U1Ptsr52bwWBzYyXVtEZerqgiLEeKKGCs/oHrfZeCo1s5WAiQt8tP
GoVD0RDJSj/4wor5XP+iRsESIbAdwbRN72ysUREh2EkcS1QyfBr6+W4co7DuQbD3K2szGJBOnqim
i9O171DkuPH/VqhpmZuySt81oqZdrtlrSgAvNn25Yl+PYbDhSBPm5OtHu9/rm7MVAYyRIfdWcs5V
cIpH3RjSsQaEqCGNCDmaxZJUdGWzgtyccG5SiJ7IxvwVnuSnq8ihqFdgPLc3W0yOjUbW1g9YXZeO
5Gi5E4DhUfn7eg0WowC0CB+bo65EgMgzgSU4WQbAHrY59rFowQRO3v3LNCzgCtF/oa3kDOTlMhLS
rJLGWHSYGrYh0A77tqGJe5md1dl+74flAdlC9NTFxl68yoEFCCxDxjS2Iu/jCfPZWWyTUL+dkSfU
YSCPcfHVzqwa4ksuJ1wgcUsj07pW9p+AYTyXGiTvqwAeN8FJdsK5NYXuaFHsgjiDnQg74bsxla9t
S1WtWXGw90SvbZ0BufUZXXvXISHgpY50TwBG3i6cnNjpMHJJirZEUuJ5W0cXuxiOH+8GIK7NYpjz
DwrD5rAsszIoJzIO4DnPFObwmtuZ614bEcBw6Y316hsdAYFCcCgxuCWj96PmwWzuFzHva/zfuo1a
8fz+TAdb+HOWre9PidSnVHdRFC2kX2KqB69fAm5tGtPPf5N5mwxCSsXfhYLaTixAIEUVs7ZSSPfV
Q19JTUE5XcZ55PXQgtVY+DffYKlyO8gcEPNdiareg1Az6+MrhiAOFYT1D1s1ax11yAu3WKl3Yna/
r+7pgYlsmjD4/4MiRR2/FLp4QfLydivqbWpncYuQ66pRMxl/ghTxF6NQ/5Nu3EPeVtxl0uAYeW3p
XX65mBeuS8EJQYdsP5jobJG59Smz+aopjJr1cXL5OmLqepi9F81NP6juSaJDO6B1+mK2iGVRDJ1O
23tgmyUm/R5GbMsG4k47cfzmkorfoG8qOQcwNDzY1gNJj20etjEek3X902taEvDlpuJYxuwOFGzb
8dZ3O5mfW/fgIFPk9bol68TrSHfBN5HJq47lUdHsIWqIykj/O4BliAcVR8RiFFD2GldhACqgaBTU
QD9h0vSg0xGsys1nQRfH0GtQNqzE+WbR9PKa5soQfcwRrN8HKhMgjmM1RENTxwAbeBd4j/y+kYqI
01iTv2ngsRJUaOJvquIDsSWWnJMmRlGL/evPqPoEZoG8TYwYECA5lV8ZAQoZtBYPTpS8XhWL1a/l
kKGT4nsnuiPt53dd+D/+euoRqlhzsg6VqdD3RlIh6+n0pkjB1wRWjTSLQVPn/pHvkHMHpX8GZEvE
nrl2mM84GCQE/SmQcaLNwNwW2XGrgvViDcT44ihmf55EwKMlRRPvvWTf0nL5EjiV995kXG+Ve0wA
U+02xTlKkj0geVfiEW4KzceGwasR65kilOqLXFZp0TisV5BCjOlW2ZXyaIeLH+WZhSo4T9OELC3V
IjQ/1DmNGv4VCqz8kOO2MmoZBslZXI11aN3+QVkwHJ31TydUFFIGtLEt3NDxX6Cpf5r/DpzVCYX/
mleSpAvUrAdmHE+xgOyPttEJ8lvHfWVWR6Q6N/3W4rOymh/ymMUFHApJDw80hDbrfeDIz39TIP8B
3np6lNRT0rTHPxHl6xYHYvr5yUmTr82pGf8uvCdKC8pgf2XJsDsteWHYyyALvfQHPExYzOQHhaTW
s6dcmGRF2jghm2nAObtM7Rl83ut2O2MuDae90o3PTqWHUo8q6uGE2GoV9SXJNJvI903vpEolV4IG
YUYbT4f9XEXtTmv0kp0qLwQ8q65uQTHBbExJOHJxvDo9GzzW6LjITkiXUq9/GzVdlzy8o6KWPG+M
Pp4Si+7/qCyqDsNVjBbXPlihqRKHiiQqZhdq7A3NshsIyB+QNgx+B9QjhLy0wu4YKr60JxiHh7st
LV0DLGYd4z4/FYmoyDbbC7vE7H9dJIi74JZ0gYEmI72jKQTlAMd4RIi2wlZt2d/QYSiXwQKbiGx/
yOfGU90TzluYHhaj+MwXwsi0lYUUOBjFkARBfPWyQY16749UIjfzr/glg8qt7zy9fvzZle2idruc
pTqJ7wbxUtfn+xvNtVfP2+yY0xbpUk1CC/jOPBIvnUhGw2mDuVSJSBlC3Uh5IN54HEWMuYYtn+Ug
SAJckDIk2SCFwK28fq+phE/wVItDGnQ0uZQuteBrhKwsRre0L6cbdkeOBPsfEVb0Mx86UDUJ90Re
DcpA6NxGQoKJyHcaJIMELkkGe8YzqXDZV0SYa2xP8R0kO/1TxigmvTermkqAL4U0nssBKoZp35Rd
PRgxZyBo/duGiLcKqZGmled7aEmY65tLeS3DWUTwc2HLTByT5+K/VP3UCF8zQqbtTHcSvc8Hi9UT
Kuzr+vqAaW2hQcZ5+i/HNRmYzvXJY2P1wCIL8jP03/b7UrijHiTndxFeFPxjQaHhtttxmEjct0DL
GQ0rhjL372UJiawyDZhlDq6yoz3CRAxt+5KBKWKu/YDvFgkiVS6w71CcSHbOJr0E4mr63TMHt7Ug
10sPJioIgL9vF5zjKzo+Mtx1lbpGnzQRiK4PmbP4dSeueH03GSaIICxbSZBTPvDJwUtvzpCrEmkP
hC91ktg4it5uiKNxmX85xNcvLaqPdwvJcoVS/hTdJMNo6A6WXWsDyim2KadhOvRX+WakhRC8BRrz
aHLravoDRhzZpXqDgg2MZqNEsjcJaBHYF2/U14QX5Vg+CpfDcYJC9r/ifXkET8kK5VMU+P+0dhhb
aHY9lHENrqjGqSOkKgvlGeJ54aSNFhpK0V8XXnhfLjK/Hmg7rwvAmqhSsfFBnL1Xm8n7BRhVhGVG
HdMxWiW8Y/3n63lFfPNLIay59CrVUXAD+2bB+MjXzRVlDQYEFQdTKYl6uljFlfD/8kLfy6E9sONT
+fjNaBc5xnDi2A5mek7hzrHq/grqlF5T0Xs0GV7DpLcWBH4xd4uyYiY6bJDGrcmo2Twy3LN5Yi8C
3jy5rz1hKFPjLAlDrR2erEtGj2IvDL4zYJdizYEEru4EXrszxQLd6ccNiv/q8UZBay/28qjn/UAk
/S+MF9X+091lTkpXah1aX+AxO4amFsBzZsKkgFMOVBx390SePCsLyDzE0qGaHTqkrUVUozblmTHK
sn25KqppWVLVpwdAidGtQWSP1WbjM9FmNTU9NjKNPaxwWStID9LibNIgXLP2Ltw/CqUx9t8Ceenc
8qmclxmJBZOZu7YP+LG0ZPJKhOSYDlEsCWoqMmPfFIdi1ZGi2wV0BJh2opfi9P+zVkCfUGUcJgyk
hEL5T8EU0MnSnGGZLD8Ko/5JYeSwdT+PVdoEPBuUsX3D3rbs/ux9nt2hQTuZZIMr8uN3k86JHHu2
7B1CgKZBPKMKvL/bN1g5Tus24zSL0tRm+efycJO0ekX0ggH5mkOoqAxwCu8Rc8ZRLSdueaLpQs1P
DZI9MmK8YMcTpTcnN5FZLSqWPlqy8Y1klsF1RbD+6CTF2d+u9ZodVI2T1y10kmBYld/tN91hw7hi
b3mZ85FWPXiQN6B22zvyw46hmScVB9KrTT53RbowsaFjaqbLSaUDh+B8GModo+HFQRVu8W9q+VV3
yRE1kGKRV4PMZlZA3K8syMUcmdk4iYAp1QbsMCJgRpRnOMTt5KssQlRDsSWSguI+SCGtQubEOUqA
gYC5rExf7+4n3+s8ydqbNMdmSTF1X8I2ag29MnuKfCV0fHiwR/NFLji/vnN5exat8oZLvxBmcIOj
5meP0CovPn74eXacyAhknZyLZUOU6OL/4lPF279aN1d7kgSXTgTJd2YB8sVVxV/t+3dMpxUmU7jB
eELquvKSY3z1wXWhpMun9up10PpXXmXpIad6QoKiRYd4A/2xVmcm6cSRrjedCp/sQFNiojoqthTk
YzpM31FtlZEJjyqvPoQWeuEE5dlRIZbPrspIdZXCcujQY7klsIwPhU6bYAa8rN+WyWIWFAwc+Iac
pZW7Q+ent+Equc/vIa8T0aL2Wc6D6RTngl4nU0I3sl2n839PRWI93pQHA80Jkk84/p48ccfZ3Z4Y
cztif1QH9H0HDIsgCewgG6LBGSEF6aSTQAiddOOuXEB0YBTL4BgyjOC6NGVULbcXJ5xrhn6joDge
jIMBaNBh6JZ+3EYH83H25ouuMnfcm301EEv45TIzAQ9FcMxnT55Be7YSgKGpOcq1Xm+AINoHZu1B
BLNxwW3S8aRKXCJgJIxd/seHWP54kV1wVlHq0wu83DuLFrQ0/OJzx7s1SgQxotMOOb5Al7La/2z1
q/ftPAkLiL0jxA8e6J0tduKa9q+H3Zw2ia3LoCjOvO1mqnJ4JyJD3Z+ucVMBqqB9aEiaaNMNRVKo
//MOfuwKyJnuJt7mELju8npK4XHy6PR+/7icxnEyn3E5pYw66Ul7Qo7KUUo+t+ost9HCMjoB5PR7
D1dDS8xoBhu4xlJV2j5QjKyORIHgzDuRe4uYl8tgl/Ekh7oAHzpjwFk7A4Di5DT2gmYF7QJnRJFD
2TSxKWLX/1a9UHLqzdaGssB5awBUfdWPcwTDgOYj91QGukZdgWNvh3k1JM2IpvLz7dIu8TrdSSt2
V+L0/cOuw7OtHO6C1fybdLjTA8Gf7JHqVBRkA3soq7NjDB5l+Anw+13WjWqhMXOmLwteSxrrec1d
r31ewV/nulnw9X5yKe0GFSEFl1tg0AWjfMCbinY8Qv9O50wumFqu3ZGwJAhfqKkjvSLOs7UNxT8H
PkleRf+XzvLkMmmkVxHeF5IkyajogZblxxEcjXA1kQhA158AWi9LTEANnZ/vng4jewjgGCP/0nDB
dUnvBU03aN09PGyPYGuc6hNirl92jV2BY1HC4CY671ZEXufp/ehYf/Xi40FYd+6NZOeWlRXjktk7
CrTja3LiHjYFN2IrWmMWIextQcxjw8pyNtLD6zHNxlHrRgp5Z0Lk+GAR/cv1+N1d/oFzKVRFPWHf
wY5c44OuRbIiC/xQ1DEbEdfE1qqomZ1jIRX21D7idOW1y4mUy/hJlUVsYnz33bNP1fj/Zn+JmnxL
S0nJBKdqF5ofxx/QorAv/jje2/mKMPBem+6WIAupciIvwTz90XKwS1BERleqsMWcmPYJ5Po2hubp
COkfY7HqdsMSiKAYmgk1mBJqHHo7XTy+ohQT5K7IadeHY0r3HmsJf9BAh2b/LBCgl+1uqcCX6P6l
z6UAseaFsPSINSOGgd+pUly8U3dkGybE53jYASoIjoOjWm67puOVEfCxqaXIGezPkLk03bYtQAaV
y5jrdmKgfP7r/Hw4RjalZzgVRKhIK8oQtwyF6kT8V48x04xchE04pwS2qz78R5tq6VeU2LkkR2vj
sEBnUMCO+YoqXpGJgK3xa7ZlVeWvqDCocamRYd9vT4HUDWt3Vxk0hQpkgAIcCFOrPitdq2/rInVt
E+hQOJGG4C55q5PJMUv36rBYexaL4LQNq1HpR5b2fV7RZtyYD0Asqqx92isqu1r9Mqpr4swYwMOX
P1NNf4KWmupwAJJYcBVh6OVSDSdIjiXMQgZ9VUFZWebwjKQXiSDVc6lOr1xPlGFoS3LgM9bZdpx3
l+gss6Djm6u5Dxt+9UuFvuPgvKOg5ZcAK8+elzXO3mDkABT7MHFCYFg4AsK2YY5qvxiltQcc1sWU
X4t8eRNdMkh3ch/1eVYXdF/dgdoCjoAr8FANGHBUwe9Hi6UVJGVnJgCUFkAiOPRVMNesH2xt3/Qe
Q9oKyqS4JCAOUT4A4EneXQ/5wjIk/OqX29BImMVi0QUan2GBBPCXSC9DC6kU7RmLqEa7cx5QWUFQ
7fuETns46qn/2QplFbhEmOSKZdwHzzobkBPaRcSDO0BU5RcFoO4un+DtJxDXRsKWkx5qyHOX0kA8
Y1a0R7T2O3o6yUcwzE12WeoYxcYoDuU13mPcm4vGYIXWX7QVWvPKTXG0DzjzLzsSBUO+9Hamppbk
KHz63b/xUAn0utsq+smcd/pkH/DgMjO4pmQoVAflcCIgw3MM71f7r6/LG+7DbDFy5bc736+WFPDA
nkFImtoFANnDa5aNNj4x7WsmdGYqEYHuritJ3n45YBD0hAoHk0qcsDuEq6EwJAwiu+dpIjTVnD2l
KK5FDlnSK1lfjnzhEB0H5unS0B/gCwNg3fDv7twoFQbLvjxzktVqkBXBP7FCMShHkD9j9JBJPARA
GvaLfwmu1YSR9y8wgxf8MFWfIs18WlZMXk4SR4yYZfWKI6vy+5V330oQnf/XJqYSr25LILTE+ppI
QOXJDs159J/iPKm1Pg801N91pf30hLYqfFXkfQ952xA2cEQ6zNCdEQwmonuiVoBed9/ejAABWS75
vxgYfSlNQFeT5d1nLL+eOY5b9aoaqg55+L1Yc+7KIoC4zLDgvOTvr9iSbCiGRLVmb+wcXdBWdzeK
OhLSge291ZkmeF0xVNnOFNGtfz5/77Gg2l/eQBu8RhxMojUzbs+15watQONLyF1rua6v4UAv1gRR
vUHNVkC51CtJhUatzrQ2nd74MzffRKwt5WWUmiM3bJQre0YlF947H9qNLGex6NInqQpaX57AD0VP
5Zf5rEqDs98aHqFArovuI/umPzR0qCMzrFAR8YpMzHTP78l8+8+JXgw9Lr5lg2auHwnxyNT99r4r
nAll8kOPpesu/emQYZuYV41wvmAg8RuFrZ0zk4IXH2ZeSEfFp8Ukm9kXo/15Aqh+YAowl6wdV7Eb
LpT53Zz3WnRdfaKDBDRcA4a0QER9gokdoyD/XcLauDa1QwbfqTvf/vzFA8EijDEiYO8Cj5B/joyE
S6wfOkx8hA6vRGb9Ge/WBKZykAGkrYjAr2lcYOHqBS4xYEqQjmSo8IXqADVO+Y8QyLss55KAA1Zy
xtWOw0Lx7CMOgFr2k2bJ4OksH41f06AAJz1m26lYEb98IbgaLpNcTajahg+o1pYb1+GsfbPWadmE
dxrRtlj86lhUdSuybZhqpll3akQVKr+aHTjJGiXH6i1V4Oz0iUJhOEO7hEbwVwolbuwMyXoliLWm
BDgvvVEklxjRl2JfNc/NHCYxC0c8YUmb3Ded0h/2/CujwWetZDw3Gq1wk6oaVJc7wryITUv5nCxs
1ec/N83ynOAWBMoi2qyTns2O9F4dtO99QWqqPe+oHSV8cFLT+/D8vEsRNmhSaImb53eyQ+0aO2Id
JpqPadOWuQVk65ER+tt4G150r/Ma0fjNLBM5JOruylwLWUsu0L6hizUPbzkDB5TEndFHR8VqZxEp
Cn+mVArTO0oCHlhjbWev/R2zNCH7oDUJOvenfZHDE7CRR4dHYoc6xl5CLrpeRs+r08bkHDTNdus1
cRwTUTd1jnjePlWG6KLQOfgaTs/+v+tOLB5FBw7zLsOexU+Otlgm/L6h9vrGmEeLblQysba+11S0
EXx5EKRdjtLMc6wskwgHHIoxxvs3BUCuyeyHmggIsgQpBHdMGlzAd7+zqKC4U5A5x5sYvlahwYBP
aa/QP6Cn+rB3+pmmo0avZHvZWh7Eu6Qo1SD1Qw7Xbt9jPNk6Ei+XBK9IIVt38G8ssYSy6ACQFFGG
TZZNnFcxSrBKVPyR85D9GGWwBOqLPH+hq/r3OGK8jr2kn420Jc3JXhuT8fZPWVogDu+6XQ2rWdXy
sZyE3Vy7qotkTs0MdcR6zYNCwqGaky8Y2DsObcKEVrDZ510Djkwr4W23GMRg9ae/0dX4WzTUctup
D1xNcCoxc25cD20/wHD1gqq/7Q0Hs5gHOCxiQ+dG9TIsfcSxyMuqrulvmutViSd3upUAfZfoYTTy
hsZeI2eov15i2ZIc4xOGhSsF4SXTS1wxV/SmSXnp46IFrG0n0RIEe4zst5evwiMGmcCATLk8R4R4
F/8k9cBuHQ+HJDPg/wpQ+0l3JVAaF0OGIgRbDq1m0JqTiua7n0rBZ6dpwfwVPTAI+1qZlBqLA/EW
m8Dza6GbU/9ZNXNm4AnyNPbCjYhMt6F+zUbbiYqLcXsLvkZOxuaffCBmtHMm5Zo21axw3hVMBQe1
qNMcchgEy8A6RXmVmACaWDNEfKEtrpDLbRvIGIkDhixBHPNvnoF8pkkhcDBZTc5e9KCWSuQlLCtN
l60Gbmw4PbVK97km0QpOd6Y1Ohd3T7RJxm9nTQPocsy+b3U126gV52TIb6LZYUOkpt3GcNXpL6E1
02DBDgNerMdK+rUNkLuvE7j+IErRRUNjblw6alObYklhlF6WfcaHhiThE91zSujAqR2VbHv8s5eG
H129zMZB8MWM0sfmtLtLXF6d81jkPPLHJLrqOtMoVm/e8AbS5zj7NgIK9o0dy9DK1xrGkB3OGD32
5N3V3kWTy3KaAvsCrsyI1DLkFik3jJYogusARLyyfIh8blhxto3YRpIXhuupYV4oMmGmXMH7cfnd
wCmL+sL7ZhUtI6Hsr3mjprq7Yz6/SuP4RRn/Syh+IoYw0z3szyAqRlikaXEF+Fqf3+VOBeQL6TRL
uU0CnCbtCBKLd+4hj3jlVb49aMI1di1KR+s0XgfEXd/L8zsSTWtfuKX5rvJgSPo7dkhSn2rCHx4M
q+TPLmE1DNldsM9bD5tVutRAKbTB3pv8fquD46BZF4Aqcotl5Qidegm4QR6VMv7c99jLUX/Abh4E
sfzvL2vBmqXoQ2v2tYTJ9kk7Bn0tFxeG583KmS/+6G/6VFfGFknk4Ma7fcM77Xgkbw3PQBcZPpAj
fXZhDN6WzuCVg/NsU2xAKB8exRoWVM02Ss83LAlaY4eJtMtkB3MonpBY0KUBHgeyckuh4dDWDi9F
IvkrstiQmQ8RSsS1o7MBzZB3fapKToMMEZeXMzcgQoxtIq2cHdO1i+U6SKrM6J6q3qb8uh6MIU0i
kNDCaVA3nJw5aw24DUyKnpwdPfuNBXUFKrLzM5JvX/2m2BgeXd6Ov63cvxTTgLu28uHKOHsJ7xK7
Dizf6Pk0ZiGiTqWhjHxEjgZ1L5FjNAUL7NEx0j8s06LAsjTpSi+35cvcYFTW5uIaXSKvs7UJzXGj
AhvVmGocLcuIEpTbBJ5krdgVUD9Fi6AGV52ZZS9I1B7LDJQIz5kLvYKS2x6njeDif/wdzn/Cu5nP
HY+zRL4w54unaODeCWB9aiIn+O9bUf45TIUq7TVtAJUMOYjEB0JCoOc5BunWkxpE8WI5whbZ0gsY
lzlospZjqKqGhwCjAUHDWus3hv3CGIRMw9nx8TRHoZO/CythAgOhfLFxj+0EWjSbJj4i1l7l/UsZ
eD+CRGd4QfR0Wuou4fZZubll8+T/rZaLUktUXNTnr00NjWS8Crju3FsSWVUzm0pF+E/mLvWFdOQd
R02mRfRuALHNopIoHGj/V9Kr9Q+1xBmaGF4VZkg3m0pNOWZA9f4fme8hnxHdc2Q712ESTNjI6jBY
8xZ7M95+lqSSb9OaAF5VjLlQOUblavTINZyn9+Bsau/DKsVGTn4MLe9t0yiNQ9n0psObafLBZmJV
IbB7tfecMd6LZtSsQQMJVkix8XCEkNk6VvfAhUvzsVcxTKk+OYR7/CFbV41a8YJzflzfyh5deeiY
xxecsFISeTtjstBSP+cajHk6fMNr8AHbmrax1/0fb5KYK57g3a/JTFINZ79rJKLGNNqPmvgtobeM
Gpcsuo3iYeJ9eE3cGRaksb80Qg7LgAfCbT9HM+yEGGMi7t7S0jMEWyEp3x20vyTzv56z6ETaW9oo
PyzczXnmUmWsGcD8KnSRZAQEYFjGVvC9/bEBFe7srIf7ZdX0SdG7++d65oVny0rrmpky6DrLVRMs
qc4lHlda6pIhnBBqY8FZ/nwOUwp/UzSmJOuLHEYGgg2ue3971ptkkHwQTz+IC82tpRjkOast1yev
zszlU9YeZrvjBhd2KfHaSMrnAd/ef2FM3NV0tthV3NgMduAN4v+9Kyof9k5DhwI77wI1F16/yThT
0AyiWoIkVt2kokjlrcOcWUKPw/v7bXdpuvJxLRyyjWkm4JuLtQVZT9Z5zoT+/Jdut63TYovHQNTr
lG8cT/iTK81n+JBcufMs5WCryh3T8+7xqOY/E0MxlFHaLwtQsP4mMttpXaT04G1mQTxkCsChqfsQ
BCKshv6uMoINlXAZKHQVjpbuALLDT+hC+k/Xyy6N+bA4rUxMSyiIiNn0MDRDWH3lJt4htVXL2xV9
+t3y772KBJ558ngrAt9O9FCuzRUkoCibNc9wk6Cq6oDfObf9TQAVvX5UR/FTbzaA38HhXvJc0bd1
2f2IbNqRQMyWf+U6O9Aaz3ju01G8Ocnwr8xiW8VVOA9v08s7hl6nKKLP+z6xZ+ko291BHpW6nOJA
TEpC1bIp0lxn/jDy5X5giIOL0xqUalGNWN9NvObR8tS71U+z4ClmDe3SK8NP7DOkoP6bQZItzN04
IsaH+34MNSoYbC2ixCglrlQGreSMoJ7iBWj+kKbQw3kB08mJn3XnnOCtg0PcdsARLgrldr1HOJ3E
tPbLdZwx0MDfW8HzWd9N9pLTDkxT6mQaJw2DUvj3pgU7I0mFWEtKLQU8D8XGsbW90Hp9fvQF2fLa
fgwVdu1mH86OYB7eR+IG5vE8kbKbOWKnKXIiBNuWE1vjDy49Di4OyY16+UTo/rWTzzp6eWrHf3re
8TiubhdXSCgzD1xzmB5U0qbpkRA9WMau/AGueEUYRXqp27q0OAWUXB5ih53fcKuvw+OoH2tw9Re3
FIFSopfoCyH2la3F7FqKNhziffQTF9OypIKfpDYageBk+DBdlDMJkTcDs1Wjk961gKTCclTCOZ9r
c3FWULDWpEN8NAs+O9z2CE8e8+wfq50OnACY96/UaR5Ax6b1zSkcOrkdzxmhltK3Z2X0znW2khhy
0YTaZu+fFt1JOHLm6tdFAhjvGY+9nGGVGDvIG4dbYERIPyvZsoQMCyzjjL23UpRIZz8MNg2M+55E
aP4vu5WqCSO6e7QLsvVWC8L7CBQVWd+quo0QIkLMZwUWxPwJ/jANvbCtkw7PEUT3dAN8fIMqA+Cq
6wCHhzoypVbKRzfWUTx7vfOsv1BFz+kzq6z6jU9HXypzfYX5O9qEOzAIDucfREZ78WUjbgfsX5pY
23tdrFJzkjluOqsrdSrhuTJUAFyEo7Ys/6QPkNj80bjyT/jYQPKVSwxAQmeZzGAHdup8M3zUO/6y
IL5HuW74L0SfBFG5QMQ/isNbHAnNBiL4psdqwdCljzJVJ5AvxEF8rmrjvE60wpiLhus9K4Ohze/C
Di/4WpSfx6WDUJY1sAVoqhMkR+tR92dRkkJSnheadHCNCoJVbIJHuuwqI0qGbFCcj9WsuGWWqyWF
EFvfX+MxJedcqmxQezb+3EfoPD0UjButABwc/NUAooH79JyPIeWQG4XvMj8JP3WMOQfFdq7EJZpJ
KyHfPtqzGrJRbINVaq5WFwqS3+n/Ly56UYVjKqcKP3WAm6SfOQlOmoQOk1eO5plDxi7niifBCxvI
1IDHaCEYESavIUePD2ogy1abT2oVyU2r4D6DjpeOX+LBj9VvunaT9xwxI/PBIFdo84tBn7HwKFKZ
UIHEHysDQ5m/D8QSWB0qfE9E9Qs/QkVDoQFikg8iDM5rhRgeSwixswWa7pWKnFyvksPaqSciCSMx
6ZsK/TS4/bvArQ6mBJRbWFWf8LuNPZ0BD8WtVU4VwTO3+jOa3Pn9d4zP8q2LbMiwy5yShy4yLmBR
QcmoS12aodevTYW5/tBNcLAPhkw8+tEUHEm6EAuGBy3CZQpzxSeXYtjdtMtoPO6U/GHInyFoTWrT
DzQFKWjveWmfwQBvywzlDFIJvva/OlDzYWuoR8Ms7NjpjrqSOfrRxf6TugbUCMJ025Ym+shpVel5
IeRIdL85QIRspcZYso69J0aL/NjGJXsx8OIOg+ThVU/9QfXF+7a1HQT2EvA1MA73QGeaatJHMYc+
kEhIcO/KfErDUpLQzf2Sgv7QgRZXDTa3BHbQUT4Gx314RqIoVSnOhDgxrGjUqpPq8zAnePiE4de1
IRynDbNHWFQUqJ74QItVkLxcyGhhqdbbygAN0X7atOpqkrLnR1jrt4WUAFtf2he3NIBCyGIHge9q
xOknbVkEc49LFYW3GgIit9eWhAwQTu8HYZBbFOhtnPfEuZPf1CsvjpbRx8bJU2yi9h5IlJA0bM25
UB7RjhNQI6dJ/ChF7VmQFajhXKKneeM2LB2otAdFuLuuATeiC9n7xVAoc+90GTtbJQFUi90siUZJ
fB4+bR2Wet3OBy9gyxrMvOEAmEY36kjuA/pWGKQCV882g3viCdHFxzWp04NuxekJNuFWqJwm9juT
Dwwddo6N8zIzh19SlVi7l4aG4VcG6GY3QEAEsxhNHU/no83M983KS+ypmJdSkPOVrgojBBOJa/44
EXbAWUF1Z7PWdr8xdbiNCrO34FDc8OtoG0IByoRT2ZPe0Bfszh0e4uKGo3csOu1ff5hxqeUMCZqR
5lSU687X+RhE6bvk9vB0NkTci2+D8xBZGiS5LXXfraIyeX94ob4vJYwtnY11On+wJ7xejFNMy+Gr
frC4DY4FmpvkFvKt8+khaQvDR/3dH+aHgg6z4A0OesmS25jp/qxbUU1Pcdn9goPKs5FBiCxuHvg/
6LtnlBH0lnRur8HKuz63z27wIie+xmjSK8UYSMS08qFsIVgu81HrSyQXeM0UcH/33WewWMJOvkKG
qFsK9t9pMJRa5m6937y4imAKd8g8CWNvN63IQZwfFhYedakdzWHpzX6BDMvqSGdXOwYLb1eTWUyU
t3j6ATED/0ziEba09RJJP20LzSnntNd0fQeL6r3F/5y5rpE58WRJ8dqoP3z9soqiUFp7w5qlHVYY
i15mMG/o36svXM0A3xTt5Sg5/291k83k3Ruooewnu5HnTPLBLu8cMooOfWLK/f84itnt7mnMhGvL
IiBzgcmy/Aco2zYzrL5QhDBDGKo9iSU/+R9agLndBaWErwwPkzVLGgY0PtTLh3r5eb6l5YfPkvxL
Q2x8yhP8Q2j03tW31TC/X7AERrvIlpev3ovUNkdVjj9TBqa9n1BxAIFAmtjkucvwAit5c8B6mkZF
KNKTMY9Mr8E86EBmmXAGeZPNP6lfk/8jASgtFGIPij68T4twCaEasQnhQOcNNy/2q0QzXONld6/7
GwKhKkkTNuMxuUGKj4aS66EmhZ/vlWXt6T9gclszxoFpv6yJaMgpoNreZLQX0BVhLK6sgzIV9EOC
XXoGv0teWXaOs1nuwPARhNuV4Zv/Ein5udh1PydX7JUnCY3EvHAws/mfixFvOJnUZ6Pwdp8hIe9n
C4S8eHrRfpxN0SBOMjFcb/G3H9oFjcCDeEFDDgtw+qE6F7IDBXsev9ShOryA8fqOLmge9ovScus4
zVC8GSuhtm0vKXKh+2cImJMLgVeBXq01lcA/qk/zIHBA6W7gJbpA0VcAZg4F60qtNajAq2MOC/y2
R7iOWM8lkRiZhNsE9vWeDOFFuwGoUM77ChBRnO+f97MtGDPdHp8Q30xlPqc7LzgkJFDGgcWXvreL
LHWEpMlcXoL59jAwxKXEZjwmRZPr9yeM8CoLpMhnR8gYsfSDyv0I7T9PFRjEExeoqW8Hbd/EdCrF
9bf4LO6AHs4VjTcZLvtCYdb8B0ze2qf6t9wl7/R2BUmFLjfegmZBgeFs6k4eWep+tLs+PhmAkRRT
RzcngjpByVt383jwKaLgiR5yW1zLRLZy7pVMMsDscGeP0e9erx+PLXOyI9Y0t6tgOsJY6QI10Rwh
H0RImU14dHJ9xQ7eMKq7kMkODfzDWAfGksoZfR4x3NFb5LK21K1J15Xyo7JLbnbjnIbguUhvHHJQ
gxwsnr0Amc8hgss3swihKLsW429bgtmqfmHAq59Wm+PMYFasP0WXNBHAfmLTm9inOjLF8qSJhMVC
o2orhHoZk9aX/Y9Y55Gn1YLu8IlX1uQo6BPAvYePPhV4qQtyvXwIUoUIHH0P/BZH6t5ST9I1zsZ/
0AOcahuu90jYRw8JKTNxCfAS2Ha+cngVJK4+yxDGTLOEfYbPh1VQWPdbBX5p4US7bvuavDiuMduv
8c7rOnqmCMR5FBB5ylEo10WZQV8OWBJvBNNhSEUiDaSdcZiKZvZZl3jE1Mxyz9DzOePD6qJ8S3JG
nMqTqc0SDY6rzB2O38km40OJddyc7IQwmzBcf+I43mVwkC6OYvOx9iczGZtoZsRVsrbXr23Y4tjX
KnAN9QXViunFzrzzywdcyrw/mW0Px553YTHcNGEJEloSGiAcBYox6Rjjsj65N7WbqEsrVOIWzxuq
0e/X/RtZzy11Yu2tp12i9VWkoEPufT7laiqpZ2GyGpBJ7bqpTYSHwvsCbvWWWnSRiMtWX+eH7q+d
VLsYDyXteUQJ4Ykaj5GnRSO/Z5VCx3xBDeDe1Q1ncZSGhwGqPM7LDOaubbATxYXvykjZCHJAKdFE
NMb2A0wErpsZGJn6A4WENNqLsd6EtB4hTGtZV6gLF1zjol7QF0sUXU3X9DDdIa9U1p/tz0Nfk6Ny
tT58vCxz9br1RYm2Fagq9Sy91+kARcwUDa3z1ASEZUdLknLKq6C/WHSxdf0aT7phXPIss5Es3wKp
qtKQwLhMXzfBJ/iuA8WKWVsHBDa1Ih9zQjibo2vTfOzvmZj6YusYoUlcfiditK2SuhmP8ziRsqky
WbQit79PL/Ufn9mdii0DkyKdJqpy3tMbgFHdmej+vvl03Fe3N6IPCjVS7dmwMYvy3VzELkE9MXC0
kefTGFi8x6adZLs+X8852srOJaygUGKdxH95KBN5uIqLo0scOyVoYO2vOm1yhG0t6kQlGQELsG5j
6EV0beToSr0rAuyTUY48S+jWo/vcxYOU5Drv2tU39h3Fqzl26PVV3zVM1h6prcdGIgIrvFRrn5FY
B7umH79ZMmqYb3zzABY4t5WG4K/YWH2U7BzwCfFszw64YM4g4r9ra/3UBql6ypEyo6A9SESloJ6Q
+awVRsyhMpNAKhIy7+Wo/I1CgoptqTMB2SsGeKRymjyMfAywI8YLKlJx5O0PmNajL8QB4vhWYlVR
cKMCuu1X/uuYYy1cK9BD+QHQgaZtztUALkbCaXbCIUtNUsU5rhAgT1OXxy/e16Ja9MZa3Ave2Kaz
VfP/dTbOhA6GVLTZbKRYW6c/s8LB8VxMCNT7nClzLvlwkA+ljTL8GIZ573BoClG/m2yP+jlKPc+u
BayuHEliv7XpmJ+yB1JcuhcyjS1kyYxhdWLYGq+TgluJl4TmCBcbtmmjtMcP7UR9xtZHgjmHVxaP
4WMMUGwl90YNzK5PE3q6d1/nWgF5UX6BNrLwasgFhDkG3dJ3Lwz+048EtmMcr0rlHo3OLVLq00Th
tlhN+it5/lgwH/gkKPqdqUAt4OnlmP6FddFP8aho/v3lkgbuQFz/vHkygnvTmQqyBV4Eu5rDpcn3
yzE9e3ZNeWxr7ITx+NFnEXzC6MDA15/qa2DIebTRKdToR/j/yo0JYMHy/r0FJkRIxXCc1/XY0nDA
opzqMUhKNRrIIxFLxp0Sifo2vBRTahU3EUIQx9NlzLhzy+e4F7QrWQhN5Le9Hicy8wZiqmMrckG+
4IxR7EnM8DtXn/0uTsh4+NF54AHwmQ7x0os260I0+jo1UZ02YUNgI5PqI2qCdO2Xt7uTE1naO6fl
aRcDYdAw4RYQXqUc4SUTtfZ4DxJlpAXJ4D7+9QhEChniD4zlT8G27Fq7ULkoWUOH9SZqfSPhSpld
VVSpDNqbStFhrGdYsznAXWQ+F1pmpv0hrs/UhEN3GkGGlz7wP5S7waSSvia3ezpXmhmNZs2dsTR5
mnRhZh1u4mAmp2jZJLNLctIxS9cD/xQNYzsT33DQdouVAMzUlUrSADN2gQW8SSQO7nnurG8yKPgZ
NJcGxU5jbQfkXL8v6DhCQh6V0QdxiXMNoStCPLhYW78g/ljfMoMxVwTCaz68naLIF6a/2tUf/B8P
Op9HdfTw2o17bkBnsv3XUcmT2WiDjpAkidWLRrOFittJThOhFU66/tz/rbeLp7Kav49yR0Wt5YKS
FqVd0OllLfbpnPt4Dux/y3SRBYkYwNp8InzMH1puD0t1WriGPWKc6AWy0htS77oR12wDmt5f+UWo
ujQAGVwdcINa0/I53e3DADipSbdtDOnQHN5p+XrW/Ah9aR1vXwUncIiM46QxrM7nZlXtIF8b1YyP
nlFVjKWDdmJ2lXgftM1faeTExIVE09wcyMwN5Y8m9ltAql9Kyu5SLEcnwG1IUzq47R1t7TmTQCru
2QKeqeOTROafbEi4AT4m+CutgwsjSIvGMOC4yILMwWxHY9vfg3csuJxYXzB//6/NvqD8B7LiDmBy
CKbMiFnYHsyD8+1S8C7jmCreL5lvYWeXZcyXdMPiI41OhVPiKCPL3FNvIzAC5BeVI3w1Q9QDwKjF
LkKKlmsld47r3U+JNATDij7PsSIDfFDGDn+K6FpG7cjZZx0ZOLJ6dnAg6o6WaH5nbm+dxRH2U4Hk
yxh2zL5gbafF0MPmDyagpBynbUrjQ4CL7oteu3V638E/FpRLJ3I8h2Al5PkwKmCCIM2BKIj9TEq5
Nv3QSmwaRCETi7Oef2dLelTfX3B/6xjydRGEe8IahYdATWhNzA8CxgwnxCXgw/2H96oRW3kc44Cf
vdo9FZJ+QcxYImFOXqogCzjdgDRzw31N3RBTnX5Z08lhUX1ok6n4qjWbRJEKl7sneukR34tMSQgY
TXEQUJXg3zFbwB1YHqp9UCnZBKMCmWl5sARo9AkbLinIFnK6oMQQ3wD4VPiEA1+agX7CI4sSNc3W
96WPDiHGyqcNsnMmohwNsqJOxn6F570nZQgQ/hl/gRIBCCaKmrVAAOBetA+t05vXhMYDyRVL7p4D
rZ6okO1uGXwaGv08OpSA5kuIdOOxUTUj+8OMt4Ln4whYMmJ5ddTAKHfErW13C7sIIiTBFNqla81p
gBp6CH1GKfqiF+3tx5B9F9o5tp1NWZDUseNgjxk4SBZD90PQhKvhffpUgc2LouQaZDI+LDEX8uGZ
5MRoNudmTguXnptkeF78pGOki7WBv5uA+Ugd1BqLZUmo33Gu+PbhZUeNQ01GQDQgi5P9sW2ksBdB
jvhQY1MbwbrO2sJfUSMNB3P3dZhcJlylKVBT9MykaT3ObB4EjjSVuV+zKCcdnGP70ra5sHhngjPI
OWMFYPF2M89V/mhkTO/zqWqZJIruRoWsMTkM6hDCXVqjZ+iZ/T0TMgVRwQX3yFRIjbL84D7vhBBR
xYKepCCAkUUMneQYtbj8UELkmQIggiDpYyzCR9l/7kGrhoUBVUukDXVDxBx1lcHQbr/vmQpdFmy9
uWMGvOnHYysM/4hs16+i5pGjsGrSfVKDf2VjiLfOn9nnfBp9xdP3tC34Oo7Ekqk21bw3tKg6BAiy
FWfKYKpdKGXOzigt4UNo3FNQggzL6/ezaECT1PnqnK/2XTyT/Pe4WbDQXYDstq8SgAmIjlD40xP5
gTx8KEnOmQSXfoC3MNuHDQthwb0Jd7WK1QMJdFLdhepM6uW1PFphDFsPWwIEZpMCOiZ9Ajfhjh1G
kHzINrmaWZi/JaNoB3GLSollAEtwa3lyNdfVrXUU4sDe8sFdlN9X+zz01MUalRBhuAXbpAfusMmQ
+O7iZmL8sOuWt8rm+F5EfrSeUgB2JkSxZw7MePN5tYHGrnVUl7r3dEImXPipWfmg5iLd4S1jRvOJ
FI6fxR/f8dFs31WlYgHfkbBj4cKtz0h/+zfQ8fn0ORgl++18rtq8QNuvA72HHuAGESke02pepBuu
xCt7ESj4gDuNYP4kItks+FuO64OvFeImg+LpTKep/WrlHehuF1u393GOQ5oWXhvGFKOhCMRq7Mcf
SDMxDnK7ajUUrqlSTJcsj5J2M0y1kkvb6qgWeWtoNGYazz2Q/INTlFWJmnIsirpwo4+RgZx+HfKV
J8CQFOV0EuMD3Gbejm4VZ5pNDuE1K4ENIls+KG4nCw00pm5a3KfOa9qVj7pksA2EwdA9VOxxfM/B
PipZEw6Xao1BRUtXhOAVjxG/HI3A4BLjkjQ4fVXXsGrw9TBopDYd9qAvXFqqLUzyAivPuuwBVIc+
LiqOS2UGrTXJCpH+uxruS87ntSvoKJDRD6YSCpw50jUyjneXyj0qznBTICn4nMsM27oeJ52bc0E/
OKlbBNkJ1S+MSgSPNCb22uAfk/p7VKplgEhjyUcCgcqKnpQhtDWJWiprsaEK3khyXoBN8jZQSHl8
0yUH7jXBgVSfhStogYQpSruJ8qa5mtRYQicCux7wcPVrI4Ip4HMrWomeWwNGDp+/L3SwHXrKR1fQ
jUnhoEyJW54ye9JS4cQVLtU/IHfZ5o7mirldqx4m65qIH/d4xukzGxG8VK0TbdCD+8p+lI+j1xtU
tOR4mY6EAfDaM6pk0EJgPsXjF0AgAhP8zuDmyvzDruBfkusjYPsoHvCTfVA6PPfmuo0svYYo5ypv
0mzQnNznR21xDT1PQyzr01tn+HdMdGxkszqRRAbdu5NoHDxQz7Ay0UurSBCzrXjikWjMQuoljI8d
fLkHVXwIxLuw/hduV8MTKffSGTFxfeRsq3O/6jAM/0nM7RUqT4q20BLRfOaKRp0mFZXjOPphwY0b
Li3d2dHeo79nFDjp1IroMSb/U/V3Nut2EzEJomtC5x3D4LGojuFi0roZQKkQUwl2jg5aHBy7vXEB
rm2Qt0yQOavwMMKfUJym9QHuvJf+27vi97LdXQvbu51H7j12in1QsoxkLu3k+apg9fL31ONaIucG
2bHlLyMR19oZXNIF6NueYfqt5njDTwokot0M4FlzikrAtMbOfrfky4YEkM+WUNBhhpBnQtFrADOB
AUAc3KMPji+MKadaF6anE6+o5SafHa0UwXga7IWbPOzeqSNyKmDjwRqcvQDbvcCaec0awBtr9bPU
KROiCGtx9j1PNIzSjBYmO1EQS50woWqix4CZztL3LyGKnyR1Qis+qMAPA7mgDYXVSSW2R3vaapRO
PjzUmvO7WU8fd2burnWnrAqLz7GS44nPf7Fn/rtttBoB5ZCM2iX+ATHQQ0rMtlrzQmeg2GPGoOHt
nwjRTVe5PVTiExsJAfxOjNEjVGYxvEeAny0DNwF/w2b/DDs3hRNj1OnLq1vliw7n77A12EI0b6CV
NI0zlfykWlLTKpCHtM3+fGJnaVHu9pLIpaXcgEQTkVZCPLnJ1oSmdK7pLRMVNIASWOZoHaZWyTr9
G12Vs50qgI6coOcgNrSDab32H8x/bBKTF8Bt7bYv3fkAogVs/wBgPKoy1fQg8OdSS+eXFa3AVPri
e8pRQSbwGrf7KsnMOTovXBP9G6QMh1Eg8esio8oI/cE68GrRcW7WE7p5q+h0VoG3KVeL3Oq8UHiw
hyA8Cwa7fOe8icTWTUtTHrUJ3mvmc4qtuw+2kgIaOES3+No6Xv9GjomPgpeBEjbYqLy3fGMzIKCK
dn8aDAqk/t8c4Lh4WGcKPgk0Fs69U5x24InAfksC/qJWD7VkTauKi2uO15IfygYsNMnbQGH0RGIi
ZUtdZ2cvAHa59ZMPAeRDOwHwT6rE1LEzJi7cRvq1jpDv+dpu62ybrxdxjHMWxyut0MddlI/Ga8qw
JOJKIrLQ+fkw6wilV6vQHeJYVHdBiPrigamuOzXukR8cZQabYYBJu80c7N/5LqI6cWORWSVgEvJb
MM4TY/ax588ddt6uGNUsJl9a8s15DbHsIAiJ5fVGnPw5VA1DYL2hsBwyNZljXsTJgNnb5dstd0p9
xbxh1oT369paUVIwSHk7RN837UmGe9aaixHzA1c7RWYpXzjkzWREATP7R0PltLwUOJGB/gNP7lv9
6vDZhT7MGYMStzxKY4k3dwXRjO26hteFpAi8+Kk9L3nkB8dEIsnxOMNXhHJ0WYsMKEIUfd2K74ov
BASISLTMTTzTWXBqDwc2M+xjEM3pO02j0vff6J0ksKszhFBFj2hg5owTLxkI3Ws11Xu3yCkSyyy3
VFbuO9LhV+lqiH85a83L2c439vKViYNBhkz1MzsKxHuv4ah6EG8fDj0SLqpwxCRVnHd24L5uzVjr
FLSSCCNtpTFOMpke9eP/WlGUrUiEezxiZZ6UAqzwK23w4Bx3BAlkFdUwRjvXRI0cIrcwHgx40HLf
5s4TcQ5Utj2dhovv9Fn8wQP3W60WxFSAHc3tQcp2W7a7iEg3pL1+XbqEc9uLVMfRxnahEDHFigot
+9DuBePELkfpxU4tgLW8SyPuwmDGurdgL4XJZ0OaNqpmlcKjREL3tuUrR5hGFP0/oZBKd5o5mQVb
ba1F7MdAkxo5Q7anDKTNZaXfzXhUB/L+O2rsK0ZzAatzOqPV75a4m4PwlNbNNINw7cdNGqLWGwYt
xBd8QbCKBz9+Ml3po4wbpJ0TXZwJGjGhpULGAru7EECrNUpKfiV0ldPMx8xYlOQVHxYivzMGKC09
I7ztimzrLVWmTvazHr/+vvYbiyYO/7yKVBDY60mtLAaUvETUyXuB10rlX2LQLmIgiq3CWgTKSf+Y
DjvzB4mH9V9aJqEF9FlgOmoYZg/cY2JdHMv0xb1aghsBrfP1SgywByoJ73QkfSRYIXXsM1gdXYwW
lurUBCwXoBKP98496T5W4lFC8LXecYu7r1xjXYUmCFok4Hpb9luTv7M3Y6KTTohmYdlYB7YF9jR3
a5ybUznSwTQnrEZaX4ybwryVZm9E+rFFqoTbCuRIjgV3rO6PJP+OX8B3UrSvx+cNZL49O4+mrOdL
PlBwHa+j4jrmapQmecMxRPOThOT+k04sc/8NODeMPhQuL7zHcpNj3c6iQSqdlhJ2ghXzMV97ithS
4iVD5BrEs7BNXWnrMw3YsGl8roIosU+jLQDktgSDz1O12p9aEfehKo0lKYV+U4SRTho5sWqlmEWK
pYgzKPO1EkenSTNPj5qHD8CWqky0VIosuGqGSHG5T5b9VJ+KLvQQFqepTqzoxlMtsRz8mKMZRBfZ
gud21KIiPev04bPvyKpekxrGIEwLB6Yp/BcE4y+JSB5YAirmevnXRs9WKE2elVmYYHfyITOi5ocQ
4lgwoF7sjZTlYGoRUvYIr7Mxjy6CZjal4ctJbHHTPFhGzXo0LpFY6xqQNBP5gS5YAOWXxwxuEp88
lpiYQM86mDddy22n24B2w8wzDB/R77CXJ7CJF/x9VbxbmNuM8OVhAbgtY3SFZO+E0R/T4hEjRXHy
nPaldIN2DS1KMpLp7C2X2c1csEuOvgxL3MAZOxeMLjQxVH9zuxFtlT603p87LgHFxYgTwlkvUw9t
WxuMWCF2yNVWyhO/VutiRqClMfGl+wRTRMDdd0Lnx7qtL2Nq4CFeffqi7GO3kj0wYcnsGVUsFkb0
uUuVi0KiEcMnJoCh5r3Fc25gYea8pIumb8LffU941X49vsPperYFa5vm98t5PmJsEp7k9L3vWQbW
xCWKpgu/fCh7JWQnE8DhJsiIwTXASfr3ZQoRC7TlUPpS8WdwIn4jPfUktjNAYEwW+w4S5ASoIpSR
G8jC4f+7xeHD9dfQTbj0yfh6FuTVzn3Qyke1IT42UPAMrSvHg7c5xx/9X7E1MtMXRdDYjzto3hAU
12PvRlSwyIPkNBaPAszl1FpJtIehQDoaND623hpQjcQvw+UnSo2qsnWqLx6QhwS4oBidmFSZapvA
B/6DLhcC6OXsa5eeOUVg0z+HYM6dYaw9Z+OOxCDdzzaHg2WORB1Y+UPec8Pq4/zips9nbcchZgcK
TcjN2WvMZnErzKNHlLOOuw+F3G49nn/srQQt5gEnuTdQa6ufcX4wXaPM9t2z7gigzIwo/akHANkf
oQSufhA0AWoPyUjPLPBkIG/yYu1BYVgg8ebH2/lGU9/6SSotV3JDzT35QRhOZOVPibyQ1K0aAYkx
CdZ/eaMknci84jb8/YO4zlibpFUW5dZtnxj8XzxevIk3K7wrq0moBHIDvOWVFN6mzzUqOdAKOWzg
y67mn8B9M2riBFYbgrxqDuB9hN3CA70iwzgYZCKuzDukzoM6YxhhZtiHhIxcBtR5l0Er5SCLjY/K
4pVddGQ3p9IFbjFsddr6bh+Nnmgc4JfUcdRa3nXbgOfl8kx1/ZnbQOMptxsyHhLxqhj4woyAqWAv
2D9a7M+DLTYISW/3hF2yIu9h5N+KYH+sWwu8FdzIqOpk8cj2H56mDbHCXE8fMSPUPVYYJHpo3crM
jztocEH5elXYGEC1RlBBGqIWMuF/NDhjfJZAh/3uKBKqln1mdkp4rokERmCYrDHhrarEeDR8xRdR
UvLcbg2CaBVkNGwEXnn8wYec6OY0O0BNWSbmzoO15ihY59viVFU+KqRJS61K3LrUeIhNTVbivzBd
Dyvb3p+S18idGsNDOR2tAq3uku+iAC9Prb8jgeZ+5NhvDzTJEvyLTdwskJV4J6GNM7OnfnA47mml
TWQwEyDVrL846ZbuZktQRFsjFgPHkm9D57xQ94rtkAa2UfyeUSyPQ2qCRJGiGEVe40legMEEtz6p
NLZ50iXCFmB4tP2h6e9DYyFItPIo4ztWCREBxEUz/K9QEEQfLZQHt1mAyV7W3IfjGqfYSFPq8lXd
Df/rM/Sw1aVp4mEzuRru+M01nCKvto2ATpDfQ2G/7a1GVgRk93r0kJ69AN3ueD+iHbsVNh8je9Up
b6HQHdoe4Dx0Sd0qReydvKfc0NIqJMHiLsnB+BBiptCpiieJ6yo6+MuMhr3/vTmmZMtu+5m2DkEX
gfbt8AP9v71mS1QBUIS5CwA7sTdOc1yQ0f549D4kBo+OO+r8ehv2RXXJdhDjngWuavEkqHH96K+p
Z82RdiJnVh/DWNBONfG/jUdgRXdVEHdLztAixxVSQ7bWqDCgUfm3U42yrFgMyGpXCLsQQTLr9xlC
eXfMk368SFlcHNW2gUodeS83CoxV3XgGTc6upmWHp0KOpV1ercSEx/xEiT20X5urRUcyI315i9zB
iY3Zpf+IYbPIaeazysAsSbslgCvX1sSPk2ZhNhYVjsOSCmO2399Xg0SHGrwjWRVwtbfycvlcT7kM
LKa4MsNGlPmnjI27kEmTJJPsSTaEfZYbJ5BWGy88SjJmiQjZEWwTvCugKdIb5QWmZYuRpfgF0KAm
+WO0yAgDWf4GV5vFlw1BNaWtmuwjQ2iEEjUYV0uHX5VOtSLQkswg0RSZuN2gn+yTwLlHUuVWGyQe
qt6prIJ1ucq9UmFOd4XvVC8305P4FlFqpcdwNY+dY9+Nk705hYBjPSz4FbHlpfrMwuN8/Kd7egx4
VgEQsiQpY8Yc0Jqw8dpl4JFKPXI1dqiAZfWL2n+K7VmduhLKxLBBgsULpbNxAwEb1aSyBhnZS5FL
x3MvN1hsK3nuKGUkphsDaYeYpuH2+tI/t1QOVLT9JnE4CaEGz+DGdRtGEMD/Rud+cs7Xv9ZRQiJq
f6ufI4VY1OwF/qU+1uqQqWs7/gzYKy5ScyAz9rINdJ6FMbWBh+DP5eOjwISSL6jhS46RynCqXuFO
rfGME1VZh4unzcmY2a5JjjcS6flKoALr6O7/L0OuzPFrc0rBKamyFpbjm9yYsKa4MJS8OXMIS9Kn
j6ncL2A+oN+ZEuyuloR/4YZlmAA82mDqMTt3hL8fNq9qUHjH++hqP21Pqw5SrRlyd4kjMnj4S5S+
yk4RNTQLezdKUKDFtu4H+BY9CPY7tKMWP7L6HWlbYH0nxHy8yUrVeX+pWJPrG+KP86kuSmfwbq0N
rxZjEVw+l6ofc0tspCFXYWWo+/T7lKspH2utJ0RYLCeRWY5c2FRiiyZ6e3I5w42vcLfAi2HeqbN2
giutQN5fxUWFSHzyxLaCuGBSEriPeHwp8QiVKgGCJJuIg1iVZ1iZ9PkjNPZPVRPmhhPhJsbi937o
TcJfCsXAy4T2c/WC7CFC4OfM8y0sl1b0oJRjM2MO2BnTku4sZacV/IYheH+kVBa6cro020SnUfC0
FW87U0uAL5E6B/4UHugT9bI8GgnS9EAxKknUnw9LLuv02ZGeLMMcEEWlefI8z6VqefrnaDDyt5xn
LJekwh+G3PbI6XR9yNYfKNFMUpmgU4IsCIlcpacG+MuIr4ruIytuGIE7UffputwOLaDgxSRLsDFd
gY79YLGq8QF8Q1rwbj+g6bvEhNFFkzJPNVbIoCHKSGwVIc2KA/ujYXDszHML0Glc+7i+d2LqiT7U
/cpNGPjjBvxoeNu5UStGeIqoXTkninMlepJMW5nLiFcUa9hAq14PpJALt59JWpTe5zTGUEsXqL6x
3zYB5Nxc4Q1Yh7wLyFCowYfnRRD/0qvlVxa//60sbLbiXJSkWdTsQK6cqOP6ppEt/D94sG95S6Jl
lfUVHd3GicOQX5hkRWB6ft9yqh5ctD5tbKonfNvzVsjyAxmd8wWRUTC+h0jku0mqNMZCvcXhUgx9
Rsk26eJoIsEtPNEd4dAA9U7WgOji0UQnGgIUbHIi5WmlDDOGkXeySPoSpA/LMoHhIE4GI3ROLTyQ
sXvipTw9VHBFUi/4ri5s7THwCF3zgUCPFBHRFSxl1C1aWHBHZodbleeIXRvaoKup2jjgXQ9wbtcw
QaeTPxPSi6G391td6Ro4EcFZeuzwMLaVN5mFlPmX1Zd/kve/b7aiZLcdd8OTsx4Qfj+0HzVwnlVf
CYxiYy1eiEidj+swpNnVzKXLb74LGR2Zahvte1IzqBIq72bk6kYH2py2oxwMmkemwzYu0dxAyy4+
uOkwfMY0DAtysW9q4yykraMD3kSsOH/gz1BvitevabEHlRblb17DaQ+FWcPvrQCc6VvTpOlH+7wH
PQxR70jgmyKw2QT3GTiwC28Ej37ZjzCd+381lu2L3x6vqCZNJBuFh5iJLt41o+mpqzZbVFtba63o
NpzOMGPw0FKo524uu3jH0PiL8SXSDbeezZiTBF/XIv2KGNi8zkFEGvPm/dlQYHOQS8xe9uz1KYvC
dLINTykrZQkX7Bk2kjqI/Alz32jGeaPBl6c/kd1o97LbyHdxJV40dsKdwduT1jot3XSoRLLEfbEc
4HSzjzXEj9EAyTA6tepzH9kg6S3nprR8wjZhpU+8wM30dQLV4nm+bwfJjqlRR+KCDDOD5V5VGFJw
RbsLcPG5PAALnmMJ7+uYkbv+P8nr5REGXZKTjCmKESHfFCWxFTLSQaYw9TiSNMcDDz3x0qmU5Rw8
WInIZc5qWjWkrxGUWobsIn4Wk0np7/BVFprt7zOpNMDE39YSriGDXDT1VnBjtS1WZl6l9SxIKmK3
D/TcE5or9Emy3ezsmIVpcljUkzJzKhKqCafweZ6iUDuX9cbVBfNBI2KkMzCjREc92FOIBQ05tiF4
4jLXEI6yWkSd900GyqqUeDAGttnSBKA1lXfa30AI1FkocKhuG/pq9NdBtvQus6b7jszRHY/ONEmd
hL2HC72pNxTeRq9uJlGR8kUEIfjvalFsrup7f8zzRT9IHSIgop8s93+lTo9Cpvj8XrSjgmS4Yywg
qCXKDQpjgxxo9eh96hYYHOif/yciCGsBjQiO/HphcoQ1Rquafbg1WZZrwCX6ry9sR0kz0H1KwZdk
+ne0IhZhlWnWj1b554xSSVahHRcfmW4TDJJVbLH+Ej/oW+ySTQJ3MmjCC6ZIlzqaYB85paEeVEbq
O2ZUvgnSX4TNHeHt//9HZIDZMd3ZaRqE8HbDZr8q01Q/MREl7k04wN7N+7Eaojx09Y+zm9XaeQCC
1AvKk8odfLvF/MB91B3y5gWE5bH5Gy+ocqYsDJMA78q+5axg9AvUCPggWSieDfzYi59uTpkF9Ckd
WMZeG+Orq4N24nofN/KNWDfkwUWZZ7nw65IIj+Wa6jgGqaS/W9Cm7U/qPknJf/Grrec4dbi/IjdS
TNXAHO3To8f3k/xJNxxquKQ9rPQf7ty6e5jg5H0QQv5Hk7j5GeAo/w7c1bsViZNuJK7S7og63pxj
x/UOEse61HwROJKZqbmdNtPXSCjYSRhtDWYNnQ53WB25K7njQJ1r4rF/hgTi60xGcqOTMhHkxggO
y19EoTMcv+lWSlF/4h9PfdMZCzLs5z8kHHVjwejp8wG1yznL28h0lUFckPR3GNaY6BqU2cgfUdGx
eLVCRpnSdVaxyBt+8j5+7mjZu9E7bmKczs3cL3jTq54sLv+Bugu3nu3B+UO0c6a/2Wm7EEfqpet4
8ljsfE/PEbJPahO0JhJt8IC1vKlIfZVC/iRb45Vr4pmjAJygTvp3BO30Ifs6LDx+pRrdiaWkEYw2
luk1Cx88VMHV5k2Ai8jswRYtH5K4pKUxSElyJ1XbZIve6atJWQDqTNjmcgyrC5NGY/PEv/nSqFDe
YMdDWijT3yMtX+UxeNM0x1XiR6n7C2BvVOw/Wy3p9pdsn/kCKE/++5gS/MlcG66wVTd5UiVIigsZ
Lv25WIqkPtIpqizmbj20WAEdO69IQMZ8a9zdoKQyfffM9zPmDoVVFLV0lPwPl5oI3E26R1AfLirt
UZWMHnT4sLOvJbySJ89SdbtnJdCVZPD+fNvgJjGytjbT1xBgyWRJ5B6n18YbU/dTyQDlOCRTl+6h
ivUUEAgvHRFh0br2bPeXvP2yS49CTJZqpxRuM14FCGacfCNh0vBznNhZBMoirRJLQtvD5EQGNa3g
pug8jpPZDM3n5iftIci9OCku/TnGU9u9UbVaSO0jlAfPkuSepioZX9mQbyJR0RfiBNV0GpIK0EDQ
gIXgtjyIs7QyvXKwm30cWw1/faRGP+UMyUZo2GyuRKHAZxLafEuRj253dnxWup/uIBfYAbaf/9VF
0UQqjQzHTwBC8wmWg0bHSiMBe1v0Yymtxs8KiJUqnei+Un6TrD9SYC9TXOyMTDEBM+8fGn52hrNQ
LS1TMaTzixxOqPmDsspKWbNAEk8RP6Ke9Ieg0He3ms1/ySBXPZDWcbi5GZNDxf44DXwILvnn21+A
fUuUKoW7XOx06l0EJ/PIQt1AHn4l7urn6cYAYKMzJvbd81CZZy0M4JbrPTXUJyTPnr4weocNM4Tf
WPnixVQSOOtVdXC7oucqVfzaj6fPvVX3jwprDeZcl/t+XxfZerpgP0uTtnJKh/5E3i5+5n8TjiqN
00CyMh9r/et1Zv1l9x0x4Bnnu75AivjmJwIPO5OzoatNKlCQYrt2ouxL3F2fmgyYFSPMGe/d3IHL
g4PZazvSNzXwOXe96ieeR6BG1RtCSOuE7B2dSjxDQqifPasVFOAtHa+hqL+pKGhGqVsDBqxqkTYb
OS1liORe6l353A7jxUi84xAbxQ1Y1GzPn++ryyLkv46FOuiuYtKUYtGXR1GQMLRHGROz60RuiLgo
815IwQI/x4Wb7553SV7azAKvHCU02yWSqu4lMMFbwTCcGyZUC38/9cJFxHqZqYpODP6cb+/IFadw
s3X7U2CELisp6te95qz2YqxjTVBwQhom7RYm+zdr3RsX7asMWfZuWmHFulSG9PznrDaDi52SUTSP
6f6GE9+bxwnaccbJ7FoHgr3r5woUPFClZOMyCyZr5NKw7ZZm3nM5YqqxMvNGAtoo4ZxjVOhtMspE
0QLyiDksOkeNLMTVVV9pn+Rnxo0yca6GKxNlhTY57l2rI3RgH1Czo5/6qaQ6Jf2aGrveyNxPBR3/
702vqalv9dH1AL3Up5YwXpTgjOhkoEs/RQTx8/R3fufRRQ5RuUeIElY5W23h/z3tOc8xrLloVrdA
v/bJo6u4xw5q6HKpeS5w59CCWJPgaP1hTWhg7rB0D+w/0Ekolfoc5UdQOQ6at20UNNAqlyBlhcZU
Mg6Xrjez8sP/tRxiPuJX1lN47dfzNk8sFeSpOqABqUyoRXGTeQU39TL7PHMhsyzKL+/8GW9Axuq3
xSfH2RgieSUQv16COKqe4OKVXvPofUwfeWmSm5xRKgFZkKJf8koBvOkAL2V9hB6c+f/7G6icr1zj
SBRXt4hzw7YkaFR7D5zECb1CnM/PqH4vraLMx78NknqCITc70ufUxnqIvnylaaQJyUqtkRlKIA8t
Z0JRrO/jZlfQnkdRzi+VOhsy6WUSoBQLJ9oH310ULmlyeqaBFAFK4cAUsH8k7ZdSNvm5Jg67SuQZ
QYZzybB8aZCw20zYMC68OGyqyCO4BsOryQCeb9MxfnXir9Ceq8nD9XJMjJFGGIAu8m0S33K98rW7
8MItEv1FVO00SATiCrHHH6omMwx4rXTHfTJxJbswSy8GGKXrXZuSnhXMBDYRhj6GSrC92cxRPGp9
QkvN+O2xY87V6jb+B2zxF9TaIwfsyGsAJuFRQTaWoOdA4pSuEvpiu8pzgkTMHOFX1kB5n6+TKeaS
ddFB7OzvM8I5BVSwSItNfaaKXL0Y8jtUuiBRSREUKe0Kf1a4Uller6Ugpop9VVUD9WvKt4CnnRFh
OFNCMQFGPIT+x+iByo0QiOiX2TpuT2DtSeIT17b2K4Qz+h5dIXhBpLRxQJnvlVtGZqYLmM4BkVdS
p85UAZzw7Ns4BTzoq4ffQOu2972Q8HBIQ7uGCsLUZ+EPpzSIZItONUg0mpO4G8s6UR7k8Rgg/11W
aSWNcP7rdWvk6E8pmDutM9txG4Z7e3XDWjmnZFvdwAHV6P80pPKZyFqJH2E2RJV08d+fvIOgEigW
xDI+tlKpT2LpA9C6kBkXVhYRGZQiPBZlAW17pcyLEEDRXdLUyU5+NhC6jssYi/0WJ8jzAdZpI0sA
HS7yEr2Q7A5pIRvCmKBfa//gq1NlddNn/kSO80daG8SBcj2Q/L+8zNkPDGIaV3/kn+JSsV/0fs/o
RJAYsGKxiYIZHw3BmUftqBcGs3qvL7bVKLtmvU7UT+3XipgkMDnz8SbtL+mEUwQt4TNa7EzSCuMZ
B7KzDp5ZkKgHrODzd7tufMbrofVhj0J5hqKxvhzncNjk1ZUw7fy0JkYvjwwzCWzwgiKBuzHrrXc0
10oIrmVVqbesuYj2lkxUZPIFw78vFFexnhbepxVs/frLCOyrYPiyyzFsKeRJMO+FccF2lr4de0Zi
hbiw014/tX/A9KCm+506FbYLQjHI2pGlybojOr/2HlJFMh6coogwNBfY5UVPqg5OEUsMKdcF3cZd
S3Vjo6JPW8R9pmnWqqNkjoEZOuaL5bzDz2GfdlIxBwHpqMnssrfTcU81NQyvXBOTCqcScKjOCbBS
CdFEKjny/siobWn392LOzI3bxnuIymq6DO4uZhBu4P9pjj6iNcyLjKqdRP544/+cxZ5gsYp1WoOB
Ocg0CzJvckmHKOaOOzEFBdyNYWHTTRaUQwjp/+FtpxjECFsCW1CVT6xFNzNHHn86BCGCSWXpPISy
v0mHoLhnvUaNwZYyFQoR6LGLTeJQ4V6WmzmM4p6tRIghne3ibIS064Qyao8zS2S4Rd1kyxSnlkdK
is7MKFyObxd+2oC7h37GN9qjWhdnv23AX/5DxIGZj4zP1662TYHIxvtcJsABWcynl0/2HDc5sqxl
MKkPZ+mvNrz5X/RbJrCcgwXBUR7XNCFDZpm0QILjStNj5K6Yx3b1Jcu5mpIHoRCHH2/3xskxuO2a
z9Mp47wjpvgtdjEoenXqC2Nrq3MZ0gzADoUQhtC9MvhSRDEhaVWIbQF4/4+ZENOwzbtMH1hzGlya
/fFgTnCpC4dUiLNsmrWI0mBYeItFQ5uvYVYrzdr0MVVC131yl2KMoGOBnYZ63FhoJBmU6l03c0q6
8YpVsQC/sFvCSFVWE3gi5aH8kILRhBxoiQno9r/+4HVUQon9GujjBXWgn3X/xG8fApywjVA+gyX3
7BLNsfL1FgkWC0l9POTFLwB3ZLgIK2NlEYfXkTx2Lw+zgKF+jhHEDkqJIAKoTnHjoC1LgDWbjga8
mrZxlvVSVcxhaqtVdo+RMKCmywhg1jwqJtLrY4TixheshCXHp/A1BBGMDxV2QlqJsssDaSIVxJjy
032VdZSZOcTR9jBLoLw7F7HOzrPa+Y0Ux97Ot+y4kzgB93NM1Ce4zg/oD6dAT63LXWJlVCVAK+Ng
0krlNTmN7PI6Rs1XMfc3PY/ksc/3qFbUE+iXopAfCOymi5pqmS7SDXq76PSyDOkQ2r42Ux+YLPNi
NGuIx2sLL/8ijLxLzuaPWHDmbSd5ghpkPoOjucsJwQTTI6nNfkOHIWLo+bLR448XEEI5SNxV2uyJ
RgHs6uUo4WF13GcFv4UpG+nXKGia1t3wIvPiA9/rbQuKCq/iIitH+K5sQlwhuyyBVI8qcn4ADLgL
5x+ttZR/PoPBEOWFDviosQrYQmQ/Nlde6C0XMCp6hAD4HLt3wrl0BBIlSNmsGVVXg/uqSnSrPyyn
Cxi9PXiBS2KmhyA2xNpfsWtXlotmxvNA0KjJyuc6BLijfTSogCfJNrD7NWyF3C3pEOXFZF7T0svI
izyG/26mIx/aP7iwaPe2WVmGvh7Zh/TJCV7B3QCcnasg7JeFs0EFccIrV2VDDY3VFVQugUTdxrwQ
q3z01fcg6vrxfja/9z4kET064KonjQHKnb6cycJq0gkUzMRQ+dWL8nJEsMH04GoYDYOXXFUfZ027
/97thMYxSyO4l6BthfGIhNpHK1iu0cjReWj07r1UTiWJizjnRzeKzMGdoKcViFGBghDH42kds4Kh
pa4G7s4CYzWWwpskcJAOoLc5TCajBL1fbFDjp7PeZ5b03cknvEvUaRzLCJ1dBJ2OlmkATN/DUks+
vDPsUCqrondqlMGfLIm1gcNU1KKu6c5mk6IpXBXiCTChTGMXRFX1Ym2bVTW9Wm8Hk9dIdzD/gUt/
9p2Gv4Mt2FoeQXZysFu1991d8fyvBqv+xLGlMHpnmqgWEuzO9ZABD3nKHh6nSitaQyT5ixOA/rIf
WBHG0iz9fX5zR7KHHrxc1eQiyeX+AMdiga7KwMgg8juDrwfvTDC4ABIkTba1lovTKFd1txHul535
ZsNGJvhQPEQSqXMCVdjB56JAk4EStQMqRP4J5wwBrg8looVzYam7hK/ocqqRvhonfY+6R5ymt/A4
Cw5fx3xA10WSEld+hdBmzG5IUJG/ZaaM93y6itgsRFlGIsPvs6ebQcbktwJi2+agcHFlY4Bb3NGW
cJ3XcLWQlRLW6fsp10VBuJvgRHv33gN1+ZJZQaLHTorzqtI05s4RagM6icZte3UP5k8A/zZX53zN
EtQYz2ETHdBfeoT4k8A0WM2yqhmG0CKhmmM+QXuW0jsUdhGYUpfYc/Z0lb2HGu6roHmztL03uaGP
GRp2mQXc8Wsyx1FN2UJ0FLQLNndBUnXc3LBWKoESYjr/zi5keXPw4eqN5L0MW+eTB3h+2FkNeyJr
wGmsmsQMemGmjKDGDC/uNSUIX0TndpT9CJ+0evPxxTiB25rp3dORTRQn0y0L2GbbQ3n5CO7dd6YN
sKXkL7JDPxdDtILkZGUodJnuTPBIi8B6kaILNXmgo4KFusmIpjva32NURKYi6j0a1p8hgPlx58Mb
JMy+x7+DSXlR7igD7D89p08cFWIQ0Wuc5RXCqq7gs60s20P+fEciC8CHktTswIDuSxuAUqn2mM8g
DtXp16QseV/7xMtUjHi1x2Yl9qtx03hn/FLHFjoEN49uC57qUSo4fJh2K4MAQ80bJkfBD1mzBw==
`protect end_protected
