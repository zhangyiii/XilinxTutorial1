`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 88208)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAIeqKFUGO4yeIvPz9KDWAEA1+ZJKoTrshAJ3xsJapha2SVjfJNU69eRs
6iDzH4hh17a+LMeXOmU0YWV9iPgUD6LCkn8uLvB8MHPVPgJFZuuLJyLz8J+rq6N7UDABCd1hFfyR
mc9zMLesQ9a6AXtjZeZP6zyvsA0AKmrsn32TV+lalyrMA9dZ/shkK5YY1jbZaUgr7wg4bVghkHiZ
5ZtrnmturqwQtubVbylgbRKRVK3x/0IaByAh85f3rxA3kW+lwJIHryl7J022KCZMJzEdLVMwYtmr
P899h2v32Hhz8FuF3EsupXe1go8qitdv27BW6BzrqWm0JyFSQywdhTtfjSx3qwpD3xLsioWS2cns
TnLM9ZYBzuwicONRqwrAC6l5fesiYZgZ3l6yLkYWBQLJbEhXcnO4GIhd5h4O635H/yWF9mxhO44O
FpBBtjX+eMh6yCC+MBr7bGqfROB2j0slEfVBfoXrvgq/9VEjz2Cw2+RpuU3R8NRXA9eBsss7kVc3
JEi8FxmoxRsYqmGY07SqpEySEB/93/tNPJQotPSnAfWDPVlF5Vr5NxnDLi5UtX8e0VFoKHsud/cj
yRp8TLK6jHnXVXJnsG0HvU2DH53S0cGTBsK2QZcBvBDFP9U/Gri1+9a4htQpEkMgMSajP4Mscrpj
4ABg7USG4tH6r4/p8knDlg7wMKLzmbLDc/8olAVdVEeKwc2fwjmjPbsLntlYi26diT+h/5pjnnh1
Z+qp1IT2pysPI/3MGTXYJaHNVt+rr/TNJfaCx4hVqmYpR41GF4g60VD19mT918hSwwXjsau+7VMP
KZAq6jdpNjuJVXHp0pjqs+Tzo02zGPs+YPO7mxWXSQ/n1JjG0niab9OUZnaGuR6z+d9QRQpbXQzW
drOQ365Pe2JpeOUlfvw8dTTSEf8Zr5nj8ZgXvJvvdO//5fVGWdX1y9wes5mk4EZJuqYcbl2otovT
0NSdYLuHlT/Qi2x7KduOqHX3ZzUDKmBPiLMCR4Y1s5gcEElztqt+98Jeegec9WpF2W6r3e3pvfyz
jgRM/qnw372WHoWACToprjuSdvNsYzxA2wLCfNldPUjqEhowhqDPcDukYCxEgEE2u3fDr/vBGYvE
KHiytFTaPD/M1Aj3tMgXiaErHNWy5DSSlgLZQt+QU7EfqF/WP4K9l0DUhGKC92sqwM0Ff2f5wJQ6
ODjJKFanhRrsv4GvtrlLmqJVeq79wWBQa3AGGwLvm0tY5r3kVYeywK+nW9XOnkPDw/TyJQCk8i95
a9256lgvzDh+V+AKkJOBulZKod7Gd+sQSdE8tL1lEK8vQZUZm7+FKZbSlhVlcb8ZFswC3Zvys0wZ
mxncsPIKl07py8MYdrKR4cE5nVr3V9y0S+/Yk+ggOyeqbP9GBapceAVaK+bnb2ijVPvwxeryoDmZ
KBaNScK6gDneoqzXAq0iXTlVIYETs0oq03sMzOSNqh/RTc8SkAxTX8rMgJuFOdZChpcCgi/ViD8V
HtTEhSHx3ODcNzinPRSt8Mmwn3QBPdTVtLxN4oZ+b+zYY7Iy6WG6903qzatRVNeSqCTz4G1KDH2q
7gvZQ/D9G1iXjk4nRCPG9rH4Q1Ny+62BTHP3RvLTLpI1fPwuYhnXkjod5daFQup/BLvrqGpViFx1
dls3/ybtWDpsaiutzf2H4s94jrTWh1m3foeqxnXbKoB5k3KjrUulqWG8MXBfrwdpHlyEYXpDns+X
fBhsHY22W/K7Gax9MNd0+1DE9c5GvuQQat8epxbfXkng1wgoLggaDjHw2JNSpmMRVLZfDJPVGLF8
/zatUqHSPwGKj+S1/zHt0Nf0e1yK3AywTLgEus2KVROr44Elv8J9y0tmXblNn60EESa1JSEcR7iE
Y1uSLlAgyBWB6yk6p6W0/UCpZ5f1tAwLn6+DgfoGz+0h21sZLWiQemU+s8LkUevEI2hqZq5n4h+M
Al4J0wf6zgUcwNCxAekCaWvjZPpUpofw3oMppQXFpnS5qlGsRRpfWTqk701lq53eCSJadTfZC5qt
KG2Cw9yMEiWjtOhid8Wlicd4nlwuNoZBX7qr7xGDu/VcA1BR8cUzFHVMtZCbyLcec9n6Y8ekfRt7
fjsGT3hJkHF7nNkOp7/O9uGaFqxqd5i13zCbV+wU7cYiz8cUMP6ngf1TZbzuHX5L6p18j8M3glty
jznYL/gejO6ixOBG+SKbQ1GxKgNLcO+HUvdnN0RQmD8HGzbD7EtiQFyC/sfF6PSB8PiyzZa2T33G
6JHQo3hBDAZ2uylT+xBnTDj/GiTqYvHlPCDSGt8cg/5iuAfEyTVBEhEyQJGHMvHkDfzDjiohHQpc
EET9XMo52xnbDPj+q7EubuWo/6JB5H790KDFLuk8JkFGvTdNSGViAcegRhTVvMZqTgyn2WV3Vl+E
hJuJXm0N1COkGrx1GKKxGtOcHFEStDbUfn3cD778rBcMW4+hvJyI0kiKAP7STEvQ+5qHaDVy11Bg
wWkTFqoJI1jxQjX/WgJEqFFILZaQxRt/nToSp6qaGRMqebwTVsjuc2v4+M3VnsTzQYznjzyzfbTp
O583KtfAQynUitn2YGNFgtVtdq+YHgwfSmivFGPc4QGMEkFX7CtF4KYqOQNA+wBXdsKeXY7+JQba
/lGHIcrh6OD4eOdh35B9emKde6tDEtx1oP2RgY6aeVs7MaqQC44xt3+7f2sl8UucmEliIStnL2eN
7uWkInQYTZSw9wnAx9wB8mlE4w2/cI84uts9RcKsSFR3YiA7N0BeuySfDJeTbNiUkLQK8Q9BvJNl
5rleeIpxhpvH7VQ0NmC1o6ZGpzqP5V3IN/ZsqRhOwFbJ/DIwxNeSa3r+0hEcoGzxWQa1fMgjMnm8
TfzLgg1civeBMmeNF17BTmP8kbRLXTU4HsIFlfv1+JfcTRLwEnYGEYSmgxRkAqDKLDNTToJwVSLi
jm+kT3PwrCuaqrDl63oy8sEP9qknT3fqwlmsCq8hkvbPlKmB5HFh1bbtF/Ht5j4b16W9VhTRzCzI
K4uMk74j48I8CyI942/oZNQgwl1CGI9L5IOPDAl/iAczLPPS3m9VLPT/6XDuf+RWKJinktU3QkWa
Fim0nydc87eI0MXJ/emTZd99gHtS8XF0jUReERaM8kpXC5pdSQimK2ZsVuCAsFtqNKxdBhkFVDHK
Jsm32yUoZ7pK55IMmMvpJ4m1JHHXM5t6Pxm2KLzqrk6nBz635q10m6zHmsz7unoTIJnZM9KilWot
RsjA6zHjOmFTakwA+iA8ZdahgP+pIlM9fOu2BOzLxB0CeQ6xFGjOeQA6oh7ceYM9YSEsPGVw6ZTa
ttzvLO+xQkP8wk0Ujxuic+zRFSQz+BJKrvnndDUrEfdSbBwDhFdHIbI1qA/2PEqRqM+ch+ReEXkp
qt0ecs3V8yZ0kphQgS2kl72Wb62k8NTnQyLNrMxqCJmSv7tciFr3iBpg1JB5yqNMiHF57gEt+/zY
ol8cbsBcMaUYaP89AfKnsV0+zfrbsO+UNpoDeylbh9S3C9GKxLR4wye7wSNmlFE/d/pAe2BmcoKO
g0kS6LXytudqpJYCDo1//78QdkBtXBxrwnDlPKrH8yxzCiTRQxf5lfbEYZPYkJx3BKBZOtwpPMUm
WTjSYCDB0qXPg14+/nDOtBaHdA9ZBuWwSEuP22wEWtdaXp45I8EFiD3dwbThviBADpfxycwylQMP
UwHcI+NXt/ZSQLihwsDJ9pTd9+x7fZPVINSmc51ZlNiXGspH7rHX5GofTfVB4yNFAo2dP/y/dvcf
1KPhTkdP1jcZKjiLXpG2kt6mUYsN4JNrpsrlw1emXd47MD4m8iwcUB13JW9JynjD2ixI4pP+4P0y
VfxNWiDHf3WPWSUt4lIdAmLitX39BL5yPEh7MJdbs+Vgr+CVSJc4wf66HQ836qX0TE8tMzWi4XWq
aGlGt6hKKJojUvoo31sn0zMNBYNQtAIQguQDR1ucvINlP/YAlgrBuYcjWMorHzTZRF5qknXrvvbu
nPu2zsj9RSscz5h3oF1pMT7xpBJYftQWfA42ZLjh6SdKB29ov3Pg7V8L8+04Au3y6s3Cjg0J1Kh9
Du0j7qD7tGEFQNrGleuS21AefuVKR4AuQh6pceBtFOEssFBxghE2ltFai1R52VcBdivy0DJrWfNG
AddnIKziaEJH51OrIkZUjHPzbU5QxMmy+GGxESq/T9d9PXF9lxHfzkxV1Mi0QU6H49qY5ZbbOzk7
TOYL1RQ72Nd7cmtUsc9oy1tCwKiVnVYBToqzQkkBZLWgIp/r1CdUDwsU023pRv2iOkUQ3uKlJ679
c1/opM2DANWptMzTeNSOoj3MSet0gFl2umX9FuEigdyyeJFzb3BwDY2EpnHCFWR9FVXSi4rsQQvf
ACpQKKMZJKbQKWgY2jUHEjtzrJaaKqGb1paqnVdueeyPLUDXFLvoPqDSRnSvJOs4GAmlJCum0Rcm
Qk2cltoY15QY+65RWGxTPhdMQaP/RUBot2NyHUTdxQKzrbhjPm5m3Y+nL6etrgtDSewEh4kP2mA7
yqEXMJ9/TZRPqth7Ep8l83qFnv47dO97c1RDX91+otFtRmPMklPgf/RQL5oDKMvtjAqLDCRa6184
B3ruCGCm1DyGo73KjdOjzsyueMwN2FlpxepOZbyiEWEHLhqM8vqyDA04tLzAYtmIKrLRgY/rOwfz
wKtoD96br4oNaeGSQNiBfTW6wAhKlRO4teqwCPReEPH4GlnbLrl2Nm/G54W00uSpzLuL4rYG4xRm
zcE09OHiZKhwHlkH9b1uSE8EIqhF8SaGlJFIjlA8Ub2rdUfrIK67YHCdDvzsjXbyJssgPgXe4Vt7
6q6LO99MtVEDAp+mjvBM4YUlm7oiv0JWJrgv0MHclttYs7GPmwrIwr6oASRKyoxCRx1MwXwbM3LK
/aWEnqrOsts7w8TylC/ENxFNxdD0c2Wucqs62kux8/xPND+qkao1UpBsWHxjZLyaF9LN5VH0aOHb
Zlazysp/05svEerOCMMqy9QTYdCoPwA/FldGpYv05vWhvpzpjo6RA2kJSs45xrGno2pOeULip7uq
yxeyNx9yVtv8cRuIq3AbZUcwYe/FhNF2fAttqGxU9Y9men0SVdPes/K6YEee6MVis05qNQpptjbt
IZQlgnCbCcw4Fc9tiC6GMbL94dljs4CoysnHKI22KC6WEN2ZILJpq8zTX2mPgWrZ7fWOURazEos+
eXum2wsJQy3zgez9UIsz7zn/5I09n2BhN8NkdQS39I0hdwrOxyMALoAdQH41cDYwGnuiU/Huc1ng
ioxik+N6GJAYGVm6tgo1VS4wWt/8Orajt4ZSObS5uvzpqoYbzQnCz6DdsEinpxzVsvhOAfg3ISe8
DECeb6c1cXhLSUQgJCGA+SpMFVMFk9jcvOren1/4eEVAJSDltgUISBGzZFR/D36cyryFenhel1QZ
BRyCQOIxSGqgvSfO+5j28CL7BsaH+m6j9rDy/VT8SSMk9kc27pm0aiSzA6gfu4ZaPGdderCkJ7Gw
xI1b8yEe6rXur5yqY/0M/uz8qK5PEyLTxjEBjX/L2KZoNVqVoHGEybVZVNZCOozuLDtz6mVTjXZX
e0QtU4IjM1cRu/Zr6pPgjJG+at9uOY/65Lh6OeoN38mEyTH4R69InGiLkH6GYRe26RoqoBa/d3zb
NJwYI7SOPCMnD1adP2zNDtXsrwJwDqvsezs0cO7oXXThnYGvp4znISUMQKGxmtILa08QxgXtJ5rQ
XgtiyE/JEpuLQg3Cd0RWVkLolkvn4B7O+QPtW7JLtJvLQVpPKPJoZCMB+rIMqxK/yv6tlAHpW2yQ
+hM/rkbBH8ZmPKv1DbJaOwDzvl/3s/R3MvbySvudmjN3XKPhaVdkPztgdFJIqKhZ5YqI5M6JBGvn
o+BE+U364ihqGaqHTdCSyud5nUhW8obWPEKq7PdFnh+wlsW77+4v+p9HDfr1BKjK7srIEIb8NXsD
wDzrF31L6NoxiR0ZdqZSvk7GEop1rOgBnfTJp4YEtKFm6Woq2w0oLXhDtbPO+4nCUEcQ7/nJbXmX
2gkvkMBT76X6/zVDOgzCzXfjbtpdsSO+elDQhnNBFlMrDxSY1nYFdKptxSiVMsvVlIdF5S+IQAkS
HSmNSmkO6698B4NSLnyX1ocoj+FdbOz9RX1sId95WE+1QxUIb8gr4npulSMLh8Q7vYcWs9AnqTSt
hfhSJB7w+KjuMzOM1nA3pdXY0vi14EGzsPW8fWeFpTV7sRcRywaYIQoSVAIdyNIbsM3nyIcJ9fMM
QmH1K92oMYfxFsXej8aVjxukiVSuLy1qMXVXp5W/pEdMEiX+KpNMhSmPiHWesGPxZ6wQvDJvPoSO
KiGlpZmnmxc57pzzbNFfXE/MQEqE64w1xvgE5OOABguKLv6ElL9Qrn/SMIE5fazFgecyl0mpX+4s
smrG8EWO7St3u7ucOUDokAFDCIzHZ5sAN7nHXjaK48abr7ZDNyDiaUtogARtiParQ3vHdsAvgoNe
tseKPqZkUEOqfAySYbxZ4wzeLPAxVysm1Qt6lok+IhQCbanKjx3c5fI5Ad//LJnyoLUJdaAuPwK2
G3wwXgCNDsvERtoWo/anuZLvklvi+Nqw/euCaA2YEDpaWDP+owv1vckhlKNIcfTZA8EnRJl6Wr7+
8/b0/3Bc0xCNno/YxwXtGXNaPm5gjD3PPXx7UIdBjQ6I9MyIvRZ8rVS2R6d0o33N7s9cT8d8XveP
k7RAfNfYILtoWi8DE2/xBlEfrWXxaDtTn4p4/tNmUJQTOKxmRt9h7K4NT0ZkCkEfyIkGoS92xxSa
jxqc3wKGWrcJsro8b7x9Kr1LOnVmckbJNJroLT+On1a8lrvBbPUITipaRZgGyaHWSiv82GrSuxGb
8JNIRkxxcl5G6ou9H2gZduBwAZ249cZ+WvrmPj0/Bw8zJU4z9yGzLjeRPCgH3mtdBpyYXqVyl3rW
NLh/MvltBTfHlTu3SWHg/SJOpYNETdS5F2cFbK44FgODAjVQBrCbKiqFSHuGpCyH+sYPnhHhfwKH
l5Vjq5HfXkDdGwoSl3r88IUawJM/B8cBZtHAAeOb+GrKyJkhTFHTT+/u1YIXz9o5hoIM02hh8mV5
Ux58WFKRVQ3Ob9mIVNwuPnB0YaHO6QYeq1DUGZyWHlkPjRgMGD+lL5Ky5e6wJWb63tT9XG64vsgA
cFP5AW5UP8C5VedboxM3uYYZ95RGq+h8+pLLEtfgYcOAosegxGHw6jEzmRPqIezU/w5+eDqs5vOW
deqWOmDipEatSP4dSVNCtZYj/+ZZRYXFxWuutmE7wzrxmbXbcGcqm47TND06k6PjKQMA9fBoX+bX
bOFpcQm/dwCu8vHP4q9Kwgq0yYdFr2RGZMMmXmEKIDU6IGtPwMjq5sQF922KeOtTt1IxxbrrKUAK
ZBuwYMfxnETQeT53pdyNmGbs2YoMnW5u8uYFkT9M4BHgiXGMdT/P7i3GX7CDgrOFMLnsBLLC6Zm1
3LEL72W/KpQVpi9Pf9ocKDLHx3itcxCaPdoJYjgoyvFnOAnqe71vuwcQvnH4Vzi0O+fs/u5S+Voh
J0Iobw04nxboqEKlYXZOpKFPMRwhop31e80Lxk/hO7XTmsBvI69Opn6WkZu7FbSfL9U+ACRQsDND
tbPpA7tqWB7JdOfz0cnP6k2IX5aNLM8yzpaSTz6FBULqMzkozJKXL0swAbwmoFIHdhes/OK3Rd0Z
bkRCPED7iYGPSzHC1vpf+GutV2EX/Iio8STS5HAU1XwouV1LRbur2lpRdoBTUgnnnsemUO+qXWST
rOxmmPEvQdtbsZDp+OvIrNfLv14NE0kt1xDifitTApDIz3d18buaPM8xWgAby7gKv09BCisUQ/uU
MN1xropNMDPv9Yv4wvjA5LpxaiQGH4AIwB2L1bnQK2lD6YyXAPI4C6BGGHqkxolGX9qSceJ8Xlmc
qOhNKqo021zJhKnBt0jSy3p6BGP+SC9NIRLERB5n6Ge0KXD9QSQ8KdeqHDmmBIDLnOmMtM/Z9/1w
O9WWPrP1WJDasgJiy0ZI4RbkqgbdMyIlFqexphrAQ8pQFp8wRWaTfWFxsngB2yvIQjnKvIJsPnHT
Zz0g+ef8AjGavXD2eOR4Lik9J5+5nDd3ME6Kw7x4N+LCBzyH8FYwibU093wPwX899bGBgX3y0Chx
Q9bw41Z66JO+T0sQtpE9Y+5OQ815JN0ccWk9Le0EBWuoSp6SYH+61f4NWgqNoF0660j6kIPo8xXP
mNoj0c+Mt2Hmzt+rDeM7gJQ/mMlWK8rF530dFFMett4ByRY4L64dqjmJNQGdNYuGcnSKS9OYuT/W
tlNd5LpRCl0yUwAf91HGvpzjjtIoxbn8qn2mFTIox5FqIgD3YzQGCYikE0NC8q9UGR6F0uh7cSO6
t7wZK6govW6+1RllNh3CvzNCIxoA6cEqWokxa1I70jXVUM+vgKJ5M7fZaoUAZ/IXT1fdAdQl6c7W
ULHOpmsFDiND5KN8JXX8H2RTxCcXsvZJhA6sMd6e7v751u3uxjUyDqZpI+NIoeJ7nDUPLPDk33j1
6fJCM5o505BdqjDUyxPD1ibtCucgFu2vP0do5uYp+gevdIzfGTji+IO5seiQ84K1UdMrrRqBv32R
wtGbuoJ52nBl8oCJeZcTPEundGDANbxsmhyFSZHZRSb2Zf+4qxsg5kG7HSkLorucUlYIA7iqi3gH
GuaJf4dRbYfKCpv8p5vS11S7FlokJQXtqfNrC+1mW+q6sMDtjyMygXVcUpjA7cmn6iC79vXPlNBG
64LpYDMyJQBnqob+jCl0La10OibNV941/s/Rd+OFz7xT3jOYwh3l63J8LRVgYxxh4qioK5/eNb2R
fpnehLG/YALM7j4iF1rK+qWFvQVe1+Son/J3Bwn+oXS8Hx6O2Fhvymg2A7+VbzoPorPxvMC3IdnO
sLOxssy+7757zl6C7sCNmkI6RvFvjZ4HmjnUCiHrA+I1p52OPWKscsHUi7OZekzwSMHr3wcRxrOZ
hRnZ7UIqzXjGIhdqiiBJLqJdcB7pQEX+EQFjUCWBkdtnufhiBnWO1gHZMF9/mtfeQNS8ef+23AEC
8tsfyGGMJCB4hARK4WrfjCP/hYXi6tlhjRSJ/eo0FBLGYg3fvWjsFWOVbhMc9RrFQsBxi+6Xygc0
JLoYJhV+wSjIh3T144cHtQer/4ikeZwUJ/lCcu6DPYKLbD174KaoQ6hSY5vpCTPTL8tuLQN2ZyQo
jYS3ON2kl+HxC7Y+5P8ZUyr4NJ94t+4XT3qSInnXSKE1p1/QONkjTH4sRQV4KZjS0rcVS61ZHDEi
3fw3t6wl7LQoqW0PLMlJtEhyZ1lj2DxgTt4rszPuGNPdxlMrPh1TP34oJW0XQrQg+4rzCHhjLwpT
Y7eydbX5m4/eBUph86NSvHjYmSgS/Z//gaLvrvxrMbi88nvAL/gVi4VNGUoAeqX783X0HCsL5y1/
JeqKTKym5UcxphhwH3tNwDaPBu8RFkqQ/KJscE3hM+God/vK0SrRXyn8E45RGTWYrB8zqFFhkbV6
kek3N8wIfb26DZMDc6jnBzsH1Ws8AwtbVOts1p4vjwvVvKkSPbTYVYe6ERKMEhRZ4fSlOq7YmIqf
wQ339VZO6ZFggt66SXKqrBD0i8xVQ4XyyjUBia2D59eymnQETov1NqoTi7qaeb2yZ/BiMH1YLhgj
B2l04n/Bi5ZG7D1noJf/vqL+caJaa3Lj1kHG9beBf32OW8e4X+HJHlDSxC8vMvexsQsEgQRX0mRe
aHDM/B4nnsSoFo9pMflXCgVAs0/xHasFFDtByT/1Ab7DSJzw+S4gp4Od6VgAtTlGi/pc7UQlXjvh
NzKU4hYaP/lW+c9Bl18n76sgVVN5wFyUPWjLRYDGYovTBXp3h3ZBWW6LT7rslt8DojA4oOVPAgrJ
liB2WUY/y2i6qrF/l9m8d1ydKbx43mtxyDrWseRuZU2snclZlZJBk0uoJ5cUyrmxuuOk9SPAtiN5
1z6H2Rz9dk5j06/c4n8Fm0QtNAks6uQrNxDQoYAbpP9l0M6GgL1jzOTse/qEfALwHLVUiCd/WBSc
E+X32iNT0ethhihEFCQUp4/s5knusjUPaCtt2VMi8Kw3WeXjj4z6kAnogCatyFIR2PfR3TSmz88I
qqPJEfN4sPNbd3mh4+uKjXwQcyMMY+ZWye5z0wrARE1QqueSPpoIfjAZwmAciT09H5TCgmn1PI99
5zXXs3u/kgM3qXR3u7Q+NT+r6I6uipvqCB/mHkzA7+qp/d9Ysj8Bdg/4AGbqyhP6oaohez8YoND/
BDL4l9gSQUVXnr0+i9RfziJMIoShsela9COn9FX5xoK8oVcNascxqREg5XLDCWCkynkfe/xT5snO
LpmI6ynRjfrjmqnP1SaQJj97ckHZqtU9Y3tNUHOJi83msO227Sko5UyppkYo+3livAKznC4s+fta
2tsBCSCEUSG0lEynxxECcg2uh3KJcp9b7C9odjky19C4pysHnmkGQWhK5m7hoihCc5SHZgqC0rrL
HTgZmDvfFyZBcL0qzCc35l/hZQcoMddOB1efK5JxcD5Q+eA7OZYC4gC0sB7Svs23bQyb2K6x+kDN
Vvjq0eaRhRK8nSrC2oDpxdU6A/41kCHt32qxLsDyRECklVW8zlM1Izpc45+C5sVyzaxqMqRcBEyl
7Z1ao9eO0dYc+GEeYI7LBHEuQUw53NHwQnsJmmOukOk7sN0WrHykV0vVpkMgU9DrxYgaUTpeIEGr
Fa5ygH5bPyKfULHulfX8sjgz/imBACKB0JwtEf075i4hvlv2HLZAriFrhc9IyfbvOebpKr3w7d2p
TAe11OSBOaByHYAjFFpwG6633/ROV4IwwOG7If5p+8ZdXVQ8CtClRfB1drZpOVjsxz5pzltA5ogw
lNz4Aa1GLsE4Y7H0jYSiXafUoMyUHJti1677OjUsi80EKBFmbYHdM2xmpEGyAKE6l1RqxJytEDUr
R4T02xbBEFRay28nCgTc2R8EfQkZajUWz6miZRBHITpmwOhFLTEoxAF+44RFzxgYyUskFaMh9iJD
2AH3AzRuAkMHHHVj6LeKdEgoNN4ESvgmD/5hvNTr3Mx53SU5L2LMGgQ8hmdKdx0Cw2ZFTkX3lGkF
bhaLjOzOrzz9QqR9h+jSPmKRtgWoD/oPsw4cqkG5g2OuUGOaJufnSbUYGvTca4NEU904pAAdNLnT
Cc1SxXedhe44WrxWu3TqumA8LIlJNdFjanMCSYJ0clwhQ8HIsmtosV6bbokJ3Dsy6jB+/ZTZ2nup
74+JM8nwDW9JxJIkAO8S72X9twpi4fTDojwyI+ONowFBsPozIrsYBy9SlBkcZyMKPdpUkMTEib2/
1RigwNanbs+aUws32Ktk4k1IkmjTzLx08iosX9EmeafbCM1RBzH6W+yGBrrEn7F1VJMEsorYHEHX
Ccgg7we5J8d88IbJLza/zAypUXf16+1yLz8/dGkVJ1gRbqoHamopjjtPYvL+uvnG2RqlWa972ncn
Q5BF+2zljKCtBeDKUOLC+kA9MfjXPM25mtGt5cdOYltZNXydvjH8OZ++jgYJgVRKaxfnyZfJGSrq
nBw2k80IaqA72zUEN22dA5y2gIG8FdblDr5doriaNMV9i52BH/FQz/+zwdCvdKlNq3sc4/Ay9+Jh
esYcN0oufz/ztM0EsgUDmwxWkD9/DmJgVkTR8X/7n0gEICbq2CHii49/N0RMNt/g5OR/TLYaKiI1
91kCVqmjMK8yfZCdH0MZK7DOEyYcbBLikSF7vuRK/m2D6j6TFzKaO2smlBqHZ6lJfd1hYMWTinxW
X93V+iyOnjA3l4u/OEMoxgNe6ZDqBLdxPdJGmw8sl1RgaVXpCFM0mIl0JwIq8LcLr98IKLBOsfaq
UK2VRK5DQjwU3wTVCPixVC1M1W2IWNG+Ck4YXuEOqSMe4ee5RRYustqT5y8K2TkqLdPukqHEWyMY
BCEYFq6703GTHksDau65Sn7DGT0N18oIK7Gv/UpzP91ATp04eN9AeB2FGNX9AGx4cN6GzBxsfv9Z
/luEQkp5qYghlZZAeOE6UZ73GZe8BhSFB5D8b0oD959ecbMAvAkhZN0jGxzsfil0pEX67UMgnLnt
FoQzhjNmJIatrxhz9bdqCKcLzAAPAehlIVhiVujWzwVUIJ8M+gygjN42XqhGFMh5Z7xq8iZTjboI
LgwGer5Hj+hDsOkDx4c+D6O+Tq27qHlAGmJNhCM7+SRiyK3vYGxMRVpOOHJTflO+hpmFYqPrvQFn
HSjSn0GcelQF3p/oTMfN74PvB+rHORRZwWVtt57VVBlUZcND9Yw1TvBCjBawIzXGIzBZT934AyOb
AyekXmWHg9UM2ocXqov6oXyY975v+LoD1w1H79DAmJdqJkpOTz85Bv/xvhiDI51wsjR7im3WdAQD
Ev9IUS9rUT9wm8jX2U3YJuKhYjkyQvZHVCaeK3IZ15QVJ3hvpNxVCnvc/+lV39sQg2SuTd86Gh6M
xPldkltFAN0u/JW7AJY5fNRagRkUtSDX6qaxvQx310RObIgTBplL+Xwq+bX4L/20mbeWIEqTwXE4
X4a4dUgnhPpyx6lbJGbYvlY+QBvnYk/WukHb20wdwSLKKplXbwwXTES2sitXEAwvEyxZU6hscM4H
hpHK6WowZyvTrlZCaGlD3BvDwrhAUXS3XQZrBlNmmqVDnCpJOctoGAYDXdiWg19kM7RfN8N7ECtr
35rWikwsT6AVCJY9MCK3s/MCuI5fhZPXKIlcw+dUAVpI0oecBsgzic23pesMcpTdX/ydrnZpynxy
2M5+6f7py3Uidiy2Tux1OT6Ivox4GiWN7XXx3Ewl0tN9oPJbrm7wAd/kkTOJlFT9rlu18yypnwDq
671IXLo6viqz8sz4kIJhI3YRrUCgu3Ip8q92TsrgM16NI3BOMeR8XCpKQOK42iM+TO6UaETpN/Xo
m6K9joEZYmRrvnxGsvmJq5vFFRLycHVbw8SW3146ZIo2mxp9I/6rdILu2nmCTmu0BGhRcJU/EB/M
JTmKcTl8CwgXXoCiyzmRgSQHPQbMhPyXyz4ecvNUwE0rmgOLAWh/OC7P3AxXZc4Ld2jTHestmQBW
HbLYrj7BVaho+vu/eyl1QaNslMRWR51j/P8OCp+JRvrKZjDm3WBlVSO91Kif6ll1iT8eh8DWMvxF
uIvCB3L7MMWxLfYZflK/HeG07Bf2FIylHWxYteUKFMXsaSDavuDfmZd0xlYMIkrH/QEAU4ofnt/F
xaqlEWhdYvu4DqabRTk3hBo8+y42xUHOTfg2T5oQqlampI5ixChBdFbO+VtPVN8awhqbrUCxXrm3
B1PGrUf/VOyNOnTHUC9wCxYZKcSv/BGjMkoiV5gUq8egz3oh8aVj4ayDZXHbSYukVnz4Irjdopaj
IOXa1I93+7MLGvDwLL8QrtdgsTg2sF24WtX0Ivp9yrPi9sqdK8V2s3uD6LXahY75aRye4925YDvy
x5KZ5QwSuJKrJKcCYP57LAfrOu3/T7DHgNsE9HsvSxIrrbQe/DiLfOE5AYoRnariV81OUws6oJuQ
Akrua70J0wa+5A230r7847jragluldYRTqfq5oFMlc1cRfde3zPPcbTTscX2ifcyrozV3okhraKc
m5RSuYyrlGklurpGUFFGOfFAUWIUJIXG02hyp9jE80EtKg9LsU+clDogH+CJa/hmw5iVDEIzIr62
6Z2psQsJzQHH6N3D/nMpO5W42bHc34oRFn1yfTYAUB122oBurR7mTVit6Sl4rNtIA4PWiCHkhPP1
tEw1NVG0v+U919mNO+cVUAfITWnzxgv2vkap/fDpCgF2GgqgNmPjZzgrWr9leI8lEW0saRiNPscx
lCDlfTnNrWdTZDRRz68nFKuM/JYowiYpscaLDKVgDzv/moB6nJOAk8Yc1LT55THFdv1GCpxK/Yab
uPWV4xceIMtfTQu+meyku+YEBHpVqFTgp9ebW6ePe25ObxM0lkAD9LBjdB4JTiS7uAKM/RHVdYvG
/kecEEY1lKEES1p4YwHq0R6CU3d0Hq3a2SRKAupils8nJbRyGHYHZ4fiQJimMhur7+hPAMrrfjK2
155xsovRG+HtCUUbbjvGjuOzuvIj4JNt+CbiKqTn9R9Ogpu2AYoKeXE+svQ8RMCkeGJ0ai08PcT/
f87eWCtvTNialWYZIlfP89BMpyJBotCqPH2gOVMJpLLBrOILxFwQ06FNGP3Xs8lnFHqgCDBm529H
oP5LCjDqfFczztokfXqYIy/PhWKbhqK3l2Nb2RePHGFK9O0HiGPKrgddBziyTupcHX2UZF+poSuC
VxpSRVqrxjoLwT9M20ziewCpr9WAUPw7LaUuKrC9EiBZy7GTki1YIYMYb4YQbSoeSgCZ67jBxcFE
KESerYF+GpKPjlXNFcMW3trPDRki47ic08V3dWp8qCN+bwumFEmSgVj50OS2gDX54+1OaT/zhQMs
Cl0CP5ZgCoZmaZes+HH46OUfJQ5mqCs6IehnWhxnvfENBPOH4M2JazGSOjzSiCoQBRwfbRsJ409X
d+WGUqd7S4UgLkdTlsiXkpwktliewLLLpfm3M0UXwgDfoT2ywB+e+DWfJVMEa1uXQWRhFEPYsMU5
YAHZ7/zASQZpTGhX+Y5YkJm/rj9YRTsXQmSg4OH9NDdwZ1LPrnJaLrVtcbrf4Svxbkj4HtXlUzDR
81U0gIeUWxahq2buwmdPd4YJVu73ETNGL2CHRQOvIrUKz7HFO5Wr0SOl7obSu8YT1GQBvN0hQRib
+8Hx79CgzyVM0GTRBa13BEA8pKt8+9rLkl8n/7r8XBiBEA4oHwr86d2X4vG2Rf5Ps0mTCeca5Gyl
OT/ql3JSNtxps6BEmLgM1yd0eG+3nD6mabFRrq57GVBNrsNYkm3POTEhMnXhJRkTT4XUXLe0vb0O
VOHJ+6DMXh3p0QTbXal/8G05OTXaDzJax9fNPnt0VA4bFFtEbUiCrP02ki2srwTaWtHo07tQ0hoH
WEU+PHdV8iHe2HRf12bln3LTv0OYJOiWzR+DVG5h+4RoyYo59NhmWktgr1mylFzbD9wCgWfPtUE1
YDxEkgJJxNr/9CddS4+W2iV3mnyHXQykzWacQziFVxOKRiAh7cv+ifVCVvhXjmn23X3DfDEGEHYF
tTAMBOjGORlUGRSKY+9jzjl7m8WZCnbViOEQ0j3S8ueIvKGLomKGWbDjw+BMImfOwwqWrG0MpOyh
0rpZajcVGQ14SGcZ2of7RwhIrQUET67W+Lw5w6N92A3d7RBlUpqks/uFaPb8Jvsz7JhQIfr5E1oq
p4vax7Fwv/rtV6a8zulJH723zgMj7gbriANX2+Xeqf10gmFQhiPVYA/c4Au2GCZO+gmqWak6MXR4
f6FIHul0AlqafSDmT5ifpc9784L/dUoy4vBcrTJ94ciuSgsllzBZYKQ2ImCcI5Ro8EREnITkqpa3
z3rheozBkB6LN64pdrUs6i+an8FjpPvSstWPwtIWVv3lKA2FgNZbuLcd/533n0oe3OPdgJsxzjTi
kK2lcsxJJsfd7PSzYn3PLLVWiZlQWPI8iaBAhdnVzEimVbuNVPZNyADTHiHckvGTA8lodbXp7C70
91bUJhxURZCnI+XqxfLqg2Ai7zSM1Wg//ZiqRaj6s5+oIkftrvoyj6QtqWCTGf5gUX5uR0/3GyY5
ap+Mveg9cMDsEsM4kejJlj+hiUaffd9zgcg+x8y43jbdVhc0TEXpYTZstW+pQVLb9GwDXWST/2lm
0M+UbsL2lMCe1IulaFotjCTxQoKcZFTeicrMW0PfgDqWpcCtLy1i7TqQzFJf07o3UWlw/vX9McU6
VQAuPLm2m66uz1mcGHRK9B52x8Ps22fYDIeTIKiinhajrRSTIg3TOpBS+qVmPoPDwBWMJJkpN69c
NQOaCWXR5N5i40WVKGZAHD9pdRZE4BHb0yycBMDIOxXrAC5UdIelL0Gh5V2WgkmE1SEccxe3p8KX
xOkcEhNDmKrY9NXnZceQQ7jtAsHUJ4FNOZEID0Uz11VWenHJRx//gPGuhXr7xfZm/0Wo/cboJuFj
UZirkWMrCXCXIX6nM40fSAkuD3CvSeJFz0Pxfx79a/3RUSR+gIBylNulWIioiKaCWgzrWPBjY12L
zUIPB1lEBhNaPRSgORJ3HGhEDO+3UjOLQewuMxRXiqxYeboy07QKBgm6CxshmhwP63ZFWA1qstV7
dCf997ziEp/qzDGzd6rOS1bQdLxkaipNUY+Pu0hE1pdWbvOC1/IYr5P7eCrml2VFstJYO+AVbdVW
SXGdIUoznLhJ+mrdnT2W3NoB/JPMCh2SKtU6nB/Ifk0y2Q3S/exPd3ph/DZyWJG77TB3JSPN7Wk5
RY9kCNdV7YS1zfR4v+AGa3edMK1FigkV/v6hjxpfuJ0SlMg0f4GHXlNzdgdB1gT5LZxOzTMKSZzI
k40ZYz1nhnbKpgNUFGV0xCdd99MJvDNdiDVDEeG+j4LyvhxsPgz4xMX4Pf+PY37gkKAZAk74gY0O
gvxBMPZSOgoQup7XQdRfhcRYR1pe8CrIrcRu5TQykrG+G/e9HSBBMmkFK4kxfXAtO9bO5uEJZo70
r1cUJz0MvAu3eTHxTy/J77gMMJts/2dXQiie9efcUmnI4oJTGp6CVAN4KqAX1dWjhPunSSH8+YkH
LS3XcqDEb3Uh/w54UibKpaVbnykA4Q2tGnubAmBW4PXDtz25VOZtvp966g9mzo8q55IFQHUHYX5Z
jguq6tvz/VVidJVP5LlNhuSUIsMl6c4Z1F0E33vqv+V0uknoFUwqpI9dYg01IgwVJbrxtK1CovaI
+0OH8+vJgYaA/WUDvlZClpdzUGZm0JAZRuS2FdMgMsYcIdx+excqAIkw+c0p6lknMnEzOlFeI8qX
yvpZ7BmKTSMbH4DebS9fzGOwNMd2n3+BykwiKoijgVCbuBDlbu3vhlbD5X9bvxEmCY/fQ8RS+Air
xf2lbSTgsRRUnQqgVhkQSC0BD/xmmr+i3r0ognhkUda52NverAcoldH9hvlcFgaX6rg5ZdPgwunT
4UiZRzb96vRe1SVzsBWFusKJ3EhqxyQ8MCNPgGrZIqS0znkCmZREQYUCwh5rvrkj8LXrFA7xVDRy
qb8Tot1mB0ZhrAudqbaqUK+BFg1JmtMreS5qL78LmsAAaPmCrtodClYJO+CVnAT6wRDV7RrFOwZN
9RdeX0I+zYmlget9A6dihm+G0Zh/EWuBcZfOvOWoKkveeDGax8MMAXbcL35T8J2gWRDXU+TuC9R8
aVW2SV2gIAQzhkk/FrZQO42zSS41HEBzGW2p4HLSXy15qTJmJWQG1Ze24I09+w5ZjdYaxDhYnLkN
FDtp9NKRSGfmxuSan+LSMogRtsDy78VLrwZ2EofLaM3LOv4Z9MHOOvrLsiU9qvaMiajGLAqLI2Pf
vbqS2BZGh8olwyxYILu+vdpYLn4QsgK5nuW+G1zwneKSLegt/FmRraxEL9C972f6FPsHpSo8Zppo
HyDNZj1JA07BFj3uNNqDbPMjn83voyfw94Ypd5IH5QYReG46DIhgkdU+QScD2VkScXWocxhh7zZA
j7DNJyxxSBBO/ikKxMS7Gj1cXzN49L9Bo+pgUO40DDcxbMezGrY5hu1Btho40j3vmiRSiONaaRp0
yZN6IKEdRYLBT9miRU9QDg1/50HnWMb0Xv5kO6qTJnqd5ACPQbiQZwoIZAClFDd+p5WR5OroyapT
EbBFCGexT3oTQQiTiSKMzJWqc5Z0JO1FxJ4hNhrFljEgi+8GhPdOuEfLu6B2AP6cCtJNRo3swtXb
AcF4TnKAorsMI/e/iM6eW1rXEJ8x/uNGys1bHi1EgwuNVlXbdk/OvabGE3JQ+1S2vOdiiDS2iFzI
Uk8q6e2Wcdbjk4HfpnBEPgm5E9wxTONFp7mCswmENaltDs8AlQxt5MpU8H9+7mvtJKuUoVw3va3E
sGFf3ucDx567k2YWcwuGCoyjitCXfei+UZixDn0olZE216LaqqXMPMDV5aZXIpgxF3+snyAPqwvN
DfGLS6xYqL0gBq7ZWRUGGZ9slSgbTA4jfQF7jc8kN922CGSxC+Vnc29SierkhDMP9FO44joPwXF6
gKCZ75jBcitcT7Gxc1VTFuSo9+Xm7qmFUDRuJpXT4Trf/bS42K8CJgi7cFWNV4kB4nEBstXqoI3d
6xhnGOniXxmMcj8SQatGmivFCeTRSiFtia8IQ1m6nqLDmW5PKdl9WMLeFcAdn6JmS867RaBkOdVC
3y1jifKCg0PWCyOHBA1oUaALIEEO7kAa6zZU4UY4Juc2Prt6Izcm0/1pR7fBl7iO8hr8dmJ1GM4h
rHDdKlcSF6LYw/bSJ39q/VrPGce6jTruy49X9ZNkJDDaIOa7cBug3VMl4vdKOequ6Z+N48u9WluC
u3kAI6XW48GMRYFqxchp69ApoFGks14c4kZt7gXLEVCCNpYOhp0Q3pPQtt/YXvOoCVPy1ourIK8d
XwnYchmQKozs8ZeW+yyFLUMMHWAoOzhxnpjTLRUeRa2oXHZEOBqUuCnwGQsUivREEysSIGLYtoOT
m6UWQKWWDJNCvjz8L9jTfMrYreLxrzYQyrhej1B+gt2H0BDmLuIykeqgkcD+U4gc9qkwHAaiQ68g
OPOuUVk5aMFT5iYx8j9wvO+5lbOFXU3EyskNeHFfcgTkgaB6VGiSA/lqM6mdCIfczwg4fAWx3ZKi
9e+8sWIgbS32WrD+We1MssR4Wx6hYU+BA3iBLs6qETHMpwhCc2VXDN/mYU3wLpGQ5o+kgk+xR1ms
ZdH41+y6gTFIkkjr/TIuG+4qmqQd/nCLQS8KAp7I05aCiH1/15CG/QmvztaIK7ZqHKcbewTEoy89
4YN20vtj+89fcV18Fe8/k/ebbkn5HLvjZByP9IEujSmP0pZCANS3e02RbhYHL+K75ksJAum/+7Ov
gIN1SxfJfEK8/xXfRw0Ii3oJrLyME+/obkVjLwagsEZ4yLHrT710M91HeTBevnPSO0PeFpxib2Vs
gopd/q+n7Bkqa+nnfEVb30ewhhuH1pp71r0Ce8WwF8P5HNTuMBNqSzKhWCEqvT8NpDOaO3vZFLu2
iPgqLrN4Dp7BDODGEeZtd+h8ilM6wuD1yCD7xxr6+/tQFZQ8ayuLhzneF4L5eJpiCgb01R9qdE3T
L6XIfrC1Wl/3ofy5P5w1uJYa13E5YW8pmryUiTp/boyeAw2ZYH8OofA7TDQhhoEbJywAErdp1SSS
NULxxGOqecR3e3A1WvO9KBTzfBxkmnIYsWYzdjPF7sMBI4XJzPjrcBqDXwMXa+Cyv41fG0xKiQX6
kEduZl+9fdN0tmowK3dFMjZumas0qCeiyDbk//fY6WLJ+h5Ncf6GiEhZR40Gx+6+mpHWVuSpUax+
ojZwDXQYs8jdAggQsm3CD1dxhIjq+jqLslyaQyKcl7ICWW3vuud0KuP/vpt/vJ1tywIdYwOwI4bg
vYtn+XIF0BqOaQ7gYlkFb+dvGdZVQVpOUYwUBzsi+lOwZ8TH+ftvLJp3DhDvthySkWeIJgFaCX+P
MzwGVoXzEGkRvym5eKbSHPVkbR968Txn+0rXMinlZLOOmTv25rgV11AkYwPiDai+6pNkHYQFiuc2
OYbNNtrsXI+KvAWO9X/+VlW56COQQBIErZ1GEyCwMHAtBHIOnMKC8gM0aCT5v4wHW7ig9D9Ynsic
hKVn8a+LYlda27RT1qLJGH4x6kUKiJplqRCQDsbcnCGMXptuAPG9ilFAHVkZapau+4sXhlFMY2Va
dfGKpEL456p2NuaZNFcGmJwS3P+0So5c7wiEOyzO1/fOx0PmgEP4ZF+27N8+52UelyCpODA/75/J
Cc21qpn6GVMhGdxOkX8NvkQ867uYOvlu2ZTEXnWuCeL7u+XV5JJHTZus1qrzFv1sDGSOKwouXFXt
I2cZUSjIldbfGTDkDoiZyHy/Q5g6QYuIz1BnxGPGJVmV9i5WIUwXseyHD5+1MU9CLtuNQ6rHdUjN
eUBIVshxfTh+AMd3wxRuyQ63CxoXCliWMwmKliYtWVdPhTmEsA2yR0DM4UdjlWaDIr4x+NGnHxKY
flzNJj5x9zB0OiRUTOzT5SyOnQzJhqrFtBMoZZtTUKBXhmAhuIM4svBq6qkDsiVp3a+p5p6VEgCW
zoFtEkWj5q5F3HJOKTW1ROBMpAJ3nTDAlv7//NOcDLH/CWObyP5vkpjlG7qmnayY0K2cFgfTx/x1
4V4IxT0A3dmwqIYkomWzdsDYmrCXDzNMajRb4l845F9ugxqMzaPSDfVOP9lpGR0FSgN6QR/znPBk
HqsY96nBOUciavbkwfXUMN2hkWrT9ReR9jtgbIatp3xFGbH2asV1kg9B+X5gAYD8lW3xwBSRREkt
HJrkF0rMZHBI0DRiIQEt6SebELs+jQki+jaip1jypnbV078Ox8Pjuk0wzwHiKVTD8oGfEz523HtV
8eFwYQ1KsclZhUWwB0qogO7s2Gp7sYEyAW2csER/eCYayQ/zNaPE4RM+E4IDNMOeXQGf/s20E6pj
lz0IMRFqs5oDbWvuMPL6EahJnBAtm0uZijV8lnt+Z/2Ww0OHjejNpGpRUTfTQ0VjZ/05xsYdDqjU
teIrFspfimq/xCt+WC+kk4yHFlnucqHj/VX9tfmFTIjDhkynZpge5DUHZLxz9NLduZwaDG+eisot
+rQxvdFTgtsiu/LhqgTe6mljBmNRnO8GflL8u8zJkfC6SgFgbyrvYcjJurU1K9SXg5qc1LJrce+6
dMdYvnEnLUA89SAy1PRRankUPnXaWjnJFnB6i79rOo607N7aV8o2MWuksIeJ58bNTFhvu5s1x+Fp
nU2ik0vv4vLLR5A86HuaFzsMTrM8uHpqsMCMWgJSSbnOrjKS5nOi43agKj/qHt3TtvRi3CnyX+hM
62KGZCXtW7O2VTlhY1ujQSv+QTBSKE87Jy04ZG2Ov0DsN2BXnBdu/rghVxMcJQCEm3Hls7nzbEIt
S8e1z9vEoa0tCqd/CT3a8+NYPn9ms9MMEWtiyM9yztLrF/NcauX1D1scNA/uUU0xSySlALEYfExZ
i50CM0w22/3Ja6fPWl3VW2q5q9wUAcwJ8NECFR1GXhHZcvATVRpTI/veUUyVQnLFOXxe9mSL+CSy
CXSyAvn7VrrECMTRoKZCg1kBEPrfa9hQgxtvFdQhSep7cSncimXoTEooEt+TETAZkJBjjK9cK2Ct
KvuciJSP4EFruEV/M5hxmIFKQ7fcCu/ElcbABeGyGJ+OBqsAf8bY6rzmbvJKuzuYA67up0oTJain
Lp/mdj6DAXi4sRfYmajvj8xYBJIZYnEe4mtAcA5ZBWg2vh3CHdvn6LbaI1kOx2Nan/NoWO1HrNil
IzOfqsxdLgim2lKLiHOax3X4cyVxFqkUyFSYsNFFWKEv4UcFt5/bbIhZfIgTDJQJW9T8OxognGp0
MB+57x8cchKoHpJFQO+fKHnNY/3vykS5h17o4djfYRY8NmK9Ey+1b9ogPx0k+4hEMNI9erZcDg7E
XUgaFdL/NCe8XKIv45O8ChpiAlcYzUhIJgFQC0udCwMAnt6p3Wfb99Zq7gcXNHLIwgegoOR0tnAD
kStD4EleXXJpTAfzHVceCFGS2kSvJko454OvNlBZc2v3noBMyaKcJiAPeXqa0lcxrQt0JDo0ZC5u
3l8XWlvO4IzkuU1nrJyQ29jkb7N0RJuMMJAYZIe1kVC9RqQm4D65x1VH8KtJs4u0TceybU36syge
6qYE7TqmAPX9oD9ck38B4PJgfLHNCrATjSLa1dlmd6n/D5I0K61m52upKVmOzsMhpTkhMQeTmekb
y0H9sfV6WGlPfzo89knaCkK9J5/bXOkR4Bn3UX62NwIOUt6P99MHVjrgwtXoZgD5vlZA4CIaXYnU
UlaBRBmDHqZVPCweQtRsQxmlJCmo5CNp1zY9azKDnYQNCWfsXvpcQA6fdXTgVrQqzpexDZHkbgZD
zwS6bnp7RbGapEgTOO3L17lQuRcHCm9Fft5fDmjIjDe9pDgaHvtpR7drLzkfqkcOb75rsdzuh0oX
+hpZA6BAz/RDJhR+SUXw7z3o777Kc17bl3YHLG0K2LWdLt5cWwa3IBzE6L9qZoUlOHQTGCjMo4aj
Jil/LK0QtcQpZu1PmK2zQatLld5UTnQV2vQJGWNUKly2MRRwEd32VsnyGg7wgXEPT65v2BZ7QJsv
T/HG3EqAqL1+3IRPtM1xm1rgxGUXVzZHuK3zV38cz4CZcjaYTTqOIHOc4O6HB4Ir4L2thYnh34x6
ICvRTf4KJk41oAeMngKGclE2B1L+lwmAqzKYq8H5wQ+n0WLce3jsomrQHYYaDUZ9kVNj72/KJ6CX
rAqabICHcxeeV1iaVha5u15Clhu/U11K+eCJtXP2dreAigDBKrN+anRR1rixmVm6qfQbciVFMjCu
gBxqCAJuzOUTL1Hu0fRk6UkjjHHMLMyCuVP5Z84LLhts22FZ36J2VQsJ3s6C/o7Xzq9RCui7k5CQ
5PFBT6+aAwjmBUWq0DxVGySpJRPQMlUnX0HnmRp5CRqSACbfz8z/5aHmU74TuTmdCNd9M00lfpe6
/Lph3JnfrsFXYPeRzBFsrrNE2OCBG9czgt0vqZhPEzElyWdvCtBIHxdgFYO6lZLnHPt9IMTmD3uS
/n6urihElXDoweKIQIdwe2eQYx7393yoTy7au673Wzg36CnZdGvyesAsqvFL/9A0DdQs3eeqgUCe
TbDrr0I3hLwkTK/jRlIXQ6opZHtzFNicGfYhNianvhN3EuJCZxbw+CNs3AZeEPgiPn1j742ydwDW
NHdUC+lhzHjkTrDFm8PyNhbttllunnA+za/kUL6vm2KHQvYmGPjRIAQO/f0MEK2MXB5QLW4F+lS/
MJGnjpZiYhIPY6sAYQ9r8Ab/8Vg+B0NKyZIt/+lyxwEc+Ad+ispOl1IopPw54CzCAcgl9lQsRiGA
3fgiULI8AboMPnSZrE8gBrM+JvzMSEsLKnKKfEm/Xzimrq3tvyL6BWGIO9Dz8sN2E7YzSzuHf0Yt
TOf2dxy5fK+zS/BMABl707UhRdw+yIiLmvIgQixmUBUaCgi2trar6CSDU2g488j7m29Ej5Y7k05c
dkv6VKDrlHHD4+R14Ht96TSZDUvINJVcxw2ZjAiIteGntZW35U2yuSClCDDpaaYCpLEN8An+r1R9
rP8vRJ0xm1vcu9cahB/7DiOEW8ceMNWPxMhNZxTGmCbCtVIxiUWO6Lb2Zk9ZSE1UKoI6etieT8xF
rVYlIFiYnq7+P0a8IWvmMUUAUBpf2+R+8YRY+JPNQzsmTBAb/Zf1ykeenaZY73Eam+9Mb3osGnvW
cln1UjbpDWtlSdQ3nmxnc9HJ9arxiZt6+agtkS0GdQj0jHwI+S74etcR/ak8ngdZZuybU3bWFiI5
iS13WMYUtvLEDTiN7xeqaSHUFf0c0ftDnh0a3/YE3D3LFDEgzEP//g9ZWmIHX8u7bOXsxsaKHJq5
nFX0fMbwkH6Cw3A58bHNQFtHisHC4PVOetoawvPqQbWD8V4cTnV3RR+hTvijcpxFogwomaU+COSn
Kq7iqrACqEGVBS14KEGoPo5FlsBt4C/55IAsRKtOb6ln51K6kd/GQbEgXNAAtKijHRqbpfx4JVod
PN6vVTCzIaKbI5nuk7J/G0/+ONiX/R6YAeOTfun5YRA8wVIlpk+u+NKiDrwqqDgkBG7TlwaOe8bi
EGgHyB8TinNskGT/eZBMv9xkiBSd6i/G/XXqAyCofp+UujZwbzBZV/Ci2oOrYCbDR66+3wjcd6kE
UmFSIvlSpX2tDXePK1N9qs94H9q5Diz+DTS+35rzpGtJS2sT3E3rEXswE+9AwKDTHpqF6yakgZJR
6+NyTVcSfr8dCGQAtH/rJ6VRWULPjHyaacqH/UZaGJJCsk6jQRNx65bQFti0Wi9REcWjdTGBsx45
kDjDXGAZQ+XbI6N79FUn5qQFuOziFYuDNIrcZEn9NNOdo949c0rms0+6yMy6SmvrxDMD+U2xKMi5
MvByyv3CbynTVlnuQIe1Y9fg53zhBdugJqL1fDQlQFWFNRsFmrkoS7lxwhyOtlB0YeXIVfeAaFda
IHyeqOPl1RWNCaxVGuSM7Jf4TqZoqujkUJs4Is9fPGn5MdttEzIVJwcI/Gf8JVAibzMY3LVUrClS
iPyCpeb3qq3hal7Tw85VlZ5IGx5e1UDyWNLLOshdexTptLce7kVK5Jysj7PlQdD+Fe9lql+Pb3Lr
Gef0Ia30JzXoXj+Rx04cGz71hj89d1yUCqn5kgXlk2NjokXmxC2FuEJLee/hLRSzFauFNquxtk8t
YuHq4BCR+bNn3klnmJXSXx9uAklUUbMwqrxZsaMZBvbK4Z7+4smNA4sdASi5V0EDlkF1qQTtU5zR
/G+lXYBTXFlmaETfwvL67aFTu2lPpsTuBjbO8q+llDbvUeKnAPHAhDBbrbhxFxGA3v7vNcwVX4Wl
IzI1b9bSXdv7PO+rHE9kZYoIZPHdao2W9Uh5LZ2N4ga31UehfblwxZQqkicn59rakQgl+3kpdzAd
JzbsDaw1zNn2P0aWrRUALIlYakaZkpFER8O1F0cdVaQmocXvuXhd4IktRKSNCQxKISsd/kmIejuJ
3b+wYChUL58XB93cpoHzlh5EPA4ZZ3cmxIpDoWIPQJYTaTPr3waEJ3/HaqrdV1oiNpsp+tW6H/lF
9DC1BQWpYGacUJDkcbdKs0oDh0k+sdapdR5ElPuq+jNZ33PZWJGOQfd3m55bc7ncegwN6XVmAgqX
E4ePaWyDu+yyw+WesBrJViHxWx2Dl2NLBco684mzVM96qR2oOGSbTXhwAI9axlQJpKbQwYhQau3P
2iTs9FmxKU5opm5ekDVfim6+Z19AtQQPOE0KqAh22IMVqFKXp9lI+kxG6Ukc6q9gjXVcsp14DPIv
BLb8jPgDa/ybYYpSEBNAqY8oea3bX7YFRnzaSX9jbc2VWKCeLg0uW0ItJ5vvz3XBhiQo1GP1hlac
g0tVCWn0VlcmO+wdqBa5jruduKwXpY0CscDt3dF+JNmY5UG+dPSsd76mr/W/tKxqn390zU6pIfnR
Aklt+I2aixT9/EOMOVNlaAC39DSnDcPif2qtHoBwSGXd8AwvQSn7UBcKJ+htLFQFyvBk0zKIGo2u
0WENZJS5vOTNYniV1JiZCnspge6bn9IJC9OvGIekH3mtHavrg6TcsqAozytHdEGG+MnedHTHaYVH
1UwGszIfFxjbXdtEH2ohSsYRrlYMd7oHi7zFwl5NnmOQLwJHDxKQE7ZSRmGPm7GBnP24hLiXkXnT
10gA4qO8wBM+78Oxp/KApdNllThNO5ELxI1zPnZslX9OKgzHcUtbZo5eM8Pquliz8BkCElwnTfeX
Ja44idLIJbtOSbAUNLCGJdK5FgfuEmfwOaXUg2ubyTPCM2U5mnZXo+ad87EdsU4B76EwPVHAcF9+
X/9ibkJaI4p7Kc2PWdWwBQqZhbkZtfmOmqXtrydl89AXp+6crJWIasm+5BG9g0RWDljN7DE3zMHS
axsMNDZVx2s9O71bc7s294GUKyerwjiExD4jTZ0o/zWOXY7kcbpLmRo7MovjM8aEGfg0Ssmlbzrr
IVDyvjNQsRIsgLjR84Kcmm8Z/F4INPuPI8ceX2uxwwR0MiNkjwQ0FhLYSTPMJd6ctyB2jt+WtmH3
JTb8+DUsyntFuO0zFN1cJI1AHOpnQKExC7s4bCwdBZI3aGAmZ71x+GocHzzrZL7/uTngGT4krq+9
D17ySfG3GULC+YR8OCG/OCb83ibl+L/KMuxJXEF2CGsUbvF0X1wiSe9FNCBeJ1qKrMDjAO07t8rZ
b2oBErRTT52F5Am/4JgEbt3mGirKBBoul4i9/HbRsQs24DcrZBOFed6WhqYqVQrHp3wms0uOCIyV
+yjGnVLMitPlDNz2igH6L4fPfrJsUsa1fntkrZazuvKxZGkcZ03xKIFiJZvRMpXGMGCWOGYDnyal
PrAQORfqego6we9DF/QCE+bjUXDAJ9w5j1QNSla6aWKcg/Ef6AJY/Jf/Y6lDqAzeG7DtJKkih5IV
MjAl+Vjnl9o608dav/TX2eDzFgGhgQBZSc2vQYnkZHb8ar4NF1w260Q/txae/qbs+PaddLQKfzzn
MYSdZ8nF0w/gsLyFDAQgJxYUMmbkeM5Wi3Y2sjtHHpHZCEUHGGYuiRK6XCAngVfc60gK2AoK1G7H
QdC+KroOUAIiE5uBFmwHKVcfZbNa9MCGwvKkf7ZELuQcaJlXE6WecxbF0OPa7oKbvMiG7Tz/7OpD
Z+EeaI0olFhx48jk3iEk5WU8CJjyQF0zhogi2e5EpP15R6oj94kz+t6bfz+DcgRXcOqgwOms3bm4
noKuCin3QIg8F+ByWhrY8rIt5H9m/XSxgEGbmtVfVZ1Sa9dzU6CD81qC4OPCAQfxsyAkRG4ohWQ4
zPa6CJulsCNFWl/zHUUIjFF3ViMOWlBLcb2X6kKbHUT1yidGj3HLjzDvCEL71UjFgglkvBY5DIQg
uzo8RdDw3pAe3UrgMpEcFHKULLAgKxGPgkUdc+VWrxxgzy8sf9vu1qd7pB+WN4X8sBnoRvVThJb6
sWWBCHnx91d2QGbKFsfQrUHKr3ByUcfV5I3xbZL/5tMwy8Yt9pPGDvK+gDslDw72w6xABFjzbwxN
hiQbNuyHmrY7iCML3TvCHKl43qzTg+W6wCHIWbz9IRurUYk8R9sGj5q7Pjno5MA5AHZX4vj3OLNM
pLQYrHLZQwx6BBXtQC0/Y0a4MXPQkdArGC3Xhb0l6Bg898ViI3W0abykuGB4m5795kr3M4nbVdIz
ZyAyN2eMST3JUsmXw9NZd/zHLAkY/A6P85FlN3DwMx1tNXgN5nmX6PCEKHRryxcUliSvXFsPOrpt
lNLoJuAyWviP5AgugCdjw8PeV/yz6Gsl1mJ6JPyZP76tx2vVwOAlJhzeZKnfxJ5gizfvHWnO+yv5
qVV+OpsUjLIB6CSCitdqhSIK1p9d0mZCRNfR9Jvi267Zux2nmQKRCdmLHppXamZRvj3MwQLSNTE2
YYk1lYHW0zlGC3X3E40jEr5ZPlDY7YG+/aW1tgA7WDIOrTREEkywrUm41jKrogNSTwFUZ1vu6cTV
YP5LmRrFwnYteYKjed8OHpDKTHx842D9vPTCHTnH60bbMOmCkx/Fq0wGagdG63MG+00OqD3nVnbw
tJRnMzfr8l1mdAQsA+uADXJ6ZgjYvlMb6ZN2FRSFYvIGPooRxxiVD9uxtWdp9UqNKJWXbn7OLWdW
fE3yRHK2ehf6DmLVbe4NXABklqjDW6J/j567kHAnE84NoqpMLTdIooY1aaPT/BtLqT53BL4d+sje
TYCqiAypDeE0lvc74Gkako95cgsZbil/XdC0d7AVvzDzBiAGeQsQvyvQqJHjYX9dWfJOW+741sY8
IobxCYR0DPT5JdVJUgb7i9hZ7C6i3GfdSaiRzbuO3ON30tcvnkclyY+w0D8k45cTRyUO1ob3sZS/
NJbQ8J6g+TuuFRExCsl2Zug9uRPwJIXFjgNWwY7gOHqGGJ22u/mY7E7N9GPrNBVKHZmf1DaMLfCD
ISaXqjUfSsjGo+yZoGOQvkUHI6gaKrgX5j8xZlC731hm4wOeTK1uRCBSxRCHavBH/kcsKZvTchL5
4GcFnytwv1CGe85wbhFFyzORLf2FbIw+g1L9wVXmctMyof2RwHoIA5vP+dcua5Ryevy9EMpUD5e7
hc28p0FrDZlxQhkc+bIuSfHIu7/z/3eyAoLR719tvAjYGWBm7FyA148jqUQivsBGQtf0ar3Vovll
lFlEqUNQC1bjUYKb9cgQ2S55EGts6vsxIzFNkBN2++LEwO0/53Qi29mOzH0AjJlJ3WqPzKVZC/e7
+qsElhYiWxAk/Yjv3NquTIzyOencW6Sjoy+jydaVK5IR2kwfKUWrOyLkuxNZCqQUUQN3Q11guJlw
+zmilYaXz+k1vO0XWtMOoIxYUEgSbZMFT/viLXWtcRHe1pL6tXfWIZLyBtXOeRP6FJaqZstpOVV7
SGfcGnF1gbhuDfVBG3d/4S1LSxL6nEhTcwlLWWVdjyx5C3TUqCi/VGcinv14NOP70QWIIGBOTM40
0VsSNaUxUANcfUfL2XOqyynKdM7n5Yi0vR0Sws2WuKu1DLGRqGq+ORRuVUe5jcyz5hrgffxdjRgT
qjboWp87bZx9uvSKGvryMB8iVOuA4tzthyOKi7KLWoZgQ6uTgEhCwBKUcMBVZsxoDDUQa+uZ4jgL
PxTV0QqhLUigCFr1xiGNA9vnEx2C7EHRoOMOfH/5oCBnkQkqSjfB6GQS/e6V/jhGLNwCfWWg72ad
GCxp8wEB1sqHLr23GViY6CjUS9dEbEMfDZ+TofGSB7+Y2G8aG20oRYitYrGRRJvsBhaHtKfr33xx
WChfvClnSGt+wRrBRyFbb/efBgKpYazfrhIa68N1lLqgc54XMoBQIv3mczSquncfrKltcQDenWXz
DrnztcrGHRqgbH/B02WzAipu8ea53GSlGm5ype20oaFQEy59NTu3qnnxEVdxXbefIce/wTpcEfWy
3MVmsZZvn0HNdpdEUAe0XLsu5zTjzPJbk9q54xlitjGKW2DFRiZx3wJYp11rU1t2fXFNC3q2jWUJ
3J3myH+XIZVsJCbt+2lIUe8YjPaeXS3HFDWZVdZFPos+TvZKOV4BjOT6BXDx8qI2Jp0ngHEXgsst
q7cXF2udEC696Vrd8QIw0fx8v5RYa0IqnNsxUFPSv3kMulTFY1y5K1aV5aLbyxEtyJCA83UTge+N
slREhWOrEalHxkglFfqAraz5vK9boLWs2rVYn4PahomM/6R34YvADZuvQe/qDOflGcd3pnpePU0s
VNaAfUBCFRchmm6xE3YqCgd/X0KtLS6cWJGv946xlEDBkxGapbjrI7rD6kZF0i4LsEtz3CjesUOE
qMIwPKyDlM0uULaZeU0nCbVHCU68XLF5H27np7oMPQ2NDk0rmctSNK0HuRI3kgmrquMe5vXjFN/h
NDWRkGnwEj9d5/3tlFeC6JYBCw7PsM0f+W6nt8K/KcldUd2jnKWzMAKVXAPf8FE4V8OUfGc0cPsb
bkEL9j7719HbXAEntQTNhT9Uhao9IIoWVzvkOv1WnB6/3nA1AsNtbj42Act1bB0AluwkHPSt9tuk
aLfObp50UoaFoSzMava9X2u4muuYM5YAyDi2TT6SiIBggEWOSkGBXUpdj++QTTt/BgzYOXP/mDZG
2tPDk7Rqk/8IHGVxXjkB6+dQopCsnj7bCjBnQeW94UGUskb7Q4LHaCRyv90kplYlpCL6wwGqtYlE
eXPB7qAa1d7snZpURRF0bVHXjhHOMbD+tSIe+//41UJSWWE/GW1d7ig+3aJB4A5vZEnvKd8oixd5
DOpuhcJ2Idgtw8erCdcZ70hFnbiYZ1t2ZdhaT9WyzpWA34W8GdJE5C48xONKYct+Tr91QMU3FQrH
G5oNVmH16OsgEOezT65iYVm6ThccYOCDKjGLIDEEiuGjDqWBPL9fcA+zUvcsdCwaAl3TousW1Oll
cXQ1d2DgOrpOz/HTzElWgnvx3QyRFTyyT+uB3RxTEEuh5xw8ysmxGJ4Jfz7QJUJsmasB4VGSNbqs
qW4v4YaW8JRC5rnz8zBtYUoxpSXxR3gvv1QntALOtSZCPpgTlEAgEDXvWwVNtddAGwrK082HafhF
G/maI0b1CzbAjsiSept7xowkZbBmdFCboIPK7ABZHQabAeO5uCjaZ8d+bozeiVID9MZ1M31hCYex
tYbInoJnp1eLv/ltr0lqJQcqcqqFExURT5XCwOO3NVlTg42Vyg51LFC9KvF2mLzGDGIkOu6/a2uG
Tni0oFhHdOn9U76mDlS4Jgfs/96eu3OGK+Spf/ICom0B+c71n0BdkpLiyAA35u2iqkQnlB/nF0ZT
s47l3lhp2ht5xUpm8myrdEYcpM7D+RptYmMQxBtu7OgTQUViF2tofFeH+3DpQb6FExX1qhQB6ZgS
DSGOgJIN2Qx18rpNgr37at3UzeW8YWVHw1QpSNAC/NRHYIZlp5nHFQ5e1h2+92zEJPcD6zCsd2mc
YvXRHRz14vufJwnx8ejufampb+KRfHoiAzQqWHj84ldWWrPP7ctbXsn4hoDJV7FTACk/NJR2ppPj
Mcdvlo814hDoJtA9qwQARCsoljf9dqWLI206J7e8YVAfLJ8qEmneFHigzWI+0nH7HdYR+ONml289
FLJk+D6Y3+syFXGUAOqaPjaIJv3yCwugMvJTGvNiE2necKmrJVVIJqfhJYMrmcAIqfO2VhXc2ag4
FCcWoV6eov2Q+Poo9AwBcKpmEO7HDInETj3isf0Tcrh0ARue2ne0+txHbQXemTuOZ2vjx8Sp9yP/
y0vZOo0yb7gyAOIPaZVrm7snYCOqFha892F1NS6YmyAAQv0t3lh9vUFZNqFGpy9FQZeR6HD1w1x8
saBAN84JvozDzl5nlo7tmhsPu6cveV5wR+e6B7porGdBgVoq6ZRrfJasIilGOIMwvBaRdp8F3MW4
4Ul6zryWPoKbxMVPalIkWNDwX1RjXErZPdmyXI//RvLVbbeynq6D3Ll13SfVDkO3NiKCZ8vceTLD
LX6P5ixESQ3oJCP0lvSYpfDm8yYUNIUYLkLqL0x4YU6PLqBtoxSH3RQdVtiQ+fXk71m2GgYszipR
yYPwWY8ZEvuv25m0vhU6fLH8Ullu2ctYzVd65cLdkh3pOZCPE84ifk7aMXRWk9A/1//hux6DfLVI
UwxPozGz54RqUWG7RDEhOx2+onZNCv9jQrQi2IPgaxmwu2txlp88Z1uwN7kk4foM+gnxcoMDKNo2
2JcP1uqrVpJuCxpMK09yUpSY69pJJrFkLdTKQujjsnsMPtbBqOiLXHF27lIvLBQ4cm9XHKz4LvH+
1BxAcunc25gy2huLNZW9NcpRn9lpPyNS4hyXpO5tQ+S0GRxJdXTb6pqc/jBUZdtxgaMTZhsurv39
2nTtByISjUBVJOtGx+Kxj2aPc6DpXD9QkdZbqftz7qY6amI7v3hSXBj6tR29vxCyunyvmPGrVHZ8
PX1aIQIMABeW1pP+pDyldJh8CHBwZ9JrHBnoGVdn/uxiQ4vCz86A0OTvQ7p5I40peMAoDBzUq2z/
ALFdLFeszcTjHyyGlnOO6+f6AAZByAALrKXp975mVTum22gdrLff5wVaJ+Tv43+4FRzwYoBf7iok
buoN0wa8VqcjY8QfkJyW45236ZLMwOGRTNg1fD6HGYFMT9VlgTOKQiqQMBF8LnXBvNR7bUorJCw5
632IUw4XQmfwyja2HHN0HTJen8ufxJ0IgUfUMi9Ulz5i46XvVW0io9AsuWaq+90fvKJePdQgGrvf
mB3H41CtMwilkGCgMES60N7howzRyTCjK8MuE5ArgmZX7XNodxaeCtQKZRN8XUOUo8YAQiUbE2IT
sVRD8ILzOa/X17SGWbaJtMFtoq14T+16UOI6SkRbYbbs9yVF52Mv8MuEdRqeDfrSTMyR4cFWShIS
aDJorXm36Ld3MaOUYgbMi6q9FiWCh38Cqr3UMlx3s9aeWn2otTfttufzI6WlUsxR1wy0i6XnNa4r
AFLTxbMtAuveJfphGHoJHPQj0CVPSBlPTmNl+jii2CiTapSVsjH+PLizo3i9DSE8hzDH3HrGMQCa
Yl/AHGZKMxDtxHY2Pj9N2pVhmty5yxrGaC5/ImwG1EZgk6dLwtUb7NoRGlySZWy8sGDms+3qqaVk
M1nnIAE/w1qs7CWWpz6tkKKG3xmwAdOcCX+nwNQq5K+irYDH2sX7SGtiXSRdkulQsAGdKRzT5DWk
rg0wrisbMmnnN+hC5Kewya8gmDWerWpfDoVbiiZzp2C74fw77noyMc6URIBOU4+omIivO5GsuDA/
niejPSCMkf6dLYJZyUciC4BvqpRnnPSuZITOZ3OSrXEPo5x+nGAqxQfkXpvPsWHLkYg834OL/Cpn
vosc/2INT5Po22rKXRp97FLINXis5CyjveDXuiW+1je4oybkqOxE49Kw9rOFmCbL6KjemJV7Jz6t
bn5I6OQDioIpTEcsezeMM6KsX/VQUelsoNToLHR7D7sR6fGOBNVbf7BCjchJqmiyRdBFs0DcfLeH
FBWA3Wcuao1oA1ZAzc43XupTZY6U6cf84xIaVY6rtZeSmUb24CZAmwuLeCjvnp25aHjMoO62HYm4
lB3AINn9qg2mSUc3C2uiW2Tcnlo4IRiHD8fb4Z8kXo8Zi+4DyP9j6/+20oYiDQ3FNQjdpKBVRGhA
Ugo13n33TB8IjHubsDbwrdUjg8AaWzCbZnkVXa3N3doW8R7z4ezBmT0WlA/4OxlqzDqc32csAsWN
m1ASCtvryIpBbIiUARyfV2ygs9UU6BjcdE5Q+F+Mts+bV8mFk4DWHUaFpkVtQ1Brj1FHL7/O59Uj
3hyX5zdOy+YFUKXavd5el4lrKbVrDW4zy0rOlOMVFIZQVQfsLPtCIdlaE9ELpAkFf5HIVl0RPtj1
VHYKc2pnuH3WYfI9xi61rUigaFHs8FBW03faYI3hGBY5+ha7kl771sw0AJHxE0Ejqg2D60NU3gjc
0hNMRE6OZDKhO4/uUZg59q0knky3umKjGH5atvBGeShA6Em4/XkyOrQRAln0tanbEpDGGV/ZEjD/
qnUsCpZyuz+mijjTk3ulSzQEPnPLJmqezMHGW/CqF5TmoMB2psqQ1mDWRc+GwoyqIr0V+q9u9psp
qKblOI/mDxDjfwdzH2jotsfWPXKAIDjddBxEE/X+CC5u+htA3oIey+B+W+ojbi3zIM898NQWKWzp
eVAixlbb1kzoKDlvbcMxVgndPV6NlTh+qRCogT4uUH3N+XgNLI4IhbEPKbUD8PvD8yRgduZ4PldV
cioWTVzEvqinhsh3TqQwgYB5qROQLVKqJYhEuSTM61tIWYaLE6sbDfqeY3ET2xnK5LQDN2enLeHK
kolgrFIN0yaEyn7cI13SRHAV04vifTrHkMQwX2fYfY+yQ/0sP7JEFZF1gGDt2tWoPqnJNof2kUA/
cavQNh9qOr3TCsrBftcfIEpCfjrR7qwUVfirSAjqZAqSI3/wQRcPdlD6GFEBX5VLhy0kQ2AZRtrB
bvUHh2oRCYEUZtV1Yjw1hNJw29gs3htekXqMykAzgCa8TkM3KZCx5reUh2lnJTrfPDlCvTgiKDZB
RtzVD2MDOMTdCv1DHsymmjBJquh5TGtaZV08LaWH4Vb/Td6203wy2VG5lZJKescmZWlK1GjyCz7/
Fz+lIbx42oz3ncvwasLd2yi8g2+McRciWMSd9WwMg4R1PlS+EaEvoJYhzUc/wl9Ll3+W2gtatHMG
7nj+eT66WfcpCAuLjGzZTFBjFs9q7O2FR/kF1kOZ7QXHLfWCoiM+CqC2LJ1/uq7gPN/Hv/C4L+RJ
dGXdhQY2YN8ivEEqmqJIf2gqD9+Edk+bt3MH/gZS6yZckDQKymdeirLcffwG/UmYS4fwzlDsrG0t
Ej1ZPyb2/sgxMAp2WEu3zp18YuBUvhxLaQfTg/OKeshLglBU6q5mfqQcL9KEb3viERSuMBjUn/kP
esI9GsG8Krr5rB8lXqyEOaiyVzd/SOZS5kcJJGDXlWlxEnmN8huoTJ0Q/jxg2E0+6fE+Jw6860kt
rWm1ahlImflZtFHnhW85iFPK09Xw+pHHjajIrHpXl4gSjPD3EYY8mbuUxeqLYTZ5nfNfjbgV9Gz+
MU7GnLMv1fcHxL7gRSTkLr+jSrFLOg2trOjf70SOKtseMs3rptQTBlDSR28cQPBBWGF1zSmUoS7z
C/4tghIDZYSbsCH91OJCb0qwNbE2kG+GQfJD7aWbFEZFps0JCRT598aAdeSLU3gLBJVPPjuO3GrK
hLLGtrxWogc7brXQq08hmhzAEys9t81aIDC6Rk2edBtlKaKd5QslNx/3uW95hp8bOIo5BRFdGfET
yvqEV3Y37e4PfnQM9Yj5PVaW0mCMimf6pgNKrUgclA37SsPjNYbgDt/fz4904LGkjIs5aLGQq05B
JErvs8AK+EHVBcHiHFGjMBmtLwrdqDgSO6ssRjq+xr2slqtzeK4egKBeYqRd+eAekXqEMyLye+P0
+d3Bt6r9N0CA8ctyFqq8Y/CfNY16jIYPTzqfc+45s1LqheMKNyK5L7vHYWPqwoERNrLgOryuTis3
18pzYLNVDZbfc7z5bD7VfAdv4gfdpVC/Uu51blvnLjMGLcmLrHQQxm3InRmsddhImvXr4yZv016d
8T2Dj0aZUs3StawO4pDzqCWnhlKFBYzWqMP5hWbdKSM14VRI/LCHtEI94Luj6DHN1AX73AwXLnIl
TcTr5hWv/f0i16niZrScDzbv4GvegB5iFQAHlofoYTnA2LurZ/lfrf/+vL06zI4hGKEnSobJalq7
3nhhWtq20lsjViHXoPxSmcTd0HVrdkaQUD/Pena/AQYYDumhUlvEb22UMBjR8uVAKYztx2IEzmEM
CJ5loIBH1+HA6CQbIOAIBOzf9p92r3Ucjv1O01GCDOSe3Ka++m4oe/CYBpXMRwTmERnGxIlAM8j9
jOrhYESCUgPO0/+1oTaCv/O49LQRRwdM24dKEXegVR6R1ckIpheEU2FJr2VUoSmaybGUAeDk/ja+
2siQpB6uDy6aee3nMcPJSwzVvAu5qCtY7foQBOD6yTclb5/aVlz4U4K3REnN5SADgm5FVMOsX14R
IbfZjErPq3HAxXNMEBEBkFknNr6RdwdcjZ+8XJAjLis6+c7cdZA5r13uEY5bZ8Iss4la72d316aN
Wbo+9iMM/YvI7oI6dE5T/j4FmX0yl1IC6l6u+pK4r386ffIy61n4Z7Z8VFXDbQw2qsXp21QJSr1D
z1OZMcu0t/BoB6yCp3B8l1DVkmKuA8MRnBY8hU8YsNcfVx/fnJ8bbDGiJu0psW9MI85N2fRhqymv
mqjYJR9/iJnalTMyQ5GmHltPFo6bkGj9AhF63cI0BrH9Jf/5O0D8D5Of2I9TS9649sW4nwm5UdGH
nC9Xqm4isbs9NgwIH1pKWNHouMsBob+nJCiKUgTvjJXUDwZh2HkQXy/gNE7it+pC7LqPKjltCrML
2Sy/C3FJPA3TZxG/ToAH2hlYHBZLBIJ8Zqvq+oQkHh1UvXmtoX7cM/5nzMXG9POD9SpjqGSlmGtb
LsFlbjW2m5yozDvDh53neawqPBdbw/us6KfWokB+emxH+Frb7ox8MZJbuL/DXEc13NSyo/Mf6Egj
z3oerK8SolqUWPcqWIrjhmARgqxLtWPPYPi+FB7UDBf2BU40h9gX2QD08KrIr1vHLMwSslCRJy2J
9j2onhzULTAKhOCBKOkCp2pPui+VQxj0x6RGVW2HuRJOVaGWmawOb5BTn9FVhRlTVL53nwmA/Agt
cOuxQLFZtkKDHBpPpGCEbcJb5B5C7WQ2bkyfuBu0j7si+Mb6L1LQdAy09avgkHjG02Wnq3e4Gd53
iQBZnswRcHfHDlA2JJ4iTit6B8yQVFfQIPNDg4bHUrGDqISxYGLNNG2nBuc+Z6rXd0p6RBqwMYSv
umLtQTAAF70teEm2WFmpKGtqWB2b1TxmcuaN1JNRZo2/SgTjjcNSIHXyI5CO88qnX35rdA0JgODF
4vW+1x1QheYfGmqn8vpRdb8EHQSx1MgAW3U4mZPASqmi8qPXmnSAVClw0v1xrvyP9WyjuI7EfoPi
A49pvLDyJGPcdDAxYNs77iYJlsnuKu3KAWXA50jd4rSIOXS5f3lxRIejk4j/uVtD0NCFqmToQyEm
yY3uewXxWURukP1hVElmqkwF3bHJuOxVYsOj7I3SpEQLwI7Z/iIMUbJPss+NX3/ZUub3Zf5E0VaG
OGRwt8uDJCwADessOyTv58JJHZyQVhKCpQzAIEjpbA+BS+FkU+iJ4PmrnEDy+gjSKCstG0/Ss/B4
s4Sn3nsluTm22Y3w9fvP+Nc33Pjkrs+48wupB6zOdC2xIF6/8VHwm8A4cqErIY74E49A3UXCnyS6
Q3LkVPw4/eHdxAElKqLutzUmLP7gzswWtQG7sWA4nB3YyeZMpkiN/t6hi7ZDPyqopFzTsOcKJH3d
y4VQ8wCY0TBXtKk/vYT1ofcTDDfG/xxF9W/eCc9vIN3hRfMrDJ3AMBRS8pfBJMA1Qg+KvbRAePdS
1vG1H93wraVC9ZM/H9J0ru9xT72msTYVWTUa1m/THTQssXPExHNk7OnhwA9M+vTJgi0T6lW9bCO5
eYGZnyuTLQRo36yH4YLiNDiYu1otXN5qj+LokL4SUud4A2d+KlkJpVdwS7Es/Fa5dGLKyBANUkAn
DpWaDyKcLDOdrI7WenbFKdVyltQN36AaZfPCs4ORxOat8//OefNrYNqhPfTy7Yi2iDFI6jfBtar/
qNhtS7G5tQPwBG2ZqEda5sLHWmNMCab4+RrZDObM2PIoK8EViyvOCYcjYOnxkkuT4xgXaeFAMHjt
S+xm8YQTxmeNwsqV0coooGu8yprRUy6UwoQFo0UNz0JyUmhzAnaM+F75HkC3wtj9ktoxjan+mcJ2
EB+KLC87x4Xbr3PHlbqZr463Tn9B5CtTFMEqoNTQ0AJx3oGjtf2R/dU8a/84vq8akXUB9EVc5gBf
1R1jmat8B2FGTkU//VJ7a0l0n11162dk9xFUod8lCg3z+I5b5zbYjISQKVCMq9lWEj7hGjLhs7l4
LepTVcSxNYuZIoQjdVyGMqmW6/EIssDZq4elKQVcvP6ncRGH4uLtg4Kc6ZiF/ru8ayIzKdXRe4sL
JmAuaH2/oyr1s+Zi7btK1qo9MeQVkA9UpN4Hz1iBftAiRVME8I3atgoq/7kDv4HW4SPHWZzpNX0Z
hFiSd2n993dzTXjKeAygpRb6YnbBH7Mpjk7EeEsU0Ve4bpgge1/YzUKzuqDqtxvzdYJKlfTenLCQ
iTLZHwHO4qsRu5U/OgSUhKElfIQC1gU74rwNxco8dy1+5BgU5KXNC1sPOT00T002zFLVs7up8TeO
3W3L+gpMXkqvx1QFbT4y95r9u7BNQsd5iJp81clWpMeWay2jsf1ULyT0XkxmR5xJq9ck/ZSyRMg8
g4Hlv7jL7xPSylBe488zXqQ4tqGpLxMucHVQwc6g4O7xp4IGSl5FpuyeC8L0mH2m4LoXtobzTWku
kvVAjBW6hTQEBKq7GbsWMj1r4vquupWahO9a5YnwmKKNZRYpNXA/t1dL1C+q440t0VhWmc+LJeBw
LxweO0Sz6YpNhQKOxn+X1+1VSIYKngQONMKPsVLE/7rDyMJfkVgRQAoqXv/0O2OyhJGAf3CzueOr
mzKmzHDB/cTWlk6Yb+Pqk8ATeMwgKnHBLmSRiXS6T03h00Xrd++k1eVnvEzL4yRYWrpsTW9+dGJQ
lMYLTfUfNSX2Q/qhtlXKjWqC4sT1oSn3ARTPPy3CUTMn/EOcAiq1LkfXMNhdFvboXy8Lu2++44ju
66ht10FHU3OGfl0A0t/PQ8QzuiE46+HlDuCmrSZ80maXSg6qxHTq4IcnM98Jsjovo5i+nGWzFLo9
mXwiZcfK/PZBJM4QhaoLr9SpW47aTuKShRX+LnH7icT8N5a1q4QZ/+f2euWg85i5KFA5AQLQwPux
ocQh0SdM+IV+aHSWy76Rbh0E/827VHgqL+kKoV+ctUcNPCjtUgnNcR9d/r36Tualmv7CK74FSrN2
4yRXc9NHi+4DY/UO0Blj5aRikH//n27BDR+jDYJgAz5IwLwANwHkAU9NcGlwZF7BzWus+dfhkgO/
b9t8/L/hS3cMVjelLMFCL9LSGDBV2/qJaEdMO2kHG71u5OcFOG7OBxaUAZtmC8oljllLzfGjmMEA
2in8rxVtptQkC9lEI5rb3ff272qzJeRqrT+4cX/89fwTRfxinLyJep2Qs+OamqZEfNkXK+mmGCoU
0jfsxdogV/hYXmeb0qLKyJJhdgdKnmAPA6wU7nomTO5JbSpKUCm1qj4Pcn1oHoYLpfs62a513Tyd
RLb66kfUtd4h2Gwa2mY+ojkWNJI6ByOXPSgW63dPfR+DNmdJNwh+/3UjlftEb9nVenBfZ9z0h524
LjfJoMu+Og7J3EmHSE0Oad1Du0l/fJz7T7QOfKozZWRtJ8dPcijbe6WZ/kIUIB233BOmyQaZ/PGH
XiyiFY6KWzJkiNavqrT+mqi2OvbC8pZUkAt6h4GO9yoTysOFToyFg0SmslRmccHulkRCBr0332by
n0WtmzODCcLsON5OQfMtNh2NxlgraBYIy1Povf9+BS8N34Wuo38S8955UNYbKT/oj+/O1OufTYbV
ZC2S+1KNCMaYzkBGzYNHIohddQxYuWCnBjvl0sjSIIMj61dl8S73oDf6Yet4utpuXI9PLnrUjPkG
jCpzh6Lh6y5dUH+CLtDMN2yId9CLTHwhihjS0rwo0VVbv4p6wuwktKLsZ9dWoN5quLh17whpEbAI
UpOQD7J1LANFg3fNxVms5/sUzio1/0mgcXha9Nu0VRSQnCSNRvdUyBvtj9jTQe4rCfXUaKf2uhzi
GYFj8vB6m1JDx4aMJ1dbM4wGDURoDK5b2xzhYI6VkMTAtce0YTINuEifXL6RabuCQq9WBy38VYPs
s0mjH93LvIRmv7Midm1zv+/UXBo5Xj1rI/ezwhU3CXOglTtF1SC1xATZBVVLoQwzjVUT/D6lnFm4
C5g6xNuOJzf8lFl3RXuQ/jQiZOKJfYiIdal5dXWRZkh3l0g6fTgogdkFj1oqncFvBQ9MCGvDTjmf
Kj3Ls6mITzo1uM6xEbT7+EMIZIdUlgTS6dM52AMYSImU3lT+arsK55imGomOvQCPCG8gCFn2owLS
mDW/QqNW+uXWAYKdGXFs590u+sJ2GXY5cLTEIpFSV+5WhqYzvYjYvDNagFwJNtu/9ZrKryAJAJIi
QPD4sT2rLjgag/5I9JggRzzosGr/wIPAbbnlXgPId+nw7kjuLRzkpnjrnPJcHVTjRk4bBZCGEPub
4wvf9a7U3wz/j0UyiFanwhtgnQogOC9PqJ5EfwOPgYVXaVrp4yRAgTZHyOqNaf7U7I31rJFTJ8AU
GUlLLVX1jvCOXQPLEVf3oBu3RsfCxgNWgr5JOxYgui64sDARAkTTZ9f4G8zomW3xsJ+gsNFa0Q7Y
NMwSQS/hxiRJFmjUGgw9/6qqMmx93+hiNE6jimYyrE2xBZsYW4B1BUKftYBhT5o1N003ajUoo4Lg
WDSsI6f8E4e94owMuaohDlRyms9pvl/aqDhEPR1uRbFb/SW3AskRuWQiKe+eomTFk6Do0p4Qtvii
P1iK6QylP83RkZJ/JNOFz+5Hf5D26RFiAzN3U+MkbxZmtkMfJ/Nx+yIg73pQsEKHfOQ5hDgp/QH5
4tMNCToS0wd4vAP6mh7Js6yoIP9FmrejKQaLVkYnOaWjtNfBNuIOxGQaFPdMu8FqeXzY28oWXJUl
sQYmgiQKdDN1pS8xQHaH4sVG1C5aLktoVyUFfh2oLVrGytX/CL+2+r/j84zTcec1MIk6YldB8PhE
MA/lxtG4pOeBKEPomZH1zwU6lQOBtxqhZaW4HUcovMb0pEO5pfWY3iDk0thbR7Mcn3dW+INmLmmW
OX4UQbBfo5zfkq5Z/ZoUfr/a+DhIfNZkt+n20qKNKZsbqY0CyDjW6m+xVdOMhdgHDjPXRDHDR6Jx
fQeJqUIxlZFhcJjA80Dhpc1d/VkwLQl4EPCnCVpNXWNXsUj4uuAbKMwZ4a9ggRmfGYFlX9gh9asU
fa+xbx8olryKFtQryNk1PrNnTqy07RaTpMXykFpQEA3Q9Z7aBrhA0qbdG5OQkC91HkAPmvR6hYZb
jDBP2aZWleLZlwT+9hBJ0yMhiXAjMcI3cP5kV9xIIegWor4M8PTL/BerGyfGLH0RBSYoauJc+CzH
X38ga/lE3/8woMD7cf3NwwkJtf44W+iDe51kalxKSjxhoweBcaBazpWwzpRbhkT/TWMFgBrus1GY
Rp/mvymq+emykHBGHQXTjBsvFxWWyjqbL2txa16hLc9QJvW2xMRM61KOBpxAt86K62kGbyKsSPf9
wj0Iy0GcyMkffa9KIckkeE0n0s7xctQQQECxR3goZ3ESD79uhgtET6B5088HWOv3NQFD5sE5+mdF
6bq8+ltwLTjvv5Ml4eAbPXL90UNY6RxdjadTdFHUkxyatDF7PCY0F1HDi2eX9FEej3neTFkNL+hZ
0iFgvKxPahM/o0zaUWcyQHCm/71nL9v+duRkwJnr/vPezhOrCgkgYg3BIIz87lDzA2khqxsmX+y9
IXkQvfnyuLZdNsW2mgLATzBOH40NCdXRXVcUWUwKbq6yTI5dzxKEHx1NCOrd2AlL6dlwQgEJlaHj
QBVIAyqialE/3u6gyiU6hCN2ZscgV+h5iVFizv+CYvXgChlwGWW5lCjDpI1IP4yK13PCvUXV6gUJ
sSaE5NidftymG3R6blzW/LJ2VcZUKw2FcU83OG4Oa//niBNcdAuJ12fo4jmcDlksSc/C6iKbKd+t
VyxnBBVK/mgdxqo/eU4WIPUuNJ1s1CZIm03Lw6PiJu/ofRVOwLFE4Ob1tvNYy4O4Ojq/r4DRufJ5
E4PZLr4Z+Q9ikLglgOX45IfpAfywYcsLAlh889TO/BvdZntFmwXiYhxe8OfyV94wUaIdQZvo5M+I
+ftSA26vzLAcaWyq03POyVL2NKiETfl7aC+BItV3nMT4vP47fB+9KVG9+Nt0MoDkQ/HguecSx3Be
PNr6bYhj0kXhu5kjiFmJljTmcIYWJfZ3AoDmT4bskMkRoPWWRfHpucfQWV7vhW7IP0vbINr5rabR
BwPGCKWa/dYcjQHLuqDzoud5DlHSirda0US1vLPtPhrHJU9YIHgrcU15Y8KcySVUUFhSZaj9Woss
vn/rBnbuR6BfLC1t/Az+S5yeMbno3GvUWt/+4/C+JobMvknFJMeZiHQSZf/fnKKyFbkMTG8TD8Kv
ax8pDMaZ3cYtPegysMUJ2Ct5OYREAeKawYOzVzus8h17nK2wu0opZbexru00gDJ1u9qhGLmam8eB
0TqMwr9bPgjMQaTF+DLeCwfpxNqTRf0rgbeyuEdh9m5lWJM9wMmhXHsuKRhF8EclZdx8rQVvaacE
h/ZaRLaS6mBE3HY5c4wkXI+ekGTBwQFB5xb8z2Vfx24X/TCkM6e6YQpu/TKLHA4JrMyGGMy9JwdT
FLovQESGOmrTAhY6wqhyKCRdHgW+kdJTwpl1TDUrOIF5ywn7/UvUkHLjogzgfcSlOvXVnp10/eEq
uC0MpedGmrMLINpU+taloBxklLNzm/bXTowqV+J4MsgbmXJeMDiJGGLt4EL/zN312Km8KGot7PvJ
ukqzsJOUphykZ1DiRw9eC+sBpZgGWpVjB5HE4iGl1ur6lZj77EEzzF0T0L+0Ftdyem/tY4IsgptU
+0IAMKDhvdSHrx9c4y+upKrEbexXnzeQwmbg6DuovZXu6++Yy/s5z5Zsal/rdF7EL83zFjfVqymD
67E2iz292ic9fAAhRiYojx29qj0WnOf6AppSqTNXj3twOCXKX05UEaowGFfAMENBfVclZMwttAYc
rugDXrShFMDoCZO2uiAypqBxO0gy0BzBvEWaMvXmF+Nuac14NLkRVfwvgDKiFQSXyVH581ExNrpt
nU0Uuo5LEQnaVfYVclqDwEsRG/2xmHbDPZMjeDWdWo6k5fONx/NozOLlhPNMCmsynxIV9tmhWz4C
01x8f1KfQrDGzq9KZKCiAjPbWs5TkcZSGID5wo5KQFhBY+hRQci0FoO/1drS/twlwkZeIi+FUgRT
b6gvhwQd4k1L/omS5oPPFHMDm9aNkMRAK7FYSRgZ0WaZQOyZ6VnnspUdWgHQraAA5ePQSBlGIL+i
fMyGY7MbRo72w4IRs/lrm71pnXz+5gFaYZrunqvTwqsRe2hl05tskt4UDo1ibjfBUmmqAZJztu1l
dfGhpM41dssoRF+q00um4wkWCDgPNGT/khAglAwRHYs9fo1m1ULSpDk81/x1Uh8DRXW+Lq5R6ICu
3BIxmaowDklMIFXPN7YlNerNkQBGCBJ0AKdnofvVTDNlq46o1+1xS3ljHGN650a+OBcFeoqjUK0r
DXWUZCn3qi1xLkfKfW/RwHVP4AnpPQY/lZvigKW1+fsckMTFXv4O4BPypdMk0k9lOz4B2z11Jogq
rOLO7kfE2pAkaK/8hQWXd5SfUdoHwDcNVN3eq6iF2sxPF+i/m1GR/OIP0OQKRl/TJgpKHj49DZp2
c2aHvaplMifl0wHoK4DQZunB7BjxzPLeJ9SjhUQ2fYxhZouwAyAgeMqvxQ02PIxEiqp8Z7TOqPY4
zqJR5VUuw5mH6zAYQS/EoRbbsDQ+Dtr8e69sqbOJftWUXRuS1qyDgf16S5wqr8Sqtz3+vMIF/FCl
ureU68J46gKTMGb3PMWxahLaYowgN7aD8OfcVWJZBOMDf2/bHFXB1wnXaZJauOcWNrP9S5G/COBF
f2YK1Ntq8fwKtiBoe5IDivwa7h10l6LkhcQZLvxN5cVc4LileyIWPz5RZGq5q/od6NwYNc5KvK55
oy6ikkLvPt9ojs7l5OOQmSHW7x8FkpkkseYeePc0AlT+b3NbgfS7MrsqRSgxy5zUhhiEEGiqkTSE
FWnktKipKVtmdkJscZmXbLjQGS2XNbgpTNoGFDHHYd9lBFxTvIxSnfntoP1y3H9rLyfmvQoZR1bU
YZCY5F+84Fmng3LvTMDOqu5PFXFXF1hS6WN35KPrw32JHRKmKYuntU4EZKUVLat4lE+L+ssN4ef1
5HWj+yxFYxwagXoZdtF/qaS4NU91mNH2hVX9ZuZnIVI+Py9ewSrWq+uMe95pRz7AG+BMZVxXD688
Dyh36vij/K/XK3ON24e4aJSQsp/fhnmLwMJ/U/rGiPcd5skY6TJcik6exqrIJniAFteLs+zAEQVY
jfwgUotEkOawLsm2zj36ESO2qWdESTwLmPgo8Ee2j7wBdSmrIex6FDPy0euyeGIjCb3MikQvE/nU
rkYd48eeBn44rmv3CID9Stfgzp34ifwfMTZgIZmpLnccbuzY4eTX17Fw2MeGKESXgjYSZbT+PRtx
XNWMqjE662G4JI0ViCBsaaYGLZYa2XDLcfcsQ/upFAVRFnFg4R2cmE8ZAQzWnSU7PwPTNhkLLp4k
2T0+yRh1uc6ya9wNO2nZ16X9ye/5uRYQ/dZQB1Jrt/ch6NkPFpJYsl+Fs6PUH8yTYNraPlEvufKP
JGdEoeyakzq6nwRfPy2DAMTP1++i6ywHCcpRsZBKvHZBcOVpmMpcOvUWG8Nc8eCATEmDFJEGZkcd
610CTz1NdS+oQL/mWqAOh3PjIlD+4G2fz2sDw3H+QydMpQYz4PAGN7GUVow5QeDqwrRaTS1N+ZhK
6vlU+xpqg7NyhYNvdQWyngptcI3WlsqYlZfBvN0VLheeHtNDXvVwCIN5axuIixa2eEiqRvq16K8H
2Zxg4+IJwtcF5QKsQK3mcGcoUVNliA6P+fzXcm5vwDEJO0fyDWGvMf/g3h5YzQR6jlu5EBi+dklt
np16D0PcmU7wJ8chMz5dnPKkuCbnomSKyCGaFdKg+0p2Y4Skdphx2Sm8Pw71Fulb3i8tOXgT6SYR
LYFYB9vwHMqficTgxaRMMpTFYqvzVbzu2SxVZCInAxRcYGozbn8mCLnf+y3OiBSc2+dNug1qGCQ6
PMZzY1xpmb3lnFZnnV0L6aZZmH20HhzdTkbYEPJzQO6lT6AI+tjwcR9nwldXoXekoq6W6QK/pN+l
Be4wTJkbOz5U1siwo2BFX00a6ELl0RS23x/tYfaxGMdue+mH6l85RRNHzNsIbFdLh1LnyGDmdXKS
kk2Ac2nMduLtD++E+c27lTopZBlyylTb3Uv5FJ5+pGSTUth0YAgr1DOgISXyx3HJLPkFTu6BIDCy
gEozUwXofMCItHqJ+VSL9cjASt28E/+CEdCGdujJeVA+2+SS5OfNkdtE/bUwQqijR9iWv6STs8Wf
mz5iQ8otZOK6SD985+Fd1Px/SKEr7aJDIEDm+xjtrJSQN0tJ1C4ouDxvD6tb6vUiBLTG4q1jWmAm
QJEciutdB9YYEAaolKuHIPZsgBxuKA/rwp556TX20P8pu05zjTOBArJWoAVcYPajyQhIkfQk62e2
q0Fx1ELMzuRm25cnUXGrRUZe0CjJRLx/m6UjivPAR8qQsLK2b97eWwobqy0q7qHFV75KfWkaiPcq
HgJ8s6JZIbkyEV60mfdrYTHC/CT0tN8VRSgtZQqZO930ketQdZbCMaBsO0zX06xUFY8OwtasvMCb
ai2mQLmNC19JoAcHZPNzrBZ0QZ6PKUTi+cby8Eq5Tq6dU/dbkwz7so0TQTN2ohhQh9nMGf7f5AK2
fDnN3NFdUIGmreecRv/0ke+cLL9GXV5VUORPjeMGsOoOb/NEPc2GXFpAP6zUinD0yT5bSD33ywnl
xWRh/uYdxYRVPMh4rgjqk/bBfGAVO1RcitDn0LUXFaqXlrEVfvtmDb1hd8oZZgB1fpeKk1zlXD1C
MEcI7KdrUTFuaj4KwMMWG8MEv33gJtbF7MXAx5UN9caW88vt8/aDX/Qm/5Oe0ptm4L0Wfv4XGr8f
upjxdpZSUP6MxaCHU7kppD3bCNMLm4HSRcIN7y9OiiqBlm1E2n7bgkXtR0/renZBahKvYrDR60FL
VKT9j+p/avfeORo2OO7zLoZY/nO6jz3M5kTycTWngyALXgHq7FeUXZWvQQRY3KQNaXME+K6X4Ci3
jc8NH1DWKPMV1eKTfdwwaOApkq72qRBwsUOjAkPwBOYGZnkndHSKgq+OF5t3lh2zYBwU9xH3TEgT
B4c7L3znBiLmwgXq/zMuxEB6aYXpDF5Prqq4SP1XRnVt9VCKNxUzQO7T3Fz3iRP4+DVs/KDiIqnT
XN0s/ONOIIVDbKQxgJ5r2jg1gL0OlQm9hdfQ9/GZZK3jwJMwRcL2LU7T6S7QHY0S2GwcWrfXpAQO
90dcqpxmC4aMd2rNrjIF5rg3UnxLsHl7jkvBo/j9ggNucy0EL3b5z2qncV7gyeEH80pgMviPDabf
+dtW/NErRJHwmkl7qJcM/F/CEqbokdP5CiDN3fAVzaTCN+5u71bETPvrgN4Xx8WSK6z3YxuDn0X4
RCS/wE6xoc3Tpl+UUNSmzv7KcB90zsv/MBPmW7VkzT4I0xZ9bHcDRY5ZcbNU47nzwZWk1EeT4qY9
PZhN75vmDNv2mY7A8iK0cphTegvFOhekVMOYq/3AZJEqUH3mcgdJ5GMfca6ngDqG1XLqeEzupAl+
z1aDeMxdxuFUq1nQJAOFSbSsKPaa8p28f/Ld4K5MKGo/tGeSeuHK/7MK/rJCtOd5HQ+ivLmgCVZN
G1T4AjH8V0hkUgDz6DK34INyOsEGN732yXbhT+juJPVEUdmJr94I3osjFjPByQxpHNs7IszxS3a3
l/wVbxzOPzaPCtdKF1IBq3jOegk4taHsqIfZl2AqUckiygPym3P6d10HgH8tC+ZqAgRBrVpr0TX2
uAKGVh+XrV8IUAMLwoSDxS1LVOmHZjRXfC3+TT+W70QmvI53bwptLqnj0lSbS4qXBXUa1i6AOtdb
br1i4ryAh0c5TAIWSZkD9Ef/JNu3OcN6sNSHNipEDeF2nmJr8kzZveWbPhcaSvh/ZnivfBiS58h+
RdwANjAjWuPtf0v0i7pf2wT0hhTkoOaetDLRonYe5jC3c61d2w3PO0kf2lQ0KbnsyMLKxv1kvNzv
tPEOwWJzC9SqLBp9+ZtB5lJPL5nqgdLGX3vi6MtjiLfevNvsCVQJcnt6qmhrFVCaXqZV6i1c7yf0
S45ImKGHghLxGvWkJ+N3PJ/HCxUjWSSKqbYHriSEhruv+lDqEMN7U4e73Nk9syVrY6lIde+dDN4t
ziaR0uFMYt0S0akr+M2rv1nlqFrAeLEa1AdqT/czB6Lb4vVLzKGlvAMq8YJp7cM3R9gCFn02K8le
qN5e9X2mAXdHkD1OAWAk7i3BE0YmkVWPXHwEMe7q9tRYzbIsawKS6J8YRvt1j7/bxEJD9pwKT7Sz
cyBfa99JnyFFm2Wx0uQ8mjBISEsVAACwSyZ5BIzNQKtGSDrAvAg2LP5DxTAzvHYqr0AdyBkZ4bqX
MUItJnzk5X132k6FJqq7sgq2ylQ37/Z20oqBuYgAMvRvQTFXwcOzAaXcgHq/6Jbx4nZshyL7NRxV
01YBaL2/RVQG+gV9zUYQDAVQMK3pTUTTf6CVFv9yRQ/qYb7q3D2k5J7N1D0T4i05Wgl9ujO+SOXT
pko+Ozxo5LnDQDMykSs0oLh7dwM2Ep+UEHGBAC1jFzaFnOLl2AXQ6gZX5+eQfW30SjTPNU3yLuxE
8e0U/4Hg+8vJTVJrBgbOEiHFrLHsGeTDIB3KX3PQ7N25p6QKL3fM2NSlQwEdKxdBUCDmZG99+t82
y9YwfbFh055sSHIzRa5pruFd8tdPEr3jnyDG3zAcKhxbvkG2pYqEqyOD/P9/X7z+U8oqqP95T8QQ
hq1/U/KOfskPlrCni2EpuyZ+6ihUTn9sEI/JB+IBQuOgXTe/eomd3f9PK5/di2Cw/G9fP5E6hzWC
02rg0MUR4+KEVuPB3/VINpJpjCJiTXiqcrWmnOHaPAqIBzqVVO5bRwjpb6blzyptW50O2Qd+enao
EP7wXXdfUoATug88uhsM3PSSdasmjwfBQL2KBWVLEhCE3B3vRqTF5GZTmX8uSxRA1aEIHZG2/IL2
4euIvtPrD/f1PGym371rK2Aea7emil+nspPPuL0fRQoN4UpuUGfw8JlW2i26TF/FWigfdntVVGU9
/R7lkXAELZNDwtd+twmDMESPsVKhqRJHwk+2YvGMKp8i/Z/8CpriVaP48wCIDJ/AXXvfG9GknQtk
ZrZmdg9UWLb55HbjkjB0SG3iBpgZW1vzAmpTaGftuKlY0YgZt5fSA8nBqmvFWcT6xH9gyWtlVuc3
M1KxqEQGx1UsOSc92MKoR2xanbAvUgvBJyNgLF5yND8ppmSlnDsb3YsxMe4OFNqOUkRtCXZe6sOP
/OtyVGtMfLzDNrOrYLyYSeKE4d4C9khSgxluxMg4o3OR01NtgQ672pqUqHhBGeO1OQjLzY3j8tPh
MnS2qWUkCfBMZO56EvfCHCnmx5EUh1/VaRjtt+ZnBytkLRsUr6GJwk4Xa8r65RGNwfrOtRRpH1Ig
cipkjWKfuKN5jC2COKwLOWNZHAOjsCfR7ZqgssYLHmGkd4rw2Wj4AclarDbCLgBtzVIDwFP8iJ6J
aY8PZrxYPj7FUgEM15GBg7U2mZFkZ0FZC9hKg/gOLPrHQvLCLEqHXobM2vyijFD9OeJsFRtcoE8T
E0tDXmQzRJqeqtNaJh1nRFtdfuliJLAqe4LssfwIQn+699oad4O7mDj/46fvA0vVJXgLfipRnk9H
z7zQFqF3hw1UpI0jQGd9ebBIMxemNUGbF9stazNG1sGacfyJ4MWtfZPWG9XCeun6XOp3K5lfj4/k
GM41eRx58pzs0Jg2z7SiTbRZDD8sZsz7KyncogBczae8nw1g13Wyyx8m5Tk8h/6b/IjuSCttk19M
OZMA3Gm5pXlLSnqr1C23hKDH+opH762XeMdZhLAz1SeenBIf7reXt7WzZ4B0aYePwu3aGfqkduLr
Ut8NVffUSpUwzjDbKDhJluWj+D7z9WhCSB27zxoctghWgp4d1cWJcecD4oY5LH7YoEzsC71BGPpr
l8dBFEP1Fpqfk884P0IHu7VZ0d5w2OIZrknB74IDvCImLMG4P1UCULwHwOzcZ4sDDEPE/p4LWYG1
mINF74dGm1uaPhEihvKXd322y+/DOV+OpUmH+fAyVTP6nBDNH6K+cnGllSKjswczT9pGEMHO9zjD
Oof4mDRwkz8EKOiohaQ4EwboZUdYJ60Rdf7ZWBruidVtrgFihIXKGIYAlEHc64BQj19bMu02+Yrh
dHO9K/GdjpSelLEYCFWEdDo1NBPtTX110/3MJzQrcHY1ZZwm9lN8oxmKNt4bNMcm7s35SQVvN3Mq
IOGD1bIFbLTConQtrrb84gfqPd6j1rJglH4YzGFaT8CuaRTHyOaQGzraU82J4VkF0SNvzzjPjJQP
v4dumAIEB0usR4a40CCrtg1Eq40Q8Mp83v69q5oTL7VewsvDrSnScnqi50t0xPaCTD8EMQkbEjHd
WwNxpMLtyU+cf7kpgrYHS2bIx/G95q6W2JGXovhRnCMtPfBBX+I63AgHrbApkz12DVQxPhpLvrhg
q/pPOWZKXieR2MgJapwRlBF7b/KaRdN7K6lqYXfcK5CRT+7sjO7s5KdSKueVbFsVukJcNeZalILT
i7IS1IVAJlwgoONC7mpsn06j0xrDBqHhmRzYD8U3KMbbo01erNLw7sY+m0gD9ZA3n2ZXsq7ghQkT
djZCO9pzaAYUB/pvUpUQ49SaxcnVNR3dczXQEh6c+zCHBQCesUekwHFiMK1tUd435ltY//zZs5iB
VcbSjI/GwQYajzgQr7NVsIhjDOqLcJIPIDjGg9yDXUeJZk2vtumKc61H4+T/RScAGs4Zks/TEi9s
LxCwFDX5YQPeLGPd4btUhYlfvayAUXWB/wiDj8pOWtwpzeUtz2hX27bBUlNN6wyiLHbfWXZ9u9kH
EW8tS7t1EQu1h8qEvsm7UbgoRjgx6vDPJ9aSxGjuNnlyMHX8e9+ZqYXt+KwDNUI/3eWbcQjVA12N
W4QmMEQRoSnqkzLzg1ROSKfX6jtJRztJyPTrJRhIDN2jW5J46KpSNCO/WIhyxqBJnidY2D1dwdmW
eNPGmdoziqTjJ8KUhGHedE7il2ZAyYEj8n7/ltd8okoQ24mjUWELWSNGEC05ow+dECZ9tU/naasJ
ofYJGWq7UkU2wPe6LDioIhybiE13WPlu4SWH8zB4Mf1HmoSofTD+xkVo4gx47mWkSZnavcm3YeER
K4HRs3G2HmNYsxucUhle5fY3ACpkVy723lPUAM+HvpOgO/FXKYVJdjNqMnFFreseQfHziQNobx5w
0A1YJEbO+N8U1L/YKDsa7A5nM3MhWu7jXq4Fj4sIgc8FgnXzgLEkksPdYC99eridMZZyADpR0Wb/
6JRtq1AK+gzy6lUBlu6fzUiySc1mJRGmIE9Da6WwCS7XTISUMsqm9LbnYmOzlfjveDtOgTl+kvAm
Dbx380jzDaP3woo1qXC3QLK4TsD88/B0l3byo4vGR/q8Ud1MU8CFfg0xAOgsNo0sO4u2B/sEVK/i
NoE854O0mO42p6v8jMF5/rgeJzxA4C6YvP8+1VLF4PdH8CgxpH2bsOx7h73gzjrAWmYnRQPRzv+V
/pLsGk3TeISXv/U4/2clS1/sXJkoltFuH1s018Tr8n9HZdijOop/Q2628US+4pPQPdWSIC9x9Bqw
bqVaHFM/SSsu687W2A+pTMD3fUdk4UHX6Z5JRQESizas7m3CL+6ZgY9DVsECuPHKgCHbOquJyA0q
Lo1iZq/jEVWvX1qLiqTzBYjLhJ6Cto4rhm8qoQhamemnN7gYhy38L7fGfAct6d9mlsK9EcT8zDE1
6eFyMCftgRaJsCEX2UhZqMHbSTYeSapP31ZBWeqFgEZDxrMvd1mT089L8QiXrjri0VN3UiOUwsQm
BYYf8M0gkBHbxedy4ruRgeyGeeBvNnTS8AZJab+lnlu7Cd/qNoBCbuOVudazFGjVhXteEzWvn71s
Js8ldiUV7wXcATmfMoYX2JfgWSwCySvV/7A1pmhlkw+k4ISw5qsBHFFTPQECAly8CBhBk1Am9AMY
3+EFfUKhuHX1SCvPnCMTsvFkDJGuQlLIkxpV69s7g7LCDCjd1Ycvm30eWBtO3e2HcE/c8G9SRq1+
poHlut6gl/Gp9Kat1zCw0sl0vIqebFT299+9143D81giD4ltC0j1JR2ueODN10XzZPPSni1Th4Ys
DHnqFKBeFPrzGtrhFEPZEWKh/3j8vvt0NWjjKpYLxSWi8agW2Mg772Y5o9Cmg1DzmAPtzYpiyZBL
NR1zgHzsg0R1PP1Ckw4G6bpSJc3pM+mpH83Q1C6NxaWG/N4gnOLtuw4LP2DdQysWOa2E5oDENdNf
dHcePx1emc5RcechhR2EVXgHQTRaXLokjJ+gFm5JdlzqYcmDreDiq7eZQt+ZsWI2pP9aEEeWZzKg
nATH9Q+SVVdzQDmIXphRqHtJhgLCJGGjy0q2u5eC0MBnvT5a0EdmC6zO8Z1BA+uRIcHLuz3/Nm6D
XLkcRFQaiPWwBqPRYrfz9a6/ppgtQkaMNoqBNim0YvQrJYSB6Vbl3T0Ptsfs5rOM9jf3VF1a1VBQ
gnoFCW9GZd6tXvRpc+yJhUML3CdbmNccnTZWdbiwly01glGxkPayKd6aHSs7II7/cN6rToZUpfic
tRXG8nKrHpFkKSDPWHl1CTYAsRF0kGC9AAKuXnYjc84KWPUf9OD0qeEJV2sYPuCDM8ymqW9etyqM
zpPspLuNUZYPRlRIu65c5oj41hL/DzxL6QKBevEnzSEhFGajlbtLtLLNzoNLaNmptYUP8DzcsLGC
w1s/dmSGY7PaFVdqVTq06FuXoqLkt/2HmyJlRUYzuTi+fqjvwDBGaD42HdoDnn985mS77HJCM2Ug
hcbt7Dn84YBRZOkqTQvkL9RQ9kuOBLX+lJ7iU8mIJb6QReCko0diXPbRPQDxe5viwd4JjNARPfBl
szqZtEuDp/ztIw+OxaiyvsTdDdO+y7ErA+APzSHKt/cCoDPvFHl1X0xg3jb4H2QarZAvP0X40YY/
M6vZcP2N/LFBNJSs/yGvnPqiVHEJlNe//YcArlwgRcXEKKhsWMcevODezVcLAQJ5wrYPobkmDime
Apoqw86SYNKuNI63Ca008ZdbxCjsF7Gv0X8i0nxK7rzBv7ri7bzlh6LOenIYL7RVtt0YzG/v70kL
yF83fPkt46WQe9NQJHI8Hb+HDFMuw4NUiy9+PQcRBRsTrf/lALZOgMlitlwWoLzlZtfuGZ5QyboN
ZRwQUEKbqYTapqsY3Hhdaci6Zm/worX4/KgX03HTOxHKVA2dqQCgUALlLyBn5ZlFQsZudGrptDPr
A3j64IaiErGzBtQvneGQdwZNVFFKU0Z2b3UM5rfJTlolrSrc0rw1If0oTVYj3ZXhyaqtT4bx51l0
fX0yDGHZGg0zuuGTeOgHfeT6DtjNBNTkTEQhXUnea9F3cM81MXO+lc2+AdzI5rloTzNBYsQSMH5K
nFvCAzJbLfRbJZ24qf0zKsUTJF94/2q50Bb44io2YdP535bPtpdXHTRanu01RsaVqclkCD5s8vQX
DGZqwhgQ3JTDf8ggr6ZSZDGQ/jcSuLNLvEv5mXqDHx3r1D/Gnu2Z7oLh4XKPXfL3kSQCUul6W3Xd
fzk7yvPdOj45i7XN0YLZKpsmO11jl7zxdr661JEc1IU2a6bKwYYVvFXLxbdccrUI63H6jI5algd4
742b9uwvt+t9So4Tj5O1uC0tFjJgh4O0yj2ZuKeM0Z9E8t/UD3LKOKs/4A+z5WYxM5PUJMCyN0Df
kU+fDDxJCMt5cVIUZBBqFS74bGbQg89cNfZEzJWlG5mg7UtmFJHZA93h6YeZCNLhOHredgKezKp/
EsbQykv/vFjP3IqHLqeIA+6QkvPpLwa0cK1Lff9p0Xco7vHXF6DR+lXyIq52noYgSYL46s94NQDn
ad8aKasPTm5/jNnwWQ+tWug9RTymu8k2t4UeDeBhJsoe+KtTPBmvjbJKRkR1k1EL/bmZm4US3Ubl
4zMi76kzuEiCU91/HJwsIDQvlIMLxChOe14dZuI4f33GBeEcRaxzkLCvjGX1hlVeRNPEcNUG/s50
YefhjJW7zBsNcrcMmP/DmUjyc8x5kuHlPk1UQHIoFScb2B2+0gY1EK0cTM5mCfbRLJ8UBc9RQBG7
8MKq7kmdxpNBa/iKtrJ4pyGZMLV1QV1wK9MlPafxtXJQXgTW2SAOKNVfW7zDv9eyZkAyam/MDr65
XMmU9U6EIcX6fGSlBETcEUWaz1Dr+PbFxunTnssNjle4vO8sIu0l44uod2myLlMWk0JpqiAd8ol7
RKCK82XDd6gLAMtkZs6wsnxr8HxJ0uxGFOXPMUHSiEjeY1NZCubeoqr9FT94y8oIqGJge6rTqjRH
bh1dEDJC5v5z45hjfXjgn4ieRdRyZGZRGVjhRcNrmB16e9Q3Mw8PDJgPT/LPs166Sa5vhf7bFsBZ
5pUEC2jToA3nRGh+w78cI/hbENRnx1741fGTJmIG79lB3TmaYIEKGPHbzIxd0PFQ4HUYLh8yRC0i
x3luBbpDhygVmiBxBry6f6bXRXxVoM++WJun8z0sCaeFqFh2GPWxPTuElJi3LjvJobh0qS38bQzn
xcC+160cBtJujiLi8aby2Q/poBykIycxwyIv6w3Ix855kMsJJs0b+0qH4HNhaefnzXRp9rko0xMi
ipiQYfvYAoSlRAq1l8nMvwB6P8pcKp+3JdMcJzsC7nWQGIViHEnuf9vs2T1ti2MyBSKfxbUWVj2S
ePPKAeVUuBuemjyGSFZgBxx1Asg9wCGGtzHddxSIM+EiH9LQ4pNSZxOSuieOfUfM5d+s8rMROnjy
bJro6VwsgQ9rxLffXZKTZOAGsrxT7Cp/eAHkeZr+s6EWklaXg+TsdNl1XehlnQneOhqMzwyhqH1O
PIwuLCDmQV1tcW417hfM1S+mWtlGBTjvGrbI7og2Xj+W0NosbRZ8piJezz4HG/C+LGYDNN7ekKaP
9vM1oD4Oeh8LnR1E9Lq4FZJ6xeuoUJbFLBOR+CRXakXY+b450DrSALMF/lm0CaTnTD/BKjBRnrXA
t3dI5lTgYU8qRoQ+qTXdvn0x+LsqhiPQZfqiGwZRLHxJkqCc+g4wqGVvImjmxmsAApSbyFfogn0P
10Wp35gaQpVwvS9iD+bccgjHDQTtFFVuYZrc42IAFqypPWJ1omQA05z79V8nYSt5p1mLsKHemh1s
AXIBtAWqrAb7lA+Na27Lr/K5ee3krOwr/BOdsN/L6lMmiLXobHrbfzFVAedn9tKUbdEuXwBSW0zn
qt8XiiLGqJBb1I+oQuNIgeSkVi1sxCX8Te+WWJuP98a+fNo7IBZJlJ28+GH28IodQUBH5UM5lko2
UlEKlNpvE17fvftx98kV7aRfTFgIgOpLLfUB0OvgLj6Bdnrk0i71eEJT5j6oneVZ8++yJiH9PTfc
N2mJfxD5zL0AvpAZ0c4CzSS63aYbkffLafTFjTvVp1wvQLipAT135IUYcn1aMFwXnXCJUKZCsANQ
D4mM9X2rr90h6q76Kwh53MeSRn6/i6YAc9VbqQdFVZCYnMOV9fusVChTmLjWu95zvylwizySTnS1
kizZ4f/kA8jprguI8PfCHplbdg1CfWW/tORl5yFZrHt9VLy6iJ5ZWaUtcF427TYgN2HqifwJLqP0
u8p/1VYGSN14O5zwesh10V/UGrDDQEM91bwyj+OjmsYHHio2T6yKD2tf0U854Ae1FWQmNYIFhiOV
mlro31sZKrgccwoevivZBZD5mMAvfSm2LU3Q4mB53RZ2rnZjbcajz80rgOiIpEf2vjpVkHSK2VUr
dgahtDI94TxiaAhcI3WV5aqYFsWjcEnTSiQxMSLJ4+LY0tHYCoVg7jl20xudmaebQajLoxBtfovx
bBDIx8RpJsBe0MVwCaAjd6Ix292Av49EHDgPGrUxYKpt3nigq/1dS/Acm13KcKkdfjQ+H1zcmuYR
0ZkD693TATqe8ukWSozPoJvKtJN8uY4fe4e0s+AvbqLixl3/HO3G6KIsYsBYRG5Q4FCy22RY8yqd
Cu3sMV9glwigDkk0+C3r4bofN80FPoq8YG46jsoJKH9is4rQuijlAQp6zKWyPnR12LFePXI048GC
WhiVzYZmCB88hAMcws8RaQeDirZX7c1O0Ro3oh27+OXb7uuPswiMo9HtU0kEEmHBt/hhcIJ7CVYL
rXojSXDxfI4JjHfZOZyvpBlKCw5L2pzIZBkM2S+9aLx2mIueFVTmzeQeVwAobAlQ1R8Wfh+hE7F+
wETyVRCCApSWGXTtop4H/i/DR1XjPWjoU5Lz8zY6alxQ2h8KSRluwU7bYPfIPxe4kwOJdLXx7qmn
OB/x8qG56hsOk0OilS2hqMHKJ/gcdNahYjX753+3D3MTQ+xxQ3NPJF1yUJsnbFKrnLFzZm+wstFB
kdQ/ee6mwrv7c//f6UW7eyI4yzFtxYVH1zQfEhsEL1HeucRpL+Px85U55mi4mv1tXY80mlFuFoi/
DyfGX1lWPY3r7IMDGDSU6K9PVkxIO38qOWvkLzdyoul92puH4iOiireqo+k9JQjgIBjw55xGuirN
0PSlrT4FOpCRZTC2R44qDp8ueJChV9WmJ2E503Jr6/Bd37M9Nh2P8tkIhtbB5h4wygYh9oZ61qZr
X6Agb8iIx3HlfxEjMWdMDa2kBzqeFt86JjFiq8WijEbttUbhqVwicBqx7oR2irtRffOacEFGZJYv
Bd+GhmdG2h1a6GeogU+Eo+BeeWD9wNDYAdbJqH0kzv2YjENMDffqfs8mtxYMfrzpohMPc49Oi8Fy
vD4xBPTnkbvORhhx9rEfkzYMUnzFN5pCbNqgeHAnWcw5hOv8BUyxKoDeAnAyKV+yWHPxwCskG95R
vzUAMa2DsdYSFi7kIVOpa73A4DHJ3CMsLk7BFCOZjkwx7H6dhB5U6yEqJyMGPepcoEd4ASq6jh9h
GxiA8cRhOiIbio0vqZhQ5cXxbQcI/+yGeEQK9AXy/l7e51Otuh1X1DERrNfxYeiCrjZLkG9rMouZ
ffdmOy9jbtyX1ahZdZjd9PIfi3ZI7IaVGjnAJ+EsRNdq7eGkmlViEPFdlsPNVSIWrzLc4QLC/BY8
+4/s5rRa7OD5ucAlpsmucvX70zKc2WMKAAanfcTc6brKz305tPQEHNEa9TfqF2rkCrx5mMjJDDBO
RsU9WgcHLNTHDkOlR5vBolZJ5vIMi80WseBqyvdjjIPYMnYrtS2ZbsmQtWQJxOc20v/smq80wAyP
xBfOBnN4NBwJhL9MU8mY7qXm42DKE4iyH7ScLs2FkxXi8mWNlkPTmAmidT3iCsrHi9gWx7aGFM19
slA2LnECI8Vh56zczqnsovFV5qrTD1Oey1kdsWE3XuC1rQPJ6noUwnps+1M2Qio8WTBNIodu5mk+
p8IVDnrTXqajJqgo0dvesohsC9t2NoLtFKbC6SWkWQcqOuHMUIZWBHd4PyMqHxNXexTnoE+Jc3kt
qSZExCCQezp12gHPM1tpVGLNLfgLvI9Szc8Nv5FRbzIXpvKclnrU7IVqXZdPSCf0QX24fEyUJ/c2
A12oVSwsW5/2VBMyZK5ZR0ZPLZS1HSFM+jBeDT2yl9o87M2OPGsu4NMyeY13e90pOoBWL/MYbZ2c
+5khomjyogQwsFwoaer6hU+H52rEPZd6CHMOA8y87wUOw51k5qWSxCOlr8J4Ezx+/uEetc2HeWZi
pPJ2PPW47JMP7WwJYHRoUYeD6wEn6tbfBpS98ayrC1iZbQ6fG8T9/EtNuD37VGWgBVqvcz3zOJ9T
32/1XETRpVGy4gMwPxWEVDOPeCGw85Jqq1PVh/3y06Tl7+DDVMWFWtQjzItMsusBKkIaww4B8wMI
B1djtUrr2ffk9flEcCa/iK3ybWutalxEIJC6azwRPmKHfwXGAUFCmcqmh6J+G99qVjeHhLj2QJ6k
W4sRWf9jTU13l6CcP2XgGAVPwaE6dXGbEytv7/VqkeZOBZ/3lFQUWYifuUKhacVCgtK6d9sitO5K
fmdeRoi1Cv/NNANwdGgSvVuXuKr8uSRmGdDf+gJCEIArYtYzEeX2t526aNCD3uWRkAgATU7KqYwK
8kRNn/Pk+9ST/oezWKV9O52iWMvyFli5CI0ZLGtZuOnunMYrW2EYG0U047g5AuUxr0IjLMlY3leR
x/b1dY67fyFiJCJqmmxzvnVmGY0UveUZXZKdAAan3zePApoXXqDNyKXW3vdLLSp2gVELT+xO8UJH
ZeEifjfT6QWhenzsH9eCMz49hvb6h03glnxR0e9SjIciKeZX7N3lrpRDQxmqNNi2qnQvKrdUf88n
fl8a/+nvMJnydK1/wXVzJDGP/kEr+HlmWRidNZz0K5zeHN4uWQIQHNinH6tBqFpDhcR8PpF5KYBg
WfgnOn3U8WkSrthl0h+0AZT7eAgHg0Qng54cWx+LMKM/Z/DXdRzwhogvnFYcjYDWzNazST1bFdHU
QsCKHkzt3jzFdml346O+OMlTNreGnPvtHrfCQwGfAkaRJpyo+8xEuA3fTu7K1czHF8ul4/tZNux3
GDBsZjwnohj0gaHtJuVgyKpxHGkOZ78e+GdchcXHKBEOCrNNJ2Tk4iPFHUlbEXmmpqdTxdWfkQGN
/4w/ZBlLN8Y11ewXijZSgg1jJJxgzSn83dx3Om3DMfNEcJ2jVQaEvXBeL/66/1RCM7K6/o4rdeAE
4H6ySqDqh1/Ifzl711yBCayiPnCiyCZP+b457DYSj22o2QczZuchKNAc2hL7Qp4Y6ZK37P0PKhGj
VKepILiPK4VF54hiU+j+CrFcMWW/64U6FodrDaV+ZM+bSiWaZLtTGPxgSzLC0MGzrWxvCmNam7Z4
5vcqChvCBenN1cZ7JVehusuWLTDFUyKZ5+Wzs3APpufnPjIWTPaMgZXOI5DhFTbZXl7ZasGtRJKg
dQqSXHPGKXbhUuTvfTAGMZA+Aa5N0VFPuSjGUMVpzp7EhYf3hChvlG1EKNH3GJRxZX+IQ8dVfC79
sU5vrVgN4WOh5moswenn87SKAWA9Smm01tub50ppidid2MGMQhoGXptUomc9X8iVsccUBeofoE4E
huTGiNZlj2GMspMfTAsDxFX8JpqY+9yw1ChNfN0iO8xlEORIBrJuA5ReeOoPrdR8V1RBL7YS/Ewq
nPUO3bHSpAH1EUq8P601oLLA6ezQHZ4ugvNBmu3lMeq7nGJEofhNe86cP4PC3vmt2T6zomn1bMQ3
i9ek6cFOKoibf/ssqId+Oj5j3v4aPuHLOOwoMF323ra2r4vInRPtccBVX0pz1mWlPYqExHWoZ4dH
YNOpLY3dezpAIrrrTAWB/CwN83nX0EmTxz1g/YyAc5QLD0Cbu5dCEjG0FP3riHI4gwP9CcRjaeJ7
h9phEmSrJ+4hE6pVe/wL9PEhIi4YjKwokGGOuCIOmlFR0zkb6ZgTBQMzBVp2jr0LK9aPX5Y7534K
k3gc6r/mI36ZQgDhHZOgar/K81BHF98TheUlQaYALpr9EsQd2an3F85e70QuINujITUW+89hpojZ
IMxy8H7ZSpfxxbgKwSqEnXKpn11y8czXAejGs+6QXAQT0EEUWRzod2QKbew6dVj2uAd5JDpJQe1+
JJHiZExETmAttgIZ+tlEKG+QHK6shOVAFmpalFN83jdyAmEy86L+MJGfuOlmrXIYTmfJXbOFgigj
1olZXo55/Xi+2U+pxTuJbxYN/SGwVIyfH3BRphoNmQnJ7XayttHX15Ks8EMje8lWsk++XIVYfaaA
mmf703CC/SIV8crXiLUFodJ1HOPCfpM8L3XCJVG7un5Cjpf/PorN32EH+oi3U6P6FuQXc9lR9qQ+
xHbqngfq+vEg8O23ZCLwCYoXuFKf/icrwt52ddHY/HUjvDB3ugaq1OjCD0PTraN2I8s1qLNMRJK4
IqMbfz32v52M9qXYMUq2XFhIDOqrpqvfg/KO9bpPw/pY7idCRJeopHs4HX7edSl6NrGIOwNmWc2W
z+mTiGpyNqyFCOhj7nYhVDTnphvIpfKqjl/fmqZZbm9TZhXlMSPPFl6eRpzHUr6d3bo1rbKtKhD/
bsZHbIOdGHBvYrHaKd+Zj6jWL6EwxPcr9msevmFtQmuGWd3qtkp6fvJLoZX/MqUF1G2WF4Qct7JG
k1Cw//VsOiuI2x7Xc7qcAtdvRdZKw4Xj1L94K5WuhAyAuBDz+ve8L5/Hzfo1xshaWnmmlA2lDRPg
SOQMNcgi7byjpMUYNq/9LwfARrjQMPsxqxOlrJh1KXKakPaidlMIWAOcfFoHeF0+Pw8f9MrDLmXe
oK8Oj8tDHwEbWQgyjKxqF8Dvvoaeid6AY2x2+L5zLAAQlhccewc5ZW21mTirWRPGjVX9BGjIku3z
vYtCXXIbxs3OnbRIxtP8Q19eH8CCItkN/FVNIM1i+FbB2QYVa+9La4svdSJhm8QSyp5M3Tvcmfr+
/jEpMbX3f3YHQFEc3FP5Rh0qASaAb9RqOboVG8b+Jh+w6hwAwm0f0cJd5WJBqpZBT425JpUIFzrS
3xMLXz8t6L+5P66uzn54RGs65bjmDy5IJqEBnmg2LnvbVBMvOmzZDFEWWM9KMUpb5/MwtHHNZlAL
UNy4DYLuvm7Y/Mi2mtWJGui19EhfMhGILAoElkGUkpDkFIB3TOtNbz6XrjTlodqFzf0NRs/5Z6Jd
zjtazp4fvGekPfWVL+9IOM/fnKQ6XvJ8KkHq3p4G5L3s6TCpQq7Q+kj2WsSmo6mjquvb9IacmCU9
SkIyj/n6QNU71vDTNSefjNiZ0KCQf1rznlK9QSj9b9OfqjpiB8Rqv56FlYjkpDuqRP5Mv3EW6oOk
zR/lFk0YNF225wUaUvV8UgnITSB1bunmRQj90qi8Z3ogHW1xsyDB3AWSbU16mvYdmSkPQTEMH9BG
FYb1pFW8EwZlCE1CYLcCuPR2YOPAR0roU7ktWRBDwMDko5mGjGC8hJUfzpPNkURjseTvHF+9QOG2
ksUQv84M8gNdtJO0IqKklPkjZtwODiTTXdgi1hp8Jooz48Tuhqfd1Xv+f02VVZ5MeRD1qDsgfrlN
Q5Ga7M7y7Wx/6lhswTOG9jDOK0pXpJx/HHBY6AxqLAsZz+pJVkNcl8DOQ7avF0IOG1Bf8UFRzBQp
qCrmjzOdyroMlm7xN1Gt17pPY7fwDhJbzIl98uJYCSfKk03Qawq5deIjv2kh4lLwoGEi0rpoXc56
zMCjZg+5EvayNKvpTyskhqPTBE6mJJU9HgfzUmZwZVrfk5oijRqcZxUo0QZE6jwbRwuOpWqXw5gF
Reljixca49ufda+IBp9yR7vIuuSS0kUG6EvUmiBNDbOXCtvvY575z0TeqQ5oVIZLR6aY7cA0pk+8
MYtsqjyJMe0+fs1UaDekVg0nwriEEA4/rsG3PwzGDi+3vdZs1kUmXR2kfMVsw7tmTfyeehT+tKSx
ywBkXshRWVfXUEla5ixT8Tnx8+IIJwJ/Ji4jr05tqCvUJswAkbTFn/NNPpCNvdeEjDkD4yK90dgf
8A+AVQdLXBBCs0bkKZm3ViHtASEebWuZrCNvftI3lTVDVjF88XxKZ8j5nFaCa/V0bIG0XSgqDMcE
m5xn/qPQ6fa3CFojc5NM7zaVWf35GTZx3ud8O0Gw7nTSqbXLOcHw8wl04/PDkzDmPhlPLYgrouTY
vGaVw8sxEi7xYTpHZiXutPUE0WZpuGIMbP+nxZ3mznJZLjR4xs8emfUfl4EOAkO06ncqVkBOE9iY
kP4k+AxVWdAWx7Gt5b5Chy1SUp7F4o0apW+0X4ZIhd8bZU5yPdTE9uPSgQN1zrTpIN3lwC/GmFM/
k0Qqj/0BU5qTyOvLg2dSA+yCsWF7ShSC8ZKnM61e78ohm74qCsAAOihb/Xv+ZM6SOwnKeronrwVz
+qr8XMB/U8F3bdXrElHAp842pPQBdwAmL8ROgXg9tr+mUyL5LaeckuPD132mGO5hC9Z9nB71VpUc
oXdKz/hT2sJY2MWgrkQcDNnC2wAbUJL6RaQ2AZlwozc7QX5WpuJsevhNaRGy9eliq4cj49wqYVbn
6LzjEGWj9Rhc/tBWzuH5Hru4yaX37mJDXJYE5U7skwbXnLKk0iJrXvEcJw0UAaGJc22PGfKotrfI
7d5I/GYrlK0J+Z0hJ5mGjCs1JcYhVvgIHIapXDJ7osPBA035j6TBr+GMRrYXWNjPtrZBWrTAxe+7
0Av/cESDauU5EmHlOTKvNRE4/mhI6rB3YHkbwN1wSNnf0wqb1fjcpwGVJEIOmXVnzw1tma4VCTDZ
JMYSBtZX8gZrsX+Ee/Muhhi4h3w7xqjFYjkf75GD16jAFgAvoiltq1JQyncl/uOyHIyWuabLo49m
weFrda7Fa5dj7JMuDe93mErQcDb33JgtvqGVpZGXOHz3KlD/6p1aIZQjBipNKUgiWBvuA/M0Tn1O
1Tc1UlkWlHM9VoRR6wLwJYfzJsFWn+GYGwLEOuGOtydjbYBD0go3VLNkKxB71e0N4PU5FHY0UasZ
kPBfJwCOh39xQ3iEbxsfzAWR1wa2AFIJLe0D/UM0yq4791R+hCyGC1Y68CkKjz1yXhtHEj+QJUb8
eDjHM0FOhl3fHlmZOOlyfmb7BrEdWK73r93kAsQ6nFqrC318jLm2deuL/XTw+QUrPNZR8OCqwFgl
NSJkI/bjVBRGW4irM314FHMEl4llfhif33CJJe5c6U3XOWaTZ6noV/GwouDaurasZ8ZjFgnVmT+2
v5aGR4WMopfkPuxThttyk4wgBiOaH1L/nHWahQUawPD+ZXRcbz+CPX3RBkTHhuGV+faULe/QB1Ny
R6RAiyYLkbtYd3Y4EFQ3A3KQZ1s3nuKYffzzKacJZ5CiO+Z1NI3lWWTS5N3FTOvKmOSqoCKTJLdr
3dYOwg8pcOw82Ax74HwPZfgCzBhHvRDBlvAm1LUNID/e3MFTbnDFxxV6f8m8DS3iZFAvM6C6bner
/zuryvZif+tVgSFd4AyRL1BJcwZZ6s+hUtaXBQmq6vs9KhqVSgEdWYo3PYy5FXU/1ljSZG1yGqyH
m2Hf3TgR0wye1yHu9JGKFeRPH5j2hPLIAT6L84OJGeyMW/zGKgzsbWHd9nIQ36pwwe8R+kfEqQUo
L85T5z3xUw25xxBUJM2Vb5kerVg1MKCTIUEf8YqncxcbRPispEkb6xLQWhW9FU4nl6515TV/RiyF
u8iWFzut0CV2BjTX+wRzQ4mjCFT3lsLYRkroO4wzy0m9Ti0UBq6xfp0b1T63z/QGvQXfn5AEl79b
Xiy35AKr45VC4RYBI0Y+pgDVDCOKZX5cdsrDhQHcdmVwXaJ5QrfzUMQMvp2Tn/sXF56vAGNSNOz4
7JNWACo2HhCuhxlWtRDTPuyNIC03QOIdyvWjs4hX8Znugt7E5tgebMfVsaVCj716Vr2If9IEE2Sq
jM0U1Wk+zqLq9623WzH2tjPdNFYc8d9RLtoYpgPVVAA65v3XnccE5NMLSm0OmDJysyKE2f3MeQdo
tzhgLuN21uLOiUJrwUA8Nmknwzu9l7vOHOgKCmE779UMkBXg3adUxb0AONhwQuyBFC7TBv0nOwUa
juQU9TCpQh5DPWgTI9fi5VbvQlAJaFGxWav4LVf0QFQRXEWO7+igPU00P296/7g9yMDTPpFyIS3L
3ev3gK8BQY6cREVaV5vPCbIsQDRZwD8hF7KeDi4NO+qUnHkxUvN0wDV8Ds+ePU4Ot/XvUcyo6ZO/
gyW+T660PhpQWmdQiTZL22Y0t/xU4mWoco50ds/cop1ma9Cxmmc1qoPQmH4VZZdWD7wDdXaVlVOA
sNSE8aEQwA7Zieq19tdznEAxovaah3Q5T35cRC5pUdW3JD24YtOaFk5cTPddUWzjJgUBsOF0OYSg
35hamxWud3OJGXkXgqvBfko7L/lZ5unuU414R83hfjDsakOeZCLADZGxETFqy1+aTV8poHIo/Mmy
zNTzVPNWidXvg2en+hT6Y+mmKXLzL+WPEJLXGzseHSCk19D/0MMkLEAuaRpAYDHnT3XXRcKMlos9
eLv0WUGmLmvnXVigJ0rNejTdZBXznFc+GVNqunSaKhoPmlXL/mUKtop216L6G+Cpv2+Xb9eTrLhk
LXecTaUVI7YwfSuwS77j3OMnlE+T71q8wfVaxf71eOnOeh/pJOKOSfqSDxFvZvL6h5K1cLOHfZn3
uJ/2ZWmzFU4xCzCoWNb48eAy22GyCq+5korJKU06OJzMtPOVo5zpgw6uS2r8XDM46RfLOzloXPxr
nA7DiyJZ1wvdfYfnFfPEawaSoSWzw9/jvT1OPsv/1Z6bw36J/+6bTJt+YC+Epz+o//Vwh1gtAkLt
jiun8PZgKH0g18hPZrqjdnELARBHg/kq9k9xaeZMlBHwOBbHgvv9mYYQEQq8KITl0OdjwmRn/Jtx
390OKPlrr5Xsnl7VWyAxkMcBFCzrQBTbBd6Nuk5YOTVV17OUbVdeeTWmVzaRHHAc+k0GB8EjA5XP
KdXQAfl2JUm62DdUXiPLx0bf/a+kgrBCfkH8esg5erMBZGxUmbJBRg46UkaQMWDdwiEVv5VR++8N
sxLujy4tUkUYCdmlKnb2lB1HulEZwSF5bvz+ngydK+YJF5kR3VOtieThfqEsTz9y4TxFb3wxm1uU
sMPJ8f1tF3m4LIhhgi/OvCaFSR0yw/nKwoKuxOQQTYeIrkQmMeVI0jfYFZcWWIahuFwV/qMgbSMK
WNmF7iKS12L2DOPzB3xXOE92BbBx+/TRRJzt+E02zO29MDt3X3R/nTurVtM/yK5FyM0Je7CABL9p
VrHkWZzRg/qozg7yFqljre9/TfWJ9o2f0lgTLlz8a+ZptmcDoJs04IXTejksWgmiZO5GBtSz2gGT
Mi5Ql1CIfMNyW8P9rSgytAQBqC/jUnHcRLrJFqH+D1Pt/Z7UWJn0JwPLu69N1eESrOJ6CzOh3Q21
MKxiYaQ0QJ9d+jDAJiOXB9Ajtc8NcETHbyu6KUfFGYrZ7NOv6cYFq9tvlUZZ11Lwe0R0qjjH7xqO
19ehsg6kgubq/svxRXoK903B2XP5PWMY+e+Ghsslfnt1Xvg29vHOMBvvo2XzLuiYT84BHAIPjm5v
EKwIJ42yLiE+PmujvvdpLAKECHJnBRoo9a0mopDGD0Acfw/zP5VVhJVW0MQ1sp/A2zeBE+KNy7RF
C95+5bwYRVWaDY1LKsafbVbKrAjmjL6J5ag9r9USfDAMlLj4O/ZV81U9jM0zFw6pcYcW8PlfdA4v
oD3h0JlYa90UwIZbqFoLh4EU0nUmIgxPZeb9vbpO0KIgwjgMScuvv6NtaUQ5MJOBOy6IclhylpZL
j/+kDo08yTeV1H+oHQKVEtp5E9fkNFlDKE9l0NqhpNPIy9cx3oKOgTnEKSXTV3OyCmxRpLDpWBHF
/ktmhcEdbwjjo3A507ulKlngYgsoCIuQMqylksvOJH5ZqOQjU76RiUiuXfPFS5FVOHFSVpCF9g3c
2OEcATqt53pnQ8QelRIhS1PUxrr3+Cgpl1T8/wP3eyL6InoT6Xddmrsp+kaxjmQUfSsuNReHQ2DP
KOwxLjhvF49I2qHF3hiuHf2F7NMKOS8ak28F4EKbB3JAKOG+63WxDxIOHDbYFeA7GLbdbp9yR3Qc
2QE3LalhXc2BqyjpxLdyanveIIr/t5A+MLJVnH35gwjJibjkGDgye35xGaaGzku9fv2U3VckJXnb
D8hZs2UIx8uUgGtucIRpEwcEUNp2TdQVNX38nmSxWSUEOBSJ7scznGjb4dP94hwB4m5UNH1sv1Iy
Bpix/Ofev1vWHhZZ66cW4J+eQ8FUXfJK42bxN2iC24IZDitxnFQWQHZ5U+EhtcLJURuMDcDt3Qzv
xa9fIJZWVhYvf82HgSID3EvpoINPxVwEepav6I7QoNx9EW8+znmFnYVC/LHemEB1gN4JZFGK9fRh
T99eOqOnctEzcKW9zW9Dlly3I67uM7Sv1PlffAmp+P74QIbFpKxdH5nZ6NeOuWefjUHf5z43IpQn
FxrTHlzbm5ypaSHD0JuWYOoXAF0mSIjOHHpZE46DyFqB+FLjV93B+NlZd7PvSzVeCQjhoMbmEqL+
ErxDNwst3re9T6epor1rCN8U9BDxYhn0CQxuNcvrhiP9vhaH+qGJZ1WSKGq+7ynB+xJmxwUxuUyY
k7AEqiS2spU5we98JiL9AQ3ZrBngl8rcN1o+/JMjLEda0V6VKBMxwGpvTdyMz5DeEKPaRQCvdNj4
rCivl7lob4j8SjaU++fsPJqWspCv5CIs/c6nY62qwk+nLjnZhRCzFKR15A1SOHJE4+WFwqi0zwYo
e8Rc9JprjoLWfz64M8Cn0seC/hJc+8GWp93iQRZysTTX1O5JHOySoyaS0fm6Yz0QQSZkdC+1vXtX
fq7xT2bBkfBKgzaJPPfWmOTbxkqRVcOlXC74Ze6ZbOacTCY2fwslLmLJWOdAg9pmr8BeIH4AmYc/
3bf6SjgajwthpvZ9Kr2g8K70fFOIdcdXSL+xygzpU81Ht6gS3U78U7aQ268nhXnAsc53nKXkADCO
sV0XH5l6ly3FfVZszjtcAn3QL7zT73E/IuwRimn6Vmnw0wfOp48eveANK9i8VL689XprMcdZvFJh
n2KTxPqt7yGJkYz/a56lhlZT3bN0YyBa5JA1VjDwfPeoIzvDbUZ0tAwxHW08HuxJZ5XCwRfoKeJ2
SyRy6BVUi88RN0WkvQG0uOGES1ZZO/bFvUwX9Acl8SR1SchbH0taZlixekI2nmuBTg6CtBI7yy8v
kiPztH0OKhqtaDukGZpOUInGDKsvKrKfPYiJTRi/UasyRO4izI7bLB4/uLifyIST89H97LB8a8Ft
TU7upiRFVqKcj32YEiALwzDg5Ir+0qMJ5TrYnT1z1p3WDTBArahxKav4nl1G1ezaLDbGK8u8vZni
NfYczksze8HNk++3e2WE8+EofBIHXA15hHZTL+H86dEJCJP6+7hqZdV1jB+YhTHJCpm8r0ZsrAyw
Jc7Raj9VNdbvHk5dJzIK2TuT0/jgn9jz0DKS7k8eQ0CCA7LBG6DbuNcG5Tbw6bApCMa6h9I3oFZM
W3LEGiiGIQSBIwNmyWulIVoaEPl7MutqjcaWVc5d4n5cjXcpFZRnc4pSLLGpTs5QKvLtVV6Yj80z
CiEk6NILUgbg1beQEQVbJGdK0TsbS0hNArd29tLKXGWTn8zUxtEe9KShS7DBXScjXaBcAxhNzVPX
/1bM6r+J5NvK9ERs6Hc0nrEwh82AO1CmE3byGbY4Rq5giUQ4Nn54cexwAur0ULwZJoSU5cCW8mo+
Ir7wgwFQxkZK/ms4Qpv4qDcgvqsElb5EAdK5HiE2AbWw3GAFxhvNN80tFhSx5H1ZcGspABmaM1yZ
ds+CYQspbITuIKrfBaH1XxsDEwB3hOVRjLR+jazc/F2malyOWoKVR53q2iU+1zgeCHlx7Z15Lzs0
XKcsBokpkxX7r4ij/I9GeXjNIyr6ODTjW4Xw74hCSfjK5Hbiu1Dso2twRpjBrid2yR8BIQlWKcpG
V517UuZ4E7+pptVJLGbUK/o0VmG90fl0MWFzv8Z803dstcm9FThxAcmlkV113OfXVb6zar/+citz
jj7asWx/P9Knfh6tnlaLaBdNImJ1RwM4BWTLqEDALwYfr7ZyM2CawivqchyKDUp+vOJEfrf/d8Q8
itRPwLkX84eOSQlqpQR87E3fkYemqQS2hLueQoLIF3wjG/1EgD0+Vc3xSodmgGIneLfaFCswht3B
jHzqWR1exfexdjuoh0/PI473m2r232JSMXeBBUlOCgLD4DOCb1zcjqT69/u1KYgVfbRlXXjFgfvF
LbaGLKLmeO4Pc5Ll3XMpGlU31ibHKywyJRZNFtT4xxkUeOMJBbQ2WuRzRyv/C9xBG22/W/ms37IH
YJUO/T2kyCLuLZL7bkfzheFFHf/XF/9v+KltNB7zAJ3oTvi/0fyQfILNxAoMdFn2DK2uvRSvXc3V
sBc5f038zxw4wPqZXj4Owi/p7eQpTSSGdbacFhliejTQ7IGD99RfJ5d4HeThbd2Wbz+p92P9z5sT
8DwT8+ppzoFVVvzj0V/x4+nyUg6LkjohOQO8d7T5wcVRG0aaiSMu6wlYgY0gSecZfu0gMiiGKCSn
PcQcdOHe3ZgDTjx4stRy3C9bCTHCSNlZxe3PlfKbVruMEgtdyIBnV73Nh28vmTfhTasJWZA29zEB
xebn6PoXkY51OSC7MG9ptGRgHoH4jL5HqRBWuC3iVHOpOtuMKK+lMD6By9VdHEwl3KnbeVzjjmwM
9kp/NdhXHzo77eXzAVuuu0rizrfw5xyTA+iXF096Li2lGvplO/pQ414Ii51njdlbnBc61BPGrHdJ
4+Ew1w4npyMhQSuMMVvg4P5/9QWRR8Ce9cS4LbAJauBQGItfaRq3sFcpfoKMsOG93lSl5A6SK1XR
8f4dlMZ/yfxSzKfrtfAiqmVUIwl98CuUbsnP5LqoxVVuYRklwVVWMKQsPvaiiSWY1aAD8VJ6jwnj
0cS0Sh222lqOhYpRKxpA5LjIYHNuA79FUJZv2xhm3L2KGmqjpMIyEfz2GXNkK9kL3xOj37g/QeWg
yD1j5tqAcaKC/sf8grOCRupV6zJ+nrfsQGixomdkXJMnMJbe1L0r8gtZItDOFMnsqkcjBiGjV3np
NRHT8Bso9uPvMe9CF1KCoddSteM67uKm79eM230BzqxR9g+m5CDiiKilKvof6dS2uIin3CC/vsIG
hn6R6O7Pjv8RZFnfvPgJqR6/a+MkNApCQJAxOZwM1uT25UN3RSqCMTQbcJs/o3i9Fjh6CU/NwDeR
ymE9uZBTp/zBAEPGXnR4IzlEeba7zxTT4z3GEI6fzLvctE9+8L/RmtXJo1kxrSJq6gNthZl+m/Y3
zj151iOiuSg8N0GPXJObW4lDFw7LgFneTd8owUfq6/vFiBhuaA3w4cF+6wPD9XjkkWn+U8kzZu9a
jUIMR7l79q2Z7mv6m5QUZveJywbEjVjpn5d08WpbzwtslIF/x6SfR2QbJvUt9G/IG3LYGi/L5vsp
BYh48ywhpOEm5EUdCN6HaTjIvZiX4H65+KHMKtGoNbsCcstEE85dryBVG16q6Wn7G/eGidJuqBMh
LmjojS9xHEvXu+K40lXTC+DVgkkOjObiRYhPWrW3O5zvMN+IpFMu4b7oi4wA5GO+e6PU4esdAf36
lAVXNWn14bYTyF5gCoa7E+ku8f+hSYwDVSrzCcDSu5DyqLffh3rd9MoYvIZYpYLR82kWhyPXDl0A
Ij6fcNWj0lnbchAfLBtOml5WhzbWs6kdtWBOLdhtD8LG5oNndJdjvEkfB/wd3EL1pUnfCiGgpWF5
14LPGdP4vRkuVAh8bIsJ/VFfR8IeXcMhvsqtBuTsVhwgmc+etxG0MJCN22jet/Smwb8nH8qJq20j
/gHB/ceiDVaaP5M8sFhmr3A1K2IIPtP2Knh6OvbYs0AgN0VdBx3NnveQAmjDmhPGK4KJIe8Wojrs
a1NtuKrpQjFX6qpJQAtbAg61ZpA2xESmLSX1T3iEJJ4N2Y4uaaQuA8F5/MGojoVUk4Y6/QxXqTWg
7Wpmx2kTf0idRUNTymjKQSzci7NJ4L+kS0SQB5HXzYj27FlRDxNDrKXAovtQ83Dl9c2WM1v2V1ud
Z4/2GOc552tfHoSONoEVpTuIMP2bsJB2KZ1h2Z5kFVYvsrw7aHuMDOuv+/y7HWVQisaaPBuevhtF
xbWHiCCMJGGL2G79Eq0J0TjzPIl/IzJ2wz1Yn84aMnTjBS0AyaqH3jCFPjDjY+mHCrGAWahKgJ3/
jw3PMQ+5PNp/wSz+YRw89cR43aN06909/gwdTGKJIF2TyAIxJYeu/4zGkxWpJ0RWHCGS/BB2qD7m
U0h3OefeowSeBnHi6VCB3iB44ATKdhlLyt2K5QgjMMhsHLLZqHvPecR5bCmug5RwjdkUcwrqtUrx
6ixlK9zknQ2rhyd0zmRdizc/g/MD9eY5DSuRAoN7xA8TTKzUQ5ec8h8SGfLRag4vPAhwDP569KeJ
QhXC+pNNAtcmgYTGevYkW22nhiA19ttVeYWFF/ZcLHMtyzPpuGLHbNAXIsdiwMEgiS7lNjYlEC93
8/MkZ7lhUqoMwX6iuKoDFk4O+VIGsfv5hNvQIDFff13uFkbYX4ymlXoXeT+GpHeDQ8YkB2+W1Ekx
e0rgMb5HBlR2BdvtsoSbvcO1YHki4418d88+chc2xrybiCk4ij/9fRGKJ4LAuQ+On2OfQXEPHhl+
zP1Dz+LJmR8nmwM3TEQxhOK2qyO92GOlb2EQUrsOp0IhG7nHblr3sRb66hisCT/ZoFKI6ZnjQPx5
vQjdkPW7N96at6IoxT3tTY+IowB2gu1F8jIIH9Zo4BX0jdOFaye7IDqsu9Dj9IXXWP4QstNfQTHl
k7TjlIlUTI8lzAlpBAq2ABkRjcbxw9fDRd3j1VeL3o9SH38HvcgnC5pR6z9HSmQLv/bCOqo2QUWb
K/SVzt4VzrZew9qMSvbhpwJE35kr9KOaQEsXaqwhfSus+7zpkTdpBnNoIXog0+TuTE4tMbBcT/5N
evv5FN8DOqQVbFl+9zECtW4nEtbKo7lPuYOAnTLZUXFS2vohD40nCnIqRCB238hL5a8Nkyv3mRfv
CF3wvUM6F7fivi0wowhn/mP7bB9HnsKPjZeyqCT16D+lAvY/RqnUkumAqS99N+fGAKd9WbcCJ4f1
WXY/FvJwyb04SVhscjObFC6BOazpwFNDMnW6oGs99qsYj01fxOBjXVU+tOeXj9stDY4ZCcIulrUG
eN2FJy5I1PrbK5YaXBIMuZFTkaK8AH30z9uTn8iEMvASPCUT0GNWQqqi/ZzTB4dhC8S3fX6wKa3q
bdLfQfrdwSv+O8y8EJCQRgQdviXFJQhuwQFKMoZ7rgrFuG1qcIjuYnYrDRCUKwrptfdZIoLtVD1w
VcC/gzXOXXGeP9aAaY/BTQ4OjggykYJgNleyFz1CPlblI8NEpnwGG9GFP29pz3g9eLcHyxsxKu7U
99eoYwTxDXO70fRkmBs59ixgo/IHNrMKHe0gNzFEIB6W5zyGE4JlgJG/O0uUtYP3dh/nZC3hYHtl
mPAKWvn6YCiNYTRixv11WSRoor1145l6+3RclPnO365XHyGGMkfDkVc8sSafGV+QZgDm5ebV+Gje
t+4d22mIp/n6jqvxAHh4/vydmmuXiawFqII5cfiE5Qk0lxr19ObuBBhuYgiXQiL8+J7NO1qGNMqS
+wKop0FJQIHHdrg5nWLmwqWXZMBOQYj+lG1ZjxFAPNRkh5rqj4L48HQML2kOrKlJedu97QbruZYa
E6MIndr2QlxKoPB4jFD+QXHcAYogFFarh0cYMIIRsOJFNEiqcc74vgrOBvasK0oxlHrcn6WcHyJX
A0JSUSF+AxrP2fefTxyPhXc7R6/vhYNgqAnPYjTwptHLzLZsQR8Xqi0DXmCenSquvklnN9Gjmvcq
cgtyiE4rJybeBMNDc8+AbJC3p3S++T4TMd3L5gec+29zAJQm7p7TBCitpbkLnGtawYovAJFSqC5+
LZxtJFCZ40DB4j+TwVyBSlTMd/TIrCNkNBzFajJ4i0yz2dyR8rApMOwP+80FJ+aEz9i3tY5xk2Ar
wjsZZ1xkwlxNf9exzQXrUQCBqzKzHlxyz9EkwGm+xNCmI5fB+nA9oyhDM5CEbHd4tQXFglJsyq1h
uJftupSpliwctv33AEojfgZOf9JNWrjWf0CVYzU7SvjfgxBW71/bG7Kq4DVOBfpSfCjHiZdljDNz
e40JGn0sSmIaY1GXfaq2XOExZUprpbj5O42vbC3wEuxtE4dFoBkbhaubXw4vZRLkCE8LJ0MXAOYU
Ox+Hw1L0KVhNbQ1kNb5f+vFb4/cDWlgfRnTVrEbaGPkFogTXsi/w+CEzhlbm9csozRXfwNS9dWXG
o8eh1lWJZTMZC6YfhD2riBB+F3pelxQyBRQQLdxBnVgiXBdkghY8Um1zlms8rhmQoxT+eYjdhEaB
/uVAWS6iUXlj1PAU7UhOiXh2D0BoQxGK4CwHeVzMlpOzmEShEz37/ZoNQag/zN17Y0ywuppCDEN+
0brbhRjK1YR757wgXm1a97tT5ZsoR6+jZZFxDi58D8UXsw6Tn0GC4xu/GTpXEoUOsUb3GsatIn2Y
+13QyfGGDwuaaeWuoqQ0h3ME9vT1mmEKeZQm/k7zjjtCKLhTOfHhLU1J1vCR6pSNngV3NQ6UMNTd
Pl0e1qM6KOmTeWkv9RmNnCoISw1poxJYXJOKByoR2VTGlcl6F7iee4sgqb/pJN7s8PNBuK2RmWOY
Sf3Z3Q11T7HFpVPlKy9lH5rY1u7wV4miXhTcFHv0Lpyae2DNZhealM0NtA9J3oZ7brCp1OFPwKwB
hq4RZ1uR203SDjvOtRrZKBovhRP8O0AkpNHLo4e0boVQapLRQnthAxnpfiJdFuarvCJDR22utUg1
QuT4o9uHqMVOVN5HXf2mk5ehmbNTnymsGtG2a56bb8rkc2trHxunJpMVOODSdtf2gv5UFIxNOuuE
M2jEHelaaFBJQbmu1/8VaPca2+55b19HX2t1kKJrOFBWO6+h8TpUnttDOPPCwL5/NZm+XrHknQR4
TnojKvLaHx5fjCGJ7nSqUISMjvC5PwPWwWTdjKI/dkcl5ayVTQZsRjMl9J4gSX6svOSfSlw784Fi
hEwVpBU/XCicXqVCV4VKrMQECKjkrAn09srkX7luNyW8by6RgMewy0NUqQO0wS6f9iEZgxJMG0Kw
kTpUiPZoLJXYZL+c1tdXSah2bsakmpA+7j9LF+D9IRzwxCa48qp7cDRjIcVS1eXMtoPsN93TjBYf
kLc+iEPUrADe3JcBo2eodXm7K5tsTxiLby2Ch1Xv47wtl8a65FfNJkirCwaSMLbE+PE9LOn9ziZO
x3Bp7lWMkpzlDFIXaO2wL4bf/bFp4pV54uErDrF6JGOqDWscWyK2OXHUgwx3TESbxTqKb/5W9MtR
kf/yXVBQNhvjaUFZmJyhEsc/5GFDNfLbgXVq46JTCfD/VFHJuz1ZBNYBjy5hEdVTxJMthLg1za5E
/UQrwcBv9rKVln8pkCngx99KZMq6tpQpvQBBfF8g5wEnluU/9c+ZpG+wnIXWN/zlSEh3xLTc8N02
dehZJJ1/Kv664UpIOgjH2JLVLJ7BvAaOppfqFFlFGYHcm1CQLnrwWMuK5wk11jBTFheOw2hIcOWk
WvB2dA3lY7AOdUnZzEwRww2yqrx+ssXwbNVHXjFP+Xvt5IA2fBTwhJsseoGFKHc5F6/1Uzbp/8bl
/k+FlFzK6VPuHEVh4lRCtR7qQ99MHXzeqEWzYDZ7tSyg4hr618fZwR3IWVmlsDpGkGukQ9cmCD5v
f6LAOaKEAmmEvU57MzPaSTlp+m5okIoMaZ519Lk20TBwKqeassnyJ/vBKjONqJorISOEqzZ1Q7Pe
r8lz0hwGMpDrRnr1lESZ0+KmllY9j80QlFebLRjdGZL+9CmJgQT/tZ0St1oOueaL+Lad1sbhH202
yuAcev4S9a8kMn/fGgSEVDljk7+ir4aZ0HFAUkaxGNZb9b4PmrWZY4qDmwmWjF0B8SvOS23ud/7B
zg6C7rsXS8r8Nlfh1mIeYZ6HjBLmWYADWSVo+DSpt/QmSm5fzeqqAzxhPQJQeuDSsVZPmgV6FvHE
nGJ2ackH7R3hlYG8LxqiSurJMqoA0kQDfHOea4CEYlPnSV7hBr0OI9tVFFQVmUOuGE37V1Nrn7u4
OdHCJfiehthHQwb4qQNgbR5JEvWmFzfiLb/nLA2+bWL+6S05mqnaQaj59GVIGv6E99H0jdT8Tfoe
vKUJKP7STst0bW0GYs2pgSUN6bOVpLqmNT1MdsEE3AxNY7EyEXBx6gJVt4RTbfuVI4zpxUeezQMs
ZJPVK3XwB//zJtQ0ELRshNvyqg8RbZu/WYwGvKuUr0Yd25vt8sxpcbiWzrTwfvs1Ltg8o5aUXUoO
bA2s9NXNgx7yvsxaSY9tZYkNIlrnDXYC9vJhMRkuC348SrTR5VRwUS89gpEMe9SOXXKfucFrnRZT
G4s9yDcvsWgiR12GDB4XkBuDMYLWJfQCJvTGGbgX8he52fpew0rtzB5QUeXVJpT+H8Qn4HTtKLkT
NYq7gyNzKGvTRly61v+515BaLiRcE+r1B0QCW85EF+lrXjcI42fvHoVbICkOhZ4L1HDp81yLAv/Y
mgDxsr08aCRRVbcfuM0yDVow3DC6j+ci6PXb2SMO2eYZSpH+jqpk74BkJjml3o/iYnFTSKOxJenO
dHnZdGOWGi+ScJhjtaii5rOIyV4/jTVxXgMtfyuFqggm7GBu1OTT1zp8YyKdQ5xQkaEZUnCjrBLG
KWFPNZmx3hxPfNZfOs0G94FyOcsKkqRZlgTmKhaMqNUBy0iwKLDRWog/GNSpaxIEYuFv+EoAuzqW
j0YRKmdDSgoYxiV71woeiVUj9JC1659TtJ6UvpSqCK4H7OEwu3V5Jg7U7/ql+U5RMwxEVGbOUuj8
8n5CZdAkL5dgXQ8bR6qYn8YH9+5SWOlKhk3GyRxXu2JRx8fb4bey2OF6tr4GnfYP8LMzrZmKaW5J
M4CHif/Xew2h2FyFF/Ic57BoAkZeLIGQUOhqBYKzZWSoWoUsGd/f67NieERoLA8pVxq01xK3+3MT
X8RN293At+yyXfTYbWNQO/2vVRx+7UIAK1DIqT0gOnfgMOl/ircgOIIc7bK2fYk2LqUnPNZy0kEX
BMNVt/jGg37+BrFh5pCURtOoS63eoaBJOztdb/W75VB068mFIEct/UjcnfOXXlPUI+hNA4Z08ksl
BNXHazY4P1wl4d3nNd8Amrej/DlV2EoNFk+EE/7c8V6po232Mmf/foJRv9o0apJgPha1UrrlhzCA
teGJEAk6Wh/D0RNdK+YhgkGqTQab3o8jd3Yl+gqYRByztXiFGmhXUiJAGlx2ddKvi/8VlIVKCd+T
u6Y++7F2qarq4CtkV7gxNkdCN9zmdRyf9mNhEVz/iTOesr2EmN6JQOU9lEqkgNGmPgNd6O+2w18s
PCQh/+nzII8aP9ZgFzM62nYgubN2NDvpkpeSeEkliCMup8EcKhwYXRTSw1uzFFnJTFFmtH9ztF3j
0PjFE/82OIS1N4iq/Oe/c3H9wxo905chxVvSsYlkEjmU88upTCXkEk9A4IbrGNKbBv5ugs3fLIxo
mdfSPNG6vceivwzpvVXoB9mszMjUBOvZw/2ftWgVIOAKSvQ+PaeZ7NK/0wR1xgOg/TfSRirK8JUe
Wlfgh3pRSkj0zKGZlBCeIK7eLWs62G0VsKD7Yxb5pVoYu1sXSD4EABU3Hsi912LY6F5M6yL4A2ji
TmI8iyipSduPxEAi4F0KZtsXbYnAvNSQ66tiHektFq7yzC8lGlyWSWMUwjSfjnUZJnESOEnyFxIT
2FK1AhalCVBHxzRzxXywSA28TqEEW9W/q9tUUA4Hn6sLNVIoipQ3EstnGEDTz9KEIglHXPEGGsiR
FYMSQpjVklhzaITGfl+vCtSuFJi67t/86kyeNyi4i7M5js3dzhTlyBZ2+bZl/ZA+IR2sdT1uguss
SaDRC2NMdkKOqJ5hlea+Gb3x5il24nRKxZlHLAbpWBdvFYT2VmDEBzmGfrfnyWlRZ/4PBslicoXa
Pg1NGksOCqpuWJmSdQZha/Gm4RRENKKq42xmxi53EX3CSeisZJ7NW0YFgsDFY0zFd7KdhQTs9zr7
DB38KKCfrnlqoi5iWCzoPRD73vCVQ68vkbf5fVCCZajw2BimCN3wb63H4DjkPcDYZef2zKrUmfpH
XcWYdWtK0V3nVbhsKbcUlb52T0PjWVTlbgvru/UXw2l7+t1RbzyoNSSRyoaDSc71NEP4eHdnVsSA
ivl6UIvW7uL140pymMN7Zi1v0S4UQkAU2d54eB2CJRqOydOwozcLVgBZSs2FLs/Fsys+kkpvpcQx
DAin7KUpw0d1MLthFae/7xcl9gVREK4EF0weV/m7pSYXcepFm1h5LMVSbFuADORoiXit9s6ZpOeP
k67mtndGMDwXjkLy4QNdI2n8unarLm29i5NeGQhRudczVZnYvRL5tfXfVpOYDEcD8bZMmBB8NBxv
fZIszIv0fCEQesXi3cknKKw7p60R5f+XbfknxaIVt5y2Pjn+Og+t++jKJ1jN4JE5JJ7ZFxQ6e5Zt
jrdJagq2af1j33+ZWVE+LbYhWZ21CInmkcmdqW0eDO6fy95ZTItOEmtkmNth0FES4F+5RnJI2AyG
WgtONezhYz8c1K8Nzx9U/Wab6v1niHD7kevlkcT64OnmHeGyS0TIQdM/A+UB5Z1jwBNTo4EEgxFU
4lGY3Cs4tyG+qRnp+BGIUriUmlfQ5eqkRUzwmjV6goIHtPk2GuFAfes3RnIlx7SNvNRrXUhPd9JZ
Ue/ShVEigQlTtXesK8q04EzJSDY7kY5JYB6+/HRjifXmCLMGxfKp+Fwo63QDYUSzuUeY6nKjgU0U
D/aB5R8Tvbi0nNIiRrCB3rZy25NvSP3OT5htii8HKScu4wZ+IdrWeCGnKPMxF6iHzeM5olDW4ujJ
DFX+Y3e2Zlfjq3zt2S1Ob3H15WstXgA9A0VMXU/COXN+kbE5AxBBwjIoo2CJyt2ZGWo13K6A84iT
xbp99Ct3vKuvifX2RTeyKsW6hZOYpAMR4ID3wIzPW2GHderbjrmp0NfKCNrpLeE6sI3odFiJIhcB
mzwXTro4WRwfsN1leycGMEaSd2H1YYAuIqqv16P2odvh108D1WZntuv/SI7Rgauz7jCDAtfi6c3k
uP2tHoZ8yrUcOxeN216Gw1TED7DmVe5w/A0C+lJoRxfQiAmgKnl99w+nkeg6ZKKT1DY7bh4Up49F
IH5ewmtJJZEvzSx01cUCMQpe8G5pQozQvqzASdU5+JiYcXyLvDA9WlQs5KnvhzeCeUEMHWdQhY7k
cVh/eEU8zDVHaqzTZTXdvW8OGSy6921+BIGQkcKDI+dEiKioapX8/pRaRuvu2+/18HH5eSIbUZxU
6Kx6etaQ6RFDF79Yl6czmjvlAzMGLp7xN+VJ6zI+EK/g2/riee8+Is/phALB/za4l8WwuGiIr8Zx
tAx3wA54iHFpmogIcEByyBRvT+8K3HEVKJbof95M3OEHYg8cc6Veo8XoTUbMJSuCRiuP7lLYMLMp
9szyXZjj6qwpycS6KLy8Hn5a9fxBGS3VHMuGt3qAGFXX68LeSyhZfO3O90uDDEhWw3t3g9tB2VGm
KupnZlFZq/+7hW2AwpwARgVnQ+nDVIILQ+jt6iFzkVHN6bF04ZT9mjwsx41yaNabEK/np7snW1+Y
pTpUcYR7Evc+80IkBact3MpyT8Ag2ePLf/Dt1RGs1EsVWFakMVT9h8VW1oQpjOx0k/5oRBJ0Qz7F
Du/5DbRgg5PRkQ1SBC2OgneopGM9YXPnCkhIk+4GoK7PE0m7w7guiBxHZ/CLjmFNXWw+DahDYtT5
B9IJVXD96WLQju2mYQE8uUBCBxukF9rMwnhFTFnqOntB0Tif7KrW45fPKm5Y+fTHpGiKxYJ8jH4i
MZWg5KOM8f8WGrHf9rhe0qlu46NkRlKoE5tomqXtG3Spt/h6Zk19Kc072wEfMygB/FTvRPTYn3Mn
9nPTsAvUElqpGcUSSePE9z4zNPQcV1v80s7OvzEqA8HD3/w6a6rH4NG4DN4XRHIYn8xmcvUMnSzw
4BPKLvj4Sw/ODrV4mIkcNVZzOHF9FFzJUK1nvJeHxs9BgS7s3807jhrCgd1FjpRLIJRUlo79DHow
vzp9QWU/UQBAGSkQGZlDueRI5SoN+BDiFuB7K8RYDNQ4CN8dOpT2Qg3+QSQ58iZ9Cbca6rg8ZWNc
bGOVvNWEye5n22r9BkUs7hN6GdfLvmwVJ2ta+hr3xFiz3qaH+PJLqct+0bNAmlsEptjk2elQ9fy5
MUbnFIsniONd9UxUajScNDdzVVRuKIY8Ez6/mw9cU5+Akcgn9Cb3Rb8DoIwZwV2HwfUttiImnywr
NXc9YRzaJpBhynCjw4mRgz3UId0tKxdrKRwBzBBV2NRJEjBcXlb3+4is7TK2xv3rKjxKzIw9fdlC
myfWhYOb1M9KpyH78YgtpiGln4HyxIW5ASxsG1YptcYqyqMWC7W29BxzG2aZME1EPkiu+h+f7DfJ
kBBnn96DlhkxGlYjNzqUF4wa+HPVg5RsEhXw8RpuBHc7DqvocZzcCRygXD7M1RohhnDH83YDnY+k
9Ug/vGVpHvJiR+7UTiqJE8YnUsN/+ituiFY8HT40AZJxWv3WNxIC8FSEirOUJZRSxaFWx/nMJrjQ
ESGHC1B9SUG8TMrtjsXnLLxVR/9pJ0JVxnRadv+2P59eHrTilCddZnbYuLgmHSLraNTYpUCx1Y33
56r1BQ7mBkqBLnh7yGmHyn+XiYifsGCs+XS0fM4N60XQaPkBdMGCvBX5nClqauvol0pS/pb36pQo
d8R1uWoX80IQhwpbRGNzNPuoVHKJ1NvDhpEhziIQTeJCcYQeDmavEK80Om25K16DUXfS+RGWbmYR
Clys5DILWlml3E1lT2Ng2cOWgUjOiussouG9Ov1Sm/0M37yb1H5KcRmkcU68E8ROaBsr+USaKqDs
3S3wxYpQxMylqzOIbfmvVQsVDUhY5aW3/K/95irgMCtLyJaBPwdyY9HblS3JEczMzA9NQ2dH5lCg
xU4dTBoYoV2IE9ZTeaIMN147fMstY59kkCUt4nXpPlYlUSqnJtMvr5B2uzEMbVFoOrKCb6dgPTK3
wVfV1+74SweiGi+RMsYoBEQssYRzZ82tFxyp8shjisbKd0emFsEnCGdjBogvQIOXAUT2VD9nXjTC
KDYsg8ObZBJfj63n7+xG3Os19hHX+1y5DNTOj04S5Qw07Oa7ffmRhBJ2VsBcreZX6TWtgA85Jvkt
ju2oYVIJ73FqnH6xZ/Gk1F5SVXAZuzruqfILF0hszCHzjtQ+9qD/Q3KmaILnMmGoUD68IGKw2vi1
p2JtYvGI/MDFgYayyi3TS9/xevV2z/S0CDT7z/PdQujmkyIHCEFxAPpU1yaRKMgQwzwYYy8+v7bi
3d3ENVB+ABF6V9VKpNrNQ3NtYTVqFDiCYsUwrDr1YtpJ4ZGbQRAJZP93euj27Cclbar2etSQFn5+
rKQPG/UTOqMw4ETCmevRwXubjlf7xsDb5jmtRlyIErNDnlm/mvKBCE2QGRk4mH68I6my8tRCZjqW
JNDymO3vOv3xXbC/LkC/fA4mNyoy7fpcAe4OIt+vCAhU7C/EOF95nV9yi6bymymTGD0lg9DC194q
xpK5Oi06DHzJAuFz6lg+GAahLFNGfEcK5qezJR7OkuwT8cxQc6Jy1BGgz8H3chzX/zhrBX6NwVWe
AifjUgIe0TyJvxVwCkzegqOapMPUk3UD7pscJE7yuHXFk2Bu/PcIcp37DQ7RQq7ebJFiFMvjCNFh
+UR0jmNkQMoPCtjXyN+mwN5TubMkpoMkikxxO8N2yjO2mqToVVztDxggfNzurZ6W6FpEyyc1I6EX
h2CbiBCPQ0yKZAl7WixZ4E3Ld1xR2kAQazyA2mF2pnoR07MC9gWxgX7nlDefd/5O4f320Sl5SQVk
lwEUbKPwZa71ASPkgfTVP+n0Ph+v2cG13LIG9s13vmk9WqAAn08c0VgsYO2Zgh9dZ94tQfcJimfH
pCbaZZ4Rpj03BSZHDMOrzMu14KL2k1FMOBTAAgmv+2G/YxJrEOwNH4Owk6CENnkAU3e/2Xpycboy
I8Kp95GPYfRzmXhF2rT79zW86Bv1fAFlQlpk4Tht31AbVVlUo+PKfYMdO+Tghl4NA1omaZselEfv
vGp++o0aI7Ul35XXUZ+5K6ta60LPCBeCmMQLuT1ZiKLmHgNTnptVe9B9UQ1S0ZWp9KiKT1J03/CF
j5pTVfjRqycx/PDNwAyBPVTwbFJU0/lcxTu9hCltz14eqUYBddNFpwqI2u1Z7unAdqGtsTUqbkwZ
4HNPelKNtUgEJVK7o3mzVzZMJ55/X07dpHS2r7LYJU1iaUINDB5NXXkAD67p++cDjPD0tJA9TBNa
u39pHnEqfyUekEQDII2mM447E5TkAK3HHuKSejVF/MT+ee0fu1lJQ3XNTtIWwpYQ5rX3/44RGk5Y
M4sj9LQGcUaOirtVRYDN6mETPTqpNzROA8Ph5MbRBSffLqCiqynf8rDKQ36nhPbXuav2CJRtCRdL
jd/40vaAwjj4on4lHtiZJ4/80HCyseaptX6jHtDBN6nHEZZ7fx3D3Y31Dukk+zEqBqKtj9lvhSTi
of6AAmow2+Rcs1gIT9ifzzwd4nqXqv+IbyDqr1Py0g5bZQVcrT/ZDUIlE7JiYYK5SlLnfSNfoBdv
k/5KvshMuOb5TDK/r9zdLO7e/bWlnRgYQmV/C2Oojfdx2Ln0pqKv60ocn7Ztx9c2Ow6A9SQAAHr9
1yhWcNLMb/r5Z3m6oJ/Q8aA77NO49LX9g705uM2GuAKnbOI3R/X2QPgPCD1xWg0qG5yir7CnwI7r
l140Y6riPuQUaWWX07SJqHLgDaewue9eUruPrShNsyfXM7rP2yAFKaN0VjWV+hZ8c7jf1r17LUzd
ddEG4hxPcsthpCmv4ZNNuwmVZBtxMWMdFpCFdqltKaYXNKGU2akZAZScdqgh9ea0FloFB0CcC2WJ
0ggphohueySVLty+Y93XaPCR5hAmSAL2Md3xbW/2RcYdBEqLBRUQ0IJiJ2y4is9JxBhRh1zENen3
z7kbQP+DGgmAVtWnr8C+qFiiha/NGYYsBx1mdGbs6dIC0xNH260KKjeY6yCduU4lQ43D8ghUi2S6
97XQA+sNxr51DnglwAnO6nNW2YEdsTTnPQ3rbGLe8QoIa6WzpWfxpRPl5dcSJIBWBhh1tw+nwuU2
4ufHPQ8GLV+vXXqU1CJfpS6Ym9PuYnr3Z4VjCWetWS+5oaWbiNpLQLnQQLAvJXqJ8utQwvSXpOO8
g5GhgBkUbWbVTeL4ZyrHhZHygFS0dFgiwniaXmSclhhu6QVL/EgPD5jO0XGJ0uyfhzaP6IVc2zBZ
5L0nzijX9UqpjQLjTHpRbr87Dce1unYmPA3k/GKq40L85Buxt2GrtBDm6p7nXeAag8qmHF8PJhyi
p6ZLtAhYF37+wBVWUC1FAAyQiJhjP2zagfAXkauV7yjGMkv1c4FanAMNCZYKKhiH+ZN1Lr6dV3aZ
o0YVOw6MqYvnebzWFJwgjQtrbkcFvN14nGEALH1VzLWOWELoY2bD/5y3vVZWSaf3N1vI8WFITYOw
EE3+WtyWz1DYALveVi3BYtyYCZiRv3KyMpWw3QoLabEXo+n4rI+wZ9CEtcWJjbl2Nrax24qfRo1O
NpdFo7GWA/HI6PYgccLchFDL4Jn+6uUBHSEKCpIc9UyYwcTH0awjtNN7SDXsPsoq2ILRpJ9DDMKn
YpUk4P4EYHalSXA0bl6D2o6ymJtIPDxlgMh5fKndv7PPugk//xorvDclfgdyOt0Wga7Ve2MyF2OD
qAh8xdmxTLbmqq8eQswhmI62GhFFWw5M/jgepr1tQ/JJB4ktw3wVFa0S7P5r6BezhZH/W7W6L1LS
Jm2NCXHm6pK+C24Nfu/gNOThSYNJyBYk8NuAYrJXulSVLQzfGHt9gnR7QTYD/s62NmuTO/LOV7A8
AIWm1Ky3Jm21oiaFkGum0LQG2P830WYqliYYkDQ8Uucrr900ILo78Wr0P8sjEnu2aOmSI1cJ4Jwr
mskZunIVR2yphHojy/xTIyM4WgdSLn/ce2ICaNQf0iW8U3anL4UdcAU9+aWStfki9tWI4zLSjVN5
PLaTvyQtFlmfMjx2p0tK0NSjfMZye9ApGdcDENW7QGnamHoXUKhOFiFWc9BtXEw1gWdvZNOqfXwb
PAZGF+vmcvErlKU/eALs3eYhD/42b+mTOxCIISAz7+KcCa3PK2/ntsL1fkhhRZLM6PKBcjITVu8B
3MorF57vAcBN/xhqU3wQhNuZZ2OTNv3aF4kF9vtAbyU/U4eJ+/Hjn2YGL+YLROy4nqT6Q7jOPBrC
PnTG5+Won6Uoy4U1PXj0Eru/LeBVVRwfc+t6T+/6wrWGJBAWZdfQgQDdoBpxc80FGVNVgbJuwti+
AEzu724tgeltXWL6lMuroJ1E40CCt1GVO1hzrMlX4QjU32NVwVInIBRYdlAEOIfpt4y+aDrW25Gr
FmheUR9h3pk6QmLduCoZ1vf8BYZjTXLOYj5yBEhN028D+lqj51Emj+Av8Zw3pcXIKiMejHD7vk02
uRMoE2O8dvWy51pIow7tY3p71wydVv13mKxZoEBhwpkrQ+ax2URNePvUNgaHdZpSKWb0fRvFJnhf
iHcIsh9Gypaqo4Qr8iq3YaIRSCqDCnsWp4oTgzrD9rA3LC+7ip9PjW2rDwk7j2VJodvCqm5y4PLY
vWS6c4WNMX+EIP76cTdpvlpLL8BK2EjX9gcvuyd3xcewg7LdfdiwiFvd4OuH9WXIIwNRhaNvvuS7
bUOhMHp9j2Le1IWK49/tEjlNeGqZraF1O/NIGxxsQ700V3JwHCtd5sRxxUjpvgOeUzZr4U7WEgaX
eXw4N/ZZ40mvrUfL3+CgLlhYwma8lt786YY3piLbLUfqtXgSSNwdUxz2ROBYouT5txxJaAOqHEK4
hWD0HpiSlXwTgsaWSWtVcOioX/Y8cRwnx9LWiBQ8vhNg6tFSxhgPaeFXjnYJYjWvof/6n9My7glw
d01+e4MV1n6doTX+wnK/BZ46k4NILKjZ4GqWHoiXM0UeAuk7lWPAMzcJpc/Ch1PcL3z43C6BdRYx
pxpEQtShyGEieNRVmxV0VCSG4JZsxLlUOcYtJIL1d8byFe/HofRY4LD8wag9ySw+w6GRcWFSN/Lm
tYRiREtzxcKuTn0SaZaPvUsrL/pcJF5xVYi+7ca8k7x96Z77yI3yIduv4GCFa3MDqdEL+l86XFGk
F0F7nLp0C+jTDrtxbbw9STAzp0rAl4DkWtiOpbV3mEylmMH3tx9PhAlm54694mAeygVk9BYnKylL
0ri9lWwXPSzvmMqOxzYyiikLqL3nB7YsNVN/GXNibt6EXj6z3JDCVVIxwT58WJJg7msg/O2dHYuS
XZ5Z2BzTY5vtP5dbCDfQqydfH3NM3ssGybaZDVmFCSHJsKO7Kg5BIwCmN5yjvI9yqyzuggcsyKng
XJHQUqjuDjGyqnsU4f6iJfVDWJpmLNI1i9yr2ttRp6QtW3M4HyC1IGGyYYD/Tc9zUlzayn21WY/G
xwwNa6GCpYPmhvqpLCQ0ZWRkXPIfaKs7JPglfmeNYhDZ4hmNGkB/OoQrJf5nE+IxZv1qf0fyVrUZ
cYWZiWFlYlaA0CPJB3DFHwD4tFgqY9i67rPRO34n0gd9ucTqXq7UjArcIv/xIVMsrRMrhn2mRlLL
inX3RaQPfV6g4+v/h8fUloMjugHUhYAK+7F4v0IdtdVeGff3d2vXFYkbpf7vFLnH3DhEG+ijaES5
iUEwHgO1aEW5n1mI0mOpyOCQKLhYi7JJVzXY0g2j9Lnqjs143xonJc6AFYDv/uxyZcFFjVkvaYVo
UHp1BResZmfmbdjz8B/9tKBxABlEp5G8+6gcpQf4ZBwIhsJCZMopTfD9uqSBht5+t+XYdYrnNU0W
gBpzcIMUapzHUbN4hCTafvzlblgUeClzljjkI7wR4KxRN52UdEIFX+2WQQkSP6cQs1865rU+j6pH
OBKm06KH/si+FyXftQ3I4SUbxiFeQzc25NxN/vORrmNjf7/hRshhb0/S08PzKDWSxpzcpfPvlJaL
B5n25ETT5bqv3Q5sahvaTihfm08rbMo3Gb74y1Fzqe2aJPmXpfzKIp7NlS0gleaMNVuw/+28A/sH
N0Y0KStJW2fpyI1PpgxYvWbXyioJOcNsQX77+pPr0Pw1TUAnNDQueQoSyuZ/wQfTr0U2Pe/a/DS+
gZEcCSIjEbhiQDLxPxyYz1e7NIP6X8N+qqHTB8nzy+bj/JOepR4Q8iHOz547pLeZBPvp1u8qoIGV
iv+VXS0tckgKKz8EYjPblQBBqQbrwlMurOL7UfV5WKlqaxq3fL10JobH4YPxCQR0jCrrit5G66xx
2XkXLxmscGVVaRZpus4Jm9+PALeKNyhXgeSw4wjc/oYRzsoBCXvXyGwsWLwY+N0zkUW6Yp83r5+0
pOqjIFkUq9cuDu+Qvyi2Wj+tB7bAlxoADqhF28APFuYOLuFXGeSliKAGv0fmYU0ZtmW0Ow5oDEJY
3vtrzlW8b3iBdOE4JK+2sFmaFBCwhVh8MISU5yMgVs4tjedmrhyojy2hrD9pJozlTAk8nZ6JvFNv
Z5zKCnbrKO2fAgTbUoccrh2ECQ3WQxzNu2YcqUYJLB21V1pyHxDJYIwMBzKZKnqKu/L+1ePLf64h
mIOGcd5fYH+1YknKwDAiRPMZpRjQicKvY/hdrC9tgBAoxFO9O9LhUHA1grokGtHAcgqK2mzzFLOv
3W7eqXwsec1oUPGYuYA42Xx4eJp7fC0OCUBMxBF4SeZEQOJPEGCAly0C91D9HOpLpRI5uApQ0Kv3
oeOBTK+jK9UtyihXvUbdCWs/ulqUODzzU7hfJMAHE8cA+dtiHMuzplp78TRlcdpLHzq6ktSUBEDw
637vQZaRjz9HFOIPaNIuoVuFY9imjciCBj9jON+zu0IkH7aad6/j84F4AaLoG6Bu39DjD9Q/qcRS
iizJ7B7VLS8/Zl2AcUHnWYEMNDiyCxXdpdzcRjTE5rMyjBD460KXONdoOn0eLtCK3hGzVNEGLin4
x/zFji0EBgzxIuKh3L+ILl2pk7ZUsOmNhPD7Q6oOJ2pNxDs693msQJ71qYWjGAwtPMTJaWscBLM/
2m31kYIV3wj0qydBB2kn/iTXNS3SBoT0mmZNnbV4Yg3ZNMdX0Qs3K8wOmjH+pVId2ZoUevaiLM/H
v1Wq0XTNropztbzF9T4n/XpN8XU1VB+CelHEKq/uTNBPnWe4zl7rVW0caboiuz+IqDgRx0b4FiCP
rl44Xe8cDi4Ya0XuyFGBJ0zd3ajeGXV1fVJGnRBrDJyCjeyzseLuMcz6fPRypFv0cQ2FEX2YMkCu
3tQG1eQ4whJgYJOvUWSCBYpeyWGjZTX0q2OSqhIY42pqNJNs+vb4SiSfwzhm4ywoMEa2AsRmRz36
FPgl5GbMRqDunTHmUOyEhZdTURLts8U6wBQEoErMmNAHPIUEzdpPmA7ffwOkbsVcCoNZQaPtRn33
3+us/k2Dl23g1v71XrH/hbGFR0DUH9+kN0LVmop15QUqu4z3Ji6duKftyc2hT6wxVhuA/vTivq1Z
HV7pERyrcwEw6m7fXm3OPDNNeGzn5SVukRiJueEdAE+0lJ8ZW7RBpqBk4U04tB853OJjG1Hc5dPC
r1l0miqmlzLaq4lxG2Rm6h559iRvK9gVtedRHNwP9AQsgfeOzN0/13wvs+KZEM2qHkptrYUcPDK3
p0Cscjba4lQBrmllJE/5HiLunP03+gVSbd7igWTp8ebco5PP4Ql7stXMtvvu+jz74cxOywIosbdS
IvSGG43AeLc3A43GFW/HNWPZbxG+GdTKifIVOy7O87Pjf9DqluuyjINJtYn6RmQZd/mXkW07D6IZ
BY5Y0kRvujB4wMAk7nkVmSOfMhMTgipZq0xoeCBbg+5+UT4KLRz4EqikDHIf+gAvSx3ebI26uxtJ
z6xx5DusTApIKEatMvjPorm+HYzxnJWPM9GBxAk8Bpq3UybUNTgLWCCXWsmt5MvPR30pMd7adU97
DGm5tADTe4kRD+Y5cxcQ9zq2T4dKCaaghmRZ6bE2OdcE1v5Bk4gh7kjvKfIXt4QKDEAZhSkZTws6
g3TiAlO1MOTYuR9dtOVcwN2hZ1+ScMr3OGmavhuQA1KIt6vXhF56lJ+9OjTSvVf6mWctBN73bQA+
aZID5gVyP49MWTk1uNBr/yCQKIY4XSkvl+4ZcgYHaQhJN9dtZdwKYj62909S3gw8a1WP5ZMGvCIu
x4Zl1T00qV1FSkP0UoJJG/pLY49x+IwoMmYzc25ksy0fYIEmokbie/4dSv3lV0TH63azJhxCIiYl
wYYfxXWoOOZUz7OInHZUnjVCEZNzn4juqG+Uj7uhKe9c4xgeNr/wew6l44YXoLT+j71jZ3XdWzys
fygUNnKlZ9rcV2txDgiapou2GjtVQ/pMHzry1cgZWwMefOVn2D5vc85DsC+JTLj1sJoBR8hapkwa
GD+qpSYgOczVe5WTplmmMo3z5mpv3cWtuMQ+X9gDXzT0RBDRLxMo4lpuI4jq31AzoUvlO9hVxud2
X5zmCnnZGBWWXOFPMdxVr8X3YCL57smHuJOnJO4uGDy9s7/Ml7+QAtsXpKBAhIQ+lrNbVBXvGQX6
aOwfdINgQO7OpW/2pNq5vp06AXwOhV4awqOiT4QIKoGgNJL60E4yNfEUkSFPWqcmcYCTXUqAVH6y
R2v1+oBjq/GSGUGXdUtJhbIv1SWNNcEEeazpMxKbb7bdNn7hTGerIM/8175o53zsRcqWoakja5G4
vmeq0hLqdDw59TeiGee+OuTS2MVqohCl6Qmj5oEDJKe5CSaFtSLicBy3rd+ps9btX5xUslzDPpda
dmowaonOcN/fyCRSwbR27NgxfdQifgHPYDv+cizuuGTAcb+8V/uvcoNyB4cBcJG1uBb4tQz3YXXe
kRSDqFGlhzNDN8yDzR6Ha9lpD647ne3MDa//l1A6Ibxz7H+wvNkO0X+7iM4qLz1GSn+5wImeKwU+
YHTv6B6Pa7Q42KidJcg3EVD04Fsy4izhPu4exNZWoZBoTztGQfDbf+JASauFzvxXxnKS/7znnIiZ
26y0gdTGkMk6A+yXCURQ2Myn5dUxw3R5y/aJMWzXRMEhAiYNByc1pfkDIMOC1Z8VFfaJHp4UTya4
nt9huslxoGoy7i+/twtHahkOu6X7xo9V0zwMHbt1h1JY8wkzjmuH+O4Yo1+z3E84NXcsliHrBRr+
+Zk3Cbd5AhD5cVY4PRFFtu91ap2p5kIHy3hwWjYSSAdyWlZcg/FrOqFR6W8JYsdFBpIT8B9FBTmC
9LMQRBEXjnnGX11uejFW+I0C+89zoTxV6NJW5tg/swTXO1dqvbr6tganHxq3OcS/xthKpYY66yWr
aEYkicUW2e15akoaQ2uUEcpiNK79O3VjPzBOKmtXQcMpnRwjMkJo4k86axgnJByAc0akp2KE7Rgh
D6nRNYogOhEYCavisncJ1DP604gXdZBHAcyyl1eimiLCEfZWL407nz/hs6/J1cqU+RKItjp7PM0f
re9Dt31rR2wzSrUWxNeRKWsLRnK8sIEqAADzziSa2jIcqyDBn4qBdCQMn/XuyBRHJWPaTT92WtMU
GTRvMjuW6HsbLmBjCyS9IYuTLICAvF48bqY+XyzhFPCKOSOkFZbsPcOJft5uoOpq1xpKjspo5eP+
LPkwDX7l8f1+/9B11+A+CFQ+4JkgJPoe3wTWTmNE4svRdqjSSv8a4GvS7ZomYXkPaoex+KDsG9Mi
EcIMaK63FR8OgNHikkSZSgUF5kNjwEjsbPhMttSg3SK6Lw2z7AzC2UicOgcfkjZc0gc6pIGM7snC
9pz41svXjKCiOEBb1HgFzQ2JcmZiT8QGdXUDw3Yj277/5MSQrxYdJiYDK8f193MsXahRTIhn/4Yp
IeEgsYlt7U0bvwO6SjCrUQcFR8Uv0ehkA7xG5W6t9026kmFO3ghvcL7qo5bz5q0S5pULtESZxe8X
xGUSpk3LlWiO84iqNQckSN8SmOffRVctWzBtbmiEJ1GfSapsCmsH8UcElQZ11DRG1ElzTqqQMl2N
3aF+6jyAXDoNwHlQtei/+bxm5yQaMthg/DrBZKYetiX39bW5eZ6XZ75mlo86SXvGEbMoTpQcyhHA
Vl6MLTQmbblYszFvk5LvQe9oYED2qR+C/J5XC+xCZJzWXaUPf0EZneOuo1qz/3eDHE94Qv1dJ0JJ
5uUnTdUDwIC1xbyniHqhb5J4ZUJHTFlj7scAoZ+TeSrfAuq1oXrzLanm9gELgjOqGL59z0JBuvue
3H45zGqgonYHbpbqKdjuemsry93XYdWtiehwsAZ9YF+5Yw46Wc1i2jrhwQSvepRMe0eTnPGe4NLn
vVSygS80BBg1AHUTcGjhFh5j4CeHMos6vyoXN/SjaGCeIrPbfHJ8EEvJRP9ghnicHsQ4W1FhcGjG
nFz5UKIfZnr6syP957ZzkcfIwBdYkZBZN4+DJfpGxDHt0SV6emeBhtGDXGU9gv78o//UpA+32e4o
ihJw+FXcsHIh4i4+RkpIgshiTbQaLykLJ4GPeU56YuCxBdMIOwVlslxOBE1KhmL7CKpJv7KQXzF6
ratOZ2ESe38epUP0K02Hq6se27Gu2K252HbHi1WtRpeG+JXHwJoNl4IqDA89vb2/Ex3AlJuoE7ZQ
OLUDntd6dNnxdKs/3hWQQ+HWXGo5uK/7O1vxfsD37CpYfmFPGDB6qM8wGnhcZMG6YDZ0nxcF9KVW
o+8ZbJKq0H4rT0dON+2+p8AKKpCijDjXvki42AqIPga78xe+TRnU3rXsrgxhMQs2aoXkrCJkezFL
sU4UFuxszn9660jCHUG77IppLlrY77oDG0xHcM0JAjSDAWAIBgpWd0WeP5UxM2wLJVU8YLM6c7aB
xhxNk6kROj0L8j0mXH202zFJivkAYSpydY3zG88LL4giyB84RaZhY3wMCsQK9LThJ2eMpLcYSa7G
Cuqa+rBXH5hm6RA43egQXKALwUOBtkDPz4vl2P8c/5MlwYM8LSDpCohfiOQlHEDADniv9VaYrpbC
fU3TBKL0aYTkiMRqwl53RbPP3C8sLTTxNLtKEJKRcm/yZ/mxGoMnyvMj6q0Ef3bxcwUOfRq0Y11f
/EkfVx5osEC85xQluR8HAFhvl++54N8578QWiEzPPy0zX0s81KfNWjfJfRrxMiQ3dyxLHOfwhbJo
R/hY8QTCEcR2OtrxZR7ECYZvnbxsX+KtunJXp7CXXyiddNTiYS8Ajjv7hVB4mxVQ/hXDBn7Cf1ce
379n2gVwdW25r7gk44QAQXoDLLYv7OpRez7znGR+XMk9ZcBDpyk3tOUFJ7SxpjZ6xTxK7AlQffmC
kFN3Zu/biiLaPQO8meYvLXHoboUPOaAZfSoa1zhQ6ZknR6YrO4vmRAWWt+OwzNBmtNRaUFqLnpOY
CK3nwJKwLKBv50nzRK4bx6MH6cidjnC3GjhoTsj7uN/ns99+f/4ElWccCGudIdseUtHK9nVz+n+d
UF8PL+2Qs4HMwsCkZUJ0/IoG5JF5Uh5InC3dCJNjiRudpnaQ51USjlkng2ftk4hqgjMIcVkMLNqT
hSSJdZxYbZmIZQxlI/KtMESHjokNFHm6ZjA9k8k5ACEpvB0QTw3GnSzv29EFuX/vLpvQfNJCG7Lh
Wtb6FjYoRFcNCsP+XpkLnbDmOsoTX5uuUt0I3v65r0FXxoWudlAvsisuIqrelai2QjTcrDJXJSI7
oxOkjVXsrdTRBpsPded/tHXCCcPDP7fdpS1Yrz7svsMNFtmmPRuoPDzdswtfcKRKrXF3lPqc6ouv
EDKAj7ECwaiHjnWDu46G94yo7PouRrzeFy4rcIXYBGYc6SuE4BbdpKwbCAogyb0L8Cl5hYrJ65HK
saPa6UEKhKY4klDL3VqBo+qEujVx/t0N1svYPKZXJoymhWghK7HiiMxXZhgMagxhJlmjhm/nOgV9
Qi5YeaYYqpkGQIsbe26gclamNaYiCCMYr+WS/nba51vLJ5NqJ33lJj0Cyi4psDbHyXDpQUchNW1c
mM+Jz7CFX/ZBwBqaerR5Bgd64jnOrvo9Svifi4q79j+DGiPhe9EECECx+a8LeAfnDvyy1GTK3Pq6
9dUMPyh9ZwSX5k9D8ufa735ot5xYgtgjh6rO+O4b0AHIFCdAUxWyPfoYo5WX7+7+XUis4oLqvHXB
niPmANoLBql1eZTmgbM/CdSNACBgIPQHVUOhpjWU2/GuJOdQG7OLjWhR2CbRht38Ej4ci+zErKVa
IQLCw9XohjB4SRRy0kPZw6eiqafgeZ4nkvGplOzYowpEQSxz1Chjw9tlKntAQBUfwcWg/uIBRyZF
17xLl9Y9+5qei0aTnIvANyZGrxg74CzonL8RLQSg+VdlRx4tyVEamuLtV4hRlK8MqESpBP3QHaII
uRaxYEpCWhDQxXZa8/WKHsw55mENF3fcGBa1n5QSm2dpsgPXyNv7nOnvIc96gXDkdaUGxW4CviCB
/fUea5YChQGr8Zt/WsxD95e6X9hbh5MCiayswQ79RWQfotOsPOPbcepzIfnY5kt7LvHEyCNHjKKn
n6YZxhP+38OP5KTQhZVx1mXug4rsdHJaoPSHaWZARG7YtmE8gxLucSKJr7aojQlvY8pU3kS7qoAv
o5noU8dVA1l/CXPtniqjdTjBioxbJ2VTjESrqsh3PsNhVMo5nHnYT4iJPMp4dzyWmPFVpIfJDur9
UqdLzIIp56tpW6rU6xHCp7bq51VhtX3tsImBKE+znqWH6vCps9f2cEC15h0ktUMVt1ronU86akVv
0g5Kwybh76EHx9BlgxHtCasg04b+qUHgyplvY33kDnujlfbkYHG5rYpDtqjMFIhyXgPwJgEb30li
leip8VtiO14jAMPcfkpKpYSdrpdfh+uSJAaBnf25Aa6yg1fh0pP85h1Y2dM5wKCrcFuagm2SKg9r
SYoSg7MdRNeOjSIoKMLGIp5wUc+5IGBh04/DhGlVDXcP9sf6Js8/KGemkGPVdIVJj/g4m9kYP+zu
+R954a4ekewCGynMRlZdAQv6qV9+jpS7qnBlA1IJtqrTKE0DV2scWAKwTbbPGn9/vkt4OxgEsk60
l3ug9FQ1TPXGg5KB3Wz/WxPExbR7D3F579zQvfF/nLDgG5hrpX7QhxcKh4IH5f5izDR04fvgE05l
N4DTrNELJyrZoBWjLp8fZ/kJ+ZOPPHd3xhz86LAcbYtbO6VPQSNgixMjQzxhWtbSkox0/OZ3Ug92
ha+okt51+0sIdDCmdJxjergQoy1IPz/yTNMbm4TzEDzMg1B0Z88BWEaVXav5rlDA8Cy3IUedrz0x
JaolV8MUjyb5Sieb9i6pMt5simDGjCX8YlxwU17wNcVZNg7/YujepmPTysbExoIkyx6MPGGiRqTU
C/sqbQnPccpa8Yt234s/5MSjUlWphtNd+e0g+W7sqQgmv9lPao2xiMaojujeTzfpk4mfJ+fFNUxV
RIiIDLCJEH+nD+Ny9oYVtv3kACHCYoYb4ICPCo4aq8yGNESOHk44j2cEkb5VF3NNiic5yfdgi8Sk
6hx+jyrFwD5nlkdkovrTNeGphgPMacoX8RQC1WuGECcg8V0eliVlY9mDoI0eCSST9lMrQxVoikCG
esFqSgqk60elJvMEN6f42iSy3YM1FkYwEc9K1M8M5kpJbDUq8mVnwNwvLEfe20KmTZ19mhBUW2tH
w0DVOZqYZFx/Dc1WeaFDU84y5r0mMLW5ieR6zc+L/orMKFqng1f88PvuVuchV731/rOAPjZ2OrTZ
dsZRXQ9ZTTHUL08hb6+4e9vqwivggQcZ59AXSug5zw3tM1rlOYX9NFUzorvL8xjPXEA29rR0LSP8
+HDcuXce1yTJI6VtIMWRzsLYjS9jLlzu4HBRylwc+1q9mRRlisXcZYtTz5eviCY2YJIM0ems9lzB
h9kPMRxKsW2UoDF89/ccgn4vMEyuNuU4WDnyiA/JzmQ+cvdG0+zkQBLVP+nZbbb+QdxCBdIaBaLN
UVCwIU+Mty9dRRuxsfFzn5a43iclT0xpot7HgPhfUcLgEuTaEYYBXX3nQvdbQtBGN1dWz9bIjTvc
0A/lsz6ct/ycAaOfUnNlD3xtZzH1C9KLEuDmqAcKM+NQOxbCpKpXN3S3hKEk0bM7bpnCIqEaJjYl
qlcUtYI5TKbispVXJlgcU2mrlNVuCm5xStjzoaTkaF/8vqKeJVjK5eDpolff5Y79OYSclJAxEBry
q08GkGfjI0Fiz3QckRx4/tgpAXVsk+Lig98d0A7lQXSUwXdQ40l9J2lFmJyitqt4UxeyZ9PbGm9K
UgckoygsjM0tJ0D+5WMDKAgoNlgIUnLIb371Zk8SsoIxwtVvzE7mm491q4E2LzTAdpSKP3PMVGMr
4gOU0W+2TdkEIWbbKvslRKKaM9qLE1qPY2lMCSnKDrINU5wD0S5nAfWANniODrS5qdyoUqkbjYYV
e03DqjR+aFsnRMa1k+ebKfxfsMPwhxu7Hby85EPLQFn7QI6MiFwQjmizW3id2EbYRu//GCxg6381
1cKUVWUSJ/p2xOEF2jq20hoLTELF/v2zOY7WkhXmdIKslUxIkXJdwqsaypZC6V5D51D4LhcAhKg0
DjZKpLt1DzNPuRh+YYjDsdX01cQclal1gOmE7QW3KTHDBdUkWRtkkq9R1WgcVDN+QLRYk29UQK1j
1SF8zC2o3kN9QdgsBAhCOsdsVez0DABLt7pfDXAP0lU5iRMltCz2bZO/hpVO5Pe/KGDHjzAZJsRd
YF3sQ0dvs2TVsL3SbuCZ1HBPExiPSJFGJqHaSGl+EPNlwwHunkjjAdyAC2MpHtJqzCjb3n74pdxi
sPbrWFW8fUCkMt73jqsyCWEwYp7I45OUoO3ERMh00yqMnga838yKghA7GvTeCbDLAJIqmrBtXxvW
blEEVAuLbzLjsRdky3zf0dVXESa+D4svnqaBsRnDrNnp8eUyhqgv58cenM46Wil2b/fBY6lBCXwN
j6PLfPCy3WyEHvq7IMp0o+qnVN+gAU1kfhwQPnrNGeS4yDRH8Z9wGCwwF4/lBon97Bm0tYImBEIw
X2d0xFn6SsmIb/oNzJ1DVwkoAHFSFmq47SjRrKcO6Ynf7F0G/lE9+jzgoMXARWzDM5B/kclB1nlB
WWOVs/ML6d+x74o74ilCztFqPhbQzUz5Q38ChPfczbIWpzr11nNI/hSYfzcwsTPC/FLUZw3a4aqM
SWjUPgX9VwFdWdvED0md/kVF7dU8PygA4Mm66eDzX2KmjP+hFkr5WICpSJMzdGrSfCjWWqUMFYKW
DQOOR4xIM4O+r9rUjl8fY8Qyxzjq2yqzIt+JiPOmaIXD8dxj8y/0CxmXFUvwerG/0/Eb+OK+UdiD
ftMx392agZRqlSuyH9x7oe49KLNP/Qq8GqwnFL0zgxJvvncEwOkAXKrqDmpjDJKk6+M1s0j1lwJf
XwFdYK+1XZVdqMchvKKoRQ0TVsNlTNl+NnU7aSCIqeKSfG82oQZ7nomNhMFdsSeOfaDzJlSizvVK
/XKq8iJnIJkCkhEj6Pk7eTJQyx/eZy9D/PdDgArQvQE94i0WqrsJzgggz6f+XdL4scrKy8NzA1ps
/1hJnYUmSNRESRfqQNHhnZS/KlC0yHU//WNAQMH2Gk3KaqsHLW04j1+EThMuM5+0lNTuDY7CjQQZ
NeMmzokJKCEyP7WPNQPpIAbfR7/8EnGgjuLk95h4KgaVKb7X/hgXM+ifVQ9RlU4KOqyuJWolskxQ
4vI8IrCSb56W2uLj0nOvxaN1k8lIHwS4A9ecmiLTuajvH4HfeiSJjfImbZj0zgvHoT6mYuGJszlX
OyR+9SHagDtleTDH/Iy81kik5Mdp05A163CBxo3rhG4X8kaikElWOW/EriLJ578oeSQ3wQ7mKhRD
BLm1Zembj6R5Ps3TfBLF7muLOAqQ49pFHrLV7dKln6MDd89yqMmbeNZflwlx8PFWt78GKiiW7lxv
oVfheMApJHUvtQ24Rhol4eY1wGIwcmcCuwVNUJS+NPbsstD8K652i6BZPUu7XUkvNabdOKBTjLEZ
1bWHGbBIgnUqFHWq525mIz57XsEDbhvslHvKOmKxJGq7yaFZfVx/nbbv9JWflrJvvJMUWhWmrLbg
99SFDs/Kkj02tyeC5s8jF/Mlb7y1HOKIoc3kXBfX3HTgN8Z++dySAtOQhjr8g9/N0ep66mjOI7Jx
JSBPTNl74OpHRuPwS4aYxiI7woxCm26qNKNqtL5f/kC1UkteAJSgJ0PtkQPrCu6eEynnDPi5eOwA
hdnePxNVM1CzDxXnHUOtC94uQhJBrACZxV5UpuPK8B67yHcWWRk+smscBpyX/X3+nTy3Tx9j/pNI
bIRpEQkIwlME5xfjtueTZ12qQkDkzRmPKs+6iq0SGTBR+fK5WLD9ps+VmzjpFieYZtJP5IqE3TBs
rE2Zbg5CwUkwnDd/XPBspxIrqIiI6+X7Qnl6d5QwV2ID2YYl4hILrcrvjzRYK9/1X2VOVdKs/DVF
NDt0gOIHO+ILlRHa6Lu5K/8iXwhQJUBoMMWz3VFYsz82oi4U6YDnndxiUt3JR43g6Bcxn/LQggJU
zbIwpoDc96B955yTw/2IHnRZWkfBhoCnq1tLaFp+NsEIJoGswiTIfXbMafCifsmQw04IG+VzYpge
BzUOprAQP2cz8KCWl2SFf6w8iH5yBcjB1JCaKoAVMRKvZVv9CMUDAZs+yNWjbp5gXthVM4m+n//B
Canq5tq2iHhE/boh1ilVfHx+b92iD8xFyQ1vyVVJASNAtuNypCXynJL48WtfjSvgXtSazuxqnZp6
cR5vkwv0lY9AK876WaLZ2kMceAxFb9AQ0Gj/6OSYsINcJrnB7LVML0+psYL0YIHiB7OTBuZyix8T
o4ZdcZsnRQLz+eb4/WbCqqsbBHq2pgPAFD4g+epJx06hk9UWTALG7DQKI3Z60FNGRgiJSUS0YPR0
y4a66VQ3q0P+5eLIerT/67RcKptJBT+yVLkzRU0m7ns5MuadFvFrcprNllQkYl1t6lP/TLfGpicT
RRTzBiR0lNco+09hK6Fsgz/KtNwohuT+aJfGe3K7tAFohXW0Kr//fAGKWl5e/YY0Lr+BglLuvmwS
KpIYFuVD6l6AVFpfAakBiK4KeNxr/Or3W6wI1ftVJID3HWeAqo3+eyNqKExE2T5oWM3PgZcHMRrT
paqcoZEoaV8kGtOyAPgl4r0rm1UK1oO3r+fpMJsZABCmflAYB5qGoLFJP8PN0qXdwor/Q7PpHZ3/
jfdMYbBGXjgaexmxax3rm4INJ6cWyIIcYm9xZz9F5WZ1mcUZx31JjoCtZHP/Gh1RWMrnvOne6C/W
As75n6Iibkgw3OGy8IfWUt9rn+Ntcy46hU57BNxunXmaak30SYNqNGoPi7Mxnc3Wiuhk8bhLryD5
yTSzRpVINzQVuikBeWWdNCRzUdLdYKxzd8qGUuNp9pBfP8NFMMFo6LpQJy7lhpUoyQ09GqarZ6vb
pj2HwxYnwlPkg+m10Df90eIncC0Bfsrk8ixT24TMP+cfPVKz90qAsissTYkUXmDpCKvupGsbWEE6
dnDSkg2nMu5KZtc7nualEJC1G1YXt4M1FE8+L/S5pEDmY4bzDYj8LP0MCEj7EVpKWuNUjP3sZN4i
3n0UTbQqpDgz3bckyEqeLFR1XVWV+Eb0aw1eqa8557LajWQXVgibm2MLg9XYzoy1j7QNlaQaFrzw
0r1+JngF5ZXiVpaiN1Oe8ctzXzIhDIs1OMyYbYSkpPjW0y1Oea1dMOGV71xuU6fkeeW8q4SUM+Vu
bo8MQfqEQWHm1aVV4436acKTXTMv0Ug+Vq508N9i2o0F9TngEtIDmRL3EVlyl6pK+iBYxJhMf2S6
ctamQqknD96Yj+7Z0CCzkP+bZYcgHG/l0DF9EZ8OTe5haYun8F5xbFPUSM2pGLkASKETTcfMTt0R
S6BDjQ6zb0SU8ec4VK2ER5dotBsWlIR992/vzYjXt2VSfl6tfpRSzEe3pv5Igiy/8Ewvte57GTUE
VTcjhz50ejpojUnYGaSDNgbrs6jyI8FN8/oW1LM4NTfcTSqlyHrmMEzXBwf+g+pwC7ox12+BQ9/k
EqGl2YG92h5ioKr36heDsdbJVSG0ML/ngnTK+JFn43hn8wf7/vMPSywACsOmWulOIvBr7Fucle30
ZSo9tH/Japx2gMgVsTlCpNTecm0SVKcXwDHsR4Q9VDuj8kbIU5qs43sGb932LhYWMWEP3NUKuZiC
XwXwNbQvI53DI8QeAQ2lnmcbCNshV7jxOjCh+/6UgVoA6cj0ToHCNLUPvcQsV4O4M7ddPo/WVeta
CM1qcxP8sAPgm3LZDqauXyUEJqox5/2vQCcLyLacOnXCem/dp5OA+ijwTaaCljcLEL1zB4Mc8BFx
BWxeHo7A5m/l/+G7INA/uTwxeLo/3VKPV2o+PPeu++VXcy+c9jTURTSodjK4HMGMwoOl6qIpR0v8
DtwajkuNpD0xPor/Ga4Sd/zQU/eh0/6TP1gZU0sPHmBxRF+qwxqLG6k5HAwOk+UkdVPZtZK6o8mP
+fNWS7Bvl69JSqpjUpLYuqxYZTWeExAQ9AqM8kjVuflR5oVdNmEhpG3q0ct1mR7AWH+rYlllSrVx
ULZLWjlRMDQC+E16Z/CbC7pZuyQZRAT0Fq2U/MQf5zWokCKFV+5wUZch8zjDRuSREb2K/fzxhHEO
btylMsPjXsgJ/ei+uiRy+Z70ehxpm8638dpvQemZxe7g4CDX4iZy3afUOQowv82j/gFc8SWjk9NP
0CKBt2BaRXvH5otlGh7NsqFLdQR8Qz9zhGitG31L/yAvQkEh9oUSpaYKnbWPerAOPS8qRAoc6esS
dCqw6sRCo58B7C6APQ0tG2ntL6BTKAW9suuOxLotPLhtCXwJWBfHxUPcK3wdAl7dTWywLiZU+chf
TtScExVioatdK6E3lslrdea2s/4EjW8CuUG9pKEL7Hs5bgGMnDD5hsprDsXi6EuQtHeXzrt1r/fE
7iDow4shHTO1+m/7BX4e63fb1wiGFjuErI9h2DsMjax1MlaYf+V69FCae23lYATG2BZlXsBDbjlr
Lc1X3wTGxss8CrqNOiXzOVMq3CsPICD8MyYt62K/mUU2aQhkJ59Fvs9YXYNrLDFX+rc7djVEjrwy
kUuStzMBMeiQ7NbHTr3JSYuiMKBUddjlfuL9uP+bLiU5jJYqvf7e6sxYc8Cy4jaWac1r83UtNgRl
WuV21jmZ4M0iQDQKPqeT4l8RXY23DJiwtg8wtf77F2ChMZZO3GE+estW1JoSAxqnyCu8mpP0TYfY
0m0Iqcke+fVHIrrgQ54OJPzH/ULRNpq2xHHb9NVXfvycge1W5NNOmV3xcAubv+uqX5xM9sLq4JF8
R/pITS7LnbkhKbCNpThW9bHBGrc+cpNLHvFDSz4LYDbL/I3rJOSg7cIwjT2g+2tWMB9FtiOMt2Wz
PaI78BuPOqdRv8ZbChW4vnK/NkV7S46A3O0Tr9OT89Ri5bOIqpg6eQVtiQirlIwWW0cO3+tQGmfx
GkqGZd9UemSL5clluZL94PdAKYyGP8Mtz/FWEjFh1TgeouWYDa3RoENYuelFtZmZufZdkftUgL0A
g0goCOLw4vJOTb5M7hxo2ZSSQXXrUZLKDHVVxb5fd3KSL6n9t0MNodcPO4OZzJYK6KbXnY8cEX5E
qacfxnEGiJNKHlwUHy52wYvjD1Ea+bM2ap0BjttRRiJ/AoXdbdsFiVJOMrF6NKQBIzqNhaRopUck
K74lMU5NxZakMkEAQXsVIvtdYb9eOEICGIVFOEDYf2LDXJ8q8yvNqzZOVXmEN691xmtiP2DlIzBS
bMCRmIgqQmKaqJAZVr6qyy1qGpMjeomN6eTYc40axRaN56wEHRCrU6Ogoer8HpeMPbl2HeT0qMzs
WKfcS7him1CED1bB4od5vtJ+0IqQdhhA8puJNJVFyvTh+k0oy3ewKoETGknWlkYbkS9HVdsASnAd
iaaib4C8EYlPgMj5Z9AhqM4bZ366m97qc6mV3VBW72KWLL+vJ1Y0DiwRGlvCwmVAWYhGPqh/98Uz
yNLc4PxXt7nGKFSYR+OtsQaf294twfKC1X6avVxXqpM1ISKz7gRpfWevTLQIWhVqIOm8gPF6/T93
LERyVdAGTlLB1eSk2IWg/1c6CvdQI/94WQ2r0lYkMK2ZYfX++E7TEXM5/O7K5C9gCee00X1dNNr8
/4BMgqmfJGLvSv7rAVkEuCx+vUyP54c5vM1UljmqhMtDNGz9iqW1kSEnSJNG/jbYR/aW4vWcYzGf
Xxz67mUeij0Yrr397s2Blo/dC7/1tfl64q6Y2JgUsxbJGpku0hUhbPN5P1Y65ImazMNR3kVOYaW+
t78bpHLC5guqL0qlq/NsjkAagAugTw0iAvmC+Rue86Pi33iOdXgM4IJ9lT7OBeIapC/0icHY2O72
MtgdWIG7NfY8rIAkdDNmugnj67SrRyewKIm0Mt0mrTXhdf+19pE4KDoioq+DMzfQyUQBtruST/6e
qKD3mdI0Hmk2QeyC7UCH9eRQ3KoQgVffx3K2E8eCJVPSa5g+YdMegQFsuUzO+3EgoWPAS5R1fjXQ
bVEidbHRga7Ekb9aR9lBce077gdZQmMHl3K5ANyzYs8SPt1kjkn5SjBp6eAJm6PHHF7PcaYIptog
bR84eDkb7MY3chLRSZ9UuVtbCwriTjPgIbWAAHQK6dB8bitzjV7fnAVm4PBs1/F8rpPSh8ALgUHT
KTsO+pL3mBPNCKFnDpFkBvhYb8gnQFzpmweyR4xTL8K7Qn0taT+blBnykS6LJY50qzPATCVcvEMT
VL7fqjf+JGozzErCivEoHRE0Gu4YzK2FpzNFPKdgD/BtJ/NK754ieE99bCtb50Ad7Y+6uvNfSB7G
qc9+hXO+sHuSYtwkZcbpnzr30YNFpxL26jBEg3PSFQrNFJTKFjje44eg7P54tzVTjtgPe2MQ8jjW
S2Xrru5lzpykicaFQRaMTgMq2TvBQ61ljFRqYlYmTcDGjEd5Qm7QxQjIRWkz657WU6Vz2oCEnXcq
LWbKtbIVdPNk4DJgW8yjWE0wrk/lCxlOSskEoee7U+Miet+sjvz8tPoZngwan/FKjAiqQ3a6/rux
DKv265O9DopwkRJAmHSqm+9YPEWtutVC8OSHgnPrpfoC3cHxWElJ7QUr3fmXymokTzG3eV/fKhc/
P1CH9Bx3IfLEfHuewjf9JHCKDLQI2bzv2BGadrJZQ1Y8ZGvvQl6rGB+XV7D1nCNbb/nAMYfJ/O/P
l2cylRrhcwxXnRI7AUUWlQxaAT7zdfQJGL5HF3QA5n5P1KbHCww1oMXh0mTdLDITKeTwEePkILsj
1552rALjkOwWYLsIUtSnbjruVOJi4kRHnTQFQGEQU3eG0CLU1tMZTq0pK+a/j+HBBO4rS7KDxzcw
cVufDQ3oDB8PXlUijBlVGVaiuMsWXCRFKBaE7r6RMPml4z5xVpAP27gXB+kelpQQq3otcjQ/4Ziu
++i+2V06k9uvKrYa0sGAe2r9yOWBtraNy8MddhuQwxjEu+BRws5qwpXHSj+fJdFdliFey5Jb4edz
k8A2UVmK/WAK7tCN12lc52S1rtEMHuqW8FuAF9IwJPDASVBWMVdRipC9zoQQfZVAPilIO8eEOmHv
Eh1RNThn/vROWenl+fgzvmzKgAdArw4SVbF3abqyS1XU1NnAxR+c5EugJSgkaUYYac8RKvWkU/qJ
orbpSAfhJd77MxYYQbUy/qo8WeRkVvvzdGhnxG5dFU+kt/YVltXHKiv+u+jTdRDV1Ywnvan0i6Na
qsW9s5meiWTyaaxfh9QWDor3QCzSrXvIftGXpicx2BpUXrCSd55COK08tARGapmdIyWwAXNOzV2U
HYpgl/P++Ykkt6qy38NXIVVWh9xjaEXqMLNOyMa3aPL+Nvf+4Shs+nlWK9f+BLz38/8/J0PE1M0Z
ybMr6MD/pnjJMkVow4hAmv+333PO7MtxvjE91yfAJGN1E1+modbTSsY8JUH73q0BitRkvpI7BXbc
4Bri2UxUntWH7bIL2mFJLAsVzzzAOULLhIIDMk2pcVN2yHGKViQGFzghKKPOr+nghuJcDzazoxIQ
oYu9AAjwr2ymPOT6vY0mF6C1m0UsAUGORM0E5jv2f4sb61/hkIPTEp2z4nCQjTZjtYsDZx/J18uM
otkay6xKEtZKuQwygaWDgdY+82lyzVWwEbkzQKLl6/aQAyGqDKfClhvxvMIMCPsdjypiyvvOZuh5
3nS0jvHk4hdyaMcltQhrrSVGXs990FE+d5+LxdAbC6XkTZQRIRGmB4VL78IuVo/MCZwkyCTH5qUL
Ga+0Gp921MHW/PyWgRB6ott3NnR9YSdF0rfPvqn2SpXZIURk+oZBcjZmp0qdrDoNN2w4mAew8qEm
0Zaf4SBLnCLN0zZl4yuQ00YGlQMjHugJWQJzfNY2rK4o21y8kk45vVMndEvZCQjYL9UMQ1Jj7j9Q
FRpu0yy0hNMIF3NPliZyOhYGzG8tDOe1NKfpMnQWHRZHrBMeLswTSZk0MX16/yCs4LgC21/H4S/x
/pfV3d43BjbfnicUmn1w6uM7T5rr+hnnOCpUvD3MigheyFTrKJvPMYrsd81BRkOHrnXHVhwxPerj
IZX7JPPp/LfUhCx74fVbj3E/9QMKDZeHO6x30q04zEk9swNEM15wncIGZBxZjxkpzds1TdHszYAF
tSwIM/q3kp4M20KTRBDZpJp0pZG1isKCwvFOEaPUP75Sf2FRU4RGg6CEIReedCaB0mUuOh/hkwDC
oqRvUzsfv7V9huxOqejsw4Xuva8jC//y4ssihATbVArKgny+6E4g878LY6JthRY7EyhT5sx4iWV2
dKzUri8PvuXAe7t4uhdN5DPB0+277crUdahIVj6lB456MT3OQXFevHnvnb9DrMZ2SQ1Bvkx4Fe00
0JffY7Z99MhhwVzoaxMNwpmTMRAuB1U+MW/FOuP9u8ErhmvKPE9TV2eASDLZ1nVoD2qPl+wvH6C4
EBWw8DT8c69jQo/2u7T42Y3byGoEVFOBAfvpK0xg3K96I/76ExcFeHtBRdfjVIwpEX399o7qrL+c
Ry3I/Orsc5PdOL4563utJiCkC7lY+3beQkzvN/Oe2Fb67IV06L/+3IonIXlalzmdOMEHF9Rr5GIQ
hxnc5iew2Drc+PJ2ZN6lZaByyX3P5NHF2OI9pottX3z24rfQYIV5AqUeaCTFsGc9tORSZsfsNms0
i1s1/NC9PLPVfOaD0tkLFqagaFZrxXImnkCYooEeIBBhVtjILA6cVKMu90CN+ul9q47IPaLv31iT
7rmw+r5oMY/FSIfLy9QqnaIUOkIJMiQ5HgLU6QiNCFdKAdKzne+BD/yR3u/nNBqqlzqRgT2603+o
SXqfz4lS6SjN4XqymXK3EVw7CvuLqR40fukTjLR6UKjbmsLAfOyxrleNR37d7LwL55kW9bxgidcG
sDardhiku5Eofch2H95CrwXt+eNX6tTYBHuQap2Vb+shsCvWtFudWXRMleZq40HtWPcd4AhVKg3U
JBLsuPGOK9cacDY4H9oRTDEGhbZPxVZ4cL2kgS+9laPDxz7YdFP/y5lSxfjNUaabjr3EkAKidA/a
1OhzA0aU2oI0AanqaIREW757ZwdLo+/YOyZ5nmiWAM6B2yTeTzoOx2PfQJ9G5iTNDJ5Aonm3E3gN
HamSvDtQ2qNWbXJofIhGA95plktaq2tL04EjB8Jbx5McoW1koFSiWjY7BMp63GNgYuFke8o2eQ/w
0B0Ec13QhKCx6QzCwkUudzcte8mpEZRUlNoXemba7PWUdDFienOZNw7W+9f/Tl+soyHPD2OOlsct
ui3QJSlZFXQYIg6NOHZZ+yDp4s/PBVGBnOg/+WkCtB008oc6biYqKe8PUuEQiJ8rivOfHL0tfe4n
kZ+lTAopigqGB3q6bAhf24EKDNpXS0/wKwlknpPjZVFdPGwKOmYFe/eeUFH9sZ+/GMpnFYIePhWC
cWHfSl9gieOXcf4u504TTZ54NKSH3lwudZxT845J7ICE/f3F5NvypiTkR4G/s4GkmjU5PNQLKPmw
1xNqFfgo+axArFwJpJ5wb5KyKguwt26TWoryCKWHcxNYMMdy8dxAD1wCbGuVyt7lDPVcpZHmL5DP
6lguGefR74cYPJ6FHF/q6/M4SCxHzIHnFtY0TOwGxeGNY6ecvJGtoEkAKotzdMJAnssrkRjkL/r1
24YEtYOIeLn0cloYXAzCTpn3+RDN+paU3inLLICCA1qkzpbX3urydMuBahukOITjWM9P9n2d3nkU
3OGX41JCCzmmDL6TbVB6VNKqD7IYVQzIdrQHjuQ5ju22mKHM5JRRh+cnK4hRKIODYEaD3xRR9JB9
3wwssy36fcFUuPhzwSq97Mc/t9xhyP9pZoGiZjP1Nl6rgFqkN1sjjyjBY7AMNUUIBTdcM2sNYBFA
vR6ZY9aebseU3xoK2usGHpjE4vPq2kA0WsaaH8sA0nSk+TWEwE2wWri85XsifwqKHPF4+9w3JyN7
/PcGb+wlvDKN5Z7xLutgW69LQ6fawhPhFrCR9pEkk9UZBl3e+ZRuz+XsVewitBmBYzJG4nlPDz/J
OIjhMWyISqXBiD/B4fViHAY8u/hSIIXwy5OcESJIBOOoCkc8MJA90xJj4oc0yjdv4AaRvmY0BhyD
YJdD22krFaEXtehzcDuUAQAKsRx2NNyJ4jyrqwQuriCPwvahFqkDvzzlLqEs92X/ZGKEM/HxtjTF
0fjwV8U0Tf6qWq17DmKMB/VpLf5xiw6564XmsaF0ilCl/8IUlYwEz/3wxbUHqsEsChhGWzhHewOb
6pD+Ynu0Fk6QVfff03VfJLc7vYYx+yOZC13tvvtfPgwDIYHZec7hFRYqOevjJ2mM3wM+X4vY/R7M
bZ5W+jnHLZwdw4uAgoUXuxffECzA/QUM2LfWzz/wFL0U0uBVIl399QDuceeNJ65cMA7nG6rd6rwB
Y7XVqsBwoY6Z//3yWSRFSeOBoZT4IyNz+GgZfOnYaCzhUqR7EroZ63lhBESNkAWRw8Bs1DpfQwdl
ZpPSlk1+jaeqjMWHeeFpRC8vd8MGl/wQHU9zW/+VRztgqloarHg7wIVEx4S1tgknfyQmfxphvoT3
ijnvFngoPkK7k+QCPfcdeDjwiwi/TUqdJHFAMaNeldCGLWxKG9GnU/8gTOa1hjAe6/HqdZpDYFeR
Td9clh939bJL/ycc3q2R06ZWW1wim/qyeLQcEvoSAR7tl4OHkW0B5Fcz0xBeqPoNtmtdZWPH4067
Xno065pn6abN49Kd5nFvAGTaFYM6FRFGl5SuOx5udOOYu7PTsUeVgS7wDz1GMMNn9lB6bogijx0B
BEpKQW9+MMX0pSIp+veWqtEiHehazOV42/oSj0V5v3o9H5oNf1s23w9bl++BEEyLJeC9x19oaPTI
Rx2s+HM9WJ5djLV4wt2UGQ0NLC2Ye3fxKIy5A+/a6hmPRzqe21clftfdOw9LeSkC0G30fAXW6h96
PVhRP77uJvdWpA01cp7E8YJnE/fI+SOj2eCmU1b6/GDMgzHRY2W++W0yZflJR+XUFEbv7m2xZQMm
DSb2zBnMjPR+yDN7Hr4Gt6qoduEycGeKC9oARkacIhuX3ZzVB+MyJsWfCjG2dRQXFQBxIZRq4+97
cGLafRfBbrf4UWeXQsAqi0VxnMVoX0btAPnKlTlq7bENn6eE4zP71ap+s1KU80F6Fj/3urjZHFuU
MZs2yhCKWeeqIq+AV920gfy9C59Bya7pc5OtOq09fRUc5atw0HjSkagM1h6qo5xMxEND4XrvvFkW
HxN/HSy9TdC203hk68dva2z2X6P3gDQf96FRpLyEbh0Hy9ljY05Alloa652lFIukVfHLYbWg2+9m
ET0pXuxW52yHnYJqL9X6D9Zy2WnI6NSKNQOEaUw9qCU56be/znw36x7KFcfIkoe2nIBVUnNMSUxz
+RrE28g7ZQMRL0GYfH4Uj3B7/5Bs3L2CkUmqleZb2UnDmXfz+wHDRMeqU5KCKMZ0YTk7j/T/eqFi
sbwfoLi+1e/cykVk+qr+b3+3eE3Y8apnEzfwHDKKjlBRiSEqiXVjbPzM1FhZPL1m27oWRo8wLQVi
coEXA+Fk9+FPG0fiAGbHUmL/+f4rn84BkcqhABveNQ2zq724ANY0wLe12QwPwSgm9jHcdd1Qf4aW
J/OMRjVxTH4KTMAfAed9jykN1isW0TVvmZscpmdvCBmzq1O3OOAyKoQ+L5zFgZ58UCyqHiuRrEQM
b0uui7SBvaHnVb4nXJFff7fVqCmRna9qZ3iB1BXqvcBXDn/DzSjmx/A20nhwYAFYu9ezPZvdbNCT
fOLDJVnLFyv58hc6mUmA6W1v5qID7ZCxYAjInCAnIc3xxGtkFiR357meFRZdLwfV3uFGj7Yd/MW6
oHlR+BXcmvsecNpBS44z4IussNqFsf7W2rubtLGyVsmSyhOqyv5l48vFv+506KlaZPQrTvNl0kKU
RbfaD4fNhEweIt9Zm1LUL/muFltg52f9LfEI8q4Cdp6SGszVjerpdcInkpDS7otM/cDkBmTG2/b5
3D9gmhHKJXzOIeANXhN7sdzPlz52ZQV2DvLamn0JA8ZZQoayoq5XU7Wjc3HzITbZF56+U7SfHaUO
EcwXZ1Pl34Dd0GMB+tD3myne0bSLAPm/bKNa5cwgVORXMDUhZP6v3ZuWwZphOoIpTdHCVitI3iCN
0L9BclADL8vomjPSP5I+2Zf9RBt7cpriGQ4FWBCA3NHOQjvEJ3HM1xI/osZbbZrFQvMzH0LdBqF7
mBCUmV3z68rWZdwjWDzzV96Anu3suJaOHhDeaM+2OPPEUgtcCiC1TLSWYuqFthDP4W0kHL/mV5jo
YHI28WXgoocROw7EVYcaNprp+ftoaiDZjwVqF7pK0/LENciJeWLy0xXwRTilOQjiiUk5dv/hdX3g
bM1SLrR5W4+6nSm0jBpX4B/39kCD8Z7tTnoZNVYF2i9TIc9ei5n+ivWSJz0SmyAcRTj78Eb0ENzp
7aVWs0YuozFeFiSM9oU1I8bnR7OF07QkZQ9LzmpmLgcFgb4b8EHMwBTnKd2vVVfJf6Hih2Q/6si2
nvNnfQkL2o7Xopq/tL2grtkXkcdFHp9YfZLe0vW7Cpm5MRJoJ8SlHzxTLgm98F5mg1N5NYE18bQH
Qs6/+23oDwPKxa6iVb1/+FZw/ubnojEGwbYy1CJYD9T0U/uafU+Opn+TBQL++p0rTXbONuxQYlNz
y1bqSsus8AMnh9oxJuxiwasx5QK89RcwxSr8QVMxB9jw/fniBilz/1sZlF+LX0YN64aO2TUtFfAS
ikqbL7p2F1QT2T0zM6KUcEsyAbp5tItUsZiOVzjzqAzeAG50ZaVKuik22t0nsKHH9roV3xqpMly9
KVoz1jGDgNXNJI971D+y0W0vcT1Wv0+2H8W/PuZBjz/+6GcHVLbma1nx21rOhc5n0Li6/dh0dDD3
dIil1liRE0RONpGUFW3SOfite9O3wRLM2N+KBYUmpEGcDRa8V+uii7yQ0JQ7vZcqow6Tg1zJiTjz
VBmTqCMBuA1Q06OCXBI+LL4Rf/FxpZ65IqWcbOgIfDpaic1h39X/iSlFgwehbiUzSfD37UupN68U
9EKsbJurk+lQ2OBgP1yNlH/aqJA9c0Q6asnMflfV54zvHN3ETOe+OrNqJXjBro6OesWCZgbfSBqK
Y+QZkGzYNaZuF7OEwwpDyjmrmG64W1Iei+PKrPoFQGza3TT9nCZbuk8oQMqoxxBozosshQvNG1wn
dlTBIx0jCyvsmICqDR0tjDbHSKgyk9IelCN+CQXRHAm/iggZFv+n96FOkKofgbGGsfwyl5JBUK+q
1ibsSf6rtnllUWhTW+g9l34jB+XB2Tc2/ay4RSG/0cWdDvogrIy6Yi95CPH8dW4M82sz3Mf68JX8
NpZlH0eM3t1jYu7um5FdPuzrjoUL6L3S7CgQ8i1m0u9EuKYPt6GZ5UbswnKeM9cQKA5TRiexg/kM
8zF7QFb/CtMOyx4pxo1MUTKmePcKqkJO7gRlby1eeatQhZVTOx0styJZ/mxMokhFZ3N1ceWSn7FH
rJAM315j08PdQiHnW7YIVbi+4gnDPZI2F7SiQxB5xGOe3M+P1ukzaWRnaK6NgRNBBxsp/Eq5EIKS
wedYoGhk8hl/I2cEvshSWBJgZ1YpVkH/BwO2A2iI6/Ood6sLVTYkqmhyBemeuXmNaDaHNiLwv6fl
PR08hKtpA/CCkEFg9KRxacA1vNVtIUngEDDXnBbZBQsFRQOpZpoA1ws2/PyawIFZJBI6PE/iTJ10
/52E0JoM6bX+XmtF3ZC6fcjLqSlrS8NOYjQxaqwDa7RcvfAokaQHG/U0duQQ81vqBQq0f6J1jYKJ
gf9+gonmOj6+HDI94zRXVAOsd3WsfOEuG7ZMFtXzZoKSyKDVe8kSZ8g+7Xc59IdfPntrRyPXlGg3
XH8cNDA16HzPGxDPWjbnsLDFV6kXPFxLYySK4WKyDMiCHALzYZBLgeHW5aNrAZvB9FVevMfU1NOr
dpNxK2f5rhqhWcvfnzcpaH574asech02KURG9jF0m2hEc1a3xo/dG8KVfXMwPTdbiKWQfgp26aFj
kLP8RTP5HxpYPPAEFLhk//RG6Gg0ytJfXQZeR3ckemuE3Iv0Xz6fatDBB9FbIVyOzT/EJNHIkuV9
tLhaNS2GVrvdBCiEsJ6NwNyCxwtdYbUz/LivrC3Zfu0/HOESS4s4tpvZxlqRF14qgIZ9AZRJi6f5
f+kMOH0c/EJbkWGrvFThPwouYZD/mD3zjGe3K0LpAY3t0roNvIpeBUxoBxfah+HfPOVcMLtkra32
NJvnh3I64Qhfy1s+ZVsxTYRApITsndxcEt5PKYG+ucsT+OKZkmUwHLb+fOglwPo56hdhMSYtXlxF
stiFdxq3jNlRoThIZdR1Q/coPhOpYz9Tk95+InBwRXbQLMgxX9gr4Id5062oVfGqGKHN++XBVKgd
3i7ewa1qLwzWYtEkCXSgJuqRVA29W2U4m6XujtHZMmhHEDwf79LG+VtZcZgnn3ukArk+pqjAWn0z
Yaa13YjlwdkNw50weLOfK351vXhkHaCMqPIUPD9rYeIQLBy+XRxCm1rbxwRH2Lb7iu7H68mMXcKO
MOruRLQnXxQ1nhmWSfhN4fVuRltVFh5JCxnwgtTKy0SS6oW4ldAE2cLGARXgR+n8eQvyeuHoCn/i
UZlJqd+bhl/h+BO01dEL2pRgri+HphYEEnf/FGpNuu6dCUOBY90ljCVFruyTOvOt3YueMHZeipV1
vufnxQ/HfEoA65ejUWsjJa5dwc8VguJuik6kNPE37Yrk6qEs+UVlyyXYuagxP0ib0/CZLhrVJE7l
q1gc5rK22JXIEhSRT80c6nIornOnYUnmHDQRdLQRvjipaFOTqF4z+1R2Q8XqutG/Kete4Y2Ht6vB
CkLRl33qXmoJdp5QjgWaZQ9hcxd5bLL50ryLbxbvCqnjVMqGkDwofmYTN5t/2NdSc3Q5x4CFuiSY
R8K/Rs1SU1ksue9IBmtyJbTTia4KrJG1uchMQNBjgLh8oxYHnj3tuumfZKcKpoUZ/A2XltmzsiuJ
qak2nxiiJQMMFFcLMtt5abQ+2l85iMv5lrTcYZ/vOGOXA6k6G1n/Q8ESk/8rZ/72kIlzmmf6XnLu
kz9cv89Cym0Oqkne0doErFz9Zg7i3VLICQFcGKN0GtC6RNLLT7suHIRhkICZ7tW/lCbgOEcRX/SO
sK4vrg6SYgVxAVpJq2u0QoOuwMZE75jCRxnAlMyepJgoVGM8HXI75RBRUEJVQOUFP/4I+fdGQtUk
TMfMX3mfmH1uS41NmMxtYF/kWIrw1spvdcXnHavjSKEzhJSPTPAWLVOz+qc74JcwU+WXUAZ5Puou
D/PLl0PUnjyiu3zrzSnWShxqZ8/2Vx6H1RpFNPV7LQOfFss9hv1b+HxIasAhwex0HOpqkDJK79zj
+Dt9QKrfVE2Ye5e3fcGyYIrqO3NRiA/+ogpWLIKfFdUS1ZzysrSGVhS+MvHn5tN/sg3Du0QznE8o
wKRZMjjv3OWqw0iB7TLkSQxf43eWCJ4+7w75XCnwC3sQR3MvHqPDV9cPTUmEOYkSOF/z2vUJL8uN
p1KFI3GziI/a/bJ4DOQu9i8oJMjPStTdO69ojSpkWc/KBRt9L71uaG+xlKFuIKNcfCZiyQ/xnMx0
j1kCgREgR1U6Xa8iIKor//oHdolDcNfYO5xzAvBcCoPM/z+LitGb/TnWQ4JXYCE7P6g8H73QOp8e
n/DF75N3On3+uAxsypG20wgg+JR1hmFoLbsiOLoQ2yqsw2FhRp7KCEokQYo2mY7LK1JJzljpM8Qt
rn9diZTC+4XVReO9sm0/unnP1odswBz42rux19im6baDMoOloWc3z3auEK+oxvoiNyQeNNx6kpU2
dkbwyvhP3GuTv0WUTozvjwR4JDVJpdjddXQ12K8lK5w3nkv2RamB1tGtsJaj5oVNcUHb8U475v3t
ygXeQtDJTuMWsXKn6zHQZCxBEHA7BuZB/o0H7OdvYbqMSQm3q+D0rELlOUo5NIN1GzAjUkMb57ir
225aBiTfyYWds7gEapt+ibngu0CjoYBng//9oN4KAytz+pzSjbbmFOJAYGKBtKlZnGVqrwP1XQFY
Zc0wh/J92l/ZBMY52gFA71H55HJFLwSAnoFKFDnqRLVP55EfRdaCMF0u2NVukK5/vgbvm+CdhQ+L
QEA9/RJWTLI+feYo090ttMehcQgXIpdX82wpIq9xbMt1TRV5O8uotd1lfGvHlEQL3GDdCTRTkAp8
zJRtAYMl796ccY92Tv57cWeMKEiuOHgNwix/W1hdXbdbmWAYKs9rkKppSA90edHrOb26CKP2Fkac
2BA2Lv8ESAtoSfpD+V3jPiYM1RxBgQJLiGdtgIAAPcTOh028XhIiOqTXPx58LB1DcXs0M9WU0kOw
/HOHIy9nP93r2a4CP6BhksKkORLa+9B3JYiZC9LVDUxsFurbdyD27O41BcG9aiFb37Ccgkmi4m8B
cSQSiiF5BfgYj7grAeCXkV2Mv42tDXCZKJjqHU+poeM2hyPQN6KKtA1CHFRBIpwa14koue0BYnVy
PHu07cOJ70TussFEnRNwpMZK8JMubiGnnGAUjFZ//TuERQSoBGQoxMJ8EWxnxwbH2nDRl5E9rNAx
T3WFeCKm3Al8T4B+XefxwhMMPwYyEyTokYQsZKtkWBfEovY/OiPuZ/u8dWvaXGM2H4fr6VRHhqtI
8EPtH7lgnGvCh4MNBhushp5Dpl1dwDaienRSXYtrIPdOmVUYUM/nMgBYV+eORRkHwtA2IFe9WsMq
6YYdslyBB8gch8sL5qIdpcOo/LM2YMRJd8Doxq2+jja8K0Mix8uv9IHROi4dNWnkKdHSkgjnj+xd
9MEwbMp61qZZONj9k6yrb98Y6xSHUTzqE/2yYS5cOSiYyrks0VkJERZmQV7M0WQvUbFKtNeTyZFK
gG15yEzsBs9+JSiMrqX8MlGa5xOQB894Y7ldwfG3vktR71S1d500SWFyflQLGEiyH3w8hdETlSVI
mcI08CEGfVucp9AOrtDPEKK2ijKOfTVQGPd46eZbwgohl27gjUGSKayi8rpIACL0t3MHM/ojIH04
Fbsd99GcUi1wNnl1KrVgSMaykcK2siygLZNQZiq5S9LMo1jvxt7XPpan0n8qPrWNv3waqLPu1U69
SlPZ7LQrELiuQkUR9T+BZPhbGbPuB/jwqS5G84V4eBdTRux8nBwQX11BOYPbr4Rm9UIyo+1/cPag
8EYF1kujqPCJDcw/BmDZRNSnnhDsavT4WFw7zpJnCO0XU3f6WQ4NqWJg387Oa3EjdQlmO9e3bTVo
IH9m1rc295gYy3EgaHAqssRazJVUxmIPjJ8smTNvXbZJHDC7pmiDoOKu7MCeSV5/nsDBpRZDhsNC
q70R1cioZt55MduoxS+YgQAlEct+QhwoTtDu6rengpzcS4bBkhgxsQ88OoMAytZ3XSHF21HHGG0P
TffzDOUcdrzyL/Wqkaywiwotp1Om7lj0m7ydtv1giunjXkufc5VoydJanzwzzQ1T3Tyn9MeljMIu
I11/gg7TVloEGrlBwVoMpi4MY4q80vvH4TNQAtgfcXrEl6KIUPWEytKXaoQ3AUIFttWqbDOetBGo
Ag+b3GirYQ94QQaJ8sz7DgBFdDUY5ezNB5dVC12Xz92qqbOctXyS5vApLyyc8serXtQhbqNlor2B
U7IRMYQyvuOOunR/+wbaf2YAfPXxGxiZYoFEP4DgWB9hbDczI+uA0PHCAhYUR8h413hTJTN7putw
Du9c2wiJCu7X6r1SrRBH0nnRIG/RdDBz24Zjv9mC1V56cv++FlpyEifDWfeFi5Zwd4MYl59mr6Wr
Fn4JUnY6DlBc6r9Pm9qoIONf4F977fAmmfTT8y4JNUb3vWWkNyPgekZoErE9NJIrwA579cASFZlR
aDXk4iS2vMG16FlFrruyco3ARi57X6j8uZkzGxFTGaMb7GEua6t1fgD7CeKc5Qd74+b4EYdoNmSv
3dylAKwxEQc+cUXRFikzfv5HwPul6vbuLLbhRB/mcGT7WRMNM1+Wus+Ip9FVSjIMN6EPkK6TenSH
CK9gs7/D06D8o4zRcDPHZJgzK7qIR56UmrlIY1jyOmjira2oushGcMAD5qO7LcpM864IvOOhvdGV
nYTinLEDSdmlKzvbcKBZRQIS1IMdkF2BRrjxtG7EvoYY1OT5TxRfqZeiLCAvBtFeWMXkp50HdJHU
GS/vRUsPUL0S0zSx0E1wvklSPgsXPjXS1rCfDlJYQGeFjtSwxEZP3ADEoJAt+DFTG1g/64Hv4jaE
Ait2CHdv9hOuqun2a6/kDD+osD4Y7uSDGbNZ53i/e2lsLNtGtAqxBGe09KnzvpVHEXvvN/spKFiZ
SdjPuzQ6d744NUTHGuPdzQTeJPukTDtLpJP0/ozE72E/S9Uge8QL5YepQZfAEtr+p9gumEAKhT50
CmPF8WCgavLCjNv0odLww62cCbRyuxMBHVkqW74amrhSZjPHkMxNd1SQYflSdke9IzgbsLcZYTvR
P27ue5fnIW6M9xZQm+KjeUwf4MG0UKo5Y2lt/7FjRPnC0bGv0e7vk/m58VjiRL+ocovj2kZg+tlR
sV9gisGM5GXdrXf8DXobdpi0JXT11Ck/u1Z3JHQdMPGJ7xPgHwXVHAxVqIGOaGAsdbhBba0dBzEJ
ks8iGvdDYmVpYEp1MFkMKIIpiIv7tqbetLlQWuhsVwO1D0XOb19RfC7W66Kz3c2JP0IdnZgT1ORz
cYZSeRexdgbHB7XEpLQ9zWXQ+7WMmfYu+n7koRxLojYqPnyIrLh4tBtSlg26yqHhDeoxEfDoGk9A
vzN6XuwaG5YbCL/tMtOXbymVcVx1pbRBB7j3QBfehfraLyW7S7BLip5ZGLN0V2l8TXjcKDP9KJNP
qmoYMZZbPTrmcMdTQ44p4d0XmONAaSRAdPwBlxpD1wSqbu1fp6gS4pMK7uE5zwhZcBuocCwl10AD
Z//QvpGueKO4MbIzL79RNf4oMzXW9n/HSt7F1yOZubnCHVebXlpWHpjAAELUMgCjp7tmI7M1Rnu6
cKTWShlbStYWK1gs0Zb85w2RbBTunfw+L/iZwx/3GmMW6Sh40fIyVMmbtIRH+aOlKq3TLzCZVHPM
sWqEd1/WNxSLabnYnfro6Fha2CINOVBy/IUn3Jg+9dD6/n7kg6ANn6uLH8fSNA4Ko5541xB/QzLh
zK30QIWxlHH3/oVXIM7W13YwCwXsy68fONvoQCQQaR2+hMa+UL4Yqj2bvCX9ezlErT2lJ4NFcrgM
Wk5E16PdmblW1WwXlrFLG9UNoADK2oflm8xP5vGlQjtqwb9NucQuHGQKCyzwB+HtXdVhtHS2sbUP
dsUA811qX3Mc2dmU01RDxCLrLoFZsRSLnl205rvvftInic/i3y+kjKAH/OvucpuYXhOJ7DjPhvpJ
qagXbzu2Wk5f2cs2acaSvZWDiFCTMD4nVsd5xwEHVHJPJOwsxXNYaecqtTIf9YFYAwiw9l0pjT1D
BTwFs+3iLHf406u9/5d2x4F1nLH06yac/VslYgB3rITtfCe+tTNMXuZEshVCBaAjFvQCVG1Kvg9H
gCwUX3sreFC50yEqC7WkW3CN1k15Be/5k7VFNw2NMTBk06VUjfsIf/tGk60uoLO1gfrvXMOgngw3
CH/Cbxs4MzrMXfJlAC1GWsUtY7PGojnLYZPbYJITw/HIJ52XHl5j0FHwdmymF7kmBj2S+nYvLSUH
a91Uc208HvGErPvO4/Q3TVn0TTTaXJyCLSHIX9JeWx+iFBCZTlDBP+Hwm9sQUfCwMkXYi4xhQvWY
8GxQaxJVk4GeoH35TBAQMnSUoMRHlCqTzV/leAX8+n/L/OJvtHM6+Pp8l2I8lr3wGVls4a89BJ+C
+3+a+kG+4tbA8xMHF+Z54Q0hQGfJb+7wDMoBOqSqG/E1ViF5MoYJ2F1roitrQ6M20OpfoHxm/uZI
OwrEtwVdGBz7CwRBJoYwXcv9SsIubfz2vplwXccizA3mAolLEHAerlxIYVTGLQtkOCm8Kwrw03Zk
EWB0CrPMHWwqjJ0tPM41euseGEOb+Z5UEPfC1pNTiM//BmrkyITb7bBfdv1+27jKEksndE4cRRTD
2sROuydDFoRh9q+wbdzix0iwXeLKUwiQyrvjlKW1ThIzQNb+F8CYb/IfAc7W0AsADU2T2xiPIrm5
xBaM30LZ+o0+86DXhswp9kUpTwcHr6EHrUfRXUlDVD/GS85m4q8buwmzQeyHvirFqwBXJ1cg5IWW
3Vl4xDkH3iQ7cFknCBqFZLuSwDAthc1MtJPZglvdy0bRTzhnvi4PbCCRzSPI6jcVnDNUCD0xxQZq
36pZsefICn42BfDFTGAirV1gEPy+uifZQqmy3SCmh24OsW1tpJA6OvANWVfk0TQgUXqLNiOYuWhV
wuzuPl1EZ3OnxhRl5iRIGSuUdiD1RKZTVN+ZDfu7d+wFIle1ilHobWQXLtXrlQW5ChqcqOoSNTMX
ugjtv+YMlSeZ8prkrL+yaYU4+ZufSJoTxN4pQFjFqL2hTfZMLiyZZTGPfm+jcA8ADsHPaEpOEOEm
weMUm4krjiWSyt6mghvOsUiREoSXQOwIBU9ziseIwh3nZ+JxGVMrKRr5giYpTxhLEhaVwm/Wh4L5
upByOZAkZFKl89Lfr+i10WKLl6QXbVrO6SwMn/B8em+pRY34IbGIx3LgfGnjtxwvnX+eyghG6d8R
m9X6HHn8z4z2hf7YqgSsNObOH18Fvx49yzaiAIlKoEcv8yKMiDit6RgaWO6eUgNA3QGWG4yfnWVG
ca8LKPKxHEWOTj2RUcOPo9iOSwVag/Ger2W+k+1/rKjYZecHXxdCvSWfQDHPPkF2USZOhGOcQ29g
bqamWrWbDRIKPEuv41khw7HiGpSISPAesumiH4+BVV/fJyD5JiZ/leU36lJCJGCqlGmo57ynhkC7
TLG76x7RFLeR9A6whZT2eYS3Mj0jBE7dCcmce39MwOI2rGk9QCpZW/jByKi9VFe4aheZdPOxLPqw
dcFfMzT6exreJi0MZ27Y6KKc//otAHBlAp01mcUZcdTJaGTcuW9z3yn0XOkfZ5s0awo8VWfuUnAU
ZkyqQNYy+d1/DBKt6SxdENMuZlvGdwfB+hoS7LAHqEZE8rSZ8lMxPHwyPS6jf/zF2M9JiQYv/wDv
Wphe/Y7xLJBFoMP5hrVuHaQDdlU33SJOEcm3miA4pmQXPyqHZWqECpl/j5N4FPf0UMlsPmjeaz1G
HLNMSdbSVf4kmizXX+QCUwSSLtAkLG7dA6vEHqoLWxa6qLVeN0bkeqFCRgXqfFt1evafevn/fgPj
DyPFev+dO29jiazIJ1MIFNjJukHIqn1iCj9BeRISw5Zlayo9hBM6vl/Ha3WJcYpSAJ9Cq19i20B4
8QcMp7gKN/sQF9fnA8Xtakm4MSii0oLf8qngjqGmZY8D6DyvrdPU7dBTu4r58Yy4QuhQJaP26BMS
5yLnEJ0XiMlqL0IK/YUBHWQD8lIW6/O5R4xYuBOGRYQPhJ+GfNtS/Db9xVb3R81Xh93LLdXLGQYg
G7ytblOaFW7/l4SKI3j/4qaxtP/cJ7kO0A0I0dfUkU39pq/Q3M9WCeERuG1zZCWgaK2EQ1ipl8ti
zLOyZ3Blka4PNJFMR6rXssHH4Ix8McEw0nsdO0UuiugYCnrAt8LUAxJ1WzTVyag2VGbbZeMkoD5c
CBMfyh0lmuGknup6bwaIarPoDd5Kqc+Ye9MJ69cPl3KfGwqS0CPBn4qvKPkk4fJV+55bfADVWCkX
88xb/VfMHXL7tldVTl0DyNl1FYINYSKe7FGeFXrJLbXOCytzlUPpSxXWkytfTZrmjSMdKJ/1UP8R
HPD+t4szWNkaHVzHxkrhzo0qsLm/IiOuHAsdPsyzM+rODr/VyeX0pIiinhLingqgHrOIGKaHyHWr
Xcn3Y7gQ4fuDJBp94COMBle23bn1eHgaGyusm+J6Aw7I04JRIcKWcDF2IhMcCwDW1ijF79rPZEP6
pXZgi7Em3l51bi/DdiYDVCvciwui7alEy0WmlyOsHlzIOGxabenb+LmVPrPGowhzZhCsRkDFq9qt
9bDU1d+Rk5kcxt3Z4f9TentFT36SilrIElOOH1LnsLy1hhnzoJlQ07Yf0UpSRgnD3v4ood9fpUvX
DDm8pzU8CuCKGPKA6QAy6T3TlMROXiB6uajYwafc+0rxpeowy9SGes+Prbp6NzftWc4NI7ft77IA
YHpdf4cWPnn1kINy5vMc3kf8oG68p3gEAzpI+6gpyo3qi3+8SqFwjHN/ML7dYo72fbl6TOGD0y4J
ZOKPQPTUIQoVBix1kOGN3Ovl40QZdVyyLGyd2bjZGtHqZhUJg1ncIJjOr2LsVCAyMvV0u/jXl1VL
Z01JsnP7H7S0Q41YNcyMiWYfOBL5J5ZcMcFsDrjav1//5QPwLNNybf7q2Jxb2kU9uHeNxOaxdEV5
TD8hLrogVexovU8At9EKKywEHXfBk86QNz0JntNllDZujYJi3SY8vcYHyuOU8dVfhsjYiIPqByDM
NgNn/qmNIt8OTmxJ7VNCbE7PJnK2JYk8Gk3Qd25ZXwA3Z3z+MysZQ0vO/7Gt4ABpdATueXfDDYA7
ozqh7klwar6ASuSl7hflSGdaCh4LqM7bfHWzn93uh7SyPHhmyVcUcpmdi6rTI1Xoc7HNK9iKilWD
1aXNVU9OIbNkjLQtU8RNtDjb8nUcJwcUSJ6MxhZGW2sNGxKasgSGdg5eyJ+FO3xvLVgGLbOWG+Uu
7PcIXpfCg9BNebGz2HIN6A24R8/Kx3Iygrvuwy6HCv3w57bjcXIQD25sAHVd3XOr239BanzjtChu
RpSgmM0RZ5EzEQyjHjNrWj7kthJmwUVZkgQIPPpEnLAO5ZkNoLYIAgBJCYRiEOrMymWIGkEI94Bg
R345sH9BpGCqwtBegXHspidt+eIPVdW7cJU14FTGtz2cacFZoI8pzS010R0JGBg83tOn/avkm5lZ
Vv1eGjf5Hjdt3rSH3y6Hluji3LVYkYNxTeBrxascVZPjWdp6KMFFAlgg7qGu/RqS6V0KJ96xcz1k
ix/sKgkIIKUEWvNEiJkcJhG1pfVBY69uFr7/qr0zRfAbY0pXMtEzIlX8uU0IpTKmETynlgtCq6FD
H4vb+Fv7kiqrz33BJ+hU/hNJA251j6cgsF/z3iDxtsZ3AIfdmzm4jxA1OMlROeogcK1G9If8QKqV
/YceW0n3LDE59gBpLD5MSXStOswQJl5iTZOPe4kcKRWntHj3JFBSmMhG1zMEVHstm9WCB3iSuTvU
1LPg6uBPNfMmNEftNCUzWjtnb9KNqb7hPPMTnzydwOxmEL/iVfgTxYLbh1L+QW0qEmh1GA1QD4zD
649dswlKExlgNToZmdhgOgxRjd8517ZDqsb1YR7WY9rJHdCL0WP8vlR1+D9a5xV8ONzCVsCLO1ht
QBrGBvnmF3Flt5jylsfZ3wW32SEQPc+pz00vCvgycG9F/k8JMRrxkWGqReEx//fo6/qajMqpbt4w
JZd1W7x4r1vi7sqnZtXzdGKED0RNFZFhNMHge7Mo+QkWjK2JvPlEjlOmIyekqD1e6WwQkrFMx5yI
UM/9ytTJdovASEn8jZK30OmoqCVZl51mDOSrofRRiw5SqoX9qQM/UIMC8McHDS1s5qsAt7TBMw5m
JpKVizpM2hwXL0UameoBfs0xQsxj+MhNt/eUKX1Be4q1AqVZJDBS1JH1UmnzxS1X8di32o23AtxD
NOfaQSFUJ56+vjpYmoWq/k+ZB27EZaf+w2+GTULoEgAlnYil1WdD7vxiCA8u/ArSLdTGaXpIbX5U
jBqWcMMkNwEgGyFMsTgLJaFZh4oIqv80Ui6Uub1tdyhu1+0CYeBR1sfsflnGxjUGeuJPH5kmNlVk
NC8RDtbfTtMmwJ/CzkTD6fQnwOkFiIL9ZnS1n5H1hihUPY/xubmYJ0onpKo1+ztg0/e32XiOlNH0
MJA6diPic4Ea5HUFB647a3c1K4DNthqpIR7EsfUsXsVPOw88ymi6ITxRLOlCpBLy0oC3lEoXDi9Q
6ULF54RWfBK6ZB4DiSnVqbiMoKs+aedWjXO1ei3vt6wccGLMaU3t8I6nQxw8kYqTGzu1iE61CRY6
4+b1EUM9vezmyE8QGY//FjZFWIQaSg4v7+mc4i6DcnsY2BPXg/JjR/rHK1mIhy9JZCBPTAlBiOcj
n1cARUIda4flb8MtMqfytRXfEz3FV3WD5X5KltIrptlKlBUlmKv0gEOqNn2B0F2mk3CkKHJUpMgj
jNysYYI2CorIqvv/WeFrwYTmmeveQmZEVie8gun9ysvj92yTcQGe5Wxs2jJr58OROoatWFw4A8Ig
g3CDTz9M1zFCGvMWMOS1lSVwSv2nkRbW1JqGl44rDUpMYLdCXvF0VSaHJ3qDVYB7dlXxDCpK7slr
6MDzTu22fKNMtiv1C1p9p2dnhP4R7TXEToGslSC5PY9OOCEuGXjpWJziGw2IUIw98iEHghwMIEoK
P5SsvYmQzjxEZo7l4JL1TCXvAxcL4Q9yGXUbFlTOw4VKB3ZqwL+AvGdsUn1NMUMsLPC4mimHmWOb
pNjq6+pvRGAffvtAoXT9mSLLeWXeyVOplGTjbj6LUstqLVF1qSNXbwhElTDwrEF4ymCNODxNGSoW
DeauHDUQmXBmQFO5yL87tlMJkfXd4INSTkRbG3Et6uh5iFH5emjWQ6maB+hyctgkxCmobCRoEVut
KJP2oca3LkDNJb8t1JQgXdCHywML99v49iUy30Lpm8Wc47j4NeR6X4BpbhHJ13o9ddJBpO6fXrvR
lbK5jArmdjAZg4l1EzSnfn1HBwxqL2ATLcwLoj5t8XSf2c/euPY5N05PH7PATaoqiiFAS0rb/dRe
6MSVBNGZWWEWXtIg0tCmohQ8WH1Joijh9c0w5mFbNrZj+qostawGO/1P43sGiB9XhBwfC1iJZmQG
bQo1KyPOmgWUVRkIjyOu3Vfi1RrL3INVgHYwrl64HfJCZTJ8pOVn2aytcwv3AMgLmA3hpxYWvItB
Nntk2VFYSUPkhHAtW9ZL57EoeS7ulumNJ2Db+y+Fv3vmiSWNusnD52Auu7WLqJ0cAhrKWONDVXVm
v2JOkPl5avlttMrUGbWL/oPjRgGYqMmoKIPWE6eFTVLbI1ouwuEVqpENnaOloox1sdJdzXuHXC9M
CfmfHqeowYq3kHVFkOWwwdxpjMspxreCzv+v+vC62giotBD7WhwA+rAZtKvvfBZmHycXzpWOMRLN
R4W6SBquJOPEpy7wBX4WPg/ZqXU+zRQlHvYCegNxMjXR80oyAnhJ2kQs8A1qCvxUNzupUajYbVUD
mvMJl4A6EV9QeOHV/89umApPx9R7ZxdX6dIhsC8CSx0Y/SFh4qzgGLxjnN0EuTcBXBovosuZgnRe
yyG/HDWTZKAM4+iSac0sWAPGaKDhZEgd/bOl1Lcq+FC1S4bC9S4vN+6M+8wehTMhuj/lSxdDduhE
pKo+akdICGvmTIepGiww1pXQc9zMoz7oR38aF0WCUKEsm1jT/2goia4OecbgdGXJ78YttmYF8q/E
KOYC1AjrhM9VJbjboNEOFjBZ+XQE+walRlsIQf1n+IyWZlwDFQ5aCnkBi2UeEpkOP7kpZMDIYka3
bZQNcpwQO7+qs306DQVi6civ+OzYcnmoBbNUGF7AQD4ENvuyFgjmS/MOMSqO3YEt20xjLr+xQB4d
1L6WChZUpv+FFvqqzly5FVkiP+I/tKPgJGtPV4hDC7Z3X/7gfejNGKMTaQAe4F4XuxlCmWd4+1Gj
iuVK6FEaxnpurnxwGExbbA5uxJO8oG4mP3ZeWn/1c8nByCxSRITli1/EZQHzOH211q7kaRTF+fQG
vU0gjEtk5eaO3bDDO1UaScweznGJeW5Y9cXPl8jcNY67F1SVlt/Oxi4lwdXwq0xmQ//XUp8Lb0BZ
17lc6VU2v7iVkRe2dkZWHRApBUkDJ0e88x1ak8S1embBryhL1CpmNo3qHrEBQJ8l0SS1b+NeiCGO
dd7pUDSN959skiU/t1AKjq4shHnr+KYVR24YHomKajZ36O+Aog01Ry1FHDd0aFMWkpP0gyJj3k5t
H7Z13GbvjIP5Uj1GZFpjTfXWcPIGMUFOjL1wZJNJG2JoJb2NUhhGM6uRBgrMFkBlot6WxpXQOL/K
oBwUrlJmFhjywBFnO74rBGk5xX4/eIg30DWzqcOl/inI+6RV6TDQeZE8TL2XHx3ZRY7x5A1YWkwg
NuNVfNMS+WJkWWVQVgRZioqwGbvuuyruD78SAg10Fsl0mH5SxgitOnRpNIHs23jMKwMQpRKBUeOQ
ZDU3KQxJrJQZrVgvkWdsKc8cf6wiPZXLLaqu0f6spb4R/sYxQApcVDrv8jWqgXZt77PVH7C5ET9k
lpKyKR4fsBpJBQAPiPBxO7Ysi5NPcPbfqiiY8iA7s8YthcPEgPRqI2YQNBVO8gkb8taHaANFon+l
bzd1zqzuWNwnf0S5YEI7J9mLGvr45QNwuIakBI75N2EJvtzl9pHRvObA6+WZdYOVX+AXTCrinN2s
NfKTl79yuxaGHMf7/xsUJpBiZFt8Pb8JrZK3rpaHeAWMGPRSJs4+V7EDO+gguyhw57YQ31WFPCYC
UtSjfWF8B5NFJ+79cyDS+zGBcxro/81NV+A+/X/OrvaIoEFwgB45SFh+Rsydg62O0IXaJQoSwtri
fsOcljNfQa448IU7PH2P7Xk3TwYkaMF5BLWZgZpxPvTqYWC0sqzsiH0RWhClMnPpKfEE3iuqKsPe
9lAkai7eAg6VfW3xWxVK8ldMmdqA7a8DuG1N+SvgU4S1BTNOJafc3cVOuJkrD3YOCG5LKOq1MAfZ
GuXTJZ5s1mV7XhDT2BATXjFwflIDTQq5PPV1+rwLobK1Ab7Z4561pONh76DR5DFpIvpjNnvPTl4R
4BXzQedJ16g5GoUlVv3ePfa2TSKTYLwXYBJU5LCTL2462sAI3o2Nj3ZB6ME3LoWeEy9Wy1iVHo5a
KyiILGbmCFjxe5tgvfRHLZs2ACYjI3RWZ08AGFG+AKVyjTGTq8/8yFV3CQXQcwPLcj6jnpAM+z6A
0QvaNAZYApHdxTqkSTmB6m/w2gparObAkJoBxm9Y6zX17bY00VgayGv3engTTJ9kErMv3YTwupqi
F4I2LyGpGFF8JK5sY+pOA1dRxWxEvMOaEhWWvrtyAVpuQCEDTPUmbH8XdT68t1u/wrqKFGaBssRy
c8r4Yoq6dX/t+DuJpKFjGPpQCJGF3Ri3R9FLyCNoBfqiIf7R/BG40Oo33fwf0uyWy2DM7zgfJ2Zb
ceS1L+xYraEhN7GMekVz+lEc4Tdq3fnmnmKuRn8=
`protect end_protected
