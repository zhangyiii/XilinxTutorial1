`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 213680)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMKSJF4ybxqqynmhS2QDZyMorBy
54EkT7C24tIue/c06suXs3UM44KaSZwanj6Ds7qCzstLD8HfTAIM8cmwiPzApSi5Wn8H50goG918
3o5HesA/3EKIZt0Ei3zAf6iRvyu192tmxWUgV97Bd86EpEigRmUBpBIh0CznwGdeWOyqgw5z3BdQ
kVzRagOiuzT/nTpbnrNrg/TKDVss0Tyy8xLvxB+T5STWtljqGHI1NmMCaj865VkcK4XLqvJVZmx9
kPM9fE/db5Y8ZnDeGLCE38UTsroU5wrBMlaInUUXeC3wPlgRza7UQJdCbOzQK/c22ZojBw65JA4Y
hjtW7Z1UILp+qO6d3JjJx7qlCrkBWW4tIqhaAHp4hGDUQO6beI5WGMCjMFhwbjY6tAU62Is5jZO3
lysTuuqjWTACglLWZGGi9TPECKsfH/ybT31TSxV4xpVvzmt5UQetkBAcW/5Uab8cL19qWRJtFLjX
hiQLssqhKJgEabRPhsqStJPtttfw6HLZa36BXlH8urVMUa3iUWovsBEdCdwGfL++rtIRI3Rt4DwI
uUKhOWWWHlG8LTL+e9awR4rW3sm885oPgVG9wIr2g680oVr4gZtGIEGF28DG2gNbp0x1bkY94+mb
PYd08ndqeWGeM2JwZyQsYkJ9avvLRy2Ot3LStMCpWZ8ub9E0X7UfESlJbk2MRGWBAHS/cG4VwYnk
wg8/CdqEI5Iq/2T0J36/TilrAZ6APIoZvWLUaEHt6P2OXR/HZGxuW9Gw8zf2uoOHM2cldf50zBL1
NNvjUpIa3ZeK7p1hyWtLaoBdNNT3H03Igy7LdRtAtb6tnPEm5Zk/uurzlQaM8jXIRmeURxMo5PML
cQm+IrlQkrlVtLA0KQCjxcf6JtyqFJsi1cKBbtRMILUkejj8i04ZqxOqht8AyY4JMycB49yMc6GA
ku9ZRkVTH9LhOwYe8Wg7UEwxJCAEyB1s8gV0EKSTqX8PHHoBlHFQEAJHdbhoQQP6SMkVdW8ycmzK
0qNE3I3dp7ZzCEEDF1Ajjdk1/ljWt3fXMBOsCa9QJfYdbZFtrQdpUYKBwTlE3hrriwVmVuBKy9/Z
EZTe3eq6k6Wmxyff9Ot2El+wvg6e6tWX2dszRQqswZ1kIBDlRY4B0YtrQLbEUI+xkjvu5Zh8HRg0
bWHGEgPW6McYisSxBxyEJWVBz3pAoZiDxnldVctIvZ3psGeyY3LA2ANjMKJYM6DnVBRVqynjUSTX
FA0O5txVtZDeJLKlTazKH/l7YnPcmZJCux+zhdkL43/1E68x8eT6OM2NFG1hxVco4WU8MIyrJxip
GQz1oWdNSlmnw3bw/TNIvGu43yoxMPjxJZsH5kX3Y25Pt0vn6T82Mtz4UCYaoYsazAiwLPUY/1vm
fQ+Iltt7LK+wDPvfCOL4WLlgPnyJiOkWNKtZHnroa517Y8nsSe9FoBneWJSPq9ZTjcuM6OTE5oV0
8MDg+gp9piI4mA8KuWSiIpqWx9sls0zX/rFoOaMBAu7o06IsRzaC/k9B68fLXTvN3NtJjR8tMC4n
L+irNt9D479+C4Dj4yNAjWOSB5McbVYAFZ8yv4hIn4Ilf7eNrzEPnktCwLIsqSTfK+AdNud9tdG8
aqK0cMDeFiTMKbAB1H5UBmXSaGznhoZ8hLMf9Y+nUJHDMUHcDf+7qOcxlF5JpJDvDnCx5h2LkrH8
kPruwiB04VhyP/nQgJ/SeVDapnKAEWA3plPeKQgF/HCDPWN0Lc5V73BY7XKQOF52iU4ZV1Jr8RMt
NlCYuzFVFdo4Vk55Q/oxhtit3RU49GLicKPsMNGYUxXWagqI5gfhFVONu6LahhH1ZNFoD/ghKFRg
EDo3gqI+M6h/8NTsmcASekQKovIlwiIuCdzalWH6hPnH8U4ayBAlH80ykmcG7MMWzmLuHPXFuFi4
yTwuPJmk1ArpzSX/zCSAGP/fl3nnrNVy5QXzva4stZzQNnzRVTIAvZCzquvrb2AO4LY+/Q0lvWFJ
31cE8IEN9sFaeKfhC1T9SFDM9fjM8i9S39lydH/KD8ai/CUkg6qWGKOcX1F4Tq3XSYEcQVSPvgfd
+OlmBzTqBHghpgw1UwXXZy3QO8o1i49l/C5yeOwHPoA9buL4bipOnrNpQctM6cCIMTCOgdWLc+Kx
xFhOUbNsp+UTLoZT6cDso4admu/5tiQSsu0oe1RHWbgbuXangu7nb9p4t9/pR1NtAjpBXu5T86tT
flohZfiIf7cHsuQiR04bQlQdcZWHu03vK5Gi+KZVWGDaBTTPLwQcjzn3v4l+RKwuSGon28O9zuOX
Eq1Y3HuWIOIz7nE8gnu+AAp5K/h1vDMWGFcgJI0WyRL7Cu2kc2xcHq79ninow4eQN3bXwAR2Cjra
LrO0RptaEHUQNPvXEf9DxQiZlL+mVU275+niv+C8zNxfwog8OwQuKs+UjAIXoCdV1gg8p1r1w0Og
2tgKo1wURiNGKt7lwx0Sezpj8L363qzxkX7RcHkl75fnUiDRCjLzVOzn64yIsd3qrHKsgchoTXTg
iB7bRBPPZRpH52ZpsTPGcU4J0GvNeBx44L4F7eHS29M4vKYP2jwCh+IdyW3r9Ygbgcu1kaAwvCOT
Xiv7Li3AVb1N3Sp/L7/DY7aJPv87bfhuZlmQ4h6nci/IkuL2ARi06lriDUR8mUUzXqZgI7Jsp+r3
8EhAIyX2LXKeTAlzi9RtHK/MHqWvSMYZj6kEwfTCb0QrfIpJWSiB/0Jo68P97187MCs4vwFZY/Kp
mzNhwNZ/CPJqD9mUkvF/htmQ5kYL3VSE7chZQRynVo+EU51iEs7nxNi6pPM4Wm3L5D6TUXHNmjeo
8Fzf86UfOZglhPGooYBbuhzOY5NYrx67XOgcaebxSaqYqh9GZGUkzGq9ZjNAPyYWMftVhzy5wQ/X
dw68PkuRpNccy/2zHb6y8b75YvZeZv0GBevgdBK2cFWx25uuqEA7KOZ3VvS2klQYfLDKy4aQqNU3
6q/aUMtRDxdApC/7AEGGGWbZ9UQdw+N1ysjiWSBXr+7S1iVLxzV8Y64W/IPa6irq2hzLaEA8tdQy
l9HlpnMf9Bw51k5neBZFwR/y9QV0qpvQAqzuQ2Szu4qJBYn9ActRTr/2h6Ya+tbKliZwBierrO5L
x8wjPIpP/3i2chwHmSYv8vQgqHmLQx1pcHKmlHcNFJDxkgjEtjCTSKUfA8rGc4Rts9JlatYPPon1
skgUDt0mgyppqka4SynjvlokwV2F/mbb5jMMWAuh9IjFOXePA8UlXEUDBiNEAhPIWeYR3BeINt7f
VnR4L66Eg5/FwUlxu0zFON5z4iwEC4WY7XQF2PjBhKvn82wFurzViXcXGxNBhokFiOH00RcKTa6E
mQXWNs/RK3IKRqYMo9ghIUDXg7kpSwbeecUxgq8Y/igTmMIXcnmtGhHSPKiPNPmciiPuIqDTS9hN
GgbMicsO0dHSJf7ZqcEsfQyO3rzDltcd7oY2wKc25FOsr4qTMzMwGAWCKhjtantmQzMdZpUayNvf
x+WypHYZzckc7r+9R4tf7lEGeUTHFiGbi1Uy1kDVm5fQOGw/pIvdF75g50qH46Y/wjfzuAWhHhy2
tVi8kDHlgf9k78zVQaN7T3EyW6teOnf93qb67WBZSFnkb2SBd7qV6lZ+E2frhVSz2FKbi0aazU0m
N1+UP0OBg2dZIJl4M/GbUvoYWgt70e0XuYB/RUzMJdLX7lHTex6L6CHsiy7pHmZg2IElGKM+Wtsv
wygrilZ2SZrZarced9+52yHkIQ2jFb/8sudNCWOIu94667xIkiQLEelg/LyhW8a9d7xFSwY/roi1
+cdX12kM+ugUfrph65bSL3YG1usFza1TNV5JiqC9PzvojD6LK+6PSXD7tH6f57CpsDOfjhh59Alc
hCuV2PP7csKyaHxRX7di7op20YXvUZErZcQ5s63jsMB9NjIzlzlyhaG66GVlnGsHeZfFTheWuQdI
UPy7HiKu0H+0mHOaV9gFeNMO4fVYnzazA4Echsx8f0JFK3ssuCMhohxDmTFxanGAJNBPwHHeXD7B
Kr5NJxZ2WmCeHxg2n9lpmRZB1xdKW/VmS4BC9cOPQUfNZp9Xwg5ru25Bi7Yu0mPpfu1oR/9bDNhW
BNQPrSBpSXdz5uH2aikkUJ6eZEf976iB4MXVzh/qnAzucmVwRFJi812lgYKHh8vAbE+PfnAnvF5h
47zxJiiXW+euQ3ZOY0ookmNH+z711jeMbpLnKnfQbWSRoQYhLkSpU41IRBaE5HFQHalB8KaJGcoI
Jdln/4A1TIg1o60+WhG/ZgM70I8M8lrp6QsEzY7Ol7A9Sy/Xk+XKGyllVouNbupEcP9KXrRiZ4yU
mtQprUzaIlQNYu8lv1wU2e1YvCF6LZlrAPP1iF+qLUSmLdVW5FRrKBiRwvMwDNQ0ndfD80MoKu39
9j7e7C6MFYB8JmqZpdrkTcu6FoTWzHEmqCbND+jv7BPyptu6gKdeuFd2lILx41FzZ+uMPt8mELcL
Rl6RUX62NXpjbfrWFv2FZHKFZMorwX44/Td1X6dtuIBu/7zZFeZHnkBvnGLHlYdQiIz132uFWZtb
M+0Ch72NJU4Rb56amPVPxb/FXfYLEBgTxDOe5ll5VIZrM/EtMqX92n4JFoPWVOdXwz/DuwmM8jCN
yvhwKWlJBOaY3OLZDeypq208SO+7oOruyKEP4HRjt/x0mvEpYrk0FdrO1Vnj370EA6M6nti4HVj3
/t8oMecC+Yqc6ULHmRRa89DnAqtAhJujBS1JftP+faoU/n+NRex3zoG1lHwJigat5+l8yA3GlTy8
YENfZIPOPAj+TNO4nfDF15Mi1AVHYY5oVnefNmYrAnxIq7xVa9ZIH4b/IbxdDNgK8DvM0wV8B2PP
OD80W67PVOIbcDTC0XUpiVFL2JvAhvU/SULCxoQWovk9NTNTbQ35VCWsXHepef5Y9BFdAx4S1ONr
RsGvqLT2b+XSxSdBsCGV3MEErkA/4bDg/esgffGztkGNeVaeUPMYemSABkPSRP/BRFMSZvMCPhLU
SF48ZLlLgUX5JW092599HzNV+QHtOvYDJpcPhTaK5BspcBL7gFlasl0/PFacpZTfj9EoJsKuePBM
OB0SQMZcaNpdS2aTLeg4ULyKjoA5eZxZHALlWCUI2TbjNVTe+GdEqsqujW7LoUSLBa9VdhZXI1Pl
bhgapq7F2onHy6y2OG/c0zCR248pfeHOrJlPkSaukytNBahVUZy8GJmvzje2/GpSr5YGhWoaIFT0
FqpQts1wnA6NP4RXX74hLzUoGJYjCcD7PnoMbF2Gu6ObLRY1t6lGqlft+vqbpjZp9DoLtp3PLoUm
mjE2aQ5nTegPFZMVgBz25hOIKQmwehL8zYtnjzSB9ETAOE1NeKLikot4V2dTNjdSGZcZ0HymOobJ
v9F+K0Eg6m3C5J5IW8qE8IwmXQp+aoy2gXY1y2Cno/mdADkxJey31/mNCMB1WfBQv+9qvG4WXTSS
9BEzg7/sP6/V8wg1o+K7CbB5tADRt+iDso72gmvBRXQcOYVyl096ofVEoXQK7Po2fWfJtHeR5VUW
MPemSLKpPJIr727QfVqLqkCyB0rWL++Z+WB3L8NF+SVIkw2LKAWVNKdgL68EDSClvlpKXu2ABgiQ
qeLr9aTXOo2EjudnM4EHP/2Q+HBOOe6ZBcAMrgsc6c4jyJqCazbSjJwnlPS/Fwcm1C2c+UTWGZ3F
sMrKVrC4WlMy+PxzQQX/vG6C63VlFUElQD1pxrUR7BiPXA7AwZq6NxD/7z3oSWIfYOfgyQJ0Yehz
q55eVpSLgDVeE/WKXwNXGAwbh/PwM3IdZk1a24LZEkMauF8HymReu6neLSOON+fnqDUoeYUNVVF7
039AMh7BF7vWVm9pjGbiAq+mFjn2t0ofNSRY7E+olh4Xor8TsluzGAqwLujz6qCcJtgfqwxG95QL
8G0KBpYnV4LZR/bi69eUu3/H1Y8rN319VBbT3qMxYATNd1kP2ZfOh+G5sQ1eEUgg+N0MyfyYcdlh
GsQHvbyzxmfivZSBHJ5Dk9JAhfENPrXr2Ca7StZIbIIpWIz5xky49PYpNUHacwfpJ1QfAb5t0rm9
VT4bPXzzU1Zigu+K3ETcuzhJHFHkCXr2FrlTh8JzKl2vuTXkQ51fptkSEbqj7FddeWlkfAV4KTaZ
iM9j/Eg9AvJBXUePkx99GFoJhhlZchaitAeSthPPIOjUDbGzw2MZ+6KKdF5GVIrZP+942OGRem77
z/ArAuJz8V3bXEMX75xwIZQQAYIEOgjuxoQYUfaq6fvdQmF7SMZ0cDpOdQfjKFFBRfE/lJR/Mkzb
UAX2CXp7XIf37Bf4Ne6IIm3RtcJzuFAvgjCmKJQga/jIeqB52Ir0XBuGe3kSPkekmfTAvVgDBsan
DhiazhqURt96GDbcLrYZzn8pMFcs9NJMjjPibHgIe6MkeBVvjLpm8rixbKbkqXsohMyVFSSrfjzj
+DggiJP9Kld9MpcacR0UtsFh3HLl+6WUaL8DS67/0wN2JVVbP4tNIuM8ZcSRwRXef2lI/Zjy3SRF
nZeoGJAl0Y50cVlhqqTsVZ5dmJZKM8GSHAosZ4sBgxhQ4ouj9Z90O7FK+7C5qf99crsFhA4tQ/Oq
8TVG1RO74pyyKtYZyBhJYYmJPT16Qch7FgAK1/dYP8+9l1gFzZ+fP6+OPOwSXRc85mVJEwCgIiIu
vrtlL2CY7XZydCx+qg2gUeDjj54s6G9+YTK66H7xk9SHHY7EzihxcDX+IwkG7NGbW3EAprc3ebgo
SDMqT5bC8V0dTyFdjJRmr8XivABEL9B9cW1lGdDE+Y7w+hkJanlCAAOSVD0KAWfvOdaASXnlj5Jy
d1BKOebBDrg/g5JPc5oaAENWp5/36EUjxecG9fIZxTUlFQlXzGb/okNK6ilN2i89IcnkJfhNxT7o
6sn+rTR3p1DHEDV6cPik3SfEXzQcX5/1IyypLMMLNcuiA9ZaC9j7F8pLoIg5iUIfJ5w4gLnlMFbL
iejUmRLbWiAAeVyTVQpCW4Nq3GZysJfbR8eb9jnmWRjyvu9wPgFavTPiA0cAGf1Af9p0kVTh/xYR
gNkQNuFxseR8IyB7sOeTjDLaQjpm+1Ry+GfPsDPDWVChGllJnmBja3gsa14Yl+6D8zLdn1w/Qa4G
CJ9CpVyvINEksXXBUbcUTvy/4eUbaVV4CEKDllFyxJXE6WDl/x9O9i9yQIoQ435XA2GhxtqlawVQ
F+qdmvjeQJojKeSKL24PSw2T3OxTlYpgPutjmRMx9fGE/0pqi9yi2trmMK4AmJIJwJEATLf2H04X
s6MFNOXzmmDAIH+kTf+6GIs0wa39Y6iy890pBqNCExFPiGrqorphsyuHLzN5YVYVOIijlKII9ORB
jZ3SYJyByvWzdhXJSh90wTOJjZy8mTi94J2+ZuL++QsIgWnYrEzoZuSwBmRXo2Pr+EiiqYceA340
YMITPVjbProlqfDIMNzFgQH3XmPUm6/htXWPeNT+Nwb3CpxQd7cnY4jqYYaZ1A4DMJK1gzTzyMs1
CvWubQGqvTSDstcxZl8aK60tIHUB9HqkuRqxmFXiMT7A4yfNizWkwh0vNAa6kiZoZvJnMvdrsTi+
AJPi8ZsTyOu1ihJGh7OV/Sa8B9PGTTYSIz1/xSGz8vRly6V12oRYdW3j5xwatIi79k7+XaqbedXZ
D6Mt1Z2X6vt85RGV+smne3yZtitNNG0ZGXGqwDOF5xKXB2YkjQISkvXkaRkVA74gitLwiz/FR3rG
G0E36jIuPpKPP6sf+PhwUg9kGlmTQ+4wtabqfrQiStqHMUx5Z9t4Txbn+rtjWRIrhcnGAatuVK1F
UUIvnu3W/5tIwPKFfT5VAGpD3tZvrl+3nQlsveBIPZDv25z3/rNS/9KTKQnZHVsQc7nARelYd9zn
i88nGzvx3bL2eJlWxOgcs/bS/rH9UYmratju/UzOL3ZllXmzGeakTLkzlmeUCa6NCdtgJKyes+3O
gYCr8OZjW65tys7VflJn7bA4Le7aI48pyf3dJheo69A1vXqyD+vfku0Zte/0ZJ8vP7CSm3hR6vbv
anJTwQscdH0JDhr5H+joE4K1VXcsQ/0DznoUU18oM5hlYv8vwVsDlGmWsaUXLYIdPwRjG6OynaHV
dwsBDHuQIWSlPVpsdk/PCmvQCu5yfisV04iHZsBMtHCXJKUkfvSTsScTNL9eCm8LGHfDU3YgmX1D
r4ZDZLh9VJ8DakW77eRxu216iVR+/9xBiB+HFk8OMP7d/dPkCdPgXouuNOtL9+j1wmaq/DiS+94l
6aJsz8CJV8kJRS0zqOB1iR3G2wcK427wzi2rz2IAJPXeYS4MXQNYUlLlpWqzw3/kjdWEPmBOsWHA
7IY3T9KjNr30K5jDsV82T34gE2bUf2553q1FPzBCfDPryzGQWVXBkXKtJsRxv0awXL65lsoQ1snD
9Aa/WaOq46zv0bTRBmgxVpJwF35T5QCyL/iz3V5RVlI/b8RVUzUgvJbEFgjM/lHLPFDpXizHhhJI
cveGy+JZSaXxOVsJ41EzjyLpyIyXJiLunDG6DnwLFIzidEyboWqXDPWJ8su6UcvOI4hSgOMiII8e
h5iy4ExfcsjiF2sBD6whlGqGPyIoMHTPzW82WU6mi1w2i+73noooWCmJ1VlxEZt21BnOaTNbSOhK
CW/GfS1LuT9rC9ibuL6ClaH7sEH7mR3LUWz0grwPFv9uCLWeQo9wdrGyTZZGT7bKxkzKIHTImp3c
1JEAaOcqZqFBVRvgGUKdmh2Ss6R0CO72RyLbMRIRdMXHOb/rBqYmCAJ6FXIvJgRRQohuZyxTtv0Z
9aUz70zl6W/ZmBNwvLUIVyec3yI2WY1Y6rv3mbuIaP3pk7cPcrTctgsboJJNe8F+ALiO/+c0MnqK
6+s/mi1Lgcbryr7+eVnGLbBPqSkb/QUdPTZv04mSa3U8g30EqfaCuUdnsEG6BXL3qSS5wuiedjtF
qFsa4Xkn9Xh1AeB4Xa5oee4T6tmEwjMofTjNx4H8iKakFkHMSCQGJeNeaj7zlrSGux0yB8cuhAsA
GXlomF0OpxryOIekZ8mqLzNKn6JtpQWgo3aZglGjR2EXx7wrtmfUn43Vsw/DeAGFMljE8T2uZStb
D22a2rP/y+Go3Xe9N+HG4pZlzPxBCRJQXZofFnv9Co40B9Qt8EMdq0XWRD9Hz0gz4Y4In8svoyKR
j0/BnG7rJYrG8l9/8RkuHz+uePsHJ9CqrAMtHte9Vo2tJRYYTGGdVQrxOYRHsImWmo8DAw0Xzfyp
qeXJikIuS58AvUUNOprbjlOF73KLtQkFcCorUrpKhR8KEbmlZtIoMZOgUACtqRynJQXgSuAO8/Zz
2hYejHRMlyn5jQxg5W4danp3x1VeX3QcEx+OOCJ+xAnm1OBKr62Lp/DVH1OySZIFy4z9n/SAhcxE
8fqBSo7OIiRNtbmXWfP5Ilk+ESeR3jk1PHFJaOJtmp5y7d1cMGGuN9AYzAOzzYBadDx6T8Ab5MZ4
QGjahv3bibPqxz5Fi65pBbCbtv8K6/uhlgvLR8doYQues3EMZfBv0qBDRF9q2Z4y0oK+an6ShJYs
n2Y4sI+1ti5PUi9COWkUc2uscXRi54kVv5JI3xHgfqpOMIRnyKmtdlf5IKpQqmc2NSrjJWtmf8uk
3dIniHM4zfi5KoXClvb/AjktvXRoLH1/qbGr7HCqJl43XCst1qCP7LvKkq/lb5S8BRqlFS2aPJyi
B/J/z1Th7b266bJuafgcR+BtjH4VReLxJv87b3TRVOaAQylj55NmJ5OaiI7nizG3Wzh24drMjkGA
s+4tioA2epUyQMqJepqX0cSvjm6O7K4Ba2KvDi8d7jJoEiRTYHeblgSZ7CNplECZsrHYu7dN8o33
19q8M0RqVlKx0dy5hoa695taTxjVTmXEUB7ItOZKMsUF26+m12kAliHzZ7IuM/3WVntAkmn7IhVv
UK+edwdxqB5C3kZPTKOquoiKditzrrwAceXFBo5pdV6f/MWjVSfWHgysu82DaiPSZKmwWsMOVkWv
afhuxX7Ctkt9eHFPqoLBibL+FEm57SVNwTdIh81JPDhCL3YvUgGKurzgQu/dfDY5UINY++xq5ymP
8I8OM8gCjPQfdY1t2Q9GAuanSBs2h0E0kH+CTzWVEtXD6ADFeuqC8MBzrcW/le2I3dQKNSl6IbK0
UjvYwiqg5e1mfVcqsOsk0x8w+RafEmxef5U/5t5nA99zZNyFKTcKhtHuXylhUpUaXBb3Glo/TpuK
baOM+pVZ2XT+rANljjE5KTasyHShWQuqSr63KEA7Im9EdyLbH94YcKmuXIjH31ZqFO1s6c0Ikhn2
Rf4c4HHA75TkqsFtWdccBiWk2Xz6d4qgrEop4ky7ie2irUg5zMRr+HFzJAJibNXNbgv3YgpIYYNR
AMBQrQYQ1XezdsXGET1R1rLVFaLQs5pm/TTQv4WlvjorTZnZoAApf8FytIOXvQUGgGGB+LD8OfgL
hGbqbfH0p57W0hRxsGQDkpD14Mt0qTUqNjk5nkDLsG3B8smxLA8NiridnGskVLTZnxHZdgJWD9s3
65M4TgKQxPIxPoE8m47C+tjG5Ppz0ZBDPaSniapoa0l3jHDXelymBaZQx6j8MwIXUModc+x5M3og
Ze+pyQRVruml8vdagto7+kgIKk+J3PCxovbK20r3JO1M2C6zPdkeOy4LqpmmVuSwIpeQcpHLLt6Q
+k3DUb5+tm6RIb5T+HW7GEYIX+rEV+4V6hTI35n41NJC4Q2iX1A0VygKU2/0lJRUB6YvmEMlI+58
lB50cT6cOmegZ+P5ZPY5GylvtbVIavl7QqvWQgn7V792RphApFcf38uFkRC4phMY/6Pd7NRIWA+D
Ep8nLwwSgyM92yHOIEP+cINo8b3+jKDAleS/O4Q/UCaDAo5OhT4EVUcWTsAdgfTL0bIOLdXG/c7S
LII4qjmbgIR6Hxv3iEG5cyz/Nr8CQL/IVx5q/zbT4WLbgXf3SATKFj/E6ATdCwhTUgtmnfVmyXPJ
ifvha35bULganuJPL1ct/EJdfj+g1ly9y3+ly0HCxa6eDwHaYhVlZcdEKe253bqaeJMg8nczm75u
rIh/elTMQ431bsvGwTpE5otbjPxNekd9OGPy9cVeGT/0J102ZDV2vtUs755WSThuFNtc3DO4hh3j
nVcaP6To4cuc3FaicFUpMUwUCUkiLCLKu93cKovNwahEk0ErOHEt6riLrvTkiHAaXiZ5EExSZV+S
MWGU1AgVD7rQZ7P4IjWwpZpNRAbja9cVU4q3efz+y4NL2uFwnvPe2pxbOP5Nk+DE/OqlO0ZELHfF
XqEsGVmp9+xWF1W2DiaLTUUCULGw2ir1/ZAMOFu0X0L6otcghT879p75GXU7aYphlXMqtyOgNKzZ
JNdOxFqQr3uyqpxNa4bX/5l1BWzeiTnx6RaYmMZZeLQfrbi0h/v8ccv9AuVshG43mwepBH3gO6kZ
HR4yU+VELcd9O8yZMZ9VQjB100fIx4PICG8OmAYjRji3509Nd/fpfsLvpVKmqP3WwUUOxRhGBsBv
9oGxt8aNzArYCAmW90MT7Bu4zwehT7WTDwJM0cimrbq8r0/AXkjK3dBgOK3iqz7q0r/hfXKnhG9M
r7wrTNep1N3rPq2Tgaw2B3OyMMzYgfoOMtzHYqMBgKdvvndjsmvXksgObtAp7abvtORvdwK8W6Zh
wFOXeCA4B0hhKQ1uXpfYeSPe5N3d2FSbuXHMIy2EggP5gjVIZ9J50X3GoSQwnLXgHQgk0HkT96x2
SG5RUkpcbSRqWESj3X0dyzK270veQDLQ39n3IKKkeIAHnCuBGTa6AEzLRsvZRP9tQX117Xg+80Dr
ekv1X6SxF0M8vAZwlZqZifUkCMEIrOl2ebSGBuk3OGgWfnh8x0IJYHmcPwN05kzMZYGXFifLiPk7
/HE2l9ptAtvZvrLtd1onuXGHx+pLKAuXwoXRZRMy5Gdc8h59NCs8AegyAy4pWtfUpPt1xgse+W0V
r/msSQEkDZ0ewMAeybV1cu9WZVJBXc0nobNxYWTWHdNSVHrfDDraPn/Ew7a7hFsLbTFk8819Hnkf
nMNC8FR2BABuKXWb7+KeQfuqqwRZTQ12qPLhv5/7oXZk5+XMp8pyAVKeGLKwZJI3A/xY3ovXZ6/M
iU3bcmNsD6iyoofy2jQdWXp/R7o0MIYJrd/LI3Iik2dvosGzBh/b7VCXI0ZgZJeeiUbHCDRTMZwS
X6BrUMhSxa0pAINrScaZzYCNdhxaIjFLL58LZzq0AC5Uzg8Yu0CF+GyTUjGkD4Ibae95kUj6+B3r
u4xtSLNGwUDrzAq3BS9LMS/iyIVzf3SAnF9rGJehcLFNLv/Xm+ld73gYnLVRcLXBt/AtxiH4DERf
Rd7FV/sOvR8P9XASE7+8NaRnDwqLXtpvdODjuor2HaHmcmtCLvQulApyIpMZOO611+iK5zjUx7Lc
9a2GeyO6PnOMVdvO9WDeoZSeYRP8qWGtHa8L5QlOOpLxJJHLj1RT3v02UXEVr1+9XcAHZRzoMJa+
5Iel7FbyvewVoKULQ5Qm+e8TzgevIg8r1j3cTaSNg9aEdZLLwNR1Dh3407heNtIyQPNBZV73h9N2
oyQRG2VnS2inFK3kOvZzVKEInln6FcZYxQMo1fVTv7+diH5yHS4wFkJVaDJeZlHB6UE85V5pgU8z
5xQIOxA48qBqlVpcYMrbM/xDVT0W+gYyXCl/T0bMuV7C9F39CScPxkw6DXCTVDiiNIIgUNgSItpH
gOYDYF8S13QpH8TB+bEY4fic6YKPrCluU9ykbrqSvhMlxoGz9QAjFd8BpGTEsYFqs7y7JpJdLVMy
2bVBEq4VbawXMtw3LAkxEidErNNilIHdxFvmc0Os2pI4KGfcai+7GAhKPtE7f/u4a8xE/EdPXDJz
r3rRze5Vtr/g2CDXSp1Q38190GmJ+agDi3V6pEvSKCgctbhjTk5dRWRvF2Vz9MjCdXV2A+dw6tFD
aH1K7rF5AXXUye1hIEiWWrnjZJVN9HEdihoWOu3DvtzVD3Zhp8bWYNhIb44W3Y7dwvjNKtgNuKbM
Ep6OEd7Uqp9h46VJPgADiCD7N9KnCywd1wbebmegSVWtTjAP0qV55OtcHeM9yFgDwT5KuGOsq125
V+RU+4wLOn7HLhVQzhkcS3E51cdSQDF+kpZIMbzehs4q5yyyag0vAYtRjuxa02MLjRB+4v2mlVy7
KiVHp0CqMkIKm630jlumRrIRvvKZbEyXMfVVz6gMJUrAam/jiSQ3ePpEXBdY2g9J3tfK6hqUBG5X
0vbRacXE1P3XBQa6TufTKjPmlrJizETQHbMGW2uf0s4dUfa/nPTZkwwhocFekgdI3Q0IVN/FsSrf
os1LLsGao0ZQOou9BBJG7i2eswa32JVGby3/fte4oBHG/wGhYGXjK3KRiV318o8XxYArafcRkkO5
Fi4GYrdTaz5MPDxv3rxKxi/lgcasuhk4z3rxWrTsn9CjiC8wHt5+P5K0iaAJkz/b6bFXWer0xC0z
LIiyboHWZAst4VvZcCrXJn41olIAv8upXb/o4WSMO8rPkQSIEGScEZo8Wgx39OufnAHvpx5RzBTq
9fpXg4hboxgYhbfFj6CxaVaQPMg+W89jRnG4f5gYcxTiH/esG6thVyqZBC+y9Ei5WvZ6oSPQ+sRH
wVFZESLUcJoRf72NCARcaar1jByt5alqU/b/BBsz9ZMgehK4dszwySkNc8Uu6JkhDERozcjs6qg3
TUFsMNKc5v/hKyFgorL10NqPUTPv2wkaOxDRkKXPZXF7WKH+kRS8Dq9Tz/Y/OW8t5iV5caJ2dz/R
66KkH6TZcYdsie8mJ9sveEah5fLrwE//BK9O4DmPq0Z4dXVZCaNT6kWqYW3UcsBZciCEycKHE7pn
LwxgknAaJAHW/1M85BNXtBCmvwKQURF5+grZ6dtKfwd0M53b3+aDxJ6G5nddCLeNpGAOu5Zm/MVs
TRNIouJ7USLd9LodozodyO4ArYzWQ6M60FaIrx86Z6MC/hFUj/9b27gaPwvUHv687RDrh+ViYcoh
EFV1RxUTeeW9qZSIuq8U/4fOTjdJdztz+hSsN+t7oFBFPsd+q0iwqraeg+yDUJ+v1wF6PxckMV89
KCob2AxJtypsyP8e2+duJwG3LgsweYjfBSHTgEtQW2kQhmYVfzqfZ7JhpMB4DQny1cji5eu5pDnS
ty+oLRsm65KC7j/Bz7zTK9TgQ6GWsLWOcQBj+g9QQ2c0utqpWAaiFRMbzhx0xg3/Zo8xCGj8Em3T
JYP4XbE7nOwQRcVPGHi8c+0XYXL/AZsW5C6z2Jkh5WlTnSu9aVn0KwZx0jdFjoLteZJVp4RO3C5V
0us+8KGNwGFaupVnu7g5LEf1zEhjQkofrlgSV686hOG5ZzvHw+q15/quM1g/jITADGeZcrXWnZaz
umdySWy55l+bV3VDs2yhiQcT8xWtssCQoOsaKQd1QtrOjqKaa5Axp6T9NeZXDSvknzqBwByjI3Rm
sq2IeLJ59oKyCtBuGHEINClVoSS9/weBo/FSF0UmUucKGYGIPqLK0F2YQt+94A7iBARXg9TB0EMf
jobZ1NfnPxvPFOQsgAsIWisfQ0IAOa5J+LAUEZBRWLcl1mX44VcY8zqX/CulHFWKqJx/W3YVzIpa
kKBSR33J1A2gbFeHAV0Z5zsy5fpsmlL+Bs26gs7f84BtEbozwSOnPpGMuxyiGTNzuqhyyqBeCOXC
FyF9eH1vBAFUFRdSUBf3lpcpcSi52HhDpl9uqFsOY/GrOjkMOs0aTSnjh18pKolGdnP0MaDbgQwy
bGPseqEx/5vcQj6N6uq6Xw2ffNVmSrnwSGspGHmYk7v07wjqIzCf2wAojBfVzz2ozNLBmo1IbQbv
QsOlv5p2VGFoAy1w0yiIB7c0MvYCGAwuvOwqytr8a+56lUSF+y+cQSNR3KS9DiBsthBFjh1uJIgK
AkMfzTtZB7EBIEo7w0n2H3e7su5Sx5LTztUwHcf8CCHJBjAoT+sU+cTPSFo8Euru6ytCmKxBJ6wA
cVXWUM47lKgE4flBk9slWMWO5Utz3iBcn3wsH8lqDMzzotTPqLKnO0XpEVBD2Y1PnrxhpK6zScNp
yw6RpVMfTfPoT/FluxmxEAG7YsXshPXotwwoVTXsuOaT0HVVHno2Ukjz8/2PvkzKC+jAYy0HX91O
Y8DJhlu/R31aGLy0sUPLbeo4PYUtOXcqnb1qkXwIJmSmrKgPk16R8YnpQ+ADwkRaOkC5+0aqBRib
EDZQH4oR3Ch11GetwJIj4lxTbErFKhsmfSLvh3snPNKFN92GLKWoQ6AJuWjezR7jV5kH1CXGOxGs
CzkJVG2qRsluToLkLZ8pooBMtxGMbecoiEm9v2UrKPG8RT14sdgVU5yV8y7NYTdAXoaui9/MehxJ
yU9SVomjONl73W4hcc2I2o7AiXCn+i+wcbFzZbo0V3M3VYXMMxbuKA+dFL/8tmpK1ur7NFcw112z
dHJp2SPw5LFkEkotXYmrrEYDyZHKlh0h7MoIlDxb/aed8Z4oKHbISIXJu1DNM04bRWuv2+aRELRh
UE+mnGsxhd3ob488dIutq1IpOKllR/qW899QMZAo3JRZAd5CpRAL7tsiCIlKBDHraSu9HwS9ljJz
Zp5JiFqW159z00X6V9/57v+DmI3s/B8iPd0yYTJLYQdll+f9UNcpj3I6/meATsI+M8QmmYn82zd8
EDpvaWO+QaLUJZZOl/uznfHQO4J6cibyO7RX2yXK+ssGxeaXB04zaUv71IFI1ZVOz/OWlwYKClmA
PkFudbST3p/Ll1zjEQci00fRUN8VwQ7WII2+JWlgnlG6y6BW2A2fLfZNGLxD0tnRcaID120e/UJn
X7hT7flow/W3Y2m9Zb2PUDuv06ci0YMfOrb/RCfDgUbNlrcrNEd+ntpMViu3ZBGKNBJnkqkBT2Nv
WWE62wR1dtSt6wuVXR44tQgdHkJm1MhtOLLXN13R+/VR/NVuUWvkcp0gbOhqP4pf4wug1NJ+EvSx
RLJJRj70IOw1K/fVZizh/vS7XIpb4X+danNA+aRe7QqOh1VZhT+mrvHDdJxqsQ9JMaAjMV0iDCeW
VMrQBXBg16srvC8bDTx5zmAxzFU3EBXxtdqRTd3fLLQkTKJdmfvhZiRcb71q21o6vzGQUrS59GwQ
yk2KgdNRK0rPUpq/QqgADoN3Ngi5LJpNekfCgfNaOFMG4rpmR3pyUDrumeXXRUsoYxZAvl4E4qix
70/u3DTP5a4ZWcJTehhSeCQqwj/imwtUz7B60SgSnUm4uhlHn17IJA3ZEMQP2viiXX/ELbMb06LG
eOV+a7ssyqhTs71zYrWvCs10prRCaaYvCjXsYjUrgJMHnqUMrdkTTkEnvPEbhyS3g/A5Kh6Hs4N4
hD7iwUjnSaNLo2eXqve0YpErQURG2QgDs9WnZQIswmXGzqlQUXQLeqqoPYOtGoHvbevwQyTJv5X7
+CeNEF9lKP4UGj+PcNxcvo6j/2WdLpSHYTrASnqgrP/mLHZvP5sJ/yp5857H9fmtpSDWj/FIuH+K
FWx3iwDU08eiT2RckPcy4S9Fn8wMhjxF532XT+F5+XMw+jC+vBaz44HkyDfG1COvaUDGvde5DHZ0
YT7eSfQ7UtyiqI9Z/SGxEkeui61oWoNJCp7cvLhiO7zA0AhIIAuDdZOgX6CIfakqmm3eZsnjCpVG
Fe5t8J4hGNjM8vHeFegdtdjJDzzMxxeVmi3DZiqOrixmTTL4I9kXkvAP+0gW0Op8QNmHaAaoDaFL
G7L1RebE6tFF1qlnqHFcmv6RPbeMC66JY00di0SeSj865Rd16qjouHTwujrewroWLZws+vWB838G
VJN7/VoS6VR7BM1iroZB1DGM2ylxAJ8Um7SguIq7viRlRjDrxqhVxONYK6WaMja7k66uwmgc8/YN
NMiVAN5F375nYqTiEUsRUMdfpkL1TB5NFBcNDjOhvehTw8JJXius8Qgy3sdtW1GCzL4dsR/zgZug
7+ya49bmRG4OXWPk3fhzAJ48aJ9KTPoE1USSjfWVo6FVMsJhx2EkojlQuZpC4t1ti8KGoCzZK/uU
ACLfHgEYbLPkG5lOSYuWMpnauTq9SMQlC3LJfPnndH4fWezqlEvtGx+FHV3GQwbdReckNVpbwYx5
uqyChYi9GtL3bLT6IkowB9uFfYVkUNT4IQVik00afljRU/9bgsjUbREjOmLPqO+SGU23UCjOKiGw
c0M23IEB1cvxB/q/J6UkpZdiYgQryxRgst5tGAucKNU7pwDKv1sOSD4LprhUjuvEkNItc8ISjlEK
Ke2FXOgFtAb2nVVmAUQx7SktHRZ7Y2ZwGZIVkXSqeMlmMztRk684Gr+9pWAesz2Cl8Xo9Aqo6ZdZ
ZBHSfHlTbOks1NQalqyBAte+37IDC+sBCxsjOpeIny2r+BSegZ6QnzS5iCklTYGHvvkbbEDTPbGs
kE+z+MttvG0/fZq+n5MXReSNBH8vBj9/D5By2P0a86It5dw2m6BNN7Ik9althyE+bnqo9wJgyhu+
EDQMDkEeuQ0bn/wTox1ukp9bxb3OE7ibK7Wdba5/maptvmz0po/NUJpyO0autCbaX1GetJkHaNAW
M6qVriWoRgpRe43szJpPVLwSiPORz94MsohEqE2Nezyj6seODIdyId4uTt9ZLfSbR1boDmRFgsE0
Jcl+Gqc55GiA2tJ8FxNmPcBeu5UdHm/JxZhWUOmdU7fCmoKA3HGaC8yoynwpAeeQEYiaJGzEms5j
ABrZqY8FWYgy6RB/4zpDMbEfEcecODeAeFAdK94EgxzbwoqmUuICTrbSxLrsgnxs0GBD2zXCcZZ2
Pk9z9XFWq3msIUbzwocjLsc4ib9J4CdY8KM4UGioJYh9ONYveDEnZI/Tr0LtGgy2fOczeOhkSr/g
0LaX63Bg/ohlH+H1NdOdNZj6ubgj8Su8Sn8b6iTVb+waaIR8L2AJ5GlojvSOQ64Vyuo5L5kV11ko
YtzXciXovxINFW5+jJ7upLzpf5XTLfdbStZfQ6xhhxng+7K54fpUOAOiozmIZB1qoZ4ccoVye2+/
oxPEUHc8OASmoHGfGI0rIM+/HN01TI0kRKB1xDxyk2VwLj2bvV5vkxqTg0B1aQt/gF6hlrEjTAF9
XvtnUbWXAJDvrMaGdgDE/fjtKvvxJke6o+PG76oV31PmsyMMkyrOe+3MUDT4F6YyP4tZLTZEMxPn
O0dA+K/SGmPljs4crJ3Tvg5nV44w/WYDJDxridRefQrEeaL6natSslhytTyW6eefDg12WB/yVE8v
7Vdha5uaF94OesUWHHW4NHYOIBGLbyvYCe0G5i5numQMNwFDqINEMv1UwsGpggAe/ZdkfHTgtUcO
etIMUIX21PIx6tPtpU626l2BzCNMiSWC4zczSSwGrlgxO4i4d21crtQXuM/+i8spxT1x+dHj+s+A
r44rbSJlC4b8EOle0C5TIpaUUTlazolmoyMKZtl8Irm8MhQBirsME5qclwUvSEyYzZZc135RmLFb
1tFdCnwFMAgftQQJ9jmQ9OJaj9Ri0lS2olNnCnjjrlNCTJnc/3K9ikQ5XSYgsJ+9545pMCWbfMh9
wSKSl25W3/ew3E5VP+hn4YQDUvp9H2r8/36zwSCcjNJ+CBQVoNZziq8q708LUJfuqELxQTehjZRn
XZt18b0pQ27AzuKId16Sto9iKiU7ec9ZDiEI+Pt7crY3Y7kQE3ppAijuq/jiS6GBq3qeYroeKhgQ
Uhc8VRkA/wgeD0WSQn29QYKk/TNUcGytQbLcQJ1PqYHlgrf1F27/7xzOVN9dd6QZg5ULxlY1tqt2
SKu/QZZGKf7ktvqXhKJGNXWkZ5mYrPl0CDynJOd7s3S5L2ee4luNE8Gpo7ZZtEdapS3F+vhiRk/z
oCRtVrFMCR9vBausb8fHeYylm+wja7LgY7FWMEac6OhpKO4uqGwyDUcC+iCbeNZqXgdjG4SUzrdd
Ob2jPpXkolgzaLcu6U9UZPTqvGDo4PituHjE+q7+sEEd/dJl90+FBN3mmLP4u3kO/vwjj9LZiWPu
TejezFBbDoVbwdL6p0HcjplAmXt7sD6sO5UM8Twgv6vWDUzIeaEUNVDnBmBtQ2+63quMJJLMacns
MZgKIQCm8vE1v84fE08IUVsh1tUC9HgNzaPWev0lFrF/vMw1nJEZavQenGIYh7RL1THSxskGAdqD
VhW5E66qxtfwjg6+4LYpop59Qo5Dzvax0qtb0+KP2YS5UBDvmvSgsE0BqQ1kjALuWTHdyiqQhsvC
hTdyeAQ7lpgtQC07mUO2YgxUAJZnsPG0cXfexKCaXDgjK2rW/sa4EDYJFSGAwR8IvmaoOX30JrUv
3HvJuJT0gpGxChQZv7HTDnmgTEHIFWhdaFMdNKcVnObYxjW45PTFHDduGlq4IElLk/+GpKENPtHA
ZlHlxNO+8VDx4Zk9tKw9wk6EN0ipwexrdmAikk8X78q//4e/q+beQ5NGrdeObS9Sm9Pub8u2LdJz
PhjX+NitnFtoTjttTfp5glIpqkQn8OmGKyGBpT5/VT0errcDjta/AHJWTqxEXI2AtVYYJw4u7hmu
gVKI3UgOwltg68qbIY40YgrBS6y0jptrGKbJqpl5PxJEt0hwLRDuGLpuaeiEs/kLYsWYzI0ccLr0
TV1d0grVFMHmAzSnnHI1bzgUZAkbELtkrha65SUXjVvBwXWr8/RFIw2HFfBDgylWBoRWnxBxx+l5
XU73tJByQwJWUtsWlgTjBbKCAlZTrOQtDI2+mAg5KreYbheFtmJ/r9MictBRf4YNCT7IlqRmN9Na
2MFmPcBZDk7yEj2NVlZ4xjErXjsn4EfC/aL65I6dlVbouhqesBTY7uJZ9j/bpPjQCg1nEbAmMuHl
n93DrMiUEBMbRRU+nvpEjwVU7a00WiY7cPH2U0AYYpnyu8vP0kOBoeB7PAkeKK9jH8USArHGUL//
7Tv/EtHVOSqbIJWsmD7VWOTJsKzYJh9KZpM1w/RDVBLwHrmiNns8NWqv4aqnQUf5/9Mw2rzxWMyw
Xsc3pUKI/VixwcfI36YGjA2/mb7Lg71jzhWIH1A7LWOfhbjhYOBfzhd7ZerNFosuCrmkkUt+nG7T
0/rv3F572U/LHkZxEYk7QwRplIuzYvsoSrWPJxvTw1zgF80DhcvQ+fFvgN7jp9C+dGuw2PABmvZs
cFDPCoaOd2D+RewWBcs76noFllXmy07xgH8+ZRjU3PY1ryb/oW1E7Zr8MK7ueyxBAIDxH2FEOg+D
v54d5fifiktDbAfbW3o4BIkzmMiMYQEsMR3ZLGKG9m07cN9vm5xr6yWu0/HUUH/YP2p0Uu7xKay+
FZOWKLvkWHCLkbpx+QQ8Nmeux1/OvOrEl8aD99uYNGeFp14EbeMrwe4J8Od1W/4RilYSz5iYJ8lk
+Uz9e/OLLBQ4ma0v5wORYSbsVksP0ejJdUAn0VTUT73Re4Vhx2nu9STB081JXlSANU5/SW/d77q1
ZT+t0z4G8DB/Ex44rBQiivZOSqwl4JOIe+efr2OGbg2jaimnPtv8F5eAxZYbrEK98iQ5a91XiSLw
IJ5bgvbfbaGzlmbZCSIuggcPwZlLEJaYdJmYm4e+dEkbziLchfU+guENJYrS1f7Pa1Pk/PDCTSXB
eBevwYb1fOQEv9IkfkcTtZVoDWb/xwQzt0OgIHYkXJ3EW89ws/jz1i3Pxd7d5GolO+y574WCOP+f
DoifCMKEcL01+7Qd4qa/sRWsHjwlZUiI3xpexm3G2jQw02Xh9sbbGJuGgWLECL00W6j3oU6/MPnS
Mzu8JxtxIWVfpp1MNJicwqjzwSfHPvROqVwNN7EtPSE/ceA1kIVM/gsWLAzVWjY11regAUq/W0Lj
Wm5YihHXlNZk4VgcTiPzBIDk5e3liOqkHut07I+ohGfq+cGQrmj5OhGwHDNUWtMM5jEASilYDmG9
b3ZJf17dgU8jWwmIVPDWfY/JmoAmGasV/fTEqME9z2iO6HZvX0Mev2UqVWM9BeXyozqyVjTvATPk
1k1tivQMXE8gQoZOz96LiRxRGwKPaON+Qe0LNzqaPDav/mJ5TT2ZKVM6/i/fT0/r+lzf1wc5jlhh
Ya7A4AeB1I61Q9R80BcZUmqhDcrUa69R6lzPuIbicZOot2JZSXIIwWHBy2KRAwHFFjbohJOK/WWZ
H/l6j14MQYcjx2YFmO1kjHTLoNt5uNyKQKhAk+UZMJJXBPV5/F9cRi1sMD810jRdMVubyukabnrS
q+c3y6AljiCEn+TBX38z7mavpvqwxDzRkbvfTpXEPFqcGPw5zXtPSES3ORz5qVQ50CRHIR99hii4
xrWo6NRAsPRbs19NLyH4GUmOfFUHpvbuK47yfiRGUNofvdv1l7/n7BenIm2t+YzpOg0Qa+8FDuBz
uRvgPjYYOHRrEpD6lo6XpIML7lAoIao0oBNEfcT/rsuebUY4GU4M4zOfcb6kAUp3ikXnsIlboWRh
l/XvbsC0Glbh6suCRD2llF/5GbPUveSzXEjv4PmuaJ21U4oyRB2ghPXcMgmakKz1iLrlP1W2R02C
q6z6eQ73f/dp3q8NBqRc/MdmAH9YhyRBMIDvk2RvbdBg3Cg1FRYZSyQus0ERaD50B4tgraramgC4
X+JUzy32EEc4ghjeN46LTfOy0HdzGFn1ObtyvCfaOKV+rAXjcCBB5o4W+DfYDMflkDatsmoyHX/c
Cv1dUVAmmA40DiJKfoNNQ47U0QIdiPDiSWu8VknoQYOMZQCyjPWoKILcQyQjgMRfGw+5aP3CLfPI
0j1HtKLB3GnPo9clgrn1ELihztl4wmTd0CbfCjlLNHN2N2/LRq5gYy9klRXEYjdqblqasMUnrSzm
4CmhGXA3cOgAip/4guoLcp9ES5DwvrXZcDDW/f2hOw8PSgP1wOIcRGZ+JcnOgqB9jFNjUAqI5l4z
pTIfJ7NqQsLZAd60fUjV/S0YEBA4OETz9SIIVJjdBIrvevWlLclogLIKZx0loRpb2SunqT2LUnuf
AGmPgu4HuKAjgGV5AT+/eJc+mLXCOHFx2BqGhR7bJija30/POu4db3qrS/rATkiWNB6tIbJeVhoE
ZdLxVHnuVHLsHljArsESU82FmZdeTWgwjVSWvmUJVa4V/ygh8DFF2fMFO8ZSxbwIgUmj7hFRt/b5
V/OEgxHcqdP5R6G3kQsmxEEOqsbNj/XlHwAMv12vueV1TWUTwXR/zp4kHnGoCkhB1bZjkwD5oqaW
sS+zxaRY51840ghUxSXWpY9DJJkqG7NPwyvDqCzChBGMjjQZydZEoFgqSIRTdkLI5o6lHWaPWJ2f
DLmI/hrMBgLADecwWEAfZW1VqXbLneCBpKzyNpTcXS//aH+GJ/kuLmriUbs0pqPnlNRjfryiUcYV
zSWRbyDw/KqUnEdxlTSg0hGRH9d2GtnPXIQ5IKGq6Y4booee9qBKViVnTsZ9Rguctx/aLg8kRSwc
0x9+ZyUr3uWXUnPP9snL9kqpjYKTikDCgTFGRokHU1vHi9XhYq4B7+uYMt6cN6iEZ1CKKdFE8TlP
fe9qVi38qyJLAEfbqn9DHfKrCoQJmPUsJTCGy0o9K3aASSctkb00C0SediWMYw/AAUKKqzoifZnM
n4b1SY50Zgi0pjw/jjdDAxic5IvFEX+YE05DFGw8jMcCCOETWibARxQiEzy4Gf+eAPdtVwbH6Qj1
6PLGWOqMFRhlfyqw43S0pj/rLibr4FJchzLf8/Tgg9C8Y7oC5X41Bd0Zw4ZgR7CkyULwabbmfgDY
y77M52+muFaR66anWa1NGm9mf3/cuwCuXZ/613e4sCFceWVjktO1Dyv8KpcEv236AF60m/5mXkYV
A70XJv5jh1QocK0di/Ssc/VUrOoKrOnc1cDMvZypj4XUvwdoC9WtQM9xU7rS/J2LJ2aFayxWVqcL
2tlR8BJQRz991lymCo1By/wMWdZKmksiMQqS5D4sJ395zXufWrQs+fvqLw4WHJgdCifP+kN3bsS4
QSHEQkpMxHp8sEWdbhZNk659moQdR2FLk8GatK6CMtji/V0RsO9IVIUr362b8zpPYwf03OynIgHp
yqYUdmsTx+OW6MSUhp39NvStBMoyUoGD4QRL/sbBptONv25s1xDiTx7q2fSEWmVqRtIZEDEko9la
/lpNK0sX7Io+f21cW6zfzOV524myGYEUlRX+hcG4LYJpjXlV9aZguIOjQd0F3YCJU7v4sHPApL+z
UUf6H2Qs38Cr3/UAEDrS+SGLY4TV6+PpQPhVYdBMNCp2MrA7KEKwK+eZ0mUB40tsLTPTaOt59TL4
hmey8FOtSRAmWvOpwM3wTuLXY3x0lExr0Jj5NEWVPx4Zf/YuVqAEI5LJqZmVIT8lCD/yPXLOHV0z
n0dYshRZ8YXDoTd6ZkYbeY57/5TnVtdc/z8q4rWymuZHWKS0xjSmhMk2lHITLxaQAIFKH4/imnep
3RUkWIMNcBSDEgT5T9wK3y8YPGsWi/VMYc/YB/o+DQxXMavlKzrkWtQzLlMiNEapwVit3aqwzOUB
59NxG+nzYR0N6E+yfNES2JqV/wW8FQ3OnA3oKT08wSK52i9b0bxAmau48eNpUE6rDGtGnzDHfDbU
GjrA6a6mjX3HTw6DFt/d2jyfJ2eb/XsttWSMI2/pjkhT19kmOQ7spwBR7HjZrzxK9IHWdbDNYYWk
/SKPMlo1aL1baauVv2O0/iMMuRhVPmBAp8XL+cSBIYDPaak2300lIw5eiyZVCmEUsqLeerW8FzCr
92BN4wdKMmDDW4eCl9BK8emlXm/wHhzFnya7vF/X31HkJjaCp/XPxjdUp9K2FwtQqNzMBSKXaNPt
87Yk+pf47h6GPWbHuhtjmCYl2nunaeqZhAhuq3A/j7k3M2Vxx1zZfnPSDAT07C4onDApMC8subWu
sy6/MDkBlCCaksyblLNjQKYRsCd1di0c4SiMIufIIShoTUO34jUgdp96bF8c+Df8XzDFStQmgbSg
96sbMDuKu9QLe4govpkFHAFjWP0CYS+6iQkIAkdl1eKeYs+kd2fpOJeOJkOfTJc12KKJGar9Guco
2e/mc7JhjGxrcVXeajHBL066VJyXn92drBr4XVMz7uWopuVctrdh2Y8Bzf22DTfosl11lVbbY0oI
L1PGz1BAggNzG7GNY36f5AyDP6IFyWwfsXAAIcykObd2hFoLQ8ZW/WEms+RA5uLCmGQO4OoPD9ob
HV3I6EPFlxg6HVfsIV8YWb5G3njTD1b9t9dSWxMn7LFdvKBLXdWT6W96HFm5Fdp5ePTeNgC/5gPs
4yuDaxSJviMOjxNCBDDyiAArh2bhK5OxXCy+y5ttVotYAQfGz301UW+ikF2YRGcFSCjijwfZVmRo
t8EuHLNNa4u2SI05TLCTmP45pv1Eyk0BRsQEk4ro+dvHy/c7J1ERarad8P5DZtKEecBvkOtgjU3l
813I31weLYAoiysoHB/eguAQLi2TuQFq/v7lP/Jgbm7YXfUD0j7e3T7nrJjaJKlOFMI02oprxxji
g3TNMXkNQZm8BQQDh+S7Fds2zfsVGUIICYH80UGXhVyk242vp5TcWXfkpMLj9qoHaXiq8HkRYswD
oaLSYACbRUYrU/n/2Ygp8Tawiy/GkF5uH/SjxOyjEimoUfqHEOvzBx2M2XHs+2jQyv9TlSYEA1Wo
eAu0+JdW+IWDM8hO2N5NoYmL8JdiiXkE+EBk02lSUKYzOuBJap+luEHFp0T+NUSI43zGj6eId89z
wg6n2wGP/nJbj2pO9fi6HjzX/EpQgrFbaORzEoj98ILYXBCLKstB4l+gRT1yKvRP9Oq9+tIz2/nJ
yrAsdKCcuBq+GdYQQmZWifGw1VRv07Z35SossmsaVklYVkor+vyeYBEBU/HHyELuvhMrTOzvTy9C
7rlHryDwuFA3pgWMpwGWucOWi50A2rbHc+z/unKuTNA4PNYMOl8YmVxRkOmyNB1tHtOdUPA2Pp3k
QJGg6ej3M2qEZ5bmMgE+l62OO/lZ2xC300tRghmj0FAy6TjITodD2TefBT3FJIaztb6fLgm2cBMA
bRSD9I0QEcpKfYfaiby/S/Ydkt9Bcc9DZgenKQnqhBCOnZqD83qjgFS61oOUPjkTfyU63Nj5XQzI
BsQ4nP8EkiWD1OAzANvVwT6IeYbHxjIe0iB84JY06Ag/qI3/OqQji0ajVXpadzdVdW8qIWgZgvzs
VyDrHeVKxtMfzxxa3ZcvUwslyFr9kCmF0AzHWZJJoOVH1TBRCQ0IEBRh8Iu9GIvyu/Bn4nSqx9Dg
p3w5ufS24R0ZtnTnyCr1JvxQeUzblLcKjhJPuYCN4CjEAPHj99TvIynapCGVjhW69qcINFITe4Mj
nW7fmMD7jds3qq/a6eD//WY2+wVN+FLU1Nby9qg+gDmUI2N4NQzoy3pgXJZY+ZKlHUxH0nI34b3S
ImcX7kJZuPykIZP3ThyCjVyE4RHjlrnIz31cEBvMpM6m8uz5tYJvIl9zwxLnV4F5WnwwMaZiLzzv
0RWYGgoJWFqqNnSeDoIKsyyit2gefhustq+gePkAhlve3I/Hm8SxHDh/wNaYWzPZqaAzDI+zbQP6
uca9Y4sU6msLBXebMRO5gu6zfPtc6aF0WjgqTv61L/1gUSvRbg/ri7koCZyDG/tSCH2ChOu26Bed
R1hk2IieVraif4g6QAWQD5mpg68EtKpzpCyBYzenFX2yvnDtK7C62clQUfrpSxHTc2TJF4klbJyj
4JSqe6zY4rNXiAfs91AH9qHA1AeAsv8caI4ewUgmnCKYo6S/vEEV16o/tV9H34lZiRtQdhu+QbsL
YP2hS6PX0hsljecsWslYd7TzNulXHTxUFhr2lKzA7BDtbOp1VBALcihmJ7fvLVmAVybXXqr9TZt0
jzqGkTPvSAMjGdoo8TIJg7du/DqYe12OtE8FLx7v3a/DimDnMTJRAdmjWC9pY1tBOEn9gLx+w/EM
vFp0cy/s7ZF0Ayalq71vJAVjtSlpkOBgtIF3MPZHcDAaE7BzbMQ/Hc/BwQppT3BFYwS1lmvLiTMv
yUxAIlJJja9Eg5amxOBN1hpNkNMMclUjy3b2K3W2dIoM1K+64VugdRONQWrxPuNPPupqmefE8k4t
yP61kiMI9WrX+HWmQSBgTP3u5Mgs2qyIjUKuI7di1rhaDPIrvRNJapEQRH6sWp2qy5QxcomufY81
dQIj5D2zoucYx/do7Kh3E8CG8b5g7uAc931xJgWV+eAsRFORuTFUAXofK2kBrEqFOS0RUEb/aMpg
FCtA2SshXEaHGDGDzG8xcRy1t3UgQOMi/UqdbwBCgHpsuVTNfM4DmpJ0876gLk2w69iXKglzBqq6
hed4Q7X30n33UdcbCBH5DUaSaE9H9ipNod54eQjtQsUiLaa7wQshQSZTLe82AHd28nvACXhrnK1M
ODpBV5uarwX7TkavrFjo8Vl1WpnBAL4/njqt6zYy3p0UEzX0nyiQBMJ5ME+RbFi2xY/jweR1WbQO
hUK6PSNuZ8Ez3kIZXBfe5ChH5k/t/4bJFfggosKWeFtxGFaQRVPJYUdF3hpm5Ei75whphBrrNiQ1
uRxnUBtrmGwG9W/b7JDzX6kZkBNmt4Sgoesm/Zhdz8uS0sa+jcbYGvhqD2/nEQMkdXCN1Wj4+fbn
4Np3zuFyFfcDB2Z/glb8NLmpnK6BFTxmdW5gIPcfZ4OplWP/Gje3akRJjOLkljmMVFEXPltsLbSo
iRZOtKabh0hhMQWeGlG6vwSKIRjeT2xqBFwXgqx0NnOdNB+d6bHqgdW3lny5kY47lCRT4aWg4jCd
3cjFKoyOqAWZelezEiYRuXpluWSj3BQKDLqEDIHkgqcX6LsPFM0aSffMzNaR7K6xXbIfBND99J+I
oiLr7tSUMLV6fwglk5Xjk/R0118odMO1QI8Bfoqc/Vd7rM2pdpMnFpv4wcmTQsIQ/G0c9u269LEM
/sF2qsCPrsxj0a2HIwHXUoq5NmcZ2uAyXd9D/eNm1pFpRhwrOH3GeURhSTTdqxC4nhhg5CB0EuSA
wKseYZmYXCk46R6pLK2Lrx9+fl7bvIS9LAqr4D5RD73OrZ9/HuOxMOWfnCcBp0Q55hNoN1NZQNOy
GPTtWFqmkEv/kLvoIShjvxpyyquLI/VAGWz8sXTHTy4hdd73CJeS70SVNG1995lfkiVLir6gCj02
TMzH56rUSzUfvZ67NnXc9qaPlzlVuVUyCQk3apUeJg4TTbJ3D0HPi45vROLk+BcLGYs004QSFsh4
MUYHg+dSAhQsSDO6dMgnZgiYc4TpgI6Mv4kEEw/FLr8k/CaPWLeFXIDMJ/tO5kjrAbRa+OMoDubM
A+e6aTrknMd85YuhDUsrp4MpDKFEl3VrD+F8GNjc1Pg+ErV/RmKda3oaKELXtdCLGKkCT2IlpSoY
5F2bNIEmqKYMWIqyW2QX81+FByiw3rKhjjuz7PWdBfUQQXtN8UEqJ0njoOs8YBLEAHXhMC+5GPXI
n/1htAQ/araug4shCSOV8+5ioRR8JsIuoBEIjUptWurL4CaTubVz+AYin506+2XuGiHzxEv2x+wY
qCoR8KMsWVlCAJ0r714Glq6a1i+W/p76WItjS7XUL8t1IXsAjHiR7RfwnoOuwOxdedUZWKHGnsKe
SLd4aVfX6C9uREO1Wh66ircgu7UDIIhaZkx9BnqMEJKte+tfe9+dlCaNVgqSSV6+Lp2X9m0sG62/
wZSjEtP/rXAhVbPaCNxL7eZvM7wclkssi5s9nGasKZBA+D58boJ1FEdtxk8ll1519MheOhujnlq1
TmFiOjhZMq7JXGUqrmhHdhRzX7csXC1NTXe0vQA3VCPye7i6lZ/6iMeq3K5LQnnjZkdq19tEWIVU
Fh4haYKErQdeVxD+M6D/hKYLPsvswObMnTju0ouGxfcRc2oSSG08EgqXDugtM4ynlO1C8jyk6lNW
AHFykyxTOLzFBNAbBHEeH1WYPBgA118BGlsSQMGrawYfcrKdJuZmGfmeTUiV1L5W1yu+QtELS7Oh
84kXsG1nYGInS9y4d8zGl7DQyHPeFBpOBk/oJDMAN0+iBqqFV5vNUkdxO+dhPUjx6dinpjOCSLLq
3LxeZQmo8BP0dMC+GFBLqr5+T9IBvf7FmXN3nIu+WniYG3XNjWoByj4+e1dX2pfGtg3uzM5YrCnN
lEah4G1cW9OYTX2Nej+RecQ/iIgummAXTdmSW4CAPDxxJrurm8lgwzXS8mfSLyZZGUUfbO4rNWSZ
37Fw6lZXoziiyX/OGFtPbEELvOf6wC+v9H1zOe1M8MJ375A/SwHlolAfhydDMeUMmF/rHG640crL
4q842AgUKzk2dGOYP1qOBzQu16oSqTMKJAE7uurILoZCWIuUIajwc1GhcyzRabFXogj3jQlWRUGn
104jFDLrrZ/tdONh5kFJ/Iy+gcUHEO96uvczvl9z9Oev/PN0iONSRotiSaSvvVqMtOL7qY8AMqQo
YXsFmpj45AhcN7NoyOMkayoNAX3uzzoU4H+bnoNFfKK9ZGAUxwJ2hZ5gIrMG2ls/SkFmemFcw2er
F/rkKNVUZ4j051WLp0P3MkidAWPCB6Q36l3ViDlNrtrQJS9c06KCSotffPIsWUO/7DP/5/qcdd3x
C5LP1bKcafzinmklvJ8FIP4DcPjSaexfLbw2zXGXyqkG4CSFKYRyXEEr5NiZbBYQ+bJDICKCKZeK
21VOIz8n2YEohmFA1j0ThTcNvssfIRjmzssDBBpw1acSSTh9NCcHJ+hufZqGhKsQaRl6FhZGlD1M
5l+/psXKfzf3sFe8nnPgrEXUqT4sNC9szazFi70jayy++dE8E6i9EkMnoDYwRHTljKGSFQgT8Wi1
jvFie9+fsp1B6gLN6j4krwbs4/7ydcOHrrbd8AL4+P6qwMCNFOg1S2enId1OC6h0S8TPNF+hOArR
jFKtj+AglBpMMpqfUc3KF8Ilv1a4MtEuXaWpeSUfA66wuB+3f6Y4dz9QMHyQqdW7YYOXyzioC7qE
Dx4o4/G0zHuxg7iYOQ2tSxFfavqPO8GVSPaXBVJ5uYJWH19e/lYPdUSn3ROmCAF8FDhMtp7GUdxR
5t+mXb2OBUxPQH0k1sWyziI+5uGg7yQgz0M2z2Ws0vQts4zo5DnnH737hcjCqSPbliIoCrC69rG7
pARN+B0ESw8yFBl/JOGcQQxvJw90JSU9oSy+AeK9nxowayuUSb5tpqiE0o4vDhFcH/N3COmfHi3W
gz68PQCZfmFM3MVCXYzi3SNDc0oKWRL6CysItzk9T6q9s8wI9aDJ91ws7H/fVtRxwf5w/3+ik6VR
cx49dIOVpFXBKXWR9VApxqsZ0goz4ISTOB2MFBBYXc3QtHdY+Fr6mlw97HNuGqGLizLkPjjNH7YA
kc+eyNowUwRkiZUePb955Fy49+9dLd9NX9Zuhe5uEUh+XfufOGhFMgT8yJxvX8lTdCU2HwBz26Se
OCazK3XQGRpSR+M6lt7Br+4/Tm3JNfAhnkKE72aCGwb1AAVaSlUyoBoTB94SmVO7mcoEsF+Dqfuo
r8mnmlAxEsCvJNHSU8rl5t8nD4l7pzIif/f6EVqIsr9+dVND+8Q1KExjeEY1QOePqqNwv69jT8wR
X6AVasPSZZzfzgATSnZ+KDRd7rGhupJoENq9MpeW9PV/OmIIxCloHy+lazthI8kbIT1d6kNM4iLt
W2PLnBDneY2fX0NOxgQSL5INfAu8DPmwy23EfVX7052qQeaaJdYsaTCIMHq4aYCiDhWekc+lBZmj
rIm6DoupDHwzq3ZgdNKTCluRf4w9k6oC4jBZ/O1yidDtCfDmuf/FHrAA63qVeYmhvl3PEDyxWFHJ
B5WS8+HtiI2Hd5zMetO38D7Hwa0XD6rQqk/2+zG+/kXlrFxCPI+kPcwZkWFqVYMxu/yj9m10ZsOZ
krjskoh3Rd8G8LHxtfSjk5yQ5gyV5ugtxtaxsTdgtoucEQmd36Z8/WbdhzwPqenGchIo1Cg2k9Gk
CcH9CO7FWi0G5lFWOEu4WKN73rgFWFoz1fIgw7AXiVdfCD2REQGnvKU4YnzP+zxYf8N5K8h7WVyo
niehHcPK3CBKgPD5fDL47k9/c6g5p8NwCsJmC0h5L2qxdon2BuLT9be7P8SqvojGTN4KU9IVtpd2
4wFmtV8w7/vIRVzI9PyTbxs8i+uSXWqr51Q+ah0lsziOX9qGAYOVp/X8n/M21M8rWystk9eVf9Qy
P0gY8cLVFxjREdk/f/8DRhovNwW2msAhKj8fHYLBdcMhG4hMKA3tkee/SiElyazv1C5JhOWlVOV1
+Bien7ytoJH639kjuXhmtn0CtG6dcCF1fVVJN630JnI1UiBCpbz3kX6qexLeq7teKHpMfc1jAGyG
6IQ4wzUHdq7MIgX5o4t4yOTaaLa40C+/ewtmR2/Dr3QnNwrQIfoHEwpP5+4AiS52vAyw/MeG8Rbn
7PEZ/jUR108Fx7HaAmRpwJClE8Q5T1CdEQyilobMwEq7VbRj/Wt1xsF81r1Y1xUdcgUj44mJtA4F
zZs4sU7b78GiUAuFrIysWtmmkpiFx1WHDQpymPjTofNEsjXMF0jET8vhiV2rYAbKtmhkbrzVW8C0
5U43x/Ko2zQOFpz2dtU5+LlXE8EVuzi4aDzNEpZ7EgdWb72riC5R7PIQxTPexnA3het/2exZvKoB
VnaXEnrCPdtQZf01zztIRXcNZ5syWHgP6vKteFYAnvmpigRSACE92y2UOoiX7H2EMpRzUvYotUjO
nDFGCJ5sfWTeRCm9xt4FgkWGIAR8k+5Df+2ocfaDm7DsJqZyvSE9yyDToZ8ygo90la3B07YolIed
bBS07V4iesTsRGB1ZoLsrTi/tATbdhiykmh37TvDyaiY4tzaEusN65YcxjHe4IHbM44Zse81JO0m
50AApPcAoDGBj4pi8s/dKo2D4STRK08Syh9iNeWa2AJ/65S4bN/1vWE7pdRcEJ2UKCFWynTxF21N
pUV3CcvalX3rY5WMlULqD8rkI+900P3Wy6Ymt++KMvtr+9XDFFIXwsVgM7t3zdqLIAq8Wv4dtlLN
8CYyslKDqeY+7aPWbIfjxEOK5rDnZnOD7XUnQZVyty/cKdLzrQrYSCHfyWheDFJgXfKxSnlLJzIi
LE9K1O0o6ZoHYJTVuY4gs4lnAMMA8VdhsoUK5xuS4hK2wFlYzcA1tFf1nIx6+o3xU/c5dpnIl17+
7S9JSjaHXL0HO/WEl/OkCIE3S6lmJGrVpjcs01VywTnhuLBLYSxypjoE8Lfe/ClAA5XolveFy3NF
zdsdXpFqaL5X5GnNnZStt6ek/k9UdE10upPLhIL8s1t9n8CbGMZKchIwPBrQF//zsNE1kX5lpsup
r18mS4IMXHObhwsn+P9RNe5tQ5K/T04x3b4V1/HWsrOA/dZmSu3v9pbzWi+MSp9fGLk6d55Ua9lB
CiBQWKG2AmWNx5YCHSp+etLSiSnjLf0D/PFoqHwBYRSGmYOTdTSSn5jmdYsE7ibOosQEuvUyuLWa
oSCRCvGwgbHQ9UW+CdkE4OVEQ8frfVVYR4phE2GOUTTL8nOaqQjJFQhDGQTeDdFkg3DYfuA56yjN
RrADqw2XEXYIyayrGWSCMk3U/LL3rLQATkOqrAkye+JYGzU5NIoV+PwtaDXAtfPsTrzq2pCgtDVP
ce0JEeo3SanXFiHPtSg+h5YhLgdDkfSIOCcwIaBRQnR7+Gxp4zMc9fd2o/0dJoOgGMwV6iUFt+UM
XiZXqWucF5rHBqsHzDNKK6AfqgPnz93o9XXynt+A5lmN3NYoU3qu/L8OgGdcIB9pppXUVeeUgIvB
ibUOhk9dKO01rGLv5+SMiez1t1oS7CL6P79tcc0X1CW3JWWVQ8b4p1p2zfLr/gmZd9NCqQuZG53d
HFLEJy9SfWAsndKdAdbnLhNpmckJeqUydIFLBpIKRvdTOPaphBtbAE4xn5hv/SMHxqxN4n7cO+J4
JCrXs/R6vXH1V+QKspsx5lZN4bJCQK5sKYRypTpb9U9w6eVEQrPi2bKv/nsNEpvplQyQV41MT9JF
lguDh7Fij6Z8tNPo6jRQjcGd626pIDnzRHiftsftWP/UP7azEYfDnmbcXWLDzNHtkLPzSEZ9QkPb
wVVxR7AXmO4u/rdVACod9XsdQEbonzNaDL3c+3qQ7VBMpEdjey1Uhiuxn854ffXxWPpwbBc9D9p1
S74fs1vHM0X+p1+H4/NLWt8lSD1FwgtfATSWf623zAXks1nNEaeGdFeYoD7Sb93ZlM6rveHAc/26
kUgjI6WT8UYqCH1drNick8w/Z9e5v8HKIyGCuoj4+fDQTI/cGTmWHicX7PVtgvJf+n/X8sG6yTG7
1zTsrsN451I3Aqx8UGpa/1I+ZtmorGjH/xXOdcG10r3hqJRJEF9BkmSLy3qQ6KYhkbjQ3RE29pP8
AQ0MprGtmtigT6osxZ0GcTWMxmg/5pubfWLAojguv7CjdjcGskZeZKJRU6zlPLuHUnKmN+xsBCpa
YwzjV+dAb+5nn1wb5YSJjjByp1aRnkHzj/d07GDO/NIaFgH6yY4sq/ge2fU07UR4THEM/7JgWw2F
OYRJpPlCjbgPRfG5RnoYvVt66/VT7tR6I2qO+XDF2MfVsruefoga5Yvnce+W0y5B1rHq5YcZkK8u
HQdk1lzV/aRkLLQVFFSVFykjQL4bZXkY3mBjrejX6I03Qczw7NGEA5kPF4DdYkksDXzq4zpqhxR8
ulqIuiUKHPGZdtRkR38c3EOov4uU+67SEmFE31NmudCfZwjwF6IEzFu9wMHJN9hncxIcY3kuRaKv
HrZnBOVegDMuVI8eEQN4b5IuoODGtd476RDTwUPTd8YYuFaHGdeItog1hrPH6WhXBsa+ZVrkYxz3
AP47D2Rn7e0z5Zjr5ZTUtSu/5t5Da1XpqJakJ9x3iCQIXT3z8axgq1AdQMFMwlczwpa8uolYWXAP
4+gGHjwNgAutOKU4g1F6BAhI2oZTRPQiDjgHnv7Az6DSqUIh4uUNMcTkYrETRI9RYODhqVve3cA0
thvkLds708qt2lpV40+dSE+NMQEKUaV+UXcqSAtoUGCAhPvi0rt6YuP/wBH88TeENGUNn1BWLeGz
YSlTsraO2Jkha3ZXlmCWNPRn5lkDXu4kkuvadRTdopf3RqjPFCtQSNxgUdeeymQVkAYzCl9Uoj4h
WumLXwy02Prx7eD58GExOgDWz8lNtJ+cVEbe2htiF+OtiRE0ErvW4xbCgPRn39SdEaccJaD11Ar2
STt7DKbjFm6TnZEcFrcHYNL2Z0RaKa2i5RFqQH/gssOo2+JTSDB1B5MVsXxkBnK9E3t7XmqF/zyq
1K4RP9Nohuxa8W76K2WuWZ0+tA9O5NuhJSd5cv5N40PM9z833dmsn20itrbWYW790fyauwhT2+1L
+t+kZV6VKD45pdmwxxuyzGtabCAr5b3kxqmOPPkax+PbjKF7ET30SbtPMDm4XhN10Tjp/UdY7eSF
oOQiSJJVeogWkQdJpOTL3+vgoAAxcCl/bpjGtlgkT/764rmurSdRVACPYO1yxklVLcNSaopx9Kqv
B8+PHOcpq9c8VVr20kD6Az9++RIvrkQ6apKPcafOWmnHV9MCem1a/bL0FteKglkoMCYbjjWcPeyC
WcXhGPNGzx9a8t/uQZOF/2h79JaHYzupqi1cDWCje+8pq+y28ih7Qcznqg3pdRt0eJe1ImhSS6eC
GieqvmDO6x8SpgF6/AGyeMDp/OzI8DT5QKrw0B+dzOf2Bfa0od8AOg5QGb2H/yqymKaAsEgsblgZ
QLLCK32+OaXJ3TNBlwrLq2K2pUIu/H3XXLHTqpw/IJMRbFJ0ExXMXIHONHWzITif7Ea/XbcpI+gx
scRFFtcDi3p+85qz7AFmCgR9rpIkNoZ6hD3E5IW/IJSHjyoxSHF8CED0oTaQrsRJbIrxuDYx8KHm
uWSqFaZEAa+6D0C4Uou1cVZ99B9DEKiV0kSgv8hopB9+fzkLQYLUWhD8QPfoFrhQlUprOBFcnW3g
5ywCU9i5exDpBtoTMSObC4yvfItfFzam3bptEA6/dcQhzl0D3jzeB1H6fT3iZxWMZJLXX23wqjYc
L+LlraJgQbW4M2EBTX+nZGJjjNLk5N8FPA/M9SVXHqtgDDdQJaGdRSHK3BMybl9LpzFKyrE6ApaW
3aVCxcjFLRz5RnYB+Ff1mKScGqSgz2wNvQkHfvFAvBYhrA+ycxamoAxRBwQ+mX5hFzN0afz81JdI
3/7tLuCReyDfV1hgyokOFzCo5AA23muy1SlGlpwsgvSlF++mR6v6XRijAFGI/FoVyjL8zkNgJXiP
V5+CqNRlxIgyd+hNt2qLE8RxSuz1gSsOqiCz22JgIz1KkaFWmlXqG3hNK4VcALFVAomepHPzOicx
Dkvfeo8CTMMPS5rZiL+x+zVf7LiiNQvQ0lGQD4SrzFft9rphybU5ZmXIKRVk3udrdJg3kOUMLFLw
eCtJaRUjfycl6nSwbvlWNtgLYbsJjBNvSLamC9qbX6qaoORzklq1eIh/rwA8226/EXQSJVtqD+AT
Vdu9dD0ycBJwiaZawnvNSc7KfkUasP75HPzXxIna9lOda30j7huH74aYpGj9L4vXl5J5gPvWw8bd
/PJE70DIbg2X0iTmahyc7l9NeX1SbxSKy/111GPH/fgdKSCyLChK8l3PfKV0hFTWmw1BG6FOGVos
Iu38eZhy5d6rQMsiB/EfgkPbMai+ijdFycaIsrn2dnYQ77A8MlMFmIrXCR172DLOuNgv133hWbZz
HNr34llnT4bDcjX4wTpsnSzdtFXILmQkjSYoz+qlZH3N36fpvluYxLFXxoLl65PBW7LU+UIn3lR+
T7SldtOBdORefsjnh/YjH/hJmC9Ou8ab02egZ8Mbn7xmsvRwDIrHaSsk2GPAdHVhMsHTIPFsbiT1
d5Alv7TyDN7744sRijxbNE7QAfrIscnv68p/M6szTe/rRkegWdaAztZQ7DepnKwSEiERsWMQ2mHU
vdxJi9mEekVihNeHADY7orEoynWzzswVZdt47Gt5B73kFhQflK9GqOgQ7QMZxElT6zsvMjFRIk+h
xxoXF19gKJmevGAwC92n+ZrbnFKFeTcFZoOXGPZIPYiigMI2vtt1dtn4dJ95KVtYT1V2/qHnQROU
lFkUl8+n2tH6jqMFFcyccvfvzuXBcFWUQ/RN9wSxgyYlr4BJzhlK89ym4tjfjWBDVkN6mM5+K3kD
1L/N8h41hr+6Ipx9AbYdylLnxShsGdy7V6wlyly4LcYUy+Ja/cQAxJkSBfnAv9opeS21zmNkw+c1
eBm/1U5hZJQ/UQRl2cuQj1AA5E3/EJACLXlAy7AZhKHYFveuW7/iSrfTapkfmfUoF/JpdeIRqP8Y
HsXxtsQ2dnheWSsZqKkp/OmcZpXZm4cJ/yOCRi8w8mAldDXYbrXN7NuwFUd+yUJXShs9a+mPO25R
olIZxm3+Jrz989tWm1AKt7W1qxoApf3CTTRw2hIC/7bS8Rqb4oQTFNY3futsopkVq5iGdtFknTWH
h2kc0Wpmi333SVDfXiD9eataL+DKTrOMCdN/C59BIuBxMV38DImK7ZiesSkQEHiPYrH+tadE/DKJ
YqkxCaDAm8N9C2r6TNYz64QaAlDpvOgjbulRRdu7m3j5/a7phk1tmTwkddHL/7GlaCfTQ+Q3SSot
AawNCw+0CJshyUMLwX6J3ZG0fUdx//z7Z513c3xzmGfTO/+9q+il8H/LzOhtmUr7z7kDbbpmwO/I
v6maaVznNbjkWJLNyuZMssn9DnN79OIMSLudqCxGRHl8BDgdNDPx1wP6eB8oHNolfK3FrhvRUtad
JFBu/22V2cr7eypthoTlirSqVYdU+MR/NpoqDCgVf6zFDBBoctbTN3at0oKeeBa0dtj+6TJmRSZI
tdt6qFTAPln6lZpcTAmQ93+orCK4nk1aJvI1t8HrWWgS5NI6d+3ZQohdAEw6XaLVAn+kK8C8yD2r
5s+B3dwzPBuaGpRAUS/+1ZoOFE8sDnjKdI73Ji52jpGjRd8NSQZ3K/1vSULGUCHtXrDMrGBSkp1l
CWvnZ1WtFqg9Fw6A8wV4F7e/cl1uZWxsq7wJj5O0vkEAeBZm2P6YGhFutLkYpU77ve1CrlcKqAlf
CqLxPgXMF928FH5d9UsATapaegAbLWdLAfrnwWLcNH8loJ4BN8CzYkPNLe1D0evZMyoR5l2/ESWr
ivcN4qMpZ1CxyANmZYi6OmHgV8olCRC+GubEbDn6rz0iZpbAAlXjNdOoxXgdw1LG/IOJ35DQVP4q
ZiYxXL3Qo9oLxC1bZIp4wt+ygmJ9yLLv6b1UkTq9OinMnLc8+YGInUsj2uHYAV2tdWdMvb10skGo
kpZ6tFb+ligO835LD8IY6o/mIjeEPyddqE+HFQRfw9YteeafwjGZgMSE5j8kfBUBFLtyediuPMos
W0PX4CbeeV5/N9H4iaVasPaLlhrmX+ewQkLL9AhQvX9vwECV+/NepGjZP6b514b2IQ5GgVa6Mmj8
y7/CD8IYfF4nSPcxLDNS8S+qInxhYzTYBtSswmJJrq+bIORNEIIATmHDvMIQWc2iOblNhsdB4HUz
CRYl5zhMCn6kg1fkxSMxIrfaYKdZy45+wTIndEX4sAAc88I43ZA9yj/xjNoKAIqzX83ygQs/F/ha
GKgbfsN9l7px5wr2/p1Jnyz0Y0QxIbZ1FpabXv4hxuoNGqOhS+sdT09DZP6JSTTf0lo7ljco/cAc
Wit2OlhWblLf85u4+r5jnhV+ulZCfZdBqdMKvzAKJk2md9IabdecQVfHU3UaGxgEcbVYiogTHGlk
m9sMzlxyz9Emoie2ecceQljwb2uve9AprybTUkHrddaIZQ+6+ScRz8TzzqcNgDZPYxd31TvzW4Q+
cZjqsTRcLS+Wi0rU3YTUXbdUM53ZceBRIx3TAy/yTXyBWddiP+lZnZvY8TKSjzXSJMusRuQLrkhw
lmGN8NSEKh/UDfvE0wW3p96cgaWP66rwqqu+TaqokN+8v82PSU8ZQ0gOwjY+PpcKZvaoyttEWr52
dnBxnYMhlWZlSW1QUSpqJPWzA/f5dG1Q3likFXVYCRJvV8yQ1L02tddDB6PCr0gEmE/knOPkxL5W
hima6El3gBNyZHqM67siXvFxZt6dXnhDuG7K2MWVYU5wlRVqu7PG5AOQABMjgNBT6V9hr9RzLmiO
+5LYcxpjQ01YW9lKeQOiIlebmG44bY3jG5ztuh0bV5oA5OnaISixkvUv5i1KFo3geksB5JvIJI0r
cD3ZTpAwo19tPm9KxVo1xOt6LCacgemmzwsnCA8o+KifBqTSGyQ6aGEfTDYfEy/cGbgfglmdOWFf
y9w6kz8xfHYWHae8C7vv0DGwOeJZHxjcR3wJclSz0vvgffelDyeSHlgWJUTA/ABfUJp/BckF7kUZ
h0RlQVBeKBDyf3og4DXEuFwiwec+2sk84QDtVDVw/J567VjUdzqiHd3rdjg6K0kZfcVCS/lVig0H
WfackODwG0nUsO4Kk0TNzwTBGoJ106hzaR3Z+O0b3zvDMJ0sY2rPLBy9Jcb8ttkNrRZ4CsDQot/r
xOO/UPtviXG4PXYHvd8qemx37Ne8+JMGsmQCGS9Q3EGeDITR4wl6+oez2q4IIMMeY7FfLXjrXdBb
WOXFDdabp1Qvwfg6IGJ5TF/3wVQ1uBMTpIy6IYHgG/sIU7LEeR51A3RbbQ+zZcjOlOJQk44RBWWD
MeuDpuiWRXT3YwZoEwLqT42pNMjEdq9ELMzCmFfa7QVmOD5cHjg2A0UTCel/4/r2Sgjh8U/64V9z
wpnqCcjrU9oHs3Xvld+jipdeHRff1IRPujiMFdahDmLPbugkM48JiaIKj6NZN7GV+WYxBx3VW7GS
7zPj67FHwXu864ZdQxB7kNDkQV5U8PvS/y2z6iybSioO7RpROLFiCoVLgkof9WEylUVjelBN1HRj
viPC9RHofrXE96TfmfIDgYFaO+LJGJW/sJEEpsKbTkyjFRjrP1djWuadNoAXPDXqxgZAlSBQPcTh
+XkdtQlGhdwaQtN5XAUX3X2UFGWVrmhoeWvf7sj/CKcPPyaIoyOrWRUdPjX4usXM2bD/Boz5/C7p
do7VTAmyvkO2PXHo498TMNDsStpqeHaPcOygLI+UvEPDNeME5abv+4bGvB/0THIodnzVmsGZgbDM
1AoQrfyAM1ceiXCluI14XM6jmGGnQ4iFQ/p6tcY8QPs99pp7OR21oPmiJjYkeXNT1FhVdjL59Yoo
QZ/ruqtZzjkjlMl0aPyXKrYPKtZTn1Qw5b/2lpseqRyxbqTVijp5GW2Z7eVp01R02oASjl3JxOkA
cIVo64wJRooS2+4NMdUFsyM44aB6DwEZLsgD61n728kdwcH7ceosEJH/tX2VIU8biAKOGMY0lzrG
7vVvof7NujzTzPwlFRsHIsspLQ5b4vaRzfeFRXEwCmJYOjIofZDSHYf2A6A/0lzzOTBhgsHv/yuJ
5amGI3Ff1wYrnPK9mp3Gabd/DatYhANF26Pw13UBdll041JkvJIuc2sFLsC4KZ6Q6UNUdQu87lLr
l8V2YW/BWdaXzOCgqBJozCD4hm5xDCOmUrn9p7JKEmdOJeDL+25Y+fKysAzWpMjNQy+xkCCUplM/
qwAgF3MVawIqSz7hdbAMwX1tgAusihSU+zScFYebjQUdt06GKh9WgjreItx+8F7i9vcJRuI5hcGg
jsr76JrQQY3mwj7z7etk2257xHQhF3EN4EVm4a6pEKpn3iJ8cqIlzQaa5ZegvGsn4p3iXcPcqePj
KH3tyyHXa6Q2obr9VcFAjZw5ScMp35bM1TkSX0t3shUi4fYgC3x6N7zjPM/SjikgnatqS77zb7em
C1bjRWUHVToHPtHrCIisL1Saqt/pwVS+kywSTtMVQmHoiQJi5qwGNsbyMra7A4eK+o3hHqvY3fEw
hXkv8HlfQGYnUiampZzB1o6d7lALK5e1mUoaa7CjITRqXF0t2Hnrpx5T1oLT1H8WAnSDV9CtOfwE
bs5V5Pzf0a7+g/aDV3fzBgmArUTdBndVJLRxeT5WDOSpG7/5NzeG8mAhsVK6qM31qWAtWVMYuUiK
UhdVYRQ49n2CQacW1PLv7my3gXZykW2Ut6jpfS5dbBUfQBcchkytEFxKkScE4M/CX7IseklDm5Hr
O6ogIHSO+l+2Qp2EoznyJIN96Q1u3CK50JCq7JuD5ofrC/KwlbOBAwghyhm80u0kMqDUbaLBGbdD
1Csx/i8tQkZLKyC3hzYputMgSCRVrNKcDQG2D7SOLchvT472cJnyGlsDbZhLp8cMP/I/tLSgQLl1
XfoubvbBOomK+pkYOemBVMDqLkqGAXKOhhnVIyzllTfl+z76enRJ6RpWcgGuHIYY1/RVMBE9AjO9
owLj8E+L2wQs9tnvmQcJq2JI6nor+2bZK0o1skRk6NYYI749ADodHzaRjpmY3BNwD5H6yw7lSFCf
+30VoHp2+5dHi3e+LWPlMhfl4sBjNATGFpKGym+god2iAinsLPu0NZI9Dkpg4t6obnJQDCRuVTNM
uI0KxL3euASuTz7dYv89Lcd9AJnYxPBiF6qqDFshoT0hPpoqKJODnlW0VSVBYTAjf98VkLlK4kLW
QSpMl+ue3VnymXR9M9IkSNCB6ZGitd1NQFxUisUxHu5AXTy6I4NARTU3Nx3UO3PM9KUGAmh1czk7
E1JQRiyGBJfLCo1GYLZVI9KimVa+LLxFowR7NXYPRODNoqk9Q2AuTGdct5S8vaAiLFW+J78ltVji
eHrtqh4s8T3vklnfh1fXZYd1BvXhDhv2f91GCKa2Qf8Z5jXxZuQEI0S9nkLky5IAfRBg0BLHVh46
w3vBoNJZeTjMGXnrT1+HvP1PDzoXZAtzniI972GUxmE04NPL60meBAGJ1colwgIy1OJKEClGTcQR
RXqtVJSGgGPcBQPyivR4rLn3Y8v9XT9UcgobowpeXARM6XmqkPLyW/4fJ7NaaUfXbBdnQpGrd5Hu
geQejQuAdDA2qvtQn77VOpDMv4fhOq5Byi1nTtinz8+jITzBswelYjXeXzOxcdp9XZK9U3WZN6Vf
f8OMx/BycuQz078rGbBS7PrZNliAFQWgfjk8aAvSUAS4xf8V4QIcT005ZVzNfvzll0/bL9QJFvZc
v6CohXR7gtNF7bVNtSiN/djlG0N8bwobN0Gr3W6642q0jZec0m+wyuu7qaD3vhFVyNsXUu8d7Axy
dUSXmReIMFWiFK2dM7fxagjpDASl90dSVKGpayXMbvNc8+Z+FZ17jDjcEpAyso8BxbDdCyQtmOaB
hu7gxjuGsevC2OjEF4+BtTiDTMr5A/2/IChNuIa6Ej9NsipAU8U1JDVvQTJqfRzzJsXHwV1A4W/a
pTgbHxLf5JTKAKKa7i08Jp6nThMa2luU/G3SKottrd+ct4JOF306AM2+9zuo22Pa5UzGFoXYAzjt
55F8yaDgjeJCohKoyMGIi33bLrA9pqIA39sGDosafzkt/Mx7+bz4OT1T1YbIez6nWgWpYg9/f5zH
eP978NIZgF7KnqfaIqK15yc2FZi2/kbro8TuAyxG1DcQRskwo33OpTfA79doXv84YXUd9Jj0vYB+
fOzTYrpTAeTFFnxyqnToG5//gzwf5szybwtVgxa/WePaRU5Kia8f51d+7p4qG+7cMN3sFwV/ilvC
obEZX3/NSrKBG124iMR9cphDwFmPJuRMEo7hYxF3aNjo1XYW2WHOz2ATd+5qEqHxb3jXngv5QOhZ
2Eo5L5bq6G1Rb5YNCUP5mVRAOIY5EMgqHVOLi3xsAFZ23IpGoVAeGRvHbZDn4CM6NRMONrTK8Cq7
5HcRUPmBMEtMBLlo6ZuDnE2hAPWTHq2A5+4yTaw9EWxwGLZ17e67HWNSgpB6w4GYs80m7Q0YFyJ4
KK4dDyNhxuo47dm4Vnk3S6b3+NGOMO3i47d/jvHr6ywM3tSBYZFTziGGMOen/GtAX0R8yO+UT6pl
LyuhG9O2G7U+vD+IMlud3/li9RlLFJD9TSvIl5h7YFhvK7boYzXU6oM54afUFTq67c6lTi4QiZMv
DSmx1q7l2PnCKIOaqx0387NlbocxFGxc+/6HUFiSnle62anh/9QvaCv/9BX0yG7Xc5q3aiXNOyy3
+Am3bcjEFsu+Aqu7AxxXMLN758Su+bVQVaUWRS6D8B/ZFycRJmQ9ui4fMNCWYFkL9t3SZdftYQlQ
ScZXfE78jBlBdUWDF3e7dSUVnecyz2S225sQ1U4kJkwJOysS83gwilyKdc+KYIyssI/T6grNFG6x
eUA5j1py4kzqTO9lwFaxu9iepAjZ/rz6fHQmNZif/zdvIfwBoKiYXO7hRPx5nzGI335o96cx/eSe
eBBmQiB5DLYx1AAMrZzto7OUaqHS1sBofhNtQ3DFRsC8AfLpWztPWvCzyQajOy8Kf3SW4STOyxv+
V9Rpf2dVD0KkpciX5i/uLS6SxW5IsiLq36zkdcIBr8KZQqQHGKG7uAOYOJf7OfFDXiTIqc+7cDSd
fciUqNK1Tm102YhvTz+DdsB7Z/zYaVVqODao4IIoKNKm16pj2WPfHwupv4J9zoiaax5uhqB/JFsI
9yFvUcD7gThgAfkSVgC7h4J2TkPdHWNZF4trQJEJpiWuqimpYgkcSLPdE8jagvGSkmXtPxursiu1
0TmDtDjdWma4+WGlI8Mub37er+txwbsILbDoIabalgd3FgxKiK/6z4q5WLotPIjXaa229Fpmt2Wt
GfWFdheRSI860Q1jUKth6NGyVJMyZB1O+x88eqnAnJ6awy86IuHcSVJvzViCaTeKsxQMNlcEFz3x
JjuGac5TJzRejZ9mLBAX+eEbrcuOuXSyJ/ws5smTGloz42JoQQEbH9uHmFeWSr4X15ugJgYVfvLB
Cb8uORKTtvwffMWQ/N6yYM3w+Oc5wEzzSK4teYxDuOP6+U8X03ngArfaauAwR7mJ6W6syAm3RJjI
n2I8AG2rAazZhfiSfKd/d1ZwwdTW6VB+cPrE763suzYd467ZBKIW72kof5Sd65xEJttICn9pZMiO
d/bd4qBQZIARBS0OoUjCZ4xPKuUJPQRE6Sl20W9oLEt3rLavJ1WFWjYZ56AArSUevIZqejDWP1r3
170yq1u7rF/IKYlOwuChLuZrRREgX5p8lRmmedbYH/T89k9NC15h7z2sTOzzm5f0FO9bOurJwBow
oown5xuKWpyCl3SR7GP7UnWs4JwJpqo52dhpAhLYqiVletLQN7BsH9uZufr+KWnFpBR5UNi40Ehz
agR5Bk246Occy6cKz5XkM1rs63JppEjOODi2T6XX8Y2Koe20Hk81SwnQUKcYjhMCsnN2swZCg9BU
vVg2yekpzVRYZUhpU1i2yj3sczGGqScLgBb6PbAhfapupdyCuiMJtTitn/fb6mVdu0Oki4n6WPGR
ETfFxa3r23EOxraIIweagz5H51YvAaWwTlu3hvMUYaCXfRlL7rVAgBRi4JaNrryMMciStl4e2o2C
HNsRBiwgFdDM6yVYrQ7gU9ZtKM4w+esoHr+dWS/+/r1aTK43emZN9IikMrPSrXIqokjhtAzfqWRi
7Ms6Iun7fIkDs+eOOtfEbUgNABCpXGm+ldI5eOD71f54d40cQ1oY1JRnUfVAXJoYrtGIXJ16bCOv
O3Ssg7ADj4g/pSyDy3OcQaPo6odY/647UTMaB50xR8N9OIX9L0K7BLFDDtTAzpeXUxudp4raX/Mg
Y6Y/V/fgx9n+nCexuF5kZ0VPBiBsx1f1r3uBrdC3xYwmrtiqOQvNLUM4hhGMZyhoxVWlfC4FkboB
kmYnwHL6y7G0CbJB8T0/t6N+yTC28UGE+lS/o25/unUtlSkRR9gu6Wt74iwBKFQjvLLx/xL2vhBN
B9fIbF97rUd0SB78bINfvRzmOxEFTHiWEX29SVk4q24uV8MsHtpvl8Awk6gDF6LehVmZD738G1Lh
SGTbngyj+9AExiZvjVG1PmbtjUp8JleW1FPB7p3zbWc+XsSqHbygWJN+8jCW4U9tFcUNC3T6E31N
JBsAYbZyYBUZrOJqiAuN2mbROniyUnEvcJBkllKM5xtExBtizenCZJFuOtFMF7Du4sOb5RjKfkgD
4mjnk7Ex6QGa7aIf9/1cA2inr2rO8dcLNlCuR9nBS1OtWLVarr9i6Bv4JnJQ5b+krQtj1jVnf/rj
LwjxLInEYKm8U8PhYGYJh7MWfZFKoi+YVEVETLk5t3uT/TCVGMJZjMbqxtmOI8mgixQQbRlUF1rT
5Cv2riTTrCteoLxtrCwPYaJVSCmLqhxM0QPRh2afTB5rugEVBr5+XNoWAlg6xJBqYV75gcrPZ/Ff
YmP4xF1aT1eJwNdbXLxfQgND51hUchpr8uUnAyi60R9MWugICQWweZLtNny6ChU9a4kSp/UR9XrI
ivS0g2hzpyWJVnnC38i5bI42S0oABfcf2WQVVY9Aehn7fW6UADL/GBJZfp1ulw3yTwsmDZNSG2v6
d45re+ot3wEPDE8MDkPozCxfsH/eSe6WjUI8VhD0YlDFC7HiYanNmZKRAJ4gce30RcjFemJNsGIG
7K3P0GJ/KkFHnstW8ngwM8BLMYItN6jyjA5WU0+lETxIScM0LCcMCRZiHzJcAu/nv5xz+c4CwvhY
vscL2QQ3tMxzf3/7FvW9csipcxJuQFpKmuhivouWM06H72+tx57BUMUVcfgZ/STwQ1OiDZT9m2uN
crovlP5GfEb1Ah2ElwqWIcd6VWwCjK/HYu46WrCXh0Lao/lJEnpqm5rY2Run/oan+ei/Jwfv1KOe
bYXQcOaXaXxiBIyZpEiLdV17SN0saJoEa/6PMmud3odMWXYMMC2W9xtz6i6uy7VxC5+HnBe+HVm9
kapQ+6h0BCVkz0gSlLQ1AhgTOeq2wWiIGa+ymaLXjmyHnsHZbfFcBF155zzNr3u62xxrBhwZjqQe
JRTMapyfYC2sZKdUKFogDGEXPv30rzXd89GD3IiBSgO5pepGhUkHDeCXhGDByyX3vJykjOceb9vD
FjpGH2e2tP4l+WzmvTrRnBSbwd83Y0xmd41MHj8NZkxKskdcPIRKiyR/WQRwEg3EfjL8SUHlZRiD
yCDPg6QAbKVh3Mu9k0QBRFvqzIpwzQ7rydp5O8WTe2t2hvaayr9+EYuO6JPKFrGfZClbeAUQdxPF
Kf6+gK3KlPUOm4vrXSALIccMzGT2/lqEK9nhZJInuurgDXH5FkschuZK2VN8cnr2Wjt4RSwtzGnQ
WumUk+UJJ+VJXuAPtWnAeSo/SLWtpiu7wo04XUdf62sk7bw/65pc0eva4+/MVMktx3/hyvtba86s
C4PSu98vc8gULznkv4tfeia0xf1rHFheIwkHPRZhDvX4lTIpihF4Boms3dx3YHRz5r+pNclDxQ+y
Qr1lwsop+sQY9Q1VUrdSR5RCDxTKkB0HHhZuqKe1Aq3rLGJayJ4RBlJ88fi9eyY3TqJTZ9NQ3tZ2
a2r3TmsoQUbAQkvO+tAGRhoCdX+qPvd5liHzqD000l4ZqP83C8C8+LjEiey9BUxvdPxkAOT++fIr
LHmLVRKILfguCKf6pqI6DK/lPHiL7zuP8n4fVNSotnGrlL7CgqU+nk1n2i/yi7CIqaOqaSVrqlJH
afpSrEH8tr9XX3RGvpi9BJRXz/I/Yx0HfWMvF2lkjHng4taGBn615ip5SPMR25t9KMF07yeSbV00
Z+b3RDzj7Sw9XAf/qoQLFDBA7Hmm/rfkTGXxi/viEHKqZyDsn3pkvgodbYs20xw2NdVkl8GQAoaW
38ZBWckIvyPtzIOXZnr8JiSLmD5wFH8JQOL0Jv1zFuqnnsHfSsg16xkdLGI/tFeOUD7Jlv14DxcY
Fc6GRqypodQvkQ+JHcwXWGI7MtVSgyL7iabpGlFkwir6uTYV1lKMjD01CKuXa8ctFthwHWOEhP5u
7Ocdc1By6jMH3qKfXSnYlz0phVMTT3rEipqQAoqILcAPoVF5iPvOUkKBo9wcMoq9XP31zJD5auqi
0vRp/xDeud1p33fNjyjcz8hww+QUapd9f3tQz5H1+CSJgR5PosW8mPJwiFIsaaWcx/2ABcOTQFRs
mzgiVIJn12j5UUvbDZmh41OEEtPjJz2yjL0AGWQplKHPGFoZmBjM+3gHvcqkH7kKF1qO93QfPZF3
VaNZAWdyUQ+/LQre0R5FkMx7WuP89aRAvBIp7rxNWRkR9y3KYL1NtFp9aZ20ynIeDhzayK3AIrhH
lMKH1mlR6Bvt2x/Zy+StDCsFEjgf/qetaweQoKL1/v8Ps+IkHmUZrIV8ispZd4ZdPpHmzktWgzb3
pHrcr4AlEYloS4xVghVauE9YFGeUDn72xcA2ILhnpOiFJuw4hs1i6kbUR+Llx0O3hhdWbIwhV6VV
RPlzktn9S8x8eeUgHZbygrUFlXnmEEvXAomccomylalZCvt3R5/u8Y5i9Jb2alpPyWRb9b3wsqCz
wLr6ip/VSMa3bsZoOyypNkWSOde1H/pOfZcpM7qwOjNPcmk/+bzKLrpgaCsMCADBI4F7Dp5GGNEX
qGZVMwso5nMlEMu4VuoopKRW1Sos51btNpQuvHCWP7ozWJ3jt5n5hrS1xTvGDG2mYcQ4wHmlIcWC
eEj8O/jzyRlmZdrc4kZnygQiRw6uOEMC721N0XRm1FK1v4Uo2QKXiTdNMsxFbLWdcnfR0cpHugvP
eygn/qG8ib5+0BhK0opgIkkig3Ir4Y2Ji8SnopjrE9rerHWHD66pTqkmz4VJdTVj1NlurXioUlCd
pDdnOTdpVikFrGQee0Go2Ub4tur/mWkugkIiUsgYup14MmTxSGhEjYzsyBfK3GRSODk9M6dEO8Ag
zu/zjka8/bc+eIWVpF61fljXhP/aK7BQcfEIKby/eEGt1YftgX3lmd3V7kZRztooxs1FtORBPvpA
L7AceT/nRIYAm8LqsYVeunppx4++xGoyRvC+G+UCJLZ8A1wiydTL+e+oSXMeACBDy0uzMcOg61x8
VmVZ1Po5VUemB7pTtlnbGrL4WFZueKpXMR1cGq24Biarhqcqu40RRcOPYUeu/OaRmZqVQ32IkaTW
uS5pl58kwJZ1EBos/8XsOwSG4YWBBOR0ShcoSUcvJ/9mvVVK6gIRB3aS0QuRdtmf2YiL9cBoi0uo
QILpASEJDvMCaVfm1j/8fU8zxoIVSOtInaaw68kxsQA4Gr04bu6i830h1QacRi9JEoD/3TGu5pVl
LWwTYQAn3KDtrL0cdr/x4ncBU0Ziul1lg48dPStscW3SrqTdKCNc/47jiUDhDuDdIlsiGF+N1ncC
gJkEP/gJuQJy7AjaQIWZbw9Pv4ZrPMkDfYagaDW24RiNKW0cK2f5xczog5V82ytsVtPPvVW9PaJo
DhGrx6UAtE4L/ZcN/TbQijUcElQmmiaBNLFWS6a1e69Ms9J7VIom7UHLpBpxUvYdvEPHEk9/Om69
lm/uea6b/BoiDl7ignxub5XuCrP7zobaF0Kn8ECpRGv7KmC7cX/L/ljtI+4WKuaflCZgH9+u5jbi
gwDrBrtmG35QdgjxFF7LwT0qh6I3sW4N/ffenAUE452CX8hPK8EDadS9/k+9q/697GyhSBnziAqb
d0fWfLRo2+qlATjHQdE/tgtmUwMOb3896tuezFZmZyIoDdwCjKn9jiI3sN+H0shaG1ZqCqNWrBGj
I4RFqWB2kJefsouPSRnRWIeFSJgNEiSXBosmHcE71Fu/k/LTEN+g6USJ737n1ZxKZLrDZS9vv3EW
VYDFAjeyG5T2XjdtR1Lte6xvzpXouLA5vjQySyU7zfNoYoBY4sziSKhpL9QLraanx1sjLenz7Ef8
vT2YhE54nQQ3kkFEudQccjZeowMTsbQzmEXjThGZi2gXYgrrJ/W4BFAqDIYD8DmsgSfW2WxJFFBi
tt/mWnaCteT1vcPYTM+onoffCfk88/Hmu3qMj9uw51wYfAagIsktz0yH6q0scTPhndVZ0Y6ZZ+q8
z4l1W1la6VFDR9ahYGqZOqg7PJ/MnW8Z4BWBLheroinId8blohm2H7pRTdanl+JzLia9fzpejaYq
km5PYp3mTQFXK+kmKxHyu+pSBe222nMWHY81+n536rrmBFQC7ZEcc2kPILT4epopgWEPu1YEbLmc
MOFePfpncKS8dvJjCtgNb3/FzqJnJUViGfHg75BHgzzYPFuAK7BFzQ+1nH0hTRVOWwJdiemlF9mh
A+z3iF4J0CWU6btFr6EG8kSj0zp5JWqOafLPP44T9Es0QSHbWn2CS+/vT9IpodPOznuEKMM/LfXb
EyydJXtan7LNCCpUOplIPAeBO7N4cU/30uyMtwFhxd9664awIEGlAMcJHmGVyVi6uuHdrGsHQb0g
rey/sjZPssPgxnm5elgxGUovKqjgyu1ZVxL3v8eGqhRShN1kRFJQb9AaISUJ8wIIrBPqeOiB+tmf
Haai1oP6eD/Jab6VSVJZOscevSbHtlz3fBYUpcowBOV3lpaEWE26aEp3s149G/ifF3h3h4yXlPJr
X0WU4ZVM+SEwHm6CK3LZHyp9Nnb+fuuIrsfXCtucPtbstq0pyvVsaLTfKWt/2d9X9T7WSVhkw4hP
CeFmI1xIv3FoX+ICkoTZ0+Q5+bR/3wvHYpYJU2wHrUe5fK827kgXYljANLsV3ysoxt7MN8eRsTxu
dzSv62ZVDwr9ZAHm7pExyz0Wc4WJJhy2FI5JcNvsQ9yY1mje9RUOu+3K/cONHbu3eH3LGHPGHG74
RZUtacPLt1epKFlfiywuXo33Ib/PYLI1yTfZb6k/Z1PyahjjRfSEz0yXAVJzW9t/Icv4vGVwXKRF
Jq10ZyH95Gkut2NaM0Fb9ozM2Kp3kOjKOEBXgsSEfPwXvirfxwm3xEdU0KXGFMIb3evmCDCI7Qac
QYvrRachTaw/itO67x05DtcGu/oxXfHGgWOARi/JPicIscaexrxpSFGgVUZCz6C+ZHUYl4jDz4O5
mCY+Gxq7Oj0rfqKc7aI3yYk4K28iBRogdRi22IuhhTcf/03UmxoTtKsMp0zS7geMFJRrg6coIt18
M37DUV+uyl1BeEmUIqu7eiUjIIH5bx7qE95NKaAw7OMLaGJ+V6ANy6aGGfkcYrmcVfWmBZxMocU1
njNN0UhDGdmxKMmWvca3ciyGBl88Zjr5upT2DyCzcnzCjeiOlQAFGWBcPvQq9Hu1UyDEs1Wzv4wl
MP9/HgOEQqLTecXnp4F0hw2ymhKmIyA3ymc9ezHHHnIrMBOy9dmqcdylpHJHySSJI4Aal2d6aLqW
uYwn3C+xnNfVe8jj2diYJt5oQz5KrXJdIH7YeMNFeLWRMq1PgUmJD6OOiv5SwUq0mCMY/Nj+OS0u
kDSNegmZsY9SMiAzkkgqqizUdidR8PP0lbTQbSG8RLUNQtbXwSFfRHDPEVFbmjfceBjcYjS3i1u9
1lmcbHU+N9nhnO/bMhcBflkTMAKyttai5O9bEUNsJ7L8INw4sJwEwjUhGD5fLWqE4dFqNGvtJ1j8
DDrlUQeuLCD62cveMpxeG0kO3ZkHodP4BwR02MRDzUmhFUlC++KgmkkkpY5A2v/PfZCDaGB7amGn
2DTNjbGB9n4Pguebzah2I8P5a8/pmVCA1FhbcNhT9zWfCeXe5bnNyONwZz5JflvkCP1DhaDHO8gc
SvY31ypPtaejiMZCoxVhePLQ5lmPdoPkFkjrZIoB9luI0lTzbDFFU9gexySkdCUNJUoO7TS502Bg
pOJrX/FCoZVQvvg71bb4y8fzv06WQslSX/6QIC798ZaFI+5JO4TOXdRg87YHFkv1+gd1EIOtXQxq
kri2Ge59TBvjA5PVe6bCK3LF/ic5vAVVwa6cO7Q3URcS40TMBJvvfvhIeNgHtIrwqjgRTNRhLsRF
HqrsMaY9Fca/+nugvGRqrjyJUz1T0uv24RtTeNta+5kJFc1y1TGIT3EVsnL5PYtuC9tailjxy/BY
G2mWPJnivsZoC5ZWhSFTwizgtLCE/o0vDv9hgs5ijgHTWM2TAAtCADZyEmKB2UeFqQyOmCx6KFYZ
Nv8BTsMkRs6h6Tgrx6ro0BNKPLU/HzDswf/Ehqv7zzppWg3B3sXkQbzGtWSY21RxtLnLjA7Cb+os
cwCo09xT9v2PJfO1WccZDywlVbgjdeyqsZLyMdAiOA9D30ICZwX/ndoKb4TWLNab2gKXWJJffnJk
LrVgCIcAqMLNwNvjt2M8wn/dqTJLt/joChwMPmNDMSa3APlPW19Vjlpi2vBFAhm3c/43uZvVeee9
rurcwJYONgl0bdh/zfPl5eciFpDfQVAohTJ7TuESNDVd7oFRcbYmtMGSICoLlEH9fYPH4bmvGTFo
3UVkgNI9yU3VPbxjZ82OxAArw/mfkcskJHxKPt92qZEtSz745Y9LyHK8ptTeFBjX3UvR9Ir27aba
LTJ2/byNerCumcJH/a0jtm63cXn1BS8U0mUWz11NoSg0n6uy0rHfQQyhibt8Zx3IsFadwCObhIhn
ui9+I3YsoXssVEZEQ6/aspDuWryjxEvAJaG/C+3lWhj7i4rl+KfH6eoiTIezgycoVPonMce2SHWu
nBdG+Hr2gDms7uMydPtab0dPppO/TkNiX/oAk26oIJnu+QpUR5Q+VC0Z0dT/mCYzA7IQMwOGygbi
K5SF3xocG++tk18x0ESGsgIg5nDZhmFDZFVwHG5hcpDtCPUWpzU0vlo571sUGLjfD+zSrKGK2ur+
nb69cHj7tmJ85GBPI9GTlZ6F0RA7gyQTrdeq0aITdat00jqfype/YlG8ISE03Gz7pam+U7Eg8WpN
Q1Oj5IaENBnPXVy3eUQKCWQdekWncTmovnHfC/S36Hi0u4Xzjs2Hu5AhExIGQe12cZRy9T+ZcXFn
gcOA7kVIfcOefVZACnZK97aiQSywX/EzWOIHSgxTsT/bhrg/f4pGHQQVrPaBtXl+V3eS9UcUT+lV
JHW8/edPVeX+a4ZQhhWDVhLlrBTsywp4ckjxJKZPTMMUIOySq+d3PZESaHx7S5cgSyIQjLh2ZI8w
9ztQndryYsevJzK+RrkPidzmh7t+BCKsDGbWIkbzDKHU1F2xqW3ffogt23hLnaNvggTs3vpw5Gr1
Yg5qoCoRc2FSKw/VVQ6Lj1T+dHX4B5GbOzldlPcWerIVIU+QlWhhnejvAf5RaRleKahsITxI+5lL
RqM48yvVbCTro0hL2Jzun7V0RKfe8BalZVLKiIh8LH/USD0pYddLWLIfeBE2h4PS+NaGkqrtORwv
eODYs/xJ1rczPNAjF14B+EmMmL/CCOp9JFBc7B2piv1D94PU8RF+d16mn62EsJupW3aip5X1PSfo
71HFKT2vtCSdyI4OAMG00tuVWM8V9xz6caoWjyvKh/8hiwNLibD/7K01ihaJryfUcW2POScYSf5J
2tw54SV9NzqweLqJ5jjPpsh0rvF9lXdUUOedzuVoxkrpAEsnjCvBPGURqWKDzJ3Kip4TV7KznGW2
DR/AyBog8DmPPs2kp/zkySgAvYxbFq5PeZCqj5XQwFwLk/XT2uKFeqgyOZihVGCqealw5tT7mwwF
ZeVPFgAGbzAkmt4no2sHeXQ7ZZfTcvwCz58mSK4kDPdSSOUgbeNoxYRJ8JCK9khKueJeRGQSvEbV
/mB61PkJ1vkqVlRz/Njk0Hp9bKSFP7sgUh9rJT0bXU0BQU26u/N8UwIosH13+gPx9Z56MxxZMP9z
jMSMhymWYBy/LwA2gsVvKK5KLfa1Nj64cWI8L9pwY6vKYfSybpTG2sPN3Rc6tOv/OZ+zDW1DSFVh
tFbyQyPb8MDIy/+7KVlThE4LlRINFxMjHoIlp+QMA4blR5j2+zq9FS+l4WCwmXWYGL7Hqm06KTNt
f0jsPdlkqCDniusARfUCM6NulhrIrGSs8M39vRdb2hY+QMxTcgilpBMAl28gHUUe47nq1vO/Nt2t
g870LmJpwonFoaCYd7Ub3MfshBb2FRohwUy/FI28cMdoR5DunwZ7V9/D4QwEAyuH3OX3of5yQbX2
6LImlDu7d+4CKZuAu+QUph0SWlcXeDudjyN5H0CvfNDUQmt/IkGAgIxMtCk8OZlRecbe8wqALMBk
rJOfUFY7AZr46YIb2dswIwQjqvePiMZK7dbFHys1YM2FxO56cw9DX4ZjfwYdq7DyGlj8I4OXUmIe
KQ/fb1P5/VwG5nudINGLyrRcbAytUuuY0bIjR2jvdi+btTCru1PyydNeMmmqd0gr6qo0xg5bYrIU
p6B2BgpsXM6o7jlmONv3tsruhveJJd2DYqwVa+ifJCouYirztuyMrHhZ4oieR6ALHmJrkIIrMbWo
IObIEW+CMdxwLlIx2IIFp7oEiLnuwE5Wven1QbAwaUPl5ZeBWIsVePNx6PUe4Pi0uc7Zt2lC1GgX
01xkTBiJvrb609jTSvyoBlbNNcEif08I9P7k7il5c4TdesfaExmfHvhLLQgUv0UEnWPvlXz1+rCR
rz/DlVeKs8E8hGRge0ZcEudiIlLI89Ed28D3QmFn7cVRrNxp1hev4BsiBhwwgrvWDk++ApThNuXU
mA91bVk2qyEtbxhggQTfRGBoElw+QtbkPt/J1Xb7FNSMBmjA7qqz2t0NfVxNiRb5ROnWQPy5eQp6
eLJLpNsh0Yl2WmwWjE7HMkwP8JYEKazFUkK0Nk8ru/xP+LjyPIvbw7w9Me7MxhF7ADw6dBOG/WO1
VsxZ2A10/jbSmLKkJu7AjpO74ZAB94DD6mFNPHy7sQ874/FWdgtQ33bqsyiNRDDrZmIOWydLC/vP
5GIlibJyD21mbHPhhRhQOFulBBa3MQ4QYyRhzyufcREHkjLLeXVeN3Gq/pYa0vKUYI3elv+JQckE
CSjHttNPwAwsUqsmBfgRnIoyE+lsaEma5u2tmbjXNXW2ChvHn6ri2cgVYK1Yv8eUWURIGColvAee
IgBO2zVReN+WOH9WBS7p/M/616gGM1E7D2lYKYLwfdYFUmXGQ6tWrQ5G7v1j9rAk2dInVOb2rQX+
hJm4LSr7QBZQdgM0lIATzKnm0MVRkrUEjSxKlNuIEqPdbn7XbkrztVpqbzPMJa9kTDYb7xg43GNh
OClmDiPqwvN9kKApygfXumD9IcNBip2rxaZwH6OuRxr/mDEvZhqKqeQR98oAiH5crUyRlCcvO+uv
+wkZLUpiZMdKI2JQMZlDYl5rHVxyDSh3W7RCiNlzAkt3jBchIos4gnALS8oN/uTV6XYKovIDeRoi
bc5ZMyREQlFqrPWNvNQ9/sn/KQdtwjfY8wWgKLBfnHbicjf+ewkTA3xqfB0aYg+xW68W4/RcX/Kg
tS3Z1vsHffRnqHnbMMT8hB33hpuPgG/s43APecjAEte0aLFeJZHS2eEvj2/y1JQNoz+2mRcoO1LG
5IYFioxeCfRnuj49brqaoD2QbmR6OiUW3n4/97uB/B3RVLeqgFIDUPh2QhLnVicUPb9CoTwi7N8n
zYnrUcShCzJb3icGPwL6Y7S/BK96aq7pSStOI8i3uS6WAFlSJY3OV0+yRkUIjJrnt8pNYCN+tOvv
0epWd7DCZCiGPx8BtCmdYMDBazjBsm62WmPlB8zNnMgwpri0PJ8EMD18DH64wqYJXRj0EA1yhwvH
mCRxffDrYRy47Z+QxeCdPdnOjBcnnNfnJyNcoaWimcPD92hr2mJ/1IyMmrGlVUM1kBVqbLfm4Jux
E2QQZCKtNJu4/ejPh34hFtLAab++AImffmTbAivhW33j1wXiQse4X+ewdOWwevcEJGHSqvprfOOY
nfASmLX/Jhj7PPmBQN0iKNmbKmaURjzbOHuQjCAJ2etgC2Mh87R0ND4W9l+rdxVupiy39m4xQX4n
RAQYQ7DvTdd9U9orc4PqOAxIry+AxkOxmkxH2QHvaStUanC2AR3avg9zURIKcm0aWFc9JuewwmpN
y6+UTnHQt19kAVuPVwL6RO3EgK1z1sCHEf9wnHmFfJ+Tzd7CAdJfVnpU6skDyRFxZh0Z2ArW3++U
IAzc/qIuIKsZNV0nU96hRmOkS2/CoOuP7g6+sNsBhx8/f4nGrNh7/EC+1jEFr6tkY3iOFdopnHWF
XHYcdISBY2WlR7+Gr92Z+4pV8gXYj+crfXmO/cVganzdA/RWNTjRZbGEjy/sIFlHzKRScsJsWcmN
aaWbZ/t2zCFQmYZW6UCw1IAktC0MmCsn3CcE6hVMT6KI2vpydUDs3HUA7UNE/qedCp5nLcPy/8PP
xPz/Sv33RRlsztbVj4bdXR0gy0st0zFYETC+t/ytE8NaPs5kzVEze7L4s+11YYigJhXltvYgHbuX
cbJWDEI8tYACjjuJ8/vjIS1CocBgT8ziZabnk7aEaWyB1mwA7sjXL/qkE5rcJVtRvjFypmI0kLym
8/RwNYn7xWtVHjxCsZRn28BPjt+96VPbOZOpgod2CXVd5eGGmMlI++r8+qdoKyiNTHz1NtNsisic
jIYDLlcOpAGc5lN1gVxP1jafJ3dED4CXkD5iILKS/ITRQuzQrPT6SIv8XL2gT1aLGM6pYQ7wgvON
ThOYhzqi9bg3B+aLosttVDhTIMzT/C59XQwcRzvCOu1LLjvecC27rWLASxDjCO3C/PpL2m03o098
eP7lg62VNYmS/awMQnpLs+NGETiicchkM/moLmEfoCg7m9xjTYeNggCne53iPByKAFQruJ76W2J7
cZV4KhZaGJmWq1KE6GhX5B9g97Zi1nrVbk0wGrV3ZtHOKs1HnxR4IPF5qFm8LoWdMOjP/xQ4qfNu
RY+a38eXN0QybkL037TEwSF94pjEmgpL/1BMO5qiFiKbJr3aKbJ1MG8ELSP/p54arSKkBX84t8/u
xv55Qzswdzcw2Wy5tD43YhsQ9kIxTjavO3HBVMRMyMnpakrNf5CdGcdrsyV4TiT8O7jITpXX24qB
nbl2GfUMy5pcDBqMdQhpgc6cp3WA57fC8xGbT3pFNlwPo2bMke5gkGzeYJJEfwLB+oNDyXujQtAx
k71xVdRc+nbRYvpP2PCJx0jfI2pMGvhXn7hAMf76DGO5eNRNwlXQmtgcVJjfk++mfsWlOAYUyI77
66IrtadPLGESBH6/Ms2WhmgloaBfz47RTLF4h5I7N015ou3LcQegXAQ8SzWBB0lMlYKAy82AOnAt
e83ipDHDfQyaSc+p6ZgyHhqaNEfUHkukPFXi7NGfTVFYmSmPPIpWd/dph6k736Z6Cl5ZyzVXeQjk
OIyYNqm/j+49Z2rpEg2CB5XiDAo3gOGrOlzbp2fPoHYxuDB9xqBRtOlvQFeTEeOn1l2XNF8qHiph
ORp/nnwdMabBjVAwK3Ui1krkqrDUJTudWV8vM8+Lv4Es6lQ200PWr7JWC6MNh0NIqOQEcC9TtFbc
tqdTvMsF94Aq5ybSi9iDICUDwk99lNOtagtSDkyIjUPGRhZsgP1VKSK1TUzULXmVsaWH1IrHGjSU
ZpFKlimR5DHiMgt40TF9RyaxlLmPcLfUa59uEzguJxLzwP5U8bolcVVHiIJ8Hccl3BmX5hBLD489
1omNP3MxphMIfLNG1vz0tDWtnbT2lmHRsf8bBKVht92O6jG283iaFRTFaOHnEvx6q0aPj0XzuwGP
QAvAA4pFMDjuaFcv7n/qvmGP8UcUJx5X9tlmKmEcYVkPpo/NvkSySF4WNuJNs1F95RxXU0+BfyOq
FA3eyt6Pm27q0QSZ+Xdu7NQCviY2iDQgzt0/Z6qeQGjn6xi77JisCpUhz9G8fF3xGr8ba3OmiC/J
YPtBt2IJlxFJRDDp833P//9dYPw/znolroRS6Ac0PC+gCj9g1Xmedkk83fMn8Pavith/8aj8KI9C
i+tp8e4mYqVcpcGhggoRQeF5HL6Ni8OjDHP78TmqKkll8+7+qLUSTNRf/GsB7Ae3cIt0u5smlxyz
BYtJ9rslFuUir4TuTHReCljmci4OT3n8ByEpdD0pHAjI1y8xg/rt7FD2x+fyFHyGO23WkZbYg5uo
BHypAxh2d4eCueQPLhSWzfj+4tkdwZ5U+caySb9B3W2oHeiBzYpvaiv5+svh8ms3tln1ou7tOZLn
eVMze64ZCmkCeDfeIce3OaObTL0JZz7zYH3zR4VOCJp/bbVQu0nGJwavlplnPh5KHINNzbaHU2mE
TPkJvCEXV2fyFXHyWmji6f7TdEgEacnBmmt6w9eF+l6XiIQIiwigIYVNlXOeclOrbN1AWp5fcxkJ
4WTtGZYe+GkD5vv2jpmLll40qGPJ1PcuBTADJG+NE7tDHjlU43X41FacRcgtbE7wnBVQSM7nZxMI
YG0G5DGy2yHuXZStkuviUbYiwWOktmHA+/MMgh83+5HY+KTjSogJmezADLDEpkS+zb8HI5RmQxky
7gdMjN5j4hTsTSO1KKwEgEBTIb1kfR7B+Xtvkj2oSQ1QHAzWlHiWzQKbsQBliXymkxSDOPQR4Rl1
6JqGnhdjOsrntb9Of1zOCROvVqaGZ5d3ZyVmyFuIlley2FX12hjDicjuikUveIIofQnAaza/Vyg7
rBdY2aufxWBwbb2hdu7MpuaapoxgrZu7mW5wXERBGezei62eZYoSW9CpfHoa7h4ghDF0atS30owM
bMJUszTvcGn85PldyWLIG9CVGH792X+VWXsnRr9xAsrI7q2SGel9UtDEPcN9JMVRNvS6Kxcuz2tL
PxRHIVCz1cvdGvlZl/dnx2qMNSu/Bxs9aNyXoJURKxIOz/sD/pHb6iz2MitYl1zrw60j2BdtTR3g
pm1UFUca45C5recOjPQ3cFUA4s+4J/yTjsoejiHZsL8XDTRqucC5prdnADAyTSRqPrt1RN2SQdaT
39iQow2ZtW/SuuCTlvST0brbt0ec6ZQ7omDKuerKPYTvXtFdkuvBDenijaO75cocwy6ZhPqCg1D5
6X2ukT1tIakme8hdkSAyJMVxobWqHNAx4yro9QGo/8c5eKUbjJWb+blw4ebhJYyCtheLsdHmpns9
8fW7WmnqWh/9Btp/T3q7z7AuO3hDBjdoWBhm9Dy4xKUSRrHY//OelpSGzlhN6QeYhN6W6yDqC7aV
pc8B3vm2lpU1TrF+scMVBlAFu/bs4SNqT55GcxQr1p6/+N0OLzju1nHJjaZuMBapDa+UBgo1aEp7
sw5eA5eAZ8usYOGHhEpWFKjehQ+0PljCqagBGsg3MCxsrUUadJJZvp5hcE197OB+Zei2y7KETkEq
SB1SNgVxWByr104hztrGvh+5iziTYnE3ww79yg0qefDmQY1BcNfGz/8MBrbwRGh6fJSh9bLZNTXL
wur5Q9/vNXUlpSA6eJ4qIRgFDUm13igGTFfoCpo4wOQeLIkpwLunjnTn9A6v25G0UkJsqwEFJlmQ
vQLdqxVpAx0xt6LnSslkayXCunsJqOhEkcSr/TMJgCJ9UIO2Y+tV094xSV0dSX01NITlzDTidcph
xVUJnTb6ANPTQnFcORTNQ+Hr19Z69sirjsZOGHF5ozlOCFBdAlqgZEU37aDXQRn3FnjWGgTgL0Tu
n58X56Ba81PZm5P4Uhzznkw6Q1lSezj46k5EQADywRH/mZBJiYE1mnXRJs8DEyjc0gqSHsBDwGLn
P4zlegF80LNkehNYACAeZuWH58GxCPuEuRpFSCqCZFQCg4si+NwJOwLfLJXwNVlxWCEGl6dZ9QEo
Wktaf9EfqM7NV3yaDl62LIzW9oHx7nssErQKA7yEsBpHxtpF7/tuq6m1MxiMQUy8Ei1ZaF84MAnV
nhxGTtm3ZeGCrloBXmHFUagloawTU1Ood0Fx1DldU4n5RxKrbBRZPw6JAXcErBPiFiWrrJSrtNBY
7paZHA5CdSzBV5s5XyK0flnSU4fPIgdE0Qz1UWte3xx9lpUa6PMGzCM4bsiXCEtduLPTS1NkQWrk
bHCWNLFuj1p7euXOPFIY0Y5mt2lEe1+MBuR2B1epSA5BbrhHmliU3pj4PnUY8pBPDmnHGX1vut+9
hDiJkgg31V0Hot46hnq/FjvTcblVlYMdFVG13daBJGrpGRAdV/8nCl9KuJwmlFc0869uu6JWQ1K/
Vfnk+UcXExyeD/xwCsaIhgL4Pf2FW0pqL7CuCumEu3S8wumKEQxnmHodWpRvEIp/wBbHpH4j0Ezm
bNuwy54bj0YCy4m4B8JbXgiHyuMpa1YoAMa4/HdZ+h8hS9RMrBcnfRP/4VS1Ns32FoDPgARlrmxa
+p3gbuhsYKgQ3DDY4BP/Tj+z8kq3w/IGeKsQcybq5ipVro1RJkOY38V1+kDnmXEaRuXvEkrMGduQ
X4mUAXndbbs83PsEVHMHpaEkttyubnTJ+uUhuL9VnoEst2BOmyzUlHrMSRBV8ybVjnAolRY6oKa4
yB9oTCPsszCetdqBhZxxnIfWr57wiEuhco3IKcuXn7SNjkyB6Ckzp3WX8lMFs7ZmLYO6Z6F0gvP4
A/aO1xqnnjQOMNhIK3Va5jqOi+MlvKPCTyAmPFxn0+lb/8m4laQRqCPuuCLic2qrmnqU0YKvPHPJ
jUPpoq+YjQ9m92hGUAGAF3pU3/dCHykTymrFHVKsqr2+kp2GfxEMSu153+bCduNqe4h5JVTSPy6Y
T8swJhdjvDAmZ9mB0Eqx8q6xeWZtREvEQb/rZDBZnevXYpuHe2iTdV9E2warbPXtEvSLL3GfRn0x
Jgbs09raovLKZyu/VTrqlWqlXFM9UitXcUTAz/uYw4WFrhnYhEjaF0zsQca+ixSA5tiXWRWVO+oE
ZQWPuLFw7ePe1lDMDz1MT3lB91rry/TdjO+/K86qmDYkUbjcIupvCOEnBaOe8aHHR3yhjk51fP7b
v6cILb5mVw5ZLGgwhF21aZ1hma/DZIGdQAxZLPTidYiQRVNhpfE7W2TRON9vW/XiI08gK+Lo9RyB
+fhbeTBuy9sFM7V0Eu7iOL5GdMmElkzLWSwAg+rs57t7EM84TtRAZHby3o3JY+Ak4GzAgw+1Q/2q
Z7pz160Y3PsnvEsSdsIfu013tmiT7Wk2bbKfSUkeqjtJGKXNgbYiUhMEZ6JqHKbi9ruJHpkU8rIB
DF6tfbNi0tm7X/Sbp8cJnFH3gZnO2nyK0FdUijbNWs1e0BlXxho+9LtqCTJT9QyEvaiADdPH4Yo1
io3vx1kzFOUtB4IO0TQc9MQG97465guoRmar0kwvvHfN3NVIk5117C6PZDjM80PhAS1vpmYLjZw1
i8euV374Ma9XyjRnMDlK1Om61JCZXOQlJre6/AZUcyBqNnIp1iYg7ThcOvS/e3f5Ilxo+rs7aQrH
RCtq3bRGfY5ksh/GsrBFnf3vMlkOzYmHwna/h8/xgBI65f4Hjey3hctdjT4p+VbV1xMpQeHLzDuI
VPUwY9ZyDPIwIoxy6q0FG98d9OXAANDh6cVH1O5thIQXlIC4Fe8DAC6M/TunSS8RoF+uPlBK55K3
Q1QMcMvXScK3Nr5b7HQyLM26fwOcgVbUDjQbnMxfLa4j9V/NilMNa4E0MKKN6V79W6+8y50rYT/p
GUDs2HY0nDuGkQ+ppUVSa2l2oustIOrIaLesXgl88jr7O9XpzpxhZ3CDC7RBjvaA7A8MtMkymEHl
YWzirEJk1HE4kQ7k6ZrxiUK0ACXzSP41vB4di3pEoFRStAjbcpqGei0hZlErHtkd2j375nG6gQhF
H94ZhWbcprRBtvBWwnOdHXi4bx90He4Gy6zgf8cNqzK0HAS3Bn2+0lcj/pKLYVLeZMjrHd8wzcMw
PQ6gDMtmpEC1d3z4+kLmqOKZNMA5R23SDqkkgmc91XS1w6lbqIBAdXzhORCBjQ0sTrIgKYxnNjAw
8GnMQPsSGVu58F/4cnbu4WTfitA7UPiDBdRNu1mImtc300i5QJ06qyx+C5XqH3BrFk0SIbfsE8oG
Ea5hsE8972UT3D3SJNcvdtfrCunBNeZ4n3z8sw/scr/Tnfqsuh8V3xQeAMXZ23+SRFPEDFPYiAPv
E81jU8VObMj8cDTBuOgM8NzUMZpy6xvXVgYmVleiGOZLP2Qtqsr/EsQSoAN9gYMhM2u1oafd/4g8
zFwn5zXZrXeOQR5SP6wXQPisJ+8//R5Jkqu+XTM7OdHaid8GCMoPTn3+Onm1g5voMnoOIvpNBIgN
hCk+Jn5RKTTuduNOieUf53lSvtzFBhX9opShRKxfY0CC70nxxNou9RY5go84Xa6wzpICqG4RcRhI
pyhmhhm08AXdWqhdCPmSJaZApB+7PptmrxgO0gTWmpGpAsE5SQTrpD1WiK4Op8mf4kRx5iPXQRZs
uiL5TewMOAmZvsVHmy0CtEZ0pqIfDSfxFl3dTb/dbeDza8xqnqAsveqViebtaWTbcReW4DJnPXDT
GQQBCoUf0+OGQVtRBAxvrARDrqJVJja8ksoEVfegGnAkO8UIF5R3bB/c7pu9vRReOOqO7chQvYfV
217H9WEchGtHSfocaDBc1EGwV4jn1YZhD2oPg8aptg9WTaz5E/+oh67WZJO0ZOnSPJ3SXLd3jA5m
MlzMqhGs5MwE+QFy9O92fXEKBLW5j21wNfZIEzqYGcjNrlerwEWkW4e93Ye/MLClx5OWY3m0tTTI
Ewt0BTpjBgVvV9qTiQmEpXquc05p/H+Yg+TmHwdu43V8dUOpX0oJ7n0EZvPzs2fbprgcU8NUiZGO
4j0oSFAWSurke5O0mBdTeNDGcddNkyoiz48vFk3R8wgo1j3OqHLUKy5kC85glHNMq91/8YDBrSIr
I2sJnJlP759D3Wv5JMNy/c6cNcTBCZCANJge9/Zqo40Y98zq/a7DhBZqjScLt60JfUeeCOK1Hp0e
qawG8ShVJdfckac1UVATQrQYg7Rrv5cnfwt87iMgURBWFPKp2bmwQ745e/D6hVbULTUxtT+Ryz7b
Jkf+E13sGd8VTrhHSzxSbR4Ns/r9ARd7iw1x91GP+FmQr0JMdmeQSVHv6Au6nvvKjaa+cBtIdWGV
IG8umz1yx0FCbdRl3N9yOH2tEBewd03/Yh5oX4oZfNjGF6OHOGu8Ol2KuAInqzoVIeqQR8eCdNRJ
KcdrAp5iyN8e3jjTsziyxC6Sn/AqDu5wOAjiHv/KuWx+gNO73pDyZmia9Rk4ofZSsw6DtbI4yOK6
jZDxRaM5NnnQsyD7+P8M1uQRnTh+g8xwNQcOwjbzO8tL4Q9peJPA5fdmSxmdpzDrRFx64Z72J5lQ
9RcGyztwgdXk4asqM8zGsZ6A9rmlXP8EYt4gF/W2rG9usy7Sum0mwH9EEL7Z1k+85vG7tSQyVVJC
CGMXrSZJeXtf9wwtbDhkuhoMYGFflLmv7PO5epumD3vbasruwUYB/5mUBEAZiJSwNZsTIwGsN1fM
XZv7Za/xNJsL3CQufloh+LAIdU1Jf1mLa1kHRgTnynb4CBn4Ivx90yKHsGjQYZ4pjsbd+Eln1mfa
H12VKGsRBNnhAgAfkX30p8lYqvVjows8KJ0OXoIeT1GspdsSS5q47dOJF4jHmYwnuOtVtLldS6Kg
OrDZwL3w2DoFSg88+6ECh1d30sF8vzxrgeuN5I0Jif6ejo8yyZF82FDp0VOIvC33S1ltoau8LlcX
FYX/v7bzL4gqlDtxuGb2TroMXdBC9IPD3FHx7lUiD4AB4Faqmj4EP9+SsaU/EBGMyxYRY3aeY/Bv
jgfAWnJJDBvuEmOhUVC3CK0/yWHw9sannuj42y8GBXO19F4h4LiVN6/2/UXq/k1aWWOOOLLMWhk8
SNNXLOBBggrzg/s9piBrk0oRsfWtSKuhU5SMY7ftqZuRnkbGHxN+FhGVZ6/eOES75++noOLWXCMH
X8aMaSaTRl87ircq96rTkL3kWcQjWvyTWw52DeRJjXcKPemUy/oukpvejItQt1VuYLefeQwZby8H
BejvsQ+t/3ekIgXF4Wqg8k8F6GsY32X9XY1Xf9UyDikiZkERNKKLYvuvn2b3I5GGEhDg2jwIzFdO
tRFYdMur+hiQDQ4vBwlVGPlmw+jMtTFNwxgOJ17RdU0RVIdimz83KO+qyHVC6X3oCtEsxvIooU1Q
HsKUgHO4N12mYJN0acxvGVm4NxckMvdi/3oLG1azLmVsBtvsi4P7Mck+7PSuEIx0AFV2MwgxqNNO
fshXQLrKu/LCpdQ5v5YbIJjwltawo+G6d4y0Dhudv+Vsvot9hO/LrrykxDMQeMuPh4tuLwumtvCK
CuQIX4mVqzJTv/sEKbzr+g2Bbq3iW7gPAUCaKjx3j8Mge2SeUlpB7jJOBICEaeMRivyWvaJG5A44
MrG7Qw7rMoNdwKRurNVUPLd+EQpytlio+YYk1PasX45P0K3vMAtdioYw5c0W7DQe3qP8AYsYZtRU
nnrup75fORKdfJpKkFlmOeQLFx0hHAPqnIP2MlgnDEacgfpxqHjg5JHXwijJ+BKQnaEqRg3vSWo6
jAmc1Jv7vQ2xHKqM+TAMS2UzodbEGqVSSXKYdg9hjesUvlOXl54YxdVaF7obRksPbh8jj25CbyLb
lWVTpDCjbwoac/Qfls/bBoXZ2nSfw8+0k1XYq/CzCXq+8I9+chnG6ODjWaS83cRUJBKHFVO8DoN/
pfSGCXqbfgJmaRMjF/VbIrmbDwRALxGK6xc5h7K8bXACb8ohOJYZZ9WkxZ5p0aSUnZ0pYjpnTrxe
scIqPVz7okbvf3RxHFy1hk8owwojfiJa4A8MD4NhDAOyjMexHeClEuEMjv7aO4fqRI+wdrFqf7cM
u+PYj0vE7n7M9PADw3Me+k1hBWJKd1rxv5aQjK7ay3X+J0FlXIN+cAzd3A2JQJsr2n1pL5l5y1xS
dyo/4MNKoYxHHiH5F4UUNchjhAWbhGKOSNYXQegsacSxlABIcd9jg2aw0YaF1DmsrYagkzVgHR+y
0TbLZKW9zh0I6AuhP+NVTIWBPkudDtsQoTTMeaI06mqrb6Pb4q+ZANLFICap66LOtpOaCNM8p5dp
+lHuvFujX1UAbL/qrTnX+VH4yv+ydYa5iNtxcuLjmHwSrWqmRa29D5wVe3oKyNZF3HeM53MBrrrI
Wfw9ljL+OGgqB96wXPndXxxpu1p5Y7kwonHG+rVyv3YViMKyFo2Q9bocfjz1cUnWiot6EHwupH1Q
O9dws1suKQDIapccU486+9TDhFhLHl9vm8H1lZBIg8JZEvErT1SfkWCg7O+/I2h1OSFG6wTz1q40
xBE87H3lUGxQwE6URJdq4MCeGqLY3EwxHwxYv+ffCWtMrBh8vFHoQ7rxD6cr5DpxLz/5GB8UrgeW
P6cChUNgf1EMucV5rCW+7H/n/JJ2nl4JdfqxcpTRFVUEvwoznTFmTVq1cJzWalZNqIsnTlCwma3z
gEJbaz68KhDV4Xbf7POICtOH9znZhjjTa7VCLBQbh8j0AmZJ1Qa10XFIjGMKA+FKNBMw7OTQdzMg
Us0p7ZtBBh0+iSdMsv9CiD0Ln6Zh2W9fF9koACxK09Xy+f37v8p9HATjK1T0qIDtXVKXZZiQWKq7
G/4Q3HD2Ffe8Vuu2eMglGpNyUsmzRnmlR0A2DDZaHvZyPiy0M2Mi1xFHtCKiJXJ1O9yHFul1ozlU
xcHyvdcaY0IjargCb5CA8XCVWEPJmPGID3Cmrl+VyyMdj16FFkn+4Nte9VN9j+ktC7WZz/jTpNoL
vgKeQTtLc/8W+cPqXhQ8LaBwHi1eXtlaDBgU/xpUANGaFaxGIE4ppaj5oor/ZUc0nnHTe3dlsyf0
clCaav/ZkET1XDBKlPz/1heES3zL3jdOZRBJDL6sjmWYkJxMzpaIIVLFT9Tvcq/RowTsjxMdoduZ
uNnDnl9sHcB7T3pfqlAC/2/G/R3B0Kf8tcgStw9D10kQGGHs2PesYfbi8B+bdSfD/Rg/j+uzzNYu
mD2nmsrn9BjQCw4C3QMCWAuJNIVxHMfIkUBQkH7rh5GJsxPO3MbMH90yE/sptE5sTQuQ4xmmGfC/
T1bxJt4z+pFimdFj64pLMYzq3dRNkrrdfFGupJEGMzRhdJQk73yt8RptxnnGhBHLkbtJSQ2DXu6v
mfdzeJatSTC8HyFv5kGaXOhRimR34xFU+LndWHgLVU+92vjT8UVv704fYD7IxsTpTo+/Amit/Gts
f8d9020940AubUkAqFne7DY5fuWKJzdGxLDQcijNrgaAFYztcZC2uVvXPvzPorCgac3TBp2qfIUq
bf4xmgFroL8jSLOosgdr837C15yXZaj/wVIEhIzNSaUopBaPDyb2IhSxyfMeHttcjJGbMJxArgfH
r9dIRq42M14OjdDxZ5JsA4SvdGMBqitGKnrdoqxEZbkBRZ8vAD6huXcwu0uJ+vAljsn1IIr8nmLp
IHLyB8Rlgp0pM5B2XtVEmRTwcZZkYn+l0lVUfvZYRuHaoXRrU2PqSUJmjQY1OKSqfhKmdEWRQjYW
r14H9SBl5rTKodpCM0MjPhlezeNSUOpSdQuDbffmfCr6NGv+EzCJjAupjfJCJljIqlUPTj5m1y0N
pN6oY2DB2vyRUooW/vYOU6f6oG98MHo8IMiaXQpsyDDUvWc/l4horG3cpsvcwQEe8qyQfYDBchpy
CO9OfRS34+IDWSc1/4+hJS6HqJpd4cNqb4BJyWf7hhCC+9tryml1s2D/8ZCNnvVooT1J5PHQevJh
F3pGCDjSH4+Adzud1/RycopgFc0wyzZC6P8A1sBbBj/pLfF0L9vxbe9rFsMZkOQMZDoK3w7EVTyN
+QRiNScL8WN9tyHE06IJ0FH1cVN76D+5ebcHOLwVCHcFzUcenLQxMDG6VOjMAPfeU05FZJL7uY+F
ZWbwvnoYRV6kZ3FncXDQ6sOp72HhhW5NVkusV++QgCPWhB0NlcBpndgeov92Zu5V5mYuflWaD3RN
api+vND3FTK5Fub+geHSoxwYlfNsgqpxnOHiH5IJoOJxhb7x84j1aJsDz2o5kWz9yX/ObFyq1aPv
4HVXPeVUc0fN62qpnIbenHcUOmedbD7jVIQQ1NrKniyrXpJWLVmQ+nQV0y3dkPA3h4XXNAd3AX0F
s5NFbnufZ1zZafrXGeK8rJxNjaFIVEAFSFX5gHWQ+KpblacW+PzL0Idl+VUiiRVpAJ3S5ClaGjMf
CDZzBNbpYwMKTuhf1CHG/qZnuLAUfPz6gSdy/bfIVaShWuCZ15M6OfXiKr0UvHxzOUbAbg3Eghrk
nAi+5F7PyQPi/5NcoTRvwsQ7NyUG7FlxIMW2FjBD3ib36Y/EAEvRKDlRh5uxxvjblccWnumPC8Nv
5reAoNN7jVKlWsn1CtAOzdUSHE5/yddXfp5FsuWsoUW2hxKHcbWroHW6obfQn/IN+ZkQrIqRNQwZ
a+0ReZcpjAznKkelFhFFyuoJqk5ymz3L31z5DRTmD55v573Y1rs1GLR+0yTGK/qB9l+u9VKt5mrF
mNN4xbqVjvRQ43wE384xldAd3x9YrwhE27v1qSpaZBXKdad5mtro5lx/yXnpgRRVPzIug8gegHiQ
cOBrcLa77l38ME34VXvJwKI++Itf3aKgJlibnA3k7mt7zAwr6xo3RhAW20UgEg3jLXtScv4rIAfT
zElwNbkNqXJgUe3fgG2k/yaIJvgSh7EcncKIpWtrF2oGLBLUsppkzBqT22ZK6xUQ9DQb2fwENWe1
8dHqd+rawMlTc/5Hb0DgqOA2dUzgudZyw60YoKCuPxt818Bfc2tqWZhyTHMnB+DODru4F5+AYHGr
aXAUWSeqDfhu48NoTH3qmUu8rr/YN5afGJArLiOAzPXOcL/fg3hO+L1aSCXsUnz65NGZO/u/i6TQ
eMF00YUgDHLtcmhrAI99KKea4qja4LeAdCrzgssclE4HtW2vmRVknMynbZsCKqsYBR74tJh+kLrc
3bVUEpcXGstdC96H8+YFaDw/U/Y4hnuNO7Yoi9UmETymm918cGNajG9wVE3MmhbOWcj+QCZm5EpD
S8oYtXBFencnH9IRfa4i46n5MW+WplJWA5DQwzqtt/84+5AlOJLUx+EiRkw0yPFE0NbVtubITp9f
K8yysCAHAoBqFxX2KTIDKDConQsq3EbeywHqXSEsdThEl4e7qcJQVmen7eAWrlLmJrAyH3TCKhx+
dsHA5x7c+urL+6qb1GTmLs1e4lOvNCdJZzXCEeDZYckC+Ab/5T3GBmyVY50znYCjRL3oYZG23fM1
PJXTfEzLr5aQFKiH8w6X5+nsuH5yAabwlexX2IBsq+0T2yHouk2zsWc3OSzk07RbTDxceFCFLnzv
p9tQvAAH6Z9nal0M92tyGJbFq4QIKMi5xVVBX44ezh2xsLodZH4OLOlY93fZrItlY4yGMTB10Wb7
nNTAlrPyPLLlooT4SVG/TvniID1XoH7sDkNFPo3pqCUPiXPBlq4je4QFfa30/fJrYi66sJm6kpsj
ztsudaRs+6RHzcrEiAP63FbkdgffXBm1HlxgtUzJeQsLkq0ynNvy+y79+tCC0/nY/XaT9bjvDHuJ
fXPQ+F6RuxZ2/f94xF8bNk6MQHCol1HGY/SQWAdb9JAywUTOqyBSkX+E+AWIDvXTmhUw6cb55nE5
QnY4ZrTOgADTUmcC/2mm6P/9C4jjphZVsYMmXlFQHgdEvH0ImNCgwz7Q2NmNlcw/jaLnpFdjr29J
l8eQ9Usz4uW4mQZ+/N5Gap8iUAWq7APzmynmpq1ObnfjoKRkCqyp4HtI880jx4lZSbT+/3hzp94I
R7MTIQYMzM60Q0joelhbZBZSMweGtqsp+s8wn3MNlZNcFPVYdNilk6VELfmNobhPxXdEtOHC7fHK
41cO/XAI+PJ2p2GB/g0wDF0lgPf/3NNy3b/40HS75tpIMOLwXOp00W9XRjsu0z8TJeNNM5uYleUW
nD+PwtZtppNgEJvJ9XQ0RepTD9vV5m3QoOUblqtLpnE2US2Jelrbpdm/DXvn35d0g5GgSUqIWlOM
VbW8qnCbVwIKB6Cn0aEWKA4uqApK28MpctUZWaN0+ImEJ1FAgbDUYQQIUxKxzFq+fVavzl1/bzh0
lWPip+yg+wr9Z39VSJaG50m03vM5gJJD0QQtyIJyNJCH7pu6P4Yhp/bLAEPL44tiI/QyZreL02xe
yFmG0UvBiD+qW2UAO3J4wfmWAyoU+AGmlab6b66pOa9zTn7GlPaVtWbQAdvh3OnJHTVgOr/mdUPP
9G2lXuZ3nH9632bYkoR2REApVgVFgh1azd4pWucQGMmhG3/4dqhtGf4MdHba+mSdogeKVwwBG378
wO3TQzC0qk1CmdZOomBDA5V7L0QhGGC37WhCwO4e7aNcyT2bogJORUoZysBN4yj/k9OFqQSOgaeS
LCs5q8g89hBezxXDBA4Sc4PwNHfwutxFPBKFUrUHl/p5l20MRMEm5LLo3DOsTWng9aHQykiX3Z+t
toyMh0tU421NmyHhqYcTeAqz6RZnytGWEcKFssjBOeN+AanHYiw+ei1i9qyx76CJRJqC5VA1HhDf
xiQt4N+/B0nffC/FvwE0SSZ/4w9HpHAqmq8gblJWZ1spg8mWnGyo8x/xSYRESsj3uCgTmh1mMlOf
y4x4iuIaKiRCedhUNE2+SMFABurlJSpYR8Ajk1PP+ucWf8uQVKpOGumFTWPXPKIQtNzIL8Wl/sxI
NzdDu6GBd2lYdu+Z+0LVRIF7EUYTx0+R36adVNb96KKsfEWGzRqMPZ6uJXYasXOlrYCVCfLn+8dX
TEPU7JGJQQcP725SP2djyYnzQ2OmD26xf9bAhUAIcHe4mc86gdrZhFEYatqzhHWWo0iSE+al6gRp
3pv9zHKe+0HX0lnxV0K1+aYz+CQolJQsuObLhE8DThatLV4kKAERelLHn/2IHSHXLilQq+h+k95Q
joj+DmLPPF0R1wSUW1ip1XShtClWjYe32bOgiEO3FyUefz9qH5Qk/dKHQVYkqddqEEY70zFGulxv
gEegXT92s7ls8B74/UO1eBQdsDuqcyjr59XkPzhlGYKBe0TbdkUC0Pp9rKZty7EqeErqeT0X00Ko
F7Y3YSnhAzV59oQDTLhFrM6EdIksZEvxb5LoqEjH9jitYlc2Mk0fGxgcM7wZP08yoTSGtQyGwoWM
3AB7qMLkF4Xh1eExkjoYIPgD3By/kyK/fB9UJRoMBZVRJLVANhYS9gTa1sMBhN3bXPnGCmeLH13r
Wqzw5HHc8IF719D4MEF2VJ5qtgox+29AGHbV6RBB1F+tEzODnG8zGjc3od0Lw+vnIvMZ6qjDJYmt
ItZV3FAkn4IlsbQTIzJc6f4P1JxQ+07RvrgXs8NqiGE1HuFjjEf45AuPlqQKEU/hgpp5hHCCYRhf
utafaEVyMNsG06uRzrItzUtM1Fjk9OpQVk9R84fCBUMnFvZtD7qJdiwiwBZGT4bIsMsfBbe4+I1M
OQgTELe4l9dnwl8VOz5/WpUs0L9iq8v8yiRjlDXT0oq+4C+EJ3kye3VhlX/XpGu4bQjU2KJXTUgn
F/kRUMrcF3NzrhRzwrwO33auX7apWXaLfU1iCmzydSFXnyQKgiateWG0jUtBfQ/gzym7cmwG2Jde
mr2/h3YdLHRQBDOswA/Anz3HnKO6apxjbx3zlC8+HgPsRCOMZ9DIHNvGuRPHv5VxBugj+yaDGT7t
g9wvQUkp8YVAquACjjFGy4Ao2UQyGcfMqWln9yKEzrsRlqtYcpShCVpZp2ahSR9vVekD7ZSJ8JEY
sABbDPVkyahdHmcr1IRqJu6WLQ5A8nUmY8mu6WJJWMiloSa3KOmLp9wiFLtz6v+8U534dSMjPRt0
EqdXyrJjpwymh4b28FNBumJD69usF3rZjivNVhNRqgBys9NtKbGA+4oQBRRiZF2t/XKxDRKOqQTn
kFk2rEaWU79IxYK3sp2nWX8SUSRRrl+gsgpebFhG6gwC8zFy37vc9Ime1p+Ru84gjkAyFE+033do
RED6L7lpnCWXMGSKe30Gc1+pX7RhRK0CVBNOfN3naqm8v8u6eABioDt0dMHhdJUMZWwIQ/A2L+Lo
yPlzo6gtx72S8ByDgFvMC7qS80tppVWig8mIjTh0I3aWLsIGvGSz1ECfniDg61gQ8K8TnJeKaA9N
9ebYGak2QmMkwau2SQ4hQGZoi+xc16Ohj4Gq5Mq8Q8ZogdlAaZKtUUwaJOpjI3bod1JxDs7IKAik
brYDDtrxzaLsg4KH4+PK8ojKIIqFBrbcY1Do4j1q9uZjuJnNPk/jlSpodzmBiJopWBnZFeaFauiT
loaSvR2Mw1xtfOcHIruy/eB9d67+D3wh33Xexv0K3WidXLorXyreD2gktNShaHs0z8tu2Ps5nPR1
FSarhd6AEQq+VvKtoI1Sz2BUYJvfla2tSRsCYfialpZC2kbWNs9//ZGje4Ea4FapS455rawIdiuj
hLraC4XyUJP+0YWzuxvxI3pW/PlDga3gV91rR8MLmJUVreFabS5dyWL1/MfFNK+Xa7W3OD3qmIAH
6XKgsXoJ56Au+oaNPpEYih+EduMiClTJ7y6ABS6jd3zkbTydMKe3agcQxRhlwC91pdD5P3BQ5Tc4
z3Dh5e2oLKAT3eCS3lO/Y3Fh42cn6LvtWmcLu+xqMTugGZPEm/Rm4USRGJtl2lFfhbwDrZYIBFC1
9lEElTx32Wfkwaide8mKi3KFCVdZgSquXYQfEZeeVa5PP1dON2SGxs/ajRBOS/CZk78ZpN0ZuOHg
5d5gef6HYrbeHJkbyMx00UGns1RefqwdM8C9pWEqrJF+SRnrNCPMP1WBykPPtJT1CH4biDI/F6Du
Dk6pGN2XPm0RDIAKg1Y8bLH8mZQuoJ1hs3zXhr2uVE/2M94nLNMJ4D+cVoW7eKMrzUViyEk0R7i+
uVIwcOLMBfQIbAo8MpoJNxYzS8QPFSAK+E0AcWr8cugoisK3GIMZofuudWeJIRt/Zy7qTZBBTBb2
3qj1gHBLq5oDLr8AyVgAFHsWNWu9EOzxffPpRB8mv0/cFipSlbJT3QNohsfGNq3D03I3Pv2bRZQV
GBv1bum+DpmF0vA+JAfHAjA8xhbm0itYFPUjAPSh+vDtg0865jxo4GAX0UBWZiLZ8AUA0vI3ZUrQ
uRHc0kQtjtkRY6KT7Ns8UontjijYIPWyLsacjJKNStbyqCapTL/rpVQII7/98sc9g2raImGjxCsj
rQpOYhmYHv/IKPVzPeafTeHTVdum2zWMeGh2mfrOrMOGUxh3hDWJJgiTZ1yzElOS0xJ3XGIowD6w
q66oxEBQyGeeYM2AfCmtbE/dM6dH2oTLEdA7Zgza3dgQznugWomniek5s3PVeAltWbUwLGiMfdui
B1LuyQPpmhF7gk5NFurewgRJS4KacpRk09sZTdPxoKv1hYlY3wkHsacGAnqtfFTSJ14NHfKOChuz
8hS+oGgBkzg1F+a3HsOYh62QWdQDW+mxkU5PwBBJxWDCPM2VAwHQaXk1GmXPJSl/7pxsOfDB2Psq
OSj7h8BhEknMiU6ypNumkEEarFPsZfKb2Q7oFWZKqwWq+8YH1prgtjQkPJRZ8UzgEJwvJ09ADVKI
pmLc+kEJ8I3nHvhKdF5oxZ/1qZ6EfRAwiDfAGJIFg4bztHUGLYse6/Tz9I/kuPC3218kfoPW3T+G
iLNDulJflFGolzyZRf7NMllVrDTt1HQdsw9u5l8YWF+4oHUpUDlNOzOdrsKFmO4wFOZXVkomOGk7
K+J+nAo9KOzMiFn//wNzPCmvrwxxa9cr0AiEnqMYqnAEPhVzQ2GZm/5lwH/7FgId0mZI8XFK4DWJ
FM56iEtltvjbifIjpzerQj+1nKSVzKtARZV31gRMo5aeUK5ca8ZH69qsD3IFO+N6cJn3tGFFuVnl
aiYnSAYdLetnld6I60aS5dDc9BpVqehebvF3qaxqMFG6vNUG8BeYxmmB/wNtgjWmvlahvOzux3Uh
QIOsTE9B+DZfThKZK/1LDsma/W7YGUC6gApl0y11q4Hz0JzSIoLwiu1XUpbo0AQfLP+ApRxPksCm
e/xf68co/wWWIgOYlu+QHy1oPMOQwa7HO3+rfdRKXdNyBy+ux7m2BT4or6AHQBPZYMDDXqv+bvUc
jnmIgJBheUd52FUWSVfPThMfARoV1DOwPmNgQQQJz3ZswcGh6ihXD6Txqw325zz+xD4VWm3Y5TFy
lReybidjn9K14ZjnD9M7BkpJlv7Fp180GlepObrQRdZlfUpe3tOLVDLHHhkEwdD9dHKftIP0Df9R
Y1NYnVhBxUW1f58ZyWRM/Fg4+fJzOkpFEtAzE+2zt5G/wFyJxs/kaM7nNpWHZgwM0xTFMqtf8PuD
piGUYUw7+fPXL1Z9aBa/a7PU38GQuoQyx0/4/4kJMqAzFAQcVjdLOFHIkoOTdXnx9GAOmgz7QMD7
aGLMntN9leYuDOumpeLWJ6v5DVODU/IHuVlQxpXc4asmJ6R7qAgg+O0gua2X6hAD8yrtWT6aK7+L
glYrjyyYM5c90EPQOna5ci5DqJneDW1DRjghtey6hgQVpKwwI9/+2KgxFL4VvBloX4b5eeLM+sp6
75Cir7g3WvgmteAmWmAEw9DtPBtWETGmHecOeRe889c94uG/5ufAm9JBL/twhh2OUB3CLCF2Clhk
ff0qK8TxF1Cv73bfy2sxJ3PnXQun9VdGdaFFB6g6YDgp4kVxWCwUnxC2IUklLWot+NWbzmh1F34B
a+8UJYPzvdd9J4mWxPloIJBXp3as0w95SrxJBt8LmvwTaz/ySc13DFG/NqHKKOgs9t4ZAC8dA0fc
ZeGOf+BuWQc40tl2Ad/jkg8BEe0ncHY8e/FyIjPnnFpnWJSrSESfKs7l7Av34w9WL14uvXzzEc+k
GIaXtIVZd7e4m/aMVVLIrejCFq0unXladjhnFXZq8RU6GZOyrk1xoh2FQDIMHptr88dbE9TmxMru
z6sKQSkk+CeaviFKW8lbaf1DsUUFFdyclP1tf1QyyzD46jsZI4S4C1RbkVZKmzed3dDyD+Exyuag
ZYd3TC3/zVySLEPcMRJKMJPFkIuahwkZm0hQih/DESps0Zn8QspuHT8xB9pXnCKjuXN3Pam9w2w2
nE5LV+8EGDqMdr7Bme2SR2PqT4TikbK/kjyctJ/MXK4ZY0Frc0Su5nfBdPZSKKNV8U82D+iCcgX3
eBRQnqmqfwDvT7/UwUkq6XbH3bsRjunZEYebayOci22I94av2BW0t+GyUMKirIM+tC9MELguSudT
4wf2daWts7xZMnLl9i3vulawSaDFeEs88YeCOIWqllrXIqeUqQqWwS4lqC7M/jDlnwz46o03nHes
neP21e4oZ0odMugLkg+8ad+HWnDeeKAS2CdNSGx9pKlGfJ/HOvPTNwSxgnEOQyPKn1D/KD47aRiO
MatFYIJ/kUBuIMjuYftjHUBvZWo+5qkQ+1UnedX+eqxNZfw2eEQfSjLLRy+ur68/mXrY6zsiGRpx
0GMmMdf9zfQULblasaFHraLuOZXPhPWZ0UYfFJyn8b8yTDfRSeEwoOGhQVIO8ynhigVJL8HZAbwn
47RKvEREZ00y3/qm+/hnfaa32yLWM9tQeb/n0Vi9oCSiDKa4ZiGMVumjjfRRccXZ0vEDNS0d5sjB
VURI53OOgqCwlMaq11ba4Sb5bTv85dDsDwUOx/ORSs7Mp6huvB6XyPT7xbxJRUB7iKDA01eIujSg
l7Pf470sUJQM7PNQfqI6BKQ9kJbu7oPekKMEfbFJGhB96I4BpRE/Qp/BuFni5FoHxr8c7iHvEoBn
a7YyMGWlft0KYnnD/MvDCf2I4eX+NZ9QHd2ToO/2Ue6VnqlJ2FYydZmt/dBOiUpwTmLThNtveS4/
B2dfTnT73EPB4aqBoTrv3vBVFcaGPay+R2fT5RX1HXyg41DgYEHcyGRbWeTBtRtRthG/HU1c+1w8
gaVf/p6r2085xWjdEJ8ieawmPrgiQZtIP3nJCfVJSGhi9CsdkwHWPJHPXoZfRqtkplR6Bysix2Kz
2772VFbTU3XDOSKUrhJ/pJSUfrs542pfPtbOa9C5+zDbgVRs3P4bCBcoKI3w2AGzKSna+wifrklb
1s0EicvHIXCMCRinQgd+9rTd88XGKnRZwYNitpeMFDGGAYgV6QrBvdtCKxJuCphAw4bWU4ADY0Sj
IckZRdd/n4ytTMXa6AU2fvk1F8mb/uusu/nasoZHBw7oGbmKff2JXhTRjN/Ydvhu7IvB12Nexlzh
/h7pSAjC2OgWILtsGU36b6Y9i1+Tml8xQECBHuc4Td+oym2pNlA16AbLki5SNwDu9yKNsWFWvduB
BFs5qtbPCBzB/ZQab2wfbc3xlntYpJff6JGF2RuWyxECUw2FeMwGVOPKiRmFYtswplpbJOrFfzt7
Cc5IztK/KkYgA1KnB7uw6U92MgJevfmVslLqvmZ/43Lozj2okD6OjQJ5CfGxW5eqULlJRn1xc9z9
B7DxPbYVcNcBqxzYDGQ/J8kDCkXPnw2rU++CDFHZFZtAQFcG8CgXS/K/lirXVMrbI1K5n/+FSfNc
f4kSd8/FuziG69ng7z8TLnx1ZJwCaBC2ngCKvuSc5zO9e+F8UAt2vAKAJ+RO5D9b2nsCHcHmy9IR
FUJQBtNsG0Wxtvg0n+cfsOGDAby+6ziNzKK9XHHKuQst6bIz2X5cIGbpYDI24F7LQcbpjE8wf9eM
yBYoazH3CLp89yjfTVA7CjY78om1q4hTFd3FQy9t/I1i37qATXqpwaGj6XX62C1OiilYpQk/eZJA
MqkbwKCzbCNuy8KQJ2OO/fxCG9QwXK4/1bAgx5fdF+PZChy9csiVSvBaE0tgZIog9uAkR7TWtm4f
ozVK4NkjfuGcnVM64mycqZtso2eLlbCSqX1pLehW7QrdM7IuP9fay+I4tR1/GPRY2Ndi1PPqmURc
vpwAlNJKH4MN3UDM85zOVKPVAzsr3ZULCsgrmGs/rgNUEFAIPNYOFNMitmEm+icyz4HgvSpYWiXE
vYjsvTJdxSs5lFq5xPKkHoG+xTacGswHutkuJtq49uoZ4G5XYLOzHtZz7PfCDjxgH5isPjrhiOVq
8y7Df1kjvc4LYhxMnet/BeRXjv88Pq5SdvD779s3CRr5/M/asLvCXll0YuGs6lEwiTu9CLt5vz2g
Ad5D/gRPk9T847Iku8mz0LgpsbNlhrLCKcVrS3UziJ4bG+T7jdd6AX5eB9kL8UV0zMGf9z/1U1wB
UOBssEz+jM66dW2/I7UB51bmDF1LgM055n1pPUqNnSbJI/lX5OB+jR/JiyUe087zOb13DgH6IGn4
a6lxdVrIAhoUypx9rGp1s0PxqvpW/Y8H344oFd37/BbMyYBqx7qYYHXSh6Z7Qr6phLrQAkLfzHJE
8gOzHggKKneerlc3Q3rQASqJPY9zIr/lAvmE+DTVqMgfpK06rYHbv0NVz2ycZ34G31nSrWsd+2c2
tdY668HNbf5nd2avL2xUuC4uSEC3gwmqBSTt2QvlIly8uBs85i/4M/WdzgmyiqkgGBPZAPFUUfwv
AjN5o/N/ZXvcaO5/qOBTymKrfw6i+1gc5o0Khi0gbghDAOGzNge5onWMNkt4eeXTPoCdEgDshUDx
MPyRSKagkHvtO0shcton25wnimEktbBCE4K2kF4fv26x/Fc0nfvv4th84tZz626HsdsJNn6Rbk2U
P1/aPenfEBOCCfCefTVl0zVXSV7k7f8q4CNPS9cWxweQIVh5zh8K173PZT5LdJ4DbuZneS/G6qX3
C5yFM77Urwagk8YkFZjkoLE5RDJnlKI3Kw5WCjs3Cj2zoJxRdJD3AL+CWIH3+yrqNfpt1SpQODfL
4t+9EHlTlgik7+ZpGVShoUu4gxbZLgEMCsqESsmqUP1SrWqFEGWxi9MT5l0P7nnASXivJ5sWbKVn
W/ns9D+anw98L3GVHLSztSf4LVFd6cuGc8cTgP5+HOpDLd2IRoZR/kB6ihJO4rAesmhqDWMZ1Jfs
H/Z4lrFj9KxkOBoVJsqS7eVddpmXwaUT7xT0HGc6FNvzd8TDXoa4YYdVmlbP88yw+IMKBtETYASO
bibPsL83LaZ06ApBKDSx33BGWuxEnNXr2AdnaB5udn4gaSlwPD7Av5ncpoZD06afkZA+VC0sIBoj
2CGLRLa3+zwPiLIzzgr20h1P39B1soZ7rna33NRF/PgonWQJ+s1Ks7DIvGyX2+4AZU4oPhd0jm5I
noCi4HN+2lI3a+pRQPVyqlv2x7XruYPwtOgVgtuiTRQy/6Czwu3V9HU5HDmSymVV6Wa9kHZp+dk2
r61W/xAj+sfg3UXqdEWi1VWafxx/S3eURzGjYVgCBCFe83aglPtA0YSHX83jUxnJMzh/XIsVxG35
V2TY3AbYGkbflLyEiWxoHxvf/aoNHUg1wj/tlANyt1a4FcVt17dBVqlacCc/I17PHyeA++e7XKwZ
dXZ8roCeGzRMjZsXGex8nZ0ZvTC4fMHfnXCC9plbrWnz2Dtl3u0Kky6+z76g/azVXRZ8dpNrUWAx
63dvi5KmiN2uUS6kyFjtBzHbNvKxgpUHxewGUWfXiv8huyWfjMAT6YSdnvLTbG9/S2dSGi9rd04B
gHIORD8KZv200GewCF0W0uci700XjD8jGR4pSIJfyR4u+P5WZz6VhUS/EWU6W6ZAJJ7J7EJjSgUO
HshVZ8SAX2idm/3RHiFsJT6AqmME7TyXZysAWxiwrwamqv56NddYPziOWzYa0mmG4FaI3Ec3Adz+
OI27wlq4oSNA0qjv2jKxAtPE0bhnlYaukPPX2ed2m3p1KJaBBRm6pknuAGrfk6gZgTMVa1q446+4
DIkS7xxitggZYXQEgwyka/mSL7LhdCWrcJs0D4kRgxSHA8kuwAOdn3w5vaCU92wpPHnTMAvEG06q
sHV2+mKf4A731dWv3uzD5wvnNJsSPOam5I6JFXNsMyBAEa9GBCfkqirB8i36/MlI2zFK8/l+Yfsi
cE7n3jt96i/1womMPE3jejGYRD7eQofoe40jndHGWqpBnnKiCOuS4+wEpJLoylQBAkDv51bl6/HU
HTp4aiLmK68pkp1PxqMt/UgWewDdanzB8QWiQb7wJFq+JeQTVU1rVr19ooAEf0KYltEuJGbEwO9E
2ITrHRnFLGxl5hpkMc2tZdlyS02Tj+Ujp+7cSd8sljQq5uRgViv9aBRkbqEQ5ACrxong5IZJ7tai
hUib8FE7AIH480njqnh58fOCvn22UzyURPMor2Y5xTCBaXpPiT3tamrSPhJxWTA30wHbaPJatjR2
QDwnl982X0juWuaAuyGAUZVkEdYgQLCJ555sko0rgb4tTRMR1fZPzxwRksb3hSIf9aGZrGnnv5Xq
yxg6sQ2u3lnWVMl9Y83AyYp5BRter7qD63uaiEe+GK/gh2xp1sK9Kxoqd8j7B6yMLhc90EmlhBym
Ze5trN1Y7ejyWAw+E8PgQKJuiVUKNSWAaQEOK0m2qHePuEFWAp0x/TxiC9oVGGkdsdJwxmRdRh+F
9xU5pBD1PV1IsTTxHnL9yphQ6cd4//xk4B1MvH4jf9xgNnHs6S42LEnsGCESzHRYpty+mAkQecUH
xcKPAabpkRj+sMFjBkByZN08G9SaQVpud/OyzrtXf3Jqz1CntqxDfJ349dzCubxKIOqLwMPzueyu
FcSF11/pXZ2emuF/A7wI+W6eBVvvw6MUTUfkMZIrAU3aSfKcRFor4Y+rrFs11Y4h/4mp5JwfmkTC
Vzy52Z2rLX9728VRb3M2XGyekX+pcx5RwuHtcqe1rgUwReDHz/fs+4vWhVoYkTS5DOOnEMmfF5U3
oOiC1Vr9gjsR6jVzSKs8fOANmXkWQA5LusH0hWVipi6fUTK8ZJkTDmjlgCqGNs8BN+VwYeYng0+w
LWKHE4CBDlw+AFlbk0ZAoyOOdWrf7Y2/ESc3RETLdLaHh5OZ9MNLu2pDUOsCqMgzbGN6Y5PxYnUZ
1KmcI8ZZGuZssH/lygctJCRBIESLNivBuAPuA0yTsyjcbcXK8NaiyZs51/5T2LpdUFTWjNjPXZpj
0URdiRikm30grnn9NWiwLZ3aqulD8JSxV9+V1OpT9b76/A9GZxJT2835G7kLehWdCMEAlJS2ogk/
rgx4BsYyjqf+vY+Az+YXwLFoZRsQuvW5LLo5FSz38nu2JTT7HljmoqfVRAEbYg20nsD+fSvDBgz7
NoHo3D5tCeA1EIwXrGlYpztfsPdi0Zr6+0A1zJksJrD4a9miGd6DHNgv022SM4h9K1BAjcjY8YcT
z8LgzU5YQB57A41tOC3XhzG6OkqGMiylypmGjBjl9OrrUD9+jSugzW1/tHKOjZJk63TOfMkCaUrc
PdkLjIddu0dQBPPP4OpmqDB90zBj3MOxqPSgy1Dyv6Ad6Kk02mIxJDataO9nU/HNmssM41qyuk/K
5Sxdjc1o/CQ+KKWvqHbQrRbuu9G8BagRTTq6fcdECwgTQwx7gHtv7jyzEw/kvoceW9CR8Hqbs9tf
RYrjNsENhxN2zhFIla2UvLk1wKMbfWJvJ/qzSZAqz+ULJaGlzfmXfxD1Yk+ztqcvlWyZ5cbEHI1q
NF1GX++VBvzbF60Ukzi10fNto43AdEGhUJcJnl8AvCJQdTuds5LOfDDv3Hjs2ACS47EnSAEBPKff
u3vnhCibwnn0dV6umZLJYXqnemioWZ3WOXCOITlijXyh7DiliJkch2oxl7ej9+x/0VaiWY9LHk9g
mut+Q1CkwawR2ByejcYYs3qXujrh5fJI+4KMba+FD8CrVH9GToUWMwPhqYA+wIIJE6I68HZxE3PW
fN9k6T3r+cx7IvmZB31tcHt+RuBAPqX5ZHzIdzjuNbv+yDoCXWu+Un3W8YbsmqVcVo0wd0GNwd7H
aIshL82Mxmn0KY51Q+RHqUxK9PCLIOPL/WHhgvl4U7ssQeYuzC7n03nzu0Pl6MlZnva5eUAAOBSm
kb18gZxoNXWy/c0Z6pPSPmBUTSTr2+XVzRMx6ZL81vDY97oSwwQMsRyuQ9SI6J7/Qb6dHzpQ12S+
RqcUavX4FwJU4WSaPk15El2j+nyxhTL7NrPfXzGsVRAvXE0lNZxD9LrEF7o5caw/oTF4yZt9M4np
65FlQAOqI0yjZxFcYj4iIzhc6u01s/j0n0DcdpAEwolJz4Q/SNraEAS7YNduRKH3ZFuATYcL4KL5
OR6SscJ46/mmlB9zfAb6Qr7DN/Hlbdq4NjA5/GCzeFFtVSe4EHFsYH1gCWKq26o0KvcKVUcCMCGq
cHifD4IZtDbHmUxfg5Nd889yE6NW4b7ey61a8O4K1el9uznk8dXOK49MzeCSyU6tNA8am1VqZHJf
NjCRh8FmyKbcqx3mLerXtb02JIdB6xHLp9p0THHhBwGlk58hvjyLm2fPsqp4AS7I+OtceCMHMrwC
9gIKXgL98nvbn8L4uJetT6sMl5srDd6zch+pKSXqUQIPFb0PgybVIpWh9QZs/CquHplvGjAtcfq7
61NhycrKKjt0ylhriQpTIB8s4R3MTcpVSV9GcKY32HXxvkuWI0oxH3iqO+CICHQcdq0ACU08fbf7
1ALyeOgm7glb+U8x3GB045LG1tlTuATbRi6hw64zvbAt8Yxbp+crYFWYlf5I2DtfdJNpxV50BTbv
Qen46ri5evSga34h6y0fnr4BlbI4b+88gUfzOxrR/cmDSK7V5741452o0KngUtlRCibDFVf9m1OH
vCm3QIKRaigDv2mwiszu+687MjrBVXG2ZB+6BDCwzUmeeYPAU+PlOBSmgnX/OzGri3AsURG2Qs5s
U1VAUO2CK3/uvD1NjXkbkeaxRvgvnLiNp6yyOfPwhMwUjEWTOf34ofEc9VpwKGC4rACdySm4QKA8
4zEAlzDlsvVxu+hT3CDw6cRuo8oaO+Cdx7vaRnvaACQGAZk9FMrciPWJzdqWrfJKo5JHo2GevaTt
0sbdLyxVoQ8Ij62ChcoUJLWt/Bce5XYWA8HDXk9oYceZaggSS9fCpOpYOqe0CjYuKcGvBA/PXpEj
m6Ua0+SSMV5A4+lbaV+tjnuIvzs4jri1qCj6s9Cp3q8haYhImVqpPfXVAX6C0OAagC7iJs8xiTwA
zWoTSv7iqkE5gg5Fl5ULOb2MWV7joByTYlS6dI5nawS7Ld5RsQq7o/zHQ+HmzL3xuOx+P0vw8ls1
Aswvof5XTcxtBR1v+jguAXBh9hPO5T4ac+Neo/MGW7jVSCJjFiwca5QnPec1e6RKdhpKo8fOCTyQ
6IK7xelWmjfsSms0ivnhCpVwLBDCfuduE71DQ9+GQR8BF8c1Qfj362Zl+QtJpdIlZI/BDtrsJKRR
r5uMvS4VzlWfPYPabvVJN8Wy0+u+7KALZgYnsa2K2ib8/jOVceQ0F1K0rE3z48w7AKDawBeG+tBH
kQBZGbZUtdag+zZORFWsxHnHUEtGuJbBA1GasHDN5P0mPnpaWT4xF/mtH8GPhAdHj1PqS5lBhIi6
eRMRwCpJYeeSFog9xAfgHc2MULvIpPd+FrikCYmumh7K1oLUIS8COsra/jstoEpFSRtNDfZGRcmj
q5O4ijB0zRQcRB7YLjn42v7/EjOlv4dzQhwHosoL16CfDrcjjqvVpFNRfl9UwCUx8WWBPuxFXQSj
Xa1F/DhhUYGoLcCxw+8GPjtK4MXgFZM2qPcEmg5ZU6g5QwTxZxcSIpSQhjZMMadG8NwOq2qlCZ/c
BLsJ5xMD1v2mDV4jkXYIpyV0lWKBTQBka5yAXMcXek5PkKUGDAwvE2NVNP7GJcoZON2A4rt0hkG2
2vv49wmHA31Z8QYwsLzgYrHie6qEDvX0BaiW9FhQvW8/goaElHW7/aO1xGFrwh/Q2pdaz9sYgb6e
PVdAptnkHpv7rbdLmKrkJEJhW2yoruuh8YauDn2hD21Rg9j4pQQ1fxv/9QllBKv59hJZm9w2rf4V
O2Wvfy0hKZ+PdAFVHoryjjKzv9RGm9Klwrdlgg8ic5Pv7F0/dMLT3WAucIgeqV9IKM/SFX5mIbRf
LUS3JhQwhFdVwS5IFkHB8zOCkzOaxp6GprP3PultsI8mshO041oSMlTVuHQsDnaWkxv/p7Wm2a1S
N0NDiJaGoX9zuTIe6DBLwusv9TbSZu5CeVF4Lhs5aJ+yMZDjuzIEf/pPdIhlKjiUtPkpee4BeEv4
veupSgkXFAJyQ/IwNV0ZRYIl7l0EU5cdObCPgOH8YG+PjumafSNSMpNesQmr2vQI8gDyjNIXHsBg
06EKPjUYFsVa8+HXLF/bTxu/iB1OnNtq8ugEnM1EMsMh0/7hQn/32JiqANRQfvnosfDV3XnXRdNf
8QLJmKay3GPptk4jj7ARCxxbdl4fZFEfVC/tuiRpPApxQKCiAFxoe1hTUWvB36QUyxuesGUmfxWD
eZElAYfytWb34fYO1eEwEZl+boybW0XK/yEycHSMFDlOsmMpBjK1pjMn1g2/1Nvlj0SOZ3GGzNAe
KXDr+Exr1iNVdsF3HJAfvTxzy+SKJi5jOAZfSMiiaZ1ktDWRIgdDqegI7AlwrApei93zSVCioUqY
Nja7XNZ9zqR+20QCLTvpNBSIk/DgtsdW3DpENepZ+zUpV0VpDWkdF2Z3QU8g/LNoruW4DqU8afgP
up9Na6/0bg3YuliQ9N/p9LMDyVMFmkssGWTSTHhhLiTu/4/SuQK0K7z70IfoHShTi9hBP9wgySE2
DOpdWL1ed4hXZgYEOG8C6SBuRumunKmb4diysqlo8WhaQavHUuy1OmH+ZsZR3RTfq1VD6N2gUkAe
PA3KMzLOtgDBlSBdgB8VEBoqpBJx6bFgjUZLQxGrENUxqB41Wf6M9Fr0uc1B/N7cNYcVbegKeQYL
jMwhFQhPXtGkhJ7x8A4vG42FarIhej8rFOOU7XVof88MEEy4DjPJLXFU9NY2V75gor3lX3gBCPkJ
FFSvLO0c/IxcP+lKiD6SbOD1v2bKcCokavagDE48NkCJOVN3+daEPGyEWaGkLoTxT5qFMBeNH0ZH
tHxf00A202P9qNLfEaWl1BWuHoVw38sr9GhhTg0ZqVbPuCb4Z4DgHbUd9ThKNFlRcVGCyj7/OIu+
qgpxlc7BPaNdbDUL75b2FaYBu+/h7tDHwRi+R0opLCa6wzpe9VP651zAQ1A8BlrpYzLm38P6yhC2
a58iDDJVT2VvN10VoASIPR3hYPDcGm78kGtdRR/ddpHfQAnTYw91IWVtVjoeeTE+g3OlbosjsZiv
ERLJ+wpWGp8Kq0pzJoK3p3m7IdGyn/bCNGfvvXBDA5yN+/vAo5oaHOoeDP6gYNlIYDhwW2iYLdQs
hBz/cz/g5wte/FHmMp+QizgHLieQVyt5CyIk0RB3nDEVWTUVwgQfPh3vpkAMiHgdGnAJYdKjbqWT
0LbZ5r/NpKl6W0ozzFxwByHjdHnFr5ogUNTUnv7ubnuvDgBLDLvcV2uUJ+QgYpHXaXn9lnAGneQN
UsY99jPSaW/8eiAMAYu6MakfiZqa6N2vzNhGwph44AhQRBX8bJFkozOYNP1QsocDjR5mcbPuMYRM
8icbyLM2d10Z+UXWUN7zKbYqsiA37C7YuZ83wGO+dH0OZmBxtv2zB4lansuovLyzJBNTKinu8b8F
+ECAa1BQ56PkY10QM532Jx8yq7AeC/cgdfGU05FjuUElie1kSCE+UXibx3YdlhtGhH6VrTAS2XWp
nGwWuKOJH8zakg/rfjbMqW943qA0ymxiP9XulWSeSUHcJC/9jbqwu8H+SzGYdBZFNcecmJs8DK9i
MyDBvYFNjJe8f4GHXtYQVeEfADn0lV7bUbg5kLlcJ9B5un0Mu4QEE1nQPBnkBwOtOyB6mkWhfcv3
dUQFSTjx43aYj2+A8803/CWrjsJYoYTyK98/6u+6f4J54bA6MxdqhPQYuo/lalppJ1w6UdXDKLh1
pPN6tUNVXM/mvjQavU250xC634p+khP6lWRTFQH6aAlqA7F0UAOLx4/lC1NgTM9z25VGhK6aEzqO
i+ozCt5cZGZgN9TzeN8B2//zuwiPCFZZqXXv1pJAVyH+qpl9cmb3saBexXoAddc8FH5yK2+ZrLwu
RDhOiThKXYXJg/mNGygY/5SQYbVn/fb4qXGmD3D6UAl3X9anGlagSrd9oxGrWYW1v3ZEFGEIHbu9
vfc9/3XYEUVqT/ju3ob5huhDx/XWAOHiqHhwQVk4oD+QfPdlERpyzt/fXZizK7KxjL3Ki9AP58EL
pOq6JIUJo72QOGHGCfJ2cnr7Q8cJISvyshS0jp9WZMIXccyChyaGoIr93HsO9gWthPUysYBa5DSz
2feO0xuT3WMAKSKiOD4nR9/FwjiMlXisB+D4R9JTOpLln8PRB3vG7MxZ6qVBpBG4NxGtPMvQmUAF
1/eRf1BEfBroYr31Rg/yCZ7FqylD3zLzrwUiz+Wx5MRf4IyLgV53uQrMWKBIyIoZUHveTcNTrK+m
QrPBp8Db0YpuTslyMym8q9Kv3aGoMOD9VkMdTT6jipv8vt32tKZz1kk1bkbCABMC/C/auoyjBfJ6
DGOHrq6LNpbYXwkVfrnMuOM6OlGPjKTSNsJNaoE1ysCyNHFS3qDnjpfj1LDMGA97hRgfR5qbxGhZ
/8YDRDy8CeQtGqveHIAYV9gwMuHtJpjg69izVCsPxyUwgxiaoOOGwVseu/5bPZXUFcMxdouUULqG
IHbyLHNx5mjfZx6l3XwKRPR/Veqrxajb8DYRqQozsSusXsaKzp4BjwVWdNyyfUhPZvY99ynDv3GN
rbOgHEtB9ogzoenACGG7db76mlhVTnwDSr4u+ZbcqkQFsKlCnDIoQqNbTMm7ICU3N4iE9kpBx571
ftWYV2906NcDdEKfIJfmIUfo1LfVLIzSVl/iCGopMW/o1QrmLEVamwgb34FIzrpUm8uUMFjYbstJ
/Mx77rbe4EJTswtFlziosBDLnCpKT5rNbj1Zn/+o5+8jg4EI3KCjSpGrPMG1NFIi80sd4j+YoBXu
vglHK0XLV6MzjaBx6DFilKl2dJsAvKFx0r/qSzftcOH5qYMT60DPTsv70O6+DFPvK6Yb5jgTGVFK
A+nuEpUqLPScG8QxUAktgezFPP0bz/CcH67qPJSMIKDq8yczBc6eZEJsILZGD6o/4vde6YJA7QXb
3J8Rhirhx047kLj8q3HVNH/g/jnKHANbehfCg2fKYUmtpQ5pdIHRHmKu609NTWEs/Hvhc2rajFj8
d9CZN3gqeGDBgFm7nvmgmL7WjZemKL+mj5XR+zJeD2fHO893DqDUT7ICpMVjowoU3uChDMG79/Kg
E3C0wRy94kHd6N7RxoOQV5GEjUCDg7BZ/l/6zz+tpm4bggt7tikFmIUaAlha6hsVRi7t5kEP8L/J
eykutoYms/sytxNujufVBb9683aXG3WMyaR0b3T5ffUfPwAffgz3rY6D9t59xvTP+jHlClrxZ51C
htn/pXUYZVZFy/tk3/4Bv3n0NohdowRiW9HV3c6uNzoRz5JEOrCKDCarcLuy3uVrKJXB598iCksx
5yhd5eyVF2sddQ9xvy2IUoCx7TK1tadNO7LBKFUNkiARkHR5AtsBzLdj2lCk2+3FGZ+/YFKJS/vX
cUgJFt/bRGPKmxESeHrHs0nIjtO6BE5/Z563q9xdl/WuegfkxQeJiy0DpaXOimtpuODPJEsiev0M
SqkQ89Hb9WJufLrzuziXDocQKe1CaYXhWIOq4PKCFRFPnB9kk1Eb3r7YTsBo2FvOKYAef/QUYlgz
0EAF7eHU6tS3/WIh0xkaWHbmL6ocF1dAhKYjpsLxBMWTX9UPh8MMyqWiX5XyqxwpujKPYD+BYHlE
dHmuJ63Z9yru09aEp86kSL+8rvSMFrsJbkwqcOxg/bK5qlPrZH14sjPMTAgrHTzYJezUfAmbj0gc
Xzmo7cav2TGxpk4kf2ONwpLpWnQsG5RwKjJbhoyOjTzwSvrvA5fHzF0hBoM8J26OaTqyRt1Glesj
xKw78ANuxa5PaFaPOAUrPDYEdzyno3oqTIr5S7oameo1BjcHImC5v+QE982tar/ehXsd7YruQ4Bn
f1CG7gr3rIdhiGZ1akHnqv5B+zM/xlHYLOads5LyFGnPyw1OJvU6zsu+eRXDrOmxctkfay8hD1XS
+RhrKJYBEHw2VsZihGYGlgM5rhEF9rppfeiRXr0zZqNVp7T2p/3I96LC6ZzJQU5O7ePxEO94joNE
OHWu8vOpMlT0Qicb6piB8Q5p9uRXaARZzb78oUxuuY5P97ksfBctAhu26mldpKXh/9gBVuOrEnTM
r1MXTucNBJZu0HuxR1pDJXetI6PH6T4HCASpCUQKKciCCYn1xGGEH522j5OHdbDGcCVh6OmB8Tm0
kY4tebWVWWeVSc0aeW8sFce/PrY43xSj6nCUJxyakYcAKpy0e03WJTkZQgpF+P1CUnTjYwlbLQaC
iz2ZZ1KoiUh5BHkkED/SMYatZDMOUJbJhAvtoamYN2P7aU92G5m70ALoHAw/cE4CAweSDLoB0h9a
Slvt+RpxiZHE26WV8v5L+96ALFAIKusPTdHcLnRnryyn2a19EPIMmr4o//v7cUGF5nlpwaeQrovO
yIOvrgg+AvuWN4kHDH5KYXqKCYfyU7oMS1dDxz6/n+x7HJe2ONiq7dLO+kB8Pfr5ToIBPC93cPKF
GGvvdXQGcJExQrTa6nQhG5Hz5dPtXWkMOK3zGVFJBnI44K3szFfKhtC2a5Ai+GSNayYXRYf9QHYM
styJ2sPDzhbl8h6PWQdKlC7lfGL1DLqzkI3epvWSoHZwyiTpS/SATR5WWKEck4ssLgMcRhw1oPdL
+IQza7VoJTPmN/pyJb51QkOt+fVvjmG5QGgqyNjPLb2UAObrJVflt51D6DGfSVKRK8TuXAM54V6g
pgf+UlPRnCrKKG/otoAZTAZQJ+cuweJGXzHNpSb5vqQmsFsvcgTFuly3qmkgUL+sjDc7tFXrjoBH
MLQvvRS7kR8lMIBqjct6ady1JK59lCKoI/oZSrR7B0i8f0vqGizWIcJSDG5rKwiF5tumwHgub8b1
aNC/4GuXiUpNsmGcVIFHrdKARtQXeaJsSqM5034dNwbUYA8EYCRMILRKXL24PznqOV3uCx52B1cd
6ISjGViMD2eeZM8lxkRYqWCeH5ZAgHxcEHLK25fr7uwQKe191TnkwS1OQQ1ZIrcxEAKlbtFX6DSi
ORAvMIv/mohqBiDfEZ9ZP8x0Q1dnQeXPXJcUX2zC5TwEmEydTToQO1MT+xy9eIkh+KjdoTzW3hui
vj57KQ7vOV04HiB+nfglRvGwa0AlUrIdCIMmBfU9QbU8Cezi8bpgaZELQQtfAvCv7V9KMDKTI5FN
ZJQ964eEN158O5eVSenWXArpe9GRJuXtqeQsZEQbTRodec+72YrcxspgnJf1JR3Zo19kInc4WbcP
65tDFEy63eno/RZuFZuR3U5yf1c0xEYQ3E59FzB7aoODdkiOdjCC+9db8r6Vl5M2b6Mlj35hmx9v
uKQUEVkD6multV54oNm9yXck5twAkZNj7mNaMrYQ9f+3v83x7CwbMV3kDubUEeEah5YqzxEzHMgT
1xwlnGQOdfpV+WLNoshRSIOEqDhcLX/nKQn/mXCeQMTU328V4y7JZJtaRTqvPS3+TXSuFi6xbzcD
l+6Yn+2A9A1ZXSPeIpJibowwLflBXl1+dXqkoHIXGt09ISJsJW6lIOiieJgdr3wcZExV/4lNc3tx
YPAGHJWIZl8nu7QQcRoyCpFSPEbb5pjbkYUb/7xtQLI/AB/2Dwf0GWpo8c+ubaoopqaBLjv+rvdy
elqztUlP2tqXWSfFqWsVBPGGFppG33nsPFlJw6Mo5IS45gnsoSzvx4uKFMoksCG5HDO/21pjnl67
58p+WnoxMn/7PigBK9POjxEE5v5fx3W/iOYqdQReyzKiETbkoqxxoO6hO/QDmgjJYF7mZqaBgLsk
A7tC6lf0gQZ6vadp1/YjXvTqoGytackz4n9r4e99ZvcNc1Q5xxoPaYrzvcicbjTuzc2pm87QV1oU
XgXVTu8fkXFxZGjQ4Va6OuNQKzxXTOEfdxuWfdxzhl3KWOUKd2ICQzyMKjut+IfbfeTc6OF8wEZv
qXMTsGlyk76uJXVMbYYgYqNf+uqaKgQtn3NT5xRlf/nosXsSYsIzqUtwCubLkpc3fw4it4gMQrZm
/AuuIXyK+McPtfHu+2Yw7X9A7T/rFDFNo5DwhAEiLzhRwHbWARxgEF6O+x7lHC1olYfmFdEH96gW
PHeTCyqehL+fJj9FXz0OGADO6R+lUueFKAqGIzXcoVV4dyRheOGxr76IawkVIMeCrfuOFklpU7jf
bqfdju3RVVhBkBhN3GQ7i/10kGAtHdcsRkVaaZYqwDRteuylrLkmyxwg0g/3aZGVylLYziN3lR7p
KRaTej1jaHvjWS3YeVb16GcWmxTuBDYWt5cwmxAuilT0nfoT/rqnRKELGn4t6IoHuO4XY2vmQKB/
ZFKMEHuuSwbXiGuDYk6/MNNIzrl0ibDJRFesj0WPCrkrjMu6EdSLWSrCMfetNMtod0vj3MXXPbkr
YFYk00mAn/+0Iw6UaesWVT/K7pNC93W4O/JQzn79xUlDCWsCLyTyl/G5AQ7r9s0rbJfHrD4rbkMB
Wa1LRpHQx+ygkyagS6HoyV7a55x5SVuiEAY531AO1uBKmKA/03mI57dzgQN1zUaGhtRe1jiqjzpe
0AKe/w8S1+P3gn/O3Nw82ln2qn+CaZ4GkD7Bg1MEnf960ZO6h3wsh0muQnEbtFzqnXZ2F/viOYKn
ndIOpTbkplb0XPE+WoY9HUpOzO8OUefCgT9d2LqaA7/GxpKiv/agQ+OEk2Bit+jwzpxu0fnOcnVZ
9RWyrkfVNK9rDncizejU01hJHZcelkvuViUK2bLnXEeg9w8c38n1RFfdfaivVxtpe7Swex+5wl1D
cDj+/nMj4XFqhb8D/raFOsV/uFTv10w+u114oKB09NZltA+8lR12kpqM2JEUPe70WznPp4A1oRjb
l5hRgJW6Xi32rwj9HRbq796xfvdHS5HyNoy904BrdT5EMDYuvBDWgt82HmjBudjlbvz8tcWARs9Y
NohSFhi5Cto/fRr/g4iNLEUmLfa6ZtPcc+76p9HLNeRi254h8bGsCNVez5ZJtvg/v/raKMkgRZfn
ENOAH4BlDx6qpX2TaoQw6TPq+EEG5BMYDQbekwHhj4Fc5z+qfTW/6vtMGkRGEvtNAtb6f3V/siVy
maHqphJUs5lst7Lh/tsIP+t5xCBjnWJLRmFwnkZmv4RgO29h2Sn4Xfcatp6QwFzN38NnHO360ke7
HPD5FY2cyOLC2JVLwTsPcA62EELkVxCQKgUmXJfnv2usBfKd+OWG646SHWRN7i56hiAJLTM21/50
ZPTTEP+mMyhd32x9OecCjMUHLyvmtcBUONkZSmovz0hm5Hx03WlwXe8dQml9K05yOdzy5dsw6Mus
Prgqio9cFsD7mmFuHa40WJsWGreZLe63qIU7nrhZ7JGUhZSgbthxZTT4ung1EbtnXdIbtjm+mfga
/unIg1eWuN+wqpt7kvN+JZ7xvy7W9Zo+mT9cQAAnIIpdI2GZdfEkWjY7Fm2+BjSoYfngWMKaFYLX
FYttFM6w8OMT8MEd9GzYsRTyRmtZLloCkAGRud5wjpno3MSLgNquSqwhV5cF4mB89VLzIa7SrqF4
0u3B9c/LvjmquwRHlsImDh73xkRK7/OozK9Veho5N6DGouYWIFbvAlCooqjEZHToHzCdiFZfrXx7
B6hI/qZb+MHxtG6bvusi7ijYhtaBtjqoePcmN8YciVW5qEtXdchuXYvhvlRxdPyEjmKUJqLX2q5f
3RkhMczgVmt1NwLbKFmDe12nGQ2oeoGP/VxN0yLqTrwYkxhuAezVFafNpFrPFOG2hUnsQrJ8/XTK
M7FBGHUtiJP7WMqeUfSSXLJLvSaUFzH9v6k6H1sw+G4vR3nl9CG0Qyjof9WmaMS7CNPbAeTdZnTO
NQJkJo0ASins3gFRGhc6HyYbolOeJkokJ7HgQHO9PSaqgpebWYvGnFJzPAxdmabGZo2+MT0ILPx3
3W8ZuprEFDtPuSUx8sHBHwnxpgDh3fDh8+KRLTHfXERfVdAMJrdH+vcH3upYJ+GxA+xFno/c5Srz
WK0T0lGV+molc7RnchLz47kUlUFnkHEznVENfeKlQqaohPVtpOhzl06Kh/QTNQE3QgweHnsKsKYJ
3Hw5i4yxdY8/V5qHFEjiz04t3C144l5eoXv38DlmlsYh8nzcNVsrMpC3sFYeQ6+SgN+ZJ/n7kIP5
9Mlfu+gxDr61f5HD4v+1rE9s60zgqYb7wp15ux5ACAiJZ9eP+Jda0GqsJtLMiHrgu9lY1fW1bHO2
0NDSkZCHumdPojibNvIpIGhqY3Le+BcT1WWBumE7Zl+jwQj3Ie2tS6ACgUb1AxxwJ/yXwSYxOc1m
VGr9MCQURjpe9Dcl06FI4Bo3q3wGDF4MJFldrOIuGLVkF0ADDJJ6s5o+xWhG/DYmh9i8uVnmtbdU
u3TWxe+iR8k5kRl53GzplxPu4sq2gvP8aQrstFf2i8jvU1NYRIhkF//Fat/Fp0XYZ2p6MfoHdVLs
8weyxt76yhxQaQL6ueNRn4FjQKvsZzfyCrtwpbJzG1FE7SHQb8gDUGcTX1nbzW/ARb3zt74VS8n2
q0FwhCxvDxBYnU+rrH8eGswvqEBTh493HNd4VzycBR0WUsoqBHOpEuNphx0MfMbl/LWrJ8v8CGvI
msN93ZASfEnNLfyWcK4k4en0+wP9BinDVhlif2erZqQqPT74meE2AM/uIlfupQb5GB2BDZnJqG6u
x+Pho+wqP33L/WvAE8f51YEhbgs6s16v5skBGVjguvGz4Vlj6fK5MMNAR+DQkTVeNxLX209JeHZv
1nwPLKubr5HSJP15fjla2R0qNf5WYOHxlyr3jpKiFzUgTPCjNCg6rEFnxCrEf8FYcFelVklLSFLF
S0ouJKrzWIgH7alCz/9P7R2PvISVrLk0NvckcyBq1t04kGKWZ3S4lb0Yiob3JQ0MZpCXdfLf53m/
WAf55Sgu7XzJv0v/ukSeShkWXpjM6R69+GFaQv1KVZr68l4uKflmgXcaMST1o94mjUuVTG0v1sM2
2bkT7daBuExDosynUaMEkHsWF+FrtbjCIkdYsDbhr6AkS/1zKhMO7uZynivJxCiKEol9hd0kA62i
XEu16X/JguPAxP50EOExsudwO56Nm6uM+LxmE8k9SOsE2AyP2Ys/mjSlsmyJoh4pm22eXsddiiti
wiGC0xoKqIySjn2gOQYPhjbR7UicWAEKqkrGoiF+gp7hwvrTLqWu2itoiQWv80wYXQzgcIwxPFOn
a4OYIsX/7EMtL4WscIHaoqrZrgsddZsVrtZNsic9rAP0yrE3tJ6SFyxcfoUyMiD7aR10VRgTTC0A
8C0/a3vqjXXiJTFy0o1LiA+7dST2eLUBgvKwcgIyU3UqzVDU+5w5LNxhVXENr6SPvYj6dX8bfrAq
rAJsgER+vnRFaJc8pJKfGmPgIDcqIuBy6pOLSJLJ9PMrmFYRhGfud5oXbb60n5BCKYHq7O0UQV3w
nKPnc+n2+LOYW/xq9i1JdoQWtgZMvgNh4WlkNisTmVkJ/WVsQ18akY8ESvsJ49cuexD29011Rs2t
2b7RBmezpmkVvO8m+aMdHOOXS7xq//qt8DZnOLJDwbum4d6WVN3Ih8LdWRNDBtadh4II6U4dpTDu
mf2GzU7PU+NsLUgNsN/gTllwYD39Qf9rVW5eTTH7UNjhazMndP5CulzF0Cnbn/96O91uMY9siw/r
tlskzZUAxNfUIJsVme/1HeRVGk0qnJ2nToj/5K46Tc/ooJy6+N5m4GcA7SAdvYPZCgCNZtntYfWt
AMQhClDbVko4cee/E9r+XlD7rX0Xd4DJ6heXzW/d5PfphCqsvrf4yhTGa4DbNkK2ubS77ghMjJPv
hs9EXq7derm2OaOor2fsk7eccz0bgp5jV5kqxU9y4RDcIn4jU9YR530BCNlsdzehHIJYu06/s54+
M+N7+aRByhphmAfGWoz5cD4j+1JBeAr1GUx7TWgC9iwpt5HrEXTO7vSj5XzxZ+opN5y7gd3mlyFn
k4z4Lyr/gdxPhsEM9w4gUAVnmR71t7SoMl6w6GwjtKtKmxlqfnyArbYsMw7zixjnp//6hWrIqL6S
ZzcUvzvYVcGy9ycXg9C/4QiUjmjOAp6mGnJCCKnmc6iMlnqxCBOcaqusM0HDc6emjy+/G5Ey6pJe
U+GY7xm1z8GClqnqIVM6g3s1R8jzpq0TqEdDW9IrxR6tL7xcTj5nTmkmLjlt9h/77gxZz7vzh1aF
+/f3tTtfb9SU3hfacIq1oOpNx/Fq6VCTc/PSlDnH2D8zejGHSeacPfQe5yf/nuskRi2fYK4eYpAm
sySUzgn2ebChIPKQCcZJmGi7DLu/1+vFijdv+s4rtBR/BBXhX48xv58e5Q5iRlhmPC7tODD1Z+63
LFmSj7cTAXnpfrUTOmyDxxMzfyDrzi2PBiTXyM7itCKE660Yfj1PAsFpErGG9B9TwKQDUVN375fb
Y7mC0y22j5VRWKn7nk0UG/iC05pc/m168UzxB483dwI+46JJyRmj1YbE2yudVbOW5FwGye+LSTQQ
0oMEJ5EaytWjR/a3AWBvlH0JJJg7vQk5V4aiGx4VoPa0Ua1KPyVENFlJa/8tF2V6KGk0O/uRK1Hi
9Iox62bLzpDFZBMD+owc8BgaeDaumk6sG8U7IkKndfLMhfROLTqXpCvVsnwSIwKT6nkcFjHv+3rf
FYCmRtQJf57FlaE8No1QDQv6/C3rBOeDu5GkuzGbkuZh0lvfm52JlDv55ggl9qR2P+S0NO4MHM87
4qjmfoOQEoXKxlxhkAq8hfT/CkdDc53JfObTtVU2TF6Jr/61JhBPuee1PoR5a3VDFf4ZeTxBODk9
eYDGb79jyCIOG8chJCaIiHadPdsGkyBE+H2Cc2z8sSNNgjMnLPm5fyU7nAUOQLD+Civb1jK0KHPb
ZeQPSNbfUdQnknJQbD+VlHo78gFGUPl+cIxQbwSK4tXTV538EnwpcfJMy1qxpQ9QNegT00H1JF18
n5mM5wHReLbJoPlmLZpkwjuBuZP2ri3ZE8XWvQh5zeJ4/hnkWTF7f9YiQqTEBancnM1wl88eDK2J
jW7ff3iqOozZRtY+FGSBlJKZ9BG+cnqGyoB27Bk1WNyFA0cFqDU5FkNcbxGmYDNDrVOg4EJrI3xW
nFoNbQko10n8PA6IY/FInS8oMMsfzPP1V0cy7NRLL3nkltusl4crwoDVEgLzB52FI9K0NX/HfQc1
VMYBCMgj5/QWkjQQkTAYUs17zhPkobE6b2/tbd2Xz303Iv1y5dAP3asO+wqldXHn1VbyrLzuU29f
JEQF6EOwQyhsDiRrGaRDzofJnfeYKaMrF5eOu17v7Dmyn5/58nI7tkbCx8jNyAxru8ilCofo/jHN
Cy7ympEcDDEj5Ay7Wcg9T4awVXRN4KoJyVNixnHRa1CUnI4kJiFoo7Uk9tDGG8CaZ97kyWLtzfwR
J2GX+pKaYUJMgzTH/W7fldF6xm35SzYtIHgfM9Y67zQ2KpDWYyu5XnN/7M5X43noK5tlE5NCwx2o
pSUtpM+RMcLBkY7pv+AX6SXH6a0aUBnV3hcQakZSRUMWwfHtkGB2ivEsbX+P7GnmgKYJhXA4t0BZ
/KHZmQ+MAWJ6+NRM6uJ0SWyqvgWOhvrZTJ9XELO+egXGhuuOaWtwbfISgvohO7WR5mJ8gPscDOal
2um557vYKVmPbe5DnHdbSAc49oLMsKxOTftWY1rezN+5U46gvlXNc5OzG4cl+SYcyPq96w3JnvlV
6HQhSgatEkKZqB0r4qlSB4K0ZOBg9yCyLh6jG45C9MRioafNk+Ll9katrLOvW1gZV2qfvma3kWlz
vJGUP6wOlpvyPDYDJk4OlfmcIWr4fMDU9wrsUBCnQYzWqxz96b/zZ8oyjlPMwsNrZawLOmROqlkl
2cSpi9OYGiUEFLtMI2TjRn11duRLoxLHOfxGMNw6P7+hlw4Z75IccWKEAaP9utC0mYlLcf0s1u1l
1765ec8jg3cBbgiX3j08DlLQsT3adAJemZybwN2TyuzVKfEhuEFxccS0eQgnWkgq96gfDIGTXWQG
ycZFucZMrg7w2VjqzBw/E1QD4rEX7fxjvgHrpcCVyd+yqmSm4SpJboUEM+BQSskt35q78qNOBYBM
f0NAm6OG1APTpU8X8VBY0MmXgeNgdl4PHm6Nb8GtscLzwG4hPdzkY9ZZXs/CnVTdO/ZHyF7Az5K/
NyXvr3aCIg19aV6BKQwxU4OqcbqBJjgcNpkYGA0vFrAqrEs1N2jAiYD9WHVTUWFx7VGcGcMvn48J
TFHkOMhX12NtwZFKsL/MJW/tBWKdo94fo0uVwVrQEHSs0NA79WsEFoNzO/Ur6wNa5kAhA3YXeHIJ
XITJvLf45TVDf7LHJRUxGVAdMkUUXyZS+0wcPJai9IpaEF9ILYw11DLtRxDrGp0AwNQsp4KuzZUH
U0CSzQU50kRdP4ED+U1x5lIKTZL5SMNLpKmynWvEYWOe9RfYDPf6ksQ/WhCFYBmginjFotO6gHHD
4dRxGW8r2NlauunO0AucUXVf50lZuw4S7R8GdOqBt+72jxAmUohqzxf37/IJxduXycG3a02S5zoT
XDCy9VCIYeMItqmWbJ+OKw9IfN6KCFBiSENhV2eTfuoh8dkMlA4iNYtNRnIZRjrHF7QTGiqNXVUT
/97Zsp8iV01AmyId3kPUel2db+MmsvKEdI09lodhtAUDnNjIXVKYkl4mee63c5quAYxg6K4o0T+n
E4NmqJZMomV4qIV7/ccgsZlalLewXOyu2pyZrvmN3XlA9wOtHDNAhKj+6eTDue25f/aZYd25Z4+X
BFxnYgl9/S+jjLH3fRnHuH6eVjjxBJbdu4LnsgtLcFuiqcZLgZgF5u6fQg3LMjIl9vkqkTrlM6Ba
ThbCRh4PBqf4eeT8vEdB+iqVaazgot0cLmllgUpAXzQg1h4VDzn81T/bx1COcePIpFrV6gJOt+eN
oXn5vn8cVeZe01EhzvIQiWPe0WOa8s0jZHLdX0rJbZZdJFdADcdaAdGMiYRQoW6tTn+mnm33oQLy
sMQ3Ggbl/9lq6WpkargbVRDAfH51mmDkqYeCU9LXURj3x5MqJYtL9oYv28f3zlfGoufyz8Ycb9pE
oRLdgkxFE+3y+Qp9E+canTDJXTQSDcBwF+znqYkc+E5c2Ckef2HQXuqG7Gvr1gB/knZzJQq4xTRr
Mk75Rs/GI8iU/m8PyIiwq9IEkASz8BNEC15f/Be3/o6mmwIDNoTBrdy+xNgg9HRzNBNjFKV4FAeq
WpTAQ3IDooWci7bPT9fKOW2X/JQDp1DdAviLmJfYsboVEvbhIbWjSEO5BzvXEjwqNOFt0vT4fROS
7EveGSbCTouPqYL/klOLuLjZHpDJBCGrh04rKFfRMGaEFYvL9iEDjHSByr0B7Zj2O8AJupXo4aPW
NsE3YCoI/fQavZf3uIA7RDtV+oWxzsKbkWzn+FizXP/puJAhRJJGSoNfAyRmUQlaLNe1Qiqzp5yd
uyneRUa+GoJ4/uemf9mu22XmqRhRi4hygKdzAhJx+ot+xiZuAdiqsiv4pDWVppl4aoF/dsM6fB3J
cAxfDgxznYknCUQO8WO2CM1P3EHNgPe92pMxyhlAGMRSTe9Ado8PXdZ5HtkzNo4A1RfuTBCvTbFB
PoaRj5sNUlEJW7tfUPLDaddnKxQyKqVRGeHuxJyXEBIZrFiOQQ6pKJGQIZn6n0wLwxlS2RVhibSY
13PaepzwhQ5BRtt7ycFilOobVk3ce4QExie7nF1DnrTK4DZ4sOUpzskYXcHupYL/xP3If8RyLBgm
K46ymaugIVi4F8xpchVC+YNcoAyhD/g9julGVNZB0BGlsTX+ok11SbbYc91iXY2LkFYjw78skv6k
spVgQDVcP8UzACG3pWr1hRLLB6VPG2DQUsGWQDe1iHEiIS0Clm8VSSh8KdMaTHhPz45Y6HbOxAb/
CMO3Jxgz9kFGE4NY5clrvPSv/td0d5PfMSV3PttmZw5CHQvYK8jrrQV9pGDusmdJnBrikDweQo1N
coQrNzhPJCxFdjsd3tro9IFthcL9x1cZgaMA45ypz/DC0fI1Irv8dQ+OPKKB3WrMbebAtaYa1Ntf
8HDeRMw8iZJWjj8+sgZPkcfUpDeCegz3ebGlw8mrJMikohkPZSCOTP1HdE5OE7CQxflfoIHPqtve
7PpRw2ucyEDgsivQ02YAWUq1KIIrKZU7mRo4z+5dQIApLQ3xCL+qSGp6NmkJKK60Eyk9rlC/xJp7
MUDh/cKjag/GiYV+8ae2jvxEXxGftrkS0dGYOivKgGK908vHHDqioUyhnQZTFI/UTV2SvkdsnauP
OOiw33f8jPgtpjbewEonc7gk3674fEFPiS9c8qdY4uirHcPI47ZoAoWO4iiTrvwpHI/rDCZ5HfXj
D0BUE9bGxYA6RKSyRLIm41YsnsKdHqExPorqPNrVRH+I1TugySSWFCI9K3C5OZOxuyAWy1391s4L
NPajdcSnU/wKtsI8TPjNlPES2q/38P+N1m1TbQim9JJHkoaWJBfbdHPqerO4c2YL1KHVTpEO/p2e
Z9+Lb/UhenOcHf98QHulxpvVkezNypSQJQ7i6PCucMyAsh+VQtczh0psh6OMSUqQu1GupDrK0HF3
Wa5mQpdUesUgimoHfxsWNxtItSj7sA1UHAocFAWPteTSWVMKH0i4QlEEql9Jlsj+7+EsAxA1G7IO
g9mXB76VzWsNvKcQMKXjy2E7HNhnYWnlociYYiQkXJ9u6UDViWFaEBK10FX8PI3KMLEmcIt/6yP9
czC6uPvju+ypxgSSd110A3CAZ8vuP1naXC25r8bcsjZEJZeKHnnuofqhDk/woUjmWhRyAJn4yIfT
PcgbDk4JCa2PUMF4Jn63UxiyB5wJI/R+YCAzPmiKMdVbU8htU9ngblSqdmfmO4pkKJnFjdSanUPR
pVYnJpM76tiuChJk/g6ORO1Xz7T/Cz9svHwZlXJ/2NtK7g8Qvt6E5thIHhuU8Vbfm4Dg0J2XpTTZ
q43jDRUgyk+c5YjmIx2F53UcAiTU42AR5iHiCP4QcXlrT/lWgVA3+Ue01hdWXnyYX7tdgsHyHmgE
womEo22IuO7XwcsVUdf54sGH+EdOimM5r20flavA+J9XmDwKXPAdjjuJRUaAOHpsh1x2+MhWlCFV
jx5T+rKGDfwggSbiXOIgUaa80qpK15T35ZWMCIXUSOa2a2fuyMqX8NhXWviSkFpkeeU6uiNlN3yn
zAUjyowCLQCWQ8737B819YQseQrXICho8sgooltFk9QqmAc/+f6JHhCcMmIrbtAnZR3lgwgTFmGw
0RFilIsTV6z400PHqWx/Awg6SeXWQSMg8G0++b1R5PrgyYz0Q+DAXh+LDVlVZ2aauopmeaKjVRT1
Hfra1u+JKHXurqcZmc05qtSadd3EVqXISRCvu3wKaboltwplwiZQp/6XkVWMNQ8PquqQQEsC6TR7
AoX067xnp4gPTScYCocXVSHL7+OYdaYXXh7YxmKoOFbgD9q9fL1GsWRX5JbxSkW7qCBTXuTU+dc4
kw5tl7Xh7oPgbBD74n2W1amAXLMtvgwqeuQIoovNJs8rYi2ksIpUDYQ6qUEIQhe1CihVNtgub7Gy
kQKrajwNNko3F7CLmQwM0Cujd3rr7wNeA5BJ/olhEc53YpMMxk2mREmHJs7asctQemHnR1kPHDwV
kXQ4lBimnnu0IjXhkhmJKYxqF8Zsb8gareegrxnUdZ7iQjNaPkfJSEYhyr7nPA0V+64ksUX7Atln
9IEoSGMznKLCfwbWrSb8OpA08gyNdcljvG5uxkwu5PNoYDrSm5PThXD4OUW9+isCr12smsk6RWKD
yk9fFzHZSMpF96NPsbyJDmzDHgt/P1Zz5e7b+G2zmz1Z+sUG/7DUrFTSerO2Llw9RjVVV6rbNQLh
tfy7qQKEVkQ27m018Vw463kOTDLLMrkGJIMxlSaucWp75hBEyLR4NoGX/vxxREj1vMls0bWh6L2j
IWd5U+wCQubrPWZKmf5RiWVw/vFiU0gae/wzxJ6SOnoAuKp0b3/50+2f5PYU+T4gLL6n3+ipL2b4
/GTAoxeOT5kf6ch3RZrjhKhFuxFg+QZ0db4jDBx0L0tYmQkwiYX1d/oG5pyc+Ps5Nwr1sS2rC7gA
YT2DQEAiTKEqxpYP9iHTbhI0svpvUKBxgdSlAU4AvE0JBOpxTr7XnvZbiukRvBKe3wXK+jMgBFf8
PUQ1Z/nim71a803I6qWiDcLqitz+TAO6G0ZfKUuDPbUA4GqAciSjIMQ6MZch2awmTfRaFTeYgmvu
ibYv4Qg62EFNQy3e8mJJo8EHqUsCJ5kpzkAJNOJDAxxFzOPlptLesh/FwX1oHWlFq4AxmHpPVIUx
wM2MnqVYB6dom46+BNZUCPz9QAJ4UIQm1h35P2DtrwFfseb/T0sKQgSeRRa345HX/7q810gHzaaN
vUxkeYUw8pnDjV3OmJdVrvrIEyZ0TUQ5yE6JYfiH/aTBXgZYGjFm+ZZ1puNIKpu8j1R/2+Vh20fa
Pp8s3q6ooWEabl2SvPFXODclmTuQzejWvFCZ27BSMresK0yffpckxS2RbUbQH73rBRt182JSVsTg
43cYN8Y4qNwikYlWUOVN+SouepYYsJSk5W+9Sua5YekFg69BjhQJ0jzg1Cz1SFkn0gPWVv4YM5Ot
T8HgpWimOUeBFYpnpr+uZ1ZbjFcDRhl6tP3lJJSrcKI34I48R3+XC2zXBnd7LCoGV5dBHptqigTj
7uWf3mURYTEYZ6gct7cGOksYIeitwrp1eh+Ll6WlAm0LdktVsPtWEdwSzb9eI4FEPstZ0qNivHei
cZ1z3IqY6gF1X1154PBOy5+WEbmkpblRcBgNqtRIJ1wg5we6btx+Xg5INY8vmNI57g74NJ9594UC
1qZcvwKIXs0WUq3S5AcHNfKsC1xYCuCCy4hiUaQlk9i/i/4RAs1URPXbIgI3gJVCttrbBqGIUvU+
Z5q7DsM4BMKH0gsoIAjOseAH+W4yhw/KUJRWVOiz8baAjvMkjpHMrwsbmDMxyeyHHRamwqp1zsh4
hGjRK6plvsYLDZ+4oV5Rt+1YjqCWN/IZwzuBs//4VisLca3ned6Hy1ARDE63n/M9YWxwdbPllFuw
5m408y1+NomInPwt7jM7iuMk08pZI2MVxNCjZ//IMVFHhfO0s8tJcssA2Bberksn/ibXUcPd543P
pB3Lq5ngVjf0zreeQcv2LXtAthTgf/ctC7eEWrq3QuOwpQyJN+1ApLX1vuP0WF4HZGcdPYFRvRRE
8U5L9IwlizKWcZEyOP2Kw5j638o65mtF1COBr9/u3fLRKeMxdpoohxyQAo3yRMGwPi4sELnecYw6
2T2Ky5kGZ150kKt3Z+zPmnNz8F8EKj3NyAopClOMRqVshDfkFkWNwOaQojghGQMJD36vpTHccM1p
rfQWtcerI+sehNi6ccwC7hXgOzpLkBtXU+Os9Pb6DKypYy2Pv81N2b9BQ3zqS2FUV/CIXGi2vJka
+/NZ0shVDLLL0zfHCAL/cg4bBc822VPDZ5jhtTXMRXNVnLPOgiz6Yb/sEwAntZCXBgAIgk1sV8w3
awrJnurnnSy+8uB0W406LPbYW5KISvMWAPI7w5Z5FkplzKC1QHULKqfgjPCRSL1diwzZeNnF7V6k
DBexdC3Qv5ahkxWkVTJXixtB/7Zw39pAxzNfIXkDLud96qixF3EloaaFJWZ7zVIM5hC3NkHNaV0x
kXUCmGHdpq3xBVmeODADhCqSQl8Dx1ObWCxggCXl6AZRB2BGTyjhhVNOXP8iiQegOzwIH8YB5k8z
r4hjdrhhSReyyQVxheDKpQFn33wB9PfOCXaPUWTqmLmAG2gMuN91Yv34v2kGxAPaCLmojEpXYp4o
u6740zFdre5a3chNYY7Ecy/Uw2Ha+pNGqYGTkIOQhC7+N/HP3ghuTbmk72DQTA498+W/rn9ywl+A
iPMEU9gXOMLOw3oz+OubQQ+15xURLKseRzJmUgpLgrglGy2zv5Tc08SIcDAxSGxuUoLUE8/OZNYs
8ew/DGkuCqPdJlSFNKrNia5ejpmwbq3VYQyBkhljBHzHuO235S+yNO548EwXr++aF+96AtVfzN9e
W18Qd+pyCYn275jFNBbzMSqeWfkn8JWBdJ9ohyoyOFp9quTbaFCsN5Upikb9K8DvXzPOwyismbLT
dihhdlaFwxB0O+wPPQRuoBElRk/bgU8z57WbCCAkEuxn0NCKoKlgkRv5PJAda8dmFJhOagRAVdGF
ZQrIDH3+bLiQis6y9S5YoXKJZEZ2T61Y+0aKS2BievEuUKUaFRXyhbJ+MaA1yR6CRvl8qsuZl8+T
OxP5gagMhQYUy/lJP8mVhA0M6/LqVEX9IxFdKSO8Z+Z01Jmevbpj2c4of3BBWhbjEVYty8hI+sIf
zpJV//OSNrOIUBJPgMP8lOIbDsN3BzbXsdzINRfESZpLcnoAlfx+R+UFKyT4qM3+IG+o5BHBQFkJ
rW/QyegoOFYbIsdYrI4YFOEd4Vtc0AJciPWyQkUOnjqrdl8QdULfYRaWn7uf87LzVxhtjcObPlCk
hPqttMewslFdnyjBe+IZxuwcv2mlxTgvw74MjkT9eaLa3gRrsvIryPJwwmpo6O3/ghdEs5t84Qb+
yL5jhVvJt/tVOalGGIVqvgZbQL/kR/VsB7mRwd7xa40j71D5xie00p5QKbT9DCrQi7LnAV7ysfAI
bDHKwnhswLz8A07xCHPdp3tAh6DdGpcbPtW3n6MNjixpQUC1NNHCUYvOe+OBH8vOrzeT+4FgmwRp
w3xYDwoAKa2UvdtcjKrlX7WoKim3yoLJjim3SnmvQzAtsPaBMJ4tJpWqp6jRBLu+1NS1vAH4x2q8
3Pe1fmg253HXdCnkusyOIitpsyuJqVi3keJErfZh/Y+QtEKV9nC6ZbBMqQIKR2XgRq0b53RWWdsm
WkWcT02D8klPvUgNs5PZLPzNhV7dgw+nfu+T9La4zdgJ/L7hyCk+ULjLtqt3DL8aUNa+9EZYwu21
iuVLNHdnMQFWPqR/zUh/CpL0w7tdrxbVg1RyMWQ9EnM3dcR8IlJJhbN41myMplsvTSYb14X4ojFL
aesl3x/EyA+qspBcdJh6tredbtd8YpWpqi7/fiHIooDptQ2PERphtr42zUDmgvPThxn5dduKECNQ
hC0R7dwTKDe0IeL1l7kpZYGs7YoY/5DtPdPQtKO0zKGoZqkVazqvKXY6fsCbePZUdH8YT/ln7qYx
+JdYrNG2U8Ev3q9yWv/tbiw0mRAJpUuHCWsqYGMPEgiOjXC+KKV6u2yWej0QhmS6ZB2+GE8aV4C+
ASEe3Ry8WjLKdQp+ySnVKUzDXxgaHQOHqK6YIwezOoeLDDjkeI/W6+nmjre4s0mlPEveRwwnSR9c
/VRQbpwknsvcnS9nhdtf13Jhgxs1XYHmXMfJXpU5rmnTqVjM0YHuWXbeGjYjp4cfR6QbZ9OpGFuu
GiSoZCMtzGlBt9um057NpxWUiefRS1FZooheSc/PRjHHup3Jl6z6Vvx4fnQAnacc9J9p5wMBAJcI
/5fjAJtt17VL9V5LxLKFcaseLHnKz8i46kqLneRBcElgFc1fg5Nk9Eh5DTww2KarEmzwWTMzyz0T
A/bi/7ZLJxc6r7tD9yVJ2GhWlspIZQpxCRg0fGlVfQXdrrRGU9cOvPnBHromj1RPN8WHFTNcO6Ru
3CTKEl9KOU6bkHdX5g/Grec53wC9GI24VAgyYRED45N/VpTCwB0hvNIX3cQE0s5zkggMFsaFlcBf
zv5wdgu7kiQx8DAMam7wg30YgErEuWLinJ8rqMFBiwvbwoJmolTwBMgx/TzyfM7rC0jjNHIEdNA3
JE9qOd0tKzcmniZJewXVrsUWTihTjEosDNOpZ9GOrAALVV+29AVDqpTYa10iC1EokGjBIbFSeHGm
xfCebBE+L4uD4aze2O68JLJcEoPPIhyyLAUF+MlH5i/JqQMv8tAKFgzREQsABULgVW+DtEeK1WlJ
HX04WW3bdgrDGGB4VT+ZkwR7m4PgnWCg4+wnSn9H+svE5lGeV4+u0kb6H9xtvPjC8QdYsaWk6k/k
ecl13nJSY9hgr1+kcwY5XTKto8veKPS44qVe2iLjQ42OKK7oWX3PbSu022YGEEfRbkJImATV8qRE
TN7OwRbMaCzMakiOIO+r3gcDE4bHiVlYstrjVcfPJNrINnuFR1xrM6xR1LdfRDkDjGmlIkHf5CM0
xKKB10HpWvJSrujvaiTwHrUjipPku9o2HkPAfspZ2iShve9ZUCgm5gG1u20m//uLF5VAHqvbexaS
zpZbwOcWuy8zG7ZIDqDi6hSo/iLmKzlATaBsgbKZouztc1wp/9YFq1Bztuzx42IGpaCSZkJwliu2
mm/Rmi523Agigke0N4COefTTbZfZ4cUnw23X8L0oSuGTMFdWZgP+aJt5VV535qZpAWxH0mAlZeT4
ORHJqpcYedepMtTJmx48h60s0cLNvFvfeOdFr8bwPGCD5nN588/WCG2WXxBKQyd6wyi4CxBdSuDM
Uy3yNVKV+jJ7+lAg5PGIjl/Y+qZRxsuTvR/xuiFa7Sw7uwPrxkM0lKZHyd8Spz2p3n+yXeBT+q3a
I0Hvi8Q8GRkLY/AeRzzJI1hhEzOMrqDgZkaTGSi4raRIOQrPnb1oI7l2U0lJhFmvfjgw7Z5n/Ll6
lumvbzEcsgCXgzlxOmKaC1Ph1e65wAvWb310QzZjV7NsN4FWTtFxcRbb+BRepdkhSADjPDW07tTQ
TNfOLiRbitqS5TbF28F/cRErve3pg0X+brogZDrxbHzq1UZvcobA1wUsjVTrG5EgON5MvfPquJP/
93qBXaa/AF/eYHhWw8LlRb9MctOYL/hTM96raRcmHaG9JYny4Pi+LACaqWXCBBk1Q41Y0kTUcO99
OmVD4Iotfcvjjn1ei+JMwOLLAgUhO18bPRCTt5Wt4Qa6DKLwF4aPXlz4lltqRqwHQDrlWl48gVDS
vGQdxiTnoar8DR8fGJJmPaZwSy693VgarR5Nm3C3ynARfWXJqi48WbdQIks+wfs5X+Ec0fl/Qqfd
XS8IelZ0nA8YLUculcZpugcg7WjgV6LpyYoowzVZ5lv+CGrbClof58x/i2nF++DrUxpx/3qhTOi3
rhJTQol64QI7dthME7nFF/gdIcpymdmVWLqz5QUQmtMHU3ZVQh1Ee3a/l+v1qk9Pc1HrYLqOOUSW
F6HkjGfwWVQsUElpRJ8HUGylZvPu+3sy/KTLNpaYBtQ3eX/fsB+T4xKsO66jngwOxNDm7AA3jH3N
ToXa7pIf6IVyS1IkorPV5WXlSJCkoHwxWawHLPAEVmDJyuehk0bRDPeickfpzwvn6ikgqJeG1+IH
GnhXCrrkddoLJfkum+TU5sVWssif0e+VsyTdpGy2DVrJdC4rxujkefFhZ7e/0zTYZIfIWlBEkGJJ
52Gp8ljuI3bDud5CbuTvhV7X3X8VllVGRs7SHzcXM0Z8xU43OoNu7sizS7d9dpFz1cDpPQDs2wzH
JQ9CDwH0+J54LFPGJSlgn9YSbDoVQahnyg1g63+OC1LZS+tUVL9OyWkkKQ4FixqFCzvRX0JCnOVr
4ZMks+2Esfea3zkiM9iMEYoLo+mww9C/oE0LWnDW4diaSzpm3GehYxpKSPxI9bUsxWRoUZDum/H+
s+w7vw+VlLMrJWRFzX6FkHjS7YKYZSFQKsM0jj5f85zatAnk8/9z4MhJn5bSrE5drJE1MfxQvnWP
NEfLZtAr1N19pSu5Ap+2AhZgXnFkjGTtgui2pbUwo0jD+KYHrcsglwt2TC+KiDqZUuWzdYIliUnc
QR4MUnBvHL4UZ6DwxJOXHQ658Cjys4Tc8K5Qlma62mipveGR7FeOnFZ3TqZ9t0VlTGL5NybXFlJj
KSB+QmXGCRlj4DsNdIhmUgZYEblkRO9pbKNwQ5A6oxYfuo0sso8IPPStjDX2oaNfnjhhdYMdvLoB
wXnlkPvr/yFQjiNyx8pnchp2ZbR7Kl0R9nSqhIydVjROzSQEFimmT6YTfWVmrILz0RKgJRIBev2g
IA/qybZv1i2FjseVzAQyJ+QhH1Ag4eHNle3MT0Knm/GiA4IdiiXud55jXub6poasI2WY0YGtH9ZQ
x819kDj9tjGnEVOE64IwwOwmDcBi6l2lP5CELRdA6Jg78GqzZeU/KoDVSGeb9RxUkO/U5ztGrTER
xdcT987wZ882CDLMRfuuBOTBuOGzM7K9BmNTeuePV02+Ct8d6uBgr4GYSmsSJsZHOD8jUXSzeXwq
PXLxjiIVMSjMI5cqRjNuvQHI+bVuEl67FsGhtS8mGZVNQep2SlpYuk6+OlS43XwhakeS+GHPXQ25
GYFqYydhgOV+qhSo4orMFKWJw5hETLEGgsgHGlfxBckCkw6/2rVjtSqHvnsMc/ArXHnktonkpl4r
21JY/Bgj/79fzqAAPVzrxkmQkXkuL/W8ybt8cVR6REjEpUJ6EfTTI8ML8eDbB0MgWmSzfe9PuTC4
HRJ8LaYGaL7q+gcvgaUaCuKJQ+Ha8Rtj0i94I2QSYbUooeJg+uGkR0F6K6siEEebp1wJyDUkxIHA
5SBtqw5r7dYr5uWpC37yWHk2xwX4i9k8lruj2FK1A82Y/vZRjdrHA6mGBViGZjsaRUZ/4ajlpFzO
lX3KQwhObhm9eT8j96YkZBYtKS8KryBlGEVaPGtdYtqNvDHlEm3/gTYM+j3vpUqdi8DcxgvZ/Olt
IlN6fCYr0+6zVX7qCIWmBJKt/vyDEWSH4qchnmPd7HRLg7vdWmopPAgPBeahU17numdoAV7cDHtd
xoidaeJGDgObAlyTWpH5YDnC+B6clbHgEPiBYDJryUCMDRtYAfBn/bKnVbRqQpDp7WYPozra2ySX
DtuVnrrQgrXqKTrB9CYA8caroBWy+E2LQdXyaisXrPV3dpxr/ZUNSBALwg45SOa6iD2rPEzViURp
cBUzJIdmitT4pn+TEyQKnBqGEYO7IklHkgwG6leC0MVvC+AmoOuZLYevSKMXBLiQodMhzHfaT6W2
b0PgtuukoqiX4hJ+6ODeUQ303lMCHFqECH9dxLakERAKK19ZJAbGxfciflh0ntyqX48huTU/DjGa
IF4tQ3U9bofrE9lvL+1DbC1AtUxxmoFHpIBpAvr1T5+qLx9Bqx6UHNAvdjV3Fn02XnCZzNijfytB
bqddDykECt2bTmc6IZiluN4ymHkwif+zpButTVxYd6tQ8ioIJSosVAv0R+iXPoXnqiEkR6k+PBBN
bdfkj9zf50pAX7jjggSLfz/FC+QCLlkx44cebAjqEO7O5cAS61hSaMa+YraupVL8lLKQSrruQ/PY
GQDPWXx0GxiSzvLLCYEE1RhL3l6Rb6hHAQCzgZc/XdfPOvUYEtGhYhZ1byVWEeP9Hm1EH0DOKxcr
x57GlrLwxcXeNddxkL3K9lkwJvb+QmNaryAQMkJwvr+ATEd+MEEwrzbzvtNL5ZZI74LWsuIZ3kq/
phGPDLMvulPH+qga3/lY9pEeXGkt2UBtJvrkQpnTlywsidtxqI5Rq7zDcPLIU2FGc3e0yjqxN24z
1ISHwkPl6KSoRcVrEMRShZnraMo9siX2K31UsaXG5fMx53Q1Tyrd3Y15hG8Rzckm2vzHnaha8nNq
ZYVlTFUkhKuOAUGx23kmJMbtZfWXK2QgzIzYZIBvboo+JqRgF0P8EED4Cw3CW2cgZJfh1WaKAsAu
iXMzN0SQPWzg6Lv+nkuc0RIcaqM/lLmRvdgXqIo3URIX7PcU5BIZqSZ+Njhw3CiGg4EKOecL7ITu
7mBeib0UD6NXpGrFwOwsMoSOuof2Od0RRiwxEAZGvcu8nFebiWK8Q0HqaqmsfBhMO7K4cwRa+zpy
S6ixcRQoyTNqoIjsGKl5Bf53x73+/gWJhpMXzgvHltwXUn5/Dqf+g1PLgC+VZJUqkD4Yf24FC3vB
RcD81nTwbypbZ3EdbnI+8vx3B9U0F5dWv7yxjHZMl70hrJ+2zTOokTp/BgRAYj3w2eprIZPO0yB0
8jW8BvlPoltjIhUi2cC81G3jabGh7UseNQ+zN0QVmJsCorib95MucRXA+fJZ+bZbZdFVE0dckoM4
sXytpC44LwAu8djeefNabxVJ32A1XfL9siQxFeu2YY16m5+ms9UIvkHFKabXh8y7WQbwmfjbbOHN
NKCac1YApMo0HVJ3Hcn4w9kp+stY0Q07kUkLc44fM48rMIIBrs0olBaegFPmsujSew62BIu/oUeW
USR5fbI3EgUoMd6kDHKSE/ZwWT8vz6A+ADECeEIfxvsoDP3uxZJJQfDStnvoGZKxwZN2qAIR58qh
LkdOrPFUTOB85Sq1kmAPUvmmkSbHyML9uEE2faQIXNxWeds1E80dnGwjC3YvcyreTRXU7vOYXEcE
y6mqEr/IqxCFECHAD0GLHpWGxWfrNlV/dUkZFhHrmlQCh/TqKh2GW3y2Tk5KcQVZv5bdyM+pBOpk
5nge8JvO6/GpQym4Szk7ThEQlY+ccNHETgrrhCKI4fGQVDIC6dpyOTZrrHoa+GFz7SSTcQGfgWeK
Y4WTAcw3prdpvt8o5aY5sm+apxORe/s7sw+hsdpZgkxHrztSSNnQU3UG2Xk1NXMApCfHSVchXWKN
l6UYKWimW8GiUZEtgoyVL9DYNKstTjSVR8MK6a2zNaccChYo99bl9dZNnCesk9Uz1yKrdCxXDVo+
K4MoyjtVJ80mbNCxraaKmS/7LaoFI/LKCnJurLUwMTQUNKI1e/eOgFUM4wlDjMKwU5+Iiebc056h
6i5l8/8eHmRGjxNfHNE/yY97H3MrgkKPaGW5sRkvF+cqhHMsZG5WuC6gnPGPt6r5v8J2IlgCo+RE
VFmjpV5tnpJWTpA9Fm1JmBIuu5t5FxseSYeaZCG3Yme1/uOHDdT7mYEKvFy7hDhAa4D7ZNOhkwKa
/pZ1OP89SQ10YTc73EXO7Ezsbb/ItX28V0RKy1bKMp8DLCkSKAhLPRsc9kPp6FD3Jy4k1HWDB7wc
dMLSP1HCbFwmbByUZHwHuPVwUD1ssmjiz1JySyW9zZYLNQYDMYVU4n/ejFaqKjoGF01Y/ejHCqgo
ZC0ux9pvHWjBOcsilQeXR3tRWJeuWwRAKWLu7RWd0AlbG71ALjNpIvLVG5EQYGe5OodDUVAgxsCs
rFXAS0U9/ZJ+PcEgqrkQC+NyYXy5g4LXCzJJwyeJDK6mo4QSLAoibsMi+eSuhaLWuhDsWXyy/NGJ
RWVXfc7AY/K/hGmlC44rTXsBJ6cW1qWpgybjzvCqsr7oDwop8BSjaUBbGsRPc0Ne9ekOqIkFUS5v
Kxji0Jo1mPOpJZGcNdlagn0WFvzYR7FqJrU+X+k3908vbHBmbHLrCPvog4F7puWsnfGo3S+2lrzs
HqMkjuOjCg8OGJN5vv9WkbaSZA91fSi6a/76Ev9J/0vRHIZ6IdzlLwtzBt4As7C20YYvFbPTzP+S
8IfpodoxrKldUQSARP/zjtR6fSJz88sRQr0vaFov5tUJ0NYakys802hQcV0Jbc8h1vJbY+5tgnNj
PKa0TywvVzMX8riSRa9V1+O7MZEw3a/IwUXoBPX8nNThpXfe1CqTkS5trex6Tg0ZGJL9Zl1qW/dU
13mAZMNra8lvzGZB9lQOXS943LsPppeUv1GtO8ZUxfhqhlXi8QAFZ5fD1vtww0mD6U3P7ChOYmKH
IV3U2X+K0riQXajeu5nC/3VAL1htkUkn4z7xSIyYVcNP+mLYS97YqJJx80T7PN2boFBa0GOuatYh
IIcFM4mSnI5xfrlwKRdVjkamnxKCIDoHzC/my+DLbQxMzG1rpCkWQ1r1yL3oQqYLBK6Iabhdtb3f
uh9CjdqsHDlN4Zy10qfHqKEj6YfqVP5xSGPFL5khX7e7dBpk5z4xKJyL9WIx4R5L/wpN4FhX3FhS
iQu/Bkqt3HxRX1RyWx+WTLHWysEasINrUoglU+jMyLzoIYEbs5zYls8anJY9Q+VcowyPgcj/3C4G
U96VEw6ZVN7N9cgo1fIysfXCXyEvKshdyHbkwv4Sg7FJ29aamcZNLENNVbRZUI/E2vVg8mKOUEdq
FTNDcm6k6uDQy/4Q1WenLey3g1j2PsQP76GFJHJ3R4YHGiK/d8+61Lf+152qr1rBbgjsoAD7F/es
tNXFj5Z0xiWbt1H5YEPFKpN7ug7qcngUX7Vz0TPwlg2nQWTsug4v1f5rMP3gz9KhEKLXi1qy34Iw
17V0WopXLJ216e/oqaEl2Aw3AhhcjIybyYOukO843qVilH0LOYV3TV5vZA7pdYlhAcBjPki1wtV8
86rLEhdEyk2w68u0z4FiBWLpH8KPamH0LwzSRLQm4fif/4omBxrJjLCfieKZq6/BYpOTTEdQYIsg
47tL9/ju89K/yPzkBeTXdDx1xDIyv1ivnktvsmmm8PAXBdRNi8Eqscts6Kh3WH5wmCMl5bYPrppn
pg9utxP1HgambjyoHJm7SvOzjQjVdFrr+bvo7jFLffILNShmfw0H+qSY6L3OXPSvBc4M1jo2QtRX
oTnLnRB4UDuhsCEWxWdkTPYGG2e3N9+xN4hdk+X9KEXVLsF/LrpLqf+fDjsdnYFT8SEbTzhkmone
7GlRwKqiKXdRwBxqPQWnfBThemOtMcqzbIe97kgcn/+s2VCRPnmGQkeLkE649zd+fIe5C6+MyedB
yBOtH5CUfnyfxON6TWlQu5XTBKRlks2LxtYovbPqqWtr3Nhc//hRYr8wmgl3q2uD8652brrPiW0F
Blf/NP5qRr8n62CFqDdwdGho0++hoxlQBdZAsQhvMh85eruUZ54LlE4PdVF6Z+Aege3+mGwdfxsF
dzxqZcmTHey9b+G1otKxKjy8cIU0o3N+pIBwrb9uMhuBpSJHdHOMryZkX/9EiKpcSfQmeOvmWeHf
Xwi9n1JotN0bmBFni4WFs4pYOvN2MsAc414fssuXGz7KZv38UaVSf2xuCF984zo8mSazaPZr5VKy
/bJKJKCMJ8AH4Wm3ClGs/xzNsW9muTTOqC2xlzDZmPkEqIgXAterQZgTtDVpIHIP3qn6HVgjJhov
iRBy7BKkJg3Zdve9cSx1MIJSdgawi3P69yJadk5agRc3qgZ/Ay6cD3Jk7iFqxJrLpTc0WPLPRAjT
b8iygqtEyFoWugzQ3ELUkp5mj05fxigYsuZeip5gGQaqSNz7WwRA6ABDWtlbZWQ0ZXbDlqGSpGQX
ddrPnn1YZMdOMyRLYGQNrKK6pTaehuqsgpcfgyvF/Joa0BLBYLzWlMCZPMrGKrdFqlcweelN6HT1
f/6jeRmfyU9QhUTi+wyYatdxXMMBzhXpYeHxKEuQR5AOGAPMM9yb8FAet4qO5utsMNkJPsz6ZAEq
rnnQClga6lwNhxhAAG+Bn5izw8JD/qjApHAmeZVL4eS6X5i5Zra82U3okOnhcLS4yCZhKEtKPxZt
pS4PjRLNapp9hqthn0CinGF8YGJFG5D3D0c0C0zahLncaDt1AjW8lDnWQnSl4KXmnIgP4/H9KnwT
XkLgVivKwpTqYrj9/Ls64G232Z6OWgSMwiSSjItwqkfG/TmYlRxJiIJc+dqH3JK8s+gJ/CZTSq02
U7vPwM3G41Bv5PUxLTG4fkbI/m/XXX7TUgmHAYdCGSXA0b0WvDkR56+x9TiR5pKv8CRY5uRrF47S
LeAaXMLYe2hQL1BhMErnz/SyMpharSSR2L2GeZ8w21GmVfUSvhXvdWYPJT1c7BPi16zOmb9XShsS
B1sjdz8pnh6JCQHbfaYRHJbAe4q9tr50DU08e0qYalhwt4cEPLyBcd2tmb64D/spQ3RqfvbsNUAg
FM0CGbDXSj1d/hx/O3ZcwZlVh9c2jzNq2EfNXwfekCqM4+33SLKxN3U0IWHfiuJGS7jQcxXOZYJV
A3rSOXKkkM8eQWXQcVmtUvSpBPry/+FRuTa4ER108bo7qb/ZKWRmWCzhfL7lCXzSVy9oW9PZSXM8
Tt/7/Zjg7BFqhgLOt0BHmP9sKiIbKGQKE1IhW9A5f3P80lo/Lt5VIYo5RDlxHA6EQIj6hIfeP5l5
NNx3ReXbcAqAiym3KHb5TyLPjUrphFjAm+RbyURsDpIaXq0vHMAzrCwQXL8Q0S8YDaz1iJcW3IMU
TLZQdeytssliXtd6oVSgAvwkkdKOawVR4MjS4dNZL7tAF+nzbO7x+f3UwF2S0Qh31/6liOGVgOp3
R1Bv0qXAaRTuymNpNZ55dVdkKEkSrL6fLJZ9FguTsgvJ8VV04a8wxgiUXUK/dpQiTylKDl8ZVVDE
VYRhEaAd4LBX19Wl5OiNN7cpCiGMZr4cLYpBOcrOK1hErGSaVm7xnHK8c+bqJiB1IFh9MCYaZILm
BWWo0nURyFXvNePmqwE6mLyvFrhAqoPS98gnGtBIuQ7zDcw/zXHGvJoQMSYXUA2585dFchXN970t
AiG51Mfj5KoPgih/VVLKTuK28vC7bOpa8w0BmYLTgS6vwKrWrRky/DWJAV9pUxlyUXeSjd9zT8+X
vUaiiGM/HVp/eaACt2NbWOwEL+Fsa/lfWbDyZD3EH+l2zp9TO2PvHh/Fllth66WYVPHgjIHFMR9r
6H67vnBuMXTQIiAkAzGRMiDsCRiGm11etC5ESo5+F9zdU6znguJRNX/ZjuLvJr9hM9cwzMg6BHz/
zOyYvrC7XPTKA0NfTVislQRNf+eyamz6Ir55X7Gh67l7VF2rpKF/LWJb5yJwfBYpGbjgDUgi0bhA
TFGNrYoLaPV9A8jTCrEppFeGoxZs+p6/WeGSdPnC7uTTVowgW4U2FoiXFEf8FTI2//Nv15U2rDsL
qzZXwNxSWVPx95BXtGAIRewseL3DYhvrvt67s+GaTpEoK/qYbyotCwoJKYWeZVdqsAH34PUBpdjb
9xYHjtSsU2ZdZPSp7wAEHDKRCk+ZDxuKDHKbqLizhgPvLrVqMLcPEPqvUbevwfWE2+zHnYl5d+AM
acOvx4P1G07/zLLmaVWcLgoUlJRbQf9a578duz70h15o0/CPriL4xXuJc6FT200sUwiFWHeAXgSN
Zim5n8BUBtthW2xm4mY7SNhV6YVZy+9dn78SZiouQl+I0HU+z6dvKHz85mP6cp645yaA8vKaHM05
cXlxszZNzxx22gQ1Yu9bZuFdj0bBJamtX6nuAy/71jBypRqUnRnL+CSFljdkXMy1jwSMOnprLnb6
Pp7qxaPdL9yeZHoq0tKP+mNrQ42nHmAaXetJGhbThrOR4MJDy2YlKXmOvCILQBlx6TK3vBw7xw/I
RgbjmG2+ZmAtqstabb5dy/3xIAsqojd+UcF5m8G/4z78WDDaplkoYpyTvyBb02Aw46caZrQAwxQh
ev8qvKlzuhcytUb62x2roT64dtSxienFSkxxBBw8snH5aDY9uFL3V13FWleNruignWK+1bP+ITQb
YeGlCF9Msno0mHDR70T2N4euOGh2Ni7x5vu9Njhms5YErFuolb+fxsy72EXzB4AqYooM6kzkGSSV
xVJ7UFeJuLTzrzAx9mt1uaJOalJhMHgg5HRqei/LBPt6IP++klBI2+FOMgoR1rSLEqVGtYnejQIT
wu2A4Gf6tCfeUs7i73bXfoyzHEJG9gsb7yAHEKiMqsPRpcQ7n/rZpq9f4N1OG1OmxX8F7CrdI5oA
kkJCEMRjSG6qN/pQacsNcTMtSmEaze7D9XqhONGfDoJJPD0ODHAUrcXC6WWQIh0n6Y1C5vpYM8N5
dPlAemg2Q1tK+GXxDucjXxXb7BMQxIxpfrHlRYPfh5nD4OdvvJATZQEIMxv9aKSqgByGRgag8K1V
myjuvsR+6gIRG3jGTRWnmQ4qNhdjTB95Cka8/PkJv+KWLL1Aqu/jnBXg+SbZ4GS43NSHre1fGQlY
9AEkLWNX8nhOOkz89vPNv5NzC5UdJ5ig2UJF5s/San8D/wKRFKHcXyO0NDbXJWHJIkLmAtlDQant
BDk5CBRx/mVQ03ctDikm/12xDdLxJhAEwtIMKZU/CRDIJesTFekLjZdy4usZ1Ei7wG+RdkRXDemI
eAC33ivPbYX2hl76uvppwe7ny8yKkcPj7K50IWKZBuBRrhuon3EwrBsVTb/Z3MYn6DqG71Z+FV+W
Bb+aUoDK4Lkowdfh7rjpZxhAAJMn9p1yxDf4QHx80pULtFehtL29DzR4xAI89V2JXj3epRl7DMQL
rVrQo7LrkEpYVWRAfsxl9ndLp5Sq0fXSyNsnIRzQ8KpCz3uyPv2LIhT7MZmXZ9JpZ9/YutaG7kQ+
gdW+BrYh884hnFblhgyBEBuTJx0Ebw8eZleb2pCnYwV8QI3ZcCvVtAV2sWt886Ui0uugsTdbVFC/
77wg5+/FYbmap+W3PlQVO8HE1kClwCTOH68ZKL2MjPDqArWzzkjA4SayVkIWkQHemnjutvYcCZ45
VvFeOD1S7DWn+EVsd/+ToNf/lq2DbeLxGx1mP+KziF4cRvSqQYxLuMQ7eJhTUr07CVKVLdzxO+4X
y5dCO9xw/Xn7MA5Me+zG+ikJdJFiLw1AomDy01DKJ3bA185v3A5GbGJhRQwb/epp1omDwHQpmKzc
9NlZMUD2YxbGIO/99aHh5Y8FbR8PJZ5SO3q34K+L3H7/dD2GWlqWzh+Fo2X9KlVWLuETcK+b00g6
FEBKXYasYI9rN6vUIC/D8LzFenfT0DNylWfhHo/wXnP4wl2lfd6MGpj1U+qXWPBkqEnuOv1qlRNb
CDIvcFZN2BrtnU3lBn7iCdoW/PAaEYtPxgLslAvXP0VIQlJi+p2txjVypzARuFVhIoCrvA8Ycvb6
AcWj2/TQR5lCRJEkzF8EdtjHUr0dpDz6YKyJkoamoN0HYRAJQ2y7jRWze0/vjtPC6ZkaqmLuep/Y
0Zfny2AxxwPQ6sjugl8CXwQCHokHgRWgZJfsfXVdZs8vdHfJZfc4eDCiLLwcpSN4hmm86GUIUAsK
gDRKFGZyamRPCeoCevg3mY/wMzXJjjIJYiwvlQx7fereNJYgy/5dwFu9zneJdhk6DsZM9RGrjwKi
EGzKuKgjVAlkoDXCJ4q06KA4I2yDxqo03zfkHxAjv9bQrSfg6IEOIxWrcTEJRlsLr9ERThstSpAI
qOpkLQRls+UUSb1zA5DpX/gmQelC0RhIv2Vio2NR6dDZ7G5Jg7aD9zT1aLKoe1GG0uaWPKPXa+dm
K/3oVvTqtdnC8JfyySwesY6tGUccAfcvf7CaNyFa/LOAHi55VuiZ4cLlPTiUj0ZfaGRf6933IgvR
ycl5x3Qfb9yBNqypdNuaeY2JRjLATjAkQOlyTWw2EBcLSpcG+K99hK2qf0RYlQQWlOFfV41KHfAR
APOCWBkdVZyyX3WhOdjzahqh1rr3c38s/94OeIjm9fZJbdUgQ4FIXXcByzws1NiycuSB5XULW4c5
taPBJALoofseQQoT6jdoseKYmFUHXvsp3MGnVPJGKPTL6AZKVWRENOnlZPqu+a08rxO3NxoX6iTV
qjmjE9RobHoyL1rG6hfubY/LZhQ00KctLUvD33raRpwkuLy7xMIwv5+EVPJQYXyxVsnhyaNO6C2+
WNgqisj7VYUKdcLoH+FRuSY42/JTLKKf6aaqdC7TazU9uvlQj1i6O/W06MdJqJuFbrjy7mfbqDGn
Cu4o6cz0cloTiN+KIUb3LlRTj+p64PKjGFXBVVoWmbDb39yHpCEURdn6ZckzD7/G8Ynkqumrpp/j
cHQWAZK6rsNVgdGtwN5LjqphClN0bgyGnEHDsTVsROl/h10VS/a84/zKUNxRb7J8oYcs53BB4kOy
gkC/kYjh8T1VTzpP0RjWqwJHN8zpdNZdCV5AKQLqPFdTn7Ej/nE9gLYjmhZaKGgTQKlU3fIV7/xf
GYf+R1sTCY76GMHIUcIf8VYfLSycAIQsFJmeY4oVIZO9hDx8Z3B2YCqKuS60lkBMxwvYm7j5o0uO
rVsbAWG/+pWCvFpl3ozy2xotGx0dKvzB+6h/cWWny6UEtJvteUpJPc4zpY046p2grrmrol3IAxPI
UWhya1/qt+YMVedxVkKE8XnKihcKIrJCUxp50hgepU6mA/0Ds/7Mil6eoiEYF6ikv2cf0DwGtJHP
Nwu7U1a68s2EoRDCSM2pZwcfha2Nn78aSN8dvYngyAX/vzSavqp9lbuXpzGpcvLf6GSZXgAUKkPU
ST1TRlTfKsSXatlZJJMSiEIsSfwOGLdNs8258vnqSlmVEQkkx70u33MysDEj1mAoHEGF+YzsdoDg
b/COjXBNyYj/ySTJ7GjuL+qI1zx3dSxoTCl/2j7StJOBMNpWknVN1mNLX+P+O7DTfbnO0MDhDoSC
GAB/UEQZv3Y+wMHRm4EyhHoIsy57lKTK6lpkxy6PDt6jSGH+j8TocHbETNXkmozHtkzuiDsqllUd
6eUyYSRhxJG2m0gVk55EEguCwoj/BdsryvZEFMM/5ihJybSovTj6Rkcf5KGGxHls1wE9ugkH15Iq
h1znX91sHguluvdIHGvd17U1J+7sbpDpdLuJkLuxkpgjf3O1TsvoA0l7ks6bNCy/LNess38aQh4B
aY8tJxzyRJ55FULHUC8E+PWhYmPfDXvPPF+llBK8jwkreaa/SF/cn+Zs5zjkjR10UjoeA4PxRyyz
/NrCeM48OHN0k7lV/Xf3NvdwZmnSRp5GsTyblwkQlYvmiq8LX0G8y8/fubF1Vz2MlP9NffSrAia6
2Am0TjNzrty+L8l5H49BIj5WDkLQy7O3rjDZ0KSxskjZtRNKdMYxkXn1HkGLOeWQb/ncskM8CPjH
sy71ijN4JwfLnovd2MKeQXcjX9/sONpX5BeqzcUX7xLIuHO8HdrEiCgy1qgwTZDdVyScnWEPNG7s
v2vyEOvOSG3kZLLp3nSaGT7IOam1ODQutmaeJpyf1WfMHhSPX01xOfU1crvBThd//OAWMcRe7G5+
VH5F+OtU6RSETAYtmteFSmTATp0Gip14KGhnSIZp6vsdeXJYUlcqrrf/6+s29Mgxbf2/6eaV+y8t
ndyr//d12L7YeCCb7+AROmWW/pXDLoD5KbymJVvwAhhoNh6oNVXw/kWtDxe3q3Bgg3tDVEOqUkRD
RkVR6+KP0TNnyM0QYBHNhd85Bxn/8fI1AItT2GFtKQMTjjTFtn0lZJ5l/EbHvCXDTyqRx18qc/94
xI7qMigV3ZtP0O6aPBIlVJqoePOmnyL+EP9m+Mie9anMv/if5aSeB3wi0IrE7MauXDqD8fAI/Ysd
D5VotMEKZkuWemOPC+q48gFlkE1Kg2lrlV93M/9l2jY1UBGi1/68e6pjU4tyJE4zNZ8ztI9NmxTg
3WfUVvbx4zNKNiYjFLCDWWOZo+WcHpeGK8H9CQD44TgL4us3mAexA1PfixPBJ3gdNGbUp7HnxqV/
dhNBuslTbtHYsf/LtrCtvUPL+BUeFo8xCTsS7s2NaJ4CpXO82kVs2A91ogNjgTaoAvfbUNo85Hl5
jNuoMjOgpmqiwWOEUWjXZAokIdoKtyHQQL/qagYDyU9Y2Ae6eKLTfVtZD+dzJ/KSZcRrRr/zSRxv
6SKvc1VdHw0JXWfK33bVXTGOj98uDoGzIjvNceVxM1WUFttoo1GgudeVs2Q3YKiZXoSpdvikDQ/g
UkOUA9cjOHWWK1h1UIBPUqERuQZaG+3fZ5FVHV8dpZQVkOqdmV6q5ULajFbB42hgg+VfJJ/IZF5T
LAwnxZX9LtPCwFWcQ5rPQ0/e3TyqXZqRGEKTj+Y+CIFfLtwE9TLtdmVQQKB94J0yONOTXcEf2dth
6WKFbARmTJhYbftsfR8gZCtCjI5bVEKomnmh3d6kBSjBajqfF1n0ssCU82ESX5VNpozKXmJ9sNrU
5g0XlFlmX5x2U0w98Y7VaF06npXVVXR0a4YKhGAW1dp24wkIN+yzoJ5OzqogqXYLjRpEg+d0fGiO
tmWcuCPZDT44Q2dadFaAJYnTU8hg1kaaL7DE4mnca+xYwwJA7y1EPeegWzYgGLh3GEKmgWjS0PzQ
ixvhLB81J+cv0dPsuyf1nVbHf4SiSxtkK/gnQ1t30IvAxk169q1vgBW+CCooWz7uii3y/QjsVnVu
tQuEgS5B/g/KLfbEAetHLkz7zCfDaEhz9kAjJFOkWKOcq+z1ryj7X88Vq+rx9Xj3BGyHXNZOD6j9
lkMgAIVUVqoFRCkES/szXcNOzL/FTRV8LUhZlmDnHGK7YgeIQLAdstVlasDs8ceEDxyQZ+p9uck3
yn8bVubFtMTlSYQgsIi/OyfITzeFBWSSPcWwgyVPVpJ83i8l4vkAZCJlA3XsofT9An6ICA35rD0I
4VXWxNfYbkMXGMXOiyGjT3xOhqsKVhVFQgOVg/vKSMPgTmP04uqC5HRoxquC31oNpDmwIp4JKY1b
xim7Vix+LqjLRAjQfiW3Z3gv6gk1ReDz2EsRjuvAq5duwRURalnflBu30NI1c9FpnRDlsNwBB/dh
0TswqkjHVYSVl1BwjudR3U65zs1LSy1hyGKt4Dkn7MusLJjCqZe+LieAcNI/mcHL+eIhWrk+Cj3f
ketcTb2CUtbYene2mqRM/pAF6atkEj3YSzrdxhLf4Z55qzizFf30CRq12l5zAQgSQLfyMwFB2a8B
7Qf9tPtTauxEiVF9tVbBT6nHXvOqdEBTh7+KCL+fL8DTgdUHMtwebhkBPPzlxjf8YcLyZtEA7T2v
C+6Ygj3SO3ype05W/WcL8fUrGd80uX+jAUUh2IHW/sggvYNw6VudCQU92WK5Rity9ioUvcyYURbI
fR6tOpg7TDzTEJXx+cToLJFhKYkP6GwDlKnwKmUioXszb/UqN4c0811qaCwa7W80gHiFdF4rlVrh
lLDGgDyf2lWfImWMmuSKmPvZUPSc53AXHwUWi26ZQledtbdJiQtTXujqP5zmp6X6iuxZLvw3XHzi
OTY8mSQGbTROXGLN8Sq1wZZBU/dXW6MQh7WZL87I0PKmWIfnVZ7xuWc62CjQ1sI6nn2qOlBAFnxZ
o2GK8TndYrfj8BxzuOUw/zXS7x0CwUqwjC7WpnCuGEx2fWQG1azNS8UvgHTXTO1KfOjcDZQTfsCV
LMSWLTB++83DAOKorj/QdrKrB3e13a1Bro/xyVZf5iYGrA9tu5Oeydkq8kzzrLyjlxhlKHbI+XRz
MNYxDttR/OOaHeAbv8/SvhbjlmoA8mo0Wdwq+xgdbcHPIQP4Px9IgJXzXsvb9lu7b2hupmkivLh2
xkdFVkAE/Mqd2qyEwY4rkmhvDrEbLGfjSMvwnzDoRzXPkfu7suJXFUvdWIZu4eq21JJH05bzgMzk
2tlPi0GAUQZ9ssJ7mhWwUH4tuIHj/gljcgJ+dewMHQGQzeb6tmmQcjhQGUpo7uYpUaVD+Lmrqusc
EP0Ic0bMMVhiZhiGLXx1kOvI/9o7t5nu7FKV7hV7y+UXUm31/nCu9UWj7cNKVfQ+Yf9MA5mfgoHX
Nh0RN4nAWnTfu3T1Ho0qk6ahyx/hA2iWRF2jxLoBm5YFhOBZ8TBbzJvwmipwHDqoigFwxXKNYJsI
1JE7cD1cH7y64KQ1aBnwsTSzEYdgDkdZ0GultW7MdmkX80WFKz8Zu09OkvSZNmkKUEOraXxvo4Sa
J09RqLqONCFdGKyP6PeXoEAo6EIxpLXGyaOyjH+5lZl7O2lRgsLEQAymnBUREorHIYIFiAc6etcK
kCS0WNMk7OnAimv2Icnde+SJikS0eNUasWku9SvNWIJqIkJZ94Ou1PKWsCbIdEshNAzcsoo06gqb
n6UN+7I4mmZG4Yx5xYY/EEXB2LWDDvQ7J+lqHTOVPG1GK403uEz8GA772uWli8kEultjZ2FyykeP
ZHjSnP2pgH8mDNssfzWkFkrqQO8LtN+/XkwYnKVQ8BdQzBkco8K8ZfIrEPx4uLVr/kXdLjtUGL+S
CYgQIiw0PtGvwLBKxon5A6WSTnUyA1lTRFD8fNbZerFsSxVNwifsrIVr1nZWBvmg+iJa24wsu+YD
0ddMX8s1zuoifjuNxYR4S/I9lwiy+mywnbw0b2mwcv9YBqN6CC4K4ESCEbG1DZmrCYuLP5sAD/XO
FSAVXJRnKWan+RdZVPrG34XCURVxajcakVZPqby4lB8hV6j2agnzZSF1i12ApNRn/ZZqQiXbFIxu
H4QJpE3iq7gRt2wzHKsF0W/d9R9A6hFW1yUARtoklIt0nLSoiUIrW/AEJ3tyZ6r5Y6QK/kLmyGS9
1STJhsyfTB5ijw1r+YNwaZ/3yfOmrJ+vb28jGg5BuOWn+zodGifojPpWlGDgrMuJdgRzwcDG/fa+
FFee1P0+g857iR/rFs71WYXKPF95PMQA1Af9L8xA/9UOOVduaD4KOAFOzWoax3+xfz/NJiaQxAX5
wVUJCuRsuwE9n2ugUB/Rv1Ax3Ohog/2qt3IyR5PFsJaK0oOsoUaAnSHIrJoRiEdaUDxPbi/3/bRD
nwU/Tqlwyup9JIh2eGowsk/HUOZJ+psPCejz4Nf8qOndtSR23YlHqrkjK2qBm6/+csoknDwexA5g
ycKU6+o3tD7JH2PTA8Ra2O+jemfB6xSNMsA8QJFhi6P5wy2Gn9PGlbItfSIb9orBBHesfUu02fK2
ECBf63DFoFYsdh8oWMkcAVKsIZuFeCc3S7zbrpejUmd/Q40m7+Y9sVx0rxvOBZtUkoogQztzqKrF
WBR3Qy2cMQJAGlnVHkhFp5PaLlX1H0re70SRkcnnV3DDSYzG3jVsZkXKSumpK8tV4sAyelyG5XUI
KdTyLTZjdO48Y8oxModC6vVf12Grhu2gC4JBeoQ5x2Gl50Yss05VVLHbWkXTjoQ2Y1vLCn9POCGN
pexZ3N39aR6tvAj5azjsbQN3Wa5X3FxFkR+Nye1Nk8OuUIWOXMHTiuIc87wOxtw5AT2F/Fw3HhjN
M2c0oXcGGS00MDusbikZVnjFF4G3Uwgij3Bl8rdJrijOB6WIcDsmhqNylUDtJS6tia6HF7z1yr39
2PV/yAqUagLGYz6/E6VHuWTI30tk7nffdvzxJyLMmwBF6D5jwpIlUOK5GMiazDLNyOdI6kOGGVT2
a2/OvUrUSaDlUyOT8F+FLiFM+BWiA90lAiaPmfCZfpFtA0MyJGU6GvKrazPPKOFn8wAKxFnBr8jL
P+i8HUJJemxmUlXFuuWR1Vd4LYayOaISih9FXWj0jWWanMCsvyty6JFNUMio0EHq0WMV+i5YwjT4
Kfxqjt5BLEyLQ28XI9pKFNm1S8dSSbEjHyGPXcG8hA4XqmujUrcMN3SGUjoLdA90bDaumwiD7xsD
qDyQTmx8fFdJSSDSKT9sScvScO0AKltsxcH1/9L4kap3yuQD1jmyZgeJo6tyc6bBnz5dqhZGA6UL
CTPMLNDeg+gGahwhFGnlyaOSBB6OjJN/sDYs6WvG4GmUAxDYM6u/UZNrLA15lIvJAt+xDJxeRTiq
kzvNv221gCfqudouY1L8T0xSRLOX9TdyfWnTX/HKfF3NkCxJBge9CsgTqJ3Ls/yd/6pjCjALL3Ky
sC+jPjaqQ2cn+FTS+TxDT/fGsTHmGDZvdJ2FNFZCDmWVsW6TpwkQJnQwijuDDEK1gvNhyLbmZtNk
VjGoCTwQJ8BHBJpoQbNpnwvBcA6T5q2fWgQq42yA/CBHlaiNeOhFj788aCmEHKF3Eo1Oif6yVf5Z
IVN7uBn0wsyUD/dvcQqlTez9NhqR/NKs+3O8Fe1s5Kz243pl2oLM30PBpxJ2JcShTqmao41wW6/k
CKnscjdHTPZGnh/YJdW4wEI+Jm4+2cDNK6mpJo+k0NgRaV79yBPXtcCzQ2Grf8NFuWRMCNNCjKD8
cNcbZcYGZjlrBSrWlQMO1BgoSbJedjjO4z0eUIg5x/0pm8D58UdH6Ga2D99LcnN/7c9007C7olz3
32yu25X7RKbx0zPJUttlbot7799DcLzGajkz2OMBqVasgpmlX2v2745wcKLJudJj2wwf2nfE1llK
RC1n6X//JBttXNI8CWeuE/yFn5cXTF6yBAyJDHbwKIucYqBKJ6wd4qTOO5x8gB61imlj4CtD/7G9
r2l+x+NoFsEQ4eMao4y1Jjtzl2aGxk8aatMMXSNJ23I9xFsLQgmz02TjRvMq660fI0Fa5cXSgAwK
HVgcw4rS8C3E2+ojwnv+KkyzMolSxl9+6wYryEIK+J4F+xCdxCU22bXYvvhn9VVHagf+jzPlHDsF
8dLm3ZKH3MBTCVqRscDJfLyPkMhqd+uaW07S5rpnWLGXpxHHDk2zCP92xdHTqb+HAeNRgu/5uD8o
xD73VaLc+rDfAIDI/7fj1zc2fLGrTEBMoIah7jLOzJyGvI9xfAJodRMGebejGMNXtHciAzEAWRHI
XxK5op+Ncj9AqK/xDs9b14gWSDhS4LT5zMmxv+oRE8rqLLlOOEXHG/2jJr0O5o/bxl7AphpjYdYQ
9qVup3mMBxyP7dcXPECYpyDrvdqKKYSVG+yIRKqlCGoriGx3Gd0PQ2WJY3soeOGkZRG3OTyY1Rme
6EiXkwzVFHG/kaQ8n8vBS58LV5eFSh8NNsy4OmrnuoUnUQkO6B3g8BUM3xbU3+EpvGTRGifcMFiy
rOkHzgESAp6XtlVV2rWrzDosvaWEnXi0nS7J6Z0mtIqES3cXXolDpjLw725v+ms0viUDSw7rbs39
cL8MJWjIquF4QwP4E0spYrCBkO0SDoSvO+OAv+GJnzobSj/Mg8hiUMDRzttG89NhrMQ08UKnGa41
+wNP8QZt+GClAdu1Tov5bA9RrnJ1G9XTcw22iDsxSI8R+guuxDTn5kbj/tHUBSXW6jRzgZiAbVmH
K/GwSw+pxejQcFBxYCcgoTIKUy95H5KLm1NXk8kRQnn7UTZpaHVzzVCrhOutsiR+M32rkATR7l+F
1fCnsOB3ZqBMb5iHGHXi4LvrGEoOYmybyp8JkK75D3+WSTc1n40XlYK1+C8EHgiIndzQeujS7SGX
oJB5ZEch4APsUAI08hoEnA20HClEeUqWOkKMCfqaERMSUH/ziBik0I+/PvKOl80sLPvm/6ubAwF/
wBsbjXKM1QVKbrJTL31Xd04VZJMZ6OxUgUhrrtI8/eKkv9mGp+LetwjXPFmU3e7LNMuQD0nXW478
1JdLYz99AKrLENGJ30OkNthwhLbumD8tuLBg9/4oqXMyPFuSyCvCXbbK4mBfPaEyJFS6wQu95QEu
vsPSVqakyDZbwAZQKOT0Ov73LbKMUExcSNiwQ42S/9nBok4ghY2C6kLraiiYKhJuG5fHnDGS9LU7
ktTcBzwgAwUCzFZ1QaUBEBLzlZpOJ6nfLfyBDDu5aYe7uBuNzhK3oxoUMDCGXLJFkVQbg0DJHEoR
TYUxphQsIONlNXy9inwlc0ZEsLDyhyBYr94EdcO440s0pH7/fhv3IW1fqZKcBgxUfUJmm2ouv2Cm
NLmo+Sk0W0oisdJpQEhginZMyCl04yJZ6YmYw5ulnaiSQ8JEo3Ibx+p6BJ+iz6WhmssXrtiNYnbB
txGCsh2BoRBJHU4G8EnzOyP1ZOf1iIpJK54wW2UaJgiGOYMaLkqtdRJPqhZqPBMQGQU95enDkHzs
SAbo3kWi6EjcjybxRKKlW9k4vp1Qpt+NMNInkgd0K78ef3pMyDexdPIWKG3jku03AapDxHHg1sZI
CqW2WhNbSTuRgZwIK/5W5cPgo9fti631P3WC4fS9lqcJ/dXTKx3qRGBhJK0cSIoWai2pkqs+VlER
OYUraFG9cJ/VqZ2DepguwGqJpen11JwtviTT7tLlTSD3pctj/bpDdXyTylNEGr3949pWNXZsVwxW
MrCric1qjr7wK7EymUgiT/VQCyJo/EhZ8iE9cySb2uqRuJeky4H8SVWFfc1h2gtWk8Ff8lZSumb1
f5A/tKmPkBcnzQvqX2d4FsdBas9Ocokxvxi0Q5KERNegJdiEZPsgjDHMl1QHb2RKCeLXxhadD+CH
O+XSb4ZQGK7PZq0Hh5B8SpqnR+5mcgRLuzEAIpEkgLjwrL4KkiB8hq2XOe56568ly6C0aRJBOQ1S
R2XAW+kw7YmnM1qk9/77EYqkPkCtYheQ3p+2jBsQtfMh4yla/gHHa+GaXsSyr8FzU/Uyh0zhhWVI
KN4TvKE8RYq3Yqkj4Q+64ntbb/3ePYFnwxy4G1Vm/IHaZmgVlVz3wiSgpiQ9ydS2o6tM498rL/51
74/jHwhQxYSR5yL/o6W5KnYYDBGk1jJcbCo5EuAYvO/m17h21eqFklODDggQf4E2HjlauUrYinxZ
0pvznFLvRVSIMolNNxmUVoCRGL5Xp96yEXwQckkapYJX8rrDi57mykequxSYf7B+xyppw5+XkHC1
K/rWubPLAKQtrO+1noyrga93mM5OQ5zNQZIKZRCAylXMMIyM6df9kW0hFmBZx+jTcrh9i0jSuWIA
9WbiYKdH3tf+5BdOo4c6FkI2G3ITRAAw9aXrdtixkgDQvU7OC1gPNURJext5rHJAOjpHTaN2y3FQ
sCeY487tl7RNqmDYYfOmUDFaXYsk1JjsuV2jQJfLEwfCYgmDmduocd4hZkaGqpZPUD38a8IbVN6j
PzehjQdvDFa5oiSdPnzWQucDDvhfNTXCX92GPB7GZOyvX30HbnPNFOjU4ek3SAwnyxTrBJVqjxx5
a+h082qMsDBOVwQBmoWm+2fMqg7aM2KSzBSIXIxVrTB7HqSnv8yAHv5M+gMPAQuPX73PvSR5z+35
uYnyUkR5V1GutsnJMuP8E3zN+2DKwC8Us6n8eD1gVZew3h3YTnvlE05QlAkVgH5PL/atRqRkxg4G
8sihMGDhmSMC6gsZ1laqRwob7uLbujlCu+2xdwSYzQ/XGpQvYR1Um/OViWrUtm3PcWQI+EyGmqfj
b+gz12/WsHLKDEQAdHLYp6PiNiphJzK2dDJV7vkAI05OK/Ue2MUB2gegJUXJYR07d68eClD607mX
uwrMsOTIq07+MWxeEEXVW/VE8+ACnLxL35OJNYf74wlJRS8oQ6QEVLxAytaCWQPZ0XqVXh09Fb1H
otiRVH8F7eqz8h+yv8WWW+KhdTEgVQQEkIDqp6uLwjzep7o4ea6yDD1JnZVq3mWfg2V42xrozmNN
TPeaQ+9Mpj/rJSFSWjQeYf9iLvxPkOQ3jIocgb3LTQpzWgvPP0xXIPO3HqY2zVcLEyxmJwrkZGYP
iVfM3jaVixtHz/CY7ph/f+Iy0gZSbBSBPlN0eBh8bXqZhrFSUfso/DFvclDHcQQ2Nv4yv7ly2D2A
MYJ5usP0zJU7Ct3+ZeiQilqPxQhmnUHGbu6g76Qt19K8V85qH8+FYHvVW5qp4Iv1AYrT8ro3xBTm
Mb4Rpg+GjEQ0Hq6Eouvy81tV/AEUzTKyyaBp+y/y+qfHnogXQAIl7brwq/kUhbRXcVwEiC5tlNqL
A2mCyKrqqhJSBeucQ+yjbmkNWXhvIMTG3D26zDc+lE7+0AAes58g2Fo+feL4F77QfDINq5S01IqH
liWk5G6iDynVl034oGuTytS4wiY6uv0Z79t7/rKKmDeZ5EzML2wnlS4zPNIGP90SbEWLM3GKjVig
W/9iazKMCPzOnHzELLucTdHjs8I8K+zZ4YnPdWN4Hu9ujsQfOLsOX1XiVMDIp/oDdESMtXbWoLKo
BLDEGqUIcRlcZo9NkJTiq0OGRopDhVGlug4eJp/AjFZeoe1tl15L4Tljp7u+XZ21QKBPWpi2MRbp
Q1NA3ZOsyvaPGUyGcaBqeUFLUI/Lz27VbdXNg649so9dZftp+nAVq81y6At3IOOY7STX0REMXDV8
6jE2zlBKPwlwgFw/XFyExlLYTWGN5D328Xn2OvnvpHaJ7VXjWCRYYDnFhVkSFrNeWTcmGozgFvP2
obVZDmycpuAAg81wC2ri3ScWBOI2JUihBrOfiuKvw4+jJlo+kWLCxhGJGhKMcbrVn5r11sLhEDIv
TlC2DvsEbaGQxC+wLP2eiXId6umcD8e018A72cdx+Mp7RkeHKJEMGKi/Je9UyeqFRnAwbKpPnrbE
wqcOlezPNhkCxNyVnFRcUWfgK/POvCSI3xeoVuL4Lov/rvYtuwPtWJZmqQYoe77R7Xam6VCFXBEp
Lma4kRWC6SUN44NasPCCto8bNIMTHXwrsqx+f3jerRDpdeU3zsfijqSKmd94w8JgX9ClFdVEN6r5
UEKEaiWFUud1di/FMoRG2Dqx5QgajpElNoYpRmknRmDOoJXXbf7qiOUW7pH5qKUeSlIpZKd6ojtH
Uc3BmazBqPhoeKErXJKkSaXvvpD29Uam+et4vvo/6ZefLzFsJ+wJCu1XBzc6RWiNmxgWRxWxpx5C
oFgiz/qLRf683I0XvSQk+wE1kyNw57ejQ5AjkBivxV4ULELVtNYB9GUvU1cNfrtXD5rU+jfZK8m4
+Sa8FqE1ACaYdvAz0prd25uKgS38wMtx/OubRG0w+bau5gmbXXbQIsH1zmCXcX022QD/+ulBuMw9
3ak/ZAMZ2nBn1SaRQKX2sR6VNS87zXCn5+JP8PsLFm1EXA5xZxaN81S4gzDCNULymPKSbmRj4Ex9
40rRLYxgeH536bS6XabdHeMulvyMwvtkc2Ure4vOIN71fhYl2cFZviI6uP88p1J1cDdEuyMaH6z+
uJXmC88/8bBGfm7Pcf5Zk+Cs5MzH4Rtong1AO6UtVwi6is4Vd32BXopeA7wYs/RlPabRgFhWgxK3
M+WEt+bITCdmnvssGH7EiAkEP4jAsO0T48ZWiKQfbV2i/g64bFOU8zDgI4LtKU8BQ7DqvRo4oD8s
76XgcJO1d2QIJNOZu979HN4vNHqSvJ7W/uRZXuXlp5vkhCIY9LEoau79/c4rVmrJPAfykIkId7/W
+oSLS6fSk6HG8yZc154FjS6s1QQwkN8souvMQmv4SgsrIH/cyvoPlh1GvRDnjO0qQljAbDsQnbe7
L20Z4mxLGPdGXlsjBxJfEHEA88YK6eXIenD+vMwnKT5WS90bjdDNo5WCwcx4ojDrQThmzxxZqQxQ
IjO/5vg5IUngxK/HeqcR9Tu17i7A0B1dehhl6deC0H1DXdSysuY49leyTLY+5jzPWuH2GgTjnEXg
Oc+yFyY+wYzZJPN+V6kgjGowtqyy2VF0PpnFOmelBi2qgLiS7+g7eLyUUuzRwzncQeaidXocPxIc
YAvt7b5/GVyAGYhE9wOH4KVtuNNp3h3oIWrGZWxLWHYtVFAZe+Q3qC5ZQUjrDD2H6TWwAIEfjyRh
M0VWI3mSUS0RfJpmzcnHG7MemfALaETuB5ekSi+2y6MUoDfKqz9X2du4KLioKBHuCZ+UTAb1XMuO
RA7wevdVM3H1wmJlWCPtzis/n91JSMy7KJdwPFQ+hd8XmDzc4UUeZQX849ndsfRLmBBV+VdGsw0U
RpKB2fw/fJfD6PulDCLfoCugINNX3jWLyGxlQy3/dvRuqaE5xr877ICb881kiP4u6RrAi68zfatu
iWdM25CaLIwIt8WEeeYSkwN0WaoyuTby4GpRSvwDNc2RRzs6BclnBassIHGM/Gom4DYVloVX3KL/
TUNuzH8XSF1wzD/U72xRO8csfzuGG5oXFsXwTMenSJJafsXcncNaG+6a5NeN7LpI/76G/7Aqnmrn
IxA0+i2nEWhEgITNIfwNNjXYnCWTPfGa0rWyvtZxDU+bKW5lPJcKqQhBNYWRKuLN/rgnXdHSK4E+
+yEP11LJ4Hsh3xYV78ajnYy6o4/5lATyR2ayML8h5DsRYvwI0MS5ZCQfZJb6D3L1m+ZEWtx+smRB
S9QkDBZyInNN6SkQR0SINbJAQcwFRS1yl89sS6ZWgqPFwL3Nxb7zFcwDZOnVXNRasG9fRGP/HrH1
46e7+qbSDu1LdpT9o3NH0ypCC5U1YEHm6XiWjATXCsr3jaMYJFHNDlZJkai00T6NImxkTidfxh6+
0qbY9Xjcz2aEYF/rQSRmv025VYIecMfCFLYd+KasHRcUeY82/ydWWFQmqoxZm4SzAgnX/Q3OyBm8
30maWNchYpdK6WKCq7o0W1JkuLsNgSpfaVE7EEdGN6rrKBoRFHOz6IRoyq28K/iwyHPwNkL4wkbL
mOwlAauR+G3tOzxKfHfBFNzd1alXPoDsbqITak3EBwZR7Ki/l2CBRNlpzY3cg4MitEOiW4tnp37N
kBnjx9rMGmhWTkU0DMWIe5NFBUrn9WaNSuwzbHlANSC707HN/7tlIqDHLwHOFBiKc339OKjg+S7Q
Le81k9QrmeP7FgpzJigFqmcfknIYfyWpxRkJnOoddDx7Jt/HOnZ5yI/kJ7uLPtMeZHt0y4/cDow4
zWRZ9xjKmG0LKUs53ybQMZ/6LppAYY9fil5UkO2v4ZKx0Z9qveUvKdsNCMPEjn5ErBrPUhURyw6l
W5css/tQobhFDRF3bx0qmoX0MqYKivosFNUWkD4OwR1cDtEqd9/z2uXdkDoMbAZ6mCH6+PrW+oFm
3Jelyxh1KTiArkTtUMR2xeK8Y6bqL7qXRI+knsrcM1lhcP4sqWkDPq3WMrrc6ol59iiEzIJxI878
Q8xAJ/nTXdf9A8Yt4pHNytJ4rXcD5w/OlHGlnlQK74d0HEH2RrvrmM0yVi1yTpEGtf27WBm3PaeW
B9tR4hiEcEKlPToYsAeVJV3XAmmG1kO4JDoqByDXu7+rroINE7sBvckre6kAHFyqlpa+m6UZ6nbt
XKJqH9+tvlURq8lJXCRhCmRg8MDNkKlPFodLjNFGyrAeAgn26Q+aklAXrWUG2/u6ML7i6FCjWe/E
zJaAehvIISum67IRlVD9FqQagoj/7HjUm2uWkcgQT3vRUcBaJcPlbOJnku1IOoBb9lQ/HF/Wi1C7
mf1prdmBBsf6tYBSHVdVJhA+ccxLYMdKHWQZytR9M/XwnjBcZqQbtYxeuv/8GApqEDn7vGScop5R
XIbHMKB2KxWNSErNNeBW6DBkX4ItQDTsP68hfHOGw+bvXbSAj0ioLDxUuml78J8UCmIja8HPTwAJ
05aRLN18LvXIBfKf/un8fMdxg1uaNhdTwcWFpBgU7CtMYNixjcwDFLZDINJaxxGlGiuI/a/gIpLq
AzPFvzak6/rZ6w550bbjqkAtS6Sx7bQ7OHj8M3VJx35/HOB1q2zf0kURGmlVVOcj87nRZvvXhvzw
V/wuJDPFhlTjaoEoCTUMa/p5ecA1ltQzkKsxNGkbPJhr1u7zT9mncahMRs1KuDNNjIcj80iGuvVl
1hiScUbEA3EazqAX0iSHmA1aGbnZtHqkUWVR53k7+Ie5LLKkJvcR9XnBJ2FOg5duWcNdKxUhf9iv
hk3llKBaJ4IMPgBbmG0abuf6kXX0moNnViXAft+ByNU7+2YZJ1F9ZoW3wBIExzJFHxbECREIXIRC
2g0iSaPJvqsi3JYX7xQaV1NZ2Wjymbv4iyTVFqzFWgVjUoQZt3MBNOHBFFjywbbpi7KTT2K4X8NI
NbI8I9XyBlgnLm0fqSlQpqFDQHnyTI+PBXOh4RFtL13pdpJl09f+wbojp92lofkqswfhuakYg6yA
ZMbu3beY6w4pj+fDhGUtbqMu2uL+eZKSYRwPb3MTPDSb6L6AYObWAZjypzAr3KjylNCYK3td08HO
6jXpeXlLULKZ+4L51LeCWtvwBYVxgc8rl2gvxE1HM6tDinYS+0FmdI5BRc+OIEyKebEl9It0Pibm
NwVlycfitOSAkIo2yxCqRBPrdEsrqNhlE+rbd3gy1Q1B7j9P8E6VkfxPbULK534Rj2mmhqrlRjaw
LtUOLe6ezTjkLTEFIKx4C4mAwgVNpvQfGd42DrfWAYK7XnD5/aHOMRiDg32GGQ5IJnA9bWMdphP4
qAuZpdmSVPuZtbROol+WQQLrnWDuBpwfw6qFuAeLt3KGOekll8c6MAH4zT7fzya0y6mXD9r45oYA
mQvBwcqu3Cd/0+yDdjwRdKsSsQKgqIrrI12XcSo2BsIBItWb50Nn1lEr3ssq8nhAPT1mTqheJCHy
5k5+UndgGrJ3SR90aTDzqAt4wbvDYbrMJK3TPMtxQ5TLdDxUOlAymdTGAmJ0+MImJZOZ0c7Qsk/k
2yfVkoyY9mMcHtWdoWAoV0B8llOSa2AuxS5pi9ufYeoQSRNaURGezyKwy22qBhcaZ41mEtx50dg9
U4yTX7eIfQB0o/f2KDaXgU8E3zLy37d94aHd8eb7v03BO2pLxSfMfLqPy3lD6TRlQia+MGc0uc9I
DxM8GW+FmyMwh7tVqWQKJm4ir+myguZYgnFF8+6e4HS6U6uZ+YvIi3v2nexgZq3f/p/d5J8LIO5Y
Njc9M3kOl37LC2hjDYSHQ1iwGkjweJm2QZXh+faI+xHcy08YWY8WmL0YT72EAf1LHzfHH0E4I3Zb
v8SuM5mOL/v20M2c8+IwxR07eV2f3fCdOC81OkmwyVkGp/1rAEyAyXMNWzhB0uIWX+lNRhgLwhRk
3pJ4S4pFsci6HdvnO+TY8m2DgTtDBpUGEA+Wq0uyxTr7JObqT/9WSdm9uJfy24KywuKNcZY17EiG
RXwN8gPZep2g9aZs4C2HZzXY6KqYhywLeUGr1khBNkJtH6gAUiHecR5i1tpFAbXF9fCzt5qVAITM
Hf2q4YdxyvdVSJ1hT77lb0rnraGdM0awPI9VLymoY7UcBp8zho1cB6+rS5jB900avpwIg1Jr9Aw3
r2cUpYJv5sAbQmUyfbhkEpczzzTep/i8fz9z0+4SDQWBC7ZrsJsLIMsgKwYZFhrJuDioU6AK7XzP
2q57AzJJJWDB4WxrQzJ7h3oCxHy4T4UTeC7ntgf3Mhj8BOXWxk/l7rcB8OFP5kTofWTP4kiGtS2k
FqtAWqzMWdazYjl7auHNyLj0oyMJ8C6NFGRE1B+4WrMWDfVtJp2CkdSz9kqrNz1IsE/t4kQB+koY
SLwloKfZj5ThHxm4t853G0+Y9fydPRKDwU4OPyZkWmYdrJOvgcLakWe0ciXXaLxUo84XEWUf/Jkd
Gzqk7dVp+6TXMvIVdxWkhoEnc9nA/om92EVI7+Ja8zLxellpTWOegdkB6nxR796Xhk9zQthdn7hh
kE+bBxl4e5dADWLOJWEWi9GlBmUAfGDxeSgKGI6qfSJbKEc7/SS2OwykLrnAXEjgHZrvcO3be8Sj
IUX730p0Kk9vm90peWwEzA4I6om1LzGkmDaHVFZh87WW1L24I9hiOxcwM1gP6GPXXIEOq3nTxkkk
b45OsdqUhiKIkAwXC0xGNlP2rbK82V/aPNHdZrLp21J6Docj5AsKyPyx1R3f1qnkbyL8w80rizns
p7bhfs9p8Z0kIa2RSMWdKrMPQvMSRjtfDruLsTOvcBe2DVt/px/jRe9X3/I/c0d00PgPJ/w90Vlp
30uOH2bAghjv3uyf55kLsT7GxgRe9qfBmdtJ8dFKGx12QSbvqD5VhE3PYBI/7MJOGVw5GsLOdQ3u
ZYylFDVMsGOjec3z7hS/5Vn1zgTFy2PskLSPMc8d9zWWIcpP/9esaMlFlJKjaxAD8BWUcJ/VfA0Z
XMoL2sS0VmXK+ny4pjd/4FI7I6XNu2HfOh3mMvfu9aqCPE5xS3ZhToxAcjn9IMnd//X62xqF4TNf
ioU43P22BIQqGNQsxnI8/Jh5KSROFU7f91GsyO/JwSBsQqVch4+s26N5qXDK+z5zowjza1kT0MuB
jXPmf0J8SBUfbAxYW7H2FL8Sp9o+Gv6D5YXGRK3r0wHD5EkokZVKjWDmSGH/tY+e/YRwEHVhsHMg
cX4a20wAf+kjEabLr4vAT6b/cz7V+tIiCI1f6RDdQMiPKpLUEFi/R+JJqO1qTpPIOpgGCAvJuuRi
TGs4W+A237DLL8rskN1qobJLvhL+l6HXIWt0562n3VnMsabvuw/yytEXazhTeJhor5H0hxigakcF
gWW8bkShTKTfMKepTJfRLP4YTlJZmnKnGRUJwn2rykvKzIy0dZNKwQUxerOIRO5TfGh3mNQB7cM9
VEKqcDSB1iLQCozuZbJeL1UFxRqtAwLgzuc2+EWc8YWnjqmJVV/Y7gSDVT3S9Lk0H6oZ/Ch78Qpn
dEFXGWiF6RkahtoaB7RUKsSo1BPCQ8nsQVZdRFS3+q++tvArr9x6zLQepN5KA+zHfw/xY+ov0Iuv
2wsXpdhtJDZWg0OSKlX+c5geBOp8Mc4uGeuIpN44y3PUM2z+RDGgcx+l3uxUu34AdKEKf2UgSdcs
LUMEArpCJ8Z3g/KciAprbhHjORhwwwHyj+tDYglJs8QYsoyVvrp+wSsI6UGnGYr0UIHy4fgxtTaT
c7NpMade4Ruo7zAync2Car7m7b9+CLmBFHgaDep2nWCJMfYrN+Fovo2x6vxFsaJyRBBbxP8ZZyYP
HI3XdRji4QfN2ahlsLCfFa9Jt7E/6fLxxMP7GN518BrBupbRD9dmLqAomFvdgbtb5vizkA1D5pbq
SSureSHzhHQ90Fu9ltm+wiYFU/DoAsjG2lg7Y7zA93XCXpOkglWUlcs5w019A2viCk5CKlzcV9NK
d0YLDWBTwQ2ibKps48FzUp2ZJ++7gZNM0NdiIz6GuuBo7bmF/FRgQug3WcK2PqNRRViUXE2Fvl38
nszzIwesSEXy/nInEaTrGdZN/kjAksQKMYRRGAdIigAQaNupIF8TSeCIf9VhGXYdQfO49unXABO7
NsEelKTrk662fyspDJAI5piaEuAMwf27KnC1DeLHy+jBOHpbNTG/Mml7Awm72phzGkqFupzEMDcG
88penwHsKocajDNHhHjFeDFDZetxYxDNNC0Fdjm7TVA/T5Jt4OcR/9MJhHAE+I1WwWrV56O6RluY
N1kPgmgi/va8SmO7MsQ23UBD4SwEdHoslITIBQWl7VW/18+yVASvwSdkwymPGaLemRGDQSf1Aj+P
IT8xini361ksTHuFVKGIgTSMZ/qUaI7jF02TKSaohu2V6kiMno1XG+rGub3ZIoager/+OB9N/+p+
NFGErFz3fVFFNvEzJhUsAQgP+U74YT0MjR9W8f0hMS33XM64t5t4wC9R9EGe1J0GEmVydJfJJDvr
tLvCfqEUywP914RKBVL0ABDyOusrUiAHcvYnunfDeCHyA0G7VHq9k1d8wNQ9kEmQOXKVDv+tZhli
5d5pFVc3yfo4B4yxDvfEWQR6z24huj0ELqaRCot831wf+TyVTYqRu3gPTYpHNFqhp1KoEHzCHPcS
3Hck6SvOqKegs4DO+7N2/fpLWGQ8YvnUJoDocCCeLcxS7l9xWQhQaPPwSkziwvDsQy5J8gcQQYkb
dlCWJsooFjq7kDbfV9Wr9tJllSBRS1bJRNT39sFs9KnHp/TP9lxDcAkxEqKPhieanVvsLVbShnsq
pK9RJkhS9/IW19omhXlevGQcCTrHhMZNgqhNjsz3rauZg7B9nyxyx5DReLItEoPNQqnchb4A2a6x
3fxRjZMNNoLd8nlZFPymFcWskYnB5jPJYH8Hpy1CbFmiyOYEK+K8KZFTTw2uOrVOxC6hj8IDlVCa
OXIvIAK6k/UJIj/ZOiyFkpu9qrKPnk84szFnyawHIWMVChUOMScUudnzUngNV+XKkAoDj9q9jSUi
7/X5Lq1UzDfblG6ryR5k5mUMeDs1RB9LGheqyu2UJ15byWthIleKufJJ9DPRD9PMz2nQXcgdQD8M
A/HggV7/gFVG+OWB7El/Yx9/B2i67kSoVcvWIzK0p6+wLrBYDP8vr3X+Cpq6EO3YW7Eshuhxm2YZ
2btkaLlRSbqt6bOyd69FcvGJoIMK/bigbR0Atxi3IVaT8lrHsqeFXxa2y8nwPjY1tqCCKbIsUloL
4OzxFsahsQ7TzwWoa9b7o290JdDVtXhZxKyzav9lqS+cMNN4uqOsFXUql1JZi/LQZM3XfPg0IJYc
XNkr+vSmVOR+x/JFcwq1yyCv7gq9NUImIWyAm6Mah9RGBVCypgkcRWebgxB21qZOJANEU4q02I5x
p9nlg+K5JCHRloEDHX7bhokNB1PAGp9dM1fzIDNjME07W3VYPni1ktPq0M9itKfvOlA6GFPTits+
oF6X1fbjZxNFyv4ru6Jn2b8yYH90Vcc5jRyf4HisAr4H815RRy6LvMgUsr7lKol1DFmRpQ6lm805
3qX3Rg3HsmQUtm2jb5TFMXfS9b8I36dg9mRL9c9oPnaIkeNSC4M6wLdObHc46/RlpduURgaSjwq2
wyz1ZMAELFUB2FCH+frtfcMYEDQN8X95375KVxliG6ZkI0FxHnzs2TppbVQPMLNyguFdEjQFJCuI
6cCcz864ySdfmGfRR7A1aQmRJnq7HgirElRJPdguFYNMfGgxitNIMB92UBjelUUQxBL1obNoCEbB
iD0DmaAtk82Xp2rNjEFpZkXxpIWi1D6NVnxLfFLZ8R5c11us0PJwqpa8NF87JawZ++HZAbjJTzr+
GBcst+O9j521Y/KWjgLZbx/0lUov12KHle1wOI1b8HJEbWb6j/mkybn825P3WensL3aws1EEtKnL
nZFvJtQV7JF58BkTmWwBRtABG3lXK5yu1AnEX8OEYmdj2GPcHpQYyfpCgiMzVEszIV48M2Nl3MUn
Oh0mfiLrbaU9RVmNrbCouzgKzYy8udm0pmUTH3i7ZxCBJ3Q4EySLL8XyjN5SrwokLlJc2GuyqEwb
f3ACRIzEUTtDrjonytmKVz9Ox+1XOWCMUDKuMU1ueZcMzTAh/zdgxos6KqIAA7DI/CtZHT5KBFaY
PfI9y7NCAyr7Z1fYR4vl+UKBG6ehtM9YEoJ3zZtrl3bwuJv9cgvqITFLWHFWovyPIzzfO4BGskO/
7E7UyUuPPu2+NkSqdDfp8zvSMp8cpKkOKYzpruAkra6FRkkolT44XY/3X61rWgGFR2FbWwD60TXO
6oIsmx8UcdYc18aWkuTH3PdTXmdOm4zlQsaMAmTfF9RlbM8fDI2Qil6E0qd5e/glczKb0oi3tCVb
FIsrSphayEVqjZF46S0gwQsdv/tFUphgxkl366ZpPBSjERBwzZ5k8KzK5ObHFNqZKP088ujg7dhj
NWgVeCHkYhlMVHaPfLCAW5i8UaO8HfQuZt9+ZTiaas8Z7I/D/DKawsH1aSW9/6yiyGOW1j2unBHk
LDgfTyWw9ya3rXmkF0Z+O5fgC5iVuETasS2h3x0dvL1LXR2xBKgTi+bZdb9snJzoWH0TKeioU4d3
Q7QJc72vEKu/ouSsPtTwf9yt3+jOCsOwfaiYDZ1LMBogjr5D9bDham4TQIVnfuhLhPSWDGCpN0GL
wlJsx9Ab5eCdrBIFAiyb1PsPSXIkH81c+DFwsaXO6lXuOkRWX3im11nBBpas87dYHF3HVepTQk54
Ks3Dlsyc/Bj9Y6DzTb1vwB4emDa1MIsSVtiuvWRDmM7OtCIisX3qB4H8Rv7EfAfKO0GTM8ruJNEZ
IKV3/NDQOM6//2DIZ9P8EsviZqMdfT0LyQaloWIEus4YN+nVwjgrKP6kclxOKlKxRJORs6H5/ENQ
ZgBZD8fzX6uvoHw022UKgmFSDHatoTPJMLbjay9wO/hEFJ9pJXhe5n6iUAILYenyIsTSrPEs5nlg
1ex5QOyl9uBvrO6SczXkQBfwIv9gceyxXLujG6dcP+zXp2VV3Q9Tj1KnDWJRAhhrXjI/1S+G75px
Hj3EugU2D7TYvtpt3cUgXhnMO9gh5HFYE4oTwzeE73YdUAPNI2R7xblIhNOQUOZjH3e6F4QJf0dM
FUJGRKyoXxaYZQlkrhFEKI2JIa4g5zNwWfiVfd8IPAh+QVbTYdiI/Z1x6CqITqkLYfnga0+oWV7y
gWaZyRxM9OQEOhjM2Fs8TToTJWiI/Fz9gjmN/8GKF7o9zGLf7VriI2JKz4jJDxwCenJxIezfodks
A0vCMBufWLLVEj0Drk3n5JrXRJEdfI2OZjUIME3xSpV6iKtqfDjm+9JoAZYOqaDAKBGLjUMizJrp
HK3nR3+rqiJpHU2YSzsVsPjr4XKiW40cRrhIy7CK7M87a0MzoXFoMK7HThSr9+rmfZIejnK7lNRk
DcbmC+Wqn1i0rcRDpQua6WNCcmsXXdhZktfzQv8M1jtirASSvmvLEdmsFMaNsDVauq1+ZmDZtbVt
F+C8G8SzH2mEiJnS/ee1YRqY5IzeFMGkDbIcrfm0QUc3j3TOqhS+jCmGhdQ1U1ODzzL3S4R+639Y
YTuPjU7+yJT9gQH6yp3tKXQNbvY7+Utm3RHTeA2zMQCyBcVi/5dTKOQ4wkyz2KcxncLgmGZs03q6
QyRrlqFD33Oc3lI2xrCGf4ci8OQ6zOrGrgQ3I++I/mSNTepEeRgPjic/stu1BetkY/y26H5BxvCh
KQm0fgyWtHZ0jQ4gP8udpDdrhYe195n/yYVhPJ8dHD/jWnLWLvOL7HeZ9txSOUusT8eUJdZ/dgjF
HA4IJOXZ02jIilcYkAYQ7u83UYRWsPMht3jWW24W0mYKbYzMRiTO25amTdPymY1a7WyPQM+zwims
bDXUrWPNG37NLCRsm6dzIG9z8dGtsCsFt8nD455Eyook2EtpBcFYWiiGmrgMvAd3Fdft0P+3zuKb
6Q7QEy63kSnzylzydEzBhbUCa7R1+2YBk7Yq/b6diuF4uI0rkH7LYEiNpyUi1lxQPoMeOzqFmmKD
5rpSDGM84cyjy3c7Jzqs4saEL898yYlE5CIQAtGgY287+acNB54n8A03iBhmhfm3k/aXQftJQmW8
zXNpxXHZWL0OIq+uY0Ky9tJLyJlSi1gjIMcHjw550TMYCVmhJyA85NVvxzwbCd1PaRu3zxhWBAFh
uwwPTz6WFgl5wkvlmog/pA2VXzm7iUTTZe9lQif55/rhfih2chz5W6ZpLeaPFXIYNCjdbtVSNRVR
ch5HDI0lI4qqDOnqT2ONfsI5VlJGU0hveScq7r4W3MWpVDQqlR4QWVMcy9DWkIk4aMQ80NccLVUZ
1U7M48q9asKtREgsWlf2GdOnu5wPYt6woT0bET3NojtNsP/107KOZraQxuGMOWBoJxsoFwOHjpAa
ZuVFz3Q66yNPWywcSxrWicfW6bBr2M/VnP0HiiZ13mhhaxuO8bT+rUwwFGy063Q61fJm2o85EmW8
qr7qWIAkRcT0yyuTVulyEwgWQ+kNcqKkadd3qtM5QaEQ9jSx9HDpZqVjM8YXQShJ6J8PT8kRTKll
KePj6XjPN17SCUaBuAy0JtAnkih+4CWDngkKW1M6CH35e2rbUeA6qhDa3vMHsMzDs27cHpLZNxkM
l0BfMmEvTw5UZF4m8q1IpszyQIXq+FRVi8Yaywsj1MFAYxcB6iaq5tFFOcCTQVPgmuGJlLCFgWUI
Vq9j2QpQb8hKjINw2CfpvoBVwWIdVfJty7BSHDeC813qBsYiwuVEtHn+O7TK05b1UKVtwKFQXzNC
lbL4oTLzR4WLm8pchanRPu1ta4MVXdemo7245nErMIXEpE5QbszcIGQR3KlHMv/Kv4Cj9mpqpUo+
jzxEGz5d8OnZZRmACBvgYg0O5FysPEybb3p1uSU7JKeUHOeT4AbvmguhXZuGtoyZ/aIbqbWZfUom
rcYHDW5LNM+FuUBT/FQr45Oh9gyyexfDIv/rNyX8/Xj7o4yiXNIa5bTzSpTabUxEqk6v66Cxif9U
JuqdriiMn9iv/Y6XxUBpTT3bC+RNr92p3/TElAN2lT243AZAH3czSMHkoos3M4ps1bs1ixkBnGX2
K9nlYOugIolB7m0/VSdgI3274qyBY286c4PaBvOte00+l37xCpxt7yDyX/KRUK95gUuDoDe/xUr0
d9HEW8PTl5ePiqknt8KR57tA8cBlVmADPKHeeC8gh9QPd0G8dU6OjVl8I2GIYhWpfaSbCmsw0sQ0
WUQfSNfYYPlZ6LftI3JmYuY0XCAesAL18e/H8ZTPmvm58OHd3UgcjdXQyWxiNZAoWEStKPo/I6Ce
ZhXvnVnTp1p8ENJUSQQVWSWUeZ2Uhkwj7oiREMroPzrnBVIsZXw+2ysxU8Nc4Mh28QzfVkvVSb6t
R+30hgkSwEEiojgfizA3vRuyoaTdVcV1QkDQXELaa1gtPbFoHwgW9mUcEFpR2PHW9QRqMFWCl44G
sjXsbN2dQY+KCHbDfP/Fs2lLztRYeKoZ7rhE3xvZ95M6jCyLgIzRqYYJCOJrL3U7iM9Ay/sttflo
80fql4uwL7vfpVDRkIqPIAGs7fXk8zzPBt2I1RBNC1MXnOzD1m1opg6ziI+TIU28G74C+YWjPzwX
qnuRWxyzPAAerCgtM0IuuyZko1b5e1SPxF8aZZ57U/z+q1rdsINw2WRgn/2LVKYL8kBdivPikwyF
U3fGib3kb6J5GjgH2CsW//Q7/38mZw4FBSKtz1C2rN5mt3JDHticv1lQzePuu5D6cP+LVTta3qw/
qAvufZDh/tZUaGtwEva3ISywtR/d7I/yr13BZbt1Ne/l5dJ1yhg04o7TfAAXMx6YcDqSC7nX8ZmU
j4jrk15CEk8BtNUPH1pMjdz2nBdO0+DFa2dTpnQHx7tlfrd5wz0jaI1RLLRtD6a2tcYVXe5NRw2A
zY2+bzUiigcFtNVW5ESprlrdMpTxjYrXfGJ+Cxh+ye+EUVfqhBXDMz6BALmkzlESZrCl9PkKVnwb
uYgOXGsoPsZ22Onk7XMJWfBhyehgcRoyFsttgP9VxWdh4RPG7gx6MVu2DAvm9MoBAbmdkuqMVq1l
YAJZhbX3OiWDkzXKWdTy9Igv15/9sA+6zQHxoC8SBd1r0sO12g30I6TXamQX9BwYmufXGB4FLC4U
W+7f3CffSvSiwXR7IcpGeDFUAmNXxzc5ERUcFMS+Kzm2NXj3yJFz76t5OHg+chg9orrbtdns5wm0
d7jjNoHkF2PHxqNHox59M1tGUYodMQKABa3OVeY9me4M4OBGqEPAbHC/QCPGc3Vd9HDPAT3gre4f
sFdtAsZthU2htSPwEchiSA41ggN0Y6p0edhJIC9rqi/xntyB6k5GPkUG9UdeYpeuB9D8tCDHdtu+
cvh6fkDfG6EBDTpReydYwOB2NMYMB1jf629v5r/Dr/jGdN535oFtGSAU/0ksSPWDBqnvLJtMJHN0
p7eXhUkCFYVBKJRWfMX4hRvOBCdtGVQ28BzqApyTi0Qzwcr/YIqoLy9JI/uMCbYc6WGalKc0bH/h
b5IV8WufEtUMD1OZkL75FGRrJIwawSiThgQA/LLuwBxBbIU1hHjGzRS681WBZcPFe0DUUhlaGiK9
i8lIFAoZ6NtPesIqe9jlXfI8pURbpMBqhMRIHc1BUckq1ggKp1Acog1B8bWlx6YonA9EXey1Kap8
j+iEn8enmDcBA/RcCiUoho1qjrZTKVIULTNYyB5nhloGbzNUUNXHypY3Ph6KLsHX3Cfx4Fx0thXI
NuoG2rIN2YS1vD1DuBLXMYWrOxh/mvWzx1zHglmr0t1JgE+PKAZrxthXve3YHK2qFuMVo4eZDXPe
yiDwzxuP+b9XxGQsSYoifINRxcpIixOgZNLIiIihYkOzDXuuNZ1pxwLzOaJUD+DOa8nMGpO0FxFV
sWNVtaZVvlRSwQjrNb5RkWcdIl5IAdYVZtfAA7Ha/ZA0B/0Tbw0Aze3nWi8zJ+tCECaeuS0igWh6
dQ1ovRpsaqiMl+/sqzTa1nujKIT6w1EMb/CT8y3a+gq+eIih8PxThNLodOIG4y6FL8tjFQQGy5JR
IgPXWB/koGHazFa/LfbakpVYQXm5KWSrJ3WcEd45lCVpiFjvwQ5QiuoQvDN/LnuK8QFbwTcMspAL
BxytkZLw7aWQkb1cXQBH6gdmmnK+E/6BarZgVPPkqt1ih5mgp/a2nyeJubx8owHxBKHnyo9TvYfS
OVPfZDlY2iaVxQTy2RlncHu91vmEsMMuzPUtFHknxsXaXlfqI89tkS8PVFJqrSi8JTiFg7be3dIr
O0WUCivIO9228LfL2spe4maWuZv8dV0wCA2zlpaKcmDZN0seoiRjm5W0BtleK1wmcEcN4DuAhUH0
ytpaEzQmbspP1X4+1SeXhV32n7QGGy7bEN92xgfuIPHEOK0X1vfTubkKWX4FjRlkYheuvZokTE3K
HAx+l9ySknhMCZgc8Da1MRnGroUDhOo5ITVsckuKeiNHq6V7aJ1Ndet6EKHuTcXmlgI8Agnfo+zw
O4kZMlX9+nYRCvDHEUAMYGkXYX6qZwbp/0bODvna3zHyQ6nt2Uw+3/gil57fULO6TmoH2U33NS4f
j/fScJp4O4N3LDDe2KPA+faDOSxp+Nsysr1zqzz4HyxWgnShj4D3+9W9+pMFryeTo+T75028W6gk
yYzc2irRJZ6Z4NKUES1QlQoySQ2n2j0v6dL4aye9hRZXlmEfbWQXB96NblR3vA5jau2MF024Wx8p
gbuFIqcOQS1Dx5Yicr65mUFU/NhPsWZ7hGC8zDGncR08xF2ONRA2ldr1mxnQC6G9Qp4qZ2dOuqH1
2CmlKfsc3w8red/xLidzHUwZEUX2UrwCJm7l0TMfyB1HTfPUb1K2d7GLdAJdtTRk+8p2hiD+Sglc
QT7KLP3HH8kZ/t2CmKQ91g4vRW0fmb0tc5m9lFF9DBbe6RczJQoquo5BdexwFcBl8/nwNp/Pxaox
MY/adBZwoQUiR/OccIITX7+xwidHsCEW80Amc4ktkD9eT9GDnQ0m0+zySHheNGlN5z+aSv1mZE5E
4o88xLAG+M5SnIrviUkU1YifoaXLrI7CONjaLvI+oCHhES/A1Bj7cfMdsOhKGLyRSBETm2je5ehF
xVAvyx0Dj99AeVDjFebv7DSrFi0nE766SRGIpfv1gZ9Kc8Jiho4Vsxojh+AG2IG6kl9K0Iq7UOig
u40MgOCpL5uzSgRWmH6ndlT5/SEDwuzWl1lv8l5H3bQ+lvZdPLeRDa8UWWQhlsjNwKvytR3WchOi
pHe8LlpEmr08VegH/ww1eue6e9Orjr/ywDVTze/OTs8u+TDFh/fA/k27irsaG+TCAJfjmX+BJhXo
pRHEBRPtCppxIiTuwbMJ3LA/+YeNub0WNikd5D/WYDrNxZeA+jQ1xgS/kPgzwI9WA7itzlVavYBk
meFpg+fKAAHuxKJivH6G1M4aQHzzMP0Clz8JJEhWZgocwZtTyR2omQ2HlJ6vOL2tPbqdBOC+/5gX
VXdS9gTQyg5l5EAv7Oeugok8WeC+BhJ1UMXq5fo0BcrpxcTVeDBVENb4QsiMNYggTB0pIpHIlV3u
DwlLViAHUVDiysdTmUdLA5z4geY5Hy0Rq0xhBZ88ga2BR/vslrhI6yfapsYfaFUtOgpiG/Wmyt25
wpwzusFlxiz2DOlT+P31B6mFPn6vcKohDucB9dLVb25MuZHmAa8Sa08X0UyzuCjarcCd5wlQmxab
oGqHZEOlIk23AO/ZUo44n5G4EFIUzU07kqvR6xpsLneA/ipzxcpP4J87KOC5xcAwo8YoJxKL70Kl
2Fygc/XA1XiudU1/SXroumoO7XMYKGtxKGamZPeCRssQf/bCQOr+5/p0rrASbOkae2cpT+26X7ag
lClnI4840jyo1tqDjSaPUbMNX5W/EF4E3pPnUwZYhfCp8+l9WPrWDmLUpfz+3WWaC0dDd2kJEuGE
WxCwvaHwGhk9dvYsxvy3JYboIT2LwPJQjBlNBl/SR5Y+iKVKYUPBx/xYV2/Yl2ar4MIsdwIf+bVQ
DQCr4uBhoD8p+NLedxEZEK6o8t11ScWvGObre7my9+HjaaukkGB0dGHsDVjjOpCXlfFG6WVEPIIZ
ZhkJ0W0uUEPWYKp6a6YbOj406BFkeLajTzvbPXV+vu/b/2MNV0PytPtJNSfOGULLFiYpdMic9tzW
RLh3c8GH1BQk8c7V3s6ujoYI+NTMKHZDjNVaOoqSCc3rAsGHhqIMLNlFqn/EvsnCurPGtelgRZSX
a/qGHTbvfjFueWqd/9LktRBUOn8grHfXWGbw3rKsVlPGNz+Q/+gwxNtey/I4C4Er4yzPNLbJq3F7
K+OVCAqGBFXYCrzv9z8e+POy7hZkR/FE8RluToq6Y3pmWZ0RRF4ipAd9CZWv3P3Q0SH1rpeoBKF+
jRqcIUon0JLzIdd2pEoePcp0RT80UkMfSOjTF2pXKvVCAIpT8NOZCOcQLsB92sYxumr4CEMwGuz/
GViSxAGVSqw7Iij1sutSxY5IErfYRG8NZbS6gAg6FoA2b5FNM863lEAEKaICJBoUnGdRaLiCVd9H
8KcW/V4Td36v/Cq1AivAStt0Cozl6EVvBk61YJ2MPw2zhlwqoysxDgW0XHNzmUdKqGYWQkRe0XAT
5zjPtdLWYZoK04MamF8IZcp7/Gq5sCKA/BaVC7dqhIjpahSeqiMudJgu8sMopT2CeMgoubNtZw2J
hKJ6umNs1PY8i5BQEjF9hdWUBlPizDdEA5RZayoAsNVu229pvWgMzIoX3CBpEtZcWtkT23KEYm7z
e1f1O2192QG4XV050/1BpJpvVcncvNDtcugG9CUpI1a3n7aZM3l8910ct8dQc181QtYQci0y4eWR
1CLmfWz9tZZwidoCLTDr59JdLfPAP4hRygUS0Z8vqbec3wEziJ3JJ4mpR+x99lfsGvSeN6ge4q4u
XMlazVARE3TOlyEXrMldcliF/BgLyE5nG3S6r7iKg+RKRHeGchZdTi6l/1lKthWjbRDqk6LX7oMV
pkcztiB19+DDDWI3UVGY3egTohDmesY3IiJZBhRCFv/N/2dAbFJ9ODNK25iUifpbJaijC9ng91+Y
g1EG4Us/ybZSQU52cOdFOWoEvRnErXpRGVZ9DE8wL/ZdkFL9gL3x/7/joxU2lwBYN44ZdKelyaaw
hShsOHd6Lx8cgtPOZlSZZwUJtkiSJfslaw7ODu+OeZIt60tX2osFNbcn/nH9qi+NQtdtkX4VrUpu
0QHciUvvSYbtUq0cB6FRBizr54IyU+IwPlMo+mVin0Mr5PMtjkXr+cZnOJurHWbcXPRlmAnS+0n0
q+TwcHXmdikNsPWNwT0vwAKuJXELWosq6bvpg30UNvYW0jA9tByMj0QA+XqgrvCxVJpeZH7HZgqM
RTSrJtFWmTCA/qqB/Cw+Aqqk+MPUUmOIJqmB6qGneqz8PP22Xk9LqBRiSgsgFlDD68NPB/kIuCHe
ZwQH1zlgLE3t8H67AoffwvRD4gGElz/p5vizCMKgi/RJ+oJNEmqL4KyQivbb+nwyLUs9mCd4cukV
2Pfk8gQg76BTBK+2pu3BHsSlf0/FJZF9pS9MLEeb1Di3oofd73ZhPRP1VlHuEDa28IWyWGU9fkVN
J2HAx8V2gvS8rwmrlvw5053UNHzPPL0sx2q3XrlzFM7qBcMmJ99fXG2FEYFawib1cLrq8gv5OAWH
xmvw4x2J4FNV1wWVWo3g5OErHLDd1UZm1WT8u2YJoBcrXquxQX4gsOoNR2OQaoOUw3YuhcGyb1Q6
qdqqYOcC4ApBkih2v7bZytH/pwNIRZ5i3CSA9ydSalVmWfFep+K5ywPir/6JXarmxZuSJTPK5awX
lgjl9k7MXR2FhpWv6AUT1yH8MTWlbHVykv7Fc1vzcZctR6KyfPlAeDcfLGGiRfCtvn2j1lZ2/ZW/
EMVw5xJbr/piPFUXu22jGjyLDjMb8qGEXZS7VrZSWUs36fm75MbFSRlqSlJ9UPS1K+ndkglGxGoN
h/vpcvHHb0HpFqpEJBVWCKE6KbZX6p+jKkFIQyznZGdNydlO/8XAzT3ES92M+PDB36aocJkhpKkM
ZUqqqO5UVp9qxhlVeghTy4ogLdMDJBYoR7PCpua+qkXZ9oTlDJmb5d+w1VmOKVXf/JgSLCqeDoNI
14PzK5RG8l+5DdjPzN6IAFBK6PiT0zVO1fsDFhnVOBwvqGRUogX9j7xF15Px13kzJeQytmMdEdmm
hhiTlpXSu12iEuJEAxTm9hkS0BINwwhEbYXcDl7EG88aO2mV8K4lPcpb+Eg8WtlTRpUfBDbxsiFM
JslEJXSmhM40QsK2Oy/XTfPByqP91r6+OtbnI8WOuv+gTVKzR816gmud6ETHtpbKeuN2EsD6Fyh2
1uIq3cFUjF7J7J7h/ma3KWaA2ECqKVHW8b7dBhr+XPVSS819bXPXT1Ev6tiIdwqV513ajt2dgCL2
wZzOqT7s6XNfyEhYwV4HlwDTnkCDpGeFwAf2LLXuRBnHlB28+t7wmy3q16UyQZWjHB19/PszqvNt
9MpX332TYfD++C93SppHHQm9ZRxLwYBLm/hEU/rYpbn6SGzuD9BmWkmIqowgqjMxqpoovc87SM4y
asapXGqR5l77GRYXvj4JW6wHwAcE2UgDt/DTDWYBi86dUWP5PRuFALQMtlt0foMk3Nn6yUmOOTu6
hIeiIEJxUopM1B7qSvsXZTD4aAeX/98qD8VH5HhCDaI4C78jdOM8+buR7VXdXjuSxBE8UjULJApA
K9mweI6EeAoFzMXLE2k9jLcvwB3Wqk8YaXqpX0bd9KDb+jhdbD6/Z55CoUI/1rjZMWSLlUCuIXZV
fQ3fo/Bru7ymd33fe86BXbJua5X/z6IFFnT/y66Z2vkEQH9uoyR3fFz7O9eqIm0MtFCK0IBjCOAJ
iwCukhVNLwD/v/LVssSe5KMHRY3UIN5ZNKElNxuylsvRnDR7PmQ8y3KRJvnDLZMWq0j2TjNYu8zG
9TpSTIA6QuSC/Ue7cfpgYiKyqAUpxMSh0SjronxTr2iDAI9tVqSglkY65N0xFEK2ZFXaodVd/Vwb
TQ0PKqJe/nHVKz9WtLarlAIyQ6Z9bcl0xc6SO+pJQtrqbzjzFNAaEwTMBzBKHhrjYEW3J2vaRiLP
K5PTKakarpXfvH9Wgpw+y2Cuv7+HXpHMO1GFZ/fFUGin0dlVGBnO6cZLumMrfNHwGwjJnq3q6UWY
jKcTxwOzsnw5IHOuklyQyoKnVep0Ls4LxHavO896CWEuK61uZlg/Vp/3jgJtkvB30xIw8ooTSg4t
HdrcACOyyQ/9gNcrK7AyFUdG+RcFfW/6fb8OrkOf3Z4li+rCU2dHMGxisuJF5ZGUPdum0BCDaj+E
kpc+XyuiZgSUOxJDQBUJ8oaIbIxn7EwSMWUCJvtkLVbjd089DXfudYDDHFIpaXdcpI4Oh0yr8FiY
fLnpp+I42acsFq4s/d/4PU6AN72rJnDKFh3/3VuiA+TbsAg+2XBksZWBBkDFJyIUliRkk5y+5EAq
TkZ+PWAPZ+tVDwlE9Sl7Ikn/DycqAuUdw2L+oh+iSr9YpURUWJWmz4Orfg9eNVJb/y0YhZ3eOC/4
iL8rk/Sjc9QA3+/G9McCCGn1LkbO51vI2l+l0km1wa7WCjKu+TbnReUmuh0oJgzOKzY8kCZ1XBt0
wKuxtdbOzeYm/BGIdYDoLSONfMJpCmkhXnsQIAX8AukMzabnHltVszvKKeIhxomcaEAWxsGVn59C
skD26TtqiMg9IxP0rxU3LCZViyeCtT/IeKhtYGIFbt+TQcSryyv2sML9FwPL0PcgJ0JrihAf2b/c
SUdshelk1RfuMCy1eZu2wAr0iobyXRT8Y6dZliRn/uON3qOYCZpsf7JViTCkWQME7JrfrTj3+fEy
o5bNnUc4xF38pTVi/4iojtE9Z0j9S+f7fCUvCHYvyw8fengJQ7SjmJk51WMU4BTOXOZAa5BtgjsO
NSRLBm5kNQ9Mevv1Dpjhv3sfm8U/G1WbvaRgp7J4a60RCYeCulSEhe1hmnzAtZgFETKGodN2+xZo
zdrAlhlEJICvCqCUF6ZJDefEBxZk44wksv9UyBcy7EFdOGeDiLQ8Tdg4L+DD4XULEyHx2FPM/Qld
ePcWEQ1bKWBJ3YFIsz4/vclKO3MSqYa8qvrIkFI8p+7EvMxujtb1kIkGobEFV4DQwnae0nX7qSCF
+0IeYnw8S0r320xRiAmznB+rjUZ9TUg6fIP6RlurvX6BWi8q9X8ZI7MFoSORAtGUcoUOYD0yHZ5Q
Cp1Q0g6cYodKTjmWbI6wW56KcOHbAu8fNrQfyzLByf5loCq8bAspEug6Gzuw0KTF1xxjheJeR6TI
tWv4gghnd3FponxZuICEZLZASqIEor7TaAxTWdi1sillgjFn/5dTiCIng+/ieZqMOFb8Yu1mjKYs
7pyGRmzVT+UtpBB1kLOCv9vWplYY7SJPHuo9yf368lLLmRLxsRwiLOl/g0JKlyAfe2GIONnCu3q+
hk0z4BVnro1k3Rh0/QN2hMJ8oJxEt2tcmfhohwTey24ptZ+SF62bZCuvav5ldfYbhFwzmERovLf9
4BWGs9UfPpSYdmW+QGAXghfeiAURozqx2Ubtp6ltaIZtjeE+3T/gUPGJKDxFAzXi3330cDj8cZux
dB+ihXBQFu2rlG/osCcTsvpnen0PqqKHmLM1SZ1NkGS62wZSo3UCWUgTPz+cvbSykRyQXIZMUCF6
L8fORaLt/0axo7UV80jrIak6lKrzFAr69j9vXJvHiCirSlu4KBj1DqhS917q6V8rH59871sOGEhm
SB5VPR0xuJhz9sGHpKX6i2oCzm/NLrYK7o8XUY4u7EW8OFhul8Ch1Pj6doMEW1gnQYOIhyUsqelx
mPt/rNyXAcsUeJJi90drGaLsQcxvqaaN87vefEB1uHl3T4HE2ZTLhgk9j74hgCyzOYvUVjkMNQvP
1JdELpFSKMB9wrzEWaQQj1AaEWyYoUPKeplKrYZ2vnduENIPUydvwKF6SahRK2c6L9xu03SYe7L4
V2maIXHqeQ8rtNg6hdrACtiq+R/rFfAEw5ewDg2x3+r6dkRRWJIbSq5BoBmUdD+PFug4i2fFo/Vr
v4di8a5ZXY2+lnctnsR0O6GRO9/2mDMcZ/hxh+jy+i6Ww+rgiIlWj3FIF7xe6fTr++T4eHv9DTJR
iE3+N/qfbinI5EMqfhbHcu2L/tCD9GHHdRySGOrrM3AhQg6areuP4qYs+afx64XnNvGiJz+P7Vi+
Wz952kOOuV7ClzIvJU8jvD9Z9Dh11sbqCRG8hNBfbsvwKb0c75oYaYcWW/1nQcDl+zPZdRlWU07s
nY+QVFmuRktP9mlW/xskMzzyHb9l5Zoq2F6lmguOEmyQ2c1C4+TEQfPN3Kheb4L+5sSz6ATa69zq
FXkhntteakWrb5fSP4qbjds9TJEGbLBZLXw4gQnwVM3K7zCOo4NUjv+juQ/+mCPqX+CjHuYijbeC
O0aWvLBNo6b5+vjdoNsXhvgDwK5neVIEJYRHVJer9U/0NPtxmaHw3RknRcIUGMaPIUbjZXHjG3mn
xYjrZOHw2E+/xCrZfIqJypvSqIIrxTcxMedNXG4SI2bTBF+o/i+HlDDcA8mmvjkZgMCakxfpO7Ds
UPIOa5vpTYan26GNvy78qjXJCeKRiMe2RDlepPxp74axCDXKbkR/cX6ezhyS41GwEIe26e4xHQLz
AGr3Fge0BTldxoyvP8xgndMewFh+nIFry0fUYF4lfF/P6LyLzFsQbwvsLHMuKtDYUuwz2lyM+0LH
ILlvu4X+XdRqRB06pm3nCnMkUC8Fhh3tDH9Gh0uCrd+15KJoA2Acd5QnZhvdupuHEa0CjM0/sDpX
HglH1LRZidGyNP1n1RsYoTWTDA4Gxf4ImuRlJCdng5b117/n2s1dUfvffom6BScbUE9Cns75SyXa
HW06LxozYkZXbesMLUyO2Ers2yhpqMZyqm3R5H0JXPYv/Eo0ZlqbthgYoy//1zhjs6rS2ZleQ6rS
pNv7TLGmMPFWMwOJTSwfPrN74KUHcxjceTXYrMAfSwed5e/bsOOWwAjHbiJidaij9SxGnrTbDejb
yAJsEQQyJFobwD1WYavrZ+59HBmSTfomku641DHpkA/ZeA8cJ0Fjv2tQzGSyco8lJBP6qyn/DUFp
nGz0uPuNsUsWhMniUN9gikbFhxCu/dT8w1h6C4C4y/7fuqfxd4pv5yIBmDrG3BrH98xd+iXKDj2S
W6tCy9yYPpUvgO3JiA9yb5T9QgTkpuiMudwqFlsbTgyPKNPUFxXCkjuLmRCtF48wQdQY51YZtxVm
hKkVwFw6L+Yx8gMowciB2UfIx1PNUJwoSQXMitfgOici5OmPp0NKTp9HktpiVfCw+U1rA/PVbQIw
1/HH3zG9nRE+h3dF6+CF30rdhBBUMJtcxCJtx6w32Sjh4rPvyL0ydBgk0tdPApnsEmkQrkJshs2C
KvX2AKQSMM2cce+VmsRWXZOXp0Sp7kvJTbfcYk1zDUY0kcGuVfe3dEJIFJt2AM5mvKczvxpmMLzC
ngsd+1m6MIulYVXx1AdMfnqjcQcKW/z0pUee0c70bgHJjUHoIYUNFP64BU2Sf5O2r7T/+uOIKtyp
uYHwZ5pIBNFbQNuBjMqCbUwKz3JYlMwx9qpY3ZvkhlKe3UbGXTpUq1TDVYn4YM0FJ69YglMHiu1Z
v5uvepg4xtSlgbXYOe0nQ0K/ljI108yDcp+Jl+f2bl8khUDo3Mr+aBCeXv021JFNZAoGDNqMXxpN
5B599zbQQCTSESf6puZk1RWjuHItmKIMRv4GtJpksgkPiRmf1mxdoVghRgHIr2BIAUYLQ0sJNVUS
bkW9a3Dg9cRSpiH/nCWEsEuXTaCPQuA/0xTMxKI48oN0bgwJaEf6ugmXKuybzXyAa2zOx4V6K1Qf
knAmD75h5vqeQVNAS49rtCQSXCIWR34rffe+vjVxfTeXZxCyaO2fp/wDrSt8UyvcnxgZ8ImJE+gA
pmGOhvRMscBEDEmQMKlLc9IDGN+WhxE7vmNdkaSqp3mzTS2lR32NiVN6TPCuprgIm5gUp1ZhCD3i
DIg39W0Hc0SWp9qNRty6s3VuJ3KTxNhXlkflTsWhLCcePSPlNOHCAvxcf2Who9eLir90jSrum+vc
/EPcbBaDSxDbdxrN47zr+kXvUyvCML/zKIms/TJB1iTR9PXc5uihvL08FC1077SedXFUDQXXuehj
ULI6gi2vs+q6N6OMHUVBk3uWCk5jMmtyveW62sMXbSG+YnvMNG6YZOADg0ddhhhPI+/MPTY1RwDh
K5sQZLLlLeb0YJBD5tyDiSJSXH0XrM7jigpm9pOvaRw9TsuioJ0I7DV9O+7BuRHBUUk6w0Eaw715
qDCeEe4mzG+3od138veYb+PbAyrArfVuwu5bY7fXOKvBs4/G/nUE/LXy7D1s8Y4U6RYUjKhNwOhQ
BrXR4rFBwH3mxX6UTc1/D8N9cVkqyykVtBqK8UA6Yeuz9IqF/mLxF08nkJeosUIXjtYLRPHD80HY
Mj/hvjjOKreYbxha044De9X14TlCOvYKY2fvPqOxel4jJdepZmkoYfaVRZNqJjx1OUFip6Gs5utl
k94Jv3BWP136HzOwmJGQmrxtO3VFVIlyKlO1l3kKYlMioZOJYN0Q15mQPXeW9kMRVhcI1IloVxze
PXKwjW1CyKsaAklcP0EBO6a2oBvDYFAos66ZcLgZcB3/YC+DIGtXZEPNNTnLw8cZOhZWA2ufo1T6
nPkqSspNFckWYKDJJAjsGFdSwn5m1J+22+DYSec4725Q6NeD0rCuG/vKfrL6miugHTejbXqiK6Xo
Y4H1ItTC5ZjkCWU2x9bJGEUvNkGp/5CwM2pg9nfKlqitcXl09GAVErzxBT641fVY7rxILq8Svrph
0lDb6WnoOphj53OpGGPJh4NgpvYZz/UhP/ZiukikvPRaxv089r3Ulw0EMiYKGNVzheaTrqfjEEAb
wWa9icYV/EUqR1sZ3ZlJpusHVfg0kRSfoxHP1rJl93wF8um5TynaI+B/lXlq+srFOTgs1xmbF86F
k3YUbq1Z7EEQYyOa4CZZKl0g616v9tOBdMxhLMuBuTv0bo448SUX7ckhacFl1uBjgSFyW90QLQtv
jLH9NbUFa3X++YUX00F3K9+p66kYgEe8nJjU4wDqk9Maa/7fo9Ytiy2hdmcV9LCjzfyhosniVFLP
ICX/8E+8kPVxtpE6aSWfAc9q0hFlqLbLS5qGJUj9xqvvzgT3NJ9pKL9t55Odb8kAK4qki3yyJBPF
gNrv7ZjDnj7Il8jylTTEb4QX2m7PBXReH6ZDqp409P4mY5XaPgODVd87gZPNQY5W5IoeeQRDqiQt
3PFMbvjc/CE/TnfN/T3iuOuQTOWAD8q63fx10bOFdvneo+tFHQouaFVs+t6SC8/5YEJNPLGfimOZ
1DF8WG4gKO5DkDXMb0S+pe8THz9IPAVzs1/fZW7DV90FfSPhByycH+FF8foT+ZhaYLidG35A7rvN
COSo76rX1aXHhJvR0p8eSXTF12Xs4e4X6ZnUZds2SDxOO+Jz4wR5FzAo01p5MrPa6LMnAHaHT0Gi
hmoD7tzgbHjZO7wD7J06ZZk3U3mEOjwbzqTPqf+sx2bh1AelMlAl0sDyGmGfbxnQ0EjqKiPMibmm
aVhKiB7Ii143QCGwg0ZRSR/9j2nvDI5PMbbjuf5RHBaq0FiuIyCZw7K8IW/DLDtq0pGB5J/wZSTG
LXYxTcH+064zI6nQBQLC0YAnorGrlrXIcGjBikiTQJ800ElpXqrWOHPZ4cT+VPcsVjkYKVYWICYc
VwViLla0/geqgObCNwXgOhL+gaY8KEWHd54ecmNRQxNh8c24/BitQGQBWg7OP5iSzfKh7/w8au/Y
TW56I/7u/xvuU3mRcttpgFomn6B3eyEAPYseNEAn1N6JNUChN7stxD1HYfDssiPXCHy/yZXNXAuf
N+BBHOIeMMyij3gn18+Q7ppxNEr+JJdcJyRyqUhpYtmmtAiE4/MjIYwnfexI1MMrgBE8Mv1fbRk7
Zjc1wPNHohTqeArztFlX/fLCvCU/UbjRMGxnRE2oOMawXzth16lfXaMVHfVcY9C64PStOqkAPNby
nldQjPAZ5bp9jzpZ1g/S7PsfWgiEjDr58mag0mu1CRAj5AUEOi2N6TTAFaIS5xMEUsC6rV0Ts0xo
aRsX5wVMtJjqJCUTqIFSbS9qZ0KRrF1W/IL0g2JyrCiLVtRMSxyYcNOoOeEEapjWG5Sp1O0nIZVX
7VCeZc40KlOlx8pV1DqUUzudivMS48FpLIF/HoN6Rp1ygInTXS37xMhTVHlGWlIWzKSihngzqXhW
T0N9NtnVyv2PR+7NGpEkbnBj4ISmiMPqgp9DYtRHi8eJFc4sqv2CDvYW81Ur4QPAn2FYo9xnPgUX
PZTCUauQU43jo0gr4HE+98VCXI6QQ52PaJkXHjHOM3lrrv25YNT1UbTJ+nrRiS+/baRXCRaGuPi9
FWYy6ph14E37aasFg5pt6VLj+UzPuMbH+7yy7LZoQATOVljU9U4EIf4UQeiLIhJQPOdfUJovIdJ1
f6Cyutq+pwATQn0Z4kpxP/jNr4fxU1KHPSTCkyyF/lRpxKqaL9GX+l2+RJWcp/DQsXxwcq/Bf+Dg
lQ8E19oRhJihqn4gUMMJQo0HDC9S0f7HUDJcdG34GyVanQ8aKlZDphURtsnJfZTymKKZQ/zri/II
QjU2klyFKcEYbfvBalCUU3bUDBuheMXSdGcpWCs8+62PV8DLgTrU3ri90ER90nk4uWQ6DD6vxsz8
IB1gI1bVASUqUZTzapZRl8JDewK1ETqNdYvKCUpQNL7eeDFq8qLETL76jIFBvtDejuktOROhAZd/
t8w9owzvk1rLFkPCs+pTH6jpLX0sGzJOA8wj4B9wIoxEwIz6dkMhVvOgLUXA1re/IlR0kueyBoqp
ydhId8U0XDZsYSTFRYp/YFqBRWI+yMTJTXJhu5n6tmRL1/x96MhTf2vEQ5h474Vn6vRQ/M68lu9H
hpq+tz8vYWXo/6diKk+7aONDyCtyoubNlXi8mmQ4WTbzo34TCu92Yc3GfB/VCTzPUa/RIIZvUbZb
G2glbqva13bQlyeqWJr4xT/V7SV6Q4/hTbBtZOmbEw7F15vhbJiR6Iu9BGfSdWrlUqDACmUpuhyK
3hUajThr0EmLUCDRR4hXcgPughfqtXFIIKIMx8k91vylUZQMUhkn2r+L/dW3rDLxYPB97KrvC4M6
QT8qAsttOBbfYWGO5Ur1ew1Qv0RlN5VVAobFGtnK97/2beRaA+vYEC7I8nqmBkshFVTVForEzRy6
Cnv3nXeYFVjT3NhiK0mSD3Borc1zw1b5PpoAEIuVqUpoyajbq04aqJ+PFFCIk7pxGBI1iod2BWWH
mKqJHc3YKwzuCR/97a2HqVkHr64x/EPWJTF6Uszkoqb3Qq5eUNGgNL4SxBtF+NHUZ7dSiCGs79om
d62ZxlGP3GMpp5Zv//DaeRkIOqno9fVaW9P08RYGXw74CA3rJYyz4ML2fqYqIybLghBA/ilQ2c5L
/SMIkziELym8pSAERCzhzYXm14Vzt1QuWXtYFIta1MBStGZNeae1sCzXDVCUN9ChlQoAxmxxHJux
qq6xFsRVYWiKhYuSATEdix7kQRy5Dp//pAkVTERVwKS5WA5LRD9NYr008+HZkD3y513Kj0ea7DO6
cS8Gm/kDGGyCH9BqQHVvh9kMHyUW9Og+5uanSX9dDpnzdF2qOwxozUz8cjTUYacGggZ9evEmSdxv
Rtj6pWgaXycpnyDHDLwzPxoKAWecTa1Dk1O+1N0FZ9kCJi06B5I3TQ/3f9cdrmtEwHNiaRKsNRsz
8VlsYnU4pv7EpXkTEYp269hcDyW77y7WtvsJQFTXIiyM0G9Xwz90Tafmh0t1LuRTCcUBNIzpp5LG
0pmeKZasrEixeM/dMqHE3R00iZq3TDUCtoiKJYVgQawMLRJEpKC5ieftKNISY5flgEUrPm2SI7xQ
5goQQLEPlGUdT9u/GWHjQv9v+fPunnxhkzB2FbbqmJl8QDc67CKcbb+LrZgyoXLYbUWQwCBi7AYc
x7D9oQenk/BLBTuNeVlIQ4yokswzkAbgcajw/Jt2sv6qXEbUo8yb9IOl1SNdTrIdwT6a2T1TwO+Q
anqJUKAUeslqyb12vRpCJiaHtIfAXEiTNv5vXXrYgyd8XYZxE/+PbvOD3iIcgTyuWnJNYcgZ2zEk
qCG6O5/24oIJMxh6L++Hk5VSRSqlt8Mv309SdgXWcPnJXlCSbKM5N6tIdR28y4YnrVxswEuRWYNW
0C7oq312rkq9yi68QdS8J1ZjPrTLylcz4ge0YNUj6ae13k06YdGWkhmEhjlW37DHIgEK1GMPKYim
5dZmUdG3ecyxAFaiOnkhsT6OsKjornm8Lf5HT6b2xvvSWSvoIe4M0iCtNXxiDjcXLxWlc37ZI7Sp
MwhbUzZwbo/Y0sCStB62kH0+pGoQff1JQ6F8+vasnfHl9yzJatGwxa+iKn0bvlK8v4ZqGoO62NdJ
GgQYGdLAz6muO77qqzdK3Kia2muX81FzDqBm3rMLqEGeSuZkdqo3ciU/ki3Aq1SsbbHFf4dvU43e
zaHtO9qgKDG0Po7v+O1AJRLkf7socVde6Xe7GPIDHNOAPrs9HOTrFIr8O3HZImmLtLbcGtfRvXUp
wF0hVk+mdpBVnzFEmOkKGVqeR5xrBK5Kmx7UhDzZalhQvJTl5tqBgeyXwvYADgXL5bWnomh2b0g4
JaTxPWisw70oNf7Km/y+SjnF8ev3fqVbRpBHUP49Q4q14/ag5cxqC1eDZaYrG9ojhMzknNtWZhUd
atcDOJcUlkMFKIIvHgOvM+qkrN8/r02M3QDGHRCHFH6Ht8eZoSLHa5STvOrO2Tam+CUIFdmBpwXZ
rdKFsNdqmuMxDryJ8zOgr80o47lfXetzpb5pC9HX+7dqfjlxkiOO5ENJexwqKiXfi/RdSWPNZflC
7RCQLf2vDla8x/SRREQqCIPFGnSsa5G7beTMyCtR7q7BuSZ1NlFQgcMOen2d3g5MqDcdDJ70L5HF
jsRDfhp8W8M2uasaLf9ANJuTHTcSmYdrAhY724ZHMI/1mwVMbTSjwxhJFaz3qWHFolew+UkIGzg3
KrnOGNomHcf9ThR6+eTc7AG9YFBvbC4PFOBflLWOujTqC5BZczj0N61uQkkpwFRblM7o6calOQZ2
zjY2r1WTNQOLZDVkzphXihyLgttTw46IghkX+XjlnaFmxDqjNZwXCqrBbHvhiYMAWXc51K3zs6jE
Okjw4MNnw5Lxwyz2c5gq6PGzZLPPV4dOQFEE17/YsRewXMb1a6SchglwII2POaytGWPAY85vXjc0
HA60jd2Sh0oTSqhHhp3vjZY45ERKPWjw1OMc4nrDysMR56fSqfhf0E9sro2BU6lPC2S0gcJvgCjA
zUKSbGO9kaZ0RrqlNOIzYHV6fdRh65jphKnZFMWbdtd1Ucn1V/EeCV1BLYTT2iBKDZwVHXl2YjC1
+FeV4nV7QhI7OvUhNbvdoxQAfPoPqDF1R29u9R0ZWdtaths2OuVaujXgC686vjEqLOwbtSEkFbf4
1yI5PVdHjs1bjxYmkL1tZrAjWMpAqqxtlgnLKvnwYgkJRfyNwqPUgXtkmn+Nnfq8IfcQJCARbqVx
yOGkDV+w/FPD9Ndtps+d74kA+NsscLK1wsfD2+bLC6ew36nnNpngviHuIWIHf8ppEb6CQM6yGvZO
a6qTFsZFfU9VvOePci3BgCdZtPlgzAbvc5tCjBVy4ipoBRkKpP7GlVJG6JG+kB5n1qpIKKomu/FS
hb8eONA+HH5ljXJ2yzb4d0HsZhMYkREVbzdREnPZa2D/phIaFRUZNI8nJywFzdQNcP0rYPkGUIdW
2BLJfaeDf8XZJR56RoDt1yGmyjfyM4OIjrm+4gWnEsu1vU5g0pGEn+CU2H9vJsigzDA4BaLDplJe
Lbn0nVMNlIS1/3LMhXD1wgB/j3msqKIjRxskOcniKu5nQC+HQN9fPeAO3tPljmNwct2VmYjwLMM7
PuZK2FG3SwhVn6tE5T2TDgaW9clXCOSTYtsYKVjD2tTnVM//z9uCUv37vQ51X1KoKER7toppmM4w
mH+MtDa++dg0dvA8CUNiYob2EcRPeshLalNaHIaELJaE9SmUlbYwt1QuA3RqckPKEck3OUs6X5cM
os5Qgmmc1OUw7yNJmouajacPbR/qMILzZ/3TvDuWRbroajdVZri1gGy9dcYy0qXBDmKg/00G0250
1n+S+V+hC3M+Y/SZmXhK6wyusoZQM4mLO4hpPDbXrbJyrp+wxEKZ2cxdMlkF1uU7nb+s+T8nXPG6
5OUwWgxc3CUY0ih5CvGkYESyyfMItX8yov8Q1xsOPOE8Usacjro89SAGMX0I/k+UYZq5VYJGLPr+
gqhGgy+7bY9qAZ9/4e2WnCbUbX8V3aDlJegPkmw6p1uu1T6TuVoP5KPP+eof6Kx9Z2ov2woiAIFA
cBgLackx0WZGB700/kLLWaSLzpJhkvSpnt8RLPVAlDllYpzlm5r+Ensei07Ce9zMODqHAoebLpl0
ROE/nYiiM63cKZQeIoXsK3HQazaT7BpGL4vV63kGpN5nEB9P6NTIZi3eckZ3t9A9DTy1WOM9HgMA
Sftju3GRavzLc68Jf9aPjVWWA2gDfwx4/W6WXiDWJyrUvIZx0q77ryiLBMjwTYj/fc2JSw9/IK7x
cqp6y58CbaTBVnN5KGtXRe1KRhuUHyI6meNooirQ2WxuoE0RoglStQPoVgElIdX6hbEXWjdyeSuY
LvGYOFJAHrsEooD6SBnUSsgJfOntk/WNY55PExztrxffka701o7LHXKAlfx5iF6uoHKZBBI0x2B1
FZi22TfcVc9vEsQseklUDlQePZcxva+ogA7rZEiHjUFZDYgmMiGZlUV0gzOzmj1y9qCKgty/Gc/N
urkfGTS+e/ysM6cs8sP8kXDU9TQU2QAvJKun8JFN7Vu8IXXAenQGa4HaFCEj6fH6gIzlZN0V4hCG
4Labemva+u5ICzbU+yi89+4rUXAJO4KEGubcD35ZHXLCo+gct84e8eMlA1xDXNtt17Ua2IdRpr7l
rQEj9U9ONeE1DSz6ezKR85Zk6tfe1WaGhcPiVUv7kZVgDK99TyZM0TkN9hpRagP8Y4uAreY5Yyse
1seC3oYetApcIyegQ/URWoVttFHU7WupcQTAcUysID8mX6umm4o6N12bxZhcjeAhknMk4GIfAdKa
CcQ84oCDkfYZujqy/CauK9Sojl/i6i7O1A1Fj/LbBD2/0cYGLbfETQVeql06wf1woNP8JRfupwq1
v3plBg0GCYLcjAfrTmZusnVnM/4kCR6OMxa/EdpSw6/DQ0nekHByn+LTCD67vuPootyzjYuKYHP4
/Ug3HVULoRxdDWaYZ+lma1bfjozjavECsJ9QKF+ZztSROsBQP31s2REePXnLa9z/WpdMcj3lNj4e
u7hWfhB6GqhYiB3mZ4fnnNk5aVvDDTSsS81OdG7+afQ3DVvtPca0EcHkyEMrqGZMY6kTVMTstJ37
HME8Lc/y4AaYoRmds8bK49RZeeypiQxDUelO73P01daH5E+orc5QsdNONPWg4NSQhVxlQWNHVRah
+e5kqf7Qmf4atiq8zVEWz9M384wt3WzJMhAU98rNTnF6c/BzPyWp7DdocO/7SdTy/WcfV37bORbJ
kzFIM0JKnUoaJTqF9kLlGUUvcPYTL/SkbBciEAzdVB5zbGONUGb89bMb6sQagAN0t9KOfUJJ3fSH
I1YY2f71DYePX+5WSeW3eyV9pBhRgo6m52iVGxZAitGKB+f3hoUY+cOyBAtFNTYdFm/CVAAp/mCx
QOOY1SjYcgAN7g5D/SMqgFQ5WOeI+zXTeVF6Txnir3ErS25BuAUb0A8Hw/RuuGbqA4bJGk6TGb6E
UYXNOUpa5Y6uzeS4WV0KgOoQoFL2rrrj3bexzbZlZtlAGZELKPgygsH/NbmLWoYTC4XdsB0nQVDm
R4KUyKhlht+uaLNJ5grVJhKsq8lsFGPbbBGNELoLZHroHKuC0xjr4M8G80MFhBoDhGIrrj9lbAYD
Yq53R/rNvp+hwRdPvK0qDHil+bSpV/MpmoPHUGeadviEvCUfdEDvHrdVYuO9c59k6nU2qx53zewW
PJEpeUx+WMqjgal7/I/hSHMVFkQ8LjaZ2A5Ksank0vJhFu2bp/aA4NVQfMmZM5WuQnyJe4p3moSs
4pEj76i285dwX4ZrkIlsxlkhMm8VgVw/JWAa+ZfiWV9GU2OtqFoG9astrqf1Hx6xmxL3HRZ9T9Z2
1tBDBJ6OqVUGjdk5JySu7tWAfct3vxAaGBVUe+IO3peldBxVJTiShd0pkquN4Wld7wOKVY1JEaqT
3KYVIOT1Cx8FNHRtTDWKpZtRgaBld9oG/TYUkPhJQiEKnUNHAM/FtA939vfgvrI4wT17RiWoqzxL
i+EGgm2IOGqhgTGTVSXkGe+ZHstGzmNSTcIIshUiDqXpB+XN0iWP2RmLkSGd3Mj2ReA7HD2GC92q
5zHr4ktubIFKMJ/Gi8p9Av71Be7PIs0XhzbM/+FrEu78EZLVpR4BDBe7x4C7Bpzm45wlighV5s3h
rBEB7SjIcMCUBJbx/pjWAAfV2edtXFjoqVDj/jfv0Z+KHbbaC3tvH+zNrKq0da+wbYbVk3+dBnbm
Y1xSD6dNPK32g14v/4SVRwAxZwUBNfwHhiMAQm381ZkxLc7vZ+N+cw0L9YzoPIRz78CctDXLUPD0
majtIy3wgeRM0b3NSG9gsgm6P+fwgxySFz1838Uu8+m1ya0hBlwHKWnp1Ko6Ng0oI4mbQ7rkqTyj
b8u1bw563UIg/zZ+wgQrqIhavhdVlwhMbA8DN14gxZxTAKXGsBkBJjC47/beOVrM2jO2YQPYf1pP
osU1W+JXlllKcOEcKrJ6YogmBud2cUltArZZmC8j9T3Vl11gdNZ+lnDZVMRIMhSAvoHaTdSYF4CM
jwDIRSEyY8JocNjsb+TS3Z7W6MjGBAIT/jGwjlH1MgN79IrPI+yKA7RViC5cgCBccBGkpfkntsdz
vTXoRnsB/EYxNd323BPAs62W+ZJX/13zsZnSMaa4MyDEjZcWDduDP/TsCI5TGKsTPGWLaVAX+ZR3
KjyYCj0+xkp52rbuXBFWKW4cUknu+xxgdgylI9wWnk2NR0nnDjCM8UA8gu0HGgawpv2sq314uxgR
3hA4jmwD9lOutdFbf8tMhHIReqvXfREZV0xiwoAKM8ALoDoH/FctjOvo74cdELiOyUWY3hQ02tOi
2nZwtadCtDdSsCQv4EQ7krj5ur8rbfCQ9oIG5AXij1rRbs/j2edbblHeRKe4fy5s+marHEVicPbC
5Uz5FzEKoiOQP0Qo1cf+7ITdsTLLmigGjlSwCz8tX4WHvUI1+pIDLQZly1mEawtuM9pCEWffhwsY
An/ynwZvlNxb7IumI5ausJVUSIhrAnnfvySztc6fs7UjkIGfa8ImLm8imxoowcO8974Q41Xy1NJb
dHOlycEoCM6ejINGbf5Y5e/vUebN7OawGMBwcpkuuAXpKsd4xwCe7BKzZpMTVHpzOOIsoMJDm4kx
gz/ZJz+kd3iBAozMuAsBhaXZUMCCac6L4+HHIFiJeaWjF/Bys8U3mLD/j/Wv71p4+kFZI8Z5qyDM
bnMOPPVKhXtmm+m1UAcUBphiZlQZ8ZHZ0o/+pyn5RAjo+iMv/JjwiNc214alZT2daK5eq6oCUHhp
RcOp63H1x8on1Ucxd2RlJmpiaNjJ4MPiVkFFcVKdx+gAhJT1g2icH9AeEBCj8BTtZQBAeHv0qCJp
8Ev+A59ONNKT4NAiBIYgdD9pt7lt9m8Oeas4MZu4uqscJWA09w87Cc3mddBJVBfttXO7GgC7sKt7
USe7IH63a5Kl64y1OU7sHumLk1c+sCS+KE6gQWl4+8qW7Zw1XrLES3Nzg9ov4tAMDFBG7AsJfWs+
R+wC/X0iSzvRNwr/sF2Nhz1U2x7d/GXTDkcGNsmNC0mca+99hKmaDeYZByaD0nAS9YY3sbX9Wy1d
W8Gcddjo+XxXHgjkK8Tv5ySnIEwsP8Qyz4HHNYp2NIXIdtGK4Z3wqJx/HKOovyVbyDe1PKxcdCCc
NzQ+SFuM9aRBH27DJh607fkeQVNKZBJew8UIhbCtI69lZFHL/ACw0cu3usL+p1kqIp+xdKxBPvzP
2yd5YdLgRF89f+BnSMPY595jZXpZuPxEP4AJ3V9p4A6eF/a9OpwVeDF4Pd8JIk5/vK1mc5P77azt
b1DhOVsLC/yRqCbZk09zsKrrdD536yy0TIfn/20k4uyLOOtosN9FJ70D62wFtKoeQNTupjJoEsIg
ZMxNuHMQC3bc9qZKCZ+p92Wy7753X3cuEPx8fkHfr9LVa3NdruHYsIkEDflFoPM3XD0BXspIF5wb
u060PLVYmTGDcaiuVQqpWHhGovjLVCXA57JZsk4oTpoCulVUsFIartzdX5/W3/95ObfgxzUfs27o
wgo8HgPR/rJVGnURLxGQ+KaYEJIg6fN3dVwC16WnHOq2m0X3xKSr+pT9pYFg0MMmN6Z8NNXV6Q2I
0cU4XrouKzTX91/ja/r3X4EpYtlizwtQznXdJor1vgAy4icw0/RxMRY+Cq70boi96/VMgJMpcBel
DQ2LNIej+zZGTBb5KiA4KY4QgASYc8pxQ3cChgluXpjCNF37QXkSwo735Yqq7yH2p72NtibPurAU
K/i//6BY48dDMzgUtG9TDB2uHqeGBROCfW7TRZQh57nN6Mg3fhM9eYb39adYkBV2tBE4IznfRySj
gK0Gk+LI4TDXnvDKlmhpSasiTnZfrLWnaB4tVPrfL27l5URlcsjDmK83NAwE7iOuRLBOiedtc1s5
hIP7WAYFR/kYTt4dxoFo04S6F59Hb0Fs79wnTv+g/IJLTtYt0uiKZQBnjNxJG7N1Yv8tvtZjnoru
iseSsX7GUSbMu8Cj/h5+fyf8+Lbkm8laFcjNZFA4AYGqjp1oqZ2+WRLYe9LR2LVc6xsr6Z1VxEcG
eKUgb2NNuCDVDSiGGEI0SqasMA21dirBG3Ojar+GMRsWLVrW7HMEYWxFxi4/hsAAA93tDskhRzUq
1DaEpE8RMZ/LEQYuVzsY+JE6cw0GeZHE79Ivxlc16CWnCCojBpKYvBtkV3f//mDkD9K7hv/p3sJr
GaIxoW8TVgOP7t39jBTyp02cM2S3S+dxaXob6DJgh0R0lPszM5X+9Y1th2Oet/+MXr49XBA4gUYw
F9j36QnfegnuJ3VKTtXZ8xjIjDYOwmG8vEnygFgkzKpilTJ7VdOJLqHWRZ2S9cVXTc4numgmYCmG
SnEAxrVE6vqPYc34XP+b7gstD0WldetLEDoolNxkdtAjSVntosb3RqHR8mjetzdDjLEUT1LDfH4/
/g8V3rik3zScUl5WfP4niVwExiN3dfz+UdDQg9aCo84SfmCmOChR7aBzW/u6dD2bV7P6ZtZywLyN
12DwxHSYbMt0xgpKKczqsLDx2AFR3F9k8NiqN4JVM698k1E8wCz/oxyJfI2ZAwZ5QaCd8MTQ9uTG
VYo8LdDenxeAYTfxNEZuszY+zf7YmWGvqeNb39PcP9Oqld3229UP5PH9gQNW4a3+++GEIjBqpfYP
DnbOT8MLs3o8jIpCfRQmeUJF1YOXP9prYTmLsJ4dJGaKiiaccPlyj9ByhrAfiyATaechdGdDSn2J
tRD3E4urd6NljAXjcs5q57g6m+zNsPTsTXe3XJuQh6BRLuTB4KbJ8rxt2rwhBik6hPyNDSMFfx82
6BU6hN5sYmiRPex1ICrCaPQFikgkpBBseerQ0r3LDGX5aoCwGCfO/39p7kkbZj/RlIaaKiAo2ZSv
xE1QyC9sU04KuwGkDfD1TrbnTuO2vm4QqqVO5dCg6P3lLH+LBpRyI/FStEeVWA6M7WqjBXfuqD5l
qBT/p81j/UfwZ8f70klA25m6siEEI6i01I9xm0HNpFlDlNLWaT3THAR4MfJ2W2SuaoysZQ6FgEie
XecYEHb0zxqzF9OOryG6nbOb16DQYbdM4b2VmQW1v1AK+W20Cn8be2M1ht21K1Mr+6InkkAT4zRc
b58raVTx40WbcDpXvm+dU7bQWw3KODovTAntsaKYQ6XDhBjA2i4rUcA/R/P1tfD7LArUMp260OxF
YMZTodS1jgMIaxEDwt2IfxhHqqLM/+8Mk3IXBdVyJz5sdLe3txEKoWrAPqNJhMHm/j4JiO2F9bnJ
M/FtBuRgwC9BATXmDJVO0MRA+hpljKTvhwRoaUtLiJt7nskU1a/m9bbp/rzLTgJVyq4XaIy7w+P2
EsrJF9OKSv0endMn6kNtUskqI15ex35DZpl1zUnFLdoPrEbvYJKC6b19B0PFA1pOVOkil5HY3Z+v
l9a4A2f82pq6kmzTVTKwAH58EMLBil9giq5n2aQQ6EHRGajVJRpnFGgGW5tDxelyNT8P494Ksk9q
WwdRuVtTJhfMps+lrIrPvSpLPBUqqg23J4n5KLU6KB4m7PEULsg5ztwiITf3fUFhUN6TkKmHKMns
B9FFSwvlkto8HI+YexHsvyWFbv88n6shk3b4b5B4BwKQyEiYOEKzq2OY5bbX22MxloWjzWcrdv5v
wb05ND1+K/AcYQzkxMZA5v1Njh41EAvF0V+SIO059uIhmM8dJ74hHuc0ekcdTHXxjoPxrK1PjeoJ
YbZlGYgaIGtXlsZCvf7U9DMqNft1yEftUiiAWAIw4rdscs/LWFEJFFWi3avnVKBov3qHQjh8iTgX
eQ9BH9rPzXkU2q6LcTu2MTkVvieE2+pehlccSOlorEsAPEa+lt4nq9lJrvy0F3KWdDYlGoDmh3NY
Ty38vWZVfqmnN1rz1gAV5CWhXpaKiJZG97+wEFcL6p0pkz3LYDj+3AyseSmN1pe5ViwIeK6aXwb1
/PGsZgKp63TvT5EFVf/VKa3hz6i7r8RMFw+Stl0zOMQOMLW/aYEDKqZl3wUu1l+EHDjXUpMYt9jX
jMeVE76K2Zcwy/IeZBaM2DqKZT1zcOQvwTi33BRdQUSzSfXgCzjUs7bRsM1FH5XugfE6/7d1Wq6G
cvtt0xIMtMNe0Bey5N9mKnC8Th9CEQBqFmCmRGBSDKRnABBFTyb5IXakgeGP8kMlPJwVQEYxLXwi
AF6EkVRlxAwBOQKSuEIl1Laiww1RtW+OtpP7eJEoGyLfea8mVDw+7GADpQjQ/f7WUDqRuCsa1u7B
5HVSjeTORr+YItGPYLBXj39XrNhnRXO4HpmrwLFu/snjhkMDuR73lkPNGvA6ZuJ8Tf7WIbFt9sdN
aNxzJPCb38soOf3HFYyKBUj/UCiRuFohvNTpJYqEIERAf70oN9q9bTs+TKFe89V28ZX1YSaEPNgT
JBtvwTmE1PC+tG4STVuYNbXQyOy4eyYBe/JYT2/YIVUPP4Fr4dqSF7J2oa35VtXEhLFrs6TrSDx/
9b3PtiJIMB0MeuiVsZsB0L9HzBvGx5saPu9Ben3PdqoYg6XugLhFQu+93xTVBiU392u3FevtOMRi
6LpMYSi7fpFmNAcDucjhWgmB3QJsvZvXLwKy5OA3dP3VW4385NMOuAx6QZ4JwyqPdLXCG/NqUuxk
XXhOkggnLQct+UPpw/U/Bjs7Gic3B/PtSg0H/o3TeEq9U7vpkrdU1nm8L4iq4ONnT3IB9NYTffdE
oXF6k6HkOUlcoeg8FxlS3uKKl7cKm4Wl4ZYrULnodDubUjY7ew4MqF1hqcV8A2Rx+qBfR0Z8nQvz
rJE6IWgoPGPVRcOX7qC/fJJNf10YdfxM6x4lwyK2z4nzfdK8OZZEt34wxqgCHON994pwYrcUg4fq
dSBzq7DEMkyP7q54yfrqQH4iwMsUFx32pasqzPp5RrS0Ww5WEhl6scBBdXBUMTX7OxzhWMPMWX53
NsHkaWEKX39xpOif1gFATQIg+fLwvYRSpwHdYpIA+m5R4xNh3S4IyqPRQVCo0kAEg4s63D4OT18t
YHPa7xBB+Rd4M+fMGyyP92D4IsGK9LNZyAD01ENxMBjMXerifl+Y5x9KZsK7CmLb7vGAdAj3K1cp
NOWWoJQQpm/Y4jNromEoTotlNejDyXBMdYlSvAPAi+IXDTiG3q0FOGoxtYQoDuB5712N6CRgX/T5
ok7zKfTsihNLOM3F4iWiyaU/Jp4a4UF3VeO7Qza+vud0VPmDZx31H6NYPUL90YfCDZW6yY+lkciG
eZN+ipAQIkRNmI8ikiusi20Nz6gCMmuX3ZQAI1zgYZUzZHKUxf6a0RrHe1jKPNeKNkgWinyfFNuo
zHkvytSNQeKTs8c4Tg29iOFWGw5Jjnm5Mdq8tpGcDhMvryNT4/zAcj1zv5t3fln/B/smleqYmeMT
k2ZZitAvWDSIgSqILtCH9Z5Hx3B7w9RrRt7IoQhDUieYs4dtBL8WYl7PRXqxaNVpJUi82WGXXw7r
rtPDYP0wFFe8sGpeRfECWudi3StWlgezCbTFyH2UdIveWscLbNS5cwKuXxiyJQ7TVbT8248pguQF
W/6ThOY0btJrcQmxSsDXodUWkG61hxbvwKE6M+Yip1z7OiK4/Q2Ex4BOV6L4JT7L1/4PSESGyRBe
GYyj3bl9Xy2DexEmgYll3HhgUiDiFUGXYt1A0GJgCu0ZpZ9R9EJZLhrOY6+5UFPbQDTd8UBIWLnQ
RmQuUkw5M7pzwvRoRf21wBI6PxjA7kpdT6R0pKWMEeYtnnh9mn9BFZVeAjMO6CcJ8QK8dgeIGHRe
VMWR1iwehHOnJaTqQUDZSM+sWoWwMC4CLUak5vQiHnSGuyJqQdbgUgf9jxT2ASnuelBswR45v1S4
8hqQ5DUXewD/WS9ReGnkZf5dyF5ftBFmzR4roA5ast9OPGTjVYE4DT6Pb60PPqmkUYxvinKldYWB
mCJs7VtQ1Wxr3hBFepUg7cSNrasPlHcAzngIgJl4Q+A6bK+3r2MYnVxOTCDu90IcJPIAUvw5zAAa
YBJBCjyhN7ThLCUigfFBm2BKP0KGqPou8otQ1v6hqsazPvMCl6AIP+xUZSEICXF4/hY+U+hL44iH
ixTMqHsRyxL6SEz6Dk9q+t557YFOc0OQLnxjxCKARQLOrWDLNOxlsppoOpgg87O9jlknbDrZE6jz
91BjZzfCnV4bx/HYTGmaBidDQUA7kL+7Wloj1+bzO9ziAIg9l4YzoxQ24kx5MqgzxeI16LvNlwLu
chKolvojhzv4YnD5l4NV10+kpjNiPN1RfwMSzwBbq4kanLfCRT669foO03qvZ8lMKGQYV8Q2A6LP
7QlBUbQZZAdfK1KQdglFrleoqjBdp3zjVvEkDHjb7Qn6kRcDw6i1QmsFPFCnbIUpDT1c6P3TNOiN
YlPda8VA6yAFU2QBVAF0EJZ7AirsGzXYMvmAvn++uGSB/hK/03bwNtBbvrviqofzkGoNChqcaAXN
B6bvMdU+obY/G6b38sE2ZgZI7q3TuBA3IsDAilA8wFUwdIpHfcmcdRD06MPsrir5T3Icuk6ZMnfT
/fSsT+RkmCjnPtdHjqZTRxH6ikXWiqAgiT6ABiPks4RaxBH3cCesbAYaFAAlumk1mfiTYfAXpfHn
X6UwfJNZ+/m3mzeWos7Q3PCXkRdSpPy7dB6B/IGzDV4Syj8hi/MBhyEGGLTV4c5jHfhjA94s0caL
hGOU4rntB1jD9f/mTRLMV78jCCqRwqAw6NXvlJ+xdqPddGFpCCZTg95brop7hfILGQiYCG5d4OMQ
t/nlNl2derblnxx6IUIBeuRC47YZzhbIG8FI13+cbvtc4IyXZ4rP0ljp/H2BDtu/IT+3X40JS0Fa
sUba2kh7yfhhQcdO5ot03DA+fHek43i4HQZsXjV0k7MYk0/cB9+rV5ZUZmFryF4AZMddvGGgcspw
BMYbEjZrRYbY/2SuDY7sq8BoQVJjmKJUepFyo4VIWKvbqEi//prYaMurRba0fTegJ/5RntbF2Kz7
l8TjbDamiAOUR3OrlTXUyw8dYVZprjdjAzJUHpk4i0WIJv6PfUHyDB0+lx9hSsCDzC1INS8WK4VX
RtpBrjID7T5QLAHvjf4nsex3cAFhChocVb79By2eLpnTD1tojHY41M5hUFwf9t83nX3yMSbuwDOi
/YfnBx+SEVPOOS/4NQXwgtVmPa3yTyacYL0z9NK4+oAxFws94fmS97l1ni2ZZTbVHMoBVXcfO8b6
yfTdqQaezCUXJDMS866bA7UkV+7aQ1crcAV+1AAuYXVo4WtqHQXBpdYUjjrFQgu9e0OTZAcesddj
Wv0VvjpPSgm+T2KCOTb/50+rKvWENppn8aXVduC9N6aexFKV/luOR45sKIsa9mm66lOyfWqyy0S0
2JrY86f3dKlm6EVYf8JAMKfY0tgkbY5bvnFQJNF+x9DH38anK193FdVsDoSzU8ZDHBUR7xtT6EJ0
ePO82/73bMkOcMVwxtEkfdgxbonXqtjNjfBonDAAR9wZuDrq56lsQL01e/rtJsCwL4RbtMp8HIzi
WA+o8MQdfzH+K2DJCAaqg0sdElrvE+nVLStgBv2FHQoILbCvBoVJILxat5DFk+RuB2gDeE0aImZE
HMbgkB16vgGb4P4DgKk810fCmkE1Y6TAjHPv8m2UkAumQernrrc2w7jaDre7oqB1nO1k91ckMDqP
83kLZf5y9WU6t6gnLHwFCHBNJL3ZyBHWDPr9aivvk0jqL4sDMnaFsw34ilT776SvHGZcR7ez4Bor
cout8sClN9vXa6p0jacs/GgmuRFcxpcxC7FnSKSvxILpuXXpHgwjVYEnnxuWTsfYXqiUJarZ01/9
6gzsemm41CKt0KgyWD4dBSp2wUvR79kXBnXhvxNp/DjObbElDSoVPeJYFLtrhJv3X2tfKvid2kdn
oI/o3cWo/GhPi5q0aluMkYAo9Ep7HgQ4O6o3NsC/IHGJNWFEn5jqbz6NFRD9yv+zdO37GqVCbAmN
iBmKbBSnnU+ARYfoM59SeJxKBjK0nAfC02uDNNN9lsDkRFQ2SuRLRW3/b8fBrmQjJJ1v82VkE5yG
0D11kL/RgmtwW7BFLlv/wcel33KuCAeajuN2R1L7wSNz0lpCKOpXrghcZcz26ez87M5FZZicuxMo
wk5YVR9X9VX74LDJzRt1hgPwlwOmnIwVjyymLq6IOxE7VmKsA0bXHyF5oHO68m7tJMdy3ZUvyRAa
gzFbMC7WLXNJbHAkTdp/FjWydElO+sa/rPwk98ToL7LZLQp2o1I/VGXQZHoQrUW6NXAgKm9Ql1zu
KFg6GF1zvI9yyIuQ8RVF8S3cVlVItDkh4gZcsGauycDJdBLGcdv1Y/3L8sEA11c34Yh+hq7rJ+s+
kHmOqzaU1u9xNxwg/+8x9BIJ4HoUu2Gk6cyXwa1O6GCfnOiVDvI2Kc4GqT25PaDNHiFO1DXcixPv
LfExyhFby/XCJcBTj7FwC+LZfCCU8chaEzJ9AcKllbeBRvHp3I7CCezEvQX+DrG1VFy3leTLInJK
nuhYmDGACaYGhRd9yJOy9Op2bQPYpuWJoK43x/OE6yKBaJ2vJCW2+wGxZFqCvvO15ccU067JaK0X
/MxesnMx/o1wW0q/WguvcPnWXEdZKXXGfiF5OzDJaNpe+dU7QyfkVQMxxCDA8/4M/FIASS84cWLj
0hPGgLel00jwESO1BOS5Kzs03SUfL/UvA4dx5g/NR3W6bv9qFRR8H5s0ODXgZNLts5EU6rHvcPsZ
P0BCSF137QyAPFHFJLIfX4hwbNmcljtk/WH+mRDL6mAmAC3o0rzUWAt6gQ2mWQ//jlHcfiRLysU9
fYEa6Ie2A2Ub1tA4pZIUtqXITz21YOHARlhxhKnTqJhIRNFp2qy6aXLG/LAHI3VNkLUBpG+UhtRM
nkFNW5FbTAokvLpu1T82lzMrQtdLy9VFGUnbk3eRh5L9vYFG6NwV3d5t385tmld4XOq9NRmYF7fh
7keSoh7I99p51Suu8DjKk2XGrNRrB1Uinh27Xg0QROuI4Q68Zzh8adlzgF39lpMPT9I0AQKRS/12
S0p6H9tJxvdUZYpMP8At+G/siIYJu7bvfNHvX0bnc64ods4ofRzs/220p81CoZOcKKYbobqivZqh
VqHS/KULFCo57fbvsHfU1JZeMPeLKOQjMilvV+4sVkpxLx25fpmH+BWi39TG6my3nq/tIiXfPTfd
A0m6+Tcvls0MQo5zoL/Uxpoo/zQYDn/Ypc/HvyCO8k4xw+lk/W/5zq/F/mX+a4kZab4hif3KjanS
uYRao43bYMAnndTKzEN4bqMZEqRpoG3BMa20KxD5QobL+6hxeqo6j8d0MCHxBYoKicvNz2elP+o5
h2Nm3lHttWkX90bigtb06SmoNEzNaH5XPA7TLp9V7zSHiQCBG/dt5dvWu8RCXMfCPNVodo1RFBkL
u9KurWpQyIQPUDACcxZoys/gZB+TIZpNPch2nPrVZGBgqARQzAcPaByKeWLgMMC+72ELAoWkSDNx
rG8bdi/Eb62sdCvGJ/NxZPJwzT7XVR+Xrcn4zGOTiiUKrGUFmFWDop90mewhaJqIGprsP+BWVkXN
bFwA06vV0o0LDWoNAw2KUlEAlLevPr2sAcPPf/GWXwKOJjEP0AAkRBBTw4TS5KoxzeGo1wlfqFEU
pu8yf+YNh7CIBPOqkdgBeXyVkxNBlLjSdTDvxDwHq6YWaH9vZqV/7c4/uVs8sJy4W0siZdaBVHz+
PY7mF3/jXOMTN+D3mHD8YlkmOCOpDFoeV+wQAFv/QeRqWmvlz00y4PeAdReGUg5ss57xhx9+SEAS
26GJpO5Nxn9aVnL94JTv8iA8AzRd230CTAOiba5d/H+gWkXfCCL26onR8HWuuSuLikHB/EyEgIS9
FHe69ysDK7bZ4OTkUxzuZ1GHJqyZYVJo3Rh2as7bu5DqKMIUeG9yb1SNnUxwNWo0vsrRfuuR6rNC
CAz1Ynx1eAvTsRa14EPnew2jmvaLyIGR7gI6djgb35xj5oH2Ab5dqteLLQKMpfL2RnzO45/RDnPL
LF1kWlR05Ngxnv3PAP9PI1U3lEUsIonPB739y6Jws01OwQs5OKUk8xVsrHw+IVWa3A6pmXuP5DlB
rmjRg2WZRC34qWL8WbxGdPKLOpaH47tSRLUUz+uhaXVEQAm1+6n3d/qdVNH5kphZ4vxWFCIEKdFS
ZHIj9eQ7xFSrL0FPUx6gOWyGiIuG//1JX6fyEyA+AQaYiM2ATnsQIDOKtHajAw25Df9qzdRjlBZP
ebGss79rOn9ID9FHpi2xqH2rN1t+qIJcusfRknA0enR/8PkOYoXzRXxh3eVBxPBGLqVKa8gOGhb8
AlrYvwpLG8WQxOn7KAwPXVEC5p3DAbDL31sau1Mu+FPYoaOpnkmXsAugQPw25QZATIi74HAL3d86
RLYe6tmqN4UmP56Z11Y5Utnz0ZGcXxoUFeuZJOn9L7FullWoBA49dsWwIHZ/3IKn1e9pSA43nL2G
ygKV0QeGmzzVk/wNO7CHiwavucvGj2+SVS539AZE779841jbqCqEMQfacOZVjvWsBVhLYyI5iVNV
vLKEox7bkjAQPx3P2YdYdPPct8iQPM5AZYRIViaSYEM8e6gm0/ys5dQvi7J+iMi2j9JJARYFTPiR
4C3LJYaNGRyLcV4Pnp298opURkZzBpjY9QrRvOYDzfSJxCGrNKnv/wqygMKRrvTY+1Vwak21Nms5
w0MuMQ0LxJXDTATgi+OBhtKKp4dTnrZfny+v7rf4sshOSKr0+dTXUedBR5ZHLnXMI1m0tUq+7HCN
UQnFPAmVCf4WBrKm7NHPo+rHu/29qV4eLEN0L2FnmAbINSn2YAc4Q1GtmB/+5B4ABxHYyEnTvpNh
yHA2reLfq2eQY8xf7F9uswdwNo4Y8VRtNuIAK7po6EPGg7++oEylfmde2fv/1CRhpDq///a5lJH5
i8NgLtJ3xdP2w0Huqbgq0GdN34DiSrKUQIYZPbR4Ea83WcbMEBwpJh6J6J/3NlZHZD+QDy429Uk9
ViKsPd3k+OE0tSxAxN+Bkt0M1Q7fdVfQifa9thOIzWHJdinaPQpYwH9vT0j+9MfQSQRJBvc+2YVQ
JXGaV//hviGRijx6T6m3CNeGdDcaoF2KbkkHXXdmDM+0AaqX29biiehZ0aOcUsYZaLatdfu/92pR
eK6pEC2GAmn+lJrOm3K6U4ZCLLBIOxKvYkWCPDEyc5VygXpToN47AKyVnO22fpMGYI3PQC7TH11c
vEGBUdldcwdUdgeZJSipxkZO0K6K7GD7aCAUbW01XALBHnozaNPeWc/nicDn+uRpALobhddSnHc8
SQWY9V7P4fL9E2Pj6kpAnPAQ2OiZ5hT9wRD5Vh2ZMrX/ruUTauB7F763HT7USUzowne6a+k9jCUp
RXCmF4cJj4TtLN5BdTIumVeMZv+Io0Enzp3v5Hz0yzc3zW36OEZGIpEudCvmAKDtfgnVxlksrJuB
hcg93bp7Ln0nB4bhrnVdXFhXGb5TdY5pzSmZDptXI5m3QGBqflDFhKJ2uDATE0wpeTYUrbU3zdbB
usAJ2LB83OtnTJd7aGtUS/tLT7T8PSYoh7D7nF3F+R+sHC+9UqY6mX5fU+xRhhs7czXUsjlLNaNh
n82F27cEWewZAY98JoFufVCWypymzkN9OkjaaAwcS6e00/DIC7kznVPFLscI4TpGRlBQHwEfGTe4
6m0hDTZD44kQZ2j2/uzMOPOpwJIhcG/BSQ87iH8J6xVjjOdFNqJNfRvyybKQx+sq0KnmXkBx0H4M
EKSI5DwQsSq/5ArIU6XSVsGe/elxISvKyKAZIm0T4eKuuezvoZ3Vgp19p9KBmPquuxfSZ3VB69S+
2jGrnxon7wnUSaD+VXFS26mmIGvNbinzczY93yX3pBQ7D7lc9u8AFuV7BVXrUZSYkWZc9qBRZcoZ
KrFKQhi2ApAMiokL3O9UoYuH+rb8snJnhRPweP6LO4JPnQG/4vo7VS+rUrzjp2dYO73VrmnF4ydX
B3Esc0UiyAJdlCzcVto8EPK9VJw1s72bYOEBdqQCIEyMe7cowxZnUhk6ZdbKg5TnkFqizcHE+pOA
z5Njte+QdrGxLZ0m3OXJA+3ewhhkPNRnENZI+46/d2LZNLkDwbrPTDGtubHJzC7lYJ0XFGbjedI5
OaHius0/9xRqGOXT7K0FP1Lj9Z6Oo6fK4kkAawCDMuoaV1SVT2IzeCdc3a0peXaKkDfHdsRAVsmy
rNOUeMF2tCj5uZH7hODvZ+yQyvnDU+c/uo2PhnF4m7LSt5VyB/AhLQNflr6HU+kXKmSH//wDqwug
86MryGk8PJ+VyPV0tXBgemdlDUkpBuH1HEiJsCD9usa2X0qzN9gn7EQdHGRseNfevNp14gblJtn7
lcSA3WspI2+Ff2DmF/8INHzfOpDOD8gGByrnqEqliMbFBxqFb6cY4s6HG+xJxO9G9+CK4clZRaEU
jVYxhZc5VbE2ulQXm7KnJOfS/HLP3/8A80RzDxv1xN1LV7cFNXpp6NbfSIblD9A8S38LCnZ2mQlC
rKczb5rtC+ibp/z8suptQQFr906xk6qxLBihH9Nwgn+TxYV3KxOepchpaLqOG2IZ+xkZpq6XyPQv
ANccCZKlyNLW0HnhEaeNi/lYQsNSyeXgvGUu6v9nI2271llch6bnE6UkVz20YNbZMXHSPmSG4AAv
L48FYWrF8Y6twVcKK727O2bxMzER1jxMJzRo8UY3faZwri4r4D1088LHMJVU3JRu0WRbmlkvnQdZ
+XjL8akynw80FdrHiDMVWwFUlAAqp6tqEk3x3UyxDSLmzuf87+JWGjMq6N0EPVHrdcK7lyEud0jw
rTLoOisxa+hcPtPoasCjenL+2opLConqny2OXi6R2/IxZ/btOgPTiglznYPg2Y7DRcoi9nV7Kvti
SHMpIjS/Z8fHcw+ugAPVk5kKe6bpYSfkYPPUPFPLaTFD7cEe+VvZsMMWLsVHEVi6cXnw3FwnXq7V
dpi87DK0NKEVHtNrCOn7iK6VSs6x5z/NdWizVfWmKkyEg+ALoKAvy+wTeMtIquS61d1VdPD67FTK
kh0v2EE/dRXjdDsERAFjxzADuLOPcNBoU7IBpcUwIKcCnb2DIZsL8j+qD0FacgDAgYtA+lXnCWhl
ioGeRvOOTzdNQT+0SX0dX9UlyccUWvDBBY9BPZoT2/6GtCPIjuRu2VD9Lo23KHmXUe01CK2/0veE
PaPJgRyFt4ahbm4yVVi6OxrDoD7+YD28TpX2w0mbpQCQeckPAgcwDuzj0ocB8YbDfWQ/O3xBhO3I
P5uVZqKEvmph1EgLe46h6DSu/T4cRVUhdIRSz7PnDCF4F35CwyfyzCmEE5GXF654ek6qjDIxm7rm
ELx1co8RLei24wva674vnzHF5AnYK7lHoruMIcAuWy/jiFsNzkgrAt9Vc30aSf9GmkswO/blYqC/
19q+il6179FDkAn8hGe/EFJWLH6IjKTKfzg3NDUIHqmHGB05SYEvjh4XchD7NKazNheiNKpoVpIC
4vcw/RZaIj86a3gLVdXXlpXzLrKiPB4NYzv2xxAh8j1Cr/vJN/KqmRgJsf712/9ycjOXcdhLeWmH
DxXNc5qX3mUj4SZQF+NGX0ZbE04qowUIcbO+gwH3adiCCFivmcJ7rM276fyFeApIy8ReUh8UFetr
vGfDRqplbpJhO9/DuEEpcsg1RZdap4lauafMx3hTh7nuSFa+NSmjLacBZQEHQYZ4gwzGKPfAwrbH
YFRscW9/21P7J5Zf220ILOJ9mQ8AV6RPhfA4Yh47E25K+1szvsCb48Xk17qkD0qY56jET7KAUH3v
0M7tfPUkEktXFJ6fNbNQ17PSSJMPH+D6PvavdyGUYXCFnrKy4KgEhIRZDcwT0fIQfZZL+LHxc4Sm
bMXXF6/3ckLY52IR/zZ0AXKsKsODm0YdezzEG46ijMzDJ3LQmJCzkRnODIuo0fUYzIxRFuUlkghn
jhHjs2QnQZwWfn7Eb1wEUvF5ap1Jtre26D0ILDEnUGdDmkGLAc/apimvM83Whp4jr2mWmhMZ3WXS
l4Mc+DqadTHAtf6t6AflVGXZztU6POTOIaZUZnTIr2oZ2FBM9nV5/4xYDQczBd0NAy6nALfXbmy6
axCZoKOGwuK1d0T3lDEbgXplIcZWRam64jwppD62dpLHK36sLwXBIsaK+HUqmVy2+0Uysy1E6tII
qBlIPl0zJsVT5LPa8zBy6unjHBrm76b7XO8jZ3ZlLzL7XkVVSdsqeDfDUw+5Ti7tIkzSj6FDcggO
srrRJVWS9+Y3uzS4H5O0apWYaF/i1DoS/1dlm66Zw+Tknu3q3jhZcb8I5bNmJQyx8iQiolqhYzIs
835BSaO9gvdvVz8T0QKI2mjPVNbFctnMa6I1jm0ryu6vo3lEEL5H9qFbpBFKqhozkrg876XxTYW1
UoOc3ClTxFzxVbOjZwLdtDUbP4I2TGcml+KFchqlvbNzOZTq3o6xXDjRTli9ofalkwwusXjj1HHA
f/ccjwthptfzwS3hnRe3a2s9F3tbS/vphor1QS6+oplgsiZZ68XMX2t5CILVia09lJ+LeWQW9sbt
mqJlnXOoxqELErpeXR+gKq7hKNmsU1jibKtUGnng6hhhOuj81FlTKmshmQWIBInbqqtZkE3jrJwa
rwSrlCSud6f27vWIa2Yy9Qr+AJ3eiI4eHWBBWt6sIqJw09B8rKix2gIZdVY/bO0CoRmhNQk98Igg
uz5uHSWzuq80kYxnG2mERHuVrWB4BVTfE+cpvPXttV9zqfpgtLBx0D9K1RUnbzAdWvhofPIUGJH4
BxVXVXrvhEgPis2FFpSR4KqDL/Iu8EToW0pz9ovblI90QQrUUsigaMpUMPfnv8We7BcsKGZLPrAx
ofP9puYYCL7gqLXb2C2I39UWJ9lJBFKA3tXmOOu7g2vvgyvBhwhMeXFFBw87w8SGdiB4V1XkbweK
EmsndO7W4NrwV1KVnLrdMo6fsumxqQ7/VrhwXTaexuOCVx90j/cdziIpvcIYQTF5G7Pz/du1N4pI
AizvWcOarJA+LminMoZ3atOYcBd+7qOoeWoQADXqLdaL6N9XrKjJ/znPpaTw0FOWk6NfaVxGuWe4
HZ6Zf4UCRAzo1qsnXmZwQwuh4mwzVxmjD3rVj4IsT1wJpxjUEmwPK5Vzu6tHO58qDkoYTFCDW6sM
8i8IcbxUZUd5yFM6lZB6R6BqR6Xm2CiHsj+/ecX0WAibvcgnOPLEVNU6qjI02nS0QQp/mpmdm7MI
h6MsThp3MGqOzUEuRMPF3dd2O9pzbx6Ag7nTo+AjMPIaKp4jvloCgkVWUwWFRtd3BUp0ShTCzRc7
ayp6kfyQqI7JWEESkckHWSwI5CgQh+qtt/hkbC7fva/kKveH3DU69ltJHEf53+wdMmINc9z5plWc
ZcreabMTrk03Gd+QvtWlJrCiowIc5BDSvco7t9+R4Be8s9UYUcfx6YhtmgBDiQn3EiuAMe6+iuZE
7MQB3JNxemO9fTIQWVdiutiqXiBMPv3WtWzQSpaG5gu8tvHl5htB87b7pwZb4x5fk04+/0ic1ObQ
niCcnkqzY56XWJfQO+zV9odbNmOibTSFubNX9YDBzsIh3PT6Kp7zxnSgLJB7dYYS50IGdOEwMrUt
siZfjcYX+WaRSmhYBFt4hUUV5sdHrYCBVjZvZobFN9t68r/95ZL8UAXA+gsMEmdFeL8TIjux2EMk
iMGW+JZ5N43J3LGhP/11A0A8WD7DGQ9wTUbQYyjpRU1eL74J9OzpLqFpAoNBxVZDdvNGXkodF4iT
QHcobVlfTky8peCMNHcfKA5lCfGmfGUlk4zzl7LEFkHj3NwVISe0zJgaqindnHhonwRDDJ4qDhsu
vg6C4huv305rpxZZY6DmQTjxkinmUG4S+Z1OWfWN6ULaNI0/91lK6p2cqUHuXTFb50Kng9id5J2h
HOw7z64G8JD9bQWCQkiu78BuqyMSuMjPw41C9abi1qGP6cEgZFi7gReMWLBsW+MoDHMMW7MNGU+3
C7lrzBCXnI+25BxSG4M8vXlBGs6cBPOTJyIUVQuKJOeB1UUg5ar34iUrXgxd0sZI/2v4lOZIG4bR
87pJ+UFMSp8LJqgecyBnrHBSUW8LNio0IwBQ/rlau5KSZ3BSZmtIXq8RVJ9LAuvvk060fmWacsNx
mcw+DgNr/XHsKNFR87r2akbtfS9x9MoJcyE2lUQyxmyb9uWAUTIqS1mdaVXTtaKz0XSUOEYqK7ty
4Es9ahq/cH9JNxY0X5tTuZ++crJL4pXpJAcP9mbNjCp9IboiGuF8QadzHP2DinKkHVJ2yi1hxRzj
YSqlEM0LQsYzCCwmF1vfuy2F3gShZDW1wsKsdwrK7bPPzfXZqviyTsIRnAcZFYuzgZirx0oXkyPb
ojFscVNSRaYHFn3EFTyqTSucEaw46V88rD3ZkP1mnLdHPaeWruUiQld4g4dHpGZFr3UgszXqwy1X
sJew7nstCR4zRr0MRQxuYHnrIAIQoAYb+a+CCmlySzD0I8YU1aCfbBt8OHoqEzIMMCj1K5p5juta
2dnJID0euvp5rYEvt3Rhi4zHXLSnpEzkuZHhuI0exboydNYJkwk1DXvfkZcyPOY6ck4G2GE5y+te
d7B2rNLUSpF+GoqjqNKdozbf0qdJ+oCdT4stbBJYZ/IBEAQtK44hZJKljEQn//Or3rrCp7puESSY
NUXHPjQo0Z0KC/m+LfQUzwo0qVHa4Sp7DBxLhT+/ixHaBX/bP3eINv8AMM4dM5o0N2PswKlXr/NU
uY4gva1RxUssiuoKXcaLrr6dxFeIKI50KHpDYrHQIfrFHKKKo7xyC94F9AUO2Ba/F50E4shsOn4W
j037j9UgP/EYaW0O8YHuLo0pizDJNkejHLN2PGlG6nFyk4zcWDlxAKfgRbMhiu/ny+R6FFvHGf0M
BVRBk03r+0wgaTcaKdjMYSkij2hor7Wih7chbqXMW16F7ueAMFl+A+q8iDYOE5XsNxMBy1wU/Uia
WMxoLzeXKZ3jtcZ2Mip3DN30CX5aHFPK+G5FEQ6eoR+sScTaO/q/UALaegez/DCFBeRzI8O9xBHn
0NIdXibh2YjFyhAxzKrS6QebF8myCUnH/RXxACMSXzXxP6z20vGgFLEhEDcIUuoCq8dL2QucfOwK
BthPquITGKQglm3YTGthfha09tuXrwaVqQhg1wjvV2yW4Bza4SgNVptNlxKPB9aQyYdueLEDcpq2
EC9SZMLQRD2K+rYa4gXksETshkBCgP0NS6bgmt20BZRA1J5bn7ee+KPtGh2lq2abg/X1CYemi9Pg
l1ro99/Fq7bA0xMqFoMCt8BeL5aVf5NKSiH8wfxj1U10FDmq8OR8y7DARI5thJlQ4OxLO0WDmpTH
RU/cAVT42VB1O+mf/IuQo3THifjoipfxZaHuRyn8gnxwUTpdG50VC3r8Alx7slQi55FOYornDYsL
HppseGX59/fwDqFTmC/t/m57QRXss5MfZ7A+kTbYt9E0DvDfWvPYqmy6BQ2c8yA36ZRkebH9aExO
FRn94x1aNj3YGoklS4msFntmZYPVHc0KBYL2+QkM0JjLloOJZeg4mPfixyq/wiNG/mViq1QQi39q
OIxiS2a3XdDPlVfpe5mvtcKx577WHjWAQBnW4ufJhc9Xyz3vbDcu2+2E2Zfql95sHX1elE/v6Q4Q
GWKBSIEkR+5HWezgXcbMFK93N6AP3mAEM7X/7LB3jnWMGjYmRvf4q7ThfqKseacPNCKKM66/SfWi
AV5LBWbSnLaB6ycdhIfgfVLZoOf9+s6WdKubIwOfZC6m8R49OSISdc/GxReVa7B/jfTpXo2ZWGWr
z29ZUiFp1D/bAKkOcmjB3R0kyoyEWxxs9pmavUuavH+Jn3Mk/DSz2v11G6jIQvmmRDMFj6q+rDHS
NSkIdDxE6eXlqyPy7zY/Xe/ddt4CuF57yPtN8zxFZsIo7AoTkje1cRdWaY36u6ZGnoTUmxgrbTd2
fAfU3tZ0i0R3IaSaa3sLSzcdOiH6JHSgJBwDx5d/DqYXuNhqW07Ns4nZfVvlQBPQQ+NPmtdO4FYj
+WXxYIMLegHJp4V6vRRqE16vugIvmOF3NkPQzGBf0JB6hIZSGmyMXIEv4OTs0s/jRz7rtHh4Ucby
VW2XR0f1aUyygW+FhlAR4kp3J+kVlq4jp3GONx1x5IOMdx1O2zmR5OMHW9mAcK1sFENedgC5thbG
LtTcUaKKDXBymuTT8WmEkd3NzN5RIAK9kPS5n/lQweX2mhvO+8Y9+VFpBP24tu0hgDaOBW/RecZN
aawTBjTPHhwNgQgj8sXA59yc9+CI6ACVxb7dNVA4RMngib1vF18F1k9d+h6Ly8bPCMot73eDffHz
FiLKyrC30IN8MTlRW2wKIYZXKnj8Lx7psC6c7esk6RRe6qdSO/OWtHeg4+/Efaon2ObqpN1gAbHX
i/3WyDqJRZUpRN8AiJgpDDOdK32iRiOxkt+irSa94t+KU6NX2TdRd9AwMoh6/gPdy67dtgqv6OaO
lPYqOq+c06U88pnFw7Gigspv8xjs8XvJPzwcP9SeNyISF57Aqtsn1yPgfWzZHxCUelIgIDpxKT3u
PiyA9IdkiOq5z/fOml3BWXggLYwXIA84IomGEiiYFX8QRkzFeI/6CSY2nYc1T+uMJQcKLkOOtY2v
xl09QRNHT0j8a6U4u2FTny8U9FvdRzZDdYSZ4bVafEUokbTHfXOpmfpeaie196BtOzoqgqt7Dz3i
KjH1APigJlxEUBjA+t3WthYb318PzX3azQoFpiVmvoxDA7MDqpAp25LBURUzaHMfG/oXMgFBTNZt
C+Fwub1vO29E9TYio1hxtvYUfS9JYsLmzhrXgB9OliJruhgi+jWjrFOxmUS4PsDgo7PznngXDOlq
yNwXANtpi6GRc2CcvhCPMo682yhKUyOo5b+/uhZANPP74UJOEo0hmuYVuAIDM3B+BzHG3IjffU7A
xa+diWeCoMNEeYIFKjnMT7tFOhhk2u8iJYQg8VB5GmSbu4EGwv/3ASizrSN2HmwL0tz/YJ5Y5Ou8
2GnN8mwgM0Gh3ofsIVwa3Y4NXUl45k+SqE1Idqtgk46eyM9HoD+dn3A24TzYembVa5y4YpHBxQPU
DS2oibw7/WX2pOlxxXWNQmfyInPDRS/KuUjpJOnG1mvz6TZP5Mjzie0GaseJ4TaTSkTsfQyLPKjE
pspjP+7V8tyekLXJ00/s7tGEike8bsN9N/byU6v0O2SYMfd9F/5Qq9JOIuwr7+oXjBUBhwGbazNc
R9aTsU9I5I6a1MpVIbGFHlH6w5MLa4gs/29OC4QpQOuCvMBWIgmUhxYsQZlQf9VBFfViDEXGTRXC
5gQfEz2ZB9+DcQajiI7xaj/96MNgVJoK1q/li4Deqn4vD9e9IWlER2P5u/ocOvsbTIU/XlckPcz9
ACQ04wfJFCnrMp5bOkol2C+nVQt83MBoULSN5RdrvOblVCNEyHV9AJI4kjuNeeAaPyLVjkjMzrDl
Xl6LHdwbzXM7Dr3YwBBvokTqhLqAZFrC8nptDEi1bsfTOf5KrwKg2UxPo9g0UXOqk5t6HfHKGLPi
k6aa45zBNn79P8UpWQou2T5lQb7U23jZMvXzblNwuwKuKHhFrpAtz6Q4mjx3xkEOmC98Zgd7jfuB
xvIhpqzaSSJJ1N27dNRA25UHh55cKnJhYoSt6ET+q5tX8avnAtfP3qr5IXBnPESil933ma8hlFEb
2TytI59N8NTRM33u85k1JMO0L/vrEyCP/GIZUONp59qfq5NyQf2ysMqf/Vm8hGbEi6WvseKxaPaO
dgjyPSrKPkCQ5MoCAwmjtiWvFL6UcNb8wqfkHcyhTJcuo2TaeUIvjsZ0EtDPJbBycg87pkso0KTC
w/7K9tfJtW2YDZUvwjb2kkZTbnJdNiba5LwTZjlawsE5iqunCgacfG9vkUm5VJ3fqv7ShoTJxes8
H0F7VafCelPlwvyN/nSCpQVxYOIAbesiWSlsDqEvhcqzEyeowneGoRjM/tWBK17JW89iMkJ3jWcO
aVle7QMxpL8hMPFg7mbuMICLY+ZKMgVC/57T1zFAEF1DiYlLfT9Nag2vvU4qrZO7U9hVRQJVIRur
OdN85N3lhWqVxRUk+bH9V5Ln+OwJpQkTHlwJ/BKdOVAb1SWKJ9qmg9gXtSSP5cw4aQ6O3YK4WKdH
5QBnGToLO5I2tLTjGwvCtp1Uz1ip55oJt4iaxDPDSrTWpbaHFeuZACzIru8T/rYfeh5TItKSSaLk
p4v6oTi9qOqnwMGX+1Ib0haHYrjDuXHmZu/CgKMRV+D8eOPnUPC5j9x7DLF/aLps7oAvNckIGMXg
pWRYCZ9DfusvE3m5lq640hAzECAK0puIF2FaMvWJlELhzl24FrYZNt9d4Fn+4QLxOG5UHtOl/3xR
fGJEOLqzNFA+HJZHnYwMZdDrwYjyLWP6A68AocZu+vQMug9R/rHrcpYcGtrRWef8NrQh1Id4eiOf
/TtF+i7Y72swK8kF7SpGN02XVXf5/QnXkpou9EEd3KctpdBJ6A3BJUjlXWzow9D/QufxyYBbPEKx
dO+hzpqXIqWLD83PAmOcCMLF4p6VctdgxsDnkeoe3SXWR+W1KkffjrmOEw6ZPRbKBUhNPGmHWlwM
vTKps1M3bS8i09ZbeeTJt9gs4SjsOi4yhYT/Yp7PrMlJWkR/OYkhctuzu/R+V0IHwbQUg4O1RjAW
tOCaf75kyqTJfzfP8G0aUxaxDfHLuKtP884/fEGpoHSxfUzHf7oQ5BMHhLgBGJilmTxGfZb0bcA0
2+xjCdhVSFs7E2KJRzrljGs4rsBktlj7CF3cSqZ2TxKnN+36MTFUM8b0O+nnhsQ26txaNY/Id0bb
+D78BQWwcHNp5HQi7opR3qPpQVjskRHCjK6NfgtmiQlbbS8zN2yzjHl2CI6Zr6efKffaG1GYJmNr
feS68xGieRQnOU/93JrGY5s2qd5+TY5yeOahR4yZbBDWpB0WEJbdy9oVI5pUf6PUPM1JTklYZR+A
E09aWMGFVjw574XLgGs53wmJAeu0dyccGqj551RkLpotgI8o/Hxfm/2Avd6aEOLKmH887ne5Dq/b
bS6s3N9BE8bIeKglmiGTjx/KApLIeo8Lz9lH5flD/BkomEpzha+RKHfIqCsn1nnNXuF5vO5Rk6FE
MierJn+T/8CD7cRXzZ5OVcLxgBEMo2PF6PbS5v6sIKQppmVHg92RciwjcdBvIblVezJfjTZCSx29
dnwvec1h53XJmV8JwaiNe/v0ODgojpc43f4T9LAlqjswQ5msh0baJzsSYpFCIb/5kkbHOJlgqOvQ
ZX3yEh5uhmAkNpeeQQHx0Q5oerzg42VG1ahc7T3Gcmkfsm3oFI8Uk/epv1eAlgVLGVY7Z9oo5OX2
ZNb9rRgshv5+4d2AjNyVlSE24ElK4Rk2MiSGTsD8QPt0j0S97zNBzANWeJ6LhkygVwmx75iGmnFD
cf5naspYJpXVfUKmigbFhCSsl1A4kCa8x9IBLY/QnqtWrxwZ5IoZ0lrqypKGRE8MaRpyiCy5kKGK
T+CAMQD0tr8GUYdkJPLiazv+pXCXadxoeE7jAzHVpoIscb2rw3rqX7Uvlt4/43TY+iR4cC3B2udT
q52t7emLL3c1K2cjnR29IMcXBUn0LK6E+GDj4iML9JmOvz+sZq3uanQud5WW4BvI7TodTltJ3iM6
sy3Xa0j2aJYAIXiZoMK6Daj4c7sdjnMhXkrD6gQYE01nFgiIT8X3AORr/vhvu6pO5vm6997RR0Y5
nMKc69LPgVvrxZAq81H5Hryo2cHHgrNj91VyK5Wff66cwIUYxdDpTDTvRBsZ8Ehi8UPPsZHIOU5b
X3vNbpHz9EjIaWA+WrRTvRcxPC/9r9OwPuAqcYdSwAjtvsjxyMnMtr2nwoEfcvgpVqYtfRyMYqtC
FP2lykIRsKyppaK5R3iRVkcXgyKxpvWlYjrVegADhKYOUFI0bhf1Sjtgq9KXtc0EkzKoKzoWywhO
qoGdkl4DnR1lS/fH02ZjZIBW114FOaaohhRj6C6/TE0871vLr7dBHX9GMjBONrfH+RlDZtClwKD9
zXSeeww9444xGB5/peT2xuUr6YoN66igFCT/9cjspR58k1g3MsyR7x9ABQ2wJvFIGsoa9bbDzS5d
wZ27otzvx/a3g+GwdLBEFRu4nAj0Sndpro5LdCt528Th5Knt8SB5Ik39NNhietz772lDBHT4MS2s
rbnjZ4sdQEQBJnpU3V4DefW+yyO6LYAHqgtTvktDKnbesw5JJ10P30dPt4Nl2W6EXLMbicBfaVwD
ejjJre57irjPYsCYhiWw1qA6+RAnJI+gFYeV3Sbt5tMPm2OwiHUuh1AhkNfq5QWfXq0Erw69MSLS
7ev+5qcpbiGE68DEk6h0eG7BiW44Uy4Qilpn5zm4z+qKcHP1sYNU12mTUpXGFEhK7paEs4ixEjVc
knXmLLy/+t8CzEmswO6p4bMiAON8ySlQ3l8xzSVrhsrdcBN4oqjci5opJLzVzynM1d3/FzQQCdF2
iVGlJoTkgPKqVE7UGwxx/rZaD0YoueGywLcz5wnNIJAwjKVzGtTlC3yFQurZIRgcdzyoqD/dSeS8
R/0GMfYMvqIr4lYdZwtq7+sKy9uXpu6v2IHCNZpCL2jbrs4qMysPyn/2hv+bhfbK3D62R70y+Sn5
SP3xBBY4kjcWOG4SQCI8FQN5zaKqqoP0lBB/Ly7uhh2otOAaqwr9vzfQbyE0l+dHeGPjVaT4Ku3V
Ai3Q9avRtyYNDw91M4dr1VlHb2LWGQWPi58IiYLavspHg7gdvzN6peuGs8SorFCkUX/ts02hUkka
ppS7fmoKIJFTWwKtsqrUWcg8N+m2XRK9Okthc2VYp4WnrAsklCE4879qaRxi8m0p3rdBr9UfVYKt
reUkluzyiUAYJaYx0Q+3I1U3RbJIA01/LLqVVIwvWRRWW6FBBhg0r8YGenjwTP28qbf94F2WhMSs
+o7deY6ebVcGPYgssgIu3/qmZA/V6OT6MtKFqJ46/VpFc34oozqpI/Q2lbR6E7SO5ZDW8d9lhOC3
E6k8BDpe0XrfTPSpqEAva4YcecoChzodcXg1BeF5JEC4bxQo+AHqRPIAvRjo6BxE19DoUCjxXexr
+LtjTpA8KrhX4+NhQIY0aVSTfIrs8l6ux5kVLGxmV0HfjJDLjtz7n6nLcCqLLy4DqeM6my4rMU/X
QlNsk4tIHtJnilIbpS64u5imc+aA39Ngg/Qz5/A1as0gCzIHfOUUIlRm5PYAzUzF2fuLnGC6HI3r
R52spUxr/zeNqKjGBwbBXLPYLAu18EUJ2DS65+Ytu3mmnI3qYt/HVMr7adnhRfZuM4K0Ks+ukrJi
Dltqmcqq0Jd61N4g5ev00G6DH/iAkV6Ux1Uv1/ZvockGubnT4KlNP7QIc5LZrsHKv2zpA9u6JzVL
tzkFtTrLW7X0XmcFXLMEGYKqtTcvTUU7I8WNRjrscY7oRolMqJa40WS6jeHx3UtFi3SIxdqhC5sX
SvPGh4E0pWVWilGKD3DHPH8anFBjGpJIi2TAMJCGj0w/Q/7du7J1ac5pAlf3mUrY6x8YEYcFxinr
v9tzSrrlYKDS6dT6s9FP598Eh5Ui/k4Vz0Oxaq0CtsdYW8vllST/jFXKUGrDE1/DbRfU2rypdc61
UfOM/hmL5GMNLoBI8ElOcTZ4y6A8POOsHl4NWDcjwMEcmTvtaVqjfg2cwAd/hS/b7RMLdiDnrKbw
EH9GoiCO6769VY+pY6qzt9OjHI8ybpLoH2Aes3gwRFKP5EQprFf3WNlyROONMtdJcprDUU+hDrjd
8C1DY8MxjiddIcvc2F5A0Q1C/64vsvHyK8DI70y6nlhFenK8YHmmPgGXJxrdA9BD8v7E2RpgWrHU
obDOxK+wjFCb+FDeHOm5E0NPgOeqyGXYNMTWSeU369LW+A7SZHbTnnFA+J930+XGqaNwcJ5Du31h
WFpyHOC2qhYqY0iVUrcteQ1Snye/RkNIJ0p+/8O+avwSCSOMOw2c+RUnHQm5hVHaBkaIq4g1bzBA
8E6+icAbnL4P6gr+Nt674g+1cHvr/6TqY/EujS7nzWakiOFb47A6jeWh0c3g/nxkmGjIDORw3ec4
nv7A72/fEoarSJj0p2NMazn1JXmWhnXxCZxXZEg1k4DgM44NYdoH5ZFolGC4+ZNlwaF1MkLwRLnw
PwH8JXdfwk49jkJqDi8ol7Rid5dtbD4krHup2SGIjZtZK9HdqmsTnVEX6wSX5/DDcIOgx1FCwVDv
cC01eZWldIniXOeJPJT/Bm1SoivfXOv5NHBVhsfjBHzJhgNK0QeJe4qhzGKyFyo7KSW5r2xKN9aY
qGRJxT4GUbNaLHOtx98WhAvQTE1QFCcfj67Hd6aJt0njumR9Vfac+QehAWREno11JBGl6rGEMarC
/5mNH501bO5+QbDQ5gPWQ6RYe38u5MumQOEUu7HFjJZUz/KM070PDQw5Ns8ygxT6eajQt2NTtb3r
esoYRlof5rZ/UFDsnm75ZQzdZdOvtUSzMwO7Ws7lzGTts0GiaaU9uWN1iusXzkFvmFk3xau694m4
Gb2kUf5rTgKkwhBL4Voh++sNEVMHyxgmPCUg+8PchKFOXkG4+a8O+kXS2qvNjAqGHP6+T2/f4cOI
ADzVZJJSAKvaogAz074HftSLf+o48cn5Pl5evh1ZTCIHuiBAvhcr7vrDwfS9/t+BHYsMJjot+PXH
G35zqAA7vzcd+r2I/P1/FmlqkkrARklok599vzICyiXTIjyQ5dLze2FF7MBSsT7oOrHYfpSAUUE1
Yo89Bvk8XO54eKxJ9Hc3s6n+x1zk2juz3wlRtNcEF/MATqNL2b0XniyFC12CgmxhTDluwXAVYS44
M/nWkofQhAyw9ac0LU/vPk/ouqThiWEP4zc7DNdW6nmCatB5Uy5R2z1DFNKRYgClvllqko85L3BF
Q2Jmdn9c9x2iYKcNI4sKxQP5E945Xiq1Pn8xk8bbTuU3PmPKWxrusv8kipM9nG5c7FGak+hVTBOv
gpv9H08fd4tKiNvmtMrOvXWd4thOaU6T0p3KtkDS7W5hVhtMAE2kiHbWBR2AU/6BRKDE/nArEyLT
DRn5K2z/NWKwx3LhSJJ/Rvd8EKkDkyh9Cnf2EIlF3pHbW1+SNQ1FvVYFgc02JGFmVtULxJ8BXeeD
NzMSMVPjLJ5ZFoEWclMWA+BFIKnItRJ+5PgB1roSw+Tw5++i2PvYRU+/Cfj5bVNPLNqW+SY3rvGb
TYCiaD2svC+dJ0MXVg7LMa25cVyjBW6jdeed7dIjHqbKfp+VN+oOSMKoO6osUi8eOZ/zS6xn8Xde
ykEIjHHiKHIDZqPir6o7m9XVvhYiors0x+5MTVyoZSxMcrv1xh5n00c0P/+54D/lGXDULsNfpe0y
ZAhtylxfJ21ttjj3W77xKy4thIpUQdnzb3mJNb7quP12/iB780j28khWX/wfChu8oJUA/wmGNzJa
xX5G3jvq5i8LVM6fK3D7In36cWza+zLGg7g5SWuEM6WvplVVfPayyGBnzStDwW8FuXBuilRp/Gqy
5K6V52HZsV+nfdeOhkWgyawoKBAxhk4pdEcOVWVL+k3LHRXJ+2NnwSpvNaieRQoz3c987VnkLuuY
mcdaO/EljPGcbHSckjP7kQRswfRLIs5MXufPvJxyVOX6MLJbNq8SBN8NZLFgQLvxOimZBPU+9LKZ
86eY7AoTN+tjxnBxRE8opYKnkIku1LsdRQiCGQzkTyOIm/V7QFmD0OC01bviuD6eXbyteEsf/5MZ
2VH+W3yTmpQZijuz2KnyF27ViCU7/0aEZEEmuHsvNLkWGcUV3Nq7uLqx+Sw5CMKI20YJmb4LcRYD
f0g4NN0bQdC8ElFEJTh6mvc3ifLc8RqvYCjUZrylvtF54Zy57dSuUG+iC23cbmBkDKgvjzaBzR6f
S9pLvFm6LgWLFOtJiu75Qe09Bp1My5QcZOs8uJIvZ1QlEbv+EQmLcZMJWllwMMUmlPBHtRY7eQ6G
kwBM8zdGKnqYA34GUwEnPjrZ9NL7LnuepBTohJpLdPzNtb6FdnvZ4X08ZYYeTcy5heW/7ouVXUWr
DGIrSoBLsvuyVYJBJhHEjMDeuygq4dhGhvlj3ysJVHT5vZ/bAybKHqGoXM6PRTZ9sVETCpO9Acfw
5QUQGCUEvzT4ymNiXbgKB4AXiQC35qtQRON9OkJfWg/fAFhuaKn5yxRkkYAldg3uBxpdIX3bIvSM
pL9EeQ3a9zfBwDFDeFeFzMKoathxv4TvEe20u9F6Yk48PIq6kCuH31hx5g1ibJnnwcNZEk6C2vHW
QIC0nXsGGOGXVJufRwbWHAmFm9Uk9MVbEO7KG3vw/cLg7MjRTas2wvDCUVHu+K0P3kpG2xiv5NqC
7bPitgUi6TaMyZO0N0B/ax0s+KWPU0A/CORZLstGYlvOaCk4G93CWGmHc2JSHD0HjLjI9Wnedu3v
acKx3Az7tVa08bnsPMn8JhQPSb0ipyf5+TNE5GZOVz2yWUshtkFFuUIo2N4AnfoCxcQII6wFcXM8
kEzxzPSOOsl0fYXCaWFq2aGwx7g4IllJEk6xsAkgyfJzo+iLpte8KjhAscTi3kVDSQdz1sT/ovRC
XkgZl2kyLcYd/uJ1WCU7Rnlm55swVUFW4IUZhIO/v3x/SLdqUUzwdpAnGAnxGn+xQtfq/cduoNel
YvZFnoWIV9eHp5h+G/xJeAdF8dqBxIT7DKkY3Y9oeL/5XMv/mgY4kg/Lw7J/PBgJvGyQlpO04RLt
Y1TvkGDZVx/KnOyrovIbpdrHELXx3fnCETugXpayy+h529uwpk/z0tTLs/UUaKhYPcFE+JLGzZ8C
DhhFgQ026pCVGuVyw3A8XHVp0hjqg8Kct8dAUCt5W/ChHD1MtahViqClaixn3XiCMWzY3yy5EzlG
velO53KHYEicAwtLLsZak+8LJNvueNd6vMKPkEoY5+XSC4tmomIZPuUrgCOw9mLqOYiiI0sefuC5
LaMuoJ8fwv9cHySw0iRDQt27aDqAuvwSbixrG2mZ8v80wwmRy3dJPBSw5kLSIJXL5oZOsSY3Xehb
DvngT1Wj4F7X4G+ohscZ3mrF2nwJMo3P5SXiOxCDkTq1sCDYIzcf/BzK57KsnJTavSj0cIB0yLcy
1tGvw1/nY1QqgkoVrVr6s9UNybEVCi5751FSHua8PevDU7oY6iEFntIODdgP9rlMwEt6GV0CkGQa
0weK2zHSsJBe31VkBQqykTddhiXgiQ5RL39808pBPbwa+E6WD50OZoQkeD7ypgAMF5W+CS0XEYk4
Hu4xK1/spPj/jwjRLQ06i/OTFwb/FNjDE8Huf36ST2Qi3B23Mrpy+FCVvrQg6rEMJ+0cf/pIGKNl
YdEDW9KQxsNPp2F8iJtmvrGQBm/D4SidWkbKpr6VNEn0ltKJRcJueq7DK6ZaJ/Dll84q54WhyMYe
SaSTLbrb/ENf4F0Jw7xFdkhPME1kJx6/Z2rc6J5XURQtg/CH/meUmi8Tp4NTBgzMuT4DSW6Ietdl
UCW0VQpd14e/BtVu6cqgcowsmQrHEtdVLm7dn4rxJCKn/P2KMJyAuecaWmkaFNSSRUIfwVFhO332
Ca9qE9yQ1wOiS72DwIEU/1Vsm+oPJ2j2pDWu1mddx/HTcm3VUZLLhUHnOvZBCyzsPMnnOicHIqtu
mBU7iEMYiCevJYmoqD9VGjZtyFEg2qoUJnLxzA46qSZJHMxjMPiiEgcWM3t9cnf3ODo4y/PRGd8v
1v6C8AHI/aAquZsHEbhco5k80f/L2QUATUogBnaraOC13BmOekdijbtuuKneax/t4AQuaPAf02IA
J3kX6TcNtD5RfGqANhP5WWYHGSZqS9s/9hnDMlz+GA5hbEeCHbfQg+GmlI8u3PJf7H72vYMQ8M+T
JeYHKlDIoJTWSgSBN9B2VQIvHEf7/5dFcD9QYY3kPQ6dqbnVxP4xk69AnuuCpsrHVTTQRZeDTNor
PmOCCajKmfGgks0Qfg5RyjJ+H0d+jsRi5O+S6EzI4r6HbUM2HzL510NFWJfFh7rg2c+Cnc1bhdN5
tUOUSk1SY/odJ/kSydWo/cWfTHRS5B2YVSyglFwixYXsJ2fthgRlJaiFx975sWf3ghmMmqpmsJAp
zMKUe46ei+bL23+c0FKXfienjUDkyj+YjfDdi1xqiGTo39mQWN9eChHvJeuK4Vc4oUZy8NJHu6o0
6F97VZsvzGhn8KhlDYDzu1vZVAuUiojWJOyMxnStPQ52XIxOHOXSazPBsh8MnVcE75mYX+Bmg+mf
QLupis7u4zdOeCGKRx3z0geu09NmsUSZj9LelYPfgqKUDGpUciWOCClK3DkD7qpwpvZdWSCBxmDJ
HrPacCTqQ/7bibYyA13sIzh2n1wU4hDX7oce/5r69nFd7YybiYt91eik0iUrmKAYiydYYBys9MDb
7j6KrB+JNs03nY4vFfQZDFfduf+HR7lKeHGPxmXJhVx1sN9dnnK8aLd+s4Zg7JSgP4CHELlxXNYg
Lj7u6d2pfaXXq578xRtwtv8yJ/8xrVfHO7DV1LuoTO4qQuMuWbqakhSVmcOI1ruo1CuyvU/k/JRf
EpvMNUOvU/7fd/uSodWP1okrWHXy+C3HCIrgskjyNf7z8fD6yUeg1LhPYz2b7V15OmqGYBqDikdJ
1rhdy0cntNRqVWlicRFbWTSsTH6skuw2DuLL3Fy2Qc3XVWHVI7rXiQ9ouMKQjC3airjuioWVDP7m
YaZqjkkmsYFQJ4pL3cxiZkSU37UnAnwqYQWNEmefKUy9R/0iJS+zuJcOHDGauNaILWvszQ5wMqb6
jkIt4jzBkCCWL8p+XakP+XhKUblT66XknNS02PPSrv5oPuIu+2ZB2H8V/JrFK1v8k0RNxrZkGg+P
Ve9Jz9K43PbCGIZxCz0HhDfkxfoUWfTA/BJ+wqLsyhqEJoc8DKrH0R0Mofgdx5ogCGatQdZSGu4S
XrbbnekRIOV/ps+24BjCy5o1RCLm8EFgBK9FceOSeOyprfg60SOrRtidGizVGSdt7ZprxKUrcP36
+bHRHudy0TFLD5k/MuEjyZtI1NSekOMuxEwsKCsgGXahz0YMOOLALqz4NeSsQeY6diadWJwGjPob
y3IJYj3gZcz9d/mgSphv+dXBdDKRyZxBAqwrxU+oc5dgYiISQPB067I9tjMUt+qxyvXxSNeAIzZE
WBjoFDpKGiCOpMso4RIXwb0gP4BLxva78oH/RwbhGp3x4tXO5LBr6ao4GGHTGHKvJperBhLufNf1
chQfmE+dIGCOXRugj4KCyM61MueUzKGdJdZLnFwITm+O3VU4t/maDWhE2vTogi1wYd+xg0GvV4dV
PiE42mcRfltQa9R7uxhJvMyrTMtRf5/b/vefBp1yWJxwAeiR9tP87gwJaJOeWn8gSlfqe4Ufo3Xs
GYS+VN0faPvYTlH28eas6/k/O3p0Gmp3pl4Ndq4xI/tBrcv7bZdQ/MuBXHEISRRdaHTXHYlaDfGX
83OA9PhTfJlI4pwqAut1y/MBsEwF0+lmzMP//ilNvv2rDEr+i0MYkaM27tAysIggEncIxWPE/3Va
pf5pEApUasWjFPPpofULl9OdeFkCIdac2DGH8mvlbLH1WMauwyyzcrW8fQfqlfjvvMsaZa+e6ZYX
tlTR/uDRf9rOKkNsLZrqneSvtvSynr/CnZGrlIDiW+wKM0dOo6Bcwoc+RvXWr5NjQO53aFuIRCNN
qSCH4GOpjU5NHdzM3Q1z1lfp2d1yqNdNqZJ9eDfhykyuBlyIQjqLrQkJ9BHgOLU6EoXtQpjIm4AN
tsXHdQUGfH8HWVc4tXugfN4DbVA8HDslO0SMfc7g6Xz92w963Gj+DkMUbv/ZsBJXVxqJ2MzUr9eN
784S7Ft+1X9/LOTRGXCeo0hDgiH78lF2+f3ORkGcUNx9MP1OiytJnLG53V/oJIALMD3T3QKA3C3m
+8ebkcOsUBTOihq3DK90ccpYBhvEsh9WZrs9MPX1b3+4plTfmMMWBeNuaK8nbSvF98w4DGHbodYS
Anljz7Vxgbty2/nT915tUUvzOvLtxYcUm5qS8BAXtSp1+Od8w3HZR4VDb7tvHXLaqnH0RgLA/FpE
aZzrmYtv1tUfG4zCkuDBP71amBE+hqJzfuYeMjkW8TSjDfdjY7WQ1YPAOcwY3WCi9Vp7T1Yz15kl
a9e0PCIJ5I1rcN5MrYvOpzYFGChoM5R8lEgD8TgoB4vNtqI6BXlFL/o5m1bMz+MiD+vo6lM8URir
z8OUhA94eXma8FChJBMW8IQfaNDsDD7DakOR+SV1bpCBfgerrjkp5jRXFTFzj5uzgGy/5vvb1g9l
ikPvL9XqHbesIMlKeYH1yXJh9nsafbKZaW73vHjS/kY4xeO0JJtav27h5pam6PkiLPkh/3KzNLMc
UUwQtKaPlDJJAKpH2cUFI+u4KMFMIxA573nuJ7w+v5lCSnxphfxPFxztWOQAfnTXLS2v1vMRJRoB
Wqp1YXGm1Ne4rCNIXLzRt9P2VvonyHOCupQqfcF3d3R8NaFi88ErAgnp/LjGbXvKlC1Mdfnm8lWr
7L+tXK6v4/v/mUtQv+rS67keKNFoWIkSviDKcdL02E7LhzqIL3ri/DSFCXyFOjt+spJMXGtFLwp0
5oXwHmHJf+u7cMPqtbd3nTiAfLabQjGq8wmog7XQS16rBC4Yx3zcMqJXypQGCR8IiIECHQT5VgLj
9ANVL1a3o2KTs9uqjPBlZi0xgVZNywKMFhiBB/sbrSAd3mMheP5Q+DaBvYOqkA6FmjjgO6+6grTq
59KyqII7Cx6h7gbmSoYWhH7SoYeyq7N7BunrhBezCnXc2bGf3KrzKQH6dpZvOZithyR2VrFEoXjW
WOp/SSulvknpO7E5Z/Hl0waPiUOLQhhF9RuwJT0bnkGbE3Iepq951D8s1TgA4fCkI4+MI/EIza+3
UuphrhS4khCDHzMH4fZmPk7qc4jJMbwEgsspcIcypeC7KOBSVx0NN2JFyiHDe/8nbnrUsq+bF/Tz
e1ui8XkUEdQkDxaO6fFsm1VXAgBZoV9loTV06PRflZgWk47rHxUsj1qG54dC6xZOxBdJq40gSZPR
frIXiHzIDRnCWIldPSGQ9J5OrrqGmQrww+jWAj4pNUCP9h3aCXOMmX21FRrgs0GxBcU4ILO5gqWH
rZ11jISVkR3IU/MS5EMizdy32+Pw6ZtxN+/oXMnt1EA29FZ3t/PGJriwu4qkIKhqc0DU1vPWO0Tt
tL4RCfRf9qnDhfXERwv3ry81/6AfTyK7btHZjSm3rmHo7Q175t+5iXED1ebVbzs7BxMRvEQN2OlB
gojRNUg8uNKsDZfgN3Rw39Zz9yJxtevck2GiezmXHO5ENqkpnW0LhNMVqkM4R+BQZOWiyNPChWQT
ynGZ9ogl72De91NR4KuTOG3giJPsXIhU0/YGO7yyfNrW2jvE03zWD0X5WWngPsyYrwl3wQkpb4yj
o1TqkmsmC/W4rs0cKW7qvcEP5keAf1oC02YwBa916CwlP/exr3Ax8LsWKUb0Ier9dOcETeKtjY+G
PoXWaCKynXqZ0zKmZHE+kI8mOEQajGS4t3j6arN4+gVKUnMDNgnf1rRCji5XW6SwB0Jn75Wq4QiF
zHzBk/haw0/P84JAHRsMsd2Z6/e6g5wN+1psNBQjhQFsyTAoRF3Kkr0hbkovG4tKKp3AYJ9zMu6S
1XEij+7L/U2LxCVDSML74ycUfkojebkBFcifDW4gUk92oJKQBGh/uNnv2MRIxJVYn60buQgva4pr
deuR058T7d/DM3CZgl6kknsDmin6Fk7IKZzgTTrmYUXhTC2D/TsGGIsrl7ZKdrMieTHsNzHOxIhG
DZ10S2LAVT6Av4oHgejUA84tXd0EUe8vmEWRkpFwIRYK3ZEy28jzNsIlvHuJDyuJO8FUh4Ngol8n
v9sYxqzzjUD1zvs479GY79SyDQfAcxapdhXPJxzM7CftqUSU5Ik0UQLrzVvEpS06vBFDtEy/HVD9
vG693vYEzlR+S3xgsKs9gU/HWAXPUKJE0PE54RlKvCGBcpK3Y5fsGg12sfgTGxgVdKzlxuZnGLof
Y/O1hupRBQOsmTdnmByIiQ6GR7tTjnph/DRAM9Eq2qBF+X+OC6mZhp+jmTY54lmh/D8rEc03Jcw1
aIHyghF06UHVEfHNCFh17IsWag2Dbjd20vmMqG8+bfJTHYCcf5YzasPy4OO7wkgLhBHsIUmWc9Um
/jAn44wuzpIEbJ9Ymdqbi79mmx+6XwrCmaVg+Z8ZgyU82ZEpHKtYa51s0zOizDAbhMyziHWlIXuL
0wAwUhMd6EDYkk86ayqn3kWk+BSQhXQsveldX7UCzwl5GIoi4aP9w5pwZpz/VOEumQ3um3cazuNd
d18xtQkd4LdotS7gJ8tTN2aHK2fMzKD4uQJn2h26hgJH0ebnYDtQb2PI2zSYWU2wcnZkqZy4NSTR
fS7VglFfe/QraaL8lnChJGqQe4ZUhfGsP/IhDNW7+UD9rOUbrZD+02h1muoC1U7yrTaTC6QRuh14
pCvA2gpRGDGf5C4XEoK1GKCToH7qokUiYE5kh5g6sUWVcn9pIFoFoJmAemGMiBQPkc0UMJVTwuLe
d+9bgbMUx//OgwqJDWIHWnLMmuW6PEDIhwRGheKStm+r44szuM2jpmBbJ2yUvfxWhPnjEj778LjS
XlrqYrED6KIxzA3sjd6d2dFAcMm7PtFSvb1DKDrPcZ6OhS5lzjAbJPlHtMoeche50lVKfQk17Ggu
EyQpAxEEsRth4efuhU5Nrbp5DvdEZdOtEpMdHfpp3R+W0xR07gd460AtqOfVmeQ75GeIgC5NFAQN
AwFs+P6Gj5azEVBvU1jUuvCcQ9cohqt97O5KwV2ZZgjAYRD0THx8phATU1vDTnDQENY+jo9RMfoX
I75LCCdBlpWpIneHDJ1Rc/49+O02So+422RNzCTV8NI6amMhizU/vsAerU17xT8P6XS0aJMaoldF
lciA0zoTxu8vIOzvomZIwvbOsEiekILr0DTZlRQKKurRzMQ6GZOmvN0dYlzaNOb9rS1//tERucVk
fCL4oKavBkZDB1yyT/ynmga+jO8jqfI0xbB2yiq8jL22JBQbty86PLuRqKSQxVb+C6WUk8O/24FN
TSMbQwgFmmuKb5FFG9c7nh13lnodWSn0UBKER3m2I07LqwvD+GcPTC8CVScd9lyMlz9Y1t8XWHM+
lWdQrtA5HyFs70f5sOCyxh+hjeTedovFuFY5IBlbQbAcA0mXe3NdVVaEhB8C2wmMfP/2vAzy00jJ
l5DuKd+a3cK7Megl+OR/4peBAypCBqUe78Kstw/jx7ckumCf3cO7+3K3g/TcjQCbrCZrlyNhLk8d
0ENkgV55XHs265DZTC8m8sCObzyrVy8dDNcEKjtL/r2CtTvxlZf5dH2CelEGHKaI1kmoHIBD6LSb
fPvnbZrbwvTfUHPiS1+p0TGtWrEptUrvoC8ouDRF0tZornW1WkeY1Iku08L+isFkt7eYHcoCkSMZ
8SIkcq0GdqPR4EwsmceqAP84HSz/TDUhP9FMcNMp8g5KaCkgOXmfQ6Bn6AgHaMBEIdM2q+FneGDM
GlRnkdQrSUkyuu5f8GtnZkzw8+q03h492kKxUB0Y0Aq//T+jePrH20v2JXgjYVBia6C3HfYhG1MW
6aAtfR65e/Z1pBvcVubwZI3wLj8ChcxO08laEHCX+yTE8+QfmwBEMsWCv50bi8qCzFEMqgWQZvOd
qM55P467r27S+UEUlRmS+I13MbpAfzBS4ZBK+DL6/VOpIkE3O/9Gvu4TXO1odLS/gnsazazeLQO2
6/UFjstVyu3P97ACZ4M+d7Bv1HPR0J0YwumqAaj69g03Bt0duZIz+0HPt8MU169PeN+xYNRAVKhF
HWMKS8yDJLkCsTGRGffKUxVDPoW3WPhxiAanUpKmz6u8KrA4edNHFmr0BU7U/D3VMuO+hdF9WB++
4kEATSlzzl6k4/blsi3oX5We4/m8PmG5ZLY1k2iP5KLScOphTS8R54MnBFua78dA5RCB+hlBDY9a
NVPmQ9IwEO38Zaud+TlVIbqefQz5cUMPAkRVhsdzWI6atYNKefP+a0fud8H7W7ttL5lfOHWL1L1Q
5DN7O+oD/tFRB46eQFMOsBZs4lIN1wuo48KgrvWO5l8QnJWgTBfprMpSZDp6rUOB/JoYR94YRsuE
Q0lrzIZGMiSFTUKN3l79+PxVApNphXl3KYTA/WL35sELqqkwMPXDY5KaueRODIj2veodgSZNuH3j
wi7aBjYLnTv30/0N5UO04HwtkpuvaoAKU/1oLyxnt1Fnt9VQmoMb1ir110SLMwy3gZJEmNmdDjtA
y9n2K/fXjq8MrmVWXoiuX5fcB2co9TffJ7ALFgZe683WNg66dpn3q6/mcARm8m/tUBVeWPG+kjfL
gZIpeFqWvmIQBcLJEMdaRmvLz0NLF15Knx1bfapleItCXl2BcYQtjXCZ9w9KVoRECvaqoh181Egz
7F2yhlnj7aG/UPbMKLS7GWtTuhB6gqjT91fyljoLAIQwkIbL0Vozl4M+ZHVpWoIgwyN1I3ujN7RV
rdH4Km1TB5t4hqQCT6ryV+SWy5Nfr9jqzNlX0T1Q/RZerEd2bLVVhn11Hg674rl3f+ZnohekNTo1
3DcDnQrcNaqxTDTW7jZn5MTdThxhpznihMYdAt4arGSjo2/13BM2UdrgJzcAXg9kLyCVldM4o/9B
8mlzr9Ikh4QW+ZADsRRwvM+ouPnSsmGj8ZTSHL0wscpV9vfcjHUDTTyFjr0FWuTuWz2WE5TqQU7L
GPvCWkRo6FiVVBHl0mLxGk8HBFQvXTsrJUT5Paid3fy4qa2DcUBOLHM+DHzJ7k2uKJ8cVHxO9ErM
C59Bptt5Xx1FrWJaBODp47UudS8+ZazuKQk3ViNE5okic8M3ZSQLCkSuWITK2ggVIKhrvv3gdekD
KA4ASmmA9yxFc90Tn3HMFH4uPlFi5txyPNaJfUYJ0sS0kbm+bPbeDFychwTBlqrSTu2bebsKdTVn
wF/DDZ5QPAO6++1L+pWiW+q6qLO2Lm59bgKScRsKq9lfsM/Envg2R8B0RwdKcpx701f9sRUGod11
Evql1+vX7pB0HfHOPasxajMHHXM88zbrFCGBsUWkZJr2Uk7gQF/qMmuwhaDYRDuYrQsilIqUcGPD
Fpp+eKC8wXx8hP5njbWNNQQ5/i8t17/LHeSnqRBPvKjFUzwX0BV4ZTgC5z1xkSC8D3wXVKInY8Z/
nO27carqBz2F2LCehIYQYS/UjIWI1cYyxZXCOpZkWAAIU1N5Nx+k9j2FIOHi01C88KfC6AHN8FIq
7hhrTi4/VRjJZfJ1tD2alNex3S8NkwS34kAhxmeuNJykOjgF5wfIzn/8MzR6hu1zKpVaFkx4UXz3
VWlhB9iuW101tgI5c7JZ5kkz81uI7Bkngaxm6bSspyLQlH7aXyJVhtKx8gy3iUcFu2QwdRRdgBor
lfNi22XM2zP4y9EpPhbhnMtCST0Biw1JL5sVcJsiEcLe8UXNPAhLPiOeaEj7mMwWK24bvLTDsAaY
DSY0mVZdpiY6xO8UxzK/9OOnvOYLjh2xukov2FFz1JCbOrxW9+/3lX5m3spo8+Ive6Wun8lEQk9J
6uPegG9L/a0whS9EWX3GYPBq9bKzaw0wKG+E/6FPFYGyiAzvQpkp7Vq6d+w1dFHy4uSSze0s85GG
NwVUeFiuCUKPy5f6XG+h/no4HIDfEBBWjcPmFdQWEiTL7BE8jbHn2fjfxbJNrhqTWFuBHNIwTk/y
lhAPj38iKWvyPgQjbGnd5QNWT4cRHtZMTcgL1WcO/Wk5BGNyJkCwDDrQMzMkQCxMH4Myyll0xqaw
9FGUhILOBkZvXCx9Q0XmjU6yijXVD1shoBOFgOjywHCYfwfvFRFlrkYboG2bAtf3oonq3EjL+1CS
aSAC2NncDeLd4lsH7+RAaNeWPufzpTnqI/IVI/Oz4x2eAGIzrV4wq1D7FK7bT3Aamd01SB1s4Q/S
/dJdkDvNjA5BRL7ISa83KTC9OYdA7Fs40TWTykJwZ32niz3GFg+WPd/Yj20jaiOTOQWakKf3Ozj8
gw+wh90dVhLHDNfnbiKQaYx2QHwBtOdeBDLkT644dYoCh5PbIlZeEgr82P/pXOrEOu3BNorzeZaX
QIvXXX2wnq2WBsmFRVt7KFX6qW9atFYan4Cqw4bZ5EcUXnGrzuuSXYZQ1KWj8RUorcT9pmAJ1v7h
dhyhxrPlkoDUN3Jvd3J2/FZDJPmipGIIKi5mNk/vgbrNrbAJU/XcfUdECh2Ds3BTtRB/8XlTo2zS
LatC2PMkHdZ/UYZc4acedgs4g5l0c0ri4nd3byhiz2b1ecvrYO1nmM2+sqIw7MXLsu/Nb4IiqQHR
GgOd98dnSpc8aaFfcQNgAPR5ZBefnAOTbIv9jfoniynToxY9qVr3Wg7WFpEk5RGJawFcAkrIwWcq
XiuzB3Vb5b2sGVUWZoAu+jjn1r9UJ0LUjBm8BfAh0CYe36G311SlYIvo+9THTS6LxOeDDdxw8qY5
r52b9uFIvfPKN2aZO6jcbykIkFCGPaT6DAzu+53Pq3bLkWfq4qJkUsT//aneFGEYcRU7TmqgdcoY
j71R2M+hkk8eWlTMklXFDi1o0+J40QPmEbm70GbX36RiLAFs8OZdn6raQA3J/1A0F308w6iiaYAO
a4yHoVaPo8CucnkOBYdINHaJw0hVzufPQ8nrFs2hxB53XjXzAL+bFlRjjiT5IiDVmWvtpKDPtTFA
wMgXPgWUVC+qf0AtYJs9piQcA3LfTZTq52M+g9mISapIsgIVbFikcBNgMXgU8x6ywE8UKUbq8qKU
yKUOy3qgp922/2Ti0VfytelvGX0DjWaeh6uF2oGc4V+dVtbV5HikdmPrmGw5Mpp61FQ3nJ+XJIR7
nZX/TnXoDs5G64L7B2F5pjx/7IzrbCroucR3wBS6LhHbNdCn3DSnRaZ3EB/49SBrTnMQeIK6a4ia
OHnXr21GqQUaI/YX53XMHdZXkTQVaI+wAHho6web1A77qwVqJxDcCnpipY3G293C9oTe4h0TcJUE
HHi0J7EhmunC8WeTxPuJqFZ6StJWorjGyY9g/UqlYj3XlHLkcW5lo2A/kcEgsX+OBrPz0YRe0d1w
+199iBIImjt+l2I5ygeSwg/bh9NsVDM8BWoe1OE1+9qaINk0vaiuMhTvldJruZ7xOuDqFlm6bKKW
ExHG/0CwCoaomIqIuO6B5LAyylKNThgOTJXYpb6T9PwMUP0yN/rsoXtEY+RfXU+k8qvybF4nmYKg
TBQ0GfYNwRjYGtxHso8J9UJrVQ0a60/mybw3ADQw4xWJAWkwj8eS4kHQ5zOWoPu/Aafyo/QsMWT2
AeKy3gEsZ2ESduGXL4zSRxstwzMHCDGHetlqpHEdurkCQIO+EaMYak5nj2Oc5zdI5YjNbKKRyJtt
YdQ6zDrwSJlg5g8bXEBVt8lJEekanIRWmHoo38ckLL9JXBrTpEY8/U3q2LZxJGndDFD5eGuNyEJh
Y7f/NjvKlSsUigzpO5jBS3C/1ys3mU41/QbLYZ4vTnrXDSZkJfVdg0e1WuAZbxEEseINZZ4lBKB+
bqxwUgXjNLTKGRf0JQpi0Y8GOi1aSL7f10lnM4EK+lFpC4cUflsAP93Bs1Z6PyehXdIGB2kkRlmc
Xw6ajs63P5NU18DO6OwzJ7CRMaAT7PwNNZ4wpptZUS6e/KWDMlKqpzcIHcuRTmhcIDjEAIzCEda2
DuFbA+X3Y7zosPNynzrLcjy39tJPDdXzu4HKegMr6ZSsyHdoxCNz+4bH40IE4TMq+ZthDbnVm1dv
hv1MIW9x56WKH14pVHIq7ThMmb+u4mitL5LswBMmp3BVWQ8ZwiuR2/GZnwpYQjnfgef2a6yOIvfL
dGQ0lRl+3r1bQQI/SZcF7tdNezsZF7fFvia39Jgo0XPqFZRa828bu10tVgLpwpZpqpnnx0ByD2Tc
owcHJkPYQTvuCwj3d74LxE4xAeVdSm0jKeBwnCNyRukw0ZCC/5GwJIcVsxvbZFZwnmA5zJNHwRIm
UJ1r2SJF/w4nzPRVW7FxfLdvOlmBKkid43JlnaCtWs1j2LDaHLq0ZvYxQZTlrSBtUO3iiWLApxK7
9pCG/9DewPC7LXjTnpvg5n646D6icuZD9uycytPDTVaY+zaKyV2tMvN+ROHEg2mNdCvypwioq4/v
HZVyjsSjUv/uYoD3tBjg6zSXMXv6xd9MRZECc6r989XmtYzRjtcwJTo7c48wMpA3TosWcv+/j+HM
uq2tnZvAVJbnLbdc7LCnAZgPuLdb5r5BHODh7sV3nbzfoPSZMzbT5aW5Vd9FkAsrd9w2ilZDOHLk
/7nRh/MTWKFA9jY6wjRwvPDnI1iTYiMxOVkSu2h2bQBT5yG9cZLRur3jAHByduIgqvsCrJ8W22Ju
fslmsyVUDeRUJJy6in1+oViwxekh+EVx/RXIZLuXi96ZKsd83a8zD9wxF3zZizfT2QgV34icWHKE
nihRZqV/StVSggHlFjZS71YHBsee54m+iESc/DnMLKxfKUyz4PeXzmfwnpC/rtjBtOyTCSaPDRKr
KvnFWm+seAtY3Q5JOC5A1/WPmENvDEaGqKtSBUQyXo4VImfF2yZmLcNXc11+gjIa4IRAoLwEq+I2
wtpIcURbDIBUzWuU4A4ZRLzVZnpqBMeRAnn9liUn3LUy4+s8v3ib2mXDnISZjF5MPsgAyHeHVEcl
1dOLEWo18lxk2Z76lwONPUInlNdrlT2H9l3XdptuBpCKm9haPF9kl/sNUOt1YwAxtgA/hVliKCmI
4YZPgfkRzg2bBasOGZl5/AdHjBvqqqaHqUcZ1y9+aRI22s+CE6qz8f3cC1AMWX0iDeyYl7L5q2K8
DtMw6UVttKlLOU5nOmqAtGyiAJXcJKP26EauT6kMtApz4M/tZtI9MDGyC8JeBMHvmESh+88bl4e9
p+u8JtDraiG6siVzsTxPSfqYNhR40JM9LFIh6oZfR/OY+IOrDSVn7KhLNoT0p/RWTCZvoejQute8
xFOSBJ7NY3tlxKpqXbkrpdCVUVDmUJNVvXjKhac6jbedmnU2oSASXFcivAoYzGQc+3EpjJNd5K+w
IMPAW95Sos/clfT87Wk+UnAR75k74ojjqnTsX5hrSfXYYGDu9mPLTMMbl+Gzj4Qlk7GAVLjBXIr2
CWTfr+Oq37Mz/SpfDtTZtp2jp22cOrzh4ctEUTd1qDvi0qBEmCjlMhak8ZzRoflBBpI0BZ0acz0x
7b8ndBkMozLXPh3NCiw/bvdhswnVQU05VtA0my722z+v7CtG2JWE1nRcSXQVFJUrGWqjid5TQnjU
YwDHleaoZfCrsBiL070hGk1kKx9XMbU9Qy5YaTOV2nEsh8QfcUe9c9EuU8rs46YctDpQPIggvZgV
+Vjdf74Vq4GF9RX+E4/NIQU5k6Pj7auAm5K5Y8T9PEd2JjnW15NUAtzYNKRDhKkyYhTKikFSzfCF
Ooz5hsSlrMPvKwP/i7/OxW9UhVMldns1rU0F4iL6vh0c3GIt9hhLItyDxB6hscT3DlIIIT5St6+V
zYDVg4CjziUdHjEq+Od8OWOlO8UnPjb3eVWMEoO+a8HWy4zQJxkJsxIaQu6wjcHC0VIXQrHICeyl
uliKHVoojFz+iFQxzOJFh2WbFUwNv/ZwpS4rUiCyYF77RH5LkRtwOkszpLchLKgute3urbijF4J4
6hGwVu0TXqi6nFKUMm5wUpL0yOQzvBShQw7kbCR0ieBOKgSw8VA77wqQ6K87tVAXWu6Ni5PfsrB9
SgwmHpAPRnEPkHXlLL/AiaRIeYjeBjAZPHspLmAPJZxDD5NTDfNABUk42rTYa27qxwPNQxB/i5gQ
MhcRh68sN5RBcoV7zQkfvcG3ti5lKOiWiV+aimTW6rT+HgodeLqblIZU5R5ULXpRI7w4Tmu0s33S
fGhqpjjc/aJWLlbr5zTwsa9XCU+VnNHUiu/rDteUsYAL/a4VMfqkKK5T5wOl7eK72fmmNLwFTiRG
6o8Xngmx/tnyd2dmP6iRKXR9YcNBPOgpFKBwAh4L8rgU8LKlQ4+EFNrd2wdSnOEYhKYksc1w1ZOy
Bfu5rPeUE9gjcyYwpSbm+PsA5XbkCdZh+jeafCPInYWtXyFNNM2K3fv02inflXUNnfXJw745OFrA
1RZcoQS51/LFgMJuyAPXzjanew9eN3OJd+bGDMpWBfr6soEWvbCqkNKuk0oHfiGgjV2WCuauQumv
fJYQIPGYr9BqwmEQ8W1eIsyl/6pgpb2ThUnRDauPVH9qGEI/VtcR9EY4VO6swbmLVXeW28hHZWc6
dC4v+Rv5EM3Hf+U9DsJirybjjPxQvSzMfIOKYGftSRvyvsDFNN24kI7XiG1N/2uX4I8RCX1L9zw4
/UYvMaPxffWFgcFCW4IknO0MhnV+7ot8TlU4GtYZigyjcpLxbq2EOd1OcdthQj1ZOHy2qsSoKRCL
+lbGfJWlotAeBb5fFAMvyQ9lqEIONCft+DQQJLH5ZQc+8A14o4tpxqo6NgGw+CBOi3DH0DAg0I0M
Ck8ZQuDC0isubxN+Acy8Sa9y2HHtQAmx6r21PUpII0ozexaoa9N5xWyyYFMwGNGG76AUlFTDItWp
y6TPKTslLn5eCk6IA6g1muICcSbJnGvbn26uJ4cmbIAXEkJlQ8L5TuXgdj8YzIWxtgVAlfIgh2wd
QXWgcFDrQPjDx8pnl47Fooy9ezG8W5OoA11bNf071lJZci/Qft3SpcYx8bsULFoUg2Z+4ZwQfwU0
KbV2T8oGmZYUt18k0Qk2Nj4EM+YIf1VKPG/dyWUhp9tADp6hFvF6Well+NUYFg7MpL11GqVYbHCq
0Y0MvfcL2jFTbyziZDz0uf7j6XjH3r/O5YRG1iwzeC/nOg3xy46KAlPrm5t6G2syphnZgN3vNmFa
3j4LHfyO2sOZcNbQ34ik+H0PXfJgDvUqnXdsuTwOrz0SjXgdBXoGJxcNQ7g1z49MMx1uXTKGe2yZ
IZeaGzcK2yKuUbM63spY2YIuLLCGjIMyqxNj/fTpOAG/5Lhh0cyyn6rjpMQF8jxMDCiPWY1aF+zO
yCrM4hTPCOYJlJ+RWdf1DNzinfszLiHCOFCRVeHh1c98P91sKJLjG6P1AcTTqaYGh92wKIf/AUA3
MZ7YaE9sXOau3baMzdB+SGPE82L+R2aTmz2jDy9CRllY694h6QyQWhzJwQZLF5SU/us60r1vGEQ9
Wr7lwx2N1BJv4SSbfExUJ3hL9CaTB311ZwaATOoEGiD9Of3uUZ2Temu18E+a/ZzAA8LO9NFCDb9D
h2RhFPegQAW0FUBdAGNIbrBWn5TcZWy8gvO9kfpcGMXxmUZRdzlelKCpPP1EcvBfLcRNyowOIyv7
+17TJQLXcNIhf8fSExts+RUXaO5YjIOHjtkp6VQUi5nQ07qQxsHaXEU0PTOXeVn5mID5/C4M6806
Zr4svvCdkApP9O8mcofAnWtrCmduMB/ZzU51KwH/vBgQ/gQAE5cdt7eG7g9+aBGJ1VZb1oDrNUDY
FyUIUULq+8iK4sHmSjeiS1b3dj98NawRf9r0/RNsog6sTZf3VPAQlL71Eesh3c9Nzd3AMcOKuTxI
/Bx0HEHPH3GfaW7xsReELVnquVy4NHcshGFucBLaVfDk79aEI/VJcamEAgj+356ANos08/24hYzp
pTubKTlMOyR6EStTu8STLE/D/P3W1tYjUVQ2Kdrd/HtisZnD66AZnAhjkWlP6RaHMBtRMsjf+B2C
WVN9nE986CSull8NFebyPjGlykscSNl4A90LfN40s3FRj7GK+N7cawjQDkCafzQTkj7+XjXrP7Kf
XvUM05i/QBNnj9uQLjBXwzFriErOKDyjJwMnXwe5rvQ4D1kDnbpWT5sBIRM11ftLEX/cjsK2I4nq
3MlZFz7ND7yfJ/4bwYLWC0qtObAM1CSHiHMfNR/houJA8A3TYeKfo+IREv4tWTwH0jw0j4Ow+BfM
NXbbtG1hPgcIrw2TWfA9cJ1KT1XRv7S8aIHHHVc7b8gcl1JJTH0g1qtCoLKdwPW+BzX22nnkAh2a
yrT+6F4Ghy+U7S0OsjU377BWPrfv50/7icltYhkwtzs+7aDjDI58GvGPYQfChYrK7iL+1bTcfDpf
Mll4j9aIemG52KMH8QPF5/U7d561+rdcZG4Rxt11SuW4Cdc3Gglaut45fncE4xIj/suQdJM63FIe
fGDPbdZ2xMMMs8Wy5GEbku2jmP7UBLBjS37Gu+MvxsEpwNstbZdgONMA/nI5KYZI31jimUFkA4s+
vF4QOLUOydRHk8xf1bACoKPe1AVafTe9mVg10rvT+0G9hU7FDdQkumLlGZY0spC3yVqceqvkS/m9
Xn9LK4i2EIupPMOZzA+Xv02ewUqMiDhI4h4Vk6wt9tJAF5xYWG7dx5V63FmDZDQ9IPWXBgap9Zgj
ZUpKNhYFLoUeozxMU6EKR6yB7DAdaS7QZmSN2vlrZiO/ImAigyRHfnb0+ycFMUnTHJa8Zi+Uu1k0
k59W20rH5w3irBLljQgsqqXd5xHQ41/OX7xPMyNyk9D83bFzue58qV1u1lHLtgyrrMolO9nLfTIO
Io1o1LVxo4a0YQdLfE1Luge0NMjp9n63epD+eKD2XCyrVeL5S5Ep3E6dxe10PLzwjfcK+zXxGAd2
dpIggveK1oV63wyWgiIHiXefbZd1orqb9LYUHaxlflbB0mK3AQ7Lexib0u/+6+OUdMXG6/hB3iWe
+bRdRTdLtarHn+5G+KHF6yqWDYVItPbX90cQVmw4lan40I2Yn9tv4UQEcr63y+hKiXppRxvNfHjC
5N/2rDWgr/53g36RxRcAT8ueLQZlVJg7JoxAujESlCKi4niGsjDbWfGSk2nVK9GCoQje93v3m7zB
kRvwNnhN0ABQbtuqJWtcBHInhhtayKEciG2+l7MQJyboiOVFVut78IisUnSh/zFqeYA/pFaybNyI
MabpRdLQzNtpwRkeS130a/8kQV0iEC6E1aoF9l4ofoMNBf6AXuqxh+77zRD0yDyFA2BZSsog2Lhr
GI6m0kZO9BJBKNsVxXV1MVxGVAeJdWq+AmXsM3xoeUig4/6rj5VXSJWroCjL2/iYtUwUp3lFPqmu
Z1ZlkVnZPQfBqU2ZkmEAcB7WV3Edh1nsRgJy7aN/v+CH2ayiMNyreXLCh8LwUD7tADMWa1VIdrTB
P3P1Yl62wSdvzdZHLDHFSdcHj64H2q23vBgbfUT3+/DtJ7HN1FZN9Lz44MFNesNLeG56jvBHiUBx
2RVqCrE9JFHBaxPW1ElV8PwJncSKPMDDearhmUP599awmEohpbX5g2IinpoFzSQLA9EcD3ctrdHC
Ne2hPCLc4odpq9MAKg0VmuGjwO4QPcu/xIPPJ9JHX9B1opbzcpz9llWIu3rMFzJdthvpzcurHgKS
5JyC2MGXZ1PcUbL1LTLiVWrwuKQ9JntzvJGwUelY/VldpAL7ZokhN+HF6cZ3F4peDwsgNXBZWoub
9kcoJWc6TEbOj8QFXMWwgDC2n+XqwO6n+XRouEShBNoOPSrLEXADGeT262IS/o5ED1Xw9rnkRIph
caOu78zhDUQ7YwJLzmcNXdYY6uyanmIUMhrW/dQBKnauijpZ/9g7fb1hsLgXwdpCLARVNnevK7w2
UOXVCleJL2/d2zRGpOvbC587YH6cvcaqcmF8C6sZgumVexswMGhawQX9hX3/sr9Jml7tnkyHYX0/
EDgM86r+U6AseEeqU7xVZw4Ud+f4HeIozZghRMfHJthUuFr2RbfaWD1ZaLtXAkZ4FlAwh/HW1M9I
4NizjvJBEuRZ7ubXGShdOfJL1gWahMOWMk7y6tXKKNFL2fszmURG6jLWQozw+o84621JR4uqdBql
V4HS1aWDamiqb5qA3aGDwhB1VgDOtNa3Qs4Fw2wH3VIkHrlMeFS4axbTS1jgwIquDQTQa62yrjMC
E3ry2dO2LDTkbzv28qXGRLH4EGKkFrHQwmMIP9NrZLyHwFAab6pN2PqFhZnBCr0BrxetH1pjo4LQ
vrR3EKRiHsi9PrSwz3Yd1kIDZJg7sPZ41kvlDmLGz3v8urS6mAGJrntqBLfXJ8OmsenpVi8j/pSI
zni3BM+xJ2WPNSJHceWnWjMhaewXGkLIduBqcXeOnK0LozXLBCehTw6HNyBd2YPtA017sprr1TVN
Y7eR4nmXSCRdqvgpa8wmv7IqL4kXyHJ4hxXoFsOi/gQUNJu7T5qYQZD6+HuJQ82N76Y8UptAPHD6
/tdlK4KA4bSuG40zJVBtqIPCICzJKpkEfUgY7c8VLej/6hHVNbwUfcyUMg+xxVh5+itKnvIvs391
wlZR5wBtHpGbmBn/ql8/l9QSmGff3GpoDNpMM6/ATcb6EzwYJNn4M6ykPJC8+K/TOIoMqJdoH5Gx
s/K7GgL5xnsqkYbDK+EFxbQrE+i3F9bId7Ygzq/euO/ETyOszPttVKqns2y/kCP0/yOFHJSVYUP+
e7gM6JhwPeyhVG9r2iblh0tC5zkuEIb0lpS8zBWuQEmSGRie02noupLEEAhZ3CEn0z5xuvBlzUwu
lNbDrtp3aUsWq78/63zxO6LzgpNc6tNIc+BKfyFkQqPWFtez/O9YMQxHOAoUtbCmMnq6UdoC48R8
jZaOCYUZmE+LatOrHFRFoE87nKYZpQnkkz2U+yb71ZgQbdKxomkebWqX1f6ITkMWh60ap0eBPz2x
qtHNYgTvPornTy6RKg0JJWJ59Dyrkh/TFRL1W9W3vHh/v8b/adQ+S7O3zKvurd7a0PaejLkSiQHi
gVaCcXEJtsDGu8EnOeXuhSeNdRt47rO5adTVKy3mjUn3rL56OPGZLolS5mqksTkGV8paWS6X9KsR
2ENldOtxDAuzhXO87VQ5bxGlljnxOjmLGQTOJ+3fnCKUjvl7NCp5dbFXyLNn3WkzrRnjabW+hAOR
EwhMgm5dm2diR/LJ7I5THuQ/gFkAqpyOzN1oio8JXttlQR25bLo8HiOdpzvT8bimnJs5+t6xFP2i
H7lS+CaqgM1+hwvGnD9J05BCkEjF/iNVw14+m1SRe8UY9WmvClWTlS4zHXRYO2C0FEjelox2T1PQ
HngZnfUSv9eoQrFtGrO7Pq3FDw5R9ih8xke20qrn6W4i1Hw1MQXKs8QNXwNBPV8L1aIJJnpg7tnq
OtwUlj7DRPgsHSQL5/aUk4wu1VqYRYpcaMuScscTiif+MXcFuLK1Tefp6Ff05SfKqi1JjZji4Ft/
5lqfCNxJ7nwLqR/JpIeYlvOatMtBMjePnVtVjEbVYhDldZxrJ8+hWZifZsMRzxwWUzztijzUSIGl
w3PlOioHadDooYHjCYXmjNAySEOyJhU1tYJ8JFaHh7C68U0r9bVSaUEsuaQvnmG/ZyEsEcGyhEHv
3RSHF53X8IgDiskkvorxpJSqOf7sleMyJSA8dayarshNmbSFjmq+Sw5IFtCUqyhk68qJ/8q0Jhdu
sTvCYVzEuDbXniM6eamIR6QzZZEPRB4/mrsuTHOLlSA/tU1Q8dYLY2uMmmfLdePDu3uM2D7OtkwJ
QWl6/YoyskEDLwIjrkDtOFZHVQya0kEJn4vs0VSBNRB4W4UTv+mKhrlnDLVXjD8cwax3a1leebua
uaFm6J7TxzRcKGKPmVvGgNA+JVlBHwWmENneNC2WuPOV87rglG9qBEmRZvvbzydmLA9cFlHkL2xD
o71vEtIwN5D+Wq+ei6QjUqDfUCoHQmcKbsVKLtsv8d2bhJXuMW8qTYll/uad1NpMbmxu1OJCdBv7
On7mxiTZqiT/yDn/oCd0x6P9oj6p3Zn5XorpRLyIxjf7nunbIAvGtIG21dTGUGQZquimW6SIqtOU
HSc3paZ4qw3/bAanOZrCTSrVW3TGbCd5hwk5ogvY4MHrXYS/awDONDGSHWLdocB3j4lQNYsOxS2j
SARqOYftAY7TUexMyGlYRem7DDeFOyGsa9eYgYXh5wmd1GwbIPc5vg+SCIfNoKQBnDt96T+yUwlj
Tp79w5TAIsw99PggYHn250Hm+l3z9XjprVgiOh084DwemuehhX+vLB9EUIrcrpt0a/L74p8WAfyw
VCSiXzimyCgegC/+LvLzTqqqgaAciDQJ/jMM6jAkq8l6Adyc/HW+vcBgyMJoH6Kt+fy49oIFvweu
TID0RZ9yjFhbrxVD9ugHRlkHbOU8wneBSZya/Grj1eEZVAeJCr94/bKbXJC0QIqJoXcvdHfcMyzg
Pcsh4+0535/1P3EcYKCkbeY4FKgRrxTwwkV9oCVhVCfCWX5cRf7g1KJndOA5lEBv4f2q8z9PY+au
RoYZoaa1eJQ037g3aF2qC+HOL7+5VHIOnfi/n+sdaEhS1yWlFarBbj6sn0NvCqqcyWXdYjLVnM5m
lcvZ/ktBdyk6mJNwfUDPtG8MikRkm8YKXSTIQ3AP0znqoUsqr9uZmVMh6BGcNlahI/ap7O13zXF/
SjRwio1VwASfFWbGzncS3GSfEcBxU7B8YT/+lXtPePjeelll/HP06QQpLE5BN8ZVAjmy2hTX5NX+
nyMnb1esOo026k+uLZQqeqTMqY2w0F7q0XOzT2+tXSyM2xi0EQfSeGDuALaWEx7xJs0krWJUVYLQ
FCOebaXOisEy96hWE4FqFrFVZ+bBKm5IT2/+xnX5dInd59p6dzjKndqjqWZOgqf85FykysNgn06S
MfnphyQnJV2nwOqzo8nFyMbnidGPmAs6AAL78i9mabJMuOC4eQvo9Y0+mFFlfAWJBAhge2Rhru9S
E5wtLNXexiIrMOTVmzvK/Kejx2EEPSsyjcjOz8Va0aYYpCIGRyUg37LvUjbE9mu5cqepAHnAct70
h/LCcw05OD072lwKD9JUBsqikxnBIB0QCr+gOkIbENfe0Zb1D/FB+SIdBKK9iq5lgfUIIx0+ho8z
cwGFka0a2rnxd65DZA9nfhLiEmIUwOsa+3VhdSM/sluMj1AUi27BhQQhBAp4Aj0UxJguguCkh4BO
VUosJ5RkS9+X3vl5pDFpvbbWzyY9gGAiHv3zmV3YJjwZxORoPbtnQwqPc7PMn3ZmBl3Gro4E1ftf
OFjASzj5zhuucufy50QkNlOx2TMRKHsmGDE6GKy2wcqeHOsnpulRIzRLVBalb1ZOg61orAtSZmYQ
fl1MjGsv4AvK8LwEBQxCxx4QcfiBnzXxTIUq0p7oBT8qoq11NgdoKSNpwpLlSVfCNVR+Dwi7ahtN
BHoLYYMyKvXpL1YTecid8C7w5RthJYmN3Qev1kzKziqHflMtykHRqfdqCTcQgZTK9K+mxGMFKGSC
dOq/yAoDOjuO9VRrAwvrdsjKxgDoiQTbrTNGYHhMWM6Skr9kEAKH+sD8D+N8B6DEeyYd8yG90YrV
TYcVz0OqBrxgSa4w7Ns6z1PW6iZByBr3XwMgrRBvF8NU+XuCMbh155GYD7LlqX4s0es7j/mms9+Z
duhIQbdEUGZo6mhkAdi8nq5QY1VNexOkJ5GWw32tCCFVJ+Z3qZw4U/+504AycxhhXHjaBSVduYEt
tHQf5/M6H7rGt6hDGl6g2w04+WOysp08oY6g8Tdyg3XrwWoxxVZFIbIqAYs+0esmJCZ15byuemy3
uz2jSw2MPpATEZa5rUjIi9iBVnv803kTqSPhjxL653qOx5LIVz2k9z9hLy0KZsauiAIyOG9kEP/c
1rOrsR9SRr2MO58TQa6FhZ+EPIDcaA0296A63ZijxDaCW4gC6IVCytwdeEWhXlE+7EuC+veEwd+O
yM/EpreeA+r0NZitW4UsftUqvmGDnH5w9OeoAEV1sBt7TIUYjdztyXG/TDTZPt1Ec37rnDkXPFEW
d4o3mOR2TiHcYy8BHlebS0uXE1Du4DwTq5bxWqzC2b8RryJebq7OidM1sKOoiHAtcjoPpE/41ETD
+khMRB3Z5G2+whUD8ESQeRUa8Xq8WS9VzrK3vyFW11hSIjJVUXEFkb8Z4ECAmWNoheg4Yc5xK1Yi
dy70waq1rHm+QbvZmPu7bjb1KIusNe7Em5Y7z7E2axhp3kESYqQXxFq17ZsqqzULp7WhC8FhH3nk
6HG8MxFYwgc4xhd8KOUHU6OYHGoRI9V4mGhnLXMoMWAhEa50+8IWAACiOGAl6jBNLcQ+4Dxllce8
61O+z2Nm/SETsT1GUtucWutlVkg7mfuzdiQH5zgtjuTsatbr6fKIy2GDD6MtsSZ9ZSgsMP5qNdxC
dD+dLIG+LPiFkNDUSZ3EC5dFHpkGITXvnfDfJwWri5UfgFnnLgp0LM0jPpa5LeY4s80fiunjb7ML
fC32mridDUXoQvvnGorCJDG6Y4at5SyiTeAvkiVs9Ec2dzHa4hagWO6whrFZy/Rp88cRzGp+1/Fz
6XwVBuJaSwRTtA4CqfBiQyUuQRPqKFpUqmGGhpdKLaNTL6JdBU4OLaneq/rAt51K43m/SYp/7eKT
KBuX2iTfuLk12mgou29NfP57QT0Jam+as/dnSuipnvtajzDcSwvWuaYO95ukcmdRCjcfSn/almzS
7qOAZQJ04muUUTG53EE/9LVYCm1QTdgGy2Cp1FXL2c/9Df9I2kuwUwHF+ODV3zprTCPAO0HoclsW
G647ezBgppCo48ZmQhWARIQ2ES2FT33RZKF3JNob5LsGEHJnVk0Q4kWsK2xCacBIkkYL5npQGr29
75R8qqpWcNUQnpbCDHXCGoeL6DggDVAV8t/AMzSqpzacdR58+oh+x1S1H9aGRppKqAEzdA+K0Cjx
36kFuPXRA0q0jqSgVOelqK0Mj9CvpjelOfg2N6Ax/eIfb9xs2C3cVJwbLdExB8b3dzFOIqZuQa16
+aTlVQepzLmHrRrtrNAVAualWZNnXQbAl3nO8OlrIph/P49WUglOQtR1NJshw0tF9+dQqxwVqjnt
XUGqTGrHQshyIcGqBGofc7bWUz2s+ARZ5JG2V+ca5oHv6e/IIkhrSnDkaBg1q6VowFBoa3+Xmvr9
PuQMUo9IvO+Fwe6xOXPQutOqqcQ5jbeAV5FLlUu5c6mn/OI6S9KaUUXLD4gYayghLX5OfFKjpt4G
IHvZXMrCVaahkDc5r8xV4iAX0CIrqASe5domL1mlxgHMzwhD23CusDJeGTvOwte7h32FLBAd+HvC
VzBUrbvdPGwWKzEkory74oKkyrbLfsZwkynpPp4/twpR6/8Bn+0GwEdPOXLzwVLXLS6bEivoWymT
VqdjK8kIo4p5r+2GGtXoVVjL8nLvtkuLQ1pR2I3AdSrrXZLDVwjKMcdtXV98FJV6abL5m1WSoeqL
Slm14VViIZKd0QTSXioaSQ0Zx9D/nDEei/FAlZbxgqXQksdlgS13Tkm/jysI9PifssnnK+ky61Dm
9WGi+tDHG0DmWsbb/vDAqwpXozNupX1h8rFNRKVZf+c/0zBLMa1VsqZK4VEBm36USjpXYTnhOcDU
of7wqtQIjsrf4qANx5OWO5UDFbfUU6MxorJT+r3jdV7KIU8DoCw2Gsj/SFLy5mWGaPgdSh8UBtDK
ohkBbYrgTCVgej0DINRo1Wgcypq6EMarhbuyNX25Bl+z/3UaJB2w1QEAao+8mWNNiskrGIqcPjBI
iI8p3URgacCrUqZRA3oasQoyj2cJI/rdVs3uQfQXQ8kUT/e2UaWp9+BAWlVCivUqmYgnZQgNKYnD
WmUb3dG5ArFhzNRdgxB66B1l1mYEHLXVr0iOylZjyNOQe0rHZHJZsYMScXZXzYZYI0lIPaE+k5qG
IzDICyHhAPk4i0znQAweEtRh1/k686vOr6gP8JrQ90SjTDACptSoOSCfG0pzg/Ogd3HCOsp+sl/0
fgTmw1cZ/6Dcc9OKFYLXFVVDy+GOPQofRajWGqjdU3vVlDxmdVNsEjMkYTQ1g7+X4lp71wh8McQG
v29zdq2ZYXMMSan9oxkSnGLT7fWlDgnZIxHPZ/ootFtcIh37piVaxSDsPm56v44/iJt9VXGM+Nh0
kawqLDen6ZBLmEyeebfHcWca20u785bFu3SaY7+61ownyMazPdhM+p68MNwVJXZgVDDupziZJIlK
qW9PFAMFLjQijUbZt+rLBxEQExULsyd4zJrkzzggZskI00zJpEN2ZzYByb09U1TW8/+qXXhpAlZf
+bI3Ry/Zh0EOshOpQ6V0bBQyxz457LXiHuWbCwLyln0qwUiRGFZItRHMbwCPbMgbI7hD+DqZwvd4
OOlLLdMuLvktSH82+iO/6baHDUsL1asKg2iZQ8KLP2V9/F4xmC/rghhb9hCylcNxXRk9iwPpzsHf
pRlmSGq/G/M2cWgAzoNyJgWpDPDbJYM99BP9PkdEfu+fH6GVSpgSbw5WMLVxk1IKwRbTCc90uwcv
MX1Vy213okRL+nwu5ZeERHP+0iS4qJjBnE/WXSDXtLvGcu7P6tFD2Lh9ZIQLArzz9TVOfx9Arlh8
vcMM4uHUFZ5lqXCxZvv7LgrHcj5wJaMQ5J8sGl3LeVrMk0IUP+XIB2pNBPD7WnT/1kPwNhbpV+sq
qvlH/0Y40Q6q9EKDb7fId5DaghDMzmLtKPv/LrMuN4WQyCvq6t/8F4XYNhsA9AEhTQvQVSbBntpQ
6LuC+NVRhcIhIg0dUhvMvM92Bu8HZMYm9PqeYiIBYQAbcGkpT/ChFsC30r7uxs3elXt+e4SK9XFf
AmDTPzkikwOTXmH83rNdLnEJjlEbXMmyFdfvBVCQ7T3Cdk0VRwkW6sNDNno6bfH9zVqmN90a38N9
TVOPM70o1dljeq3qER4mHG6AXVUwyTNmahZoUmcs8b0ikeUIZkGxK8jbH7cuoOmpZ8itP8JLnflj
lMwcFLx0pVfzookwPdB9REr6MQP5pTSHJZ57BY3HVOyYnB+9kp4O0S7lKcbDLPki0P+Uy8rYcKr9
jMNkz0LhMpgDfVDJT5Zs0mUJkQOBl5ZtzkHJdanaAIz8cbEA8LMgDPlJRFfFvq5u834Okyi7IDPn
bAXE5WvVkJFR1yO9xEI25a+4Ymrg9ZAAgoVLJwnKRCu3DjDHCgb9vcI7WKCDN5U71e/ZhfXVAOuG
RvfCQIObxORPN4G3tkMUcZW9fe6MYGFj2G02oK8ChHToDH/NpVQEXYw0hXLAUcLXF2/D+wk/TCYi
eML4ZVN50mzRlhkVytkwuFsnmRoWtQ32I425yPT1099PvlrDdCn7OriZbyBQcbPJrAxXw3pEA5RP
bSistFGTg90ikQPLZeaxYyT5By6HffItdbDhsKAH2lbaZYAMP14FEGhb8X1peCU9kTmHvlGNYZuj
+REq4Qc+sDuIPymSAT/2HZDGv+7X4pna5I7lc4hSC+hN+KyHMbPYWM40AT231EVJQFa+MTKQxhyS
Ve5A3I1A4+gJfVBNkeUMUQ4U5/scHQvKNefLZylxibCobIblJmF2gs4opAN6h7zSGmuZlITzyZ/2
3EGHLTUWIUglV6IJW10VaJU02WpFoNbdopfvslJXz205sILnu83DmGdJJbQgysbs/wysJoYFWqKs
2MN5j2kGnaV0+uQZveLMIQTS3cXdpoZjKxVBZyqu/5NVcj3FnmNBEtMuAZOmpqBsac8E6ALBSinm
Oevr2OS77OZeuSDw0QKSuI7TC6ew6Nn28nQfWlfgMJ7nsHnaASo9L9/oYWqTEUKZVLCox16oDFFq
VjLH5OVdg04qLat2jbMBD3stxZ2K7AdciRhLujSrumrDER8hjgQnn/mdg/xfigWhg/s3LuDqlXK3
DKjHp3QmNzF9QaBGcmPFp0UD9r6IEKSYdKBUazX71Qd9ZhWj9F4J5S11aNZDMYWekucRDxNONYG7
CQIAbKEyigILaQtO5+j4onBVqCo/nt8TucyK8nutUo26zW1lZYThcAu9t/fAaoPH33ENLrSl9I4+
IQ76dZHEk7WzId4K+9M2fGJDpPkmGwNoiA9mJBRhafa+cDUu9W2e15HW3Wri4BNG2nhs/IaSf9v0
R/aIhtHDPQtVbZ6mVDUWIsz2LHg26G8qvyMf/LLvGyY5QaTy9VWP3/nuAbKZ82XYV6fRnOeBbejf
Aj97tG4sUjBPMkg5Q6F5G4XGgHZ0FdlaXV315b5tTWSmjHf256kEACTW/7cKpxS7Jf/qH/mdMsx8
3r8ZOd6eWyBsZ40NGApBLQ7L3Jhky/4Zg6ccgxbOXmQzdng57vd/Z3SY9bFcyFEQwl6BrYPR4uXG
6njzdrPO1xlv9BXExcpJpXiJwWZqHl201uL/gUMlN7ShDPfOv574IzW9jUIF9ReIBkZM3g5rmSUy
OyZG4rgsgFooaxWGRztBArAUwyeKAtYAPGt4JcwNRFZVBHZM4HVqdWfmPKOvJ4KO15OFo8pvv1TV
84DNCHACC8+LDzTGE5EpINjzNZBqxcr30U18+NQ8cRDJh7ztHJZhR9ICj/bMuxzgNbyEFlXKakLD
h11th3xMacInQTGVn2zOcERgcPiJrBfUoR9hgHicfLIVQlOEvQTmGyOrkx1ZXhPmm25cUcY9WOy4
i78NK3bNhCcOZXoiRNy5GUXF96I0MHc31YB8qgAUGI5VwFPS/bfJStrXWhg1k67w4GLKOSNyMRj5
nYoQkATQgym2oEIthaBqrf8AXreqg10gTYb1/L7Dzqd2BeLUT4YZfEfINv1TP5uNh6tvuWGOnDQC
+2/omPA8Rlwt8NiLBVNKGvsD806VL0U5ukXylythnW1GHNFGlAvKpC0Z/GcdNSLNGi3qK8KZ42Fi
zQ6c3FWIRjb5igAT+tO0iGSTbXbGh465KeZ2THjfuf78gQiZU05TRV9Zh1TPauj/L2mTfb0a4Ljs
m4xRl1YesG+smzhJzrnTcaM9OYcD4bZONPSJQeTyfhvFaRgagDmh1/+QIq9v74Emc1BEaGXu3E5C
DqKrU0g8u63QpquQ49dsB/3qq2k6RB2u1IjfoCgGVQWQdHWaqyAs+Sh/fXuGXE6OUTwAdOdJBlFW
GL0XE7A4y9QLP5S3/1MDko4NPmbTBcSGPXJNzLc11YAAAz7dBRSEDp2iDE+9N5kFamaDjwdwDOUf
XXl7pbBp1t/sAjZgLRKABrj+U0yn/Ot5sDuNh3hgggkYHCYrLCVAXj7BBvUUFt9W26p0AqLohS4t
iKeOaj1gA1GVnptbVDcEYsH3qS2Z8g9Rn+LA1XAxcGPjiW+SZi01GBRXp2CseDT6aZrtn0nNzAhp
2/E6VX4DOtgKCR6NdKdIYfTo7Id7rZBXpls53WUBCcUDzkUD0kpyfGUclGey4A1LPeaXGd+DyojF
WMDyzqVW6snU3zd7Rea1dprA5Eu3xfKpNUwTsq1PH/ye5LXzGNVfCy06O82YYfaSPIcXiMTdsacf
C6NiBxFcV2vvvh0Pxd9xifCY4euwW+HY36XqR0FRSlqjnkQVJqfah918RTs3CWDWc8JV54hvxNsr
CjFECihglV+kUTu691qtBLMdtDGBbGEpe1SjvIekMSFpUQJa5Hw0BZ7yXMevwPaTGiameEBYWKXY
50FcaOPzOViu1kFappoDYsN+CL6VHoCzd2+MreLpJTxEUrMXNy15cxqYUfWlfbpSAEfu7BSPYIjY
0xXkJvTSrgH79fCpmddUmHBBNXd01wemHMCQQORRymuQ1atIEHgwJ5NT/92164TtRXpAjy0gtmIp
yKM2v/WHOUksWE04HEUQjemPrajYRZlJKdXgCAE2M+fQkSWVmeT7de9xy7O6iQkbtS+lufSc0pUP
CehGWAM9/LtUBYauyGZ2P5OussyV/AZpjdeD0mCg/aZMm5R671rCruCCkF6INEOydd2MQCdg5zUM
14qSQlCBh0y5a+oqcR2zrnzo4LRuw2xAvdeO02wfmuJlDkRM1P7Onh5O0J+lbbI/LLHYI2JPLrp/
Ui2Ukc3NaGS+4VypFvGGzAWJGpLQYLIcJgRwaPycN4l0j8J10ErueY3HhdbJnjGFNPfAHQHM2xRw
oa6NlGFmEByCrHueM8gF/v6farIvyWOBZIkLniVQJkOFYMlnb+sDxohm4I0Cwsh0av5xQaqKvMz8
GRWvsnduHKmnR6/BK/zxQ3URNgLbmOPpYhSmPU/J/ikTVFDLmHiiKEIEqXQBtSEYjYXxoFU92qfR
OH3IFBM7TAYN4yTxupdxN3t4paWyCcX0GUR3cX4Gf5JZvfXuDeZn+a5pCiLUtuo3mPKftodb6O3/
GA31N2cRkWxtvV6OE3RJiFyiU1ZyA3oSBvi94MwYHQZGzG/gWkG5P9CdvXy3f26h/CDPfFHnmfm8
g5OtYvyeXEb5lh89rtaAE/2WHll1LCZ5h2RBQxNKMDpnGO7KvblmUNFwl4ZAIA8/xBl9yDih/SI5
127HpApp+QMsKAh6uYUrlHFyDClYPJnpTrRbzN3p2NGJSLPbHm1U47tDfJqz0L22CulJgvyFTCCa
dk46Zu9aZyLtpIJmYv7DUe7N8yfE0ywYDuQAQgJYEJ5VX5SeH7gGjioqGSLWJcTjjg1DMJ0/bF2C
vLxXJvIV0jCUJxH3dtBO1DcB/JOysZHoCS1SvrrzDoKLBiWj4JTtt/tEyKvvB78X2wxALt1DG4ay
YNXKDR2pwJrbo8TwC8ZuNUOQILNJB+pZlz4LKfmj2I4S1FO69B3G9du/sMVi63fVlEM45AkkJimk
OvAXoi2zQzJfaFfo9Y23tYwuTBfv6aatlHNNyUDxNPSlPU7TGN77TP1aaYC9IhhuBIiThT7hUdIe
rpwxS8yHufHhd2sc0DXYUl9pUyUiBYlxObz5tnBgbsPJ8duj+j5gROuhboPSMGtS2VICHv46qTDq
zm/3Dl+buJv+j992K4vKRIyysZXnks+neRz/rFbZKDEGi6SEQ3BSSwXd2/vcC49/P1VWsq8g9Bhq
h52TCXBP1aZZQkLjT4cZqxO1bmXkOfvWFy35fQ5QoQOtFGLQIis6hgZPG0H95yggvhQoItnFMOuT
zOr01WTxrczKI5eD/6oeemBiwRIz124/qQPN6S8LqM93Fg0MlU0l9n23IyniGstJHJlAybMnDn02
HC2lE82HIZyfSGc90zpPXTTY+WewnzlFVHR2/FhKWnkyUu8xmLQ2KVB1hoRG5QLYgdOu6b0J9mYN
EE+K07mSJKPCexzB9qbawghFFEC9hb5nMPpispUU+20Fddo90yG1TZh3PD4QtPQfOH0aRT2XYfJq
HXSIoOqe9KqfGcX794UfkRBH86q3MG+x+I36O5fm9eUk75QQs5obF0LO0VRp2fTyrDskHmBsgQvC
3D9a30I6h+6ZUmoOvNfCBcJqtYyHf68ZYQvYJsmGAXH2Wx+z8eLii6PvVCI4CuNU8dF94hdYyyja
xq0yEhDCF5QsO1flZHH1tsRu2kEwGRUbhOxwjqp6aAVna6GqTtjTofn/nKscSgNdYjEgXUtAPkkh
ocVXt2Q81IR5IhXv7ECfScl3jfaS6NjVRFEndhx6iwifeyo3XBMxP+AvGVtdmXPFerISGyh8/Csy
9iLXboMhkJ91GAi6L96lq9FBIdoIchtJ48lm72JgPjxsr8pKHGolMtk+4qZ4G+2CVVJj+YeSDu7c
VWa6rGYCttUQ2xByRM4Rk/S72+72lgbrmQzWb7VZ+vtN142x3oaDsFUrBduhq6xGWFb3iID99qLO
DgcB+nmlrrodr8bLDwzUB2JfznMQwcqqxkHvwoLTjte0q6XSOJWDfgMt0lYxU8gQ5VlB57YR/2Y+
ol6gC5JuLjZpB7nFew/+wtcdYALgyHJs55uoBPoScfBpwH4Xi5UL0PQeORM67ipde6h9IuEFt/m/
386JP6JoiN/jzxYQIe30s6VYp5O2GdBBcf2OnEYcuZgHtXFU/CMyknjo6r8yBYUG6XdrV5SPpMID
gRLY/Tw25tt/os2uqxP0ReBLbDKWv3PhgCmZgU+ZhRoX4hAM3mgkCE8pBrWcHpEdC+AusX3voHQD
ofQVWkqeenNeq/cKNydoGhxheWoCFGbT/UMqI7v+v4OC9lFC8a1kymaVMKTB9IWgJgQF2FtDh5Ip
5TVYHQwr0AC6Lqae6yUTxgnEf1vX782A9zhH2O9p3WAKYoeIvY0glbFGnr+lD+V+yCtANxzMtNLW
Hsb3s9kjZIMOJZrzx1iD0ZJKoMI4pRsgsVW3RfZJUHxsdvVqOIZIyGfG0bwwl5a/bIG08dSsRwb4
Fm5krRfMRAj+cs5JhMV5w0F+xq4TUgwoqTuH37DoNHDRY9P8DIHm82D+Thewj+Gi1Sq6M/HkidVq
txPHZstz4FAOIS8mOscX7Vu/sZxhD3lFUobiiTzJqA7lFGfXFVHLcpk54O+BOhZw+3xBRi1CU7dc
KKnrTBYLcbQWF8Wjol09WldZdnMkWy4iQ5nTMBeA11IHH6rKKnGVnN0+Xmv69TQD+sBSqVdK3Zvy
xXqo8YqmcdF+cLlbUJ16ILJJcLJxhTkaRS68ZL/KxZIhLAYOcfnxxdMupwLQkA7IcSejDQTJBjXm
4aiJMCKKUpakDDPL50HCvAjzn5ks4oRyWuPFOadV5l3BvQ9ek4DvIHE9MGb8/5/jNlEqQhsvvdKw
z563kF+UxbnP5XR711SXZet5V9yLE12Gd+INoFaFU76S+aDueYQ1ZvfUypVKLe0HQzPBHvKuE7Zw
1bnS7e9I+vZZLONk8tgSd2zbljblgdOAM+eUvYSilkcILbUMChnbMOOv81vi5EoxubA5gl8jdUKN
lgdf1nWiV33+g715jMiKQFQ7D5+GGGN6KzPFnXHZea7P/Lpuot2r2CiaWDZ4NyMTNN+hLjD8Ewt6
EuPuAOmCWwKVryMoOTijamKrs7rdkU1eIBiQaUcyQnQJvNCEV3Sj4mTOByMEUgIA3v3Ihbrgq5wX
qJvEZ+p1UhnGs5uPOKH8tRdCx2OILHPSk1IWa9UGP/ozaeXnF1GAuPWzWSoLAmgyBDir76a122Se
i+Ks0GIZteCiWTGActpp3lkY82FVx51NsgtKWL1EPtC+qeKHu9M4dFkwGymLtEe8Thexsz3uwNSt
FizPyWOmyibVPU4aDLgxKFsWMgzfpza3OnSiZquMxFhwXBtgxQKjLHIGbeuZdToo1jRDRhLLBzeX
fn8mnhEVL9nFN5CXr0lDPTkjkhBazUug1lMX4sun298l3e6SJQp+L5y4ObhBEsC1t2FERe7s15oE
Dzkq4Jbzn5T69clAIWVDLRUu3GRg/xyBKV6d1pMoKip75dytkcRHdDCyamu312u06xYvAhk+FjEj
u8/gL8tITUDNaNDNl5jUdTxa6ti/MRTDyCNEXKOhOn3P0Ob7QTCgVyVo4j4UwoTfplnUgTBSSlXZ
ZREB1TTAC6+Y5JvqwwIWi8xYJ2PO091SdSCV7RDAu4kMu0Tpi3Y3KDoN+ieCpqlUH9y1Hbsgw167
cf7PA9/AL5F4rcIw0DUe73tuzWj2eJxvFZUansT0+RZzJtJsKrsbKQcMcTCyKp2Bx4IW98EIX1ed
WJoI4sdE/Xmm1EEm3Yz5+qyT5kQIqKxecb5ZUb8c/Em4pNnN7NWzA3WvkJZihCc1hu00yvRCsVCX
ynsW89LLgFAVu1zpSx+5IB+tc8/zKflkEpr8eV+suvd499mK8MW0enc99OLtyXO0we7i3FdAqQYl
sRs0zfAjE7DO4UX0bfb8B0fq2nzydnz3I1tqE2yMlOUykxn3oP1hoRPxORoYRTuUvpqcfwXhLQNS
ZRGxL7Fs4vzBUr+X4YdoXCiPuyL9rnHFoyZHcDsy0vg44Dez1bgNRzxsTapDonHb5vN2tIa9d0rp
8weQTHwzYVcn+LxuZa7kiIS/kkqcagS4WKrvZzwAhbJiVyuAlw8whoDink4sOp5Jb1o5HhlbM48R
dk7D9uMhWNZ5c3K7s498udone65Ehj6nTEMv4COdOFRetMkOESnhcTJ0RQZ5UzKs4YvgPUBmOl9d
oxwse4cszyLHheUfMRVQB3x8P5Xa7PYtfQcxQK9BG59Uri+lvXgTELjQy1S4zYpBqYREMocAusQS
oG/8fo0xhRxyfbot1XGjIkuSRlOiANsZnBkB+kB48eFA7dtig2txDa5g+2C1FAxhPKYqpuNWktQ0
QKzfFZIuwagGSrMKEl9XGqaci6abflcwqHtWd/fxq3oYWLTBWA2IhN90tgu+8hUTQ4JiKjqbmKNh
BWs8zm0dGheE/NR7/D3PsuGOkbreqb/XLRANpIdM58gkVbrEOZSVrmRbuLOH1SFQkmix6Vs9Aui5
AHp8w6NS8s6gfagLhdcoOFlDLXei4d4QFBEzqQsvw9iTIXM2Tdccm11+Lu2F2HgkkvfMHE+BE1e9
LBgHwF5UDi/Vl1CkNL2ERSMU/kt86iRPVHWSEDeQiYUZ/eupOvLiVkO2V5bUFynvkclEOtBNEiEP
B5yAm4oLfaIhrr93VzympWZKpmNwQav6jzWBUEs4/AxvX0CuK3uppfhlng/6OR4ABSYZgB1e1tcJ
H9cv9V2hVGcbuuT98TtEoAfOjJZasyyrh7DQmV56zPYWtip01/u8YSlDI7Yl2oJ64D3On5/di+0N
ozdODcflzpfwH0SoLNKkvT8h6cjz7OuX8fXerxfB0a1TGLnNoAcxcs8IbuJcsMmCouUiScXPB/cV
PPDJKxTz9RmDuA6ABkcZ/p5+uWB1/QKS5t04FMasd5uqGfvG6mLJV3rmgWKn65IysI7iiXhnsZyK
07SLfCfl23reZjT3I2N2Hqum6ovFc87ABtQjGo6sZjppCxnyRGAYefaZOA/G2TEyEoW1vjqs0aKe
u2O3mHhIi4ApssXNdr5Vkg5kuvNyRD2uFJ+MkL1srZfh3++mgR7XMpYlj5ox+Ls+tXZm5Stu43gQ
KRX6RRy/88M38rwO9TBrVBat/QoWRtNF2LDeKKgpk0im5EuyjBOnECqQbP6cbeIWwu69WXNqHbwK
HNSFVHCIXfc6r95/RvpEraM263f5zTy1JzVnCguSPXybyiV7ZTebezn+adxJ2neOvhZcFM8XgeFC
p98hsCcfPFEm2ZUZV/RqwP1bo1twCWXJapKhWA/aI0pfG3v7NtbvWJYaoTJFSt+hPm6ATpKrRc7F
fr8NSVtKqdrehp4WQzE0+TqnR5rIDu61ILZ1yPKEJFLKeiPsMGmPb6fPhMyEZf/1tblt5K5AvsGR
n/DO+ZOu8idpwHIZEQFR0qSx8GWyl9E6e68KX9Ghzr0TJ2tM6wfnu5gAoDLftN8JvUo8vpvvDcKP
z1ZPzQGNDCPVUPWJpSRIb9ibV72qqIofFSqbq53iu5UqSQBUaVzWdE/EPYeq3MJlFzbNWOiEG5yP
SzrhXKKl1d8okyBmdHnIYA2vNJBY6m447HxhgsmMK7W7fNwoCcE1j+IJQtD+v/oarQLXqSVjLHni
VGr44yvooQ66ZIWVXh5dRFIHBDCTdzM8i86yXrKBmADCaixknrp/J9Im90jZQrNKiU6zQzo2mtyc
J4FYk2ccDSCzz60flcRB3iQpSnwgARi083m/1e4kMy1+z72UK/3viI918Cqg3ZhXCHHOP/McIVyf
8eAqkrIjVjKR3NFBf40Cc/6plhhTn237KkPvAA9kDkNvoW0uIyahjlgHvt2nHsMIYSMhriwZg12N
LUpJLWqPhebA1t8MY9HmYdDkXjuzgBPhA+h0jmIP42OMXtRhPSGohmDksMkgVYgA9gxAhMaYKUcT
kOi9Jme3T+WqJeIBVS33ISDnLClJK6JR/wNAJ4zMc7TSIQn3TmkvaI96EREDq8iOWo5CUIqsHWrm
jlc/EpO/kLMLnPvSRC1LWXiqWZh2BSt+GMbuWp2eipZ53ROHYa9RF9Khi/Ts2Sd9/DsvoyrkW4cZ
Jy1n23ylkpND4rHGl3gyXBcxri8IRM12SrLhgrGN+eFp0oItQOcxypjHlCV9IOMFgqALxh2B/9Wk
F0/9B7L7vdkf8py47Ke0tAgcNoFk4ksUu851fleuoMfle9xc1khUavtbPwhDSh1QTWnFYtZvrtWh
QXYNJ9jokmMCsr0oWOKaCtFBPCGJvCoHhIkvHVU4O1VDZWMAaneiA03Di0B4zZpDFeW095hkaDFn
3SIU/RaDGvbRULANeTMeWB8vKpS2nC26pL+O6zfFQkWI4FJIS+apxp3348lKbYUFXOvtaePpm917
oYvN2CC6aartqEBupRD0/RrWMZPVY5aMj6U01QXSvd5rGAHfYE/HCdx5xw2XcV4k3BOW/AEZPQTw
5bTzq1ISLwJhRVWJ6zLkYQDVbQwdL+xqfUEKXMV9RNKf+ixwFPTxWzgNeb8YfDctK6tKDS1TrHjR
QYND4HoW6tbjBK0y8yLD+niFQLV5b2746Tjiungb0BJcVfyIO7FBgY+GTN7xGtNVkOYnpoSdtNyN
/3PILnbmPVC/B/d79wLl+/TJDY4W+hKaJZSZJTPa97G/AnbIh5qRf1QnGN4EM36bKIyT+f/dp7Zl
B3v65rfrCagWYHCKP2VILgNmBJlvuT+wR8WtyuQcrptcaFe+xNAlOUG5oJXb9igSOcfHjso1riVn
ovUv9Husr8vemQ+iQJsGJV5LB85a8B7V1Tg6w4mFD4IJutFChu0mv2ns6zg2L83XfDzR/LXyYvmH
PH+gelVefHMdIE6jNQm34MNE0K+3v5GOVlmTKyWN4MvIYZLKs70FTE4gQqb6sCfrJ/5YbGnAPP5R
3yzxXazkUpYjVFx2RJq6ly7V12JPCFubgZ2lMnTu8n7hN+b1WToIWvnMJZGAzfPBSpFB4vOwj1kt
x/fTRlGMti/DjWH7rk5XPbPi7A6TJssAeVuaGQV2/Zo6ZDd2tpmdiOtnNWq47u9N5k6caSaAhv2z
FEarpt4rbCCjqa+L0AUQdmwP3f2zAeoSL+BXrNlMIJ56dnhWXKluibNwsXMhsP4CoG7PDh6vQYvK
I8pNeNryex9OTrNqITYbMiwXy8WoFby4foWIWANoZ9AvUYwgdniiQDvrN7qyhHC+N8mQ32qQoiRE
FHy6lpS708bp3Bsim6byNzsvyFJvO0eFLS8GTbW9wjOjoY+lz66NuIjur8OvJn4ENQLcydCYl5y0
kgHrZUy5i8wwWh+dv196fV3E6kUa2q1BqJFcrEQdoIW+2RtGPj/c1X3XANF6RJ+miFek0gZ4KrWX
9C57sOLpEzmFWUf1GQ7YXK9TBjjAVfP376WnsCDccZgB2jaHDioyoA9+Uo0dRYi87MBbI5B1o/S+
xDCWaX8jqgqe8s13rS1EFXpyK/+cyHCLGqdqhVazfgSQ3XbcCOEA3PQNbUmGqD08baJR8jWBYW0F
0tLCJRWsMFCc3jryVUktdd7j88nYbAo1nOdv6dM8tFBfm6ToUeLOcPeXU/tX9tOQhI83qTG3cBfD
kucGC5aW/S41wm7Orx/hK6EzNn4Ouj/M8IRONF9nItw6KO/1pH1LOoytlCCr/mg2rkr4N3UlftQq
bzakaa9sRrmV1OcaNloSZ87VwRlv+ndw2lcD7It7MzuueKvfH2loI1VWGeXY1VScz8QjNQfRGe7p
Bhs1xTqC+DimVtpM/dNIU8vtQh2unFxDmk2hK1LsUadhUAoDH43/6coNby2wF8JIBM80NFqjuHcZ
sPbWwroOyKXxLZCHO6b2c4YyEE5JjvuaEjrn/Jw5LUi1PuQkaYlfT3gexuaIpTgRSc0IgkTmlADs
qQM2ktgxVKGLUxNIUeMkYAE6lud4mblBwbkRoptOJTCT4QSAYjXK7rVdgvQROu+90m+t4oAjmg6F
v5kophdYY5HvHfFfa+9JVt9kFos40S2Ishn4WQvAamXwFZjGAZCHxBHUZE9t7dSDisFhmfbtAsQY
+WCgm5zYYogfCcn5bisaGV1oa26is1tjwMO+Y25zNLyqeTRfXJTxiYgr2ua7uMwVrzn7BL/x66j5
y0IMRuunsNgbHIxh2G/zOZfCOg06CqnKWkqaqnPZ3afjbWK6Wg0v/a6DHSB8qfwQWMT3TC6smybh
7hd92fdVWnzPg8adLx+0Vom+WzGIEdqiR6V2nWkFxtmmP39Sco0iVcZ6pN2yTTW7rvr6J7WaH3+q
6ixfKJVrfa0pD1pAgzU4HJWJEP+P8Ez7Hsw3QXkjk3GLDstzKDvZU8KYOe7YGPtkjOaZWPwJyeda
mNkfgTf4gicB6oqWURu+IXNxktoR/Tyi8HaTjeGndzt9NGiNR1B+rF1Y9a6yyLmseDi2bEAS6m8w
ZML/UCHilctsSCYGhs8SwFVGB7BCK08yT/dP+MpPSZU4Iy9s1HuoBnuiN9+k0dipT1RIs+SmWKwQ
3DK+moIHSPot/PkkVWtuMhYEzSVwuXx1XFFKiSzZRGZWJFi8TYzljyFCCjphdbceyKxkcxuvIbOD
EZ1iLmo8d19o9NI/D/fZGd4L+4OzwfFVf7OOWoiZMjlOlMQzfX3A7DkozKflZ7lAis4jRiVAmF+6
BOSUM8DjRHi1qYDlcJ/bSSac3mJaerMkPv1VUigxQSdoJN/J4jp4uVJpsUF+Gh7tHIgbpD8WT+7M
VIrAMp1bLoCGRwlsFiMF0pAUDm7n1P7A0vtqre4QmdjElgVt3QxVNnO96qNlmiCouV22MmdmAYt5
QcYdq0xOXNHo5rbSmWWC6Ktb4WwX0SSP4aeoUJgQFWr0/m4LSW0sdXQFOJZ3zefuSrAobvaNjc19
YC73xWAelabwnBCewBRpiwYnMNIHZZ54rO1u1NTdEH0R5xrLaTSfhfVZm5VP7I2NaTwDqtkOYkwQ
F83vrBttjB5c5Q2KZUytfRfwp/NweM7GDb3FWbXZkF7QQ5S7bMN2QxytoQq8zSSE/jg/CdtVqaCT
KyZ5ppIWdd6RPDB2w7i3u1zjOvz221eGNzMTPOcfERvTeUFAWttEPA7yPOxqvIlfsR6VzhgSNTi6
15yzAcgIwHB9i+F7Zr45Z2WFnddcfd4YR9MCFjfO86NOtETzEXXMmO6nFPAPdGh/XcOasmlkMJDv
yRvw2KRFvS+ynF7V6N4vYWMczIRyHv0weL/J5f0Wa10p2u00P82f7tPlFJTAjffhTek2kIcdC/MN
smThJy0QC9T6+lfrqyq54DBSdbdCOpD4p5UmB346KJLs2ZmFXZfff5RuDJwU6n4d3neLW17Ygxyc
Ynm9u89wD5P8oJYMc7Iu8IwFciyfyVH5jRagJ85+Ot2B4XB0XGDovfCwTPaos11lbSzN+D/BcUc3
Zu4hyiGioxpZwnh+/v1AGs8FiN6J2nQnbQIHQlxxuSU5v5dFOm0BYxq545Hktdmv+YV1bkoVrwtA
fq8rgONXcZgRVcjp7vZiFV+lpnVxyeYChHnjhxgjZSNknZXJ16vhaSRz63C5CXMECEF16jEerYd7
6wcOt3V7mq8vY6NHE3izeGL+TlqsrWiNBvcNR3sQDdZjLZlaNs6oAj2FeBcgTTN4jYtSE9IcEMd4
QMdFnKsV9qtNYVCNNqQ/9NPwpdzQe6fveN0mAsPIzZBxUzPuyStmTnj8y4frHaKtsqkoN+1ILTck
MSGFYnKjzq5Ak6io1t5CNIaB4N4egp/daiUPgl9HXC9eKyfiCO+/+H3T/kj8izUTu6ZB4VbASKmG
qEoX05zkLMYjkDphfH3FlF+N+GY+JbyqIsU7pz2N39c3u4nrJ5KnecgLwjW/CHm7IMfWoGtqpQ6o
h8VlhsF3oujSQ6R4jGTmxN8OEb5rAH2lDqjFHC4mV83MQ4gglOUoM1lNgn7x+7JEhySoiuZtunbs
RbF3DD0r5/4wortsjfwIPxBiQmnkv+NvbBjqGe0QlXwTbpoEcWk/mFs5OrficrB9btTpRZ9AbyHn
uEIZsR3NuCc1t8IH6HYUBCdKINNLR/2JgAHAmOGdyHMZ24rJQ5DWAgCYt4pZcNgWZedSdlhXEW3A
N0bi7fy4GQoUX1MIcd70EGS9gZ4guHO0nJMUyA98WKgcib0fEClHuvW0sUWp/TDd9BeP3xOfNrTv
nBQ2az2lnwF2/k2HZsN+UBqP3TEecZmv2/UoAQZ2SaZla7E/2I4cWk7scjy3HznnErg1vZP/Eo7L
vGs7Na1QhECyBIuC8JdzgZ/O/HWA1p+i6SWinSy5LshaKItUnz+accFO+S/LbNf/H2gZYiXqan4k
YFkZSR1RfhhH/mD5kLx6DPdbu3LxyaRwH8oQM6pnHVTXmQHqFaLbJATZba4wqfYCGpgPkNxjs2oZ
GtD12vRLqNACJqq7ZpJkLVOKDuDvrqFgwAESrU4hpsn5Hw2UeZ9YC7qMZ0ZfUhaLdP4tG8Sim9I4
BP0anR8o8KPFYku+kbKQp67s506Q2jBz3xdDKtaqPt4KJrJy4E1xbgnHesZ7k3boS/cJRfL+0ZK4
MSPRCHrkb5xnDT6GFNjCEzJlS3vuWHUqjlX1j1+PbMIC15HpRORvNmE4hkt4bNXExTmRm1mWRePl
bt2bupbM9H64wURh5vik7mjgFDyWan6qrXGYehU5f37teu0Fxgkv65rUKgwLBxicIWQ+tUvWyCnp
RaYLT4dyYSq66h6q7VeFjV9IyZhqKJtvVHT67z1ZXzRmt1QPG2VCfenxx/gKj9YL8QJCvFZqUqcm
/l29DS32Y4wcm3o4eFr4Eg7DNmfJbHevM+F7n1zdhP1R3sWfEoAtZG7oiy6IW/QxtS0ZTuAI027D
/Y3l9EgNtXG/S+nTuLpxtSoU6IVn+UExaELGOxvDsJucbsm0SdanSCJoxb5rihvlCeRXeV6chTjQ
AsMQ9R3cca6e7IgpZwS6oqdjPo0ueTizL5HHgQNqbSJjKkBpuPIBQG1KtQ8kco/XG8zRttXgZpgU
+kslHTzcFZW6dYUles18v1ZDmfBTOjvXAGy3P5BotIs6dhWHJ6o+JmTEJVhefpdphgUJsEq8jlQY
GvIq5vZ3lFijaPWsEtWggfutXgfd9eF5zPlxZEEcvdAhVANbo0uYpUzZ/faFg7wOvVnMksZUzx7Y
c7FFVKtj+h4DkxV3evxdg6Elk8+eSVQcSQBBJnHpglete4Sde6LLhj/m1RPkwgzkr6/A83WhDI/V
PHDrAt4lQY4ArTYwiFx4sijm5W6hWfZirfIXpF+Rntm0yArhKVSXMvX5lz+7fkhYu81O0GZ/f3T1
ihKaxxk+JS9UMNyuzxrPMcVsDKQPqqTn3VRpFX05U7kyU7fqclOkO0lby8N1YtGqmtsmcDh/lZLb
GLVWfN+/+CmwqgUMtCsAm0bg46E52hKWjWAj/utligIOkPUgjCjzuSaf35rvgO3PkHhFIvMtsAWy
HIOwvGFXkwPF1Yx8VgxgvXNndOqf9PuTXr3LGcZuh3toZKokM2Q+j7W2ge3fJAsqhf0aW0P2Utgl
6KYKYWYFUZy+wiiIFEOaNwp1AhgpyDUM3HZOhTMq/vERCrCqolriEw2ZqcomhkLVMCzX97u5bViG
AUagg/7G7atQsp84klWisiViL/EKDa2zLvI7hJyxprcWqTzJaoh/Mlbyi4oLgj+9J3jXZiboMZO/
ILhdfuaRibnKKiz34NoaH3GoT9u4qiuutfFQtk3ywL17jOICfiH0O26ztqxEgSNSOyMm8xYSUh1T
7hFPHntjcTZjGNUhklnc2DHBmfEBqG0OHv7CC0lRULyR0uGSMhr0/QKYDonCM3ZCSAoT3zunpTke
la2VqEdxInMz3pXpQhXJwpzSsbCwZRASHEiSVbQMBfKz3/hQh997XigICgnG999AuGDVcXLqwHNF
u1NmAHaeGHXM5DOx115162MrsUNcB069W0pJzmJ9apVdnJ9rahhRx21j/VtMqfsztEh+jdPvqVxU
2FPvbYIPaOpEUJJH3MUUPoSDkjw8jHNnARhtUnQoVwWWgsRiNqk6M/4UVJcAp9skWsota4GFP61j
IX5j8eLb7QLnzMXRewohDNLjOGb63KFxDbvH4H0eRnjeN1xicj/Ri1H0BZxaglr/uVlX9XGAXHcy
CQrvE8rjfGwYSdnSABTb7dZuXmpnA/JoLEoku18wk/ONbccPRK1Spd+vL5v4vnQBJKeNOCUEjmAk
V9danFA+6tUziYCD/F/KsRecS77MbAszt2+bGxvUi7tSZkVnWv/nHl0grGEkdem4KLuGhwZlV9p0
jM8nSTIxWA2vdtJL3L0ctmlColzXM3eWmmmSK9WFYvsflHg+T9dYGze0vBa2oB7oGijXxGj3WgXz
y0kxB4js96pgYup1HVNVFpceFKD/Hxn+oXppqYDgCsQGHcXKqiDEeJ4pqr+2sIUbRRohVdwzJ0hN
6d7M/dRocAjkDL6afGn7FobKMMd9Kpt+DOyjPlNxST6ZZxwFZGR6I8BDYMdKpVnhE0Enz8H/c4Xs
6aEdkWXPxZS1t32aIAv2BWGw/vl5MaUHmVqX5sokGOGs4ULNdZmh+EdIh5uthbPAPnW3IEIdR9/A
jGNrZdqtyfWVRoRxdQQRwdfTMYDEs9a79iyVsmecY1/CzZPNe7wMp7pnftR8iTu1wAt3AgmNd5fZ
wXGc+0eGRDCVs8AdjH0vDdQsfq/BIsoN7t233wmp2/XeHt2gdgkqvNkb6gJlzqntNrxsZG39XR55
8XbdN66igAfoBS+LMHlJb+xDTbnViSLrcgLltQMeAmz/THRxViOnM/GZx0tkHG3m1BAmA29nKyu+
4ASEsQsfN6AXE4OZNLqZycMtqb7kBALMm1YABhWD8gpBUtDZxLHg45h8hETsMmEe+wQlE/JhywFe
InsGNz/vikjk/fZFil5iTBODt/gtP/E3jnPTQJQhn/ulJvbNGXcflb6LFMu9aYrewkWzWLWiJQUL
8Rc5mcWlw2wfCPBWd6apFCn+YpTkdmhllyiGdwtcKMuQE9O2Nn1LBtsogYhArhG0YRBFsB1CXztI
xlpXWXkPyewowmA2/m0JIVMyjQ3OsUitOQ7zadXQ2LrhuhR7ZDoxICiKNpk1yzGmuTH0DA4zUrev
Wag6EvEUWKOlBJybJ7iQ1tLjhHlfftNo1E/ApYQxvybFwniUSzkJ4lNmlidwBl/imkCcdxlNfYhO
fs6zZOiaUC/FQqd6yfxPO5eqtfNc9pFdKwoP86krVW/h+CLgKv5SK0DUmur4epvHdfQG/Y6MVyn+
DITZ4bitH7r2tH59bWqvLerM7OV4qbge2VdTyIPdwkWSP1BpNcya6AQ+7nEQLNRgt+Xk9GKG80Cg
Yt5tHS5+XuDVaKs/zuEpeFlF1hLC9isry/sOE3/5osNA7SNA0khEYReYDBTJ61G3h3yskCfFsI3G
3XYFgdbjULE46n2ttjMkVMkC4bGH+OsCjkXtw/8AGeoqtl2TXo3yProfgTmvW1lyXlqaXP/wD2sn
SUehlQiJrRy4LXUUFlbBXJUPwlu5T1HDFCOPmgbkuQOs3FghsVd7zlN1IwI6qua5gf8ieVS8iakp
khw3I9Lh3Hmg6QmbM+ChK2HQdG18Inl1LgiCRKhzWDPXaHvb5zPx3hAeGyVWZNA2W+TKJt6aBMvr
eOHSR1QKZcHQShb/Hv/x/AEK2Pxw9XwqF0mwUrZ6fmOeOfRb7qgM3ZQ2vpgCz1XpOjTJi5wdSb7A
a8Y8+y/A/Tjle5WNzA9O/7+LvHdBZ+e9hjFteqUZyLBglj6Zl1GsA2z/eEZ0g0VAlqQRTQoiiJPN
g47wwLDZupKWW2pghs96znRa9+c/P6SB5MANdpFyW2FXzvz/mzwnuhZdXIIfkh3J5SBGMs4Def+d
aC6opg2QykiU5H8HuNcY6OHHdMC0l9QMb4QTpntyyoJ+BHrNK9tc4elAxWaYZtCkkbIJ5TlM/KPF
IEymVD0ORtVb7cGXoFC9wv9ToF/0YS2zrkgQEbmZoGO2RADlt2SOqf4+QofBEmqHhl4MHTaUuy1R
vPTRJMdzszgOv+7U6eaLEaLv96OndEhEg6DeU2kf6vIlfT86igYMZydTWuedM1GF/cXms3n1dFhz
UCDzA9dverNRZT21w3+9m8roaBoZimptS7zT3uqGErl6PYohgpiKttw488kADy05aoJ9THaDBlIx
/hNEVecNsYlyW0XZR66+UkyyyklHa6SMWMHj8ZB63GYZvdeOIUpn2KHhJWSh6jbIJIipm1dKw358
UMfsEcebMGpx0fPhVFqOxCTdw/BKu9JmotqJtWDMPQDwdIi/PKlfZFInDBIvxkPN0pxG4GImGYAG
zNbuwJCnz2i/wrKm4oSI4SmLNEOyVgmx9x9BVk9iPs5sCO3sHIs2wDUYuOyiUReCwaBfWyiBLlnc
cAwTtpwwvFhKIA+Zi4IE4UojnJpOl+Se8lm4w68j2L3FH1y3zAhG5c+u6KKBAd48bBPR8nrzpEl9
XYcCjrwrmbFq5nCG243+H+XzvDiacnCFdPMxvLAgffnhyu+8du8GLnwR5bIbKVlZAiHIjyTihznW
EBZ6h8ttRxJ/K1z6cSWHh4CLsPgsggH/uD4dENTlAKzVxAQfPchH1da3OFgUFPTKWoyRoV/TxnSi
pWe8w+A+O4uZiE/34SbrDL2G8RNKoC9VtZ5sPrsb9xB0aA3buFZbgelAhnXnhCAxPmQvpnMzsawl
Cis8tZqVWW93/oQAjtwcOuBSWLLR0tCZcZG/iFf/ITSxefvYEV8oGvAWO+NEUKKtSscaKoLf5q9Y
9UZ6lStVFNZ1ZFxuhiTRX54wpQDvyE5dAXa90pxqWqvcIFJm9YX7QC0DQi5vso8KjJ30iL+nafJS
aXcwLusD6Oi5YOmGluGTUk/sVa5vOJpFJZHKaqSneFKW6mOcNfxIPQOaOr2QvCFY8wnHWappUZVg
LFSdLBT2CJrI4eN2pAlf7hpYulphJaXFmrGqGyK809Sg4UhwSIn5pIm6kJzthCDdgsQsf+QnjlfK
0Axu5ddBVJuCBFnFVIDPGNU9vSmUdzjEa+U3hljKNqNVpCSNh35gvPDmHKkMqK/5XFXD4PyvAJRJ
qCj7ZOdPiLZzoxY9fyFiwXqdqGVO3Xhq0FIWCmI8tBld94TL2YyTzGgHJEKMsBTmBv5w7AJuCnBr
FTD62D+4lCHFFS3HdavwqPGRdnuwlB6F6p056gxRf1ZCUf2GBh7Gi04K4KWYd5Tyk1EsaNwmMh6k
3Ozecncw/0vB69a+iqT6QWZ8JPW9CMONiFtweTpi048jCTZAkwIkN8iJvonvYr9qYzYN7JXkgPDJ
nYLEYY/Wc0YTQF+562LolxDmtN+k8QwoLHHPH8JlpMQKwbjQNY4RFMbJt1OahGU9wHcDCuE/9mHN
q3IzRgptxAENGfzOCS/7CP2ze9e2pcqTFgX6isVZ/tX+OKtdGBkiZdCC2riS9j7WclXIqr/OMzvi
IEl9xVfj6xSt/YVU5AlkoACtzTJBPuRSTcsERPnXNC/iYjNaesyKqNGFSLsJY2STbzNq6DYHzkLz
tSzAUILyIDi890MBHTAfh+FKkwbx5k53icILel4QZypzO3VAFaY9Q5MYE72/yNhu0yHg1b9Q8GGd
OhfQgcZ+fh3gN0GicWs1/7bKZgeOK+YkoeYPplKNS/d4dK3I5Wu0N7j5Uluc5mKzHKONnptoqLO1
GepvtuVwqWYgdG5A0S6HZcPh7D8WqT6C+SBeYX1hnqm7wSqoPYBeZYQjjvH5erdJh1K0eGEHpNB4
KCgs4okSqIjA+PGhLK/c574TBLaHR1PHJhj15FQnx31dPJQ6jReCjNwMDMoDkesolFGRISTWSqG9
RcZkKO82khVe7zxvw5ALcFVqCdhOBoQXfxVvoz1vIVEg1HRJsaFL/ptGidMXg4GxMOZgz8XlHwhT
tttgKzDSyEQzMckP6FShRaV9mtIYTjYPIfIZ9pNLY+jRcV5wbBqszc81njVpvXb5P0g4GjSiYBab
PtgVLwDQ//iD1iExD5k+v07iWBdz/Fwl02tBxmCTTw8MSoOM6tWW0f8vfjP22FQMsB+duay2sdC/
DrKkTtJhaUrQJ3vQkQM1pjVw4niW7I4gUix2LwBOLPrvDxjcmxfN+yJPVO2t2GDEyN1QcqxdND8S
7aZIzn6a6rdUpjqSn0zpVnqM5J9jjdOwvgCbdF4Iv/MkJaThAKR1PaXWQWdZ08alAlVTQIJpHF40
Gd6P5xA3ctoQlyqASMVOhqIbcoD+dLdDGCP3hckU7PH0REG3NIwkepOB9l71ibcM8qrW+FgifFsw
VkQ9jERmpMVW4ey4IrRelTaBJfmYeN6vAEBJQqikVoV1aK/CgmuSCIoh8jAYiasAJ2CxG7oRe7Zu
Hyk5/UQgWjj8glktRk47uf2ZmM+/w1MClIB0q2sjBar5RlGTjGf9p5jJYNxeeJa4Mfdh/rUj/VEj
sPPnIVI/pY+7z9F6v3jFBPnbi3zxnnPl9GUWG6l0mDdlXfVT/i5ello8fMB9ms+ZiRan81XgPAzw
gX3RVxrTPNpVp565caMfFD2AnsE5uUaeEA0k++5cS14aLATZEoqL/jPg2tJa5ZYgkoku9+29JVWW
6efcGq/obV1sL6k5cTJV7z/CUipTNRxTeTvBBEokmV8gzRVGd+tNlQ9rQfupFXH7/T6HpROwOWhJ
yBXyN49e8MlDWBtxQRj1gXCmREIu4Qmk9kK/XpF9AttpmcKUi8/akfilBW9A1hTSSW+cfiFXtneI
z1o3zKYk0oBBFfipczmqK4Nvlsy3iOcqeM0p9xWAk2rjylkGUflNMunmWQFYXPHDl4d6FOiBg3/3
4ATBEW5ETX0oW+K0sSnscCSY3MxkrJWJuCMmzMbKjiXu6qT3WjiTV3f+HPfNqjHU0QNV/11lwoE7
AD3wWwYzpqMrRb+T57QWBgjoQZ0FX3wMIpmL04438wmBq3Ze3sTbk2LmOuLucI5wHshMXFjhKyd1
5v8wUjTcyuTCxA5GE4oOkQ8k8RcGORexbzFOiC9wvMfmFN3O/xWE06se/NgGXYvdvKyrNKmNhPAm
jOnYjerAH6iuaA9hfngQBnXD8YWyXvUtpuG83Ao21+zHfRCEdIcX9o736+96yxztXbQFwWHWTYSn
OEHehIH9QEwx18bBOQF4rbJtCoGFNMMlutZPPrspc+IaKSgabN6ywXfpiuaZaiNUME/fobEipqZh
Ryy28FzVO8wSVBqIiXDBGrfnms3PZB0eKng44fBiYd0t1Bpex//MOWELffA0tW3W1zLo7K99zbj4
zJDtwRZJiVq6tW4O8gZIk4Wwsxr3asGqTUL2PIfZtd+yZBtJUo+wNbrnfxL9sOKhKhTecGA7gNGy
gjhueuI5EMLjM7e7rpZ175GQjZWauQqV+m8sW4r/v8auBIgcUK85EJJvkebrM1yvoiwx3wu4v8QW
e3EuqtzyUeeL8ZQTRu97CXv7qzLumnA9clL5a8OBukgeasXjQYVbFHk9E447fzNvN1MI32aH0JIz
4U+T+mhG8eeFQWwvMqF6rO7KKW4C2/Q8M5G41ILnHV6ZOuXeCDb8fSH0r4jFyEmua0pie7fRUe+r
yDSzw8KuKP2NwAnxw/dcP99lmDCIQCr++JjiHJRZeja2tqp8Nv3tJEUeebEXWamYFK+u5RQhf676
TvsvC+eNF1S/d4u2wk8eXb1driLxIhcRAMyRekmECAA6J7Co6xXi9IrJZ/smQJiZp+BD9Kh2KSmb
azPYqCXifBylO+EGzYm0p76Yq3eomEnuZ3J7fStKBE+fSmNUwqaXoypCqDnM3kPXACXdXFK6gVsL
NfS0K6Wft3NZABFw4plK8Gdncz5xZA+1q4L0vm3Cn7ECvuNTMKxFHltrwgXUmEdnOxyYGXLleMQe
xuLEOkivPd7kURbKZ60P+o9YzczZhcYUKl46GqM7Ed9lm+tFEt8+5Bmgyr6eVTXnmUaTjWOQktgn
f14d5kep1qNBOHpw21Yn5F7f2Qf1tA5ddLLbPnOdIXbr6EtS69Iduqc9yY2jo2TgHJ4KHADQ1hYV
DMwyYdsRLD4m6VY/GGuaAAjiQdfhbjxvKvr5ddGaW44LOvC4AVDjtreNfu3Tn2VSNZjDPt+isQNf
H9s6nqFRjnfXajTRy5xHoV/LIiM4UVw+CRXBJIn+rLFsdDXtpjP5C3meT/B4nlk2IR7KL+7XrLdn
Wr+HNeFSzk23f1sV3TamVTNgqkIpF7J0PBn8QH3QfiF+YxjlDPhvcd2DcE7ShSPuVxcy4QGG3fot
nhN8DjqhkjSMhyrZkJb461XlwgEV94qpHC/ylJrLsJyaFWAWrDRJXBLjrqwGILCopL0qmuUupWQN
mydRMlvKq+vCBNahj14CvVrEOJHOz3l3d+/YLY4Bfl9krI51sMgrn01AIxBDHH0GGtEZVMFNNLW/
1uSFGioQtssLh2/oIcbaaj7KHn5YKdR7J9W6gVV8YFh2CNRdMQft0hyl1P/Zeu9JFPaBorq0x/bY
eajjE15OTrd8Px8+U7f/s3CZxlneLllnhb+mDiqtqfQJFKGZaqEWn6OFHCAjrcmVHTfSC6fRQ70d
KBEvn1AVwNrmuQhqh2S04gJ6N/MVCEQNpa6e17kjirKZ3q1IL4gmKH8lSLBXzyW7SZBWk3D44AG+
sjdOw98SPKocDhlWMFG0leNqwY2m7RS+YTZE/p2ebSwHczr+q4iQ60ikLdTbbLvUnPMsXgbKupJr
95Li3zz9Emd9e3ozGWpm1jecCvDGYx/CJk3T7bSQ2pry59qdiAapetBC4lB1OuAZIuBsoTeZsCgi
rCrk2yDd0LKjJZtyXGhuKSva27Nwxh2QmhDU/vqhMw/unzyKaJixafJm/3KHMc88hM0QnhgwNplY
S8zt9wIPNrVmE3CRZwIN06oWYd8pQ6OELg+N3SCWVHl8nYgPgFWIBqi9xEa1zndJlfGUwzFu+uaq
H/wFHHk90dqxifTjE/5nDfMhf3/SyL/9BQX+c6tMhcs9b+q9sDhsDr2Hz3F75UFZx4l1Peic9VzL
knheT0VaPVjKfcHWi5K2PwjOZ4IyKx1k9O8GgtR7hJi+VG/hezYBqDccy1DtE6gOopAXE89tMVcO
08HjjfFqPH28wzvcTyvjVseWyzsEXI2fcUsZQK1Kb1NISsZNEVSrp98lzdakNGw/SOS0JtoMEOL8
tj7+0xeSqRE5nG/yZ4W+EYTH7kORaN3jKxubbuxiPqv3VVvBrg4VfOBJnyWfJN9b3CfiNmnYTXqz
n+3b8uNKYzaTUpUQ/eZMcvY1wS8qtGutJHo1MR042p1jqFz/lijmQe+Y3aSuuIstp6FGGsdATuRN
3Phf03O6lIb9fOWQ3/0w+DkUs79UJo5y5MkUGxaBTV2eVYEwbcPEXWsw4sFdIJH3Vva1cz7hIBGS
I9lOaCK9d5pu4NjHVd98ArlLQhJ9VVRjkQQzPkl0+zshK3ztTzSc7udrn54Lu/5Hq43Qu0EdGqhc
QoOF27/pnHA3S5XYAb8867d3AMhoQ4C94aGRGe4razVtvPKfhloPi9B/mWIy8EMkEEnxN06mfVK6
ZSAJbrZhdRaNTCGPG1k3lL/+7Alg7Ghp15v69Rn+tF48Ex5yG6oPnbuIXtnwWd61QUlxveHE1bT0
tBemHXW5Z1l5z4jUp9b8FKC4QrdJGzFG1CbrH+OLfzGjHDkz6XXLLmAKkg51rpmHsRAuB4W+gngu
sU9QMCTJIfhZaVFrjDXmcJ4pjtuFR2oiyXg+jMJ5Dp/+IOibc5bW3CI0+PCwGpjrn/0zTa6l4Sic
QX98AljOJpYuc4LSSXAh6+egJ4Q4MHUI2k9KKbUSxtJ0Jk18PYTxXUJrkgQNHP5w5u4XpUypqwAk
sd7HDRXlcKlMW1awwlOduhWbAAp8+xIxuNi8a3C/LBff+FIzwp39JNAnoJMzePrntzdL42E/2ue2
oZkTkE7+lh5oJoq191IdWSxvgYtqtAxrc382UoF908hkbFSXQImCGGVBSDv+t3y1VUg01xg8Miur
Nz0DOUDcrrkosXYacT7SgI7AR8rvntwX9jhL68/qCKp1x4qRgXTt4NTITlSRptyIhCtrFGlplqWz
2c/kRvZ7p+KklnYv+J3v3ZxGjYBWQahi7f+9ciIdEaSMpOVrTbCzTGSD3RYdPI4B9QTGOBuRKrm5
MC6NEGp68X0H1w5j3GHHFKEp+x3bWRAkN0JvUnqis1D8FJJRIPE6/F6ECUdNVQHCjst5sx1/1xRV
lOOj7thDo7BTJagR4WIiYVOcIHWKR6H8/S7XO1u9ed4AfaZ++POag7Ehq4Mlpo3QR4OHagKvkkd2
K3gzbIsZkRu46WUhgUzbuVQCpfTNWvCWtJ559gbwG/bKhuajOgdovdDGkEmHgf2aht901KoS6Uhh
nMHeXnaRO0YdK7p9VVJh5D81fLkM4YlrMlb/qll4pN5C+SmHIq8LoDp83YAnEZFXqT/k+i9Sqhps
85ooGT6Wb9TvPA62FGri3OiGssa3PNZys5fiC9IUbWUBl2zMFfDy5DusUkiW2B7j/efnMGLU5PJ2
Hd9EvoRWmbtWohrtU/4z23JP0vQ7gqvVx3c4AGQLQqZailRri1fBhT2/BBm9RlqBufRTiy5BbZ6+
dc4840COarXTGjk8n9hqYSSJ+WA4tsxJflM24M+daOI7zPpFXBa/KwE1jXxFweoMY6PPM5ZpfKnm
71BdsgBk+CVkvcDGZv0KRquJaQ+RhOptKla7hraDmV9pIMgh88l9oLVyTu35ux0yapZrp76R4pSA
b4hgZ6+azcIelWSKyxFUqVHjYpQFK71R0R1jtLvKLd051ZPYcNi2EFcdn5dCimPKAtkusZRaoUxq
4vW2NMsF1Tmw0yBl5ebdl4uE/lSgwKr32jQu9IsfxD6FP1yhddnbarTYkb+Nxa3RCfwRDqv6rn9k
8skzLc/76KmPpKpX6SejVmr9XTGLcEQVuvbYH9ugnZk+aBM8LuCiHpiEZFIAs/JgjW45yahw16q6
9i9Uep4HHoFwEZmA3DaatwKl/w0sCcHamXkFD9liFFFz3iAKsOQ+hXljHQSEZtMREk0thvs32yUy
D3MxD8RZ/yLccTEAAJ+R9+N8LWIvjY5qSCJlzlSGKv3y4X6gExxUjHjM3cLcdevKqmgZWcoEx+Er
ZflxkSiLf73+43V7aYLfbXDfFp4F5trTurZvEG/EXHARiuVonZd774W3nS1HSAUSn8cSBGkeg4zv
pNxY60pfAc2XWN3qp8Qk1rkIkgzrMOpVa1y2mUNV3ODB9aTCiMzoYJi+v9VWS2lRV82Q3h0UFih5
TgD8F5ZuUD+zJ2UFaujcAeb6vuhk5SUecpxef5jE93ils1MqZHTJ1Up1GBIXNtknY5rU7DGQ4Z1E
ZwtwIw83VAofv+AG1ZPzyUHdyd10CQLQ6HdNIfnr6pS4FlzmDQ/R/R5hHHeP354WNlVBH9G23fNG
2Gf2skNSC4gbyvXPF8S6Ky0X91r9tNhT5nI13NnwoQzSy5LFd6nLRvRwHBxpfxC3bpzKIhzWhWk9
tAKiCMDlzVi3T3sNnW2MKETKLPXRzoMo0sUN1hJ0CEzP2hWUi1JxsM9iCLxODvAfHwhYXEyo/GnE
8jV6gy1h79Lr5atx/T4R9YyqRdh6LCw1HsfnXN/nrssWtnYaF+Z+C0BlfCXZ6xsWFwOKX6EQ0Vz+
lLo928lbyMhL4TWibmsweyC/4TSU3iEWxMCoEw3ArVghMAZfnS89R1mTbSD630Gn1GxnGy3njjVa
aJhPJSGfryq47x34hoNE/LtzS6rhSp1L4X0TMBkQd8oJjUD8tiKOxWnA3nN1irVqpD40MzJrETGl
PaT+xM/ZGbMJI9T/h/NJvG168y/xn0Vz8FaVi7t9qGEuPpsNfbmA4TLZDRtpGFpGIhr/D2vmYBK3
pPLabotccFcLjheIciyhWteCEGgyQFsUMKAmDllfgtWUfiLrbhX6b2xg5cRB3DHGMCFPKC71pwyP
4wj/w9wZO57VdeNLzsWvnkuAZMo817jqsvuyfqlGdI8wms4RiH61PHsRCb19essSByXF6WqiGg9W
r72+sNCnubtb9ojgDxhW5qFObh0NSGsZcy9ey+T4BN50hiyVSiR0Z0owoYVx/xYbE5pggSR4Y1So
6e820ozLSyGY3VPDZ6PEt8waV1T2jhDUgBSjKj+HNrghwSfaV78N6csVgSYtnX7rEnESEzMDTjr3
fXAAtpAOvzvMxVNSxJ8CLwoGGpb2O3fFEvaAqzzJ2ZXTrj8BQZ7QUX7sbsL67J6971ahKX+6nEj2
vzGPtb78OYmbDrjHn2rxIsw8s1SzOuv5R+DW9YhW2/2nkx2zwuKTiR2xRvlyCl6SCTY9gnngJmKK
4ZWyPb81vbg4yVBAkH8OA+vqsbXt10Znf4o9mljK+hYyzUn08odnvK9bANGRGY34ebVcQ6CO+SrF
L9PAO3RErj9SapegK3Fd/s8yeziGgldtFhkoovNj2J3vWAwhagfRyL+YOnv4wofWs6l4GjXSqkbR
+ouEWKttoYWUvb1WiI4qqD0CgxdPo2h4cvwGCmkOeU9yPKBxlGXT+o8qPnI7vPPmJdAgf7D7AEbm
xhFlrFI5Zb7DLsVc8mlWwa3xyl/0OG3AL0YXO1tNSYnsQFM8hCHGicOv6MTAgFevO3CHGDxWIV4b
KE3FchgnacZ/Z7qf9wIPml5j5f9QGPOewA3JGx2CwiGPsP2vAEd2S5slloiJkZDTfmqxlDAcfvF9
4pxKMkOkqWorDDLfg0Xs+dM7KI37qYYSuKsQn2bXF5HutKJK+POG2q4hfjfKV/kS7HA3yf99l3nk
015yKQtpP7FePQ3StEeNfyIrXYAXit2Gs5kmvB3Zsh7SuhSw9SBgr1wUDrVhwPLU3kNq+vJJdpSy
lIwdwvEDYB+iu6nR18V/iVqhLkH5vYl4OmHcM2Otc/aEz+jmJvysBTIgFkXjXOiVs6XoJxwGYGtz
qNwJQstqyz3AaZTFkk2FU/wwi1iN21dFtT4nbcwbJ8En8XKRPOVCZq7ikwKgwFnSYsJUqhTRK42V
3nEgHsplgP8ptk09YZ2TrDTy/p+SeMsNlUZXrx96fJ+HQOUIdUZ/DOhqhEvCryda54MOf5mnq6ZT
bAr+qMX+IUDLAycEBEyYboNdBXxf70p/eaeaL8+mDGs8Ikz+4OH49pTQI7XNueIvMREp8Km1fdDo
XApVUUjt8fKwNXo/D7isZ3xXJalPk5drahtu1D8e9GZxMZlMjCwa8f/YZPxXbTrGh2uJOcpgX3Di
nzUyKBxuLW1xH+uEN/faLDCCuAw8dzu0JGyRIPcZOVZV1MrtB2EboCyL0FMqDAG3Z5MS1zEX2OV1
Ya1gSYVt3pKVY9ZQzt3qzF7u2KLmOQfCrF00qIR66LmnJy6V0QAc7eZkgsBinelH4JT9aLcSZw6x
09lRVRnFDTfesS9DDOyklAll5H086eLs2Yd6c/YcPm3gSkkg1SNHs7peQHUHGQDDnfoqxi0VU7aZ
e144ruQrqPzTK9t3kXcxpTC0OGVu9T11xvJZD6bwzsbE+PjwZEiPLqTynLsq5bm0qbXUqgB3z2IG
MSC1DiFSVoRz0sDwPobuonTcjnivkYgNzHkgEa1irM1PwWfQdW1wvtFlxYCljHAFoKYkaRZtjUOm
E+3TLgNcsVNOJxer6lCrOq1skuUG+2Qbmsajjt+7H2TPJHOR9k+nCYsF1bn5l+vxhjwexOGAXGHM
sC9t+fut7l6jgWUYoYCvFdPGsnGMgakDgxGhQ4PdhevmPJho50DQwTO8j0vBZIw7xk5qjl7VmblB
402YBsw62MXSv916r9c8jwRdwmzjniemMbAZXMWb58kEiBLWkm/JZa9iXkzDnAbtdUlEZ8hXY0BN
XxIYLL21DXVaODx0CjifHe9Eg9eXwuPqZoA8MME1BIAWl4T/WBrvKiPYjNPNVLQklMoUDFYQAURa
WOr66nHQ/zLprafDrmqcpH2/ZMCx6Ie7BLUQXBMG54vuqAvJ5syJYZAeIH5nYY8hwUsfY6Q9kqGU
llKk5gtCm8BTg4T+5gI9ItNXhMdbE/Oit0IZ3qP86PUm1m9qCcMemJ94eRmLXNzHFTwP1nUg9F2S
wEgw2nbltweQYdwWqyk/RvLOHAa2L8shFSAEYLZUEbbaUGpY97h0dHcw9D2/VUfEEj33SkZ5P7X5
duQFjecjhBNJWYe8SdhTdK+AUTypdFaNyHQNS034yH+rflh/uVtZ2tiW/gwtc5+q5W2KKMQ4Rf6W
ITSv6s6mWtXO48FjXS2ADcKPXAO6s/lLkzMZu/JNQ2bYYmAT4vANL9wZ4vNUjvSILO4KGOMXdThK
vezgeDMCxt8ROwG1raFuLOaFB3H1DXldOp6oBVw4F0NMPGtzhLQRiemgKbMmOf5489NQtww+/PTI
MjPHDqgcb63OdavdimRFLEObjj4i4qNXQIODC2ABxgkXOYJgvfHEFrZkOuyG1h8Zvu9s6hxgsuV6
mL8+PgO+TwZrGCUzwVfDp50a+nxrNGnTCjeKU4OUuY/zSBY8SldbKvxNMu7nqGQ4EMe7vAIvyvMp
8G3YZ5n4AlMJ8zFuZYd8UqpGxckyzHr1Sy6Nu+bzsToII6eIqxflAQzKmXJ6AStEG9n5NhgmoKoI
bJkBWzuMbytJONSshM9LU2EQlcQJs8CBU0kP64wo5PaNGwgWbQ7qsjU6ACQ+dnfsT7rvnr30Kq4R
SjKEu68V7XjqR20Vekoy0o3go2z0VZjZTc+qkMeKQwNdHiXR9qM9tDP1YD592G1hlrIxOqZH//ON
pFitJo4NaC+uU2lV5XWrsTxqrKUIcKtuVY4JYz1wsMwY1dtMWYfPaegzF6OaV8fYV40Zf5YWsisi
M1dtBSxLoO/OlPzCqhkWbFmEqg1BvrFKYZ/sy7n/qJA/GRVnb3fySn43SXPD9OOMccIC/k/RUGY2
jg68YvRuZqWpfRE9UwTYGRjUbRPXihGQTn9+2n+I3fmxpDy9fluqbsPDAVW2/BPS6Z32tu/QuYrJ
2V7smeNZ2xYzN5TRxa6KUFFhohu07pVeOF1H/fbT4gsCTPO3KbR58wrDIkHJtMCg0I5AJiRJmLaX
pDi0EKcrivdtnp9kAYw0SgHdUex9HdFZF8hr4lDRct5eqS0YS7ZD8kzagNz/kGVV+GLFa1OOE1zv
HY7cZqK00icX0Uf+PcDdTBcAfrqa02cl2D7OpPOwfvaNeJWrQQfsR44UH/JH2pF6ZcMm7YdjnLAR
dMejzX45+XdppgYwQGbYvvii9Bh80ONnbcHLc8kEUR+55gaTgGLdnM8ztZbwbb2+oqAAOCVtll80
m9PUV4/SKEF6tnQYI01Rqc6uyJo4UD0B07W/weNYqRwzvusgCOrNmUla/tmAsPobf19KXtnXTQ9W
WhedtB4jySrXzdLBgsdGjtj6wAz1NDamZK7mgZZNHhoxKYsiOHU7w7ojcQ1iqJ9WXLYvAm9vHIFj
fCYMebxrRZI2Je7XNyrPqR+Tdvye/qwfkblhWvm3Cz0oM1iyH0MH6gC4sDS7uUwMd/MQ7IOc1Rz7
u9E7GmS384fk1mo6tB1f2l0JCjEu58GPKrF4E7bNIXLKfRQz1RJZIAOEwkHPC5rtXBnN89E5Ti7x
M7EDX7ECjp02+hNDUpPmlLbgWYohJrPKuz625v4iDybMrh+rQLLSuIcqF+5gKLCLEv5qtk41BZ4E
4xO7QdFicuzcETC5nHgif14Mpm7YtyB64UAMPnFEOX59jic2J8Me3Djc5zgGL4LxrMQYZ2uE4cch
/Eyvr2vX25m/d9mel7v0h85iUFym4JVQXkPpjISCaaJZXYTnrpMeKhZW7Gb0oTsetkwFExzLvCaD
xLoAF06A+wwoGBo9Gi9pD6c8FQB5aCZndJbxB8Itu6j0kbtLdCJcWSyxVru27L3Dc8thowClebNR
JygCoQUVlDZZjl0BNEL0JHE7z+nzXpvqbZo4sQb2DW4ygdbhIGoXpnOPUctisKeCPjB0qMe45ugg
8aHxZNFrGK2/ukRIsdTgCKd7gdW30aHZStPQHxoo043dvXwFfeLeCeQYMppZiFYYAvj6rR52M8Ky
cr3fsl7LEFiJ4MMv2rWRbfZPvMdWiwR4K3BtFZNBVJer6KUihhTDMx/mUdvk8agO7GePcETy1IiG
MZQo5TH1KL/nh00Czfcc8knNZZNl15Imq/J+jEFE5/D0KMiAHq0z1VNJp1ywJsNBYcnhF5+avswX
JBL+hwFqjbZ8+ljeShmblLLTdDzMkrCJ32vai0cZLz/M2MMKB9EdPSXFuZDfRKkkWp4Iy7/JBcTc
TP3VgZ8RkWPJvUv8HD6c4EqCdWg8GCiqjcORFf7Bms9W6BkwnnuItHkm8j8OGaA3LvVMc6Mvw7F/
RxHojJNpW0AlgI8rs12Ogly47bdMbOijpy4mZDcjGWne/nEn4P/FelE6utH8mt5MNGY6Cco7AK/y
/D/69/NMFhtqHORLPVzioclkJ5nvb+QLGKuzBzy2Jk72PZbH0zAG+LHkQTTu/ldLP0ycwQIaHvCS
6RuUbKNSNB9kj2p5G0Cc+okGCX7njMrdKxyKnwf0h+of8nWiK3MFKLMRXoLAlJeu5TvqeyzB5nvV
dfqmrIvPQApgzNj3eBCaYmm0EsDi2upvZ/uDcM+dlmUp5lcEiLJJGfcTeMut0XwiEa4reV/bYAoZ
t24e7ktmi6rPN3xnA1nkjSaIthdCi4J1xMwRxXlv8cqvLhVlXp1m4A0sBFLYwUwVGqdCvvS6mavG
azTJaUQv3LUbcjvJADHjUSrh7MIGIxDtZK55cO7bBzBLl64Dt9Gh4yXUlOUzyygZReOqvOqcfIW/
wft2GosAFDTGWW6zPXe5vKJgeuD3qZCRFszno9mN0GpIMkE0G5CpUIIwjztB/e+i49aO2U/aZM7Q
mKEiGwawJ7vP3J0OmUvWFv6YO+DtIQChoBvfsvkPisd/xAEUbDcMrDYH/I1MpjguaJ7T6k9k9rTe
z9T4O6VPIz6lTxyHovDmWGwcI8giW69javbW3WvmnZeKoWpejPpaM/8qzv2f1RzbUwcElyD22ubA
083z8wvd8ehhfWT7EBsPx49LS9fMW32z2fLttMPVk7d+h4gCDQhJAtpbHXUk7ZnpLTyRHziWZoXG
MietTUgSAWJ5NCaas3ZGRbW8+5oZFPiTeR9KV7aoleWjEXGFDCB8CIBZ7Cj6eg6SVGnRwmWDEWuw
GF65bboZcFNDap1Q+VAMgRoQLclKHGUcIOPF43btaSM9+5NgOMeuvenBgW3TviT0AMIwCWsgUkKA
X/Bt1v4SehB0uiHmXWGHn697/FT2v3S3fO+KZjal04EkJ5aLzLBrD/GsObunxeyjrOfXOrJxSHRT
+kEmcfYFw9kN6uy25xUKXNNbDOBvVeaZ93R6PSHok4Sk8PcFVtpbi+GhJrfVeUvdbrx/BCfy/rpX
KWgIqi7w2gqq3T/bMSnUXGU2HphRRYAucCUOpAZuisTDsuT0Nd34en1RvqWS03Or0Ajr1ssIWeTP
cW/kTaDqWash+fdrbjDqI/l9yeEdAS1OeJlFAygXIFvsMUYLAfX9l4vLIlVJFrmcvN5fdLT+Nw1z
VOmQEQfpoR209aBMRtDgy42pJ9IVNE78ClUXllY5R1zd99dwZtHhIwTRa0HF85yZB6Npy/6CeaQx
wb9zBkzo/eeUr1ZDgIqnkg9uOVaMnyvYigzBuq/zPzdAXFi1U6A/vmKYr9rD2VTO1l/wJxTaiOSd
T+smGpyxl/6goMuFw4C7f4UNkTAGMPZbEXUkCwRDrT/MCicZfuzBdIhNN2vQS/LrKVTKIz6wpIIa
TZpFFih26r5RWNua7y8mtkZ0aGmA9dt/pHpQU6cx5mTOFZJHKHhY+f8zsizKgznAElAWz6CERmPu
tMrGP8NFmhRAlvEOAWO6qRQOt9MJ0Cwgx1I3DVNY8Kl6tQiKe+0UW/GeMndPl6Vn+vGeh+EvIN6v
HFe50aGe86XFympkjZl6pg+JStGB6HhnDCLOPyqEwIg27V+pnj/mFWIk4bQgAnjsRscQlBZgMfGg
mDACo8547x8UwSr6gVHEXKDm+0e4jXmzFFvwpgCplfs7mEMCxmAMF4Hve9CjGHeHTNYJbxaEX7Yk
DtYQyq2UC37qnidpgeUW2P0WufzTq4ZbIDao/Wu8LRM7MA7zsMSpHJlHan/s6MReQa0hWWplVqyO
dk1OKVqCbQT7GM1vMYcQd6UdeYmv0Ran1213qnxalvO3R4n9L02MzWkGwdz39vguUVJ9x2lm2JKd
+8cdrxNj4ma4L03b8+SqcSHXneiNO9bhvkKblhtQYAedsO3JF8jZBGIudFIa6c7vQeW6srN4oKGW
4Uy1CtvhV9WoF1/liW0QDjiu+JS43tML5wCBcHaKmytgmf5dvrHZPC8akhb9gXyodwJCcKVnyw4j
ptd5YHElJBVQF5EuGR8Mp4huTvXQA8egFDt81Aab25DyZ3ClSJ7w5C1bDYZmH2l86jEENxXTcBKs
p/jY8hBJnF92RJ4xVEitmiKBNH1u2J7JuAQhnZ1Kl1XD8lRNeZQUpnRGcgIOcwKP1eghLEOcjsuz
M9ztwggFHJ7RTZSwTzmcfdFzDEKYu2JOW2ApKrwmTq9w8PggU7nQG/NPGuQ+kAYZu68xCC4IkGp9
8LtccXvqqEx3a4fXonJ1vnXWE6HvgOwi7rxrN0AaU1QdzN7i2Rm4ZCgvGVg1g/DtJTEhaxEilQfI
IBFO33DyGYVGO3tF7snX1MMecRV7gwEcI6K4KNgNHUqeIQJ5NRlT5t6QZnEmE4A/Of09wtUkE0iL
EtEesY12J+l9blVsW3NN64h7BVjl+66DnHXCIjuXD8TTK1AD6DHfJExXZtANjNgzKfU3qoWZjTgb
7ecCo21T4DW9ZS3VPVsfTvLkPSWfq5mh9m6DVMgph3SEbAE1e+kgKiBdQmxNS1HJsXgQIjDb9cRq
Xc6k1kxagA7nATG+AZs9BkJKN4rMUq7jZf5G+MO1cM8QdLOW+oVfVMaUlYJF2yWS9agvNjdoSOfh
l4h31IaN/z7hh/2AlM53uunm15Jfxa9Xhu/G8wx7+aos3IDsDW6j+3uUVjAkxcQJpcs8IT3p397F
YWsy4eC7up02pVLpXQCVVhSdF3rjldzUvFR79Mksi7RnIYOSbwpxDm/x+SRmm9RBkecd7T++sWvo
quFE+QrJMdqTOG+Lm9BMr08SFhP7ZGrwZtpsQnl7z58fPbNKe4CsaDEAcEHfCaXI4r1aVleCLiA5
bgIFFLMEEu9GrM6zx+FbmZDdYZQqOMDMFJIMXCY/f1Ji7G15BG3j0UoXdq6SF50CB6EYYtOLbctm
yt2/wN5a2L7n81d8nrdz4Izlu0OctqDwoi3NBsyD3A/TIlVePwM93E1gLe2l78X3rasvjbD0QEKf
/leLZ3y9gG5DZBVWqIkNVZn4MTnAoz9GuJaT9OWrl/cV3jXoMwJGF4VS57eReW0TymA/N6O5OsGh
Yojghsq+1wgIx3y4+6yRXtyutrl/NJBTVSkBsFxJHb2/8i6rtVedauoswfabWqrEV5hN+ydzXIwl
BLlE/iKjcg5OaQpmxoJwtEjTGGcwuthoIko5UlKDj/CHLL+dBpmt+KTONA6IEIswFwYz8kZRF/LX
3meLXqTHsZ3SRtodvrsQemH5mD/ncWtztPefqmOWjViKpCrM6nI1Sc8T7VdXTNr3DKCeeRTJ25gy
Wf5GFT6beOCmiDg9lvxtZZkvidFdx+DSRvhcD/qiB3L1BGpNVspb3OEqaCRr/hF+n6CdfFM65Nv4
lyvou4lwxfUuPp1jO596gABa5NjSi8GElWgoYa8QFSJrvyfkqdyjEUuF4WN5JwIHN46cltjRhM0g
j8ZhbM+13wR8XwGqls9Hf5T6AqJXXJa6Yy0KOOg8VoL5Kky8J3r3REDdZLbUzn/jf4boMd1TGOUz
AidCSproEpSUibD7IzraoPPYSG1x1XzvBJsWds88BF9NV/zt0qaomOCzosf8K+HABn+Xeg1FITiu
T7u+8KfTCJJqpQ6pvY7ZWBVS/SRTg6Xm4ssfYy1GCNO3px521kp2bz0hERLyFXTSOEEeC1htZ6aa
yYRxmOgvQIxtYMjkNHK9toDw9b5+4MkgXU31pg2sFy33DuqT/Uto9oSBDHILnjacUFuZfwU+RMXu
aXkWXN/dZomzo8ZgCTznu+I9ORWLo/4EGAmIA0bUW/U/jFXR/JTPlYn9bRE5++SLRkpqatxbKExk
LTUFtAZB1QJsOvpsVdu0GMLSIKZ+XF+ftK/eJkZf+a00EJcxSIlYTPatc3MnTq6Kh97FTW0LSaUr
Xz26EX20kehFvdYU8jcdeoneq7YMrn+wIeMcOwJFlWry+QcYqR+knZvTSPazERmsdPkbIk8x65DK
RbAN0+U8H1Oh1CTGGxl6HOLwp+jm0SmgesRqQb2WgLomqsM7aWdpdZwaG7a87LPeR1SZdY9Ayhrf
BZr9eMvOp3QP6+g8BlV7MKfgWepUduKbkCKXePTo1xy6ezaB+RVX+PNhEExIWLPxn/WF+Dpnjepp
tqP9u+HzK+bZQ4h4y4gb6WfOagEXRDkywtmutQLyiMnXIzuB7iQd82tVbNei+M3I9qnranUdwYXh
YsNhPK5Ec9ulzglB+jd+2K/hAn6fAc8yKTxwI0UbtR4jD5Op/Mk1gnwmYuoHitDbed+O+ptYyExL
G8Ort0CDyi8VtUdweT6zsoi65KF/SOe2qj+T5/kiKkpR0QEl1DRdWM/vV5bf1EfflM+FLAiAMi4h
N+pGFAL6OI0qetjZfl7JwUcVkvAWuoGRPNdPS2xELd9O8IT1R0sgXrHDdyKe6qLAMoelAMCr0N8l
/tWi9wb/xDQ/AH145h/0gDSGKRvTpTi8ySVDuM6boznvc1lcmx7s4BtsEDOD9s50mrmNztAfE7ap
lGMxZ+oX6geoZMfXuSqXr6DxW0gGE3x9iirBMuscMMTi2/hczeVw7EXxjcZfvcUWqmsep7yyw7gu
U8/1jAJ0jynoWNszlEPMOwJR+jMetHas7tkfPHZgQju1vm8fBPhIwCQFL0HaFoIagisBb8YH1k6p
etb6snqBZEdqx8jIaL/2HN8OVG2HPBPGqAkBzzz8xUA9k+7z8YgS2yA6QkoUocclDRFK5rGwkytq
CCgePf6vTI5mruzjBXqVwEmVMxaFBwbKJ2YWqEj1MtLNd13SMR+lun+8onBm8o01wPUtUutEWxxk
zCGtTKAFZpnb/+rCR9diM//d4nfBvOAK5x0fKgU5OQceeIDXXVkUDovveiwgtTaLewE2KYDYLJQ1
lcNmUkBTo+H37scDgueIVfKpFbNM1Ft9gFyCtFdl9uqsugb9qsVdfTPqUfdKThOxOoYmIFYRePm/
O8y9/fnzpuuflVvdGYtq61cqhJBdPez3hFG7mE5SiA1mYI7LCiH6ka7Br5thd3noTFMrUnr7NGpC
251k+HEkrsNF5wh2LeiDEIQXid5jb91nQIXW0OEGZkNHSGD4p52Oj/8cg2+y7UMjVnCUXwXj0X7l
3Mac6Jbz8xJjKjM1LVE8hfzw2nV4NX5ymrvyhxnc+2hFFAchMm3+2TTqoJe5RL2BR3d0jJadGf5m
i1hDKQfnS/DnvlMhDgrfZKD7GA4Ci5axJZ0O1WJCIZJmRvNf2CuvWbMlVvQeoMkRjuyPhvXK4zE7
7oEUkWqdX2VtHgyjpxSrZ7ECwXmXsdPvXq1oG0YTmGXNs91GuN9xSX3fgAAFQJ8sLCUlmnOUXSCm
2ed7AROnU2mMxF0y2VCAGU8BVwRXE+Gd5fWXCD2+z2qkU4Df/uwuXHDA1S3T7a8XU9L4Q4B566Vd
+1IrvGT4GlEOD9NquOHByAsxqyFKjRkfAvZ5sat/zlbfyqK3v7bSC/JrPu7bBsLvEg+BHjstWRb9
EKLqy/vp4AzXdSZtCSdAVbuTynFuMlZkcTXgkH9ARZz1FsI5rLpROhs3pAxeq0UkbD4bvfYKawwh
WJoSO205MXKfeSQHsrzB3ekarzbyuTPLFL2lrdsTbaH+1Niam6toh3ZjskYikzK4ElOL5JEZT8mx
64SqtggDBpHlm7RDeAke5yYJFdaURzfGNwHEWzINa9KhLv8zb07BPRyU2AxxPBgz3PfRigPjaLsB
Chuk3zqta1p/78eBWxFz7HYYYvr7LUpe/D6Lo/BrPw/VA+jFPWlRJolexlugsBoxbvkbq1Uzxf4z
H+5s6fFDyXYVg8Xa6yCaI7AJgg16cVq/E0DsI05mG4lbsoEThlaumkM80QnnhxrA4vDzlFmZ71D2
3qZElryCAEXMJjqw0P5D98Ezw4dN6aP6U2O5bR8zF//PHWI2Cx710c8J8G6Yth16h206C4zSRQwo
Hyg8mTC4P6VWAKiRHtPBKHoP7htuVSnNVHCNEOgu5+nxLhkkO55zwl11bAuirp3HLHQxp6NgG7Wy
IcHywUPQt92LdoePdEho2ij3v73a/uXgCnmAkq/KVHn3n3Lrr/5mL+I1DKdd2393iOUwpmBiFSxT
F+PGXqWS6FnwVuBzBfVoJiSW76WJj9Ro1t/1DBzdFE74z7rPRr0XQWZsDGPr7BAmAAopn+PlztJt
Ltf+Krtx+9xDhYY7p7/VY1I8cRU2Hm5N3N3yVfGpMhi5Lxk4X+NdAozHmSgTRKROhZgzmWAZqyze
sJf1TILoKmVu5ViIDcaVaAsJEsXvSkBMIq2IsRUEstRTEfUpAZ6qHl5pr9F7fWg2/Ao6x3puNR3x
ER45F50ayUT0PrDfqXU/Xufe9Tpl3A/03WXe4N6ZZmb+rCABMzXPPFr0OdrC/yt5SByRFV/Ds//R
V0TbAyabSmFaW7aKZrdrteSzaDybCHdFzI5U6cz5cMCJ4vfXrWdn+P901tE1IPECgASa5PXk8aRm
+Zu8u9Ez/0uvnYAjoEfexBft+q+T3ynpNMpD3hfwj0AdVPJyZGQtDbLUdc6JDeKGbLI1iFMM9noc
iQhDqjprGZuxx4LD0mhKu63ivHwy/SbwFLj9R6nE6rgLn6vptbS+b0+PriGTSztN+5hUPMW11IGe
2ZLtg/Bi0IwJ5uwR0NqLEp4T6pr6Q6jErOEgKFfw99C5yD0hKDIGNPHxqxc7N56Sf6+SRHAN+Aza
M/q1/DzyPVnnGD+NQ3yAdHOOwHXxalkFsbRDRp7HQjGX3Cae7jsDQw3M29GNVn829GDYG7tPpI7R
7aN2foaAUFdRa9Hr9gOA0v0OT7QopwbD9SCf0b7F6FQ+W5TmKGUqCsv0TTRU+nVcY9KzpSxs5CZT
P8EAWBSTpBi76nz0emB0H3Ih4jkQEI1wyBgwxuAPNyTrKZDB1xJO/QHeW2HlhxlE2sjEbI9WaTO+
A14KkM9caTx9dI5XxbxqSDLwlCLXTOKJ2besS7FB4OaN3oB1i/Tv7e6kYICGir2172Ek4J9yYaQK
JRg0mabt/wv9B/o+khZl7/ZKE48gzmf1wV8EZolGOfpHHT0HueQoJzS/jKOU1h6ZJvupGqdvMFFZ
T3uaOlSW3fBZ2/jsaoXJf+llJXbUn2FOEtWLAbj5Uc+5He0o8Q9alZVf1x5wI2QCquQ80BJEya7T
tHKC560NYA7sgHf0hqIkNWitZgS/z7IQUKc3bJtxh9ifiTVtbYyELF+/6wkaSebe1WiTqdqVftoL
V7LmFx/kkyf+SBHUYM4RGbYgKkX7fVgwLMpNRQPMnTstC/nQ21//D27SnCowl6jzP9jTzuEQ7nr+
XKeB8C1wnjmV2YL+8Uvq3wqV7vyntLVhFSWfcurCiLsUbMfElhIAOTjVTCJ/8i6+Niwe+RXDs6q7
maARiYbaz1T28R3Rip3KCQGNH2DPlk+s/+6BgnbLv+aiwdxNHecY0mBSktNU1U2GDvsswo+R1Eu9
wHb236xiGkY+z7LihF5hQNtHCjBLL+Fuk9iowQ7Bu7OqbvcTqex3foKB/C1HvO4q47aTP3QHV/Nx
GAHKoAjh7wGq3pl9YYmeB2meL4TEOs9U3IpcM4Zcyj4Fy0kl9UNokqDX2z2cCpZY+8PY6YOWFr47
aa9K+JowWkgvqIRNbkKVa4BoXX07M40+wOrhWrw/Y10sixRFsv7GdLErXw5EZZOn7jVUoYZa8F7d
ebLEWyugsW2GtHadqm4VpN9wp3/xD82Jg2uCsFOfsJpf3XEpAgMTxnoisKbXMCj4lYPd3Iy2j0kr
gQ8H3wn46S6+B1/VM/QtrRidgI147gytA6EXsKa1DyE7OPZ2ubVtVhNjC49mkZf4EjyVZLBHt+NH
HJT+DhsO0WdQhF+3iX3FqfdsDIqqrPrKXN+L0duyTEZYw+aK426ZzEKNCZl+clIjjE5TwG7gBZ5P
EpCqtV2QTqzvwzTxbpoZXQ44B+rnRZML4bDGjJ8WOg0NfzDY9C8EnKzNISDZCoG/iy1Mfqz2IJnV
yOjBuzXjYHC6OhQiedKBBbONslEgE+F9Bei0fAH+WisQte1HPI7V2+34yppibfXgkot9GdP/LdAN
m55qtjIitGajEYbzyg9gzFAihLnDOnBLlQeGfQ4ZwWsoX1SXR0ipy7WlcCOWj6EXQDRaSfRxHw2B
WjOlESBY+2BobNUBLtROVwrjRJ/p7qkq692J2+9GOzl2SYuoqVrXw2FHusVd42X9r7yl8WUcRmM8
jlhQR3zaysw8yyffYJUhG9c/QVFFW135w7Dt/yFWQ8tzc3Y755fPp2jm6c53O12Yb4E5wfkiU/hn
lnxaHcFP3OqoSYr3FhYZWi+TvRCBi6SjtHK7jBm7epOHZXbbxdHRdcs8i1TKnQjuP4Hd9bVWOSqi
fFMphgpQoNWM6+NShWN4QeR2M220npCw/K7cm+/EDIi0AOkhEw3Z4ipfqjqxSMERns21yuOHETix
ZQe9a08ESdSfo/nzbMflPKePGihPJvi3Mhjyt6ovriFzlEuDzstUWuGpg2lsze8Qppv7T45WpxMC
fdiSBsy1P3XyamXKjBvofBYweA4Q1RmQYQC2PSKZpxiUfNjxhErXzDXdBEs+lK2JN0k56qC2zrgd
AvJXhjLrtt4pMAuNMreHw4b+kMzhjg4lk3pcusVSiHfp9PZEjjkqPpmaKtmWfVn749vy/rCi0gHv
LivgvN1WZSCAUkmlyVS5g2x/iCyZ8jzyTrJ0Cnuzz95qMfo7twTeVxaZwyNFTRtdE0+oAZ2c6wJr
nVyLIQlCWjtcqlvrDJDyAqX93tW8lfnXw4cUgAjA2lhJqjfFhqrU3A+8xJAD27yOJ4V0zw+QKxD6
Iu/+q1yTitdI2WkN3WfSqIp0moes15mw9abJ0C2Hmx6Ap0uOyqtChg9nFo3xsK452WrtJizljM9+
QI8r8Ih7pkrMFh9MHVvFplhDQaQp0/hF13YcBts8tMVQrt4ZY+t/e7orkjTSBjEaaVcDX3by9EIG
P9NAgwz/idDybZDDPnGGDDBnSlkuDQNziRKDwAWRjTqO++hKGCPg5p/sOF9QcKwj0AzvaBnFbL+o
bKTeb8VZlEduIryVGM1xm0PZYrw0cnZCcG1tTfbLoe4M7B8W6txvZjtfrRbWV0+IYIGNDjlnYcZK
g/kwWQtBaXnadr9bGvl1WcRnIWxZ2ik3v3fJvpW2A6L94vl9Uof3x3ztpsgtjuwh7/Zqr4m4at6I
T68hb1Fa5hP9xfeiFgf9COlMABUmhyG2aBN/fS0cO1R/dsDM3CZ2dB+Z3Y31xwm2o2FoypmKsFNo
nBS/NSxCr9DeMKbRgYvge9+3NF+jQaW2anjKiaPQyH+FLjqaqe3bgEjDW1ZphLjnb/jwkKCP4Q/V
9cFENckk/YnwBEImZLOCJ9tE2dNMrYN/ZrWCtJpdpiqA7yrXm/Fr8Q7Ar4iGUF8qMY/YZQpl/6AO
DyIobjDMVi/h3fdpTJS3dl4O4X2KKDKdifDjHRT6+bOy4sw80YEGHwONh/jMitUXh4zK7BtCTpnS
4KEgQpVdzi82jriADPcKkX4Zbj12vqKh3/o4gxsXvqX0JZYaX81lD/HeXE4oF+uGIgFaCVFLkmoD
NVr5jjWEJ6dSbiaODR/ynpN8E3QPodi1GmOvrpZYNqLGAGaafUGO32/rQYX2KgpCohYUyxbkmnKe
WirarlXxbIX1oxhnlW2d9TbdMuKJ5o2lmADH92kxGlPyHqRm8TVaiAedtDePuAOtEao2yfoD2GJu
blvSo8LOkL3iv160N87KnUcWkl5SZCetBeCvE3+yM9R/1M3+sBxFbbKrkQR1Qq6eOZEFbzaBQOgi
B5ypaesBdIW3tYbL6szBrKTs1LhyKgwIM7RZTV0LsBVWIUvPtz8YNCUzBeekhbblA2uQEqLVMJGQ
MbQZH0pBDS0/jJ5hyAAtCmw/TXjdfbD1Qu36VIrdumNabAahoNXOeQKpzWRZkMGNUl8i3iJBSaiw
VKhvpxsA6yGI1dPJMyq1gaCTb2pyVwBIUUcUgU3CIl9fJ9PUuk+zH2jdbx1xeNE3jMO1ur6w/JG5
Y3fJZD8G5SAQ9OBUrCldehdLsBlWijtXghdmsv83oaL39eY3MsPxRn5TEuNdTC2RjDOIjn+7EBeO
i+t7Cwpo/kHfYOL63ZHfs+lWOnqBeCcd5pkX60Q0ZW/JXR/wsD+4N9ba9ZVUXki2pCVm3rU9gwdr
u0J+ubDNz0hmjpLB52CG4NWo+TjOpcT8iLQSkI9/Gqj3RK7hvANvYsvwhbnS8+OODLvgI1AK4xTK
Db39tQnyDqbzvfWW6SU/h9GMcnJYrBlhiUvhzqgRkxS2dPunZGlZcpCce6FXwSpcHHMuS0CM3Msp
viayYdnCWzTkyhyI2aeaE2pNaq8lWDfWlEY+LttzdWlweYuzV/3MFNYt9h01I1+7ebZLNPA0gmc5
m2jcDEBDsGuhhz/S5beeJCSkXhCjRTpg5nsRZWOpHL8/9EtwC7rX1WGfJvJyfvWvznPF+gUm+Mmz
B2JsXUeD1sDMK1WPcrA1l7xZzelxnFf2gRaqUDWhMl7WCrXu2tGOWevymlnpb/O/E6S1yl7ilX5Z
TjNAo2g9vx3XnitqsqfmbYV9jiQRfstL4duc4L0OvmOSc73Ps9dP54mIOcGWMiUsXKQqRGEdc9Il
oUruoLu8I4WPymGSl72vA/Gp6iW14crhLzF77vZmShH1LRpIW7Zc2paEV7GzJ3B860hDhU0Bs2CW
rczu7t+9ggMFUp9BB56BA7zCpTsL4cGzSLFu87frKI5GtBH6W4/Fg2EFXhbi5U6LQ56riQtOzHEB
2tUcPWCG9Xf7hyvukJ29m4SEdoIGjZ3ijwKZftN30pN1jQC2Zi2QROksmQCxiwbO7mLXtTqEZv/t
hHf5dp8v2rKioSGdWkvRt0FA5xeZyEK4L7et5ceyeAUHL2TObQ+nRS3vX4Tu54MFdzK2W6+jCO1z
1v/6OCqngrXiuvqWiLHFdQfaauu+TGQIa7qyX2+Q279JjK/uQjFApUWji8dGnxWfBJq1QsXtSpN/
Lw4j31hQqTC3OCG9cVpPzYE31OSBSuiLpjh88bJ2yMxgnBM6F3USAZ0Apj/Gz5TPKDvlGzEMZCmM
P8qDVjpvVu/Du8lkCS95dOBaDamBdwrpzJ436zHZTih65xc2Oxfmve5tAlRupR9zDkfVcAl2djkl
RT5jDgIy2dXY2Z8uaxoNYOQu/sCJWlJQ7UzF4kHAPn/RNFrxdrEeD+sOlupQ4Ko8LvFItSq5xJkf
rRYLMQl2h6iNLvxU3RcXvwmfXxvSc6lW8Ml+rVLoqLdFsOV/OFJYW4skYKdVRKrig6fzIZ5I72Hz
M/ASIQslclNMFIlwktmOHImjvFyIbsPdXLZFrb+M2jGKB3VeWtnWsZMIzmil4tqUWw6Me2TZ0uqr
Bg7azX3FGOesQxnMZpPCjBahlZZ4XDBE431sm8ySI4cobSY3CPqmxriXUgWFncGgRm8O8s1o4ndP
nFDdwGhfaGbU0mtlZCMAgfTb5znSs0ZmN1U2ym4sQuI3TicnmKkEwdr8pGMl/kV3skMGU3/bA8Hq
bS8/lh5IU3bnkGra4AtKKeGdd4tQZ4mmCgY2YdrlbeJ2DQ3B2yEK8OQwURg6Gkp+YPke5pGMwwaT
q8s6mPxmGgCykrhsBnX6RIh4GMXvALDnT2T/HlPxpX9AM6+am0YKtfFTKLqr4RAassQ89WBWAb6f
2My7RkwWftSXDfRlKXNnU2B3XlonnKtqR33V2xHb+CZFC6sKxuP7wyecmMxHRDMfw9bcjnsDOVjg
irakL6L34hN51UBC7M7kqMdqyH/nXj+SagyKSJnibjaceQPTJk5B4R/LqTpmFu4A2PveRpySxz7v
C8H9lmCc8TtRtEaXckGmxg0wHzgkhPg49T9eE/yXgXMx6n/r3sPY338gc1dRs34sL9nzTcRfkln7
rhJUHOPtgABinWELG1v0VUh24rMPNFyHWl64mYyI7KVeqdY2/u8xZke06pPJcBtcBH1rPclWsa8e
p8Qh700dpKF5wJFm5SefvU5igIVC+0usOftcZusjJ/KMBLzrXEfxqdf3oQXXZ6h8ocSpR/GF+clR
smkV4bifUTb2Z4QhlojdgXBDuQtH6yUhCBrg49vOu3d1nGxkykPLjZzaAvyCb513gj2+ia2953VT
16vPP8uQjoPYRTgL8sd2p18SD5PRv2o+TNtfWx7zHfj0+ndDf4W4wW8ptKK+RyOIf+YOfXBDTnJp
Q6wt2sAvzZaJzb2yNpYnTSNd+j1Jx4AScYKmHItzxOOTl8EQK4+vOl7oXnGCe01xTk8h/AHdSI1o
n3C1Bg5VtIZV/rQNeIySVYHuuxbR//wXZoQzVYihV372ywmM0Rw3M19AweusVoDWEI/8sxJoeA2c
KfxU6Nhuwdb0HB+BRBCbTCT/L8TRcJCnuUOnvB0VXPAq0RwRq2TpTM/jUrPRlkM6bkWX4NKSxhvZ
+K0/TjIrSyTFXgT99YLDkx9V3qNSIB4ih0Qfzx4T6nPFxone3EoJ9F5pWT2sFz3FurMY50E1m0YH
2mG9jBHgm7X/48jQ+yiItvHLkX3dOC/t0x59fVxM6zWdP9mX0EHV8HqqVoxQQknFgbIoPrVwaQMW
8ahw3fpjIl6mmcnFCQxveHVwol5wSlkz7wFh6q7nDKsizi63SCvVwD8S4bz5ibhP6t9qZpYz82Df
qHB2FMqI/BFdpnPu08CaO0gvedaZB/s84UxC5/o+U2yNUVpGXEZs4um2iA8C8twVsbTd5fnlBBeZ
vJpjCMy4urZ5eqROPLfII1noMNtaCb5XBOB04fhYnQCiBMr+c6d723yj/xQkX5Gh/mWuTulTGdo6
bxIaJ43KBJbMH66a/7djTDp4xb53mygYd4lj5p4S8+J8hdS9mhLl0tOClod0tOsR5d1oXwjktV+e
mYsKAAbf2Er+kvDWsI7L8m/cB9x7Q0WX/PKTXSa15PSKw+jCArdcy8fljMZ+9Rn6safWKliw8lIA
k2pyrzHUAtgDQrhLfYXQgFDYizXvMGs1MBrJSNPM82/qZo3RoqsJj5WEJDIK4LkADZLQrBngH03i
JEo5BbI2X8fil1imX9PWBmzR20i/2qciul0uwe4kofDXJrEagEN0U6hR0NSt/j7TYAzAMKO5/WvS
pLc3Xiq8fEhwnergwYNkDvnProTHYufS5PrYwaBGcR+CWenvXrwfFOoMwFLwNUs/B8pYYtRipzYK
owN/xupvJofTkwPjGoUDIvO+Ksgys3v2Wkq8SigVGVeGODDuqh0vww7qr79y7RmcbJ29dTNWv01P
nQn+kyemvBXaUyxEtWtDtuoB4WEVtQygyTpMFc6N285vhZjJVbWFFLWSk15kEedxyMnw9dXNFH7h
/okBZEirgve33A7CIsV9IKN9epNC1u5L0NFwzPhPTTMmDc6CKJNPY/oCnKm4fvGmvp4VpaKtOnhV
EkG15TAWqcpPwd+D705li3PFGuGESwaOQCp3f2tc2IITJPhoIW3sp5eH/7WlBcO70jUgyrZgQ0Xh
zvBuzvOaXrqWOjqC4h5V9Ivqjqkxs9meVc7Ujnl9TPaR7DafeS9GDKKNMbBaxUKLfcS8PHTJofwL
eohJPkBpJYQPlklFQDTKlyUrWraBUxy2P1h6E1oqgGIs2WlsFhwDQP/WnL+p0ofX5u8IQtMm8I6m
4BVjFoft6PNc8uTIaVeeSX15ph46+GoUi18YN45+G56kjz43D283FuflP6CoVs8A2FZ1m18yjXS0
Y5g76yLgAFieYD5zWdrmTgJmvs4/mpCmrgk39vLqIHbWfQDC/aytbvYOjM8eyg51+g8C1jZsPlgo
mO1HupdN+L6O710DTqhCBeUfSHljZ6SmyhL+QSy9bebZjE7a8JyH1wqUKtwFWvsm0mUbSLmXwrwY
HtQo7nMTpEAD5SmUzxZnco0CyngiINWpf16qDX09vHn8JuKuOxLhA44qnwCQxhuDRvz3EL610AlN
9C56zgWdjJMlHVA50AjqYqm7y5x6uT+rh+NQ2OhJrdbCCCNPKiKlgb2oKlrUwv553bH4sgYvR4Ly
zXTe1TnoRvMUMEM7GagSrkUZ95daKROYv10DDA0flwecZ48FCwnMHZmyn9MfFkQWcHscbPIoYfhI
H9ZpZ8WW2QRuyxGaQjoCZnxKXoVZRxKcZfZwJfOqA/7vrww3FymG6/i7zlsGdU/jLc6B22LE3+OZ
6tapQP9acawlPt9hhIUHc32DwlouItQ+ZkTUY1Kcj293RtJX+BKsY9w8EVr+Z8q+EQ99Q79lqlW+
ygYQwtC0ZAMIAHPGXSRDfbXrDMaoVOZJ3qDLo4BtxYcb/ChQBQjUGpNUuyeT4x9s/IlJfbWVPLo4
Qn9G18Dg42oDr5LjKbov211I/Z/vQ9SASGN/+tjkJzGWC3BtCi1/04HWmx4CX4vGF0k2T7wkPZ+d
Bj9oyT3zbxNG3OFN3sjQ8xO/fV644E6/Ed4cZ+RkIC5YrOvMq2LIgaUmD/VqM/cq5q+KI3/4uoo3
r9kKCOmNiVqYoc25DRtl5Duhi+mEJflr9H/sa+GFA2afXlKKJomfwIgKKfM35pvHps0mUIhoUemL
CGSR38id0fiOtDRvexUN8Qi6ZAMEJKxJOPclgQb78gfrWnwZ/xGosehDnqK0p5t/QudIzRj38eDQ
iYQNUNw2fOo7WTKrTOACMs0ASJsnN1J2YE5X3/rI1Ub3GCiKIXMs+kBfLfkpUtMy+2Qi0rERxxDM
DjemOZxZ0bVDzlk33B4gO4+RseQ5XPqcMNrkLqF4tOTZdM6CPdw5u/cubw3r9s0X/nQqGRy6efZa
rdskK6Fdp3w4fYcjfXKj0SJvg1VCWDzDU8wx1qlW/bx8kSbQeLExxH0apy/CgUsHZdCSVUxVkesU
UgfgFxCRb75SNVWbRC8QWtlECttHV1fIsE4ZC07mgyMUqmO+8zCSO56B/Pin2lHTbB6tNgMpSS5+
e/bIk1qyWeZSv/4uPYh8ZNfP396O2DjZOAOOK6D+CC/eS0oWF07cK3myO0bzeT1N61aNujog91fm
p+e3BPIhQjM3k90KE5dp1/vilN1GjbNy//5kBYlRWJR8GYl4KrSssy7R+OFPRe+DyV3bjRA7kGGg
fmyexL8CRnN/y7YHWv26YdA4Vy4VxnDSb/dJHWmf5ycHSYcoWjCGB5FdttieWFlkkkd0j5Kcf2wz
lgVVc451oBaBL7wpvvg4G7gYWyIizZZAOb6R67W9S4rtUnIEZxLSVkljwwBQCgUgRJ0kksJuLPml
zbiRLK8rn5K5UYdLJIHyivEAt9FUCSnUym+50D98nA9MHg/FpdXqyQAh2KQBA85uvwa25IzX+9vr
c3zyMMPpdTyyEN0x7EP8unR76iN5hJGrsC2aOBhehAKhfp/EAx44Kp+Rp7KQNI6MJaVREjEGtGcD
YP55nfOT5dEFf9sVDobB0G2pjUMIvuhOSoTde7vnG/kjIAJhZ7Y5ZVGtEOP/X06DB1Jy1wIfFFfT
rT4/4pz95rrIacgfT7IjIqylGPNYPzHrLY0wA5M6ERxXLedNl547aHhhKmaf/FRq9NCPeyaDmuNh
78UN06ejrio1tFrUvEpAwkE+sl/6mF3UY0eAHM0+96+p8QxUpYfyv6QNiKLbOnRwEeSKl31yf2/0
uSK3mr6q1NTNUAKtlXtc2pGLAk/Y1o/R82veflzGqUELj+SVWVHa41WjRMnHIRSHMtV4hBmZsO0F
DG7Kg/telO/gB74zZQ7edyyxRvCBXTuE67qqihSuMnDfN4dBqvwyejsPFYxHMsO1BBGKGh9wUsUj
9x2rbloLT2N9eEMqhZT6EgfrDOyBViqR44rZm4B1DmfL6ZFda7YFpVCjs9w1BEDAlGMgStSlknJD
U3dfolAEYgenSkxpyoAhbip4yfekMBjxXw1q38EP3IkR7BAYUBEBfv3hwh15VG26hx4iorSc6VQl
oqAwC3oR2CfetpG0aUquWDt4yXNtHO+/YYrTk1hOkaR/gw6RuLpb/SD5kuxVwBCbKmllRhtL6Pnn
RXzFn6io+bdXBj4Ypn8kmtrKlOlQNL6lVzmW0vnGJJyl0O0evdXY2xG5JQIN06r8tpeAliyI/uhI
FM6dSW8pFIFJIY43QIo9OKZ+BxeGQl3DP8sUyGIKm8YZIrFFWVrEJvj3awPnzQcbybAR3IgzU2u/
JE26Aexdfk/F16julEUecrNXlwwx7gzg4gWLzQKR+iFqHkhV/vqRarGWXh8LjjLAq+5W9t7b52Wi
JB0j5Np0mCysw6Azdi1kPQj434nM05QvGdMIfbOjBLjALFH2LXPBqyG959qm2SRLxJ6C/4PUNyd4
fUvX1ghCFVYuDMuCQWl6sbcy62HqhA4NmAADgidJlHUAowrAuK/qXYSIH+zOH7BQv4Tsz290jsx7
HkHaE8gJ+sY6jPNhpfBYEO+j3NfltwBBHJkUHaLD76GRRG1yUPVH9R+CRDYiWuOd1kALb0wSCnlO
YYpOEvsVAW0or1Ub038AKz+IlYBhDXK2gIUc+ynoRJdircrHnsuuoIH5xMfLhRSk5DvUPr8Oi6YJ
ygLtC6yktMr7jLOof/cdufmekoKXiiFEusDegKOueYlfmsnKqXtmmoWa2KVrpNk6I/hb7PhJhqIS
+nRkUqByvNvIlCmhl4JR8wvwRDaWZhlrrC9HBPmt6pzU2pi851O1VrLPZ57rhdDyESe8A1sSZE5u
55b1VCP/dSYnoiEAaj0Q74WxCFYoo3hfB3aFhFXCtY7RChQJQ/IFIaJghjehBqthLe+gcbnwMvRJ
TLEJYvoPsomF8Mt0MXb9L0KSLsR/61AzHRajT/9+PyoWUZgWImx7TQK5EADCfDxC+ZrjrWLzo7cZ
3r//hqDx2cur8hhYOcj2ppoJzf/vngDJiQm62X4a/PVwSpRLLr9ChJGecTFmovDHqxAJH50jLpTK
G6z8CT5M/pBdCaFUB2qz/NyJf9ysIt8wmoHYkcu9tARc+Ta7EQWki7dGAHtDAiafjC1Z2wr+sTg+
rSMqRw1KQghH2Ggv4WWQJxlIU4gJVpG17NrOw/Q2GZNuAq8naesdUlt8194GQha/k93sWoAVC8Uq
Cr52ZWU+EUeb/fki9yghdRH81F2o2zA1lvZcGEUcgMRBsmmpHeT+hEM3W2U2pPwIAipsMKlLQ8cC
Wjo8sJcL50gt0oR6G2Lyl0/TrNixMwOw3tnaDBB6yA7Gw+3mb3ZZFh24Nv2LwsMR8u9cn20SSQiV
m7jdMGopBGasJoF9jaBij8QRa4ZOSqekrcRUuErY+Tax8Tv7MgsIwdZl8EVaoHsaijR12x4EJSqs
p+UB+VtXSWUGoTfxq2KrKUQbuOj2xBtKGytlsYkY6PGUX/wM+xobSNpKzDE5gmolZE9UFs5jrmmj
CEguYUwbx7zstTGoNmxZ18ywNRXuMuwSY86LxawVai1pCHNY1u3W0ocoDAkzOG51Mr2QX8wyItRK
WxrmEdgSKkh+Qj1oDOcrCz+4V3EMjHPxFgkLOPl+V8JDWKdLwabql4oT1abyYYS31p0N0xi3ktXU
EYJdTiVvd30jVSMVIV19xrfr3TEScqsmWHJXi+xeCS/FaKAkxWeEGx+zAw3Rf1DNcxwam41ex8Um
IbFITn8jyxAnvwg+zHyz4nx+wgbz9O+YWDdDz/g65enSmWx2Z4s3vKN/5OxijH9VIEulOSISQOj8
cGqxiznz6cUamUYUR2nXU0i0Iap/Y4e96B9DS5/f8ccpIGYv90WroinV2KBTf9BGi/SB3SkItlB/
/A/YjWG1GpUezEz4vtbWYOTILWckraexgjF2UkMbKW46EBicMDYe30mWIGS+wNlsPg4D37HV4fFA
tVFg7D0wLryxugm+2HuBmzyb26T9qn/kHhSa7AyFfHvcPCs8b9nwlqyYBoIZeW38v36AQnQ8Rx+a
8omEMbsfd5EHlSd356b/O05KpJ7As3e34WWU71it8l5gxk8lgEkX2zSKTD6RMZa3+aGr8imA33vp
C26dHyCYNk30+MhotRAkBzhVawwJI5XeAT453qZxriyUMvy5Hwifr79qRMezlAvbRDxHkpX1vYm4
uKGHR8omPhfgbk/5vr5U3zHU5BDfvcndDEAL+UOigmmnqjKQ5e1qVLtDFzXmr6Cem6wTM8J5GQhq
CUzcL0nSxonjwXNfDctbJWZMMnJLhXKgNguVRdw6SvLEXaBtmmVXVokvEvwOOfm0jhfvJ+wSnEnA
upKCmpZib2kju8htFsyO2tg/5sQ81JmEQBphDeZuUxMJ9BAm1gnYd0iqw9QqKwn3lL646jMpXC08
ut/h3RcF9/2oCLlgFXvqmyaskc16FTgUXpdj4/e1KyXSzOJrn28uDu7SVHxLtHJceh17t/uv9tzS
KEBt03LGQsQWDNzh0s9f2jheJC0uMgGWbet8XHziWfR3U793JKeBfeal5YfQskQ7EVyjWZAZTk/c
8Lh2oIon8IIooYjTtBcKH2SIJEFsTVTjgZD2OxqTZdllSVtxILAfSqy+M4JQ5q3aq/IhJ6wnZKGa
A0hk5MW4atPmFEQcMLTMJxC+OFayPDI7fFaFgvtZiVvm7aXU/yj6Dh0I+u4ZihwOkV/IrzfHR1NH
hjR3WbYAwazOI81xsVfx5Gmzn2uuhfFQQmNjVi6rUYNaEaE1C40k51MEkCct0Ougimn2ys+w3m3I
8uWWpxbzu37GUpHECNkdObZZQf+ha5NN7LQsfLm9Hs0dmQykrhW2+sC8bo273paUTb1hc8RwI42l
IHADsF2E3hv/FoQ6TBfIxu+tJ57NdchlfpHyYzMSyewHGExac6JM9k+pPebiIXlrEn1fTJ9oZAyX
9nxoSokZ2nr5n7E7VdUeEp6bkV9+34gt2MpM2hPtD2omof86U6OJ9SW10UsGBkg5WyYOMVfgplM4
z7Tnm5nReRnmiXAnWegsoHbwndGhodnJN5t7OhsaagZXPaezz6CZl98ZXn7rC51MutWL4IIbd1BC
HS74XcwsX03KnV6AXaLwOpcJ9cmKlI0Zg9BI81GPimNOTA0KBSX3Z2SlQ6X7Ny2m7Y1FtWNexQH1
4NwezpCBTl+B5RiWJqM1pVBJMFnQneGCsKGh8ElMPhvLv57o0AGvJkkAGA5HOzW239Rwr73O/llX
jQMKLdMMDWMhkPxLqXq2uhYglWsUiMvPbwwD0bCKPblqxTLR5nmx2RIp4BhSHMMMtko2XHK9IDkK
HSXApcZKXYoREEY5WVj/R8P7RYuH3s82YzFGQl4Df+s4wAWa/Q+QJtxc+zNztshZaTMIPpk5JkOO
+FvGIKsrK6JlhHfPG0LvdooIzTnpRuO4w6SMgHIh9KR8LpNq2g4RP9fciLGE/RIsnhRQBXaR8fva
MyKgEi8ei4+Ywx4QygeCl5rGb6JTM7fuVW2FVcezkbtcy5YHG/T77cWIPHy9FuXx7SxOWusiAwMN
ArSmuO97pJOQ1N8/tvvFxqZleUw7iWTvFh+HizrCW3aYWF92jT+NTBL+gCWwsM2P+BTvkovTnt6V
d+6Cbtfftvj0E7VsveAdldpqYzOHNJU/vRUpjTWu/GAdruTcTxVDeg6Er0GB6oIMg/KXwjiSRyIA
zIdzqV5C/IpfxWF2vg08UZ/vRhFLmbgFkqcKonQRk1bg6sispUFH2TGBbTJT5FHF/JalNhou0qpl
1wU2CyjFQpwUThpNgJq92Q5sbLyMo6wuF1POLRfxyOQrM4d/Yx54cLHKmE1fJV0D8FthWZLnsAjH
X5wUvr9Av1DWJ2fhXbR/Rr+fLuMdj/WPP1GoRYJp25aZQXsj/VtTK+prGoJviQjIih/RxZsa+Zdd
g1jfMgzEyUaoHSL8bEUMWRlc5FohkOm6Xm7nfqc+h2Fgay5Lx4LNphYN8/tsusenCt3pU9AlT53h
fdov8RFyI0Xtb9FucXqww+CfuntpSzSpBsahdF3GS2eeb2eal0y2no3p49MaQts9Sj2L8Kty7HAf
Bsu5qz8c/SyOamjQwnWptlphSZp2FdjXHoKks7lG7Ihynt332tCNVU9k6xKwxoE1/scF2nFArauF
sZAQBZ77yZvB0J9ZU5l0U0IHViHOj8vkJyTFLblQ6hNOBVB13Fy4OFVDqwsCKGKyMpkZUExDMRwn
BxeGKThl2eXUrzAT1fMyETUjiiCbE1qsG1/59NOAY/64x8IYaStV8QG3MhcpZc6/b9Mh++upKqON
gJWZhOk4xmKkRgoGtPZq5vRK3TgwRjH3mr2dEh4oSDHP5Zm4tbJMDGtVJ57bKUuv1r0PgnJ2Wba7
yeOiUkFPlPrqs4W1J75YFIvXS4R/DXho/zS7L+LhtFIynRhWBCqDvg+YqXjWQ81jMmW5Thg9XkZs
ROzD2FzNCTCHdxmhV3CcxP3G+w+/8+neEqDZcFrsbLEpcPrhmw/UfE4BeUUFaNAz7fSLFVx74x1J
kvhBvPr/C2C+qhHiudnyRU6EmprgcCcb7izkN13KnnHf6rtU2aJLwRmWUAuGW50TNlzZr49NjU2X
GVG0g05wUFfnrGvllQAv1wn9DVefNCyW4lNlqiz7ZGapDA5OzD1KTLb3C5VHRghhKD+JdPW6ZtMc
HfBYWmzCHZrzIHVMwkBBgL7AdcBX55mZaDAIv5RqaK67pvow9C33MhxJtFB/93U462iRlprCGP/D
m5Gew6X6W2Dexrza17nqM2Yd1gYQBvF+jOvNPLf89AjocQ8oLGgLJCiZvxn/5bnfnhK0ktTQRENW
NfUl8YXvs7V5YHP4Iiz2+9BP4TOgUvEcc+2lru2Elq1G0ChWgLdAssJDznj7lVyVEM6KfwNr5r9o
SvCSeyHfwXrKEt2Im4ItAukkEmDUXqFp5MPlGSRSDyGzRTEru2m5Qw2Z5c0EvcnGNAWeiAkqY7BY
eIcpWdN3KVMrH2VrzP0MlMj8ZSOO8TXtQWn5C1+owvQLZSmY9kObuyWFYcEmzAvVVNed4hQcpclC
3T012hhD8Z5cX8RgHCPSr6MOoQYcSTeJvamYEN5tKsMdv+USZLNrFEDuBPka6RGXVh/Xonft3zXW
7tNv5i/Fq+atzx/qmPmo8zzVzootFhm6z6jwvihlI53VL1BcEU3pMFs8MJqhS4r2ZiPbtCbFzhp+
IYwcwIgRhOwLCE5lb2l56S2XDUv/cz2r0K5TQLvWNhXcF8B3uvRYv1oSHDzxKsg9uT3QnXOZZPFx
c0+mcpvGLSjKiF9Gx4hnGKUSODvzk9hhURRDQlluj4hY/f+0wuMG86TCQkR6hz+yF4SsGZFhmxfF
GRJcXkKWQr3hC6vfg851Qrz8w9loZFMtSRIrCuHsP1rIrWRlmle8DqIaK3/uPVMLqY0WtmbRnID2
BfMKVwcwXhHGpyJ00Cl3jHqAsMrRcJAdfk0IGLvH3CiWjTkGHf5pdeazH6Si/H2TIIRvhR+T090I
ylChje638W6UajvC+EyutnCSNAgXeUr4Ym80GfnH0rJOC4BPKcrj1kgOidY4wQQi2ISkLcQiq7u8
3n21VnOQEYimlnggiJeok7LyYvZ9NnGF06/26WJxfajNY+qQ56ToVgSrX0Y6two8qo3jmDgwCmC8
Vut/gLuKnlQrzcgnmaUbC0E+AE401U4Dr0tDVAV8xOstxiC8DcIPKsXFFBHD0hL22Wu05cFVWjxh
slNYT36nOH/sUJeiMyMQzgvVPx9g7Cex4csWAy9HlGsXtmpC8321ziQzM/pvb2X5jxor4KVL21PM
Wfe2aIUbhUz8+/Wnp20s32lEt7cuTh0saPd2NDDPSOjlL1WsbKeE2zuwdiHtXB4sRQkKnnS3mHIa
X6cL95Ya/BI4ntHqZIu1tMQuVoit6DWlFXI6YXGNrlJ8ScXDwSeXDG39sdZZeYTy8azunvrSoROy
csyOyHdMh4sae6gitSirzOp2oZn6mhRSiwV+6cSzbdK4CWkuQ3mpajyEiEZ/FOVNTIFkE+ebozgC
M18IH7wk8+ap2180mfSIWbkyyRFW0Vt1Udc9XCEy6r1KDVf+trQNSe9qsoN3acTi5BifMnwkzjAL
akab+Ku0c2fNUEBeVlSCKSPTkVpUfYEY6UqnifzFsFhADdGH591op8TOJIh/NjkM3YMOn/h7PG2a
64z2xabFZHX26Xgyy8imMC3qvewxETEPO30YI6P1mu2bi747Kr01X4KWEAQS6RViRAACiwpRtL4j
m4Y/QfwasKV+SYIj3hbqxrutacs/+wptXDQEXfFK91Ydh3IEzhssRd9fOM03RZ8JNMgmcb3cJQB0
4O8meLIeg/jQuu23iEErDFM2MSgiW5/gJqAUyvGq8uhX2khloM1ftGyUPn/tWqL92Yu9AKCS/U38
94skFm7dh4w8wlpa2h/Bc21IlsRDVv6+f0J3H1XkWSYUye0IOMHPCyOjwL3s/y8DKjRKnsWE84uq
7Zg2Kbhc63XelA9Uoi1wx2UTQhqbP0/juiKthYK6RG5K6AW9h3qhlQwwhWWkxFHHKri7VFzJ+dEv
eDrpnEBeNa3EiBLaV/WmE7ZJgTSEGKb/xUBrDCNzicXBYxOdL4w/65qBnp9IJ5Dp9NFtLoXVRpq6
NNvDP/v3nTN/adp+rVH+jHsaBbveOaIf+e4KutAcOokIJcPJJ1mQ1FAx1TiZoSIZGgxJeINI1r+r
ncEw3HQjrYio9GdsRn3G3qimgsEj/hJ1YQNpJZlivUg5FCUdZnF3lk8HqeGRCGbpLWJqTdmtZo/e
3vau60xfgPVCtHPx5eImTc4FJcAz9i1ZrL48sM6+brtaSfGz0fxBTTylkm164XcR2CstzkeYuu/J
h99xM4GZHRJordAyCpbatPXSDaU/Yf9Z19yiQwp5vWDucdf0UYD8smp+4PJETYbaRva12d4WnNKK
/JXExvARASaJSi2zm063GAqpAtHImGTIJ+7DCKgXhPldDQ9prG43TphiDUKDHkJoGoPKCF8y9OqS
9sISH9+5QQHlshWve6zTk/kCpkyoB7HNTxXDHJN5sRFNR1ETiDMCnwqdz/eP//DPQIjpnYaR1Zh+
gjMqOG7CN15xg4FyxtV+YCHMCVdLmtIabWf+gtuHJeJnHo4MIZuNpgZRupynurTjrhv2swCVpPuu
YBiD3cFggtAhJBFTAvJZ9jiRKXUuoUuxqkPGDYHS6Tg85sMdpCfY4SmnNnp8DE7vVFmg0GVyNd9R
lcQ+Wb19zJd5NcTtcnOKXyIhZSbiIIFdbGqmbyjjOM4TBjX/yTIw4DJYSkturvjYWFpklOA5O0ma
ExuCpQeONj8gNHRmei5SDeD+GbgWS/f/fqQI604g3BfIwcu2mhSZJn57hnC9WNYcNp21jxRGd6s2
17hJGfaghW2zzlMs1Xdo0lbGaFRKCmez/JAqXHlinP/1a9CcUQd8VPpAopx8hcUk8aQNrPdGY+MX
2nmX0rjNMUu3oesh0CWtiC88hdXAh+4zTwEuzw159fRQDy7lHbS+Q3wV6kUgc1QsWI7Ob+GfXQDZ
CFtJLsfsLRizvkOLF4oCIXq7FZ6SJuOvyoxoXKL0D/14sEy710riROVsgjnHS9Q7eV0G2ynNBzXn
ITJ8sC4Pvl6ZWPRg3JuVYJs3bIJ55uC5HnmWQYVaiFYpDkSf3UkHKd9lLX6o7DYBtn/1x6RMewum
Mpis1n8Rk17eW4Zi8HfmlFPZ2o6Xa67T2hqq8Q5NzkExK8wrW9uMv40IDoQXnHQ4cvn0M6hhLFsb
TB/ZUvvgMu/SRNphnvCwcLvEfkMz5cFWeiDqLBT/PaIfVMtWtw5VVF2qPXlwsr6ROqhZlIZN5Qmb
OoM2JzYuTnwEseL6470FPzPSJj1Z1/Jej4rWJpnNMQljS210aT5FVyqDkKMjM4To0MelicJ6PExR
LP4oOWVRWQziPU+GMjFvz8/Fqev9xy35Zc/UTrMInQS29YOsIX8EfMI432vkHXHlgd7O4Kl+RPsS
Y0P+vHs7JXWFXTBKm1zUCsO82Vi5tjcHBnrSCXBQrfuMGX9P8zmVGK1CDJ27tg4fTJYE+DbhV87n
jcb0nBYLrhvpvczPegKxjB4yPB9dhl4RpjiN18n8bXKf9UTFhG+bHrEPWCNVjx6RNRc8RIkVNCOS
9vjyLyUbfTKSy1dslOlycrZ0oNmrW7/ANqQotRNCG+i2e2fy5SQpnUu5YirMkTHOtw0I7SvfrWFA
wdRUJ+CAu+gkjis48tju7EHUIcTjEioK8mDkNDjir3vKG83W5InPCzC/3vi7u3ST0arQ3F7PmXp/
90Pm3XsB0npn5ZeG8b4IOWH6o4lACYP9vUnwNhL2bejrPU3Z0kjmB8bgQv2C9rAZCc0boXRiUzty
8Be0rtoirvkIgHj4Ah3CJpEfQnJYp8/Itm1rb3tfuPVxvscNAxt04Mucd84jwEBuCUYWjNUh3l4t
Dm28pcS/98BTCjLmy7mPMRD/OyPIa6AOHGSwZBJfMGWIm+C5njQFcPOmwStH996RePuxfQ3ZOPHc
yXNfx8WbiuZZokHp+Z66b+mYq0MAa34gPi9Wjn+kq68T0jUYq3O1LCZH8e7pdTZg20a7hLbp+ZDU
6TqTKMsYfhfX/71ZU1bqx8pUi37w1+1s6sRmYlfAxZE1USrn3ypCdQDcQIMSAOQ+C25TJ9MmVYw2
i0weRBalNFa7bihZDM4ciYZBy84hAfjLt7LwcHQdRfLYn+vnXGWfKomSzqS0zdwTZTrA/QPdXS3r
9JrJmHr0SbxMJ8xb5WyB3m/QVRNfc3uJ3KF29HL7vE5bGfJ9PiRxuWj6bhzyLYcnohAWjsUKxs2H
P3j8KCLKb/WATfs0ZvkcO8d0u/gEHGcqBmB+1Q0q5LpiTk2WmhloIbPdgaoGbmtnxxwh1P28XrZx
plNr7BraU8LOlwtdZ4BJ50rFKuGJQ/7NwfmxVwERzsOF20X6Ekdv1WlMJW86h0IpcIgLSnVPQUOE
kCbhGdxJnWXQQLeMvKE1Ucgth1753y6/bAYYkV5NLBHdquzm86fwNdv8NllPf1SN/2IwAvRoCF+2
mDH3Yohq5YUNGGUSCfq8G0JELQt3CJ7qcos6V/bJI0EfHqwVZjCvas0/zCLNdSAiODUJk+9xSs9f
nK/4xDSRa6wRAUMclefkW6mH0Zp4vHCQvIT3164A/QD7THqxl+r50KVcrKpFLUq0pRLml5Ffsqzv
fGr82PNStunEyw6vbROEzp35kYCC/qT1ecUcemnM8nSUQ9MmiZRfcXb2BxMSXtPshhQZom+CYYQi
L1aKMEUBzi24n9kpzbahm69OQd4vAivW0PJLYOXus4AN/wBXgsiRMdzg0mZfRo9ivLgJHfCrf1kl
6RyJLUHRZKIwkKSoR0vyan1ru11AviZEicypV6DCmLPx04KdwOCrR5uj61vSCpBeSD3h4LaL86Gz
IBr6RA35htPkNoxNNBq9/2LITBTPKGxYTzL16TxM0vJNGbtjyhikkXLXp2np7St0OaEFPZh9mnHN
oYImNizPmQaJdWTv0C4Jq0st2qebRFNkb7BYi+5mxMln9mki4nMnPvffNCgNTP5W2UnizY2e8o7U
LAN9i02rldbeSspu2FFMnamgGwsKMpE8K61+x6+tLv5Cx9Aci7cZJw4jvcEndv1b5ZP8qaxuP0Oz
muWLdRk/AMK/BB5nQXmISrw6T5TyWXmdhHKnEOH1t5jryNbuTFi39LbPWRVYkmAQQK/x6XE9IiKP
+h6RE1qz0Q8w4XobyoJQKIXixEr90Pcij20OUQp9S813dUuZt4UJw6rxoZ2u3/3Rbi6ISO+vEPdq
yKO1nWazDT8tI3qIMBXg5e0sAaZjRuiJRLHIJFCFvW/1GQPSN/AZ+Yy4g/DJQPwVZrmV3twJJY5Z
SqekpXJPdDBIPEAETfo20XaaG+zjwfx4JVJ+JWXubvsTRymtkgdhCkyWSzVSZoNcv1MJbKIJVLWq
82r7mIPtqYmB96WBdIYgBZRVtW4D9nbjgUJxmonQDVDLowhYwuhXbKCdTb2NjQ6ttr8lgitA4+0S
xLi8riGeqlJCg9xleG4TFVceTglOZbEyIb4ZGWJQyRVhqwJAYDTlM0hdZAuXGWp6Vb17kzl00/uU
VvKpqcd2dd0LZ202rln4jwCLhi5xMDVR03W/go4fvgzehug1Opys89I/9T7CG7Oc08SpN2rsxx9Y
NxnV3wWiDv20+EYH5xT1vmj3LcMJdHnSae71SD4eTm9zdCEs4Y3m6yHoNKBGc22lIqQRhVE8YLti
6bH7Z45teVb1xFkD9YcQUcqlrvjaRyKCdO1tsWoBAv5fnib9tXY+U+eH5kyZL5zcLtnOo99lOZJa
ZQllWDTgXDjEPyBNU21S2dS4AkpqR3lKrGflConxoNFzZ0HClaN4Y8J/cgEHRlWBGcJqy5CeS0E0
O4eZTM1pGHGBlDP5tQWo/GJtJRIBhxaz+I2wWyMvrHsH3AlEXOqnfqANWqpACPUhQZfmyI40a6uj
farnlyzp9l3dFXG182wyViBRn40pHQGIbd4K8/vJ88FRIwxZ8ZluZBLu1YVsahvfMDZGJeBkaoMw
LVpnJi/GKn15SIVFh+dHK0HCh+JS0PiGJ/YKsBszn70zrQGGnx7Mq9ApbBOyNHzsgH9Y1Tjo3xwH
qToTZHLiO4QwiJoYD+efu0Hzp3lLbRnt+lO3yU0qccCbe9ma8HotQtjPU7jk20G11FCZgoMNnC1G
W3MIjuBDDxhvjgs6pdyHn/rf91bsVz5oCcvn+8raYW9KLFo6+89UH9siM09GMXAwOPmIlFERQTfP
ZS2a7yF4z6X7hyObvZJbsZnBIkaCk2cQVlJdAFo8knG8uNwg3xAjpgfWjLtUUvssUqoEZ213Xr9v
MIQJySMfiEcVR+lA7m35IjTHnHb/TCvQ7i9VBwKtNNPPeAcMnVVxp0prNFXRHivx/bgvP3ldqFHn
GfUwWxw+OskR6WDIClMGJWysp86Ctk8ywmz61n6nfFPmpyYQF4iPb+Q6jAtg0NLaEwj2NiQ1cU9u
VINKPVa9VuekjyfS47NzrMEbaeuns9Inu1CtrB/WPV35hoi+5pr3X/W/S9qjN+Caa9qHM/05Idtx
EhG32kRina3WAe+k7YirJKPnHvYBcokVs6PBSBppCYPZXsMmsXtW1MojltIFTabEywKlRX7E/dJD
pHgxUy93UhKqnGG+QBNTxMv9W/yRb7SKUQ8UEZMd+1gWRbHhsGxPTxD4pzEeOniPlxncqrEbiZbk
dhTDEjb5uxhxrD8hU8Aex8W5PAoxUboREscwjY4ngfapKvPPzV4NaecXTWXeGU6fJLIEiejtYmeP
QmyipSC2jKNbg9J/gOEBvFa/lo0ojtr6W5Spj/Q12jw+TqMo2wcZIhLYZxZj7qZjUXWxLagtECHF
APErGIvUftRmFFUQsOoTX6OZLGX9zqGFsNatA2RwyWL/EArxx133oYMbsdeMHqwfLSUDKYIIXjD2
tLP5FhZ04Ulv5Yrd1Kp/VJTEyYpSuySBH8Oyi7gOi1kDcqjkyhyNHyrQ0ZpoOhVMCwL9h/e8AmbW
zk/iMyaoQvje7LFN3c72BvduS63HU91jNl/4JXnAeVHIj4VRwo3dEfi1x8muyG3rBPgyNpfOScdX
4T2+r2AVd/kAKPAXajIo3WU1Ax8yM/a7glnCoEZA3o03p3MOntBHVM0dCa8tVTMblrCj5hLBJDif
+H0oFfytGm+z9sPrIe75Ody2aDYmDHs/KcR8okQG6ChyKUlF8Ssi2sAdba/2BUWtQBILVQa2fr4a
P4Byy6j0CGLps6qEWiKOquMrIwD4+/4wd+6aJE4KwH7KDPbYLiFau+K1c9zP4laVyEXR2OMakSnZ
2hD0rG19lRJKFowoqO44FxJcAtG19XrvJ+k1P1RqADLkyGzFjTa4rMaFzgzxxuifMMoq4EZcfZU+
R1nkSUj1Vr2N2trXP4Q5Cz+XdSIBr1V9A6Qk3thvwUMVrAWyT9JHcPLWSRwrK0zNGFi8WepqUI4m
tJJ19V0G9oPgpeTyFTljGK1GKchlLLSaQC9bDPdEbAyIevbd760/RLgIeP29O8TT8E48RS9skyQU
0/PGMnhk9LXhEITKIfPjrMCFFBKshnlD7b3M3FfIDsluycNZidz6Ycds3Y0HIemBs8+kbqTLm9+t
ezj+lxzJjAdTIl2m1XJefkJKBj6we6VhF/ltqNymxJ8Sjap5kSboPkbG2H7GbcpvqxXgv6tafyis
0mBCXlRJsb5uxOdn5JfxCSYcXx6eMA+R12vcQsoud+CmjW7XE1wUDWAPwwDJP8IbJztgAi8SiJnt
rlIEub+1zaW/2a+Qe0lhHp0fMl/2mK0LZLJnAoQn2vM850tw3aPJAwFjSfGANKQlskRKFNfI45xy
qMwpi0BfuzIZXVntKwGa3ewrc1n0mBUAI5kUX04cZtdBwujNG6F8sZFvEzt1bdAypdnvlUYaqHXw
97NZLa5SXuLkgAzKNLSM3VKtVXTmBVfACID2uVq9S2FKCwxJYc14NSFVOb/JgSKPL2QDUIK1Cafo
qyO13vpt7Upmmc29vfXCtCz1dyOVas+s0IDA9oRbnUwTTfmQuapaQmpOOL5DJt6QuSBpxPhonlai
Ik30am4FcuLQ+fmZ78ePBj5/x4T9aaDujvqtYyWzq5l+WOMgG4XdO0uXKhdLPFs9fweejgSToZpa
ijeUQW0Ziwrlkm5OutUhnaMQperbC6q+YOBS9sge7ImuNsWYg2/+fKM9s5seH42JcKwb9Ojo+aCy
EpiTjoX4TdCFrO9UxUkBWg/JQND1ZOFdibshbYymKLpHJb4+7JpLDPE1tjBIvVWz0z8pSdRu1Qa0
DpYuTaAvfw9H1+P0aWrlKpDSwdANjoEbHYFHwsIDNgtzMBJnSV3PQc/GEJP0j0hxJbskp096oSj/
suvkZ8kfprthUz0zdbKzKq/JSfocVmV9qygKhEX2EwlzdiG4c58i4ciFdrycSiiqvuz4/XRRvuRf
09NYMRZO8jTOqa+oAZyXEth1M7TWX8cakhSzHMdu7LDP5969V7zIrrorOkWny9FblU8tLNTVyND3
G0u0KTx8hhw8iBALXwKSLa1hzXfBaQpu7hQ+6nBv5XBJsP/KYNbA3ikhvWPXAxjnGBZC7vwUG/3+
yu3Dhax8SIzil32K9+g4NgLqAY8djUv/Nv4X7rgDCaZ5HIpVXkXjTWy3Z5kGMnFHYFWDr5sxOe9z
aoArcI8bBfxCiXr49nicD5nj1YYYqsdFKrW/S8CLchSzcq69FLNbt9iHaqJFXoA9xG9DyLxkgSmX
QCvUQ3FsMdNqXo4n3xOp2sHW8kY1YPMfodF23k22RPxJtVP0qgVEALoA667Z+M6CJDbhA9CfIhW4
V5AP+fEiH6MsFqvMExVRpWzLJ36VIrLxHLudOMdsQUu8Lxz/8YZWggdAjEqvAFMKkKQZ9u40kOjX
kcRK0mVQXb2UyH71IcZtlgHIyWz0Fzdk+NNoSKCgaviyg0aXWtfg0LiPYldzbvrtiGi1xOMaL1pX
YoqNd1esH0mz+4YpqHswGZdebI6w2omf4i7lIEU3LEY9L8LlyzadQC3sz+FjW2q8yQUceo7pfTYO
9dOxs6cqAJZZRXo3FCX0aWAEZMgt4VnJBF2ATr70uc0uNgVsUTWsETBejyjaIBoTEinAnlDa3rXR
ypKaw4w0WLAsZE1Wy2LcmCoSpCP+5V8khVIGyxKA1ybPZupBTFZ7xI1+oOZlP232oaEVID0Fpf3l
UOnVilD1PuuRi3iNJj1Ra4YdY8M3nc5JJwpNsFR4YYFggXmn83GSSzuySoC00V+xpkC5UwTwX8pr
7jIvzAIztV0gsXDc0URWMYAaSYGE5x5rHDCMMKFGx2XdzOpVFajp15A7r5YsMb7wFi8ZL/BWvVbK
fPbV+VgUdamJSVUI5+jTdFstsbj3HjNZt7vWUAjAWLNtSFK4tLr8Gh98ao6w+rP2Ml0p9epWDfZt
eSaBz9RBUtSXsNQOezC6RTLNrwTXH48AQp3AKRTRjhfPWjGMmlCWypszZK9fiyhbTTjisCi1S6H0
oG2QgBdGGP3tPzEv4TPEGga3Fidnwq0f/MLklQg9GbxtTBE2W3yQoCkRH3rjSQzFmK2M28awnt2D
BArTEFc4xACpZhaJrWcG34qgrzwPQK0Psa7PnTU/1LogSGQ4SkaqWMHcaUVlKPGk0kWpWUQVuwKm
g4RYvhx7aWD85ZtqTxRVwCQwWUw/0Qinq+mhwkuOb3ngaFVpF7dbgAFSBilGPq3AhDaFs+M0ktnV
5OSB8VH64QJRCwtNNMXzFNEr6GeMyJ1eJvcb4OEV0n86Inwmy38gLNwT+xT4LLpenlm0Vg7KtVB6
ROBJfU74/y8kj0ffT2hh/wQb4IkDED332g2Xe4wVR6JuAbouK7HF7nSR1aiOCP9DP5YD0v1Vq0sf
wOm8SJxvUh8q4IIIfZFKkjR81QwkKRDxrqGwkX+J0oRonMjyhpFRu+3FtFWyf/Wh5Fzv05ru/lVZ
NWtVc6vnlaA6RQaOxs68wnt4oLqGG6JS0Fsm2s5H33UP9qnIj3vrxV5t2V3rSaPoiTq7vILel0nx
x2M/OeQ/Kwke3Qf9cDVN2rElhwYF7FiF0AuORnIcrofsajdvXr04pSlZpU0wRqoGOykCgP6jJ2S0
4czUgv3nA/avOwW5lzmSjhlp3LJ8vbvPe7fD0diQo/2+g16DsS6O1aR6hjZ+wiizZCiXgKYGXLwe
2hHs3aa/7bEWZyWCQwG9bINtVi9DVOwGf9bDxsEFsZ9I4LLynKXVE/lGkMAbTx1nQ9jvMba0ZF4R
uoNlgWHR++zl4Bowtki5eumkWo41jT3b4KO09EPmFx5UMjZmb6J+3bwmOSbt1viSKhmWRxKPQDiS
f7QBhbrYhMyZt3jr9jmHWeHaxOCaqCQdi1g55/wNhz+c2y4U0H5u7lePIitRFqByQgWEc1yG+H+i
8dMa/9a0tefb/poEjGujMcL+vHwm97krTH7iJ9UEsEZLm3gQ39b1hUH7OBgwxPxSOPWmAdq09w9c
B2Hu3rGEr/mcYalcGNZS58OltVM+9BLCJPv+brcTFO0E7kvHBYzSHP6+CajM2BJ5iIiov5l2t/b7
4cJWKNBjZm+Awc5seR4VDKOq+76rxI4F4afxcC9Z8wI9vQ6bxf4TYk8etqsR741u96W5BO9RKPsE
T90c7P6v0uEKa8RZnwOHNFXeGfdeSbLwWNy0gOU+OzLBX5tGFX2Es3SuMypWH85SYawdeSapEfnc
ctIHNKISC+RkRFUt7W3C2EubhCoKBD6D7S6JWQK/tVTrdpZzkAZ4UYY7oBSYfY5yO67kVkGR9F8K
PpTZvz+62kpNl4It40xhFez1zwoVvNZJvcvg2tLI4OTxi/xva5PHxfo8SMVwicbd+APQNDeCfUaS
H/OR/PdzWBYk/fqYM8gJ2OQs1lNu5absv9O/u3GmuAVqWSSPNwO+mkuzpuAQ7yHNmxqxQwv13Ke9
aNfnFjtii2wGcT088OhYvXGTm4/bRH7J3nNnlknPwXfuyJDTmrJ23QaK9SgVBoKoTxtjelmD3jPr
yX4NaPJi2sja84yKxYg1Hfw0FboO90oBRSaA/5mQkYz+G0nmf2cBj43nMck17uMETaCfUofyM6h5
KLis0XPHIA7oRNv66RfoFfpn1hAcAu/vnHZCALsz5jTqR/S76uAhxQDAsVwUDApiQTj50Sin7y0E
iikB/rE7PsaclMe2litM2YcOnyDvNxR26jlmX5vxbDxuzqOpAdnke3bj3Y1wgyQIAFf2CBYbI5MK
mGozgMfa96fzQaY1caE/6wL1uNGEJdVNmdAYXMT9tVhMAXhMT7waM3vW4CzKE5dm1Q6vP2YiuS01
p377Aw0mSa44QJPJh0JSIgdFkOROEhI4xwf8fUddNLAjILZ9HPSeUgEMuAXkp89J/bfjIef//b+z
zjWpTWGHc4kgTNY2Cq3nZfrzDoXdk6CiXV4OtdC5UJCYEftVUXSu9vJ+3zuIlncQBnS4Qotuy0JO
TAMDYp4pUKkAkj5a3o4HkVNjePeRSQ0drC+wA4XU+msuzc8srnKXt4/cNazrRIrjE5caS6C/yXCV
psxhKZ3dgwOAHMZ8qGPJfHwrNduND6nc9hWhwmlGdPcT9fliVQzRWBUyThWTyFz4n15ibLhrEkGj
eOUnrDu8JuYDPAlVK7Vfj57uQBXzGYBgs9ol0Es5NKGf0wL1PiTkGJWayylvLOLjKjKC4xZ93Rnf
K0xPAhz9XnYyxq3ImPF8q+yVQPLuEC2jE8Hl0MDPit+u/0S6OqebcefRi3vkouLhSQ5CvNbF4kyl
GKURBmzxcRciE2lIqRDrjXhreYg24G1wQLS3HgYY64MiAGmjIzNH32FHIImrCfJPkpZycW2oxSvA
NRYAQQp5mBGdkI6vq34Mp6/WYgcmD3xnAdVkozcztVO1lK6+dVl62E+GoQyzvm/2XYkLqRGhvsul
DkIQA+4hyJs+Sdn1sPcxjbB4JcRp+2k78qqOGUmq9GlBs/WPz3oRX0B80CfMqoYECZ8JXF+2tuD8
uvynLMW1sPvVRN9lE7uxEEGlH8dRUo0bMIuOK7bntgmXAiwEfz9o7ddq0155Qi6hUYADZ9sBQ94R
usGYFKQUS5WJyGF9xebJRIWl7V1fO3HkqygsHpkNfdlmRfLHDncDH3N8Cbdpeu9PVAzofGRaxvX0
zBmiI/J2drvjWYEAnvCWtpowrjwXnUI1DBf/w6TfnYppYasAP9aKJ1byeA28babpiBkGBZD6BF1a
9oi5aZrM3dbdjACXAZ4AYjaasRnWEkcQECpPODiF9d1kpzZ6tLRIRPLVFPXcd32MMB7wvxF0Vdpp
TqDYxh8f9xxUABAOZnmMWg7H2eADnYM6ac8aCLIbPM0v+kfHz4Ea4aooDGTnhcAPCJ1p6LjmZ52w
V5p3oKP1fi+S4we6tCZxs/QS3FzBp7iSo8KEEmRcOJ6VY1q8gEbNQToJDI7vT4gwzlmkhxQhQ+QL
vJFmSCKMnnzzIzqtcvijdAHx4MvVB0TiH1velF7bAIfuUKGYkBF0jOTikxRmJRY0pSNF970p2HHW
aWwrgTcYVjRN0n1UtMDrCPmW7MuqHkXE8cdKv0lwK4+tmz8VIZKcUXk/UKx2MCgANZ+J53XmTvgZ
pyZzVzcrDJKgP4tzLh8wNwzpRiN+sjOjpJFjKKizTSxKW5V71rhIR8DE53RBI8mpE1h9lXdFguDE
C+nRLZvnwUnBKrrCJkfqHHAJheGb9CL28BeeT+ZOMaHMEtNOXDf+v2Gd7u8o0gDEI4Z08EWqe3Sn
TSivlvpn1368BQ1xdddTlHUa5y46EA0LjldAxQUAJk1N2kspVFNGGnHcOgeBGGK6n7aFK4O+EQzw
QFUlx78QnC8OANF5ZDjHDV+j8NeQWruqzodvqCxyF0YW2xFUVecAjpHYBbeehl7fyHVx+3xvrLgf
0ZE3J/abHrKLBQV89v/JR0/S4dKNAhGZHgxCNDJJ651WKDcrb/6JjmPqH8YIA18WTT7QBts/4UZj
A4vxaIDFSTRHrF3YamJ3i1GW0NagT3NaLeOcWTGfb08YDE39ehGeHTh6p4zL5N55xoOwyHSzs/Bs
3xsSKJt8FnL84IGRCr4cHltFs8s8GRTj2eoJSklkw3GURW4k+0MuH9mWDrd7vsvsOMXVGrDx8rxA
BKqWDThx120GfMYcb+wtGIhDwFFy9ZLb7TkrSC9WxNrAxukZqPRTvI+Bt5yqJvsqpYCZ2U8r45nP
QhEcHUpywDDavQ8/pPp8aVSk2+8/8LhfRGHnsT+EAGU8BcBEUgrOLa/bRQcdr2ks/m4kCl8Ht72y
GCt82Aw6dunLQkWu+Fmkm2ohJU5PdlbwH12lNaXw375Nshdj4VFhv0BLDRkgLso9CN5OSFL+49Xb
8ksIS9u++2URzzgXw5aoz01fp+DNtldetDhCXB12nu5Nw8KkjJma/LBls0+kwD+kBlS0ehyrtL8M
keY1BQP83oa0GyZs6jCDa5fjwSRBOamvPPjY5RAp8myqw4tEkRLsDzdFjwEXLVZwWk/IuyLBo3Cd
8OWgjT3qwp9uLwDBmBG+JJc4n0YYQzglfyWbX/kCPLqsHEN6TMCOiqZ3JsuKBVp6ivzYBXWiLeTg
WqH1wTbG3yAi1Y/Vt9z259QT/Tdg8nbGlx8Gx7IGF3TNljYSS3H2ryDvdqHlkXUWnTv5nGNHUD1u
lNln6/War+aze+bngpjvecDcXT4Y6qTDtTX8fzcnTMlgrY16Xj+6zwx+UI2PRAfiC5D3ZIkLCsUW
jx0nAMPHtbedwWuT3v2L+zjUV046k7qc95XPxbWq4chJyq20NGkncAjdxXFzrrBu2aqJKLdyE0RQ
UKYtW0sRWok485ZwdDRE3OcoQnMg3bV/S0mbgCNvbSg1VRYbTd/ZOVJATmO841iO8gzK2Bv0/rLg
/wVjBBPHXnwcL8Kr7I6YmyxwIBaM/0UAVgWCbX5bytggQ7ZzvSW9AqUpEW47kyxMhRhZ3dpLUj4w
nIbnbQpxAn2VIYVki2kk4aaDsXp+o6AmZRu1H2c69unkbWRJF+62D2yquBagQhvih9QBjil4kNY2
WlmIg1Do4HW4iZJMSRAKY4RaREzIDA+/f9773FPuJYIGJqTP4XWI2AHSeQRhjzWp/+KCejlAl9Yp
fDxLboAIbp6JnALWH7ojuqF+ri1klYSm6OARXuv1UtClGjF7PPmFhDOEfF6lYI+MpQDKhrnvHEHR
BnfP/bLVvZAvmasLl1ZNIxgTaLaWGiCcA722YhYzCtmQ5XYa5rrbPupCGN7yyIFImJLk56EgmMes
3TbcGgVK9t7woVRHg3omUGI6PxRBdkE7ez338KBihymXiqaTOTgPe/iqK0A2f/qp0NwJePrcx9RF
ZInF3Bu/T2JyMVm5tquyE7n/3o0PiKh3f8yUwUwnnLRUCfLg580dsgYUkfCUMUNnA5NQEx6rU0Kw
HAugI9p3/CcVMBIRcKBurPsnaTGOCn8Duq/N+Nh8oD+eDeI44yKQnyhBoLoZgDD+1boms1evc86n
MkyXt6laRLHt8Q4t9ESyD0w8NirI5iz9HhY1f48obxUs9KV/Z/5mSWbw20NVehumc5wPGaSfXL3B
VC8PDrFnWUG9WRTgSlN07mU47AtUJkPJD9Ku9JzW7fMQp5jhRe7Nd3Kdz8lVgWamBU9Ya5fxxGwG
aG6U7luzv4xWUkgkz5ADL3lvO+4Y62A03EhfOHXzmnsWNkm0/LzjVyXEeQlqe14oTs92TqjZaUiK
qTHM4kt4h1E7/tDXoa3dfxRXMmKoaIvs84xBs7KGxoVLcJMGkx8F0zO3WBRdSb5q68bpA1bg2w1a
2isshCrTaQWtzTa2PfwqYOX0uZlNmEAf5Xl1ymmS10i7wdJ7hn2KMx4eszAJEaahHEP/Va419vDs
wgZQipwASW2HP6D/UKa1Xsh63aoEqOlH0EdyXEifLgCIZ0s2a3JWW2TEjsVj/09L5MRYFreZKLVe
u1ZcS2sY3h8WODx+rnnZ6QnB4CWLOx2Kq3bC1bzZwLbDJqCZwCn5EPK1v65iDytjQ/B9GSeBDG3e
i6NXaMYh/RZuE/i5jrgvWJ2mkE6WgxY7EjitFTksLs2noQZzgyHSzceZcWwHYvGAF4Lo2JVWOwBJ
yDN1bVkYq3R9P6rzr7fOLNXkvQKjoIAVmxtzn3ruT8LFJ3ltobJQ26ZUBWV01swMG8+xLbh5aO4T
F+2VnZGjdFbJL6HHUc2TvbCB003OpvmELO2jf4sTEaie5cU+1OcIOobf8jKKWQ+rM/jpb0/EWVg0
tbvhtEi+eUXyJW8FyOmKJhh5ooxdT0QRV+Dnzq+JT2DLaX0i2AqZdZ/aCdgMJdVkoc/1lxSUOz1Y
ggSZJIDwDqiX4G7AkEhv4JUjeRlWP84OqZeG21h4MTjI7SZtnfPV3LNsfa6Lzzbe7ib2bbUxSFj8
LBjhZHAqNymII31UCGR8ixYI++yEXwrIDj0xCOJrVl9q8E53iQlwet5qOLPUlqUtf/SBLAR2PjrW
b3hxFN0oZCxd27rAMuKNMlipVX3jEp66L7Xr19RLuMuhIibSBkefJYV1V+YqImndl824OECOTzII
p/fGYdgCPWdBm28a7KronMHcaQeaUU9TU7XuoTqSlxYZH5z0cS795MhpVVjAsTRhiTEJWDQYlP9n
/3Inuez9d25GJ4ZTaHhk9nIKHHIak4spgtBWgbcZWZDAsvzAQO5Vzou3Xsp/CmiJn32y7rBcY0na
cJDFSU9mycxBheCh83eBDRQpw+xQbteQnfkyg6vyHTIaAE52TIf8Zm3JSYl1ljlUCwZzFbD2VxNQ
i6hYbioiD1USpRhXJ+w4LyQirLh3nXlX9m9hfiZ1KVVWd/rfkIkMkCZvnO2f7Kuhs6yDkybwKzc7
TQOwLrKSWQSquYA5U0M+RD51neuPcLpudVBKOQ3QIe0O74sqwdN8IHEswBfjfmxBxxtzM6WAh7de
AKqIYG6YZCCu9l0d79Azj2VU6idinkioZxTRwiauqrHiEOrmVi9Pen+OpIxFN/6/Maj9wjZP6pXo
s7KYJl6X99nWfPtFhv8oCBv3ms1CrBEF6juvfvZO8uJ8m/QKdTSIaPXmaNpGLv8n4IiHBzN2kGyD
bQ2uBlizUhuGH1ZLOITeXC97gxC37fEt5qJKd+O4sHa7BPzHLke/xwFMJrXH+r9K5r5kBI1PyeV6
lKWjrbS923/kPPaJeat+8O0/wr+ARY6v7R2q4rqYie8I08jG1QQLmrvw/A/Jb4zqRaZs2oV7ysmY
1dWqX/Ebhizz37wtrUwcyCpM6ModBH25KxPE3JlL42cQcRC/ij0xTCcJSgpyub+DDXl0/d7CdNsU
VDMgy93lVtxH5Q5bxMZ3qQPItXGVdxgnFLWjtfMUqwvI/IQ+myvA+mXO4rS7P8IwqKKcQ4VVq+yV
CmsH2zFrahKSeOJYGWFbje0WIh9ZozYJU7wyf+Cybx61nhufaSLEMyL/kOxVUPjDuSZEftR790Ti
PeqinS/9q5aRrTUO+xxvFEegHbGFH99rrCOtOupQxZIcwby5iTi0+X4sLg7DUKsRFGvr87mJpZOJ
WDvfuZMcs5tWMTvi2PPVunHpOHUdBUNLy7MALkBMQgHHNo/N3BlOD/YshrdvueSx5SCwTQKf8nTG
5hfnz0VPPcIpOTJXmyJh5W9O+hFnv5QhQ+h9bUm6rmuMfFMjWUxFT5SQogoASTNBpmGoBgtpuna+
+sQ6sW9wf0NZoB4acN8nOOBYCCg+Q3jQOaEK+fFM41LKHoU12wU2Vu5YbdLpZvhzVcVJt5mRPxLy
3bh4IqD1pU6VILNqDy6PH2uqou+tub4q8QRjKdeTfFMNSTu+u0MgGjZCVyEAjc5ZxdJOcXS18GjM
4DmaTqoiqVJC3uIqqfaih8yn3b3RjG7xKc+3PjPmafsk2PwwSqm2vGbRlMSHbmJueM3K4jVeaLA9
aFDWhPkC9jMhGakUjdA41paMUsczsIWNkG4BTmR2Vc28DAOrLqgrknTDTNGrRVoB8wggfoTji1eY
1bpwZtvOQjyVpuGoOfr7hiSroUCTYHsav2HWJqdSDnqu8eYGLkgEwph8kTDQwosdslqL1ijiu53h
WDZYPY6XwfvINJ+D/6ETQHnetI5iO8tu9h2RbHUcALeIbaVU1GwK4v7RbWtKkWes+zKdpuO425gL
FliYfrf5h0zN9+S18LOdRxWYIyjj1jThIwR4Mh4dlXa6KjvLP0EXmsi/XTcHaI/1O2WJKhX/hsLM
C/WNvHEGyeSY+uRoowCA8MEOyhSxNSvkOIhcSiK9d5hny8yN6EQsIcKK+KqC39p3EXj713Q2uaNf
TT8F+haSQEtMVZJhv5OxggTMrImd2gtQlcM025xHMoqG4Zi3CoybZhNyUZsErE3LPofatQ1JbTJ4
syd1LIgZY8+iUZzs8OHGKExh3JTVbO4k4iEpFIDE2g0ZtGIHlczpaXga6Vkh+tZvSCog/6rH6r8T
cABDc9fHJwwTsE0nqf34MPsNX79TqBaEmRlrSauQRS19g0eN35d30udgKvjJjthC0ZDAlEQwINOb
5ymC3vDEFkLOYkxca4QoMFw/4eZSixV03RrtiFr046SQuv/Iv0FRr2MCigEDQd9MR3FUcz+8QMPp
DXrhJcdezxafK+lXmdmFp2swW9+CRMXVI+HDbuMdbxAVSfaBTddbaPTdcFmyrDNi7wA6O5bdRQg8
BuvDlQE/JV6/xLc6kMcviqawAXd/Q3x++o9zroAzBDrj5If9w+EMS9QNc1FaDlqAM8OgyrPtjr6r
PMJlIg9si9ORs2smOd9O4/uqF2VtO7PCY7H2FphjIYDjkvUswpU00BRbdHBv049RDRfQXZG2LPWD
Db2Ywrw2CFUmjKLL5mVNGSoJvennzA41k4HIFUBTdHOJERWnT7Mv3qegZgBh0sw1kYXcXd/sPYYd
fJ6ynQ2OAQOGW81YLyWKqPfUsxt9tHilm7LWA2Nrdlx7/3sPebgr+4XuQlCntcekZLhZYLRCg9MZ
eko/53EURb3CJ8dWI7rr0fB8hIYtPq+u7ZZndni1DxkCkhZ6YH9h3HNRVCPLGh7XTn0UQ7Dr0Prm
KkWM/lUCeAzAU+pGvtfp/bRu6b3b6TRlcjVvDKtqufDIWtck9X67ArEKj0L4PUea1WpNvROLGp8g
b/PZkv0jC0K9QUEyEwMjM+Ka0sKH2bu7qZqffLsxsmrHC4Q0PYpN3GVBLS9O10ezQqliU4yfC8rb
0asesGjy0lVcg0ZLISSbHV7j44TPFeYx1ukNq5o+fpUAPw0zi5qygU1R7ijL704J/4XtOcmdZIMK
bEXd8i6rGFFhx000PSmhfL+Ht/CyggMalsfooDGJe+jjDRkLqJVi0V99ZvmtHZc2yjPh1AeaAJma
v0AghJrt6FTP3aIHMMDK47wSIcxMPwMNq+jOB6tvgfJbLwc7hwaERTXO/ocG62Qssjiu++Fj3Upj
SD11AQpmA5wGILz1he9EXZPrbv+ERaGxgV1cOwPbYnrR7JQalHruCKHN60ns7X/GzpuCs5nG0C78
UUMhF2uf4qU5tGqsw45jRKxbo+yaR1KnJ9SvKws/dkRKv/lOoAxAGErq56LrZx/ATMVUFJkyn+oZ
end9G/qDcg2OY9stbkc0lsV1ZqAIYukFI3M6UpRAH7lXHrm4SuQ4NKTlClAQE6ShUUWujulNjFN+
2Y/7GLebZkgi+bOvx2X7cvXSQIBm27IZd0kD5vcCouI/nIoz6Q1gLq0ybRYNPrSeWbUjf4gJwlTS
cZYh5o3/DcwZHUo6zpbpN8Tli+qu6wu3j16C7UP8t8+4lS9kPY844cCj8UC7uli+xYkpCvFJVRo2
gtVrhz1texzckacJTwc3mjGcmVunqGVWNArr8TjgqIjkMptTbV/YG/sbkI9YA//23Zhm81NpL9/i
jlfcYOMd8gOlXnteXld3EMo+Xz0BLP9mPfO12NXMeVuzO/vLYuMN9qbPRnggtm6Li+61n8jO9piw
BGY8/WVS3j2RQu39CrN4vzGeyGrm59BDZjX+8JO59wRsVAJMZk3+QQtDp/oPGtcqDgQqbKwj7UKj
VapoQPQJpyDWfLYNwg8jfrzp0lNugnzRkmLpfWw3Xhuo6zxdYMidHHmGcCO1MoYQFM0nj3fdHvqm
jb94xCn8CSq7cgmH0MR4tdf1QXyewgk8gKtD/bulOrh9PlxSRkB+TaW7tGVHlMH843piW9pB9BlW
GPqjt1Si/gm4l+C+YR49oosfq9ZUYmQsPmlGKbXqZyVXzkhRNFZWA5+OnDGKlLXfRqZijsSHih+d
66nEnLRpzgteUI5GE0hrsY/G33nwbCbdih1UmPtQXfn2SgWVc0kt1YdXIBwEHkKsVVtqWH0Z9/iD
1iWkOBrjYb6XljhYXJ68JzVZfEdby01rxBK/gbFuTYWZ6dxCJDXySfhcUDxrDdVlc5t0qr284Aig
Fr6GjEp7EeRkcECPW3i9tsCRhan0ZSdpKDCieRrxHpj1zqL3gXPUnVpH0W2HTgR8MYlN3M9khg0M
YRYhkhFOgetavHMl6OzUPqXnfxZ7KGfIK/Gm+EZlxyzxMmGBqGttL3U1/r10SJGgiE7CXPIDo27y
tHz+iqPwrRI7opY3h03QdzdriGTWjCstBXgeHjx70i6ja3v3oNUtnABV9+sy+qqXDjAS74J43iRK
IhroHnsj6T+GMhprEAhKVT4r6ZW75IZxq6KG+YUrN+3+w63mv4NdlE6PRoS+4EsfmMQq4XzchOFt
JcTmb9xxPniM4EiweDVPxTGAaSvgSqgdKtKD0oss4PqmvhMWOo/SRoiWnNuxg3A66t1Nv2zrMszd
lytPIjsEAu5wcW0i7qXzqf98sJmP24aKgFu55AgOD21CfrhOw0k75AGLhL/mm54255xcqV1jYNSc
+iBmJe+IfMqGcEhaFfRFX9Sj21o4bCHdYEVVPC1+NG0yz6yw7rIV095ekX4/2NJqtfiV4wMG/zax
aYuPg6knjCY7kM38SEXRaOTrQFO76kUHgRqlk9euDBZePdfMDXi7fQpgEBjYKkokMrCu8yO0Ji7f
s1J1fPy5ajqe/O9tM9vo0oqMk7DJdFDtgoK5K3/FNJO4aRe0ZBSlmLeydUEOdMaKmsuBLRfWrtoO
w60/vJpC9YwZmg5E12Au6+we8zX5IK9bStNeEmu/057icgYexHQosblw0zTb3s2KrTK+WLLwdU5V
JjJrYzz4cGr5D7wXIi57BO334ViXOGukIHbrfZxqFL+tb7yjoLK0pYjQQQt0ZIC9QSZOcAjwvMuf
s9Tj8c2I08MMvjVuPqLfwpqhVtFY5BXmEXpynVtvpD52gSUxKPnarjDA+SifY7z9qnMG2/dCW9pW
87ryr8DEfo/HUNXfL1ji+CrIr74mN7AZLG8VBE65VJ9tx4q384DLVwyS1qhjid1iBZqLlBamSIEV
v9Gj42/EVdeaOC2cRPD+sF18PVW9DyMyjeogfPzoUCUulQgFz6+AqucEnoTHIBs32ocoRJXUlLjk
8ambcgN3CH5TAD1WDIlJoFOaX0yJvp3hqbKIQ7rKnUveYCp3lo4ijg1iJoP/fs47f/7JXO8qhFiw
VIIFpWIq3djViny0O6ZYeh+m77DCqlMXxizuFWSxe0vOkX/t4EdRlsOxAOBfcPX+AjBv7wAOBJe9
jm7dKk2MBUuQSCVyh7ZOwF+ZK4TVxXiwT7pAmY2ll5wyWCi5omkvvbM43bJzh6o4N2eQDEQnm7H7
2MBNlNKiroT1Mnms2r1HDcK2jj593zpgfiAV5kVNMj2oogDymU4tYf0Hj5jnzaUXFoud9+Tl3VcZ
RmdzNnjPqAmdKkaW22FrSQmml1ULVVDPM0IusF2Pl8W1kSuM5VTGtagcbcszuUDPEhEqtdnn1fUI
6xwGXfG1Z+KWWV+nJDn1EZaVk6P1KcLQlP/LqiZ5fQCApAOuQt0IoGQ3PODcKCuXtiulaTazdVSJ
c+YhGzlbh8ye0wnigNUlSrMs88WCq2USBh/Yv9vdPDnN8XChks11imujgdUHZ7JRUYa7ahF1jz3E
ZCrgJfrFK6WLw2PdDVQbGp2aGLRAcrVs0vRnrJobGFkW9DVm863oguVkTtPG5MR/pgVo9CzKv4zL
ckJjeN5R1C29nOvRXUTDtpqKyo/7jgP+kRk84L0KoTLTFrOmFWmO2iH4P5B1oifFbuEHntWU2Fx8
ic6Ukis5+6dmrKHubAVuN8/GUiWvkh2BuIbaAn+vYE3/uDkv2YJQTb2JOwsIeNEI52P608jT61fJ
C6NHBMyQgHG9JrEcnILPTh5O4wXPwQqGiqj7dsAXLVkYTD8uAl5dSPXzU6pYWJv3PkLKTS3ISSYC
bpk2P/HcPbFh8a1Hhr4q/QVEWrnws7H1ijjYL0C3ynb/Abj5zVKeojrhLBZh4J+qMbrCgHu6LdDt
JbQpocuR7irCQumyxzzQpIdFUn4lRawABh/1Tq2tzf3FEcAK5vcNBVlOPiwfbBr2X3iQyfyX/kh5
PJrBjcFEzOwLKQ9+bSVQt+ZhUG+S9d0DOG540QlI29yo8wtVAvuz7aEWvrCaXdfichdaRUG2WDZ+
jYn9uhiGCloVsJpCNGaNCzfLif1DETIFsQFPTV/TCTHFBm3Hav/oi/bmMIj2fJYYxonQQMb93u7l
MSshFkXogg12h7gZbbg5KFyX1sAI+TEv6JOtEAMWBpaf3isiQkAo23HSXpZGFsFDcvj9PHPu+CKK
GN930FnjV0RkRkF2sfVSOjXYwpt4+9bThmnlKRh3pvKpDcPGh6se0J+T2TgzUT/OJK7eU4qA/RgD
OY/vAf5lRmA7gmcSAALmUXJZ9vK5RwLKRif/ykxGsFRswa8ujVY8hkeREPmFlHnNGu1QKq7tqktN
U7t13H7aUyaW6VjTiBogiegh5IaYvxOIYkYpZH7Vy6xv1BN94n7rKHGZslI3mglHkAzDgdf8dV7B
ArpV85TH2V+7s1lRJvyFpRKoLSgT3wdHXmEK1s5it25p9UdO5MhZE4sjsmgpMZfTV5Iu1Ja+3B5S
8BkWMYFYQ04CGxKkbhGI3+N5C3MnNjWN4ASzNpSeKJlpVN5j8EtT5jCwexthdfRYIfVdwe1aus8B
WpU/D3wou52er5akO5n6dkOEny3uQqcskQJbbeHGHIJgMn47C2COVjlMiHmS0739QQmK7h0HtY7L
Kck9s1Za9pTFzJlxT2UrseRN758P1T1DfCh9RCUlZcw6CRpIbgMpm5LlEqGWqzqo4DY4EixZxW8P
Yt4DolW+ZXf3ozbGGaN0FKECc71O0B6bDXfWqQZEGZTqgRv4KXDkw5Yhv/yymrhol/CrWxGa0uPl
KPd/M8r9ZWN8JcokBUcSe3EZamDcl+jr9JDNlN3HGhvSaiM0bX9ZVbY1lxzAxujbJCG5OvYyjpkM
XoH7o8MRTSYfutmLWq0vhjF6DmX63u808VUXk+/2nTRGPd2Os3ss5yxa3aGv3N5Wi7E9sJgfTh3c
Pmqn93LXXNjfhtTU5Bgy1mhgeLbZriS1CvKsAi+yCf+J1uLvyGG62lBeBhsNwKreL4I3wWQ/UZpi
PPYqCdbmDljUysorXu2pC3yG+9vk8d8rydROurTPjfdtImwy6vp3U8z83y/iMcMqBzxJW9M+h7YP
LzmQtzYl9vjbcCgyArqkbpgV05cWIHSruFgskfrmSfeBZQfULlgP7Gm/O4/a3otnahIsbvE/aeQj
Gu7xPXkxV6fbQNOxcDiftlObb6xvLkGhrKHQaw8gfmHbtL7lDHGlZQSUU8E+0SRfwqHRQD+mrr5h
NjMIXtWNUj48CSrsUdho49rxfVAX5ik+VlYweyR5rK2mr7LbmrG3ihGzJC+Y1A2dMtNkg82n6DIM
DDEUmxi+Y6Gmp+gPXyOwLq6YgwUdwCfyGpG0WRAt6gojJPe7qfdSmESd7rUn3VnkRbc2ZhvNbLb3
+rmIpopkUF3qSvZzm1UtGQguQlDtlnLOyQZ8UfaBFf17QUKLh+3qDojgy4P2FOSdTGGQuwzRt5G9
URy/ClQTRnTuJmDNKklhU98CrkIHUuwfeQUCJ3f9ap8PeeLT2wUe2HfFWhV+UNIYG1HkBNlZiRbu
sYDst6uQzoh09bbMpbnk3Q8rUxgLTeV8MqFzDl1RSLPZPnfQn3+YwN1k3fziskvcuZpTTWJrbnVo
A+qzW9GS+AXHLHyL+dwT7v+t2lcGu2dyp5LDg800KNHwOoXxkzO5fqkz96lIDow7gTIWWT79QQM5
fJEHIu5AVNalVi5k6EUGuxV/gkFe5P5dAcRxCYkDZFH52FryLrdT9HySZXpqlvtTJYzfly7GcnzC
VTPBO3yH8abROJCCtQiV4deZGfZhFMBaaf990TEwMVnbeL1oJAU4+4ubwbHLSwaTi65lalA4AQBO
jJeKM0tApOz85Lv7FknoHe1NGqPbOxz4D6r3UGPtKchQett0D90I/ube5uhwEH1EM52ph+KkhVEt
EzXYAkfx+xJEzrwHOeERWbyaRWkLvLNJk2Dv+6mIpmg46XgW+ZiL1ZGacKLLbdMPRX1EvVz5gZqR
HHsUGyIGtykk+9gQGq7PzFJymY7UJEZ12AsZ3Ym9ZJzU3Vn1A3uh/Oc4r3J3/0jpBG9as5XdsdfI
yC0JTVstdmHYB4N3ipr3BzwgCQ+3vOUipfgtJehvYT/vyEoiYiT87r7LR6MZax/MkUMhfzoVTM3L
tHohU6hiLnJ2KfJM4m5Y3AKcosreqkG8yMvl0rydnM4XGafX4lutxLs3C0FUz3Tu6PFTvC6KIVO6
D0yW4r6HW7EEfAL6X61xOB3Z/+ZxiQKbJIXMLXKjLFgZFt83d3L4nFv7iWOvWbLJlreRou3gRYKW
sBBmJTO7DTdWoXbYVDzdRYKbSU3kX1ueAv8jF6tQi7o1RnExkyUCuv61ZNUbxEuT1RgwwHCIFZhy
eMMNCTqx/O3As+XP/+lhGZjxtK3iutMwWMEOiVGHEd3VmH57mhLeL+EK6mViXFwz3CftmItaoDK6
+ppo+hHz36c5wWkCDqwhWydwwkh3fLXpaOyHO5WMzmqDhNTW9QJcO1WOj0/NA4OwOGafG+GU6Umu
6XA3MnpCfkr/1v05RNo5HbZB2WCMovR53uJNtWVJS/ZKdSzhBaIat8zJObDhBVH6E6xIiliphRNr
7qaNsEsMQzGHVAqo3vCqmZ+eyg4qauuTV0CD4eioEA14yc2Lv7pcF/kAkETz+j0TwxTlsjnW+Nga
L4VS1IyNDp+neNBT4DyMfh4Xg9FodBzK5NxIudjRDKc+NF4SJV7V/D3P8BwotPPpZEmKwC0zKIYp
OUi7SfDfnkjwOLeXSphcskRWap2nZqYLtX3qNfv73udb//7MR397gNKugbk4P+EiFfcarrth3P3d
Stn4okZLIXne5nCO8im0uWBXgYtubeyCbJ3inNa/dymf8TtR3hf/yUGEvUmYq24K/YqbyRDH5Cu6
COzKfLQ020f9OM+/VoK8qW1x7n/mJQkV975ZBwvtOZGZVjwu5uqt9C4vYI3D0KWZG7l9DWxHjQH7
rthh9czeO4tA++6cik55eFnsbEN7hZLrvvqix8U+5BwFSBFpJs33ikOj6qVdj7pS1ukpVv2EK70z
lUx+1Ycd7mhwChMUwtXGTAo0DekACs1o3yWJvemdIKJvGDtDSMafVmlKGE504TxppCbQ3byEopJK
g8v7ttCrcQ8b4NH9Q1Fikh3ugd6sKVo6kGFzRVKgOzG+HtxMtnr2hidwdOwm3Q2YCFSbACDmo2xK
7nkPSsRzYHw1T7L1oixAvuOtLkXCsjCAcakyfNsih0AYDllcgTxjK3oRxM7JPtfVkzh8hpkbUQiY
qdlQ50eSgvPENwYO7r+xS4s0nr0KYnahm5WRPwOfCzRNfJjPFREa37i2c4Qi2IV6HYKHLQzYPKEM
yP2Hpe4LJ1PWXn81ojGGPDFo5UGUcTxhaA4iXMJM55ce7iQRuX0t8Tw9kngb7W1abQ6mlF8D4n3R
kDlTzzhsSYNdCPXmG7IjxN4pe9gWKFWxkWTZSsh6Gdh51hB+OqZ2tO0OLcHG0DV9doc/GJh28xPG
gNGF/+9i8Adw7OvS/XIU03PlWhBS0GvNX01xf/M5SqCgjsNYqAE1P2fuOduXBnyZLCJLeWhRpGVe
dD8L4xN82JdrRcUQHidg48okQcN6oK92CwH5LOZxh3QlPUopdO6st/reyvzTiTCPp0CXpyFp7N3j
CTTyoBkzEzvZHiZRmcXvpAnUlbGj0jDoS3CXNtZeorLxJJWvYqWBCoab9Y6xE4wUCntE14rWf2Y6
y7eDFO/ZiBk4ZmuRFMBYbc4LKmRNilzGlOmPJx6jP8VgG0uGUYaMdbAJAbeQ4zC/nD3BekwRL98o
RDhKn+P+BkIh8dVJ9iFbOZVg1P15wR616th2FXdEUaDZiPTNVFDp1QKjWOFai0XpRMfYvm306bT+
3Vm2z1kPHCfbSLYW7QSOW1cB6XXcayRa+lDbfnwc2ziWwR5aPwZnQx4TqdCxgq8fUTLR2ZEu6dps
eqWb2rO0J6vpcRwk/WngyT7HITouJ+49+0rpZdV8BEmQB6o50ok6LY2Y3Hpq0YQW98XKdmk45mdl
j/NYFh8zXEUtgxGYBHoFkXo+hj/OtEQAdbDmxW4hKEbLFf7mglPolhDlguIiryhLZkbEFHJzjzWF
utgUzOfDcDdJl54/tl4d581/Na2OihY+ASt2IonLXXaWjOD89k1KvTbZ5P7FC8AGbAh1dS6jLzIw
H1rhy98/kGNmXbh1ur8/Sxa1IYwVDl+NhW0/c+aan9E2ON/93V3A2bz4XidWoE+xeh+aba4n8y/z
IOEYtdW/TTLzQZrMZBTOeaxpEEwElTFUPFTW068J0qcYynragSkYEIQBbHNSjj7VajwtrV/968ww
4tfIzPcSam+7my5ID5Gk0zmpvWLtC9Jvgrb4zDbsiL7QJ5NpEuSJCO6PTxYnvUgtZImL33ru+0Kw
lXGxlSIJarSUxvQ5hXC980lRsJR0qxBn7qTDQeT3hvwJ60eWQVSp9EoEF+on0nwLvH6IFXmw2sG4
IOAwHR8V5bmu3fx3Xos3qj93Ib7Cd/YPXdPfy1pTWXJAV13DOFul8dHb3dEg0ugVMNzE5pVCY0/t
cya6wSNgKvmPWFtkWIphLN7RpJEG4RIVTwoU4KGtoD3Mqi9+mYTsy/XKUu0rNwdfP686P5AN1yMG
FswOP7NfHNoGq1BSitiBZwaZPtLUGCeLRbMPs5TQcbumTXcs/+QUdnheGO3KUWA/BL3+QIHDj5yi
SfoYy31idW7jbZqrT8avzGrd5WQZYFcyiBWunVdXhlOp519q/gj7dEWEXXkd6fy3eOBMuOObH21m
5AhZuJG41QIwc5QCy5eAGd29+CjCKNR+2DWl1/itQUl4T3N/YTGXrKPsL39AIxAa31ZgwSrd8yJ/
edz2qctNclJ6VyUG1bybMd9+QkeN/ADYEyN/nT6hyEx9mCJdzOh350CyuXP5NbuMCHazzTfSBTIR
+o1ANkLx2OcYLTi4/yA9AM0vkzSUDiWK0Phv4PPnh8z5clnViu4NUrviyOVep/I4sRJojuLalD+f
y0SaZN8UtXjaERgqeEY77xXMarWXV7bsWolFmy5yAKq/+l4e0EfIHwjSPUF9OvZ3yUjffhi+V5AO
1cSJ/NVdSYtgSt8UsNFJI4bYnQXa22VnOeLuASl2jPfp5YckNkfcXZ/OUukXxQzE+wRnUa47MnMj
6MznuYgFUlXyZDXCFURSQihLjkruY21cfvLN39ooL+P5I7qfuJO11OF0TL5hBsf12Pu+a7Ax/oWm
ftub6i/BsTc7aZcVTeJzi7qvf8+wMHFMMps9jPsmb2x/66ZK3wiJa4IRFVn1+A2QcQOh5RBJU3+M
7K8aduYX/wHHLV/ADeUTpkYLRpIpDs5YKyA+cdk+V+3O+0bFw4cVtTj6WAz+ba9oKmOAbQ67pVgX
nEo29FOvrCef/G6ZxkxcQgaXjnyYSZMBX3GjZQj0UgXl6rH4+MDn7fStBHlex2zJRqLW5NHLwYzR
lemWB7L5UKFW5KurRMzwlWnx6qv9mq3Y0O6OpYuLO8zC+SRfq1KNNgiAYgw7H7+qL3GF6iu1fFA7
akkkeJQnsFrcoPex0jMWZw/UVLMl/NYa8wXQ4Kowu9YUTW90tVv2gFdDxWBX23R04DYTrk8gBnrt
vrUbkakmVKzi5S8z1EergtLDn4SasmQiOKLIE/46/VSGZndzHDO1xfOBNJNT/Du/DicWPr1t5z5h
c0ttbK01e2mpRV95uqssGrT0aFqhzUw/lyJh2H4UoXDKnu3qCNgc9CvI1qMqRky20tMbkHd++ehU
F+FgFiYGjWDSNW4YJMeqFBBVCOD2ehDHK+d8336xg/nHhRTpZFAJSdUXsoGRbC/5jzx5dZPhB+je
V3r5y/gyzq6MGnM3vZeJUbGLfulnvRxXREbgaMJEpM2aXHeZ7PcspRO3lJSAwzzgaOBrnTU9V0+S
2kaIJxQlYiMlLHzj9kv/+o3C/QDRvh5WVfMKeAV+VPshYXXiUKwASO8l0zDwHftcJAbyRaoT1XV0
fDJgYtLfFmdA3SCKoOhaKBzIC9INSJLO8+xq2kT4E1Nsj6d1qoIQLmKEsR9E6FvZm/0hg4i4kQds
2rjh1Y1RUD109G2F17kySNTqcqeR5qLjgTzrakFf1cl6ZSxLwFMPhz+iw8TIxT2rEMoI74YgVN8E
wx2DWmweCvfVOtESerA1vQLnAMdQFm4U7FG7efZ3moX9ABCjTDydqFlDf4GVQQpw+P1WVFFQrCKN
FJDCMQQkFxYJt0BmkxdThgvaF80jW9cCjlB6xMQpS2YOl18jsjfoe96bQF/4/rRJp2MUq7KarLeH
S0ga7rRzRo/XuFQ0SQhCAuNc8svw1zrAML8FSAQIiSEBf8CHvSkIPxOdSt1SWcCAbmTAS8G3ZIzH
hKdsHPOgsng8DnTUTHZPAY7SFdzoRnP+seKRQwaPUTpgix/fOLd4OR10mvxu9yQjUBHCHDAyxXdX
HqwdeGYtutxgYyuYyKvhsXZOv/d4zQvXrpOrjHdqCFw6zRJghFMwD2KuZur1bd/p7ZWry2WXww55
cVx2FDomUOO8dM+GeEBN5zc3RcpkWWaBkXpRzdouKBKwVqA6u3neHkA9IW5Dsui0C2704H0IG6+e
/4MIa5U+IuKzYK9PxI0jpC37zhstF69Dkah4abUYR3PvlkB+olwLtoIi9BN3ekY3s1OGZg12G3hC
84JNkbzZY/+uj5gov1XXFfOD33LTXO/EPf6kHl47h11ynW1XsfAuRo0egrNyVH+ATnH8H6q+3Brx
hQHDWXI6ENp3IQka9kGrf80zyOJQz3Me4zhVokR5CfHu31oH5zbtyTC1UumbCCQxtNib4Eq095ZI
3jczfYEpo1GZ3VX+6F65zzCtaTdErkCpOdJhK6kXp0r1BO9Fcypn/HtsQ5hMG2/+eU3HPyniJmDd
77ONabGtK4nYBDktNbtVSbpReztzCZQjUXAMj8CE7wKyitfiJE4moRHGYkrUiN6Uk0X/dX+ORKmh
zoWcVn8iQoZxCMEJrCEAFdtx2CSQawVU5nCchq1hTZ3WJh12+QIPtAoUs4voarsNqDEqgfTYtjvC
+y7n3PQ79q3kyaUpitp/w0tHB8tJ698t2Rvlm2T74Oqpn6LSqumthTHUV359V+YTr5RoABhVlBUO
zjrajolG/Tcd8se6yKMvN1Ud/xZxgaIQoagvCqokztHdyFLFHZh29XC8L64Ub9UdjmOn6r3fI6J9
Ehd0SavLH2IfVg5QnNCVUgGPADxjPWofhyXyLuQBLQc5wNT6EmE03dhfAAlJlewOffpWk02kDOnA
EszVpqu+M7ZECeiofMR0/ES2b1YdWUG50NiQsq3jNpnaD8nfLNaNXJd3r0gfgbsZw9CMxxHxrc+q
EGCMC7Ixl8UNCZzGD2NdIouZ2GxihZPXRGrwa86jx8yGe6lNPWiHNQx62Hjor85Pkq6TL6yoNrX4
nOpogJ4y1dW30c0Za+Oo9oW8uIwE+YJzpWCOdg72DixTJq7wzsyhxDzyPGZ0+2esoxLQFMAbrTGs
UBcSkdGmh3RJZFmotGEwsUGkPHnTEIL4iopQ/zEyloAbj82JYT7zt6vA0V8VkeTUPcuUrfvPBVZz
4MDkSC8/zz3FNq8fcsVxmcgHfPGyFLb9bIHXk3L4N5uNQndVx3q7J8LOOkQDTjCgLC4f9YQd7Key
0fgRmRavU/DMkYVigfTWWTG42kZCcyszuoLf9WvUjKtEpBRVaUnQigQCChkMl75MgkaGVgn9OYfI
LP+epV3Ok2lNEMiXyct/RRSml8g94rmqtntIUOCjMyURjS4aBI27LxFDB7HhilQe/7+dXP3JhC+t
cr2cM9yxW9KsbFPSIHm9O34mP9HDLRuGDtIxc/rAQOZVmSiQtnoDGaGJEARwgCg4934mAIBDJhIG
9gXMvyqm+RjEiko29fGKSdCEUOBFZS1zEPJpzzjZDVX9ZqhGCJPvsJAx2e6fu0SAFbrso9VAi1RK
2MblCGBs0fjbEkvijy/4uu+6OpuE8ujAW/X75zFGr7LF4/wr2SgRVbQkzjqU5I1xrhQVW44bYN5/
kfzaQFK2ybqFaS05JhaqmQ0CB2lFa1DPWlxXZ25Zb6V2ESdNhKyg3Sch27j8f7QdaOmAX+nmHwY3
YisJxAhwRjajrE0S5DuWnyhrQgWyExezVIFuCiAGo9k18TURVwx2TJaRXVF8TW4394G8cTOiqW1L
KhLlPmCl/MPDDjvem/AQD8ba2jev7ARyjckIJzDxues6f7TbFyIMy5/YyUs9VxtdkD2KK2QSY4CS
SscZmQbbrhthISG7YhukdE0JqSSzMLZdsHmP11CkN2fyFmLLp7+yXFaFJLc2Rn7PNjkZqa6zqrtf
T7w3A61kMMPT+EolKGzvBf7IcOj73E2Orz3LtSnll8umtT6f4KA/d+tF8GZfbBmOuBPvOH45SkZW
8QIoQ9EqIXkqnqoMYWSQZPgkVPvUyrzn5A5LJv40RJSFYyb4JxkIu4NoXYnDylhSv+CEoiL4tNXp
bqDp7KgIASploYArPw9xSRK33ERHSZuIjg1otuBcPvP10Xz9nbnXXxdXIrw1uV4MJN75ruCILmhU
F0LdKO3DE8pHwKhXXm1NYMT5jZPjTsXJ2WwjXSXK0Rnv9/5gvIA/9tzW6ZTfQk2Hzv3nEfZN/XTJ
Jtx9nDLirpifIZku6WOZCVcdMZjZ7F/i5jxbFzOeAJPzCmGNzbhxXNccuYGK+98LmTNDKFDiNquf
qZrOiDkcv0ZVxjlpFwUfyfyOd9YcYj2L5LC3U7uod0riTCrI01KuLt7gaCmBxJQPHgq87DwszO1f
kFpdlR3mgK97wb8Y5EScitCvmhoKKSlpBLnuCDYfxJGpdCsBmCmHECzCyQiz2nd832GQHRztJGTk
Hq1M9x4nCOsm0RrCOOx8yTYClPU+L0DbVqWkTwNYfOB0nOLoYUXKcPFn73A8yb/RP3YL7RQ6Bz6U
BNdEBELipQwnb2CWZp9rR7hKYPr5P1lLBAYxrcaqAnfA2Sl0fEZqKLQvV/+F6ZbL50li+0kfdEEi
jJltUs0WN3Wy6wDn/t3zRP9/YwBJVFBjnbou8yf/03sPElsRD9JmlKuH9ZP76FKudh+cyXjcmnpY
VZ8BPZJEyb5xDUh+tAIpEI+qZimxY4teEoM2QGOC7RQDhGQuTEBGRNjqofKHw4l/7JZ2XDT+hK5q
hhiBFqlGSEjl/N2b4t/4zS99bFgnNeTakKasiwn2pnIW5wzrEnjvYz8/RQxpbub9oXTtQGz4dwWT
LkHXbjNY0JflL5uIsoq5s44HLZcJorBzis/00fk5k/kuzG7dBsUG1bKgOhRFNia2KH6DilhRYMQh
K2PTBOdjNh1BZHwx+CDgTpUJqLQ2kgZPamOc+zEeqEduWyYDDST4RjvzhS0hqXQOQcGubFHMglFe
u7YeiP5kS2n0xnSYes8aDq4lLG1nWZ4lI1MWItqnS7bdz7yLqOnxy8GmHBVqeIIqgq2eE2c5qBud
vn4QBUFj4MNvnOvU6QGQWgJz3OXt006AvSuohASSs0RXW7WD2V9T8cJjACg2ChVLKt1V8xjxbAYk
C30PQN2YLFd89058F+izEJsbIB72k3FUTKI8xJslp8SF6zdwNXy6rlyHJXE1xpyu8zBEgo9P9iPr
DC7aHuksyQpxIaqgwtlsoOjldnmJJX/CpZSzctbDYNQrbV+qTNOOIB5VBiY=
`protect end_protected
