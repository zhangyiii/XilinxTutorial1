`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16672)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PG5z/BUIxX97bocLtxDa3aPkk/LZprZljgyNzZTGF6gcxBz
LkEl/7f+3dcASD/i/KhFswLzGDUGgblHomqjZ9xKcqDIbF5CYus3eYq3X66GQ9moD1e5S0PwHKNM
GKgSV7PfsW/DwTQQ8lUt6/O6LAy9b6fgof6BRniIqWmfrvW+2ZKDRj0a68z4NMDHdecvKOkKUl2l
nmYvQgM9b8gL5l1DDmn36eg0jBgu1UIPQduSAR/75q0CHhvK/uXzV4wOQySdWX/PgB7t0P4W06kM
tuw9H0yv21hTcFFB/4FK3niw6DY3PqTznb6vSFWPJ5Zx8lEQP/wb7zo/lEtnrH6bTDIeGRmI8pfe
7+XFP/ISrIvqGgy/RSHgixar6EB/5lYlCjnzfxg9Mw99gHnLFnnvenChKpdXxgb6seVkrPYy7CI6
DkG/B/fhxiCQFQQeSAkSUAtwQ2WgEA+Sun13gXH9rSzRsOMi9b6Jz+V0cyYLd4baZX3wdSpuukh8
LPZA1AbX06x6iayqj4Bw+n2c7f6TzisSbI8NLpb7JFF5qgdTQSlzhgLG96tstEIBGqJoazqnfHo3
L5fYCDM0ck+6a3YstV42sZZ6IHU6wz4PHavg1o83jQ2A1+kzkcDcbDGZKevDXJzcf7ZtAJMOhoV7
Ugca0G6dyGSnr1z20Kf46AlFRT67LpAtm0F8j/IY+/eWE7r2OFMVcP/wzKfDVhQlzhBwJgIZFHvn
UgXVO6NPhgfSw+2/UYUAdl4oKGc++4l+/a60i+GnjpoZPAgxAkJwdM8QPU+oISzB+fuKlAqLX8+y
+AZZpV8V1cfHBCc2HQm2n8DxX0ZkEXkPkxGXcqu2wrGKbjulVpHF5j2RdLUqRK1AEiAu9e5WP8MG
uV4gglI/g16MlKNqQqxE9Y9dzKnVcWhWUYYKGfBntyqbddsFytDaQEIpO5/CoH0fW1L/jfs9XGiX
r4AF2dUF2ZdcMIH96S2y9J5TRHS05VHxsTrap6m1zMZVCg+wgM740ri1ygrEJk+PK/2D8bjUpZDs
iBmuw+ITdlbTGvXfsQy6L0sJMUNJdN+BBS8GMqK1DNg0xcIWyzyz1ebjzBCL8lNdt1eg5rii7S45
UEC5tWFG30KWG4T/pD6DAzvsS4T44HUW7l68jEAtDYcmKp6laIDhnSdOyK3fbuonaPeQRko2ioWs
pmxp9U/C2FmchCyNQPMasfF3fqFAEQOozDMwH3HtTMKqw8XWt75SVk1IA33mqqjcQ9T9i/805RPE
9FrukpybkuH8q6HlDWdAfV90vbotk3dkv94eTb9f4i+TdIEBuZcVZqhpvVL+k4jOMnja7yi9r6yA
P02IAKUuo1+UNsAW7IhozLI0i4y06PGPIJCfJNkHDHG7UqzkD+49IWzmxk+WpOFFnDYbprW2uUOT
VaBsN4iq9GIwAplNa+OJdjzyX1WiR+ujKH4rhN6K3k4otmoxgIt6IbBkk+dNHq0yRtmlMWqt3TZG
V2KCkkwbhx01iDDeny13X5h9dbSVgfgUOzXDA9zaj3Eakw+p5QfPCOmVNuSrHWt5i8o75UmDBD4x
osbhqrWZE8mJCt8gYQVyBqqA35MJlTCFu8PyTiKn0GbPEGaWDUgR1S4SHPzMcYRFrdURHwgFDdP+
rQ66CzIcWC9eCrlv5rxD7748G5zbakWjS2qdCxYSwu4v48cQv3EVWrJAnlFRqv6vzFEywXN/nQPv
rEE/ms7Po7Jc8r3ooUVm9ekapzhiEMGF6cju/SZMetio2GwCp5F1oBk42ySUpkOulf0ww+J5dFbb
R9o6MA2bO7oXAvVMaow0W85SQtM7QYqHnOAY9wYmGOYdBHaJY5NkV1WKrnRU3bKWhEJDHhsopXiy
k+YUQAvlWNqeSDD124tq5VZAmwnUkC+IKbQCpBy+1Zo5MMOm2PyeRWI0ZLHJplnEpNZvZ3XXJyYi
qLOZeuOhiDFRnmzf3ooRw/o1fFuD56uZ4DZVVM9p1HCDrEvhA4bAB7misRjpdchkzahOgyoX217/
TEMMD8lnzqETvr/drTaMuLIbjNjQM9kH4t1xpcROYddwftX4Liem9JVE2bfDeBCwENA936S0QJnB
oeI67hd5WLBV4oNMB4q+NNBQ0r5waa8Jx/dUFdOudzJ4hU6NNpcxEJjeQ1ePARKOwnE0bpk/Rd3l
VsRXwfIH5g0sN1/w1vvhvcPI2Ygzsagm7EDIT4EMgGSCNpjjOWXKdoVZVdk0u/JUnS7bRAzi0gIF
Tv46pX74yFIZCg7yNQDQe55lPjapiLXrU6Iu0SWjErUslulakveXckZxpaUM6tEObjarhgtOprxh
Uppf+dTQ/1guWv4tYeE4aJi9Sea/XMu6I6SA0DoJRl750ig635cNpBlLhvv38ri6hJ/WWxunE6WT
2+i5e0VOjvr5RxnDfF3AnAc2PHvs7WHdpRgHKpM1PxGetcNUGsP5/znc8P43tiVIc0xK/5L40z2s
PxCYhPSD1ryAEAUb7eeo3Y1LCutlDdQ2+ezmegiilABwGcz02NmACpbzkiZuR+g1dfj8jELOkO/O
Yxa5xajzYt51V06EBe7NiEKX78SwVlmxoojSGBieKzSYBznC07RIY3dhv8sQGQs1v9DRHshIUwRx
IB33316FwuhMMWpC5baE73G3+fvRap0RMkQ/wu+28l6FvN5aykSMVGsarAAyauKApB5sGCygDdhn
BK3tvBJE0hjWjldWw8cecTwQEkzwUbviPdCpnkLafxAFkNtFCWxRTPtP7YonzXFZaDbpmB1IrOv2
WR5dKCRxjo1D8YXh3gn/ZPG6y/uzyX0qZwRBKPiLFf5ACG50x+OgbxWnOZ8whIgTcHxfmRzmNG0o
WdYa8rcDR5tmFUEJ8p5gOmS3tFIXx0G1GOz60lo9UqyRcMOvJzZCh83LJQCsyQtzVBchpXJEw2cl
1sJEgQTBMjspNPxDy02J6pAeWfz1gK9O5+6qSSuNCx5xYLU4HzYcwsEtK3hwYI67Oy7kW1kdD7+T
k0DpmJbHMDyUDGZsz9SoOlD5xY8+jYcph9RnAqIH8bUbueDFZtN9xOMdbaKv5igxSMXvO8EjafIS
qrDepc7x8eNvauatVOpFr0QAPgVZQ0ZFLKsI3sG79J6aSYBkjhrlkPvBSQcSQyLx6Q/9FA8GMAoZ
18z9tUXjXHa/5w9TWXIh8DPokFfcjeASw8W/H9TjQj2btXtCcAgyCeP8gKu/n4JKSb55D6o7YvPn
g4UI0FFjoe33w5fgOqxJ3nMPyygGLNbVAjrfJvPg3uAHqweDR4rQ0BwrI4VfYWdi/npxjE0P5G21
3PnNbS9FPZnewHQfZZkRmvIyNY7YQtwzyih1tklnYXZ6scq7oHA9/83IxVwhY5R4XYGDjCbatDW3
vuqKkwN340iKMNpUjQFg8y7Wx74odzF5RV/sQsKUS7McwVEMOAixH26CRAAY3p9srth3TskkuuTc
I9PRijMM6jq+UR9B42ePqZJBDH2vwg/6teKAX8+uEVOEX6aDhwdIcUn+BeuMiKcn+ZkwfQ72+E/f
kmQxmpWHi/fO6vMo6POhAVZoep0OXKVwIBogr696XCNPJSwUzKfMyVwDadABwnnSTPpWrackt455
wzwlI1KfKCiISGL4/w08Kzi7OQG4urmdUiBrVl0Cc0Y3WlliZkp89wnNcpHs1O8LeM03lx6Cqm7Q
VK4/thr+FROooWSQXSfPan83QF5diINKsIAU8yVq1ffhIz/7Rj1BSXJYOLO/3U1UXe22D0+Hbb/t
/lZi8gBEH9eYOQaze8W9FascY5X4KTMXgeuBd769ChXFiSLb8HSJw5hgXt1jFHP1XEOiVNXU3Mb7
svbcEZIambKIhL2S+75ZZ2pq187fP4NDDKno+Is3zJxHKLPlvSUE+EN4GKk7w0hcbur+sRjVxqhx
YLuoltfcOQRB7vrxO58KLX86gcQmcSS2cIRGDRZCx8q6qjzaj+p66YjspPU30o41+JYqXz9ECa41
meAIUQbaH3kKZCTgPD9cPzUpK6WfSXPVCvDjBXvQlH1KRuPoX7Y4gA6YCclQzI7eLmYIonHIFovl
5v/Df2jfbmJ5jN/CkHFawSl7OKJlYlxvRDguVtHhLGrfZMnCVgOZjJtK0orDZxVMRsYoM0woNCu1
01xVWvm2B/KWlZN/FP6pqre/9pAICSnBW1Y2NRyKdUSLcM/PDa7LbqEqCEM7u9nIOUXVlcd5NfVS
b5CzOLi8nRuVht/Ew2EK5Lcs1mzn0bklWgmjK/X7gmGl+GWYZ7WoN5qqZsL3Z78WodheuX+DvmQR
T+csIQ31R4ijPJ6qwqUYtycFVr0F/IreIqqsWCdE8zaPs6I4jftAksG5Y5ezzYV0bJ68tC9Qv783
xD9/sznoPhp+tCnt5UZNGapT7gsQOSm3gThRz2QCllavguGPXqBKS55ZBPGtodUVokcpch94mbYt
Pbr0K3tkV69LUeNWwoZzwKMPmaFYIfbflLxBLvQNbo16Z7L5YmIvIgRvGLC/U3KUDs1liGD0e7cv
f3kdmlWprzUTDukS+VkLEl/rwD/78sZ+KDg8XD3i6HtLZe4j0lwTOHl4TSkc7sXM1yZ4gUGKKuvY
BBqjd2jGs9Vf5s7X0KpNd14Qo+C37LvfyPjzgazGmJwV/hK+3rpYTz5cQjFC72rUMBkcpGhbl2MZ
NAWM10wTXXFgOLxWKTDgpGMdxX5DYa06fRO78o2IZRj4xy2KZveOrLQ59aZUl6NTEYpJqw3VsXql
ewk5/e1b5+HBG11fNVSf+3bjuLkw7S3nvJhT5QSdVKrtWuTZhVaX0Ax37PtSpH1iB1F/f/c4vJaz
vXuvofaMNdORJYSW7f4hygh8jHQKhuI1B0fV13zGdBm3TY+SAjXPg0Z0J4gDygS7d4hHcrY7zwet
SvgalbwsEyUdFkLx1+ahBuKaMZNfN2x6yLdh+/+Rih6kVNWnDab/6uRewQZYQBPWa2BfBzw4C2aU
TkVrMjRokQf1DFFpdtTQkixSk1n4VpSEG6FtaeoC9GGm63nBAVZ3Etw9glNzzEf0xw/DdyIhlLcO
xxHpDd65ApdDi1CReEQSxMG2qdMQNyYTjOM097DhJCYnOeH02bB9Y6tPq7FYQ4vUVmv2usxPFHwR
npEIQnG03t/oLpJCvrHFx2bSgPybCsobnvPKverd10UVNVIkPji41V5Y5QUvP1Nt9GlZx5z6PWCd
VzyGILsLMjTQ8VuKEGsYknSOwaJxUipkSVZ3igJeF1lBl/kzb1CqdaRWwS2zUWaAjz2LhLMXMb3o
su+RENqOz/T4GqGVp37uN2O/vmexLoaUSXXoAfjgK8L1PnVfX99PPy+YVFUxqqet/bFWYsY5qYDj
xB1QurRP//WEOPEtmG5wL47fhredfg0f9dPv6lHFWaL/3YZJBGb6q1L+V2gaRddiqNa3B+ZsiYBu
F2bSTGYfOJfAN74Py7M/9A7/wGJ+9W0ZwB/9vTjaOy0epSqvoolbDmE+jA7QWXEnUIkm9L9KxSjA
ZUAbGCx5bZcHuLBw++F1ZYVs55XQd5ZYtkLOuyZJLNIxzQ4OEmgcExcREmOtCwj+lDE4VeD0NMSz
56CMjwHjscY2+wDSnnZU7bgUdyAdhhbGZ/30eMkO6vhTPLxSiWD37Zf5+chJLfpeHtr/YaJdOQFq
ibAcbG/8yGc+7ZRmsYocHwiW9qZ5hC7dfCfj2QrHwhq43FSuLRFQQg/8MX16iXKTif9gKn/4VQVq
GN6E1DYthM3wa0Pa0VOpv0M8Hv+bXimTmd4gJKWBUXlIkdVAWD2aKujJiA1EiViuWhJ3feiBWdR+
+XHmpQuDFmWq6xr1pZsJAwSCIYyDjBEOYvzBKXNepN1Z9MRnE8K6FuV5mXIaaeI3FsfKsc56tf+V
S9XZQoSrKVJxlATJ+NIwBrJij11qujL4UzlLI0rJMRncEXVZncZUX5fD5xwgUVF6dYtMCHOTMOb/
ykTUhHiJb4wd5keXdPyWcnMX9mxTz/4K0TIEpgeddm8sZUvOlnRlkCFHu6V+aNnTaW9+eoooIPTl
Jd7qPaNpgP0yNlod52WwZO1H77C76EveliqG6qmJEatgxpPVfWxFhSIOUyYpOhKrXpOYyBmveFXr
YGUrZKAuvNYadCSbIEpmYd2KTiq6RtyDkPCbiU9oJ/V9g83fl+K5aOprkgaGgQH0aKUi7fh/is7l
Yhp9pYaq+JUivGVuIyj9fmyJyRzVb6xs0ti8FNP7/n73Nffv6ieekTfAyI6KKu+OigF0P5NIDIP+
uCpHE3SN+nWoOETIRtAqbdnD+OGFpp6bx2zXTWnQPfoy7m8eJG+JwODZHnYUeaANunfiVrXBKHQX
rkICYUFATm3sfS3ZWWWZ9C9ar+dflir/70MnMQcDgBLbU3/mj8KCto/uqtEi9peTEpeIGXSpU//e
hh5+BGeYwBQ+NK7gw/2sGHZhA/lail+MZL+XhnCqZ8HyygqcFRP/kN9C3eNNVyqpRy07HbPdlr+8
UpwiuHh/U2etfgjBBnWYLmxby8u5WQ9rZdH0zTHjI8+S1+0HSiSdjIkacgAGACGamKHN965+AYE2
7jmsIcbpjNVO6aQgfqxBXujCtARkQO2Zi4n9RA5/WDziVjki1YnHQka1iexFuvmyotOUaE0+9ixv
qUdZDvaKMpKDLa4MMXZVxorh7OMpmsd8NU5MJadMkD4buxXZ5UvLUJ7ts85vEJJnFvBjYD/niFfr
cCrCs8xItZKGZWUQOEp+HUIR6O0IU886ojNBhFcg9cApERWwO2/Cq54DOL0Lhnmjj+PsTHlpW1E+
emGa/WR09R78fkB0r5nNlJqOj9bvZqa0v8NxisbkRLhp9lcsvdTxc9SkaeeFG6ZD83OQu9ODtwgp
FKN1Hb54kiQoDmjdik/ZFGr15L9jwzqHOGFmnkM5kPXI12ruoV9lECA/gjhRLT7eHDfuztcckGUo
d1sNxPwIWHlJ7tQecxhg6xB46fqecnB59ihejrE/Oe49d5RXPJ9A9Otapxr8xMLjrVenDkfKQ74x
PwPwKRpn0Qfk9IQh1jhRCOXSIXFgIywfI78l7CPA39NfFHkChqjBiURrAJIaX4HIgfXvrLY/TT1V
xy6+KAwUodBJA/kNofwTgsOKsQe9lO7urIwdkZfP14LCAQxyPIGZFXZLZ7sFXRygFoLfLInt+cSq
n96asCAc0TIAaiB+3Dxxi08vXKJiBu6DCEhN2/KiMaG/lev+Mg8Aah60I4J0pv37o4r6a2S6cv/J
iyhC3w+XiZ3nid0PuVyH3kEuPoOL+bAgZrnF0n2abAz00+yC7qi8k3UCHjMXF8EtR+8pe3zB0t1L
tgAG26Ueo4+2gAe4Fe46zBNAcprJrTURhI+CQik3AkSLkZManYUfJwTfTb5Iogd9bmyK4wplGUrp
jLPtvucgLfbT44wUAWLyw63DHN7I+C5JuVXgNrN15C+wBdJTXshTCBmI9cZkMX0fGu9unBdy5O76
ZZaj/1HS1nj6Ew6r/kYh8DBvdH124x0e8pbLTgDOb8SdJPNg8eQ9XUsIA3Eos7o5rJLz6uqE5zEo
JNQxi+ScIxBqefAUtE8teuwG2jvQa/dveH+kBaXTT9wLrbN4ix254u9CNKAMy0I1xpo/JRDD7Nzi
hpgxLRHDIJNRI6vb5ZYou9OPzd/QzOrwYnO26dQ9HZ7mGc/VTsU3aelXxEoBYZI8JCk4K5jWE8Lv
F4f9iBmzdYKO2OPkpPcFEnOdYnfDus+BEEVa0W62LMRVdCuVzjpBWi7WmxoOsylV294Z73lGt+2e
AkQ7WqGZ0bbO2T4VNy9uh1HmmrjGYdyIkVPycK6OecPUdqIuN5nJq6QOZuDFajqptvmFSeG0CxKZ
d3iEKre/vbQmKJ60R5DCMiyvP+93g1DAhGEsTfxY7zfg5qh2ArVGmU0uYN5Tehq9i3jBV7Xd7w4T
GKnV8uBT3RdkfuW+Z+vmaNGL8IEe3PhCPbl2B/XXapxDwLm1y3FAJNElJpRNF+EWtIIjpJzWrG32
R3OCV/2RAdpNrJaQZ1CsRdm//ItyX/KIB2VKiM+PmQtcWMWGnUfuOpbl+MT5rFcfArs4cOzb5BnJ
NjtJ7mjqgLM2l9W829peZUkH0ddKne7oHl4qz7Cw6OisEdd4So5TlqpdnWey13By0EcrHSMQZ55L
8fl3VTM995ryHuWx7/rocXyWovRMAA9GRBvJ1oodt2CydN0oBobRVe2WqGq7c2lX23FRHxwbdHsp
Tg4kY50iD74t67som+NCnmXbj6NBrdcmSLUtaI2weA4GkcoiOSrYwde5GHEL2FhUDgOW6ujiKZGF
CdfPsilVNHizkAySzsc8qNJqcUdJXUjZXVMInRXduJAUq4NKprjVYGZLy+gsDNMLfiMOnsaj93P4
57pZ/yIArsS4sN/REVRKxygfd+bxHewx4KDtTfdKk55IpbeZqOxyr6FYpAyQWklGUCxkbvmlb7cA
IY4nvB6WautDqRhSW4fKv3VTH+1PmtNF+TDB/sepvy+DDSQkbsvAh0IJcs4DmFkBgySyQHak6svf
ssYpcfzhulk1hO4BcGPZi6oD8xsSmEWdfPUPkBXbBPoawba9UsrqxQ1M3Dl8PuloMnPE8cx4pe7a
FJ6kGlPsObhP8UK8NppOob8DD3J1dt6RT/UXn5e9J5DGYc2agR+BpD+Ww5keoXuHNEax2KFoZkb4
nu/D2IfYMi6fBPlSf2zPCxDo/E4cZdT1WOGfymI/AA6kkN3wRGvUVSgtop2JxR8jtO7k3VGUZ1D2
QXA0tuCfpN/esxZLRFn6OwYwS6r7igupl7KPmrrBub/7jRk9KtQzqlTn/SzFTF7+J1/ZFbiOjINA
ZFTi9eot+c7SA32z3GXgKvm6JZ5iKlwInRb6WfQ+SH6hGAdZGiC83uPXaM9dSn8ImdFsr/LMaOMY
0BVXu/afdKWFOPu6GjFxIzmkFIIqkKdS5Pg36HR7f0l7o4YbpMJqntv9MYNba0x8Fxzx5GRpX4uz
rJz//Nf6M++NenF1OfWRYXRb1mf1UEGiox8JDxhBYQFHXI7MhS/cbUmQGj0bSJS5xd8dBimulRNN
FFfMACPNDETWdTBeXDZkvSbiSuFLhpV9mR8rDKQeDskpXR0+yg4cCrS0wWsDRUIwVnUnAHe7y5Mp
bgW3pysZDM7+YDTYj/FrcjY4HAsYpk0GBjLQ32dXKHMr/mHl9FNrx322vW6+nLOAydhucZ1aDj/u
3yTgwPhfE4pZarQt7eRX+AjsMM74UyF7my+ZOhK1BbL1yTNcPHQs1bmXzHdtfbdvlrBgH1PEonOG
JHNGbgUboU0tPkkkm+3rbt3Du+P4aSR0HpGvcW7b0r5v/AM97H/DBQP8qr6Rt+D5Q40Q1IXe5ZpN
oyt3e4CBzU1+zaQ5asd0afT0DCAlzR2r1/kP4dpx4AFKV7/SDqmgCNqXDQ9n3CnPoZqCQd5Z4/BN
DFojZjqWCerD9UPzJR/c4p7rh6wjhJw4ya1dUajxsfyAD+jN/dyKR9wAVoRD6lnNo0JnjDT4SmnB
42zpDwQBnuZ7WCNVL3iDHivkKRmfiuiAbDnauqvf0PPH6hMVoQyVBzWuG8RbcrC+esHbnL0jHpmF
FKif+E9ZxkSNJKLzrMPwK8Ya6SPBZKNqiZTTQ/VVmlgIroxSdDcfiNd2FfMvOecTdSCMKOUPxyPv
/xGYuh5p5TfsRCxEqzDYWfOqBTBLjZkxm49vdc+OYQoZ7s5jkxOeqNHEth2EUnC5NNPQ0EoPuxUk
UkIn4qjGs4TNwsVCEF7yR66fHWLsmKLoF73qtJFOULHj6VuodLpT2nKPIeUQYkfeRI0CAjWcgxtf
w2k9IJBY5FTJL00mIzU6rzdbiyrqvJdk3LEC/e45pOQwBWReQ93oRsplU/z6pVwmCilIjNm1/IdK
dA5EshCTzs7OymTeHM97FS2iceW9yP507cv3IP2R7qA4ZAZIqo5zqz4BGDDmEfZS5QIPsH5SNYnv
s/cTYLY0cvSqHNoeYaruTctVw9qhXcf8C0dCnctrGdeCxjaGMRj919pkMAFZJ83BYMygoqQCq3rQ
dl2lPQ9CnQ20DsRzSkkFjWTTZKypbrVrnHWeCPztEAJtx9NplVOu+MBem8Dkx1Q+OwjcOww1reud
tJ+iKa6An4VDXAOA60kATj1NaqLVfHSojmBe2V2JHiVCN2+wV+EjbAbgD+63ddmZtNS5Ui6yiX7J
bvNGXNY/qYtF9M/AxbfgTeVUvH6Yz9bfll5CVhAa07QerQ6dJYQUOQrDVQOjbFIlzB++Px6RvlVx
j1xzGxyaMyxtH8a7avtv84qDrLVK8fHp30N3ykTzxOu4UNW0cijG3xQEno1wW9SHkoJh3vz4qcHW
7A9GiLT1Qu/HY/O4R+OfPLpAW/y5UJSuV2Hx3iJuwbFnfccE7cmCPc80PNzk/ZNJcoEw359drfFa
QaGQ+QEpclyA5ntbvMrSIuHZwCHXXnoIjTz5Dup8UR/e/NVFdG+u+okC0X73vjey+WIB39Utebt9
8VEbk7Gas9VChK1xUepX3vYCzT9hvS81Aezgcn/RJif7hmeEwh+xYcZLjpGTldYEdggUVw1qKtXU
gvf8vOEC1rdcUC5czb5Mj4H5Nvcvh/1zo6Q8cFgLlHR1RM3VxNh2y8igt5avX0s/J6KMb8FVzO6p
hRXa2gDEEncaoOMuolio5yADUF9iCek54vOWUqQWRlZoIJPXuohYQihsox7IgBY08Emoki9K9I8Q
YKSYXchvWJ3E1n9Yg694rZdcNk1gP7A72ZZEAxdlIaG0RpPt1/wHqjXj/sHuXuOiiYdMLh/unUgv
xNx3S/aK+ET8DR47a14AHEAh8WPO8EIP1oO/WjuynU1Z3ZtuEPAV5Raqrna13hhLVYYd71xdNxZZ
fFxmFzJNZy7JU9MpnLHFFOCqWDB5oBmGQ+1AFSYNv/QEDSbpopRV2nnuQYVX1ZmX/gVGc4KLmFIf
POm9Jb2jp/ym2X0hdJZnvt4q0DDw0f1619FJeDRcDD6yzA/FWkOJbE+nuTmqLz4qs9j5U7kJaM5z
fz1hO/rcVdk+2g1cj9foNDmCPJPrDInVU/miuDnuuDlBbUiUjv6rerViUuObYVEugqeGOag3uwbY
3alhaBM5r5zYVRvuNYbh0uX4UQBpM6KS6+juGaGgGDNYUunMJcTn05BIYjTAkNGMPeLl4m+iogAZ
8AJmo9mmqneZde+h0Ep4++kGm9tlwz0AV4gEtBCWaAXB8XlPINRX1ZHUmlOnty4RpBxJKd5MH+9y
efLBiwDPa3YiCrvF6zA+cwIAnQaeB+YEXD3j4HiK2kMdp41ZP5XbmPXjx4LwA4svCJ8Ng02rkPml
Gw9DTxuFErHbbBk7TdHDceTJM7FdHtBbAGV7LdcjU9iJ9AY/WiYza48O+bt3jJ03Q6tQIbfhV9nA
hhfm6NwmByGiysK8uai2n1KW6SHDZtCfwQRkj77oVXVhJCg9GHd3DssslS5sw9VYIcfUDfOSouaC
xUgBqm0ukl+H/vGjCvD8fD0Kkw2+djRLuArPqdNfWPfl3DFCkQIF/rRzlf4mQ8Ka2yW8qVN39Eo7
0uFA3KiUxoXETnYN3NkOVTxAeF3BcJk+8ijB9UpBb/ahedN+PzI3d93Y0VqO78aDWPXzYcR6GvRw
/8/yDyyE0tj73wQyLarNoKkurbgYFE48dg9ZAgfOigMc1UX/wb0IIwjw5D5oa6RXtQy2oDGjj9fQ
5jj+Gz12LSGmOfffJVl7fVM6ZMl1x/jgP1BU2rqoFRfY8mwNvOflvqNVjMoT9esjx1eHU8dfw6KF
R4CMtdQ7M0s/ZRsI0fs1yjeJvWrDaX9T1LlujJjJw1UOsdj8EJ3mNdsawgdQ09iyJUvkwl2lWW48
uZduClfS0apy15GSzO1xcevdPRcM9pUjMQ0tiAQV/M47wGmeWF5UxcBP/bTtLc7tdmqMwSx7qV72
tbTl66+fHJudCgEswhocdETbgyANnDDmtGELgKe8eO1OtW9T8lNNYStauKM6DHobjaV1Ip0kFbvu
FccYaqivQ2cDE9zBCEg/T5lTtbZpGOH82xGKKUEvcqS+Cw1Dbn6DMLisfQ+2sMdyUNSNM6SRicXE
YuN+Z8I6pdG/JZs/SNHKCHgWbJM/aFwMsZYH0I6lxRCuc0K58ViT2wjjqHl0tjViBiKr62ifCkWS
Kuhxgf2ZtVvqrrHmLCaaAD0yd+4zoNQrUuGBAkIOYotGVnddUObwdd0e56bakDSUVLJa2ZN5nPvx
Ps9YOKZwae6nPiHeYJidNITXYWdHpUlgBz4X+kDa0YD5TRVhCPNIsziw1CiWwIcLZvn12786nEnJ
Onep4mvGtVMskIZmAAdL71Mu4V/GJYNBursLxAVqNearYwJpmd5+YgnILF0Un2Xw1AIxxeisQDFt
Z+eATJgqwoVsYudq58Q7MbGkv8+/jvbI3coWPSZs2YVnrttklr9syaIhemv/aDA9Tr6Lv1RzB7ZS
FUT/PIAeRrcAdvrAf33XSBlFq4mtOiVH5094N7Hxmsj4NUaMbKZKXcHPwTO85tJpIoiQsNCtynDx
dJxjYE6nW7nsUq+5GmibjdqJCAL+paeq161XH4grS1cwN+jYVZSF3MHuVhCdU1ceAM5RFwf1QCd1
hZe2bSFyV1wS7QCzWQ5+hbNEhdj8zLGFziNJbik/L/vgKaU4P7VyGCAv4/E3tP9bIxaHNXoyKGpN
oiuAUeo+s1IlGYfckl0jV6QWefNZlprnk9mty8uMPtbHwiUC4/9mzG5YpzyCvxoGXQPMaWkxhizn
QT3hAb5VyA/f6GyEF0uWa21BZzgsYNneRQjVQl8wH8PNTRvHXw2l0lhlaf27yCT+iiINWRc2by1S
3ZZG7G/k0bWplEnHNGsq5yn8v9Ngw/kHQnPso0YR+cxZse/HrIkINq08XmB/YETLqxC42d4J8VMB
LcH7PE+viYQcMWHVT+4e0AESKgrta95h9NGxAvT9P6m2UckyOMopUGR0e7frfGuTThkmT/YbHh3e
VNGTD4+6rhfai/IJmAErngdboaoAkWEC1acxiE5pPkcP5n/+4PK1knXltQk1sP5iox5DliFMDmAv
Ni6bPkl7OOQkq11zIeBG0+7YAh4hze8ld6uj1eTwZTRu/g5P+ETcZ3s3reqVYdoja24ktpF8Nbb1
Zr8dJ6w3rsMzAGydUgxVJ/6XhiFzeWSormsoc8F0ju/fFtb/hXEEvKNDZMjViVmG4Dknu8T1qyWA
rdPfpCgVRxpPggyO8w+0/vSMVa388biirNPfdx6ykf56wmJrpl6hxlJtmEbMAnZOVgb0RK9YynYI
pZJ5V2tNnnywVzZpXZw5rsPEXV7dLYKQ7ys4MsL4PXayx9vOKUfc39QsLULHaYyiBOFBq9ls9g53
bSUZBRQkdaGrJIlz5F5vqSyYKL6ydXGgj4OqVb5TAmC3pwtKfAHzjmeox9LrbxMayz80epqVuJgv
QGZmNapK+LABsv/udm0lzc2HSXdv27rkZ97f1ArUA/wVMgxsFKfvocWHJg04cIztUkRhGql7VTrX
sUTYJ/qG4BmpV7Bm2T3alqD3ojlQfyvCrL3YxTWjAIMyZkbbSmWL8anv7A7BEiIr4OxrQmXT+PJV
j4YSwMnAU5mJQ9n299BLU1sfedq/vyVofNK1pFQK3/6yYlyaqXiCSM7SkVyKjpte6yG6W+q9G9p3
k0QY0AKLjevzu/IPBlQDOnrlPFXcgN1ycojFNh71Mh396AeK1LhJJmryq933GRb17kXtYXTfXQ7d
79LMcXRIimT91SRPPY+8tRknQ5W3HsrXvamq7FyRAPJQl6C3PcRr1vAoejHTWSm3J+dD7o5O+RiQ
HbfEw7r6QhLrahgTC+h714j2t7l+528GyEiJcCr3FyfqOjm7133zdf5WsEycotLvFh+uxvyLAA9e
Fj2Ddjc+7r5wLWnouwsdBMdSGxp9OqMPTqH8rkHt1Yfmuf55gvuyjLKyOnpKTLThcqlqINVV5us5
ANUjM6962S9H2M+l/J62JkMKmpbVcSyZYyXg+ydMDQXgTRgylJBG6n0u8OpAJ04KFvxUAGFZVw8w
rjOyqNZkDKZG0UtTUTcLHFCtFyHjkGpigwpbtqEXix/tFWnC8qd8zYjerSd0poDQO+9rx+9qvrsT
JuQevQLWTg8D6e8j8K/Uh3iArg5dINyD6WJTAKl0leal4zBN6Mzz6BKaV7vlE6gJowYR1bHv0/FO
9keEZKMg9U8KsdaQLy1PSRXRHS+778XCx8KIO/cCu9BW/xgfdq8XVknUSWA/Tez/vD6BpG7shqsx
GHRGCclajRZslw17HPQ3uI3agWdGHW+omLA1SazD/9FJF2cpkBFMfoby8UocAEkr1TD3/EiX1Zgb
bLpWrEHEH/F9gcNKjq6sTntOb7Ts+tACBvtGKorEv9Qm7U0kLX26SN+rJ/9X3ogWAINDIch4zPUW
xwJ0wjx46U3fUCD+vs86/7q397XL4wkjoU4vE6iuEkhWLQNQ4Dcx/wmJIuEJS0hHOSS0fsz4fBcY
657djYJwpG3rRaoPg0wJo1GaGMOvgUfRvzUJftcMFK1tiOehVLcpKbPII4CIJnv/kuIXg+OkQG4q
AgyG0DDg4bcT8LmcYCT7QbFLAt8tZU7UpT13ORw1AABRYljcUA6Lq9vOE6O95L9jZTVtbKJkgl2Q
JmbnxOxYNKReF3JRcN540ddEQljoFFOFtc6OT2W/Yn5qOFEUfa6iQ6Xv7vZ9ER+7xCRAbhiGr8QP
lyATMM2vKxGJYgkfBzLueNxwfPX6B6mYaQQy/QdJNhswWGXbBMA+aNjw8U1wz+sdagSsw2x148ft
O7l4U0rjpp6rviA/8I3acV6jFWKMuVu2QUjTBzAboY42lj1pJHAip8zi1d3meh/CfA92/hxcl7X+
QL4V+gwOL9vek00Ztg30axA0i2pX1olHlEc4sERMYjB3IQCqEnRoyki4jFNDAVQa4h8sHZU8LIM2
QNzgtyne+103Z1yrOKHs0LcvRoVmcA4scpNH9CI8fVaV07xuOKkRq0b6gRpn+aryvaIVmFgB43Aj
4mAUW7Bld52UBzYXtsXSyd9UHHeDSb4aQdaulUImo6DGVLXqeJjErLRNEvMl1xL52VNyG2/fEAeH
/3EhW5HJGNDXc1vKe4KmQaBfFPc5YYFkLKXx06FGaL/4EU3RevSsHYdZDxf7pyqfNwO88ZVZUK3J
m9GUHUbfLmTQYoXOYDWIg3LxnkXrsdYGLfgHl5TIU0B7utznMt+OUWIDG6K/SKYIMfZLt62WhZ78
0G5eiSOjq45sUOK4Y3OS+HVvHab4IiQB5hs3dJ81OOis68Rt834bkxqLHO5iwVudl+YT1TTaRcJF
hrijpASbHL7d0WqfRXQjcNPM3+YvQF4nZ7Jt3ZDZUYrBwoNwBE7FRJE1/Vr9rCNhSFE2fxJDXJDE
fA1vBgCOG6IKkmoI+RfqxB+/PkFYURk6jwnNsjaCNa4+eku3O925MN247p+eHnE9LQ1hsy+gkjwk
JoXq+irwWwSxzTfNO9lCAKMRCnn+q/jTo/Bx1TTjQFGLzsJwjetcSOofoqbQJcqjNq5uS5ZaKJnC
VAoJ83/gAVScfbqNY43MZuse39v4YXl/E6GxPKxr8m/ykDly2TV6tSWsLnv+HZy5LtFhRqyk6Zfa
WcSTyh7MbunCdFdMTFbTtiPSwqhsKVK/gwrkepOEm/ykSTxXKGbZelxyM80F9SerKMsEq7TF5SlM
EX6P2bdmE+q8l2v/xFzZuJAzfbS8/IFgJun5Ln75kezMwpyMAFXhHgBY/Q61PuDT4rysVrK3hEJq
v/9QJqcbDKWHbKeM1lC4V06HAZ7y2FdsC6aTFApKq6UC/XqyG0/GHJxIxwl1pOUT+lmvtUZbjVG+
u1iIXZZtP7SgBaoP19R2sCu6hcFb8DhzYwg0KwH31O7lHrJXozyS4DiHJcwRr+7i5cWvj8+bU/D9
xvQJ3weCkDUQuqvASe6nxqAYFsAqtcgGMLVuuWOo4fNw/6ljSKxvKfuSRUkZLiIQqVzLyanzEVbo
Q85XcJ84IXJztHwvxD/nH1rwseBxsYHS7wInmT1umY/r9ycSeVpgfTCsWD4eZcCopqIom+ZNyxu6
NURzY7qI4tkujDNDLIFxgCdS1sUeib2MqVBRrvnx1TMUetEoyHJLikgb16uw9NtmSB/Z7Bcz/zT2
r9kphzOj9aEVkUYKgtATUP3Q1QUEHnhQzrutEPrbIWUIkm/HWEDGqa1tryBgxDacxZuzoBSX4Gqi
xK4dA+mjSJ4csAY2qZNeXYv+CK7P1IaCHnPx8KUU22pSFUO4RfA/HFif0hFT1qxmXjlCRjvaoO4v
zIX36+O51TpwtF6FFEuZwh3Lt4uBSOC9G7gz51945C7dgA6VoLhd5xhYF/X+/eukFbpKdH2XfPDb
PApvs895sVzLoXj13Ml50ypyKJTt3Yf8yNccb27bUNoa3ndR6lkjXyalP2LxTkpt6bmG6onEvTLJ
M/aQl5JWvaXl6OZOnrCyMp9TMMc6f/EgzDcYRcEdPZ1bOXbpAeAv55dxXq78228maBuWemC2bUv5
NlIKLjdW4oKgGvtTwHSgAyCeGBQobTgfiekJh99jTms9SPNfwm0uY9ZaATi4Xt81jnjSPERTq144
IaQ5EPpvAYl78I5ESroqwvnk3o0L9sVLtKCCjAiO25ON3vHPo0MmTOd2iKRz4LXzw2FyD1g1MzPa
2NdqjkqWDBAGxtCqTT86r2NumKKeFCcDVwke/TVxdz2Q66hm7VnCxLFsxjE0i3PJpxS5qzhJqz46
EP4ylr5MrVT43qPAvsskXZA2yCrumXMG2rDIwn3Yf3JorknF63T01IamzUbUjEsse2fUsV0ApCcK
UQ31vOWpvgYjvlhR+hqpt6qm3vVYE49xf6jHp9Fg7Su+B498E53lQ6AZ81PvZCBmr1hyVc5uzxfv
++ekrn8E8usCQFNzpgpGNqUrGXPcArXMXc4p9yfKs/4CJj4BNdmvgqlQDpQcBECgtrQIM+k+tOlj
D5ze8HWlRUWexXIYidm1MSNcmdxYTVPtFYKcGlkF6NlBHl5RfPsUGlJN03H2waEgT8kklEdwLqKk
y8QFpfbdw83UI1CfAqfCM6ToC9aCWh4Q/pmn6pNy8g5EQ5HHTEQWQ34dprqeVyY+8mALszRUGF8x
Roj8OxRnntOl85MRU5y7y+eLIFuCDvcOrNug/gAQ8Z6NpjKnJKIqihyWnykmWdB8Q5UrM0S/SgJD
7v56awrOc4jLx4A/mD+fmAd/gvgzIYS8gEJEnmEMeXq8GlEuSzK6eda6WkA5iOcMWTVGv01dtbUx
MH6Q/3dNTGVOnof3j53Qw+MmAk+ZafpEiHaEaolHywmCIDU6DFnH1QQqKBME3XjsutwcRQbKY+D4
48ctpdUqH/woVtsO0K2IZi04ILB+YLfxRR6Fg2nzdlfVDNPesujdKGK7aASn3tMC8PA9A24RZe3f
IR+ZW38jg2B/1MarRNzPosnyJOoczZ6/zSppOXFJWkSJpCpHs1nwU1/kGq7s7znNrQURdFv2N0Wr
fyMTsmmHeLatPfO+n3A96BuwysZ01LfHCghA2iNTz185Q4At64ePJQcLuA1pNIH0/W/15I7waTMn
zUCHARiE7PUxLCRQn/tCrse40Nomc9sLxptA1QpVxZHZGgL1DE4Ej88dqTNrr33QaBeyvIyZKXkF
a4rC4JwPEjEJ2F5ipdFXAoRFhAMsk7qqlPZezTzh/G48ZOxnlAPBK54OPkuvn9WhFHsxIMu0iH3B
KrTkwDfjiMLzxFlOUv+D24mFSqVCwk/+DCV3cofbn1i1SL7Uv+vt2dC3QdN6XWqm5bHCkyYZoQc0
MoYkv8OuLIllWpedARCj8aJo+p5nUTF9BIFU+AVjRsxZmL4OjBumz6G+G1goSrop6qQjxno7UpPY
sUc+W/BzKxOsATjerZOTKDwKZcEYryiV15fkkI+JDu4XtZKe2XcfptFRQdtcRTte9/V6BJlAJ/zx
PFVGAt7jgw6niXbIhP574tHkxOHqIJft2Iai0EqSF2EQwRcwfRayg7Zv3OAa00mP78/tfoXTT4DJ
uW3gVI7jdKdpI/ZdHLbw7ScYIKaDpufwd7IqMB0OP3rOYE6uH/Sg6F5Ag0z+RhVbxBeYGQFCqXPo
GZXF39j05uAJSAbn/j0JuEHJCXrmVy19SsqLrYztSbRdnOE9tlyFFEYsCV8sdl9vGSqBG4h9gAOr
Hpx0KjFfB9CZQqSMVCvxEpYvZ7lw22UFGTsd5h/lhqYIDo8tvJFXKgH34p3y3jbxDqEwYSyVfBmN
J9AXBVzlqqJoavzA1OXWN5qyniv4u8Q6FAgaAG0J2KCSM+Eaivs9rWTpiKZtXp1N9XtLUzERDC6u
zlKlui8xafKBRsMnsbslpWl84oQGQa3UPMM+aQ6GGF/UdH7PNrrd3NaHoOWLrudsGPCUvSxYSNqk
H7oMzwzQ8a1DnmOcUM89S05TgHXL4BvXhzbanWW3rbDGzafZWl1eShX1ZeGxWi6/y56PKxvL+AVY
augPwgENZ4429crA2aPnz4qIsavKFf0gcxnlKTLP2VUTuIrHhuVnqHorCABUuNIkdwE6L0fr247Q
pPUg3H0KhpVbazTT6iORTwX6+v9RHY4Ud/fqvUiRhHZrPaprJ4t6os2Ty5tffSnAZ+P6VC8WVOb+
slBDVaCK2Fd7KGvOkh5zIbCrkPyfOnR6S+vtVN69nED/0+0BV2qB/mJjiAOji50XsqezkSbbtIrh
dxpz7n1UQzPnyunwUobRk9F45OHUqaJGQd8aH1Ztcy37qNBix7VUqmZH6meTX3J6Xp3dX1A3MPf2
gT2asvpao0l7doOAK3Ctczd3DIwOcpMi0G2TqzFLRJBkEZzTxtgsXTY5svZzJdjKKiU72Y9wlnBJ
qRqALPKs/gtcU+YT6Q54mnkoOVuIonrGfWiEQ1LRDvay5k+kcTK/+NIPWGEJr0SELrGSY/0Nslxm
hev6HBBXDvAs7LLiYBnga2itOWjeBHf9ZttfrtyeSqMYDsRtZilGyc31pdYEG48bDnOQho8f0QLE
igJxRS7aHPPoVXc4lBgZfnn/EXj0IEbEA69FUScqmh4q4qU4+v1bQ2EMDdWfFfWJB8AEMN/g5x34
0eslq30mGUG1JTypw4AqyXBbQqheICtainZbxEhi1tBr332LJ8nNY9j+1AgMYqHCO+P5jc+mBq48
qkQAcvJfW0kkzKqP3WkpYEoaZlFUz99EdWC4dBpxZQQKwCkxqgEnP8VhSZnpkaZWvgdDu2MxhSbH
XnKP1NR/3dTpYGx0ZEWvo3peYQvtcvftLCivscCKqHntRXgNYecHQhPFp/j0mx/yweP6Ta1pyoyb
d+4CC0+NhvUcpH2yrVvwnMw/heNSllpJ5+IcnsUUSp0DLxWCN7h2Q+rx8aLDmZ6YfI+3aeAoc64J
RY0Gv4vZrQKc+loTVJAu+noPnABKXsAI/iLwmxFjqgPUDlqBRHRloLztxbR38+SicFKQo13+Djep
PcLwJCAsy6EE44KfFXUhiBKPMERR4WowtLTvvT6x87uRLaDbcompLEf5yOyr6FN18jJdLzehXb4s
gYBuMhfan4QTSIZryMnA765pVaL3shzfDp1oPws0DNzK5dGsBU1Ap2PedGDW5yxTKWRXUiV++PZA
w1iCsyU/vc1icKROKTvESDoEk8DeqViVDcUC1gkaUVtiGBdwlKVqHTjy9/ACGGiwoRumnJYN9RDB
WLAzFTFh38dFOkOw6olIp2wsidMyBAdm4bsdYIpKv94AUa0oDg174ieqFw6jnZurahGV/cJ7/kxn
uWAfc6koeXoZPqU5nqW+Jw95HDgM8nDrRxtothITrl6zbOIkmjxbL692PrrX1Ufm3KxdcZAEXDHE
PfCoQhGt05WyQYn6L7rV5oE2eDVp84CGovHjnJ+PRcLiBMH5N45h5JtIzZxY/s/jfaSdhFrUqbdK
2ugkj0GioWa9SuPCMVfxlza8UuVwWBYfe9f5keHXcRaNJ5suxS0uycfBFCShZnqOyqi643e8RMS+
nsm+LKD+GJvm7kn0JIUa9ztI1UT4L/KALFAUwqab+/Y34ww9g/x1KK3r5KOiXBivfjXg+wd2o8Mk
jVEEyJ8y+Dbi86J+djRb+RFurvanFIhaPyG4ljXx/+vLMOQ8pnia0bbK8eUHmGR21/Q7FiljJ/xS
TMhIVm+0JtFvAcZsiLHplFvbqZIjQy3MrQX15okWi7yPoih/iPhhmllUk3Kh8G5xZkuGonHQwmhf
TUSaQ0IRLczv0MwdPHYqkBS5DhTCk7eRXQgDMOV5GFYvPJ1lh/ZtlHW4yZVpc1DQfHkHvFizpA/l
V0aQsanVAGLoLjoGgA6rP9JO8zzn8t2GIdQWhAjOkJfQE2Izmaoxb/6TtzzhBHwQ+2xqRqkcmw6q
U1TMEQ2Q/iESZsVmiPGp/jd3xWv92qbNwptWP+oFsKX6CjnBToae26sVOuAq1BdvkG40hnZ40nf8
m0gYJYKs55FOsYdmx5wT7Umgk9N7eUDZ3xcTuti76LeLCS4rCvm8t4bifqqK4pMXYVpvNmhmoFEG
mBXNecStgZfXwXMpbDR7PNhTB6JfnZXXpBZ/yd5cmASPyaliqtTksNjR6iksCMhBXRKmLaiM6DLM
zL+r5lkq6sshX279Pkz9BwzX63i5YOq2HqpAce1Xuq0+r5+JL/MN7pG1Pb8I/Y4NQARu1j5Ku9rv
itF7gaeqOv85Re5e6EDHZrPESwAwveFeD/94isOotTJhoGkGbjxkrbZPkPwlrD4XCcaLESiUiLPa
60yydsvAcd+x2CSp89Jp+lNQ76lXZ+AtNwOxIYiDhMl7BIqXzfnBCLyyTfGQ5TtkjOvasIGZzvd5
1fJcpsQpWdM/q9JL2sOotjEKfb2MdHE2QVLD4djxc0UTHw2td530QXrrzuXX2WbKKc0dKMzEfaDI
JMV5N+vu+pwaCdKl+M+7g2mV5+9alw/Y8i7KygDBPLPiH7NS4Fhs8Vy2nvFg8SSDy9TnbM045Hij
VdQGeEt08aHXlR9jDv7QbAH41sSx6nkFaTleqONRhcbqfC+PuILv1TcJPSSruc5G1tNY4odnI+tV
bn3ZoO+eAZei/L8jYGxI4Xn88BI2ikV0Y9uEJKigkeAsF/FjDD0vnFkrGV954BFJjsKb990ZM6rQ
KwBo25kD9K6EogdO8jv8zhwI9L/SHdgwcshdE9oonj+jXTKIJRRo2KFlbmSB9EN8TCXn0wp97tso
1cEZ4nPIW2WkL0gNZ0DB56Ngm1regEW69rdIli82Z6OW6xceqqmjHbp9CClUIXxr1C1vHboh95Gv
mCR20H4EKLO0zQ8L9Sh9Qc0Iztnpy6seOI+Pd3rfnByUxAQKWucqcSIoOePBAXuSc3slwAN00n8F
IuiifxRlkhXqf0w4ASCxrAPE4VSDntMMPXGv9Vo4QhuOt+9zGmFjjTQ/raoqtQYFxromTSDj1X7e
9A4jRI5MMjNoN7h/fgLcnjBVNwLIU5x68NG2K1nGGiNNe85nCnq3gU/UmoUlhWTEScY5t1U7HNeV
ZaNwk+GXb2uLrw7BsRwtq3jN5zJHM/M1SsXzEoyafBt46ledJA1jTcJa1R07cWZW44WEMVZx+/hT
hLCsE1vanN/A9McZZ/DJ7Jb+pPdoCC3FwCMJUP6a2gNYY4enNd6ohEcBULBMVRkWO/likhVXCkJv
1FY8+L1RAhUNpcGEVRM7NhpvLWS7q0jd74bs1ncAztpCdKwOiKVe41DbpXr2zL47YNM2gNPBdaEn
PQCL1VW7EFEsMiWzuVvxYMi2+7ZiEuzzgQh1uhe/eJJNq9JoLBfNqRz18zRVG8/JzW4ruOn4Jh0j
ph3HyvCmDQdvLLTe//RtDX1Gz+q5qAlYx+XKVNVsVBQrS1DBhq4sYH6d7kLgjCv0EiA3LSBb26rV
OxqTj8orc5oM0Pqapm6uw0H2Vg0N5urtaTLPc/nGM8wTZYajoT+SdQRbn8jfYXtoaNuU48qU+JJG
HQEKETOW0GkNUJvz6be1Z864GbGkCr80W8CFGg==
`protect end_protected
