`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4256)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAM4ZaB6gj7rLX26j3rNRVytNjfb3RE4+9gC0QNwSNkS1y/DfxVETNIRy
2lUPI4kx/RJaoiP4YMMMwjHmv3Fpa+4WOr7B46T4rGdcepNhqiC/ADVfnVw9RUk87yebzF3synvS
qKOwmFLBuhxZzgBueJP8mVxkHB1Emr/dnpQZTO8yH+ZbSkU+Qlb6T51f1RcFF4v8Vw6rLB2zql+r
TxHlgzaStswGCGT7cQIEsAmKr/BVFCOLbm9U22IutysGTTBeOgmW+7eKMwaezlrNERWu0NtO7fnr
x/A7mvbvfrLYBKQLZTHzD3xtzEgQWUORxJBM+VX5n/15ScI9+dCHJ/RwugAQovLEec11xgjXkCNd
zOtdfC4qQH6PLaZatNZrgO8PnKgDlQBRgUi0EZZNj+PTbIHEv9wNyMiiZK7cmz13Fp4dvCnFjcDM
R+e2d49z5O7ywbr7EMagQ9edvutyqQOzSlO4isY8tkeKyzDqbDtnN+6BPEoymq7PtDGcx4Uqag3g
9iIq/t7iDOY1/PNiSE6JD37WSU5TI4Z1UyjJfBF6wEz5AF7SxVeBJZaK7bEH8bnNRDPX1aTGEEDV
J+FSN6S99ZKLnjfReWNUpsKXD9GWomdX56s5ZTbQ4yObt7sS2p5j6tLLDvoIibQH2kR29nRo+iEH
YYkOWWTcmLS0kdLUinPbO9Xkoql3BX/G2bymzklwsOO8mHUL+P1AFqueRLmoAZ6VIyULVLgAWU+F
BmfcNzaaUE0tL23Iy0ILITvGDKc7PQKHKxa/CdI1JEYXSaiNSkb7K9MLxiLe9nv0nE1H9wUYgK3S
QIRzg8Xx+nlQHR49Li7ydpjuvspUHysKy0cjbNEz1Y7PB14Xk84NSho0T78poFc+dFFUPAxKcnpM
W/gbjNzlo0yzJpnTDnWK2LXWpdr0QwYT/Ugb9yLfzPI7XXisn+xHsvbjiBkpIATWPo20VRQHG8bf
Toif6JtqF5FS7R9pGvd5k5C7BNtk5uhJpa4SCBOEknYZV/Try89WudyduXk8LHFJWClnRfqMvZXR
ZbXqzxB9Z8hMRk6lJ7hapmeu1gF6+jIy47MtG1OXeayxwQnl7MVXNJ3ANdjTv/6VdVTGpvhZ2gCw
NjXEtZF4BMLviBafWPapF4CZnCWMCF55c+4JpTghnCI8rajWArgz38oOhgAOLJzRw4mGilwn06Rk
z7MsPzGHYOt3b+Yj+cSFvr2Z9kpqUdQLaP99Beqb4/LX0KQtn8gDNvwWDofZ7TUORpmotky0+AfV
I9eO7wdyM1hI5OxtMUXjS4SnKbG8e7zkxjFhCaF+JGr0z2gIPwddvhH3TdAcvzcVbNJS7598JsBt
evBH7Y8SBpc0PY/DW2t7IfhmSsUZ6xqE+GpU7YzCexkCxn1Pt8A82MV+oFtSrsfamd3vw4X0lfjB
rFApAiTb1um5w89FoIrlZ7n9qJsRhd0x+dTWvzNeNxm7ZqCGoh8nrsJ+FUfd3Ns/D5oAQ0qaTLg6
HDbVeFVLQu649+iUrWaNBN4eAwWvuveUZQHC84hwidj56vDEk7WEYWmig/wloRyC1J67GbKZuCm1
80BIq3WRpFhQTCVVBzQodiEHq3pv/tEWSpaqJEQjixMblHiBw5wJo99v7vtzM0zQZD1Tmzuh5ian
JJS6rHJcj/K71qK8f3dvhvSYVF9eBf3A/zHOUzZM4tISlr1FJWlAgLhbyRpfsIxZpy1wsQf4uEba
2y4ZO0NDoyup7uoc2r3oW/nS9gqp++b0Ei9c1U/eG7wp8WuIgmOM60eTXvQLCZ5Gtc6UXqNJCLrj
T1mffrP/WSQHjyHPggl4ZCFV42OzI4ETH3/jEqpyIm64yGd4e1cRf8ibQjqCmndOkDvKE5fQFIw3
q2HLxshp3UhxY/Urw2OVlZZubXs1LMp4Ou38s2zNT9FsLtj71Iuc+UmFIA1AvuwSANTUUsxBzq81
filq3oYg0zm/3HY3qlb4mqpFQC3H26j40Rwdevbonl8IdbwCDLkX7RreyuVzgHzuIlxCyy30WL9A
HOXflrW7qYIupxLcNqHPISm4MWISwMHJLZhELgech3xcrDEkR5tfGSXsRcnugQbjHuLWwDglwMQu
qd0Yv35264Ca0Yw4SqRkxEeB+MBDE7d12cqFPnk0tGb4bdaLbDmDKBgjJEXkEot7IgewtsC0Se+7
aP0IHFSt3SLoHAohhfakYHYN6sYWJIalIYIaHY1eNHgv5lrxkMrHCiIY/Us9w+IzSiIsiX+GjclC
B4K04ugl2IyhhASgxx8yDzFcq/VHUj4KWZ6tiv5IbtsEo0pLG9dnz4moHlsho11NLqLMjOq89oio
mDmAoE8h+hKP7h1cVqNxRbyb06EF+rFvsBrZZFaVwdXAgnyfMH/c5joz6nHXAvRUGGrQyiX/q7bP
XoA/uMcScVcXH3I2S8JMo3V+ZeC2g1LY7h6RiM012ttv5wmWQJjQT2Yu64BBv5xDDMOeP4QDN4/i
wmQPb610pgLxHmR5UBs+gkEKDdsyg3fZXCvRlZM+kipya1QUOezjcMsEDUuCpx5iZmPeVnMW2qBA
d1js8Jfg1VhZMTN28XR/fkykb4SjzmMH+Mg55/ai4y+/dM4NSRyOfX8mlJxLuuEPbp9KD2zp8c0n
TCYj6eqESMD5zC1B6QEnkpbelhqyxhCwSbMIEmK4wBEBV08511kWXWQrhPr7cy7CTCDzQpDihhvB
EPFqs7jeR14bhfgjR0NtQwWKaKukIyE2AGbhxwFat813/RQAmJ02fgT9Oz7EZ8vZ5MDdwnNB/1bu
a2Ze3/+n721LYsHc8avRU3wFb7qY8bBJvh1Jt/4/tCPOBPVAKaBIrlFXUZpPvhAWTNjwog/YI0zb
TSbteUq72oJugyMtQKtugaWoYVad3y8MnuW4fED26tMSlzkkgwaL7IbqatS+EwDpTy661MW647ho
JcgyWV/asyFzVl5PzA51X+gIJAS8oydpYrp9eopsPBDZ78D6Lo15mCLIc6emk8ZWEqo5ez/KeA9K
4MH+6so4OmcJf4JzI2aiKJJTJlQiZMp0kn6higb8bdkEzkEqIJ2Eq+qBghfVP82YsfIETern67wk
/EuLrpwqZs3/peKDBD6ANDARRDbLLYrBujA4LIYztKjdqtVATOJ+UJEQ/eHA9kYqkN0Qy3UydqCO
+mRiRLrhNKOXhEnNlVaKJi2CkQdfBGWvzC/ihIxzUsfAuyAox6Nh2XO9DZGCJFmemPNcGEqYn/jH
S06NHf9etGE/IXscZSMNV0YDm98oKjAgDH+XYF3uDVymwwllXHo2xw5lRui8Yox0NI0C7B5Cu0T4
c6czyXDVtiWREJMCMV58Qy4VMIk4oxkG7VyBZA3t9vFr5u6T8pYNp+H1RRx42/aQHkoMNOO6rBlt
Kyy+XMn2ji6m+a0VCLjR3etOxPu9udP34atSjT7N/aCOtaYyQpizb3k6sSSFpwFACa/2kgDkrgyr
+tTX2IFkqmuZN5jOypeqAMvtuFYlmZXXEoosF8jOBcF4Fzg0+LCOWUsmX31n+dC2elJgJtzVjj9A
ZmnebE13dUzd28kLCZCkhIbhs+HaNU88SdFQkcfV2/JF4oKBz8rb4yJhZcu722CmYxxpNxdS6hU4
JYSB0gF19NRX+EErvxSbH768jHYYoHN1IQc0Thwl95ilwmFFrIa8ubSUeZ6DRRCdAzSttqVOAN84
/XvsAlEvfcthWpLR7qLeCNJnRn9GBiKCu+56GST25pBCP2mZ5YqJMGZxpyM01Qgf+9TcYnvkw4hb
cMYkIACjBUbIu8U0a/nOBvDr51pZZivu+M0zg0x9WLnzu/XLYtYbUFD2Wgwnynhqzg+zzcg4q57z
Cb32kIMRlZokrjqBmN4J87/XvncYGfWLF6xYGoL4eDIyAXBMN8tZP5pJ6KAEhx94sEy3Ztp0aQwl
/qzLob97I4RqjE/iYqGyBOlz3G7E431HOIc1wcst3YrkWOO0XGVUgs9KFMWiKQ7kifvO8G3sPKQ6
g9DKzYeWI63UzWJCsCKW0/VtD6kt4Kx123JWab8wMV+SF3E12bWPFYFh6P5ReEQqNF5BQAmhF8aF
PWDgO6oe8XZ0877y3l4g9byHRGQfYV5vwtuyFLVKRaxY5D8qxCveTrKfmAAs2dGTGaZrg7VKtEEe
n72F935xvHTxUe4AaaMMsG/79BeiHGIaDMZ0DInCJf+fh7JcnG6cgrJfonLC6/rFWldcELrqfhIM
ttfj3IM0SdQOkrrjibmiN/9odQMx4TulrF2l5XOwJnv5ySx/PdKQD14D36pffm5RQadJosmOU/GJ
BT65N0szIpEJ4Y+W9BaABkuo8lJGqWPMKeax798Ze/m/+A6sngSMveKIidGLdHUq30rnMGIl0+W6
hA0Z2nMKpr67aOgs/pZBrVk0tEzYGZwVxW6p8ydqrstCKdPOwYen7u0cSgJeuownvCFdnqiBq0Ss
dYuxP+okJ5A6mcyBaP21lnpjNxn0iwyEz0xabX/lQAWXH3eL4W2xquLAozqo+THC9WyQ2Wlsysk6
DmHVAVM6mPpLTPpGnS4qzt7w/LDjMIiiY82qSsyrD5iArLL436o3gDz+jxfvdP+6ui+ZmPNhMpAo
q7jSDs7hb7qU987XNvhThKV6Ue64scOC74iZY0aqQcRr3If2CajQ1nBHK4kOz0jVxzRZzbt36y4N
UGG1QsPmSQCsRbiBQkeSPxehpB+jRaMAwuLeBbr331n0c+yBBJtCmfMGsTff5EqGZLFg+KI/CKf5
HVn44u2Si/SO/PvDlmQ9rPzH1coq8bhotQ/fqBSIJHQ+ls0zRB/LzUoU4X7jgldxLPzRlXfDaAQQ
W9ix2Yud8s85I9E+uJsFPuDbo8xIBEGzgoT1OfvcUFJ2GzJzXZUoJFiDKp7MvMdcIgLKhkDJdo5I
f3eiLwcUl2cm59fjEpX3hBk5ufu2eViP+vCyir+vUy4ft9Ipz+Ai9cFHl2NmNeiyNrxye3Fzc8rd
XzsuIWUE7bjoMweRuVD0RaEVgFWTunSDzO4LAHF08GvRSf/Vo8RFQcEfI0X9gtlsSQYxtTen4cIb
+rKDt6IHPgpXs5zp5bwGgHeG/AbhpOnOyIHq8W+OzOyz4Nwt+am4Nn/xrzCKbd92wHN5vDDf/tJ4
U8queJlgzeQDKpfX+NdTqjy7AOX+VgfJxtaxBC6SnS/O9gQ23MkHVGdaHnTW6/3G9gfNvPp5oCMY
RXt22QZK7oHetIibwUqEcPwlBVPhd2vuYUICQxMKnF1joo2JeJ5TMqBmOcm99RK43B0VEB3BR5ef
mdHjHXjfyio0PIochHwmb90sfae/VCVawozOqNE2CDXyY9sT2k74dt0G2yhF6oHzAeEYvNj9V0on
eEJ/6C4nxBKSxgO5UfyY9fX3uf/xKxm6DjdyM2QeuaKF+9JX2ivcei3jggX3RM+k8UjUDX4yCP4W
2il9fEfOQEp5Rz7o+H5qnKiQKf7AInU4fVosJ+chiYIuV48OwK7brGUUco/ACv7aA4ZBFZ5sm9Ay
yHGBN82FxbbWRfoaNqD+UAGAeK4pwBG7xbtF4Wx+qTausPtcoHrtKZ0T2qHeyKteQeRW6KYDajpR
gUVCgzYw3pPjTE3MlOkXHUI2qHmpvZzZyhqqW26i8GHKrUOiMMo=
`protect end_protected
