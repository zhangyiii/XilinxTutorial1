`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
d5VJXu82JfSwswDjhvbEU9He9tQ5/1Rw+4/2nB84LUuT0wfekcnbAADJNd0/JtXdeaCUlOw7Zwks
Bp1VvQeB3w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T1a12gH9+o/WCd/uq6lAozrIbwFwnflilDyEA/rZKRAxvRmKOSqBXtjVpxVSoEgX9El2BLPK+36k
Vd8y/iFx5HcwlteYeuYuGTvgQerRA9ycH4Qwt9s5DC83MaSGod9ecMMI8PPrmdJ+hCOX8sXwEsN9
IHAKBa7h08XDRsgW0os=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZE3CBd8eugZohbo93EvXvQkUxCnosHfYT2eG0uuvFgW4E1aUdxFin2hcHpeAodvxBTyPhYz4Lsqw
3nsUxnz9hTb8Lhj5XnlqKx2mVFP8Z35n8lJk21C09QHBGoSukklDPI8dbQUv/KxN+k1qsLBHfCBA
FWz2UAwKlgCaoOPe87s5MUwwDM1/P/D4+XgEQCRDz/7JDN7p8ZFVtltMEx51xjJOCvfGoEeTzG2k
908lkYgt+B4pvwsuFOHwC28xicC9lqwuIR+OiqTI+hvqIl3tijnK9dhEHXmlIo9PqdVp3p9K5niF
C0wKwI1gK4zk+Z+Qv31AV2g5KDXjXxSpUgHlpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1K/c2Exmx3hO4tktdfNX/hsUCqBDw6bH/vDRPja11f/SX2mhefMgy+yYp/XXIVeJlyTPI7AwLQ+m
jPsm9qUsxInkPzY00BDkxz+XjPmDvPZhWK1LaTfp3S2KuDInJ2AYP1AwgClVQtpRFpipBFYqQeNS
QrfV5V8iPYsCh6rtCZ0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z2R2Fz5uoP9gCKKJ4H8ByaZdL0II83JUVbmmEiqboGhJOssYqqghHZS4Xla1DO6PE/W7lUbFZBMN
taobe7WZ5vLL3z9KT5znQ5u/8vqZfQZBnNTCM9ij+NRl3PRmkUPrtcd6xURukGspBspXFvJDNTq6
HoC8rJF2dAK3E2hXtQ2qzFXYx2JspRBZw2ARE4ENjzYZSYK5AhF3nV89pEvyjDlChnkSNr7Ec2sz
zSK49rQXLtbokqxvvzCHRCEs+NoMqKlklN93OyjJFAIzYffS6GiGtNeycU755Cv+/fAQynybNWn5
4vdHnb+JcudvHzAJFK7/azTzKOJrOSm9uJYTZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8496)
`protect data_block
mvi3i3MBI7n8zvuunOT1BL4eDGhQlMnzDOzVrYI8XHOS3ZoKFTTDP4UmKkCCDyXvukS63/BOGJv3
NoJdfMFYhDx7pjz50AatTRm5dOIAKktHZJVnSGt5h4GNaEO2RZrMb78Xxh3U1zVrxlZ3qI2EnKT7
5LM1QOPzTANUpnUwZMrtssno8rTmgtUmBnkLkQzwqhjsnlkHGDdcTSQSED1SISsOycOAvCGsRB22
x5ukanfw5DKmUkfi4j68Mpci1SuG+kCh/xm1odcqCvaQG3qvz7ql0dAaTFvPffizNvJuY0JCm/u4
w7ZiemC6bnWGAYfhmL0Ia8wdLj6tr9vYVAbRhFnFN758s4yCH7fwkhbV8z8fpTPzUsfZDEp6lTwH
RRilf4f83MNDPE9KavDU3ZAOuXIWIVehxQnWgbhVNOE8Bj7KJElUA6p1hS10VmCKtKJbSkI0L5d2
/hJWC98Q8adUr+LSgRtVcPrv0iCUrbnjPWp2SK5N1TriuWI8FdZRrHfuyuTb7ZnGbwaul7CbmOWC
tabyA8E85BJuJBlZQwhz6oZCE+8XMyG+4tADK/k3wJ0p3QTSjs3Uy/p+NboSKvN3F14j0W0Q26ZA
NCMnW75YUTdpg/oIeMmPevG0M1ic84GmsSu6atj8EPrEtuHemDv9SeFblV6HggCV/TtuWEz+aUGE
YQcu/AVEbx3ZNLdXxSDs903E4xsvzqAZSZjBDDtriIrJxXEZpA7aHW3oMWgEBpV9lkxoxsoRvB9t
6JYxtyhGpivOHpKuic++lM14IjpJJJD1uzR6T+D6wTTdF0WfUYk5OiNqFp7Ncbapr/MLdiVYSw4d
AqcdZ7tpKWvcYelJX79SJD+uiUybxTKKY0D/FdRjn/JBWU4aashoecEoG7FkgFyB65nFqSLurCWD
c3VBmugIVloTNw4dRIgNx5IYF2mXl9GjwvwmLbJ0V8wyo4M3qw1Blx6MeXZydnifW+Krb9dqZyMp
lw9DF/LyD1kVW65AFdsWn7VS0iMdN9Bh15mEH0GSAIbNmAzUQpV2MA0q3OFnv37yDPKbV6pygTX0
3zTl+XXHLuqNyydQrNnZsRZZEaqQM7l6oHI25pbnVvd9WEen8uBPASWvYc2o+hDN6wk4urGvqXJS
9of3gK4QDJFGu0XaE9cfZO7JgfzuWJPyPZ6NJMEmCMjuPweA2vLalZDeAlaGHpj9IlvGCQQDTz97
oxSmTiPjqmFO4EPnx10EKU9794lujosZfW8O6/kCCplKL0ypepo3IDgjExNzAAUwAC5AS+8fJqYJ
Nn5XkZ0ovijhR8z09XM4nu23YOQ1W7FwjR70FGDuNobUI+wMxdKrd+IB9x4/PjhL6VveJrmKmA+4
fYQcxEuut0DNMMaCLtwjzrlNVQ+r6HaGmfHrV9YmZ4y8DdwUBFhAYvC/hvrzZtIgCcL01hH0GA/9
G+1os2KriJl2P6Q8tEGUDISIl8qD9L5M5ggxE5tUx66WTLPWSihAlKQ3lYkLOj5oeeN1DkxrpBv5
fx098bQyMf04HG/HuUJGcb4yoE5I9ECMoZBFvyhiC/H5eP116e6o3iHs/LQiKR7Q83jgaFXE4v6A
2SBML+ElPjQ0WmpbM+ko31avFQNAJJ0N1bSD2zvI1gqTzmJc5RYU6UDGIfEVkfkV2ZOspgP5armz
ai9+kNPzdanns5W3YTCAuWNVsrtMD6mN6gfFKXn5TbOITwXA6Ze++5gYnffDvH6aBCvTUZ9A7uDe
lcAxwZdEKwMRndyVZp8yRMkFEYog9MJRJpLUSZUaeZMFILdTICvZEm1lyqa3pkq/NLdwkm31ZUX4
cFE5kZ995+aH1B1UiH7/H+GQzJcyxsphENJmEgURLXd+JotW437UZ4lvgB2a5hQmN6i+6Us3FBOk
hJzhjG7/lNsG1+91OoBrWfUR7oEZaxEXNyVWHXHQuznqz3Jv2+71PKPZ/JPoFsI7p86xvgi52pNR
z+m9ynxZJokZMqaBO2oXkc5SNEx63mrDDdI2JPJD4YW5R3b15eiS1c/AHVtHT7WIHepy02iJhLxy
pIq428ccHcwu/tJkxBw3cOL04NkqsoEtfe4tHxLe5oCI4dDfi6Y1Gfnilh0LtjDHkMHijLffeGJ4
qkDhHLhYp9ZFTViE12w2beXbkS3gcc5oBtmGCG7Hk6S6RB3YIgguwsfc9WNL6YE6J+ocBxaThcV+
5ug8BB6/yA4Pl3wyylx6m/Oil9Rge77hWr2FxTe6h+WWq9dyzrCN6VXFKf9bYHsuCF8U93QIPiuZ
HNAB4VUX0fjpn653EJPsvMCFywgNL24aw8RSxa1QShKY5d2d5nOQk24LBslY5WQ8ifypHqT5TTY9
6a2N+LFZ87PK/1oEUs+L1tr+HzduBoGucLmpBXL1G47SvqCFmaUZzhuUW5fq3Dt+F9K17yS05Irt
cqpBuWgd0D8SLkPKaBI23iaRodRr04gwJkE43qD4QvrtMeOAMYmGW0gX3R3L959l1X25lN5QsO5b
cvm0ZVHMAs9cnReTJRYsZr2T2UC5ZLiLTRQuSenoyZRq+VtJoEe6tq8KKj4tOtqM0j4oiLRG3d/z
bxrtP5eDHPl+t7YbzaVpBabQAdvfYhh0tySmC9/zo4nnG6pqszTHqhQr8dZCqOLnSSknXVD+bCcV
PBQkh71TESSgc/ERCw39zUx0PU4toFDHgRua0/fLKapXzryHaybYhgnqVzEg6KKvayQ0L7HODtiL
D1sbxv+Sx57g3TkURoI+0BqkMfVots7lngXM3sjqPxiRZMlzX02GcQeW8cnU1ldhDHWhTPlgh7/3
JkSBai9wZSDorylQ+Y/wQYjnUMm/zb2IoHAz97taHOM7cA7W2bS+csuMMWHYDbdsq+WaMf9Zxlgu
GLiulx0kL56fkE8GJqZeNPmYarcmSIEhADS0py4aYojjYoQNwtNzocWgCu7PTT4/C8fjI2LjCpLw
20tSwMFOShwJsMKTiJX2j7NEH150HNUKJoyaF7Z8penkNZOnagSmwK59BFvBt7mL6Q9oqnYfftfs
7ZaJYjJaxwaIaaotXGxd6PZsB98E3XX80X+KVjW0YJY9ugp7Fyd186Fs0m5Xb+qcCEq5Qump4jI/
aIgExGXWq7znE1lGoncTaWFtWR3m/LF9YepN+ntEx0uc6uJl3tD97xIvT+TTIl9C4YzFguGoE/+K
4zjUfziwFZxmToTHpPw9b+l5tFxzAZStZt6mnUyfX5prsWqwBkEFICDPGyzOxEcKNBrE93FChmpO
catW1x4yyF8uC1Ao0w0Xbh2LVcfXLD1swHuD54JNfjEwDM2+7XGmP+uxgl+EBJfWzRaIyAHRWKbZ
6mtRf5YgofHh7vJo4dtD+ixDKnwsXvTN0H8T8C42yoi4AE20J//CcwDSnhLWIStF0Ob5ChBAMG+W
T2+pp/p5PYFew/0B1rX0vK+hs2t2x9mApwkmnFDT7GFjgLeDGyVUus8wTUNX9DPG22ETikXr2ERO
hxKeh9jugXFDzZhxjfHkoLRMobH6Ll0gjWloWkppAdGeFa9quv1M9wE2QE3gBOkCwbCbCiWkHOb5
VTgW+wcOYAfnRfkstLeDXqvhCTbn8LWMqXC7+iQr4onaylbHnNm8zANZzxxZNueZ9Rs8+Vm63lxv
xaYQfMW/sIU16XN4g68tSzvHgBYOYfoyKf5/GtmtFmNhOtgUWvcgyye6TXgdmt7ZGpMW8UV1rmTn
W6ZsiTSKBca+G0+cgLhcAxy821+q2usGVzTE7HR5eHgjuYBiZdG7Bb9nXhjZzxM00IMwEHg7DFp7
Ef+adnnMFFQttAPTXxKaHjPkJo+KBePBcYI6M69ELtsLcgCQCvYsMmSsvqsPojKhxtZicgCaJEDg
mhPYXVHPvlEgG0ZpV/68ZyRh50a6qPtqGzgGRPjbCamaZYnfBNT/eSGgxgZyYuk3wsGGWSNnbi8a
Ra5LQ6Mwsl0arloS8o4hg35X5bFJUMkJxPGAwIY05s6pNOS5QAZhY3d3ZcKWbTm/9GcAqmD4psJ7
cbmwUAurMz4Zv/htmYhd8WsOHuye4SGCIHYBwONQ9Y6CRlfTQzUSRXZ5UMADgrrw3Q7xr30lxEQe
H0UpyGrdHstEsyTLdCFm2s18WZK06yJKd9Z2FfCQSgr/TTbEwdH77KuAg58tXBmxoCvqEOuYhU32
Mi18wzHmaDDW5GTHgcjmxX8D5hgZrhBMu54LC5xDRMtkmtCvqDYU+fzgj1Yc+14woDCn8lJyGaOr
cvr9tWugUbxFYNGo2YccNOPakysVPt+NtA1ybyYO/YEPqceVnU1GH97fVN1Q8vimT2if/TutlpKX
IsFcHAw96cY3ZAYalSUekAJydNrD2KpbNBi4AserjKgyutqPb8dPgx+hQjEi707/ZNF20oJ7QSsD
RV/SSqfTeqIMxKrUNKYtplrkVK/QnmQ18t8KZSNati1Gok7WEtW5BTNYTKMh/tA2XrSq5DLqtYyB
vECtAOfABqZ5pMTmv33aQfY2aF8iWpp3ik6bsytoBYYcFzcHfLBHyHx/A1ZEB10eV5Ts09sAyk1U
v9UVglvmiwVMGJxQniF/ot8jo4dJqFr7TCh3OBYMUs6ZoLl8gzLBOHEgkEDVu6BZuS+Hr/bEfK6z
oFYs4DdAMrdYjjlBXvGlWwdxJQLLAAfPuw/1D+K8fnleWnBlcHEYa8ApM7R+/ROMAjd1dxmMAHQi
FLiDhZY6e7UxAw5A8wVgnJRHR4qY7Hs1DNMV7Fqpwsh6FfvM0jcC4PcEMTOFKU8H1fr22bqORUBs
6fKhxi84/kWqHQRf+KjwMW2OF5L4UZOIzJuxE7MKaspb3WedQnqMhjXttdpBfd/5YW0+oCJBOKww
KJskLStICXsfbum7bEyxPRvgJsLEKUUozF+6ThnAs3oC4hHN+7b21ceDKRrABMXhDV7gqyz3cPU3
Pc/wr7rg7gD+KKTwhSqEQyTFSOZhvIdN27APw1DLyHjU/MfJbF+1IJImtMx0KBpsuCIgOIksqWDC
JG1sM97UbAVqj4I2raxyirDFGWDfBvAejvL9r5NCOBPArkMuRqkLJeK2PsMUeTxxqyz7iFRfsQ1u
6NM3mleXZYAmp3NpQzBZVicYE/OoX/1a/0YnR4b7G9Gt1fgO4ZsiMQzncKPfuAhiMwWVrswiZV57
O38MhQbRF132Qz39ClXysdTkQ8ESxCWIznX7nEVU2Yc0LzyfklPRADz35io/zY6EvratF/TuTCMu
ydYm60WmS7llHiSWYgmkfOLO+Lq6/N63ewPdXWcq/wdYJwpsf9uEO2TzAQhc2MrruHMiuUlIgjZV
XsSzNTYclgy9Ke+PxB9vHH5DjIwEA8Fb/4+DwOMdN9XmZKq6rWvWwd0PhGwGbw8jWKMOyDIuy1mG
TQsn1jlY+eFTa6zNBvcgPZ4klbDy3Lak9krXxYgcAUkzK6Gj2g20NuA/rr4B735coMGhJG95H56f
zULe5I/DzB1lsM6I1PuN5ihvC7SqCxK6aK5l4CRm0iIeBLytaUjGrgO2CELB6ejxJHMBs8jEAHzK
9dCooJBWVrXqwl3U5ev15f1Ig3yboMoplk1CDB8oplrEWD4pJqPped+OJy5fvUcoX/fgMuHEv59s
TEZ3FW7fw6bNDdzjCMFY3GB6oz7hqKArNKAr0yKSA++2q/PhUoH/kBqyeQbFHWAQORekdxb4r9+5
XxnB+78OiwQ2yQ7RJRwQR1Pf6xkL7QlbXZpRtvE3H58lKaEd3HFsoSvfF1Oz2mP4cMpYXHadrz9S
fY9530Yz8jcXKX9G1/Q1VBg52p+BRcy3ySIyP6ScPgYudms7W5Ui4VLc6nl2tGos1PzjHNZFyuuv
5uCfv3+hcA5mY+iCdQzp8n6wSPGsIQKmqjAvPM/U5webcv44h8nydtYw7tua/CieLHtxH/pxlaJl
5NY+jk/BTBYai4DenKhcBAam9We0NV0ndYw50VmL1HkafLS2sl3zkRJxZ16D6UuWfX5x0TossxuW
q5pmCBKNAzDDBCnnj1wnEFWSE55KD+5ExVHLL7ZOzPNFM/rEPMH99RZDQcIQUwrjA5tmC3rblUAF
4XZdi4DfG9e7RQIPrn9R8Y672+I64oejIOrr4jgA/ilLKaIGPU5CsHL8NqOQbHSiAn0LvoUrIDag
ZaT1eWkWsl6seeP/tK5AsW/yCDqCNhQaYhwuXhbYb4caAkwLXeWwKZ7BW4F9nBKKBMF2tchjl8eW
tgOyippF2ual0F7v3MtppWyh+aFjXzauKCVNiugBtUnwqMPMS17orZ9hnoRJ/w6uCmYYCcoHBt86
E68acqDjgHoDTvcqJ2rkTBFF5AW/+iP2r4GsqGnZfPqzLT+8fpH5oL4pA8042tuHuPvIbKAoEWSP
AmqSQAxE5+/iBsiQSBKXlpE5u2ik0+VVqRO/FpFGgCgB851/67qOs2hqcdKtlPr64uEFq5b02gWy
Nu8DxWoC3yogWRNQzsdP0cEEp1obFhXA87yOx8Jo82AHtQMDkYLPBXESj/9/23/EtBr/a98GJGMG
fLs4K01qmtMCIK9bfQJqnI6VYC2QmZ9hswF9hGXJIXW0eLqzeEZgT3ICu2/+aY8DlNdo8R4prUZS
LoMspfCuiF07WQXQf8i3V+NiBJCXytVoPPaKVyceUXhd6RDI9aEmJ30k6At3xwujfsYNrBhOUThs
47mFgqb47LPyoGYs2kGwmpsVz1n14eSJeR4Yr0tcUzdfbsy3298PAe75w+p+4+2KDhP38SZCVw6a
iOnML+luPCEKgcUV3PP/NYKX+iKT2IGBQv7GGiVG5ALq1WYZv+mqcvmqeoj3rBK7cptZnIT2pmRw
raCYTHVblOSnsM1mzseeqQRN9Q/ShbG/SnikOH90LVibs93TtKKrLsvS8VmSulU61j95tYWexq2L
DXS85AD64iNShbZInHTEB7QgS66uSPnmmrGt63C2EEFvDMzo5OGOnFJMdDra3cg6VoDqNJB/ouaI
JfT7bBZ8h/wHyMTdvIdNT6qAWhXOoFeopfyEqD42kzdotqjm9VAJogTS/JtFxLbbZ6Hm/IuGlHrl
kExwpFX7QgGFkwiDw5uzzsB9GPMO6I9j9H0W5BWHR1lLUzxyAsSGeROXgC0OBAknrHeLQftsG6b/
6NbSucMVp6eJlAUagTEOksb8jlwbUDA6VwZBqoSji29+eGZxg4iATE3SKRqtBwDu+pQo9aTLahe6
E2XS05jUGMMc6FCuThmDn0z43R97ArMmlSgwrY9inMCsuv5BOpOVnbSHK+UYVzfznWAUD72bjXnK
iHXsJ24pHV7FYfKfzlVeeAh2v8vpiwojwp+J2l/DWyQ6y2kGWN1ncyHyZ9kduOS1FS+j1N2im8lo
0Nxkc/oqa7CtzXarhSVT57VZLQ1ceFpz2kWE+Yn3KfqUeiMNq4LNpUkTAN/QAIQnkG/AGQSlPeyT
Lfzuh/9LbD+NxQcC58MaLP1oacOiJ3GLXk0zmtLOWtfbQAdbtoNF2JMxQklTsPKmp5QvSxB3lC9O
atLj7Rwo4TxSmiU9v1StnHyHJrLiz/kunK9JeVxNBLv+m99gRage3c29knI/RWMmbUiVmqw8x7zu
+ndpeI8Do0zgRcL6Wxhf+srxjSpcvOrXmRRs8S+2xuDMbeZZtYTEt43+Zap5XkAdY+QPiKq/XTPz
wF77OLEtdmK8e8tVjhaPPQbbSjMVJ1pbEi3E+u6IBfwYs5ISLFfF+U5Y/kmdaj2FLFPAHuMxQEbA
WU1nIRdG+1yifcpOIivQ/zfj9KSWdwnKp3qKG4KACEBaEdayGUQq5fwgAMk15pmc7Kn282uZrmAj
ZkxxFjXJYMeKvzsUnd7+5DJGqYhtFVYbxW4xJ8cARfA7h8eqf51QxQjXEVs+cpa572x7GgfIVSuV
GeO9gHGuajv5ksCwsp//oiHMO0rllloD0qvcV94NiBzHGhDxby7RtHr0avzRGVYDHTLblDaR+SJk
Rpx/Om4ueusYlZabmzTD0ZkKE09NSkqGqU/nEBdGS2b9kfwUPqZOH803xqIlTnKXm7mkObDg0SS8
YQUShFUXrqS/z+5UCktqLDnnJWv9hm7kcHcvhtx6Ci/9IscFG5UsektTfXmuR0U+66PjoBDVbiIR
ZuQeJx2df9xbyOan2GbvQJ6ak5xxO0d4Bq7h+rFfYTZpz+4jT550y/VUs1FwNbay4oNOo5GFjIrY
T1M2Qr24PhoSvzERa0LgUl+BkYQkjf8uaiV2alBBkdlXFTr2HawdUjfh9xqPpOnOsokQoH8gIL7N
+on1H0WZ02gnxcVF/baRvP+GnuHJYXb3SiLB/PAdOZ0tp+Jkm7aF7cVSPDuFa6T2qfmOLdZhk1wG
WYnb6fYd2Pdz/lJANet6DqWhqJfHUmjTAVGhtaDi3gcnZlAcGaz2qnqosgIUol/ywUia781hlCpT
RafOVbGCF/q+s1Jfet6OFgQiIXDhsiqhXbrU78g9i347xg6JXIKgWYU77BGdjtApWsiZaNnwKjGf
JZAu/tUC7OEfz6QxgIOgKkkLlfu2Ub8lqRom6vy22RfFg7FwVIWUFyLSqmU91Cly3kYymJE5PXo/
xLUKzSQL/9Wp0vQIa8fxaZMMrNkfp5snTzUzX9gT4j9WGvbazpr7QMXJH6f66nRQfrDhcnCDVQFw
RGmT37Fc0nFbWvebfiWKxP28IE3cp/c9YIhU5nqjIWAYOOb91VCoiuq14sXDuYC3i2aZVi6CSiPj
9JUx0IojIU3KQwm90N8DrA+GVKiI1xUbQcNkmZORki8AL86xI7tAZnbs4LegCd5A1WGKOHmT5L6G
MTJ4RQ1jISodyR2Yfj2abcRUHDqIdf7iJqUaGpe5Su8Vz6eO755tjHCvto6FjqtYUsu8NlN537W6
DfiFIPl+UPz8zqlZshHr3olBjAYZ1wOZI0LJ6cOSxgcHoS0RsOq9M1p2CioGtAURfDVV5Ibqeyp6
LXhz7mBwF94sdin9qswEClzpWwr6fHKAJLqWmyimYkb/zJ6/unAyNf1rc32dLHbMDmv4ek4fyQ5V
YMpP8Ra+cq7kTCca1VNZMnIPauJXrrtHdBFuH9HqIrzynAiertzg1gc9XL26/sW77q9Q7N18id83
LpApESB/HAjyglUerXKi8wvy/iPvMn35h5lZtAg+hBtySD98L65CFEsb2YvvXqWrusEGJJd0UHRK
xvUXeterPrzguJT6VpkWPQP69ASH2Ot4AkystMR6+pjb1dzgfJ+iQmgijtPsTuxmcN8eJKB6tZnP
rZjH2MpUJLawwoTTjHIX1Gl5dlCbbydupIQRM8s/i7XfFX0JBACd6WO44jU02V8uCzIHcbkTjUDe
IpsxSlyRbKlX8lO4RImqKKhquCcVA4oWCWC2JvRE2ENxvIlQVJRlejP//l7R9ks545GKzKlG4Lc0
DyHyWjZbucXdvVdZ8Q/xqXjGi7MA4FKP7zE+ihds3pBIAQ5OkMq/ldkCRW6dJTFN/6rUVrQrWsOl
H24fAwGKMUulbaXbLpa4vJIyPOazTRl7C5fd2ve8R8QFzzBbzt7eW1v5Puv+n8lJFprye5XfSdg6
mOn9cvHPDZIIcXl/qSfrHetSWxMin4OW+eogF5gIwPOFqaoBcpa3NSYv3NJYzmEyKO3eppHJ4qBp
s4gfMn+CWR6eoSAa1mXyU65PZIELjKTt1Rc3LQGJBmmpEqHOjrJj+lySQ/8II12pNXWn2xMRSzrV
wGC1nLnHwEb1IWFX0Qrw0nSBElsardhKqHPWK5oYt1YUdHTAXbgwvMqwQdrVJ+lxJkGdtmLfY+DZ
uECa1RjpOPDqo8HfVy2MbuFYq8/W8zHRli0Ultx+Ka0lP8qDSYgGCSmkTG5YduTusvW3zwntlT8I
fulmplVDtyI5a6zK6kCjq7F7p595mkcXJsnV3cYFaaBJAAyioikSxJRYmzlr9X0O7lnoQHW1KuhN
JigyJuNiJiSPPZrPKOYYOZfM8cLOuumpPY/2M9MwfigKWoZsvAvzi5usKyTBhFyKCcteMDCT8gnm
XYVYO6JxXCOg2lY9LPwnKXyMKVv0LCy5lduVtDq++i3K7cg/+gwv7QlbOPHhQ1SEsBTcJRCEwMrt
UpBURLbhnNNpFRcoL2xEul7qo2pDM2CUv2IP6gSnqMJbWsjm+vrFYhoYDHlllVdybFWnmnocEeP7
YR43nlHLLXYs0MqYBvjxyLt++WvHWjoi4/VHw9S+eOuDnJeRJhe02PYyV8l8A2mgkyXbwgC9Mygn
xNQrtmW8EG4IRF4Jo5ThWF7oP4YOI+FeA7JBazGjbuEXWCxmFkQ7sEv+TlNLfUIrgI9NXnTBBiW9
XTF1moVa11XAo2d3fZqt4QEbb7GdXcCySz5yiAlnir6z0PIUHVqD0rdxoONFMLxOnrKyXck7DST9
QouwXIPAz4NJKHLbTwIWi5r/x8IsTkjxnnTM+msng7rioGBoT7IwnZTlVe5lkWiT7pFG1TUx29N8
J9pzEv5B1004l4bMSNrcA6xotitbMLwtZogpKvduRgDExMuzBno+WJVSqXEKbCE+/FJsNR0Dw63q
Z0s8LLASJfaTUpwIhZSYDy8/w6spq5845kYYqImbwBxDRKB28Mpz+LaE5FjMd7/4N/femGfxrJHK
7/BfnZnUcskiKQp3M1FTPn3YPMBaFgaPNCtmtlTFNIM1tkwnsmpYiXFDPPZDFs4Z5NkjEPDmN5Eo
ibxAvcXtClWGP+QwEtg2d4b0i8ywNalP23+Dr6L9poO2aaQlt6aJjHKLgQLol8ZNU+bDXUIBJ42D
XmAJRPzVR1WL7t5oEe43acVnV9Sloanbu2d+QmHI2ltv18rHwS59STYUTcYrcbjwY5m8AEbVMC3z
fo7UxkxXvTx2x7nuBVdTuPVXorSrs3O0qbF41yoUnL16dFYOqaDaoZdb+tY8EwbtM/JDz7sogcXJ
bLW1KB9kEWZtAjBmE0nBZ69xHE2DSOcDrXP6CytCgBj+DAh6pQgHKWYpTPBnkPfiR9lZpRzpqMw3
6IPcxwkGwjjsrLnNiCWzPVly+skVtWwtbRWpOPAwPYE7B99pNmLBJOA037zS7Cek+hkElCZhBdtJ
Ou4gZiWTrUUW6GbdILoYoptrb8wmm/5+Z/hV13IA6Idw49+mqdSxYgKNzSmADiR8qB6bsCmkA5vx
Q1SYVlv8qikDKOJAE2lJD/Gvo7TkBBZ5Bc7PZ4vwz/Rphku96c9ilJpg9LRm0qK6GECtDA2rFBEP
Dyj8Nrd5qJOJHWqDFUJV/rGVaydAuWJdNbXLseuegn+1ETrYQO8DK+JS9cWwd0DZNNrLUQ0RPvQK
k1ps
`protect end_protected
