`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZT7+RCzMGpoBYSuObDu7GHIWP4wbG2z0+NZPy5ctMvSzcpDtYTeVa9Rt2jwWGft47o5EJP3ckUaz
ga/PA8jA7w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nez6Bl347nb6+rwYEAGUgNCAGAzNmFU5MeAC9+3K2UzYt8qxPFrJ/SFJLhvmq05ak2WdPG0DC6DY
KQm2he2dsLt5QsRiFYmj2xAL1KdqCGiHsVFY+u/PuU8GEcfn2GTMt2pBI+06udHlKRy3Gt2+icT+
Rzwp56VKG96Z/MuGTf4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bJ23shOZkE3PVggRHLeGJ2PbG8xrPMkBPZCJ8ZYfdCaWhZ4ZYd1C1zb43X+ojqULL2oHyUgAMgSj
ecIJtiACC+HQhYS9ZAedcNObDtyg4oslk+vfdk+TM2FZF2Etrw/yAEbq1f/PH0Kn+mbNEo33Zwe5
Rm8FZ1wDWOyOXh016tcp0RwCvdj2XR1Kw/zAigz9XUFsy0aJtcUXIJIlKcvvsjSATgFtlJhxEDo0
pnsWRjWP0UYdXkfmSQNXFz8qVRQRGSAtue/7tEuKBK7i+2io/Fn8ReAkkGJiWskeE9nOr9dx+4DE
9tfPWFjj0ZgyCy6JPKhTrEZyje87nH/0x9mcFA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dilSTjuujT5h2DrLDbS/v0rUBHgSqc1odhqH2k0dTfIZcb7N2jGBdTrXFekiehlmoGDjU9sGGdlh
yFg/bT9j8pTdVb3lIkuOyMiLP0CoFYVl1z2IegKN7b9yFR+7EZbxn0N/B1ycLjS4ssnQq+SGbWl2
k2N7LLrQtkLu5td7xjU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pVPXt9t5C8qS/9IP6M6Y37REfDMW0SGfG45oP1DNSuCggimX25Htte0JNMgNJo8ar+6qTjWsopD4
IXOQzxTzbzczkdAIs6+pl9RpNOeJpa0bvybm+uwfWb8+Rcnz3NLflVxnmjLM1ayKKYARNVh7gQb9
C4SQt1FdooQ2JWlTXbp3V2aZpvw5F49u06L9Z5ayEEDdOQE/HQgnVfIryQKYB8stQTSh++L7A6Hi
fnnwsPjJQ2SynIHMSopYLmrhF02KU9HJ3WVKZ+nUrhCKV9djJvyWE9gZFn3X/nfyIkmo23lpYTgC
rYvCI0W4K/uiiwV05xGsCFhMYz37LiZv5/YMUw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
6Wo5rjfCVuPcU2g0iGcqP34p7s/KuW0ZmynWdo0NUbOe4m5I6UBm71JQObfl/N6HjzN68KxyjRys
HLuzYukGLhGfq3UEw+t5b7pMc2rhR0IH90OaOAAiYGMweA38XFIpQhPcHhs0cVr3GFS0XYGSc3yh
or1whPAdpaQazv5yLS8+5gci+luVwTVmIf3Krwh26Rh05uyNgwe8ynSuoCU0c4WLAZ+RWVeKNEzm
OOeKAxcZpTV+lLxPWyGrRsYSZ8k7SxGXM7DuzDdEzgMcUjyoRC9sGXsPogug7MF4KQwJafLk8VDa
d1Qu9WVkLrSSCgbggvExvceM2pCZXIWjV+kwdV0j5bAvso/TliOoiI5xAp7JcRWM/JiQtwzxUZEm
va4xXNxG448awXsYWIxrQUmQ/K44fcKcGvEsOt6ICbBpNcbp+r1OTKW1ogaDznO/b/us7kSJ5L3G
QqcBCkd0rhEMsDnXrIhbluW/mPi7sTJ1cWVWoK05Jmo1jF4/zRj3CW5BTkmlCHGW6OD4s+PXyDcu
8PxQBnkcCS5DwT2xTtJW+fs7KUhPDSnTxrj5riRe0QxRyHSQXqv+Cub7CGtIyevl/T2TrNmQM7J+
f26dNpmahLlg0joGoPsPa2Qgiulc0RWBN58krNCXVIZRp3L8A+qHVcgih3jL0iH2NOn8VqnaodQL
hRT6uOIyVz1Pbt5aCGiu1Irs8HgF9EOBmORWTkuL42m1yAK/uSvdQuUNDam3K3Syf8e42mTLNkuD
P7Rdkl1BDeNAcfn2SC4jJUatfLrssFm49KA8SXHdm8hdpTvEnX/Awsu5Qfvmr8/lr+UFUvfbq+E0
nIYKpD3b5qbKsYim+N16hqrf1d6X3hyqCN4kYQygPNXu5paUUREg3PJGiss9iYEpV5/RUWKoSRDO
lZ1dPb+DTcpxkLvvpyZqxlddNJh+lh0LyC1aPkizYVoM4ESXeKF9DnVK+plMG4pzi/1owMqlIbmY
n+lI6YQ8QuvY+B6eGqVcaIHTt9AZ+DK4NQdZg3dKZd6ypx6MU1xNB+uUij4Z+d5Njl1SY6ir1ALv
NFyVdmbb2Q5Nao5/XQtSF9SSXnLlsrA09q1Z2BeLWnRxxoy5KKnXnh6Yxsh19HSyB94nSGu9xEa5
XC3fHF1uYufLeuSaz0iZr6TZubkA0doK+mVjUVUAORvDNUIxEmTi7RwVZeWWBqstpWHssrnwa2+H
9MPzHUfllPLaQMUzKCW5PqByAE7s3cW3FvYMaElO1dBvCk0ug9GIsG7cUpunhxplxZv23yn2Bks7
dITkVdvpzxr9uRovzt8LjO4SzYELbTAL2M5zyx93v2aGrjDWaHcGCCtMsQOJh6biQiLA02v0PbJ5
rm234J9DtGN28nam2/0br4f793LXor7eXiQO4pLAAVq2g0ytUfS9ZI98HivaUv8reHaYKTN4IC9Z
lU/92PGdNtnci9CYr4l+IY7GbYi4cj/I4DVBvi6cLjJgbxIG42mXmXs59a64EkQQkzoUc/udsnOu
7hqS+E4jNEMFr2ywZwF+7KHA2hT2AGIX32WVlzMsTNWcYAjdDF4jcV+hW89BnF2gLme6Lgrt3U3N
/5wJn4NBMT8cezvUjLtsboueIdTmNvrDljqWTPfjGwK1PWd1edpVFAoivDDpqulzd3cPeGJYVZtv
gfL5QTR/f8FfZheQJNB6p8IZ/8N4dl4uClBQoCbsCnmJK58uxXftfUIuvYZbIjqzY1ErX2JeD5vn
M3sNvrCWvQ7NsRDBOccgVzgTN2M99VyKdbsLUo8sa4W4MdJoRmeF5WaK1BBDhyvvftUj77SKWX0g
AiblIpJcLA4VvJJ+8nlCIOBqp7Ur6n+/KDDwNBSHNY8I0g4Nj3l9bv1qy6ae/ySnpkA9bVY65cah
00tsJTpMlYCm7V3f/t6Ef2QBr5NNHuojF8of0Y52eZxtwbOwZqttcN4ApbFM6UsOr21WnSuNgb4a
drjBR66jbLGT9owm42vOBvt1Lt06phlpoUy82bXgs0h4dPftjOM4YeXEBigzw5m2cLcrEmwm+tWP
xiPdkfgnoeEHiKjhLoFhkUyIj/FMA+X+nztfjqSdjS0c5NRhhjKGHsseI3tqeADnSWbHNEctTWiq
8xVGK6w5yATLBF1twJ6HaYe/Yv9o/gJpquy1Vb4Q3nDTwp8/YEawyzEisovf8ivBbWf2qOB6xZAU
E/fJBdciF918MCoF8UriJnBkYW8r/N+VeDidUUcZhfNMhSXzuElOcI7n77MYCvky7o94hlEaAxI9
evU9MZFawta75eTDJWmIil8L8D0J8FsViE9YqqGXghthvt9xHCMuxVN506rmGh1t41DjZ293S48n
GD8+cH/+69t1eXEZAS5phZjFlZO7p33NSO0J6QH8J529d65Ih0mK6bawkWbg2IwDgzIxI8lY0R1H
szgIz/e1YzGZr+iSXs1QCK50eSMtOXLzOZyb8tGDXVK1OuNhieJFJk0MfTtiUOdsw3QsWLKc0P5A
qIEdHpkRpIgXM3AVlaaA0FxOTDRwFOBgMyNO8Cm+0yds5fjvoBzfE6g1qihoQr7s/Tw1TIYfi0oU
1ygl+T70J4rJ991QV+IWvzE58sDQbmbiFv+CpBAMJSzsgxY9QkOXUc6PbmT/QF3dbw2KMHtbXGIV
Tf2nEHgYJeKcAShIeMITe8fCJn4bP0zek/sQjsiL88zXUU2izGxbL2h5UpBQPFHrAqegiSZTMTO/
Bp83hn4NqAEdbsj5Sx1MdNSKXZNz6YEZZlRv5VTBS+2LlnP0MIvPqiZIjuGzXfFST8le+9FEjm+g
wAMjrkMtjYG2WCuHtQaJvBgiMK2ptenKFC9R/BMRMyDERjA/F9qHlYLRC+kKtksKR1PTlJOHPLcM
Q6mehMToE2oXoeA3MhNQhj2OSagBe4+tMMXL3i7cqoiZXTASsXwXrPLZRqdMP1poL3QabkB4F3KA
katYM5K0RBpaRePw17ZrZR4I71SNAdLfU61ET+BfLDXFChmGSKCQ+ahW5tcablnjWVGRXDjBi7Ko
BaGQCuWxE5MOja4F9D6NmmeM8MwmRRSXUBIxD8lvdqoQNr9F6/mxmVbNfoytQz20+MIl+ntBBxrS
BfkIaC8vO42GrepbBAlfwQyuSnvOxPP5CWAg9HeC2Ati74ryY5w6KXyqxw/+CvMhRT81MDwuJ9ay
l7JHg9URXqlImzKVCTTX8iAyA3h67OrEt2V2Q2rZHjcyqxQWDfdPfw1ZudfINbbW1LQO9yw9lQqJ
VhExrmhd2B57RR9DosdS1QXZcU6NfrTY9EyNmWGUdHn0E/eWkEYs0/kSybCZ7cmOwida0CP6u0jB
dxYuak0HC13d1Br+6WdEoYWNBfyyrka270VeKK5zchHjEPxaVgYVhMKZ+yYP9SBqjo781oAyR1Ga
F1GXEkH8OFKTvu5WKXXNVbQ9pgFG2h2JC/Ugk7vrnn5Zr0q2iU0MRIdF5mLy+ZvCKKInvDpHCier
pbKIKgDaBfDJ8DnqlI0rsyb+sWBemzNIZ4Je/crrH69s+G+uj3bdmLHyEMhaKhcGoEU157Wd5bh8
Eod2GmLSbF1FCegRhQrMYXBnzNfm26IrwoVDTnBldFPMEgtD2+MoOPx+VKEcXFjKMTrxL6jkKTSt
zEkuEwXT9f1K+bsViuCDasl57kgk1ZH08Lor8AGzabU9DI+TmMl9iqmBT1nOf0bINKYvl+yKOXVl
VNLtHCsuSIDmwCRaItL0z2CGGneELTNeEwctoua1FAeRHC0O8p68SzXJfHa4VkdKvrak6kBJnvGX
SVgZSU0rqEtk4lVnLV2liLWHktxUcRZ9Ezfb8X3twCZamd4/9BfjubpN4jOIn9OrspuqR8458qPu
bqyKCU8oAEwcplCn99fDuP1NhZpEaTxRL5LqzXvvBKDFep4ya2v6oaBcOEXcuq2L2/hsEjjbGR0O
WYA3EOcMDUHgNMm8ow6MnhmDCdRmo1Uf02eP4+mV6iAEZo7B1C37ePRYsUGlnsXWNXR7Q2onTH7M
TX5kg6rkwW/SRCu+/XsPujPnywThYndJhYqOK9EQj9wfnxvTiA+tdtgxKnNkPIiB0WORrobFGEyj
iLbHR2KZKQ4/K9sez9FOcYpTzaEvxkuo7//TZ4vIawsZ7omMz94beo1TpsxZDZrsHnw607yjcjMR
3cbmlzY9PB3lGxgs7/zRg2fQYegkR4g/JYpmS/Ns3DUS2Jyb9tiNgIJgCAwRUpsVd24GlrbXLUP4
GJgqrT1wHLKJst8EE731QmIZ7JKVFuERnd0RMbEBJWk8ucrmoq8qVtaOOeMCfpQ1ouc1cO76W7Vz
dJKKr51wvas4h4BE4GeUx928xB+As7FW3Au5/haJI060PrZZmhfrdonnEXkXxZaZ/hgx7AGJblmW
XMyQA4fDzbRUej6PLjMfis0pxb/kqc4t1OYbEMDjGpYMnobx6rtSsG4FxHzE3MIB0zy/bCyZtbEo
40GPn6bZQ92a/0qHVfV9LNFiL6gtHzUPIrMD9LXVbwasLYpFqJS+GU9ZXujoezjQQnnBqTwUUi/I
8eEaGu+bzJ0GJy9kZW3nVUro7RbACQWUAaPUTdbmIKYh0VdLXa3gef0eRvYI8gD/Yt9A0GoeVX+l
qQDFBuq4l/TzMb5JU8I9Sjo4fcDsebbOz3kbi1tJFRKy4F6t1srrXwI9MggzLs2yTTQgoG8duWay
nlAv/UCJtb3nZJLMugJCwKiX0yl9J1hJ/SSiu85EPwU4aru3CNwYRuraovasuansaBkbJBN9mD70
nQmkc58J+Qj/mk/dASGgAQvfDOV1WLtTWE/+AvRLZXHoj2tjd4Yx9RxxwWEcBox0Ax9ja++RTiCT
xhVmL2kPl58Xu72+B9TNyg==
`protect end_protected
