`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jg7ZSB2xI/J/jQikm8Zlko862zAjpKBGuPSRLj2TaHEWC5rTzr3rFiYHZX6yv0DYk/Y584dxn1Aj
ZJ3fEMF2Eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J8XF87MjtG6MD92nYNEuYX3aIPS/zAQYepXrxQuouCoZ7DifIM+PcGRYhyHbT1c+x8wNqIyddvPX
H9E20LneyNoZup9aJc0KklSHkCBi4RFSlJYfEHGi7VuQ4DoNHay9ZZOx7KnkG5nTkuG8dZKhL494
1mvb9OIoIew9S5frQi8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FESqZcf5Kd2nw6uez2DBxPYJSBV8lpPPNkL9mii7n9rOA23QnwFT4gzsX2GnAKh0RRoHvqDgwQe2
oriJIgtSnO9GoEYt557lwN4pjAIARzzVKmQozG4a0ZADHcAuh9dE9U2pgm4IYqaA0WHemsJP3RdH
ZWLIA5hjsrEEni35ostJyYxky5xMLNN1/n6HMS0umCbRhs8srgz/a5uvWD7FFpEZ2a0utgDi9MEX
Ot7P9GN3AM5Ug4guXH512IazlVntMqLUCdCGexOO2NqFhGpAvwGxJCtx5XjHjmGW+9m1bqRxt0uC
W0qg1W0dWBjrERQ1cn2SGOV3FZ9QqHCbH1eBSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sBWw2a997MC11UDckC6eUhzOMD6OyRi9hIrFSmKM1LtA+EoEe9hBOU+xWnNJxZwh5q/2lTaLVnRD
SOXNd1eh6E6oJtNfyy/eD/u9oSEqrtEAnNkzfHKZvGwMHsKFUk23bSYe/H7pvyiU6gwLB/zQXKRM
aU3uU6qaXWsFaGyQrek=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I+E3SG6eIVl+eQQNtE5uT75GDZk2w8MwukclTFsLuB0JtjwI9/9l+wqqevSEAZVNako39sma+Yy+
6sWVRLVPo7PjKtoO7mmywH+p7yQSorsf+a3ZiNjDaYRK+f9GNaE4daxPW5KbJ1GJwaVjbrTJXjms
6KviB77YrfOEwKiKJnAPEYDYIIKzPfz0pkPKCCTKaUXpj+fFxyjC7bycPwfKU244d5RTVzX4xHcW
KE2Pbl2/gBhqu0EO5W1xcfaXIFlrwR2GLFrc0Upm7pO12jbH3NSKac9EirjKD5ICy3GjrAPQM9pC
bmcrUujXKJAoYdm46Fb/QQhF+yxNF515651OtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43760)
`protect data_block
iXdONubG+SYUpFk1+3xjbTmoWUUth5YI3Atb1aEXZ+saXE5+BGO3fPH5sUZBPpBGvC0XNFvrYkWj
mKjKwY2xZcfJ/srndO8S7QOgA1cW3PGqqy5cSeqaNkpdKKv7LRMKRcNvzOG7grs/8lZMh3KNjoyD
IXsq0a+K7fwBVl18ZhYAY1e7ftc76HaRu/8rLjkxtE7Q2J9eFQSb2UtdMq6Y5VOj0vNMKtDPUUYQ
EapXijfXVqWDBMqI1nbHZOALvVCnYVQJDo2a2eEbg3LVp46PYehYmYWBNiTcT3fHf3km70lpX855
2eitSDl3fEbcoRRSxZE8Dd7GRlHBulzhkWO51Y2JKAmruWiveSfX9qxrc1J2+ns2jpzRnDbHsJzR
mH6NXg52JAzAA2Iz+0RIzyDWsYKD72UiQfEHpRNd9zHdKNpsy5rckzxGpo5ZuSYG6SC6j0QggC42
BJezzIXT+wIKKThjvv/jI1a+/VFfCYD6pzU8fCBBf3oPvXVjNKWzN4ebtRMisdR09CkJ7AOSj3Pd
t+iY+xsCZyQMM/TsdHfYDJNhZuohAtxFnA9wChQWflGRB6Xf99BhlN6gsevu9Hr8ffemU6tQxCXp
rjcOEw+TOB8t2UHDkKPFVkCX6RW8bY0bJkEA2KeuvZgVvITl4aGa60P30nSo3QN5B7/9A4lFBWlu
QmQMJhHAcrEvnKCP/tZfZ7vZ5wxObBFAuFyVU70IKOrfleKtR4AQyBlEkpvjSt+/Pj8XNxQqmGZs
QVMY2S/gjOopI3ABRCZ1ux1W7nBo1PhN0z3/H7vQ+Aq0KMICc2nwmi5CHXHoKqMjtpIsOgGc7KQx
qDmdEisg74KxHdljo3AgbXt2QR6T4gRkxfbMeome3wR/CNOPsgtcgA+cf32xZowz+agqZFwewTbg
lRzkz9HjLaktc9fzU8hWulUb4BmvF6NbHdzwMTLvW/kiQ1SWAZKD0Cmev1paj9/qI1VjQPX8+N0t
T+rFShPQAhSjB0QBqJ2iAh9TXJC2h8m0Imrxd5Y3uYWZ9EG2V0xi3GmbV9eww3963quXADHbLjUq
bCJ9488udjpodX5wvVH9sA9qSVYkj5LxCbqyKWZnvMJb+a7Dyr/Fy7QFb1ZgGOc+wTraAMDjVW4Z
VHvkaMkffzSZgFd+e7qvKzbslE0akMh3hKMgbdJgUCfBIggqz8xFmkLyPYpeOMvdr6RBqpHxiWbq
FJqrh6nyL95e84cUBdQiXCftgqZ/8fcZcq1skHoFa1Ps50vf3+Or24AO177LHyvNTMT/fwQA9Lgv
QS7/QbjAprc5BTPCuTgxVtRVYf5PJ+GUyazrkPR2s8XTfiU5I9YS0qmbgfeJdBXXTWQckffoIlAP
uFLKUeHB/hlwM/j09wvNrRKku7E5gnl32njgOZ7aHvgeYdOG9od5Crty2NZEOjNelmlzRkdj4gY7
nfKxWdEKov7h73KbN0EyTdQUVHBKCtWkHlA7QD3fTyXMcGC1Aa27S+jlvscd33xXE7jaSjq18dhB
d/nfFyi/oPWbeIx+xORSMpEce6wExHVXWRLD5p9Gqq9PLuiZjDojo1nAESmqiKph1EhvkjDNwi5a
WdnMGpdPyWZBi+TLiJdGK3vXbhfk/G+i7NDP9XfayHcfDrD/zd/C0sRs8FAB7UDF4ogo33PMPoXi
sq0MS910zI8M+8y545bkRIAg7TriOS680W5IxstqwdBAe7rZydTEsdo+gfiH5Nx1j6lpZJfNXwlM
UrbsuzUbEblYbLM6DegYq0kc9QBvuZdpN2kOfSDO71GZEWChUCvd5noiHGHlT2Qp29X9OLdgDBQn
APSNFip0ky155cne9+++iaR+x6UgpfrXE5tQq3YYHASfYdjSehuNsv0Pbg37gugk8rtMw9GTngdE
x3FNzOkfQQdEL1jt3gVprcZaJx2KcMGiAA7lgpdqpETO5t9fZzvH4rf8+NXKA9thE4iXXU6mS65U
krgb6pvJMLtvTPB5W85h0lEmPgKF3j0uwcfUgw9bVFnJ02R3clrAt8OUHUi0WuIV9D4yJuSmfbLU
zhlMV/Ur9J+A9XSNVlFBHLXrxzjnC/T98TLVguHiuv3ybmWqMk53VNE6b7HQDE+yve2V1EusTrNQ
2XaHxO/OIxs4AmM19xRFFfGROI2gpcvPfKGNAza7pwZJegt4QgBUv0vhZ5mKzq6mMrL1AeHeycCB
BaQW/kaZ+fT/JB1DWiXWsxLP3dJsZVxfJzvVD6nGx7sUqTpehC3LF/F/8Yzu3A2vNWyJvJQKeQwk
OntCFxdPgS5CnlaOOmADPf79Hc4P/OvBbuGbosmcbv3oGhcfqWe86/saZ3qTbsqF2LvQchhWT145
CFDMCk7ZhYxzG+gbinPMBf1dd9M5lTMrQ/qDk3uayyDZtBmfNp/SQltYX1WSBbGhNKrzNi3ejf3t
EO2dqcABPSX8rMTSNq17A8CvwnS0OQgiK5N5tMu6duupNjFrMZJtI2wOfHeZcGh4nk1CSJSb8Osi
YNNTyOEW92VQoiNQ7QTkyymi5xpzexvSdEeLx1/OVwHg+ZEsH4qTJxKsP1XPTESHAbvgeJfoQCLz
KeBZmZvF6lkjJjl8q12IJiBT96RbQF+XCOl4L4GRxSbXEi3U9iwO3vF8n0gurtGyhVQHXYaQ1/gR
92+RFCDYn5R+3gju65E0Yd7C3onh5f4uoSQaDv2O+vPSCfN1yCf/yUXZi5oK747SsqbOi3HhiWS4
lvQIDLVwDlKalIotk+itTv6ay0ewx1B95/bteGq2VZLUIEl6iykbH6lHK2mEByNEhTWxLrxLTY68
lS/35K3Y5ULcdNJyKdNUYx2n/QKT++1yG/PNDVGKkNnlQr/bW2vteZCqJqEJCvvlILvshrqoYPeF
2mK3a/HB3/XwlGs1k81GfI4fjgaiz7xQ1vecjhOApvXYIp5KOiqJBj4YUiuIe3DnhdKloRjjb459
PTVvyPHOIfKlJBXO+VwlpA7gkg7zfbR5IngA/zrtDheQiqQGH9VPA/K3AyFpcOluykd1yb+w92B1
WcH1zsyjSKEtcF3I2DqlULUBXDzUiSlMJUgTDmMbo3sdxhWQdIBkjuWGQkWU1TfiKjwY8sswcsqE
ZgLB1gya0thXgI+2+8tSr09byOQeFxZgeo9FysDysXa4t7y6kMUGSlAHhomJ1sAK05g8R7gN3LbG
uZed+J3NttniZeoChTgtEFM/eqkjY04Bcfh9qsJEt7IFZbnn6phXGj14BuSwtQ7emAwxbZn4nHCw
PQsHTZtH18ZAUDSWXc0x+0Uj5uDpWRrDEgOETaSRaZChjzWqT/ajoDMPGG+hikjzOidPt9/lPj9T
dTGyAcBuniXNpJcSKD8Dd1iUEW8HdP7KB1wAtRfcSOprthf7kv6hbTXRAAjV0qMSw1hWCFZbEUjr
AG9J5Tb9wC6/CcLEB6uU3ttYEhDtn5JtVOBQetD8XIBCAIKKe+68SPCIsvjd6y+XkIhj57F8XWFd
rY8j4ewJ4GSsFXtHHyW1LZdibppHRDXmld545P7qmvK/rdOyjM9vhSB2w3O39zRWlo4u288p0gXH
PHv6HeN/nPzKqeQ6ujigaYFBuq8VofQPA0ySNB9SnD6V0pPMqrlca71YhRId2+VRN/dlPylcjm1U
YG2Coj47u8dJ0zkGjYiWKx94HCCvzvruWLCyEh49owr26lk7nzO5nFOJ3S+uyzD6xtaBGX2JTe6k
Qc05xZgWSefkOWKva2QpABG7wrXcwWGLk/dewjUhcBfpoYRWdzBWk2kscAW08wBTINxUNIRhZbyp
KIs1GW7UU2+LHtb6k2uIkDCw7KWbvrB+xm974rAYaTuTGkEJeBlpdqODNmK+T2rYDC9A/AunL2+N
v3OHz2ORHLuopWy76PrTtpghyfKQMJShiMIHAxyoF0pnx6AWH0Pt+WHQ6ibFtbAlJ3OzoM77Z8WX
u/Io1uRu2Ye2FkdK0Pbwf4hmJCVOe/mqp9gm93FALMYdLCA3yTAogsFWQmwj3I60ayizVB+o1lKJ
tGFtQO+8FH6ynQSw0gXwFrEWCS1/vWbgUIk34NnX7IDyULpdyVYlcDsbxG3QPgEm4bAvkubSkrnT
GMTxZxqoINrNPP3yCBv6mpt2uMuY9n1281iEsmbCVvyZJpHvtBSXLH3h26wCQYgKn7KbKEv5u2UC
hQlX6R3Hmx0KTWNsJG2ZydiRhA6NyctpIIZIyZe3szIv0AdQdsWN2fIwxP1rxZE1Ipvdr6btM8q8
WnY5XuG2FPY9c1eCxJAOAqaBRP7o7pkA/lgMgXPZcm4MCs9W89m0Ab/GRFU3FWZH4kO7NLzg8oG6
vmG/A2MNYd9OSPTI8i9yXadwKL2cjpKaZPH/ueVFJiZZIYFZMt3+p4b9r/V8XWuort41eFfxmOkV
+iHw+o8qzcSX8GAXiMGT16k3LDa4de59GoIVILv+rFmOpyj8vz70FtLBOHrs00+li/uLqfklTI30
TE8Be6583AXGkg5QP9jCHgJAYOm89UljXiZ1Y2cSAQyE/fAQtH6oHcz+2VweFSBWgPtaQuEZp/mu
CACiS4/rTeQacO2Zpw03w5i/QGPCXBJn2ZoMkAuOLG65e31eAR/u4rHjtVtNOzWJeNTTazprgs2L
7wt/AbyE9NTPNS4kgdvuN5Asq6gqJAZKK9+u9yg5uykPI7RF0PbEUOfxVC3bKPQTBNxF4bKdNyW+
2bEIvuZ1jSeiOoGDYH4UDFq5v5ta2VE3nwXG8BkdmvQtuqjzmJVgT0LX01WMw4xVntqbTDr1shlc
QGBtW+1QuoqbdcI3J9rsReZDLpPcQYe5XHq5kwHTGSuG5nWDhxsfB8Y0MWit7FG5X5hphvKCTr1K
0Dod8UqgYBFfhdzEBF2KifLLdG7/PT+hMTvIuy266/wLt/4JPsHPdnpAqHqg0g467g0L6J1HTS8O
IPAZ8VK8CrHSRF9UfJKsPHdoLe2zPVZMSQDao0Y17p5pvamMS+9X9EGxEYiaUKL2TV6WV5cZn7z/
O7EFQrqKzqWgJV7VLwGeWmklSt35+leAyn+1YwSck+ZaoufTiApQpd6kGmGEXrrGSJhB2V3SmwTU
KQKvaQd34p0gWSPoG7ZvxSbAGp7y7/8GI+zi8oX7N2Zy/ZwgH8h9XPFv8mM0NFh93lo4VbBDVWm/
XIIMtEAd9fmEdtg9n0Rbh4taNEdrWiPiYrfxqbPwDwjVsyatSSCzKBmaPzkTJ+7rthko63bGSsSp
1dzAG3rtKBFeZbUSD7min5GXbSWyEBNSelWOnRAITlsQh7nuDdtr5PljcCBPKaHizdfiTsZfz7b+
J4xv4UDnZyCOMra8yhZof568vsy/izaV24Qm4ZzF6WJgtUr6kYywndWHmup3tXZx2VUUKGtY0WT0
qZWlRliQJ7ZTRl6WawGrYbTM7oax0SflFVg83Kq5xIv8tFyxPMdzc3fRWKO4VE2HTrNZdxu8l2l7
dMw9hMk0nb/bwiV+CBPwDWLr4PavBmBQ5zc9i0+gRB98AKlMVS3XXdhdJ66UICti+CO9xm0cYs5z
zcZ/DqIsLhVky4HgyYvB/4DYvsqVt05N0NXwZ3fUGe35NVPwDWGwVDailUD35Eh5bM2PiCgzK7CJ
ezueu3HYG7xoUbfXxgA0GtdPgKnPMaadBwgdLx5gJY+h1DA01n6tFNthMaqBY+7Ktf8Kq602+oFC
GMqq1ik5oS+xXn9EpVIPupOmeDB/5j2fuiqf9HtA+g9bnK58UaZTrd/ApmO4V4piaI07KpEbfwO8
8kF9F5Y6hhlpUiShz9n4iSXtfY2VRZYNxkDodIy9HJNZ2lf4FaahHjjmFxl8evKEzOmENhDPRiJW
p3RFGIxxZabTncbxMBQFVKISUqAz5w6vQDLaMf2wv0wp6z+f82CxAssHl1ljYnrEFUEIL+A3av9B
jozyM2EKJF+5+I820Nluq1RAkcrg8vZlW7lRjtZZqHdpHfMyN2vAIRS7aQhTh30YxBqCZE5HUNnt
5o9DndOHnu6jF0ysuDJ7e7Qm2t/OqVoKli4H+PWDNktOXN6uD2E2S206/erQKOOH3FqJYMmEWFSi
hN5xxsDhImqHQ+qr0nnwT6Q91WZY9QXQ434WYHsA/m1MvkTa2eWuMLfuXLN3LYkk0cb40tcAnx7S
KEZX+ZsLhHIfUumVGTUjYgv1OMyEeDUtZF0ATvBz1R2pKPPJd6cPRU8E5vm3PGLj/j80RB34w8dl
pRPGJn8IT0Qftb3rucTiSQMVzi1Vc7F+cprBbSizZile6yPpzPYrHvjDWDNN2h97AFQkAxPHQpQz
GZSmXEsCwFmsjodq+k3kBvhnsLCvpomzCQAk8mwEmCll/XD0XT+hdS4f8hWpjpkoibJwx/t6ybc8
9ttJRdG0ydJdnw2mfFeMSTImXijh/enChuUUgoel6/BxPCiDqSG//jg9uzIGrTMNASoY89AwP0G2
xoQOT8U1YRE5Qv8N3ZGRpklw42nvbFthkpWkZ4TztnQyFGmiMcOveo+OTqia9twTV4LHTBso38Nd
X890bpzqtrHIoUibCdz5+Q7ZrqHBQZHCBfvHNT1fRmIXMiWxtuxkbn0//ze6AwdsJavGl22Pe9Bg
RA7aWohdw7QVQl9ZWPUnodnDNxcndRpCl2Y4U+NxYqloWOaFe9GW9fHzyL6snfmI46WCuJpHEgM0
ua2C9lkd55NZjxYBoxE8WTKnBW4sKG34z4tU4Oe30m3Sc9Gt1DrRymcKu2sfw3LjlveC7glkWfTQ
s4dBCTCSU6x0gq4yqCT6kuzJOgSt+OU38idFzXmJbpLGG+syHw0LYtWATWLpJTQ8qoO5ECZA13gJ
2ArZEoytghqSS+ksoqFpTurolpn6zl5097O3HN3JIZ8mAfAa+n/c56lGJYPRW4U3MW9nRJvYEgcp
XxHZSCkxs411lYw7UdEpWPrTXxWkxn9wCaijOBfJCdeC+AMgJPcdSDJiJLbPOG8gmq1aKQZneYsZ
R8myOOfo3jP6rMD355brwtUMl5dJUQshfsh2WfErLg/MjxIOSxb7ARllTLudwn2+q+Niiqr6hvDn
o0adQRXkOhXK+9hbi/BtgzhErWrkkp2yxLQ6kaeY0XbHMGYnrHoZPkrxRLoAb44e26xFekaylGDG
IFiODZGHk+vgB3hSrFQ5I+5K4jsinXQrGxtblp1eEF7Sm+pxUt20ifBPApxVdoNXuZKv1rNTMG2h
L5G/oXHyZbTBknlzcNsMoHnc6s5dX51Ucs4Dd33vWY7q7hdAFrXO3MU/xVFSVVrq6dCEeLV0yB7q
eec/nTy0zwbhPSDqACLO+K7gmB3kXb0rs2ZLunNmD5YHcuEt06hgt3YS7xhsJ8s9VHeOUKRC1ags
KxVWvNZ0Z+fUvP1ncBz7LMzmV6J0Z/nAVuISIKb5Rl4C5vcfuJbb/okm+93FZCvU6c60zqVJpXSP
E0Rvj7bBtnPLmACFszEyqNwJJ4EDKPX81wZdLXwcq7g6ymrNaDQ31DAWl2J/HvfI0cyc2C3lJKQe
9sd143bMl4pTLcb8mf6ehi38862yptjss6/3L8WhWl8Nr3DPQ3GsHojYy0f38qTIL1al1fKh42Dk
M9q4+luZkMzeR+Qd2P/z49FrokXuh8+jjholt4x57XjnK1eGW1YsWz2NL4RcGET4lUGOae5LR1oa
gx5udepZRbr0RTp3k2Fqu2B9gNkcdstXozlrVyiWymt82GpeuQvVjHPoVz4lZ60LB8jppsvdz3TM
4I64l4RLePpY4ffZ92Qxb+pK0Vbj/xMwLLWqG7C0hbM1fMDKNLqp0yKdXbVs+/6p7X2pFTqNUE1D
jZSQ3JZO/7oFSeg9IlmlZdKN+/k0LTdap8M3T5s2hj7PCRrfi3kaT5mufzcFiY7W0zoBVm3/y1XE
57Ib8BN6sRvTes+T2NmUfwUMBhA1eGlhqBheqFeN8RbVjT8qMHUZi+2BdvxWVPW0iv2Wh7SH06au
nKGSiAyXTd6qP+ghgyipjbB7tiXJBHUiWSbZvU8aa1vPIJU9ouTkHtig+Azg5d+VGDRLCHL1lXHp
9YM1ESPJsPVuy/98YPKGFzz+sAqwa0UjX6qL4XB/MGZqPfh8Y775H2lIYcn44qyun7xt0IN7Laf1
bD4gEdk26mHb7DYNVwGlRcyb9y5y9E3/ektnhVQ10DzgSao/eCPcUhcgmGHtUihIsroUWruo4jqn
OnHak/4emeo+gKoFNC0rWwb5bvao8lPYILSvr5EoLitSiDHTCgYzcH6bd58Ya+IptSJ7YyEf4dFJ
Ea69zSgNEzBOTolResdp00+u9eHakQrkeSQKCVHcRCFxnGO3+GLn923ZomknYnRwtuQW2rvKJCVO
xpV0ql5A6Mah00sB9SIT0Gaj6M3weRSPmFcGQRJPWv+rmulMzgR3cJwJdXqby7pSGsLq/ZaSA6NM
ebMNRyLHpjhQCivCjnAF1roWxJSv4pZaOuUyTLGF2mRPixBUwkfLLOP+DMeN83/pPJ/PzL0e7jkt
2q+vlz2X687/zqH9VGPEegMsNHIJwG3Z8L7sUcDbMD5vgUvjqRkNeCBVjKg9NX0x158TF10WuZlk
c2Ny3cMDIBBtQgnlrwwdxPwq0PH8SRE0oGmiE27r/bDDfc+jG0G9LIZikvFxxjkUemU/rcJaEUyG
guFdSWstV46Mdsy2H1zP/QBjkUzDkJDoby3XQup2bCHicqz7R1mGeAl4uwRUoBGqJXN94z/Cpzw2
/Evh4GFDBQeAA/PZxUOu9H5epyMBBWudR1JHWAmVjTB59Cb318ElTz/FYtAbuc06/8QISmYFYJKx
uLOyA5VopJg9BFMfAFzKv9VcoNXVPFM5LTUAgRvyu/BCK76UwNTdJpKVldKs6eqGniJELDMOp7b5
yW27TNfEWNCcokfeERUCOAUhli2qEG8RIqkHyzk46nf9FyCj/YaLQhDYzqbMtPs6OgcVU7OtUaNS
0/shPD4dLMGQSTychS//MGIXf57wOERuiqJbTNevy1Qk8Qi6Qm7Ei68nPeyX6Ane09y36rrzZTE4
k4t7SwToiWO/bKwztegWlicox/V7/FfNcyyNXfniEZoEpukY86o3i9vUnW2D+iCgzCsUDlgxhjIP
INxdadZhz1pEtqkCariTgzQvOTKq0IZzQHhfAcCypp17VzSV5XLiJoWUjeed0BjS4oK3mBgRKCZz
rXBrMX8kEDbjM+t17R4Fzjk5SlhWslFFl04hT1pLydlUQ1YoCUChrkfsBcepJPKx21uL6TLAPVzR
o2k8+7fwoYDuTSs2UPN94+R6enxFyUwoT/a12JXNIiZiMKnGuUdInBvMyzqDNr4+G9pR886yhvDR
5wRucFTo6YEnikoVRd9B5r9IAB5eMdu7cLOI6MeuSeTYAUiL9gEYrjEZN39BYqiMsq52oyMSqmB5
ombF/XHVCy+QUKRLYb7RhHAuaeKTJFu4nu8w1wiX72muL5W05WmCAk/ZJ1IkkGkvfPHmTqAnkp+4
Kc53P/ve2wOijrcFHnXr83ec+qlFqRzm+tPvWRv4wk9lb0EkEPPmNR9Z5HUdjvnA9kJusHz89hhD
GtryYiiZMRTRM99qXhIpaGASiqXIPMoAcXDG+B1pYlL6P7IpOua+z5V7SJh7eK9V7ci3ETOTP20e
xe/SiMI0xtfVRaUl5JRcCCAqCICFBi2B5SwLmHvIWuKXugXs25Xv98sXO2V6HEImMZeyuyXlTm7U
qCJ6dd8tbXqqvgK2LkkAKpVkSFI6lTQcG6l2juSQdeYvxua2BM47VOmZOQI7KGAW0n4bW+zCvfJi
o3+L+ddBhgAgRdhBnoCiO5NRhMpFUHlqTSUq7gwsPTeKQNORv0+4Re1yZ8QPN1nQYXnec250LXrx
nc8Y5ohHT3g9Xnp0cWWS5TykoopKoTD0WaInY7aAUR2tg+9QBJbykbbV9Y+QPJJRQU4T24ed9RUQ
yHaPS59F/yHAJCD+E7W14yaPHrKKRMbz/sgO59Ut60PGAhk/4n5nqefclsDAyFLXLDEfiw52mYdS
sWj8T0IKQhaYPYDE/uAKPUVzVnaiA8cHwyw7H0VQbteIuWI/q4taNtG4fOACjUzqoawnGPVZP4IO
Jea5+hMOswO60XgZbEZ4zEy6LiVNKtQKyX3aUQyyRobJ30gprC0Dmy85vAcfni318Ax3+RbvELGv
lVIVgoL1R3Fq+H/UFnEVjpuv8WcX3o39hWV2BrRRMzwdovH/w7rRd/tRjYD8EQoytDNIJ1ZGktr0
ZJ1cRY7aKsMV0StoyJilGl9TmpOueJLxSrtvJmo3UHqLdXjTgcY09QVuM6XQ0Tx+fYv6Gp+5j9Ra
U7HBi8tUYaGzxr4vAwptm8fZwwDPCMP6WwxHuUVF6B973q7W75aaAMeweF5Df8ythfWwOJKmaGom
DPHKr6IhmBMB10202oJPzaJhqFS91J8/pSL3q0+sr7UJASRT65r4G/DloCx1J8UeG7I1K1n1d/qD
akFwES142Ux09+EQNefpj6qYiiZKiy+0esOF0B2FmO8VmAVWbw1gIow2bsQrI8PKUQqH3wodNNaH
4BYYIw/PMlf6OCAVhVFMugcpVqF/iTzc5FUGKgFhDdohFyaAb1KljJ/Ar+O0Jo9I+f2qWJOVCuQX
DF80oesDjUG/APiURCRuWLVTf4/sexFobBS6Qab+eYyo5BDJy9HcP9+9Sir6lNpCZsPvawLC4UOc
iiqz78KsiBM3sQvP2ItzI/OQVWYKq6dpVX79u9g2Kft5+NAvNspqFxuXwItCbJGB0djAcvpiLI1S
IESmXsJe/8R4uugqzdA4VoqhUxcr1eaE12D82krC/biBpK2L1rmREfA+lGtBBM2PDz06vVegUYoZ
nMX7KT8A8dnlasmek7H6Iz5JCe0jI4xNX6H00Oi174d730Gb5B41EkC6vRVZ8MJMLeScwxpV2Opl
j6W/oboQbo3ej+Smh3frsDbbxE68du6HuH+2oXYUJWKYvIvOMf6bk0dkVTAO7CJBZovM0TnhqsrL
yrJGR2bFi5TJUjPI+1K2IRe8WNX3bLAuo8zz2V8dgKGO7pxxMRHtA5kL4zY3GfhIX7a5otT812U+
WXyWrvhrbl8fjg6E4lzoCwrAMO7FwHlyRoUF2XDp8267ajZCgqvO2CHa2jO8nkDs2qId+iNP/GRO
iFoJ2iUeMFipk9z/f0pj0XAczpgw8sr1n6+j5D0QonI+LE5+6082cLbMZa6ri5m+TR1A4Sp+q1CS
Kum9RclUE4QnmB+7w7hX1x/cGP3fbPKQoYLo6Vp3U7D85BJOn6nIU2USwv3lwJ2omtFOs5SZmlR5
rYpUBk5EY+i7TnBVDr4DC5nAhDU6PNKk+aHmk8yFUhNwrz8P2QIrRG29ccuL5M4Ddm3mEtXDOb9s
OqR+2VQM89FFmV+nuDtN3bGqJ5ip1lthcllV125L0o1gwQC8PRsOmiD1FLHRYjBAVr+K2P9hdWK2
XDpD25HOTZ6OjLw2VZDxc7ZdPPuC+FCzUIddwwq9QbJR27Zdlpx13ydIaOiZnYNlhLgY+/crzogY
Lve0Q5TbPDj26Lm26XceJJHaniyKnlSVKSB8OZrMNysfa1rg0Adlvnvz5+Efs6CN8Vd7ld8ogKOx
FREZGtiEsNx45HxxyfAt+xY57N9zHFu9Cnr+grJApgkiNiaqpLd3/3n/Pae+1xZGYIfmGg8lpmdS
p+wU6x9PbZNZDa7l1dA9qJceu2jsp08XSlC6fC+hCvFnLg6uljZzbvxAfDgKjiMfBpj4z0XYBSF6
SQUrG71qMF1EYH0E10mKWklS+/X+MnKH/3LGwmeNpZgrMs5kOiI8S+akRWsCJfG23SyTolnB/GlJ
ArsxJYu5tETbxhJ+FsY0pw3Zh09dM2AmRsamV5/ahoew/KMMrqXMAn+Uxw04SkIS/dr4+76j/Ohh
huvIU28G9nCWJWSFRSMFvR0hFqBz01Xn9rzroQQYYuimyMv3KWsVnU0zAwzjVnZS8vRXsj0731iM
1GQ+tjIu0x8p5uXrAS2hrglRNtLETBh0lodR0RQYPQdumG4ejowYTXD1UMdxQxJaSh9Bp0RqsfWe
4xLY7I6Iogr7IJC0al1LtgPUID/DH6ePiVbBCzNAQ0tDW5HnnxIP7/Rr74gYvjOZ4VpRvK7GDPwG
WuLaWF3JoL1TqaeRczaF5lBbASDNeCKBsuSrR2K0DdkdY/EXO+61l92grNa/oLEtozvkyAir99kA
z+OUXmyakezZOXqhk/BZ8JKyvAhwZ+fl38UE+iqAxcglqWNnl/ScGUxOAbkyzGreBBrOn2GQPtzx
JSt4HWc//8dXYpU4c4sBuRv01oX15FXEmWZ1JvFq94YNSTa0QYcFMUYicfkyKzRRbZ/bQiLgYtKb
qTsBdKHM9MPEWdU2T9O/4ucsQ79O0FMKDYUo2BlpfPNx3ud4732qQlm5lpPBh5ogsrJ8pdzwnpXL
ZpMxDaY/HDZGfJrFjuQnDY5RA/+VoHzFNvh8w6rNZUzn8hBvc7fbRPQzGJpshssqbRWuASaYfO1o
jWdttM0pv+sF92Ac7AKWUNRIXHi/eEx8VyKJKqAF4P5TCnFL3rv8N0DxhAVoZR8GcWdyw7T+lkP/
G9pM5d6F7WMOq5KIc4JlmoqqPhQbdWMJsVSzbcYFQk6/38hGl9U4EZLJTH9olcwQGzmUHH9uWtXb
DIp+SqurcACBEISIm24t7OxajZG3DJmYDOToz+ZmXAiPmkGjXmh0irCYQHUZQnM6PdJM+yb1dxXZ
jqFxtBhJKXoIXwga9Xs6JyUjEn2atBfJnNWPiLyorEIlkxQiBdGDODA2y0W0svP7v6cXeRo/7WRN
z9NPG2uAnTQ1FMG3gQIOSQOKBfNhQB7aHUC0cUNWk4SxDNbIBLfTiiTIC2sJvDkgqDHwo7n+M2z5
YyXdwhwIJUiC+1na0DkZ8lVO9MWD+HaRmGbReRBLbmd0d4A+WmZYDQBVsiybDFeCzGuc/IqepqqD
GafH0HCQwc+VR32+WgRaU8BXLQ5u6Y40yEDYmY1lxeYbPsAAfpFd6N4t7ejVy63yPkg+tcnNQhE0
d1x3HvDNtIoYeU9YEtrZdNMWxONRclXhhx7CEYL9IB9tsx/ruCDMeS1n+rC0PxWRCnHcT2FE0mo2
etUySkfk9rrqrXuN9j5jRLC41aOjidLK9C7IPh0uK7a5fmOaArD/bFagbTNCXrvFVpuw7XdI8nZY
G3uT8JNJrYjGV3t4FT5gZBiQVFqapWXD3BgAfMRfT5g4A1TNj+qYaUteZBsvZu4R2Ch3FmDFFmQg
2rVJONabsGWDvwMsNDM5TKgkNb1V0eoXLs41UnQNZcbnhnYJGS9L4GZTYiXQ404c6Wcon+C+UCYb
m6nNefMrzzXjDsi1DfrZpxN51EF9gpn7BG445zf3Z4NIalDq8Q5E+kCl1WMtDYzoMaWe5j2h85v3
6qMqitApmNL5FjBmRahA61QNfFpAuI4zdcCuUAkP29QaYoTxHPKit5geZihgiH926ybukn3ZhiWl
vh0ED/s4by+Z3DjgvAwCPKx8fDyjP5W4eFmNNnpelhhGEcgloe5aVhFIXjDE58wMnpf6c+Wm1cTk
eVC9Us4+L+8dDI50F8g2RYUoEHcYb6RfapkG57jKr6Ed4ant5etgZywqaHs/iOciTPI/h3QN5e0+
3kh48wXNKy//lxUyJh+kkcCnmhmMk3FvS1WNVATbeEKCEjQB2ec8ID2TnieGMGcXy3QodssJpND4
mw3qWQiOXWx5YO6jIh+tgfgSHydm92JLKg2Q6dMD+A3QNK4elLYVKwvz6HpYTjFX5ZpjlqD0KlPA
15vKLMwF/MdP1svBSl34qirLjneR2TOjqOBiUXMTr9bwkJ91Jy/rqJqZlQrouKxolfF+i0TYRVJ/
Ed4b9xtXfXzb7Rpu5JBdFGyfD8eKLQBLwWzM0ray34/890mUaajuG1Kiv4drNQJcIDOsJrAPlIQ4
RKyWBJUssQNxz+mZtJGFtK/IRTvpRJYJYVBneihQcDmh86xVitZ/AwBYYeQbIxnwyBIys48ldTln
qH5RQnUVqaEJgVbCPXxa2CaKD+9+WWmPw715NVOq7IVIkTJyRYssnIVsNZd7pNWdr9oCiah1IdDZ
rdPJew1JVrEsp9iQj8ZvGMTft4nZkUo7N7knIs6KzLwAJHpCjbl8PE7wDYusLSw0rUoqAuwKsunq
TND2m5PTYtUD8tIWirCXPnS8crb8SYKXHMRsEd6EAt31gsyp0enM5tZACGM1uOvxTbwMJyqttg+e
D3621bDbysDCYk7uC29KEG/2tuCjmbeHpIpQRaTcjkiP/k5RoEL/rG4rYk/yZeZNYyCx/L4pt2yh
Pzbr4MQ9QumXMgEqZzwyvbh3c8Bd5I6BfpG14VGgbK2pwwTfXRF/OY0m0W7Wzbsa7jfQWD8Xa3eK
QVQKx+CUoqbqi/pUFo50wd/63R7L75VzXbmhAMECdzyigoQEZ9Z9yOdvGvxUKGu1B9KPHqr7EJLI
3+438k5jyTIChjM/za/wA/BPJXruqNu8FCfSWiiJKuccg1DYfjOsm0Z3gM3zgJahU81KgoSghh3y
mpn9vQ9wIlZFocL+D9m3B+LEc5ecCDrrIrp/4NKHI+6TluxoqYopJkk1aVmaUIatFpVrw9UjckJk
rkhNNdL5KjkCJyqD6VS0ygeiFnh3Na+MabLSRnFbq/+7JaaVQvnxwfUnYKkNHMCFKF5xDp173m3l
Zg1x7Uo1j1BpNWFzQJvZ21K4Ln88geaMqlT54J5Y0Po+62gtgfu7dQYr9VtbeDVFIxWqiJ9gWLxj
6NnTTKe4sNPsCISGTptSn72f7mT7vPAgcrVWgam5ICmVJ9SmlgEegjmKxu12jVWsp2ac4M5N5qU5
3Y18nUbKl3/lgvTKawJVuYJ0BG522FMPq1X//rsqOkiiB+JUi/B3vS6n4Wk0AhNt+SWYQKMWZQan
OEQD83oUCEFqHb0kLxrQptOvkoArwnp0xV5uOSE1ODbnE2hDcwPzlr9nguq1yeou1EZFAdp/+IOU
6F++ccFt/RqxeoL7RYoTb79uDHWiwpdAux37u3n2prZVtn0c1PQbwEDGX8jxv7gKDTEP0MIbGw8R
l/L+X8CfvXN8guuti2HCCQw2dLvQxqcXJwC3F1h6STBA45FZllMo5jvJjhru3oM+3ZfFiBPE1JiK
hFLEgw+k+MP2nLPk40UbYYRGoiPq6PQC/FXxYSdoxbsci7T48rx7DkP/vJ2ysotIyWo9v+KdLwQ+
vE9SGaMSVz8yV+OWcVem2wniqoa7yinrq0vh3Oqh8QraX6IXMJQjHw+hV8FDTqE6iEcHoL3jjzWo
Bn/ZrzyAFBFr+te7K+U3yCdn7VbkIAik44ipL0WIgsZUbDQ37i6c0xgWFmqETd9AwYHHuYzaVkS+
s7cXpJWvNtvsnQQxDJt1AOpLoxwHVjh4GOBsDsropvSW0ayvtY/DY8BvRAzwsWsuo+tuuJX8/2Uk
uM6fL5dvFXYUWfhV4ktFGqlxDVPxHFmkhyPps69LApmxhnNjwnOId+ZedeVm+8ORETtRi+l6wIWw
ws0PT4lV1s3DVEqMkEI4JHF8W7HXbAOV84bx+GZ1+RNxr2Uzy/CuNHG1lf0NRZ6y8bA8ppVrC4Lm
IVcKMLTSzdGZO7+TSjOAV5JDdGuDuEZB+BXxQZgKXPpiJ3Rh9JZsBGbBLtZpG/PntSWvUg0aPtPQ
TpBagMXoRW5AOwyjwfO2zXEit9YdQSX4gLDCebUaY4YUUWfe8KKgU3mt+4FpBE98cq7hktRkk353
wQAUE9tYhHykp7nkqADbOn63+knZDJ4b8C9DerTFP95IgtRaAchyuUP8mpPjdORkouwLHUVdFlL9
3whIGXaL+OG2nWZE1ZDxLfbLMx1ZQrJiJ+nP/kVRmOLxihi6CBhCU7T+rJ5IRFx+SkX73z7094jF
0ERcPan9/RmAstMGwTckjkKSsLHJYFR7+wjeEuVjIyUYpU8N4pV4eM2b0o1h3tpr/2wkZRCNE5Mt
pw4zehwVv2EmhtV73HjvF/6GuatAujtB72lsZ6g+2IgP8R76maecjFFJ/7bJ6ZPrnUuOofbg7Xaw
DumOSgxbX25mIBK+1jHZ4/zpUv6jDGl51KCagqXkFHNfYNJFCR6JT3AU5kGHTGxgFzVv0e6Jsbow
JKM4hkfBGEvwcNmJACTJyoy8IQolr6eG0nINuObYMGYOQtHm215tTATF4FYQCqK3bMmgPE2DPn++
fRA4JwMN5dF8C1przs8Vu28n8+y5KpNt4GDlx1S/Am+JcTpF/m6BjD20vWmYxTtHVujbbz1zlKSM
O4Ym89aTDLmWveOkMeU9k32FtXH/z2TceyRrQsSUFtDUDrDw2OHZp7zzbMtSgYhclNtLBmoV2ChF
6FuvPGsaTjVtnokgTulwM/IwTvXIgn8R+oNzO7+O8eUYmhwLVbfa5GU7ogCg5YrDWcueqwFHOUHK
7h0N0FI8A8b4zPObx8XGUVJZRN5lX8eC7RYH2KSXRS9DVOtW8/VEA9YriKJJ4wHzhzz1i1w/ohUk
Zly+qtqqwrYxkILEj6KFzfWRW6//FJtOSNN1JJuDseE3CRv5jIYTPr2APxIlevZQF1i7gAy3KKPG
MCy0/TF+oLTvtphn1qJo2zTVMdqoWgo84oPE3ouB3c6aK4MFFTRlzGIqPRznm2wfnqyWwunZPsoO
UeV05Lw0JwVe71WwUpJlfqBxzX/VSIRIHnk1jpzOF6prqbZUvWr+4Cb1W+vFnzIrzduHFNNq4agZ
ZjdzbQvIXemvBRAxQv4qLeSg49P6AVW34VIt0v9rOJvZS9empCf2jCk6fG5bQP94A1t0s/ZtYCfE
lEJhXXiCkB+thX2zmx7OFrZJcUF/MVUJFHCJ5t37XI8N4AMug5+OR+d/Ud2r+TOxfaCCwfndNpRk
LlDxEuufBbDfQFwitu3GKCCdlLLL8zj/1zDyjdRqVv4n9PjHN44w8dIPnxdBFV8J+3T03QcW56BI
l1nU/TTh44aTbw4OACYcvNfDU5S7bx5tLNzxQGspz6YgQ1GnrBZ9qkeHEnH95MRzH8GkrgoDtTiT
gdr0uBE57AZB5HhcecsT1X6JcnueXvdy3xTy4nW6COTcDe8DkImNWjTPT+JQC1t+1grvhOAYc8ma
3H5v+zTEsBbWbn/t4EGjrG5FRpu5RQ6rIe+HJ193Ay5+PFkk2jvZz6nWW+HZpZh77x7NpzdUTLJT
S+U0nblhLpA1r1ROMtJ++QQ2P1ZNqXHJxA/vhY1lje8AjOouSp5alO0yB/jsxkLUnMCH0B+aG1wh
LEM3O7MCBOzTzfV2Fk/uY5WPf+T5ZNmpoKpJ8Y6UPgP6KDsMFXllNPatU0kusPrABgM5JvqZoES6
9wPl3+vsjOvrQgVkTOQBhPEhHW/wZgdsQ73dYCGynPPjN4bJcn8gDQFb1189T5gSatclIBQwhFS5
k1o9RUr4UQswQbe/Yij1ocH7ICd+wWfY4itnvjq4X+bcfsi3E+W7ant0XF2cKSMy+e1b53Q3wqhK
emmrstLx4Lb+FVTy2M+m1sId2x6AwG9ITa5uX1SLEDm0tycBTyepdFGv8FtPxUd7riS3WDTCvFs/
RL6bAmnr4dZcGcJkbmBCNG8E4di8eOWaXjL52cpD3hHCxXh1EEIndncYIrYUfeXgiFM1r1hl0JTD
kHrSn6c82EwmBXZzveiOzL7VqHvtuWajPw2/aX909Sq49kLbGFEiYmcAg0bpYqj7bI+00n9+Dn1l
/Cmpjb3n5gkFIMs1a/Ncbt4ryQw2LEedynEwQYb7b3G9QRuAI9c+eNTA3b7xGVWkfYdMNWwTxfMS
3jCaGg7Iqet9xNnXb241w2c9DfDuICczhl+/TLWy4xLY4xFy6E0vBlPYtA6nIgLmemtEa1Ent30E
ipKDZKKEUrfhJO0kFxbPmOytGiqDTsKYNRpNZtbVQA5dWZqD8C0vpi1BcfwonUrBYpA/DFXwb8uA
dRAwC25H0P7fwY/MGrICMWHJL3R//ijqI89lT2JtA7emYmXoDnnSNyI9S5OmAMfGgqWkhN5ovyZ/
yVwS0CIZypEzERmI9Y2JBQVEgiqQOZkqQnCNEG2bSE+AQwfp3hL2ZqbpIkorenKg+fM9yt/5Idva
njyrhAAxBE2pJnhubNimle4ZSZCyKmdhKp0E1D6xgBh1RtilhCNpe3vvsc5kM/U1uGd+tgPTmd9u
Pk+gGeIFgOLsmmFgL5F4fa1ivKK280DajTQdCVy3W+6hRjam5uyTVnY0M9lVYeUvk8ivd/YLngRt
cDHXRUuj1tHGTwwy5fAcKAQR2Yth7xR1rV5H6ozNYFL1tKbeNNtj2yNwS6qnCLBpNZYJSxDnm9q+
hZDRo/FDqfQqJz/5vGYDPdJm7hW3owRMm8GuX9vgi30evKd3UJWgllIHEOLYSNJgK6OfjM9WjV+3
3mkpTsCgExRD+WYx9U0Mm4vidWxCbU9dAgAGHB2O7fX8bmLzoJAVlXHGRCkbppH4JqjDwl7FilGG
RN+gul2IYfrPCvC3LkqpBJDT+K3Px4ZC8t6Cb3ZqQz0B4u5E9honFJ5ZIQmoY5Z2ZvRXc4Z+WX28
9E9tG0EEVRpboH8zeULh+DTceJDY3y94Y5sdeTnQSK20QCTuqBmrXKBtNV8ZuZmO9WeC8d5d8Aad
kemNhzVcvRJkcA5SDdboph4drqTj54qAKtCOzMSbUBHDhfzADfT6y3PLHHfd9Jnlcf+MjKO1eeNu
rKp4vp6LMl7XaX/Uv74keS2LjwlUWFgSTaJv++ehWlKHqzTykG+CAZc+GSbc+1EBU6oiiOdmGEYb
1BY2dfFLIjYQVa9fOcLumQbOc8Q1uJyqlAeIOiXl0dnmYEPihuIJb7GVs50kX5lKOmIr44F3bCeI
pl/L5K8TQMYzW1UST6a3jjA++CUm94vBBnJj+7Frlg5MJ1VgkCaQi29GqdbWcN3A+uQ+VNM3SAyo
3zuRqjAPuQGR6XZCx5rnLDP5XfPHKhxDuMLdOEcMyW9jZW8nADM2H897rANPl2hJsaoRdK3iOHgZ
87YrI7lC/O3oM7nhSMUoVyUh9to3FUELj451ejWvzxSLeHphlJMTcAHPWzIC7sgIm63rrTPpOjDI
ok59P2Kzipjidvr94Z/Hw2rweXeBKrlYENn0DpEwnaZ2koDqZAXXOp3h9B3E7s7Xa3bqxpXGkOo3
j+Zz7zjVeBYq9M6UNO2yZxg5Q5ooxpPjbUoyRrhh+KfouwbsP8KCEvM+vi4G9o3/hcjcF27vZcup
yAYQG35ka7sSm12h3NE9OLynlL0dcmutf+NiWapT5llRDqE1BUt8rOKI0B5jAGZOTD9JLpMaOgHf
K4xj3eEx9+KhbmHRaUCmKfz9T5uCPmv84PeI+vYy1086zoQW06qIc7So0DeMBhl/R1xWN/BIp8fS
DNrlmRXlGnVwbbvpJGp3vcdEhSbRs9GMpzRPnwPqEuENfVWVvHgY+t/8UOpcGnNy+YKkXL6Vm/w9
emxD0dp+e7C6ZW2biuiIrTK9aBBVyr9o16Wj6Nycm95C+UwKudPLNFVjw4vbzc3Dj8+rut2PmO4N
d5hBkCmKjvE2pO/0hoeh2+G8WxDBOYnyDbDnaIrJoTLvsgYq/iRkqAg0lbtOzB/AH1yU68v2rL14
fm5qDQTF72Ry1Oqjw9lzVtBF/DCicD/SM3NEAe0ajPI4KWADGJMwp4/smMaqs9CG6FK0GyB4QEKM
TqhgcT4G8UkqaeCN2O4wKcJ6VsgJzdENo0eM868k5NSFvSpZhQoduKqwDPJvBmcTLbbaisShUHL0
x+sPudP18RG2K33E/onhTOgyyAoffQ8oTxGehf1xjXSyWtFbK9sAjxRRRGZVvHFP1Iy92tebpQIO
uK2svOri4Ot7e9KkbigIIiPAKv2Pm2iruhuE0idxbFP6x87dFnTUDo5V5eCyGd9WQhp0dg8YSkJk
YUCN9TBLEY93hsEPUv8+rFRbkFKZSI7KT0AHjromBP82ThjnaHlB6tx4vKCElMNQ8bWm52C367qi
B1YdtZ71n+YRgheXiIemxH3b+wD2qEj7xPdnEHvZUaTrHiugDG2kihXddUkWaQQNWPocpTxru0eT
4N5/mjXpztCfPCbm257ixyUKIBdNWdlHLGMG6CJt9u25xp5hVV9z2689EU32euFTqsxU4ee9CNo2
1u5JF6Pgx1Rmkbx6YbyZTmo/vdDkWCuQVqE74Rkx75USmxBe7GQOZj3H8RPi8WLzHxUqqjIMCC6A
gKm0T3paIZhMz6a3yTmUtsupE+YWeZjiWSXcbcm8oKsLp2sj43gVSDFSVFfTkRSPiH/g7r3+KMXU
g9wTPqV4vEIL04GRz0wGFvYGGNMD471MoC9WlgOvE6kuTVKHLgLhISODpIOO+KXC+Wz6cG5T89lv
BxyEZqvilpyNPOMAkjHbAN6xAgv5QiSddlHJu4inuX5c6ZWWrPtb2ceynfMDlQl+oumFcaDP0aS+
NMs5Z9CbE7s9YpvyExnNvgZl95Al6cevyNiwjXHRHQK34HH4V7xly0PmDFP3ynZwYsejCnlVrWnY
iSU/PtHrC52Sjy6JISfqnh1Q1U4/luI161sAhKw9dPQLAereXMADsH2EFZx2RqRTlOCQV/S+gLWq
HecIPsuDGwSg+m85HK5do9KTvjnR6YymJv8u700Jr02N0IuuG8xAVdCs4DoB7U6rAxHz41c3fUG2
ezU8YWhCSXL55LAV8A54wKG/Pxv05v0q69vN6meiL/GBurM/StNvUcG8VOEeC4/AbIYAbfRC01dJ
5MhHRVEOjdxnZyUXxmRJy06M7enSB4h7eKY8cuKy6HiWtSiZU2yVnePhCR5wV8JgqbQAduf2We9h
MCAReozVJ8zNhQ1SsSPfxun4+zCC6pnbhBJPj5NCWKnvynu88snyrP1t9ZdgPo0Zy6JAYZOPfiRk
FD7Lq4YUx3bbZfokiREwJwC1xszdRK61bULI4/TgVOo0sKVxwrgBfOCUId4E0wF0+TVIvId01Ulz
TugNfth9p56RkrQcNfzx6LZYOFpDCi0xcRPfoIYyUsqppWW55XIkLY2ZIHpUf7CX/argLu3lYDJ5
GVLWsbTNrzR3dRpqZJvWtfokjJr3KGoRlYhKFSdSgY5LzWqkkCMOW007xmlxalhGrXm4h59ExUYE
IgyOF8isxO5k9v3zVwo2Dwy7cB/uQPVKZoEygqb5IRvqAcynEd3pCMFTvmRZv4wKEN8uPqkQYe1g
wFgniPaL20dZ5jXio6kseJfNMqKzB9eYgB9LWToI7Kud7v/QFKHqZ7BOkS9QU6K6IGKF9CicyBIi
jmVCNBGyswqYbxosVS/dWerC5a3hXszPaBGXuU4I3HBoAFD/+FaLhKu4158tOL9T3xUlKsWBT8gk
6EmQA67zdmBcSKHNT1TjnzbjYpsyxlmQNMwwOLHbZWKN7vVZS8wxXzgvNKyrk9c2jr/9mKatO3Af
TmBfDFT6P1u7HWgJLW5KlNG4mSuyUIL/ecm1f6U3hkkI7OFK2PXmkWLdqxhMk3QnX+zrP/z71DH8
0kvmWR2acRgCD67rjD/NoSWnng5g2MoR4cdnpLcYPz/s6/pmNhHvSJlCTwXu+8RAOGiIAvYOec66
bUVEF1Syjhw37e74NBvCaNmGrV8wXoGs9HId+QI+CPScAlPTNK8vAk9YZtCbz7kjJGKS0ZBKTcS8
iu13maiY2QutrRG0FN+iziadgwWwxshTN9AEWhpbZEU+9W5uD0QplFVMJJ1J5uRMeQjzuMZ0cv1t
FOWI+o6aHnkjf1Zs4KIn/HHBlYd6755jOF4ffrbILAQRoFyK2xqrsDS76xpWiSTFsUbIlPWu57Am
ylwKKeAyE2JXWSvjhOmDPJcBu+TjHVd+LlCBwkQ+ZWH53LSkOtKo3CNA8eg+hy+wncpexn2fF6Tw
KSh9WVDFIJNcGc+l+zsSoHFPLOi+PAHrElrPA0CUVCt3eq+HAaIlSg6fNI5xCoCKcfeSBeTinHbd
Zr1OwNjNRYXwyg3N9w7QSXSF3+1Prv1Ha2UM+NDHN3iELv7ZcOauFLou6grtOBM9dZeQbzMkGI63
n05E5GGG88leAENlH7fxFRQFYVKN65wnBL8aMZC9FLUQFEcCLzcOJPuC43iA6vpWut3ZNmd2unnN
CB8YBVZ2Cvqf9AfXyo3MDB4UK1OYTXaU8PsNsyTRSAiqmCVnnkI9uieNdiXbZszrkLbsaDqLaHM2
xVgADJeZXyF7y0dJr/WRjEMF0YYZDUaAdV92atMgK/2vPeaggFZ82VfiXoO4FJopqTvW91LAzlTC
SFzRUxiMPZwqnn2jpjlk6AWwu4FPpPymKhzD1619tXTylZ2elgc8zysnc46ElNrmfUyQ6ku+Z2jC
i6cs50eb5NKmB9iVmGX/CetB8KxyOi6AkgBUNwqAJYhI1fD0fXdAkQR79ysNSOSl4urub8maAxNM
pH/+dJmOVJppyFodysvp453QjWfQ9AlIp/R5B2oEIJIAKpjyCzrws1+fKSrPmYWqFQ2QhpG7bO5L
mILKAFraE1NTuPGcLteqqrLKXAiqkjotaNEXDGI05sI4CV8jhiCNEX023UHG2Wf+HVBTg6FNmq+q
QcNnw/9ntjujodbTMt1PUnO/2/c5xiT3ffnIXjvpKpyjIN0/kMI72WGIg0lTKVby6Kfu+1jsYNTW
WSG3E+kPPUAFZJDVl3YCO7VlYHUmqvTBwqIDuk2rg92xH7WQNZOP/LWt/EA17XRnMDDczGBifhwE
aW+62YlHNFNE/uTbRqkjSgyN3Hl3tvi13EvF8GLWAcU9Z2uVxl6h1HOAnj0wXvVE28MJIP7xtbX1
8dxVnfaVseWkXsBQhxsmV5t8LOaaTtJOYvypJCQ2mJ7ysgvkNidsIl1Kb4d7jVSC8PhOoqEkfzwW
7jRbuCbfgIL6dg2tODzhZr83jJT4d2lFAl5jO+uNWPK8f7bHJjHXo7/887knhB6/JiLouNqgrOhQ
apP/PoVcNeHojzOL/CYeKvtMFLLqyV1lOR/KKPsWmcfl6x8DmtREU64JcFTfjWt9XEjcRyUbS06u
z5PDp4PZ7FXd0lrA+j8EYe/w7Z7SllspVNwOc6HcKwnafEdjN6Ykd6AEE7U1Jgjh4gaH20c8PPwv
N06pJbpmQ8FmNM/ZgSX7orcc/8qRF7d7JcFS5/azFF63RLaARST/DP2O9vmoAIx3UKotTL+Rz8h9
IDEIehkcQvVfy9GVBUTPZ/T8ObOMQJbpFTSF7Wrd17OvntHeyhhK1o+5OUu/p9BcgvrEaJ2bArT9
TihrwUEb/vNzrTSgYtdH1l4RV24lOldCJBS9LfDh+eDkNjwkQ6WETEAUUBa4Nty80o2HYHKk1jyr
SUlZKsSoauNdrFEnoCTaIC78YF8bMT7DmN9eCUG3Ts6HBwlWGO00vlUSAomDYPblRAxF2JDNxSPD
loqdlENQPdxyjkl+zA0W5AxQ6RfIU44OMHyv/NeDw9SkPoo8KSH9OlVWY4cnGF19/FQ+TAr6U+vD
dwpqzza7Zf90k80cWiBhWtW7c4vVUJk/DlFakCDgztP8FlO/qzw9Ra4FXkmJrbl7K3hvSkoXHXwN
QCqR9ez0ik021jqtaZKvKmexi1z+uDGZtz0mtGfHwlxdKkQLq1HfjlsKQekMppCOU1pbsiW1ViP8
aLR9I7zkYUWi0ssXJiOfMjN9pfFEge/83i407qkWQ2+fvsgB0GWDuwYjd2HOJgYUs/wSsQTtB44n
Hi/jd1sqlSlDg4kWuIS90urGetSFod8MQGivMZWU7cQXFffWWlSJU0W0ll0n0DF47eSU0xmsVtCp
D8Udmc6cG+CYNqj2xsorq/LTcviOKncRPiExiVS2/HLIVZGhqreumUz+VGk2oAdPq+DOXPlrdfq5
xr5Jr8qsLMCdq+vLiJnVYtWVQLUKwnirWAKrTWx+HJzdBkeWw6IZGa3nJ0Juk0BsLiFXI4oNNnqL
Tip6Y5WtVGQ1v4DyevtUDqwjMF9GKMnLpTu0V3n6x0dJzeXUVW7wzfpTQu5wxHST7HH6GMnkhAih
NSAjpY0PJlGvi0JTcHAnvnvTIiYwLSe9PmrtURqQH+EEc9i0egNbUoXbdrjxtUJEEfwsBQc2mtW/
pm/GIu8m813oulGfX0ZQmSB5t+vExD88kboLfoHJtyoPJaDb9Q0aGywKob5PU1QN6/CYJDTyHcZj
SQEtrxQ8eDF7eYKv9nR5s7ZgNXy/fx29fWpRafkc7dcb08H3bPwDp5GLbSRoiU96gtK7LrETM1hk
k6r/wstOXwgXCjF6uTFEWKz9xIySXDWZL+BczvR50pUeQk81pAKL3WLpRA3e1AW+aZuVIDcigFgq
yWv12i4/jE587phoRd8XfsEB2Avwuf6NHDA+SaJhlT2F8ECbWMZXlO5WYhXyYwCETVUHvaU9K27J
o37g7qFScjIDMSm+SuMydJWyMkb+SKSz1Ovl32jNrB9eoJWL+yboElyA8Tp/Up/kJ203pAlf62ph
fnInTiY6mFiZ4PUgIJsUE1IIHveiA4Q0XF95gfG0gUV90ZbpU+Cemn0P0Syw9spU4dRd+fRXk+3j
6ZzFvVxd9eKgEQ+dMwYcvoq37rTuMJqHqVNJCxp280BzQb/4E0yPxdXKlMXg1d9344J5swnnNbOo
uvH1Ra137dZyv9TowE1YMM7UcFUwwYSQQqBe3I+nAzlpSGQVnVesPCLS7Ff1WakpWsGE5aps2qcb
1iyZ1aS3njMDnFLFFY13NK1bJ0J2vQ55rL3QZNzd0Fuf4Q27Mwmn153COhFomusitgWhsu70X4oF
BuE/bKOSSrdG2i43xO/zcqqaTYJI+PZkoio4ommu2gxaiBJ8tjIwLee8RSlkWLKhW9j/WLZNSh1l
I2pd3XvytMiJ+XGbu2+R8kTh2oCAYkCyHdrvfQ26V5An3h3nVWZ+dFRbqF2a1msPdAo0D3H0fLxQ
4uDTO3Le8M9k942hyFPtJlchU+M1Kz5mC7FTIOmw9s0YqKX87M6k4ndmOJ36IBqzXTD7JLYjhjcm
j57AH9sPOcNvfEXOSA1IKuB38O8LcnAYEPhtLdkTm6OvdhHq2EGwAXS7c/Psa+Mmpee1WE+pdrV8
+TOhJ/XpPVASlBXrXvk5EjXDISUb4uJsmFSgM20UWXnVz15wEQruHWfqQB70txgbO74jpyQCy1kd
heGnKyuTxZ491fmlcIiP6ulHQNmR/0fzOBApFArpM6narfcPC5a/kC+R73uP9E/1PkBC06RhXVCj
vRdYgE3g3W4amSDWSc4BHZMD97HmgYDveelKJHCYx9zu+8D5HcgS+DPCE8Aa4IBbM4FNnITV7lpJ
yDxjz/euiG++WIr/GdV9JpJ2toakWt18+evmqcJD633jZ0f1/ySVddO/LGR2JSC4oOVdtooa9rx0
JTFm1Cp5OjfsnrMotF6jgNGUxgvDv/28FvVAw3ztc0rdPqq+9XsIYVRHErjUJqmt7RoENwmiT/T3
QwUdzRVvAopuxCh8Q5ecbMBSFmsqxarcXv7VZnDrq+e20iPOjdEGGkA886UOeqhfQzm7nJIuj8MG
1BVksWe17p4GfeYB7yTMmUopMoEiTxq7MlB6O8OP4b2l7dJC/lO0CMMBsR3EHYb5F/fluvqTKS//
ajG3KfTABFFBFUAbiJnl6V9Lez2yK2X69KjNTFLyHbBlZBoP1h6DLcac8LUX0CcmY2ILWMvKLZei
p+EZWruLzvJIgTV5i0JkhC5ZJHsXs29pY73+KlNQCXXirZGBoJObf0y9or6ZUfZHwt8vhNO6Qnbj
DR7P5zMLLOLSUdppbcFK7SOITrB2SXmRVi6tE8fWdphnDl5VbsRTedtD2ye1u0waIxMhZK/t+jhn
10kTnguEd69IA/ueluyxiqdMekFDPYFBqzzriv2JQ+lqRC2N634Ni576I/v6KEDqzBtvNb4DTITq
pFD/Q54uERLBMp9+GXkPupxE1wOoKSWacQwd8vwEM5WZrumm9yZT4/fqNs98Z8eDArXZ3xitIq7d
k6whN+1dScTo8lpQalDCpSwzoBgqkZSpcot+DremtkO8fOnzvsZgvN8JeLWRCxvGuTa3So6rjqs9
P2mqCObXzSsW8n2iXX8RfO36QDHEeqE2PpS1WXvfFPZqSlAkwYeVVRk9D1maGCGZSL64p+fzex//
sMRtg6iA3HSc6fHQBvFkEtZvA76/Ut3wAgGE4J+gd4n2pdD+wcjDzZoXg5usVd6MLRvuKiwBKd/9
eEXNUgvdKS7xJGmuoEeo727WIVz67K6Ai7oTAcQb0XLuokvYiiHKb8tKzHdJYjh363CMpBaS/L9K
7IkOB+KZDu2jJab45lh+wTYpZo5+EA/MQkQjPwwnzRK/C9LO8Sk2R+Mp001Dxj6c9MLKt29I6Akc
QLWAvP8uOg5GgQFMhUyGmD9mXV+Nh+Sanop/DthDYHPfeapkeZ0l2IoBDXQF7WmBHtLmA+V1ntRe
mJ35jN7E4W+OMIUbIkWtNlU3PoRLwaemV3gsfCJHcUSfR5cCtuR7QEXp8qdWdvRKxmEUZ/UmOX00
IXA1rm/z/m4TdLqwdI1AfTW/JGuJXWFHlHfQ2sXVi8DveWC619eo19xvDcVYpe42pAPoljwAYjtq
uAy+fLROWS3Q9L8ssq8pQC/cW17+jIJzEhrWGtNeGaKyzXDbfHElb+/zgNZeS0kBapsZuP8hjZp9
nDOFER63DRvaCgrF/b5KqQ+7xLL40Q8vjxKuSJBZs8Bk3r/0VwVePjyn3yqEnnG3pd54unH24W4D
KdPz4jNTswBYl37OMhr7A49u6P4wpvNYkz8AZsb3/xPJJhcX387s7gV+paVwkM4YfT/gwaikpB0b
Snxu3M62KqlevULXuHn2tXp8gAW1wpOaj/A+AMfOR28PFQVUGHc3XrhBaKJ0BvsnP1htxBLB1jmp
PHO6kvB8F+mzCDChPRmV2uZN+A1MPv/pCr4UpiJIEPEC2jZOKWFx3AC4+YZcB7QHkjnsdWth+mqw
u3eveR+i4b6wEPcL2c25iVocaSiEMLSC7AWyi3Hr4nUTOrSUzc+kbXRiZ4mtyf+olLuat/jr4Ck6
XEeW7mSYuxlIj+KB4zvq0/NrGVyG/TDhHTK/7VlZaiFGYaJNJ4lu8IPtPiAXHl8UDq5yPP/PXQyI
iPx2AiZfcK8KW9qUYeKw2LDDMzkQEXi/aLzrTax/PpbBiVh8u+Kkjy5LLTzqwEPcyoGF5TWPBWI4
zB79BuwPufh+U+MO5YEdPcUBk4cNBUBDYFL0xRIELNPk6sxsaeKV/S/3AyrnD2fLFJNYj6+TLgoH
tQJbq1JQF2GZds59a4gTNGRB+oxruCxS1SFvVujaZ538q0ZPsOprGKjGztmO05u93A/LRz8vVtHz
Mp7reUc/v037p5EbM2Iryuj3fIHcLMX+nDP161MsZR0NHkV/NWemowSUkPYffNk2aVN2jeMDLUlX
msPNp8GbjgS3IeIsAbVSO+1cXZOqs7vHCnHi6UyK7kKTfeiAS1mVFmMzUFlzNkDyLXwXyI75ak8N
32Nzz3I/H7XkBJJkX/JJJKgow+ixpXMFQqKL7b9lYVDFZ8IAMKwNR5krhSpsr8TIDkzoO7d4EDVK
fcxdoA2xqF7R2VQ4ZevdQEhpJ3RT7RNhyAa7K/P4HRBkCjktBvNeQebGZENf7v0Vw8JLLdkBPAiw
MljBQSurlz06+FPpGwtKjdiHWXtaT4Ghsw4MQSoeOnMvureFHOBsGfLHggBlXBln4nuPq5HO92yK
VpHRB3pSqBFoxhqiwcY3bQrN9lgVtP64fJI04y4GiVnQNId87EFzddBujQJ1QHTi0x5+ekxJmwgk
jU461MCc9Ecmt7kyqMN+rX62GVeLaxcSqC2hcLgPV/xK9XspDlvgEVGaRnECBpCfREGnwlM83vwi
7TiATUR9hMbiTdzjwiZDEDEfEq+ab8lBKaNs1aH/uDo3OaMgiT/VogQtGsH6Fzeco3hIVoYdP7Fp
IjT88nQiOCvN2HXd2yUxXECF2VO5gZpW17wDVypUmOgIbQncdrwddOHNrm3k6J0d9AKbu0P4rnT8
LAsRDqj8UDdKQoXS+Xq6egm4PC4O30Zf38fmFmg0+E/egR3UUHWYQs3kOm3jfs3/Bjwg/TnyF7iK
rpSFyK9pDQ0RSlcmWNBLfDYjCQeC//zz/1F8V9R7V5XoJCr5gB7UhLlcUpavRFYKWsYJ7qS8fdhF
y0UeA99WhZqo7dndpKzZOQzyN1xtOoWDsZJtkO0qDaEK4cuGNt3bGs5OJVRUVZVYrfsVl6Li2+wz
2FjCCWKk8KOQDiS1j1NcnsdjBc6HpjvVQ0rNu5Ae1DsOUZHcfdGSYJTNbnqEOA/I9rWCajbAsocJ
hjX9fuQg07l2rvOFexnJmhNJAt1iSm2as+HxvYB50QLqF8i8TNre6ahsFDdYZHz+3XsSl3l6GVCK
omz9jEMttXReqmu+MZzuMg7/QghJHhGqtEcqR10HyoYSrT+BN8ez3/2WJsVzqcUCC3kFE1rY6RxK
eUhs1ffs/5Uaxn0r5WpuFBptOJOPBQ46pSY+HD7TLnoVFoerfiood0D5ixTo6r4k3yl9KjzkAG1w
BMcxe0GDzdwURDImzapw80g9hmaJ4m+NwOovLiBrXvRabCjoAeM0+XQStUqZH/I3oLTbGbccqr2f
/7+IK5gMeOS7evg4Unkd6HE9bVoIZG59zYccoQzQlY4Sgs6mt4QyrSBRO7K51hUERYAB4ZBouqFp
38AHBjt72oACunhaP9RH3GX9XiHPiZN/c3zfEg/lne1XxzxS/HWUVTLgTVG7Aq8fOiEqt+oc+V3i
NfLV55w2ydIpheuIVXBPhveEi9fGb+iWitKmjNsky10vyorZ2Tgk7tKZWt6AKmvnPoAycvDNOxDA
Vek0Grm7Z+heuqEvlFAppUwnb2BNMJ0LZ8yMfrusUhTk4Qz+qfsh6YMPhVHEuPKLQcBknQAk9o7C
HZftZTyOQwzx8opYoQ0iGiThOiz8XP45UUuzumVDZkcK3cyf9LbePkWDRnwt8jVWOWOPztQJx1A8
km7GWhEzVWvsZ6VBlgdZKJl8SBiiSnJHq/ClKf7zOTfqYWvQ25V9T3n40w0UqPLcNa5Z4uUruwaP
vzDnRBj6hn3Ps/GXwoHv2zr3pCCxVTfKUeutGJA8G8L6j9gyCZpMBM2keIZ/lnMniyZpREnJjDRi
upBG0vB4Cii4fk3iQLORoU81cuevfsV0yvNhx62yJPYnsWnD/MA1QVoqfCvQln06Yv+0Xano3h5J
Pmx/Y8IoDyI9bqXk2Y7+weYVzmSyvG6bgt4r0o2LDfIlfnq+sqWgcmDwu3qd+peDiPzlVD7piGrl
tID1Ae4/8ICXN3csDUtvuNNiG08iQ9MXKX4qPpeuS2mD3Jr6P69WaKMsR/8I1BxPjnDG+1irYRsw
K/scDrTrQKmnwJy0+iZFpQg3I0vv5oNv0PN/dKLyQxGSH9fCOj7br6ewkCD2pboXN3quwFhw6n1O
aLPqyGOoW7l9IUPpvFu0AlsTPpBdu74l2reZzqsUwwvKhDxj3HpihyBPT+SJBqmQMZObDeQf2RYx
U5s7xz8zDxOvjDgnImmpCnQKXzFgcLojLtatmL24EEE7lWNQoybVAvELsm39frnFYZb4CGSw9U4G
mjpzw9DJkhFbnF3OtBetdCOmMGKqMBMpS21ZmR9U2gxCb2AmX+b0dIqN1qlHUTEWLHd311a+Wwos
+WRc0anN179Bg93iiKtqcgU9CF9gWu94b90TMwCyCfePHGAg7aCG6lKNWetVCc/uBk6fk4qC7r7D
JSh+R+L99Zp5ssPhTZNUguwLw7xcTDHmT70YrhySw43EhUpbSSK/rI9CheKL7McCsrgK7/2Wv0Ds
0i/2P9M0/UBO0b83KyslwXzQGgmufkWnsBCP4YQdARDCa/4/lNaX4UGBFPLInS/ZGaDT83uDNYIh
nEE6lIm0kwED6V2C75sTSOMCMwbSIs0c7Z7yV445mSOI6clb6YXoKwekNnYz/pPpBo+N/4UNe+AC
S0UzgPfn4DksOu5U/YZfMbUZ2aOAac3m19GyvoW15z8ElzVcbX7qy9Bh5KOw+0BI39SNMBna70GD
KyqXV6+93nFZS7jsLZ02Bh4+Wuky2AqU8Lfm0iUOZvpmgx2s5b2xvMH2OLdnaxIkdI1OzWd32mKv
8pBZAfG37e2HJ9Qf3KzRvYnyM2yIkjKo2rVgOabxaNcW9xgCUSIIfbJgHxgwbLshORw9QcZZsAld
bc1b/IWkVRTylkH8pbbTzn9ssEgL5OqUnAUsG8UN9gm/dONvqceo9j4DUbbk8GZWQykG/9xLmrQx
WOpITJJ3NcpCqNQK0aJRZeLdJM1dOIhKOdy1EOIYrIG9aDtDr7u2/RLSYPLvklIvPV93EOiZHphW
za8t0aoBcoreyMnwFhwzj7OuNtHk6iEib/KHW9ItsmVKafKlfqSWUV1hKBeqIyAyJ4E3PqRJII89
wxFoIafQxZfADkNQ/pS0OFn3PbBYO3tdL0Izen0KxoKweaOqb5PmqMRIX802cJ//kCbOOQDWB9wJ
MM446jCJwQ1J6MeW6PyWtKA1ZlCQ/Jm+hcZRg7WfxvdsgV14kIUfyP10mX3Z7Mhz4+Iixo+77CFq
VAQa5bmDNfaX94JHaAl0UXf5bWKelyUSt2M0TdwLD656MsFDw14g90uKejcK/OEDxKvuE5nNPQi9
tBDUbE0ruowu+zA+VA4fNzQSpEEfYTid9+9REWcqgwlWV3jE9QNpLpok6oSqNsuOiPwa5Y5MUVtl
3UTSEZ1VNyNCR3wAR31ceN17MTIIi8eEYBKcnWip0vDoNQOIA/Jd14/aIF60JlG1YdXwPAesOmRp
PYOQn3xHyCF9xFMS0IgE9bcLYbf6/g/mBqAvCNkCdhMmVgrUO4BAoEKPZvJx1dGuC0y9DvCocXvJ
b3Nw7ModIZiz9t1eB6wOVDYz3nSX+IQoeLrpXuOOKwqdpactK/Pn7ahoU3fveMEIsmFl0ShBSTAk
Quu0GRNphY0CL4ToHVGBZ67e4IhE0m1hy7z+DOOsT7Y+u/JZ+mNWP0jFRGcU4h9DnoUuyx5X4wMn
No6Q7xLuun82IirbGEreZcE+t6FDvFBBfErbuPboosdzCIGMhtvHFRkr5meVlIMk6BAQYbr5K3U+
NSIaRvZfr1f+E9DmJvPjp5HDE2wt+6nWH0FiAdghJzreorQkQiO+wQHPjJ/aLK4+rKZetPzS46wj
av2K5sUDKtU1uhZiqTQqi1jwk5XqqbNGRBC99tmIkCLefwUrG89F3ygklgMxHu/wcCr32Gb6xZbG
OP+MCQrN2h0ragU87nJaA2T/CENFiCGNbRXv2goJixK3y5JZdFnXUxGCx1wFYl1QFu+4UgxL0aJi
8HgXOuWVdOzgXKbRlsKBYqUUp/j+IwzfgTufy0tBIqVSvrqszPcVd0gjm9A8EIoQ8yvIhnKQyPoU
zpicNIiN2nW9Gc80OTqK4z5okVCnc0u/UoMzUYKB/J4QlPrleTOh2isPBDVOPqp6iDHbr3F+7aTg
hwem5i4M6nde06uhpi94AyWMcmz4VjEKzTBRfd2AEmAJ23lvFxkD9j0vPn6SvunxsaHBiOPpznFh
E2pDqV6wDsxc27hEa5RFGdBuDHosc9j/J/6Zq5itoqvgRRRKXJqg2xmfxBpaIMGT3rT2srJalan1
8Rz2vocTdDzUWBTeOcv90NdejOr7/qnGNH9J15xtJqLmIIlROvYWRnaopub+wiVu6Rl7vc+QEAP8
OH6b/bj7UdgywhjyayqMAAn8TfEzutWllqxldX94iw4Wy5B/hmTBBnnDMNzq5mroJdGqthKY4euV
ER+1M1qC6JokePvHUbedMwe9GoLNCy17YZE78G0M6JDUgsYKiSyinJejEFewBCsqwJeZv6E+2qp7
W/08s9eBx4wAhkWKiW5Yehxu/m7nq5EzVFZEASnuPktAFrmijZHTXENbZPer8U65jcDQyKZ6iV2p
AyWZdIWNE2xSZYz2MO/glzNN4onJ5se2cCUwfwhGEQ6+Io+7s53riIGdDY5WRdgF6295+NcxyMig
/yaVBWd3sMjWQ/qBf/5EvBrNv/7u6k/o0UfE7jwRzPGoCfO9+MQ6R08Cd3K3VXPVVxIVnJ3k6SXR
NEAWGipBJCKuBsCD8aXaQ6YLJZTvMtUGvZO6S9z0uqU2CzZnBMCGuev5WClI022amWqc8W7iKzn9
CMLPiyy8uXMn0RzlNz+E14xVPA60vrYxLONt0l7HxssZfGHYmwPsDsh0La80CJtJ8VhmrbbtnbFu
oVtLLUM70Q0S+UlByDFEE0gkSbAjvVvjn04LovGlgUeYRYHClWW182B3ImxbbzLFaYwRaqhn5BEK
gyhEAlYL4BTy1mSb/yjb/eZfVUqDr7c3p9D/U6VYNoOqj+oqXyVe6AKpx0K9NLtfHOmrC2aMnFXE
firn65btThdClFI9BRDIjeHlKdXebm5iNky36lED5qz3cUdXs78uPh2Q4U+B7u9kD525hHdSWHsN
S69NrgoVraiOkJ31qjkr2CAE6G+A4xIHBQqOVH1Qm59Syyzq3lnJtZVjE2120hCsIrun0lIlgoiZ
DSJdtmjICgdNWI9bx/XqaxaeyFRrTVFoUn3lJFCeUniS0lLjgd7llj3HMJBE3AAHJPVoFkvfDFtf
8Fjlcs4mOM9rc2WnSVI5nYocEF6P4VrtTs+7QEzemcsjWOq/bv1WdjWqdGuAdgr1JvPuV7CVYRt9
NvC3kaTaeaBbA1xCp7HhPswbfXZDmYLat7YUFJqcyIyeHJOlHIctPxopTLBICZM7j34QfCZ3l7Yh
sW2DxHJFgrwPapWc8aRaEWI5f7AY7tyXIYvIk9e9ClqZ1zFPuV9E5431rZ/pmQ4uRcjcn2GJJo/h
PH9pp+NFPr4mSDf5zo+XN1FwaRWPGKNghOLz9OJBYAuyVeUFwcrmju+F8vb5hAx/8ZFJRec9t9n7
ctm+2nTHepzFenhHZd9SOKBW85cXfw3fdbB3cP6eVqEry+T+Cp99TPgt+XYf9lQn1sz0lY37Rc/7
hCYFIlfc7GNQHJxTNYd7nCFleJBp29MdBDbPJAaiqguAE/cjxKINKBWl1OJIWqQsUaJ6hjm7/c+s
YdlgwEWVjJs8TajY3Nqf1QaL0NoAYf7LYm5sMWTxmaopQacNv9dPA9P16kHB+af8YZ4ytqWFk1yf
/KIb1vMtK4S7ynuIUhUrp1GWsBBDqeK8RCmmPJAHhAyTm9aC3du2PnXsnS5+TFYOWP8NoVa/ygWk
uejWjqMiLma+FcG79XTe7OFXQQ3si6TKsDQ4tIZi+gBgbZtyQ0h4Ax0+hRu4Qgwf4ZkCWcN2Fi2l
fMV2CB275EKkUz83/SMWe+8gKDi66trQnBoli2XEv04PKM3fTOnjbq7VuAyOwXiuX74QiRO0RCZp
HT3qUp7Cm4wdDjy/bp3vh1K4HP6245xJOpFUIJXXqvBEgIvXwNF86s69KOaIFb0LlKTbjAiKvjGZ
1uH8/TXM1ZH3zCxzI8fWkTF0Sj7U/lt5bSTuvfi/bWiHrn54HPasPARy5aiZODXXMDg0Z/FHPnkh
Xt3JVZm9hXKdCSAVlaACJFFAFwtbFLSPx+T2DwZCrsXga3HhTjVnApJ9cjGgpC0mcsWe1jzZh+yA
/IdOKegVhmbv+48RzD3f5SZZJ0rmD/B8OdhxGRDP3AesLO9BHLC3a5oRq1P4Pb4JDcgP7s1hnISS
fcagLJ1gA0QCJlUJz7tnBL73RmP3jcvBhnywkYcSzXNSR5x6Gs+28v2ReeGLzytv7CwzwZl61EjQ
W0l23UhmgCP0fd5LOB7HRD3uUY+sMbBhVhnbH2RiYY/rYfLv+8J1sxGzDIoZReTTxD6oB2bRr2ph
ttuoCJ01sss2DbwRF1AacWHC74Af8ajLolM5DDIhL6hQQoM9X3EPrVzeO2ARHZuogayu4b1WKKDR
hUcr+iQZXxj/HiV56KyPdJ82LL8ExkDsV6MC3jyxaaE8rxMuU33ndKoqjw/1K0d/f51kbJgpAugZ
MeSmnYi59d9HVAs3fGAufOFC5RNAE+dIPLW8bPh33KvyTV7SGwXRhhZNxDMApj7bAR9DMdQcxFZ2
eyObViGJwYj1f3VvCUd29IcDirWiL+N6fMwlWPyrupQv/kcZdvA3EwbMc+1/HUuBoFZwWjTBa9p2
C5cy9kqu9msC84EYtRlHaRqarF/Hr3i6uDX/PXhooXBde4WgtkT8Vp1MtpTarG7Y6lb2IS2uSDvN
45ZIGkwalnpgxXY7+P4ezEm2GXHQUd9iEleLOAUBfSnDujohO9N9N/xQClPuaIb2ft1LgxdVM2Kp
xzx0eyK6VXXgp+DvTCaXRXpzxuRGr2GCixfVxRCNo8id48DFGsRTAHFmhxCrAN/KkWvIY31T6mNj
vxZtGw2ige2dIuIzigwRXgSotXmUi1GlbMjsblcmTZ07v7mRc0oIk2Yp7ix+MbF3nvp3uP4oW9uA
hXhnADklZp0Drdw3eFHGqWQG1EVFlJNjb7BDI0Vj09aWCBm5SsmMgen3xm/9jyegeMlGVLI4T4jA
tVcO+Heci8/YJ4cZoqELLaGFSZXtNwY02rBFZ7KenFS7IZOJPpv0vu5t6YIqcrhiTkbWj8erUFWn
D5jtpxd4IEG77dOwKuSnOMpihR8h9dLywya/wc/xIhN/61LUV5gPeY6KevwP3cV0F3thFAwmrsMM
JfifB5zFchtkEqFvLYCt5aEYU+2OdzZ6BWqE6eyKKGqE833UbaFlCqdNUdj0P39PIYd6ZijD2oT4
PQG/6wlHfimfQaGR2AlutHabRjay6JO2uP0lkqlzHYGKUnb7BKP6hTyvqarzDhXgu0bRvqCSJxE8
48ZYPhcdrUAA6KCkDvZ0Nfp/kjtk5RcxxhB4MIoH9ebKrXX2Tg8RBr3HFbCxXb7Tnmr/KP2VfaeL
qzAySfNQR0WJodJFeMKqLYE2xGKGbU3Re0VZaqqaOy3sk2zYzg0eempPoiYrsEG9cQfW6A0Yl/u+
x2t3UsfkClAJSYM7Nv8RdNLLFRa3Shn+5KDiHrCgAwaeegt742pDujyO252zxWEUvjGwwy3h4fz2
FNr9D7ol6keMpIR3BrtxzrBY/ab8k9tc0vXvjo/HwoqS6N0qmRjXmSv6+ksCt1Qah7KHNKJ27Kv5
I1ltaWoHFc37I+lyI6fNThngYmmFjc/H2tqlG/qU2ST3NOnkGHEr/qwdXZs3S9zVZ9h+Qvfe0X3R
jlyM/pjBhtwaCKz1qwz1jRc95x7m6GdwiVGkJgMKeHpT6ehFRUfd/koOcYGh6bwesQYpDtb8R3LR
08FM8M79LWFM/wFdmDr0gRoKhvbd3ok5V287uTE5hgu4MF6L6ZUve0ySbSbI555ETIFkfdQ4HpPY
PGGjZ+FoNDGoDDXwms4jSlkVoXaz9K3kBlX/86lkwBVPu0SjCWciuIr5OHLCm6HHFZpc/nMaHZCB
BUhaCOfgnntnidh/7ycvTY7d4bt/W/Pb53cPAaFM0tOskBVqXhgNBlMpNScfvd5br7mnTMhR+KM4
e7kChYywXP5WAjN9NySsj47r+yMWcvLWAZIh5tXZqsPHsaoCF5d+gR/x6v2eIQDqwdgROh7Z05VU
znwc0AndRvtbMtBRVY09WGnfRPv0Cjp3zns7HFk/4LaCTD9Hdbn0QAVdViikSxgTmkMx832kwSG7
G+9lxKq/XkeFJG16BW71pKlYxdM5XO1nzfLFU2u1bLECa66sQ48SqKlgvED4DXo9MfOmDrNtRa5V
WazOTAnKEV1ldWLQgI4Z5B6s/eb44tcjJjxlh+pJ5syjFbMwXFQEdMs/SKpmNKDsOepZN7urc0L7
jL5sU+ZAO0eLeKB1WroXKQowRUXdQV/XseTjv7HmRt0pP8pS6pLZNR9peo4K6qc+l1tyUjsc0yzt
ICNanvMKBmOBc19jJu2jhXSq331MDj24TOYbWnsjj2YAmhUYSfg6G9m6bofh2jpS0oNDwOzMkwOc
tHAQYRwVp1BKy3gc/1e/ARuf101rjPScEbIBGujASFwoWw5QbR8hDxIF6UM1uIgwzycRUHAv7McF
AFCJX7cTjWLJVfgIgVh8dZBdrm8nfRxL8x46FomCzgWyNFYlVhCLwqWp/md6nEh3aECzX9rjWE17
wpMMp3EzvKTosGwq5Lsu/9l02Dhj4PvlKNrWtF6nANUY6qh/Nh5x0pA52I/Nix3u/mEc4f6zBxBM
SkVYnAf0wdBKx/2QQDNfFFK3J2T5uybBHC5iBhOJ2RMfkTbEW+nDpLMcJ8uhdBuAfkIAtwfgG+XI
G0WDZMljzmhv+/f5ilK28tq2bI+KdKUPA3gXcAKWoU4vokvvuINVprnWv1Z9o0SfzTHuJ3NVKm9j
o+V8AxQNFEv0BzMv/yjARR53bh98d6JgqFFRioumv1PRMVLw20porLZis2+1Mjt9C+RcNKRebZKJ
hsJkbT8wYgsZqe8q9evxq6snAq2pgAEREqGydteJS1pPM6qj6ElF2fSSlmsgU16iQcvfn8Sf7YuE
G6oTEePziVkJ4BlYEYkIXQHA9UWVHwp0wj5/RXWTBCmacETs66IDkJMpcyV0NHY/KLdJgWRcS/5y
RB9ZlmyopVL69IFBL87Q/+LG8sc2yjUrNvTQkFzIT4SZtBjFfy6CSYM2F8Cn5UNbBFXw7jWZ98Xd
v6FiRYHqKnIZGJJWhlG6bpn1E598oQow2nu23oZrcn3CcezA3u2ToJ6GPsfrSTZvEWVEez11Yzsw
gy42Jwtm1dzl0hRu7GkUruY0nXwO+Cz9zTy/LqJU0z05JTEGufxG1WJdPXfVWJ/Mj6xWAHxIUeXR
n8yVUw17oq4tFYU4UhvO6LMDEI7E2uR2OPh/tkMtq5bV6EzwIBxYF2ZjcLz2c9FCVvho2ZZJiyZR
mOjarqjoiO4FdvkHHYHLnrNjPDnnZtu1xfVDotNDQSvAVKoqeSz8s4BgkghM3HpLFUoI4b5KN30H
CaWu6POKx5C9l3qa8c25mIrtxDhPhDn3CqCkv6ZICABkPF2XtII9pUQLLXNw3AvzOzVNClJwQ6gz
1pzqfjXrklKv9rzoeMP5FNNfaoPxpdxCNGLj8nSVYgPXUPccxpGLu0LCdJD2sw/yJXRGjB925s2Z
A1tVhONN7e8n7OfaIssdR94pm3h2SVE0ProSxnRVK8xS4FXEsZ0XIj/xJ53PrIudzu0LakDhO0av
t+lEjExkmfkRGZVBzkrZElqt5IH+cqs2wApmyrRo+pTbJW6rPWovqV7zfSdP0ByLmXiR21vv05BJ
Drcif4/II4tvc6Nb1CM07zxVqP/LHzM9X7tFtjNHzWceSZaZU6ynz7o0nq0TgSV2DOAIiKhLiZZj
6pYBrJqzGft9++xKS1Pkc1kFaupfFadfrgdNAX7fbfL8ua3F/AdXnDP8xm8oNQ7cpeui0B43Jng3
uOqMLoEe6kuXLZQRMvNI2eTfRE5J0p/6gOiDB8T71JL19EDOmxxdYTH5hs/6SGAIlbirOCiz5tOR
9s9VkxQ36qMq3XhBp10PmMIm/6UOowXXFFJ+SZhqkjAeD3TpVyTCaz+8dD/dDQNyRkINlemXfmku
iQAQgxMJwdwRU3bMnQpLobtqaAU75Z8/krhMeuikE1HrPKFi7+GODeH6kUkw7DRMPDuoNMKoizqw
+nNS3ZbJcobMSg67dWGG9N0rpOhP53k/p/+VY1t7j4XLtquhUyc9JhlpGeL3KlzSeQ8W7lVa5p98
dv+QmDTP+ZYamC39PJdR2YObUPm0QFH3ZF0eUPGQM3zmpFzraEvH4Q6LNPT8f7BnZkze4kmLjbfw
xA25ovpjK63XsdOwccWsD4LbGJNjNQMfJvkM5S/PZteUoOIrrWMCVmk+BPmkATLqeCscN5cRKaVp
DFfqmr6VysiWu16vASNORKkIoR0q0yQF9ubKdldv2oLSieGFB6WCkyQz7zQ4eSOSebud5vyk66+t
AnW4XHe4M3T3dAwcSBZEuSscrWYi80XDMX44yHVc/Lc+uiPxMCMA/VJPBJTq2rwmRrhjk2cAqjHa
nDhpc2C1vcLYSaWJPCr7HcjxI+j2CGhBPnBYAAuTBeZuHWvxn2+mob1sReyZrHVAYpgieF1IN+sR
YKncH+469odbsPYHZ2OXzP9nmkc9wXr9sXd4/EyiAXghSy6Nl7xJvO0NaRJEbVx7cXfb529mfxAB
wWKNF/thnJzFRKPO+G/bagXl661bIFFkRRay8o4Q1/E2BQFtwSnwWzJgI+iwZ/wEfebyR4K+1ETP
F9rUh4i4+hT4EJEjHaX4V7ZpF0qRBzdMyMUinvjMLIyk0Iy85DEINsUNN541eRswzH/yx23TQ4Gz
xEkh+fcRTt7Q/joXDoGfnQEpZFxBeK3axhNOtXvQR0zuVEHkLsmOFalLPqi/l1yzwOjIRFu1CVTI
ECgAVODJNeYe3R9zL6CQLey0u3pGVRjWIJS7fx0aOa/zgVu2TKT7bAn8L2R4nPRsqfpFEJoLBuuq
DRxyldbQY+/IREc9PPUiyzhht92R3iqBpnfzmsTCGYmcIzLkAGxNbgQiwsmzydbuIT5YrbZdNqx/
nma04uJnBBY+3jr35yyVjSSwZ45xz9bVHqgccsuMiSxuvs3NRAiuniCxIuHazik++Ehtgf20T/wi
6IpGbu2Crjeqyvw/Wgv6ExV5M/lfZZjzOtXl34WiSYRVDDv27sKvPW3cqWCU6+TM2pGE3eVdR+sG
BPhOv3/3+OOy3geOPiPLrC0v90tXcuOps4WaZHlN5GGzXC6DYpnBNmpNTNS9vqXkv6N8AgHcFkc1
kBEPqbrVAApL/nYh/7BU6/McPUwXurjD7+vPRMLUATprCmbaUvrMYhLAc0K2TY+7L0aqJTpz4Z92
Lc9crYMOSZNd8jAPQMR9Mz9PkTWEckZvb5/jJEurhCchhSbewBlbW6OA6VHIq6EjYR4Tr24DnAtT
1vwyFyH9RXfrKG+ENVelE2Fg6eurC5/4qoAvi9wBTLYomoIkXhxEoOHV01MbWIazmgUh3vZCRh39
XlF6IxV3ixMUu4BA9/pHw6HYzoFROE6QHyAaQXqydyjzbQZ6xu3Fbqw+1+9Eis6c9oTrZnHLJILo
5x3ET/XltYJcRdkqnIcHd6+I7yixy83JvmMDMxxiD5pZb0oMtrf/rWGljRL4L+6nOHj1ca5njuUp
p1ro377HYx8cImFduRjgnEBA+7wru1hj1WCxyVOvnobZXWN3Pse+h0oSlcGly/eyoelYfUbQbaAt
VuUeVFqnMCMRWNv9mxHb8i0cgWuw3QQsdgfBMxLT19VRujvfs1j0bv/Aup5Q2dNizWkYmo9Dy51W
NnS7nLx3KF1B0JLEKUl1gaFO2GVHKuOwKN+5Axdmum8uc2zH6WFTc4d2PR3W+nIGKeo5ZdPnwqGX
BC3WFOasM4azt11Pcwy4avZeSFGPlLvUay9DiY1OjlbZph2KfKzGHRwhL0hZOQUIuSiYTyh6Hi9b
oRHUR+S9KFtuQP+Hxf3uUpATx4Nn3QiL3XKrg2h6wJNspGxnkemrHwn7dHCM0oINW4miTHfnLeSM
EuFJPmEbKi9d2sW+Qz6sfHV6i1k8MJyvOKtbcQ/UySXURgs7kpUhtyrDYGxqau/0U+Ey3GZmNqnq
Bn/tVkGwKbVMQVIpPd/dsY5wfzmE8old6eCosPGc9j+rRt4hbZqtz73eTdw+Y9w84gnJ090Y4wJz
dqKen+453BMGcCJIif4rPHIiaAtkXzmFs5TptSG4ht2tBzf1xZD5FJy2nnBaO3CghEXk8MruWfW2
CecycK0veTcKTaFjmZD5tGTWjrt+1yDHWnALNopGxVgDxvcxB0UseR7pkisbbU9rVQMDLHjFTNl5
/FyJJGWp78e7MMKXVpuuiaI1gQk5zVjfrdufKXHkvSxmTWFDu6EXVA0dcDXXH+7zpypYTSUoMWn5
T4VnUUPXNnX7NzxvGhiDYR88+v+ibknlKvEGz5ofK4pV0J04B/W86uKalLVe1X7nPdwgDfp/75xJ
gcaLHbk8/kYTlPtac7E8m2H+tLWYemEx9mkqwgqJQ0mnCvFIXCcJsshRqOuxTRVVtkTf9fjVDIdn
l4P51vNgFUDcet/VsFzjU3f2AViP7krl1waTllrEA0Vf7bMvBnMgT/c+KtEsgPOv5of9b7hMRG/c
bTBogUFrGNj1KKvNOdvgt6mhpabNeAhXSvrKwZSKZTL5l10IeV3AxvGqTFsMKHPHYrt5KczoL3d4
hOFIjTAxqyhX7LQ/0jhKXW6mWhRfKfgUUC4jb1wOCtPnqMGFvX0v6wKYOXCsuzVMmSMBuBFGmRC5
rbi2Bu26ZCy0K1+ERbTqZbI7ArsiYdb36SysJ7kaRfRfxy0Rq/T2KP0mTaqKF/b+zGbvrR/3hy0S
HDNmVX6SuYUSeAQGhcrGEnBrzLAJfG4a+K/1tqrXyI9vnBARgW+bMmc79qjgoKCAM3RnfnR5/P4j
wthi4aKokh7ovW14lzed6ZlsZX50tdTM/iLCUQp85Z8IHTBbxRMRxrBoZVcx/X6rrfmGfOFOjscJ
2TIda3bcKWkuLZA6JI+Q0aPJVQnT4LIiXBRxGuuDrbD4ZlKHRU4ZN6Qw439vYVV3NmMHC32m4CKE
v90jcmBkGvllIn1gg2OXV83a8ZdDpaXZe4laM5VP+1WYi+TUwOVQHxvAUypyuqn6taIdQo12RFlT
xtnBgOP/Z0wZ8MGoQiPFd2dCC/OPJarb9P6HlnHEUkYJVhoz+TKSElSQjNVwN2OWJ68zalsn9A7B
DCTeMa5PyLRxGNhZsiqu2U9s/HC5wd8I/ZCcOKVN+Fokdx57pfaaCy7BSFWyUi6Ju7W0LOWBcPoD
4ayYLxSN18D85jqYx/eCIk9fe6xt8EgvONg+Xw0LDHlRIPrV1Y7YnI0kY+EzflOcy4GrSxiw8xwo
LkjxuhGhuFkTzlKz30g/ltyWCPkikQqEzzVR5Rm/gDVKjVo49o3Lpcvm0dtccxxtteg0Tg6S/mx9
GswyjdgEZVn2115ugo/1glNtnLEvft1Dg0/uPCazffJmFmcupMudYGfImwPa7V3P6DMYv7dRQgst
WW17+TUrWeXilLPS0wWISd+9lYSkI3snIcZwhtT9/ycSzvbL/mtIYG5JPhcsQNO0N83lC2IkOHNj
s4f8lp9XCVBD5N6OrlxC+2xoCfyp0qWu62vLNnhytfo9MRaqucISM+7ibiZYjocMVbIHnolrhKjY
7sM2tWieZ8BSsPNXCnSq0EP5OCwjGQNobhaGZID75AqI3EMYW39GC8KxVeR2rBKTk2rUJBOf0lul
RL1JPaebqhkEvDANBC895wc8x2asECuLfd/9KIxYs0Iytu67dG8MKcWT5veFaufCjSgDBV6Hy+J0
IhHKYYo5cKRIU5HkAcs9ReGu/X3eN2Iaw0hW6KS253DuuOLXGPH+ctpmM/KLh9V5XOGBlc2SSKea
UBYGSWfXEBHzcUVozGYX3b7vkxeLwpIc4GCvNLtIAS7a7R0o1UYhGcR2faf2XldopzQ2vo3/fFHX
ODfrXs8cj1hxW7x0oP3st0h0tVLww2Jsd31iAsPgdHw2RXxWzHi/KIQqdH0N/zdisK3hzQNji6lw
XZ3wDlYnztfpDv+v4uF4oPSttl5CSTh5WgQh8wHthkxyfs3JiqDnZCSwrJ6qaPwi6MtRR8FH70Y/
XE/mUJZbEXObBjxSgZ6w2JN9M9qv8G0lO1GX3meROWU9uBqwvZ9X46YV39j6HzTGCdViaBegIsBL
Zmqi0XA0brdtgK5p0yKtFudtLiH7a0jxxU020CSSlKD56YlwF3JD1RfpuCA3J4sRdgf7zAQIhIL+
63jRTY6ANHJXDUROUUjcABr7LDvJKgFswWEZck20BzjHico134TbydXGqFJ7EUW7xpW7AVxSpu2Q
UTHJDxkUJ30rjwn/LWxtRc+/NrAf9VQW3ArcA4Feu2lFNAbSb40kmr+bZ3g7aSMu9JcLzn7fa/HB
JGa8V3FOD0EJBtT8wS9C37lQXpBs5QYzD87BgKk3++MlfY6njAe8/KnFlhwwYS89xPXSGP36851+
dzoMPWIbJYkp65SqTCyJjQbnzYaQhqtJCUb4Y3SEtN5lNun/oIsm/8VEyYtETFnJMoSsmEi3vbUW
nOMbwneLA7VFsSU0oa/UNWUXrPjVzTZYuqi52VvHciZSX3UzFQ2B7yJ5FjkZ7p1+aVLYJfvUFrug
RXX64lSN+Dj0c730IPZicglLIBrYtkfxzOwwRPTJRcwCO68QSGzmTmIbg/dKpoKGbrL74nQdHvAL
D9pkk1HHcuagAYEg10QkGrjxIbo8RtaNR+mwlmClvdiTYamN34weu7izix4hqc8pKVTj2i1B44SN
qZtDx6d/XCHy1X4QIMK2KMpHLkcvoBKWpwcjWWq9p3msztsXkgiROQvmVprI240ZlLtvFqWYb1xY
RNqKs9zR/Oid06T9IUYlWEeYelMAo5P9mCK/CcRErguAFrksnOMHkPLnElc73VUpaoBP8VLEORSP
YiQzgYwBQqH08XBU1RqsqSsS6TN9/8EaVKt1pcatVAwGlM7mZj3uJ8hieRQGg7XG+9o0hmXTX8OM
uJupsNMNwU7q8jNibUMdh+cdGzNeaJbQ9ikr0+Qljd8A52Cdj1OPVo90X4XtWYRK8z0gbq20bPVO
1RcNbj4UGFEQN8GhAONOvTcS8O33IfomGMYOqrJq/Bz7/NYqwztAkCBG5W9JVho+IvAzr0nhlNWD
X7eWItiNEEIgoj+4ya4PMiSnAZibMHKYoNLxCGVppcNMW8HBneXttoSWQc4PUuJPSxuTnO7YyRKn
1q4IZXFYtvSji3YQ2jPo/ZOyti67SH+M6diSZTo+36gai5ZodseQJ27ehEljZM6nWH2VFB6+mVYh
T/3GwcgyB/hPVtoK6oomhZc3fxdd5ZyKsoBGbNYLCCUXu4D6zex/yJ/4gHDtW1bqi1Ceme4LlyrO
EaRJqO1Igv+OAPwwCQ0kgKErMvMcJuqf6d3UxbF4cxXUsRu0fZO8DnUJDN5WbSY6cpga66n3BUPB
L2ErZJD8HLYKqID3J76+WvTNszrzSI/Z6LqOp0L3izgwpi+OfiRcK1nr8PZ+o63RmCCebQLm76Kv
oXpyVjHpZNqVlapOlUQb9vQ9oHKtHQcgh2lnQRoK3xAUEJEVV/SmFIGJe0ELrSMOolTSS29++2Hs
TCfPF5abbkRPYluYdXUlCxL1JrIG/pR3AoEuHMbcjXEqCSR6G2xsEGgXeCJhdgzTCD4E7YuMixgI
6pzlMWtvymwEzD4qXQ3WfdpTAnfvZK14uOZrvUyW6NPHLkansfC3vo12Rw4/AMnNzOxKMKI9iCxY
xraFV1edmCmX5gBAawQW0IsQyw8yt5d1925CzjBHFpdDaJNSWBYr3vuw3CQzQT/++Hh0zFDnzd9W
p2JfWkPelZqGWLUyWHtcUHlXHKsIonSqo6tTSWDzIshTnKRKwl6bb+UULXBlC+io/azf3jAJ3xhx
AdjfG954VJ0ZrIHLR7Dw9+b1tZ4WceijHsGrerOVlPwqQIwnEY1L+HRQ9O11SZYHJKrkR7eirKmE
Bl9dcB9BwmVuYFGyu4flutBSprxmYH8D+K5wcA+GlIPRIO/mnyzx3lXZgOIuKHUYeu4GF2osjfKU
jgo+suRQGaZkd0kWkNL+3gMMJVoj/wxyZodzzqhsxrmizru8PgK+1UVWwdJ+4Q+voaFILQ9ftk6l
uAIVEtZSKJu0XwpudogYdvWZI1MWBaZX+CEdB9jMp/Gphv973Us8e4som6IPEOXiqNOBuDxY+zMX
FI6vBJ4wL78rBDM+o7K+c5SbDD8/opKWG8W89s6y8qrpHF7rViRwOmJ7oqiriPxt5rogNEVTj/o9
z2LuIFvmKP7XZovDSWjPnAQb1WhtMzghVau2lgwm8S+qO0iB04qiPqPbYTLo0XnDEOl1/ROde0TN
M44XEyy6pp6eX3s3Ev+iTFT/O6I9veuxtVmGkqcsTYijbeWtyO8ErJ0WtOd55Ulq7AWRqYfVMUz7
ZSSZy/qGYq9C7DqXZ4hyVzoiFA43UTlt1Y/At4lFlFUsOgy5GqAUaq64Wk2HhqpdBpwyIUh+uA1P
0JQBAI0ERVqKnC6qwG4YNq1QuLcrrIiZ042xssYMHCn0a7KoKp/2nESldmSkqYI2aErdP3V7H7dg
EhTzOTGLLby900VxoI0kbfjB4U9o4doBz7gWgOZ5OWCJnv+fQ2KulKft0Koj9NQ1yGjY2vJgRzwR
WkqbyYgphZseQaLBTqvHyrEwpo1g4cbMgCFbpOemAU6dF7mCoLH2TdnbTDEJNJ0qXy8G2lYyxd5P
sif2PZDg3mkvbRDhvLo++dccpErfcBz+ffS2kIG5x6G+dRRh33yY1HzWlk1OVPYTY3KhjNRSRIGV
KoQoJE19XRIzS8h7PG2GKPWMTqoDgXO+yJ9cPSyCNU9mRYeItrUFgENFjcNrdWted3QxJ4Sl40xY
lxPXf8nnz60S/jneeSZ70lqJ+xMagUmxOdrE2IrItEqSH06vEjUiN3rZnOSiTUNvn0NxC5bN9dh+
dy/HcVt/XlXLPb5PAkwqP6BNHcdtsS7JXww1gjZ25+5KECZIDkrqzR5W8Nt6C0onzkuckWxcFWuN
B6GgnQGogs2/NJJMMEXUmK08ef0RjNUuRP8Xgecaw9xEpacmZgCL0BEa0V6cVBGs4e2k+jRBhx8K
U9wHVglIP2YzBV0I+Qiz6KEeOH7Mw7vIxUXkaqSwklBywgXn6+vilBEI9rFiGk3OdhPfGXQJBxDL
iIstgDZVZiB4AqWsNvm4Tvz77nRv3FdigPGOKCyClT1Ok54Qf0FBqCEyjfkE3LpM3StXYykrrFSW
su7G7eTDgmPehdH9hWJBplDUrFOBP0jxy5NiNst1joORn22n8eA13iIvGHFrv1ZT98GhYVPUu2s+
D7iYbzBa5CQQYB/K74siqquy99Udu0UNoEe5ICtCbDC54SxBgDhGkO99Tnqe/wpCZEQgktLW2qPG
bmchkjHqCgkHFB3t2W51ZSCDZRnlPgF/65DfM4R+sDomowxbOEJ5pLB81gIcpR2Pu2zgMcpieNrv
tsD7vJFYT5tR7EV9Mlm3VpEcAFmdGGfSZLYSaNiw1PHxwTIP7Hhkv+MH2q+jl9Pjv7GKSR/RWqEa
b6kvjBpVl946P07a/KmGHRQQCl5gxZyXvKWt5UvzPmija4+SugS064xxn1I5u0FW7ZUzhgQ+sBwp
MTaRxCUPPkfolTDi2qYK0Pp7PXfsZkZElg5NaXxiR/D4RFvHsNG41Ud9tchJ+eUv7H3l6WFl69Cs
Rk/8EQ4RJwstQMONGktVUQGoGJJjaRPuCsYnXHQ0db6TJNqox9cMYsR9Ns3C/598AOYRN7fFcEht
hblonGo2sYrt1PJUepZMcoZIJEHrIR+6pjcb5XK5BBIrXXMWWvgMqhvZumqUTWgKj7LNy9MBwh9l
Sv651AurLFV9afGUOZnE1nHlZrXWA7d7ek4uT+y/c/yLjZMWV/rVzDemKw2qekJtZTw8JEPxvOwn
V8uxukhxBGJdrHxsP4L7gM/rre3NnaHj4rkOVARQuSdsX48DJHgFK9Y7qRULsQTAhFryONwGeqQ4
P1NByKkkkPhiqYG/+DOjbSsHOarqD9emmQ2UMMRyr2e8i1zl5OZiJ7aXbdVAB950+bGxA7nJrnR1
vdr/BSkhLOrR+fYKRCVcEc+vZlVFHOpah7/rRrHZH5fR3PGN046M/c0n7MRrQ+v4PhEjWK8xUXGI
bQ/3rwisSJvzfaLQIvtL62rAhai5JzG3Ck3gu374ONCODTbMgrxvWOEvflgsL5f895R57UL0E2Pg
+XD2u6KDQ9+dEgfsrS7D6uELGGQIyzoXy8YRzoEQRIDJ6YKKZm9VqHb7gw87x8SB3RFo2/bTssBU
FSit8ey2xeqHZJeY8admjbF9t8kPpZeHbvEe/aAAZpZDdYKUhGI6OCOOBjeNc68w74rR3Gmjo/ma
+OxOE7agLZvt6SpShdHs4BdEUke+Ly/kg9D/VpzUxSbl5f2F0MKT/FTtC/zOV4Q28piAqfvuz0X+
DrxAwn682aMPifGnhyVNHCVEDw3ABAnXCCYzLpOSK8T8dgQD13kumSe/WcVJ2Zr6GNfsVewkuecg
zPWGLpIzZ6c9woigZUN0UiFELSAxSo3tM/mw8M3tj18fTsHEamXMv+rHFjDMP6rvbVT1DoP8BCyR
syo2XoSYGes6ZuacX2+kZZd8el199bP8slFm/+fXkvbPEgVofGptM72Az4UCgRLSbRB4g/Mb3fc/
qBNNgBFJZqo+dAyxUHPhaBk5yqd2fovxYB8Q5LB4FI7It971dvhrEgSJ7DtuhNmkkSvfKHoRE12K
Ir8cAKUTxuWf5BKd16aKxANJd2AJe9bwGPBdBWglXsWSIEC3p+cEOWxnMvmHRiI2FhgogGc1rQTH
hFRw+RM1YoRtjJwOCAos4LOAX+rzjhfAku1pfO2e5+OAuPAmoav177GRRXzXHzeJVKGyEnK3p2KT
4c5RL8PaivQq0yBoHgUva17tzaRBj/96DvEbRNonG6otrOaVthekpYIacfp/jCoGwCbcw49cZasC
yAMT/rDoAnQa3U16aSrNIaIqpwhYpFtO06bo6YAdW4yDJxs/k26r6TBM3pBbSvOMsqo10Hlh5WEh
pNTLp274Zab9kIktwjMy8fEhspD7pEbjAaooImb84GnP664vZoT7La8oqX1yyDN1uZAB60/yTNPb
4EIfkf4f+Zy0Ljm6Aue3/eyDCmkd8OSb0fAaCjNuhYtALgRFb4YmF/oqsrpcXIiPekKb7VXgppRe
NXhX+OpT6ttrDwu322Vucuk0Mb1bvwL0NzMnZWUGf1brUa6r2GfwDmZhS1V/0xYDndTyNDm+leSi
flTh1Ixp7usQ2DbHhF80elEJBgcv2PJWD+4XF6yhHvK/06M5APd1dRYoV0/6JUpQ2LiYBvRy4xhI
UA0yaayjcLxtDHkJeViTvrNd1+qBpxDjScOpqs/i8SCBANkUcLJCt/SVdU43rKq/M/rPgpClmSjU
sD48IU8OeuEpT/cMC94eHuAxf8OMhWnmVj4Jj3qyHmwQ8W44MR8tLt7o0LAnCpR4CpbBJy1U4wq/
VXshtGIKpk+s91KSVStZMmChV6PjgxDlfEfr0rCvv5Y3I/c4kPUKa7rfPgeSxvE8DVPjDYPV1AV8
fO97WT0acnVoFIBpzVHdFYQqycesaq29EtAwSNYLZkSufarAWEAnMD+YfiSwMcIpr0tc+VYQIEf0
DviXXSLtxjtDJHd58HDV4MSBPSdlj0BKtjhEnzt6cw54xgrItF6ntzpryD+mrY5og11IoOFoCFdV
yHvrrpsFSRwYEIENds6ZXSRQq+rUPp+2LLz8YxPpPJVi9AaUvtsmDrMIPhIPMLG5B2+r3lZCU5tq
TMEZm9MTtkxFHRREhWfCQoge0ip0636AvXdfXyegiwsP9nzkOKjTC1kP7K3RXeRD6q4VNw4DkfH5
PUr5GAbVxWmn2L+8sm+bxb5ENkhYzKBT407gCeQGhqFb/F58k77p3HjTeDToe48KVMz4x/k6Mcg2
aAGlTEWi1xtnsHBa6Y7xnQNt0H+EuU/RQXDmrmUmj/w6o4yG0AUOMyEqXjyPwc9SKd7TwdqILCer
hOKoRYpllk/CZX7eVmMn3vRamXji0K0mMAn9mNEAvSb7qSLIX1kWJbspfNyKMeSgkDDk0FYU7y3q
WUkQnXWFZJl7fdGUpME9Oy8+GThQfJ2YvwmQ3f1SjkgS/9nghay5GN0s1FOhRk6790b2oB0bCaQV
u3OT5N/Y2IRBL9DdUDw7PA0MpjEbT5HMGzIQcdTROMlYl+6qwwMYsRFQRRwnkHCpMIyczTtcILFa
Z2pADlTc6J1ne3iuToFG6/HkEQsNtT5Rwpij8W84jU4igwaGJtIuuozqaE43t7Nmcx+ewC4+8HiO
7RQ9xDamWnIeBL69lBsB3NmNquSRcG6Nguk4oA70ftqgQCGcNUwrG6tdDy2oeUTgya6JaBwzthFC
d79BqyKyiL2ssqnfmmf+CvRPSMxvlvk/kItc+26Yh/4m1477s8yR97qzXxLMRUdal3GrOA5CklRS
MZAPZnqZRJTpdXoQv87/YnE7z+QoQ4OwrG+sQ6i8+/czpm3zqtF/0xlz2eyxUg6Fr9PtmyksL06J
jGM8mG9+XEV9W3YS0ttMlxA0TvkLRUrG5pbhsk60DpDzGhSoQdF4WyQeRnlGwXM6zLOz7CdoUJ0z
HXhyvbNjZrUwyqYqnES2UKohyNn9C9E/EcZtM5jtHG6nCLpfAaUwsalAR4jsWefejy4KuAqBXXQf
omP/PzRsjGNab5wnvwM1z77747EhjwoM98CEEV5UFh6oE5zIi+mAp4vHFJ/nByHoTFMdOG2xiJy8
ZQBV+k+rEcM1cw8t1PkekSBwq8H6HHJXxQKMpNKoLoIJPDOU1fhl4lcr67Zhj8/WFjWgEgpnCGII
fyFuz+8rd19rsG99rrJ6/GEW0czvU6luwImKDA001ddqZdutA9WfD5/lLxw+23NQ/2m4nF/HVHOq
ZVyDjLhPjXRHHbcXznwHnXpukIR7T/uTQgLzG/KfUEf7OUukcgFyfPiRu22utBEdgOOmO7YaRdpb
ak38a8sY6OMqWISQ8C8niOt9nsO7W/iA0hoaHEHg7oNGbkwxm/P7K2Tz+I/XM7tUWUdwFC9vl/bq
c4WUhk20rEJNKLM+PvSnJITL9Uevcycc5Op5UsPOPiYJbL4X09LaVfWKCJ0kqiqTC5U6tPWW43Bs
JeAUs9nmWeBF5tN68Qsste83ermErZ11rgvrW2H24K6J+oaoL9zzcA8CCIYdqbFN/sxMEx7xErpH
PpIhKV4xQ7AObHH8eWqv7BbW6a0vdl9eg+/FljePoYLIMOio1h06alOeD2KAF0vsC/31Rv0jUXtn
ZuvDG0F8T7Vmd1ctyENTMYMI7jsJuMzyzM0OY2genj72A9kQcj+x8cF/EBWx9f82zyLb++Bs3g+7
8Vm0RRV9svVxiNqko1eeeVKqGv655FkGgo389JO7mQ7GoosnSfs61yRMvYROPJ8jizezNsurcjfn
CKkK6TDkgSth+i12my/E+OzFAZHhZ5LPvrUlTRf5SwuoVnzKlMKRYFJYFNkeOytX3NKUaFO/2GcS
W8vfdCu0LPXk0Wmby+5PIyHGpZzizdUSlr+e/njb6sDMR/CkY+R27Rrp5onN3WFjV6iTdiR22euF
AQVCJu579mCnjLjylAVc6Z7Co2w7h5XzVwMTrvlw0xLeEeC35eR2Z9HsIppMCnb/UHpgqe5un721
hj+A/LKmKCE5w8bh4KJyknSqoLpJfHtXKzBeeZv+aoDzLB9/5zasCYTLhJ370SFHgmeldqy1Sxlb
udyqASNhp8dBRMPH13Y2rbihaLijTQyO9R+Gkio4aLNBpLCiS48Ly7zW7P/RVQXaOJgXVfkTGbTO
btx/RWH+uYgtBG/fEQ+hJvw2VWZI4wL+mdugJwC4S6GE31A1+XQi97rPeczWrdiIn2Qo9UROqWdk
lX3WxIm/+KMJDqTq9GxZXtUsD9vIowsfP7dQnTzxzhHCjcAWqlApmSB8BdWVyniOBLcsEJBpmCC3
qX2oI+QDErZHieofovvZJ44JzVXJLNlUC8mkquTV52/xNosOiWblShCx4tQFkL1BaQvXxhEY+waR
Gi5smF8jnTDDdjew2SL5zNFnzKyfH43aL8hjndTo9L/moio1KsBFAHE4Rz9cnFI6eThAJ63Ov+GF
2WlN5LMmrRBBQ5MSEvZ831iGF00CJAsVQboW8cr660ZdWEzsSkfVpoyl03HFv36oaEjZOPDmlO3o
fwkWNY8Jt6JZbEHWoS+1w9YQYI/rZ2KAVbS3mDdd+nUSGF0TXy+yQ0s+YQMaDbrMofERF8gsiBlK
+Fd9VmuFBXO1Bs4NPC05gqRquezGuuvf4DRITr8bwIj1v6btMywLS4bCRCvH2teu4mwrIRbRfDO6
gXjDvczSzBDiXKpUobjO4CkXtj0N3c0gX++Ad4V6lodj/TK6jvXfVY2nhz2VaTU8S+jC96VZPXz1
E+IMLz5OwP5qHP14Y1Nl0GoB3A9a7iZuOY6PdzLOGk9Uz83/J89YtoFuKyedBIzjHelTOtCSNCPC
uvZL1w4oJIAsdqXrS0rAzcBkyrtmUIxHPY+y/Fki8vQcTpeGPvNvGMbnBymuQO8DCFL5LjsHIikD
+r+IFdBsoN2h/xpJaPuv51l9mtTxgkbI4/4Gb4OZWJsSy32PjcYEjJl6VSQ5aPqnv9SlDFQHYOak
4KM8W17gSsaQhrLJEeXU5w35QyU6istlo7qrZQyPVgMUSk4XZbQzM5BL/ZeUzxOsTPoZbViD2Nr6
2knWRnlsdZ/0OWqel8vfHY3HqfqbEW2FG6FWj8LBjfGu8th3l15vlWOD7a0DR1SxbtQ2DM7V5onc
q3yBzxiAnyreibdTs9uro1mE4+yBuuWp4Poro8riP86aOHco4iFpQNvnhiY1GIf2UZa1c8YgqX4z
eVVv68xg+5MuEKI7ASIEP42W2jqhMHO2iCfgItPhi1zbAF1qcojJa/KhKTBWvG3TBNfCNCh1Crj5
yXXjIeTkmyohFU/53mSlCPHaX9/6MIjmcIZMyubuKW5Hm42yBGDqN73WPTgiyHbaD4TGHeqrlEJd
bL/e46xauwv0/UP4Y2fPzvpQYIP/BYvjqPU4I6o89iXYRVwqZViXSVthwG8pYU49OIyx1Wq8L339
5llFEvEHwzFKzRHNwKG4/2yLXAhQNQ3gIUQm1/xqiiH0mCdte75mtpirfo6G4JWe6lL8T2OqWvZo
zOcVXCfdESzVkh8eF12jH2us7RXpAvJtcYs7cVEJAW3I3xtx4eycKnjNs5bbEUJpTyZIE8g09t+4
/V3ipg9NJ5SUuZ1GcqreVgBkdB4YCmhATJexACt0TuyQrBrGgNWbE9qBbr2KpkvtU5V74gPbE15S
cKxTjQXhsa+RbHkkAMiSn1fZTpMlo2imvbmB1/4c6uxuvE/uHCq1TTVp5jy/qR1bycHwKusiHD75
fRft5mgUQnIGn6h6H3MajzeOXsOCmMIlKsvglhki5V4yOk+Qv/YpZSvlQWgUEDaTIoSkhiIH1hbW
2jPCUCkQhx6BPU3VdIkXMaKkjcFzvj+r03hHZH3sel2/eq1Tov0tsK7ZLIULYanRd6n6QlNSS9tq
69fDfysKNFENxcBVers8U4Xg8ScJKNcD0qAl5N75dIseV02/0VOE10QWiHph+V/9Hfa2WXUTB14M
y2TlhmA76DumX8Pp6Ks0o5F41iUXs4X7QNnA/zihf21KMS0wI7kw8BFrYduTBYIT1rqS51axn8qR
80Y8sbw816aDvVankBDJ9q1UsAkkW1Sdhx+uv5HyudjDF3OBdi6hXuaRn8eeB7gE1m5XrpR+1Uue
ZYwZemVwwDwI17skUL6nb/HpeHjYhSIUMojeRzMIvKbNvOgMU5ukKsAxLW6WeX33GK59VLb3mWsV
T3jiLN4FkWpNX1kB9W3ATAOPUVgtgO3uvjkVKcBWlfSPdWzXFhwz2z8r//ea7z5iLmYhbBFvp3Ms
h4GSR6H3xiWWW2TkjLjOQ6FRJucZbi7j8h28B08XzGEN8evdgv+TaZQyqgyds7r6HSW4mmjDxEU7
ZRKoZkiXDK2GOVDFwIb9n7OqeSqWr3r7YGFlmpTo0kH6Ds6O0aP05NL187/hYpAGDSX5bChgoupa
Fwn3uaviM9sYkTFSTQYtj/gXg5OyusU2x3bIc0cgs6u6D7l3zLIPWXLi28eK6zEoEKdKm8FKf880
DEA5vCovIPvXjrplxiRaeEwpibKfKJ7W1z1CM7iL6Ih/KxXQQ72Ve0An2ATfAnHvptdHp19FgNFu
LPgiP8yI86vKECc49jytU/7F4EBdijexn6qYxqaUWduwkhvkQMQMulcsokBCk3KBsgcNyC6P88o6
A0Uk74gn1gik4LqcKFjGhfI4T6sfKBBf5P2lShhXUvs5p7S5K243Z3g/PA7qj/DdBLsm6ND/w3xg
T80qNDT//ejOeRMLbvrAZNdr1//3DRKgXvhUb3A/kO0FYpYdVkEEr9qhu9EqJzmXPc10L1XZRlW8
fLNEiC3UlgHi9sJkyxuL4Xg5NQ+9lII6gjE4PxzajMOWRYQ2+93K1Dt2LiqzdkkAFiez4mn4SRoH
qV/9AY4Imsvk7t/D0tCBovKoSWSry0+kkETqtRIWgBnRJYM/w/0BD7nkuWuf4fX6elIBsVO41r+A
IlzgZGce//OhB25EdMq+BRHBCe/323rbi2qxrkeIGObuYXbx0v3oX2PZ2YTPWGRAXqPpfOIruFuA
NSAQcsSKpB+8bgv5zzLNbFNU/eNsh6mxy/VSD5tbkbo6jv1Qm8Fk/8Knm3oxDdZb9DhHqDZtDr34
cX5CAfcRfbX8mMOoBSpITLk1cAMMrgat+5+PnW+PgsyHP1B8Rjt9/ovVObDGQqqwhzx1qDgH8ICA
ELrUV9aOJFHkIBkCFENns5/8Yp0pM9d3QZven5I6BWLVEp2JTJ+ALPk5ioenPBw1R/VF/usyUlOD
u7PMstd52tpkGMUHIg4Q6EuPF1dmUYmvpGro1b6cpm2KOAUIOMs+YA720A1cFp5qojv0XPKi4nBC
aBzbFnmXQK0EGUkzdAJg5W5TdG/uDYoq3IbAnG12dgKC6ylY8KTYNqUjJaRhLm6eABzC5PncMHEe
gopyeSyVXeT5m14dbyWpoRjqviwWTXwvQE2Ay+gDw/wCHELNDft5yHL+MXOmOgYjK140qxF9ZI9S
+RS66VrLLRcZt5Nh/oe6tMU0tGxCm8FNKJUnOTFFdy1PZ/hpdxXjFw9Ctsv+a1KmDhtlOYG8pjBg
sHBqgIKPx3yOSuRvCGAVPrO/oipTteU+JtpH5BzG3jQOjkPYGhBzaLQx/+Pf7K7nPInZeBRt27up
AqPzwgiLn2/zZzwKDQdb4dEagIDnnphM2+CHHBEGr4VRmcNZiMaxg1ZRbeWWI/JVFu35gkHjWsMo
1DPHfwVBw/pdxWKTobViT9xE2fAhU/0st/wZ33GV3Umbr6bhqK9GE4va5mQO96sKREUef4qdJqZI
qJ1RV7c25/nhzLQhRx2rWjubEG4lh2BNDDAD58Hb4KP5pv2ETxAa62qlxuFauIRzxsPgElz6qEWF
bfyjDTMJBhNN7X/5DEcEp/pFdSGZ3kYk0ymigkARS5XtuhzBdd5Hbhrf1vdfpYgKTq5tdQCIHbml
tiSwFrmRirEM+G1e4aDjjudb+IXLVYx5aBu8KgvwKWJBbftMZ4WIbIEWAqjeYpQTjXift5PevQx6
wZcoy2IZkodg3reEL/jKTUlIka8de+SuTZR89N9+YFI1gMmmOEfZnL+V8j1POuORv6cVeEH4KGjM
fyZWyif0OP2XRlZpkOopD9eOKA4ofPEm25YEv4ylHr52PqOXI7pT8LKcEF4UcLr7h2dBMYl+LfTJ
4c7sEm/FdmHUiqBbDuLa20ZGSNl/TKYOakhMMOi/75SIpQPdpXjg10hNJEKne8MGq1lLXsNIiGaN
Att11JSOXqGrxaGew/AzE7gW1OuiyF8mqAvYlN24Bi2OQtjEMZJGfwGPOPg96o0OaKT8+I/iMWW2
2vDpIx1SXSUNlNdXk89BdEflDFCxal5kUdFzrEkmdsm5B+1Hfb9wvFMajQ8gxR74sdWBWWeqfLtV
Tk1bUAHGABvkVykCTnXPH2lDtji2xtcJnPjf54s8MjWqSsm+0QxSG0jVd9rkvG/73vUmcKpOJ53V
WkOTs+qvmXzU4N4tNYl34mcrdYC9iDFOUy+XQPIv5gniCXEPtZuvY+pqb0w6xQ+vuVGJ8AnqwsAG
80HjX/oNtMiTwghivUnZEU2pT8S8ThbQNtrMcNv5KaOBT0XAq5piw1wrj0q9fpyYcmqY5cESlhkK
8BIvgivsmi2UVG4nnKC3UjYlJEnifu7oNfMhcNY7oE665ZjgkvKGHGbnkZnDBxGgapRuHWybtLVi
DXDkA45tKn24l9O9HyzQXyOLLYD0+DFVBVvzZZ/jr7WtnyWkqHKqU1kwUF5nk4MeI426Y+F4UMiq
LrkBX01jwSSGsx/voXlXPhf23DQ51l3LYuPAHiGwMcY2jRpZG4eE00FaKuXsLyNspSO5JK4DDeQF
iKMtEqGmSAj7iUoEcGocASoA/haUpsXHMi9IME1oYjJGSyJxC/6KRIzvMts7w+B6BnqB1aYUbXyK
QcExMkf/BORk+hUScZDIjVFw5gB3VrrJrDQc9AGDthgMrFzcHX7JMSh69fRuc5YsULrgErkya9oT
9w90QAwkPOKTfZhVucHJfNQ8XHSPijcaiCpQkj7+Dp3syc0T785kJFck7FW5RXIQB5Si5x4pBGaf
9cVI5IDzYykHtImJS9/sVYuBI3V292Lr2r8I0PknAjJS3Q03/QDNIFe3LQhUMPOScwkK43ohPQxR
r7CWsNoblysq0AmXedhipHHEidkiOqGUSJU30OjG3L9kEjhMtUqdsMvDVShkOkwN5cix2tN2ckeE
vVw1msyNh7xY4RRoM0ktHjspKUY3aC8AXusYwbtCb4IJKlksKUzedugvddqHs3WlJMcS7Da7vZdu
vSX0Sjw47rKiGqC3NkTF8WgAKJ7RLcnBQbMDliww/GOY8hqxF0rLDoRIpSEAU4idYRejnUI5/peq
bGfwmSXEdfj4OVf66HnAleCQczsk6RGvoDhu2F7qTYVifAmEwUxYShQv90GxMRECSFOJSc2msZMS
oDoSVHBCZRJ/qhtW1W5sLhevimHi8QM39BtcgY2MfVHSJWJTe/5Vov6sHUleyYk8eDDIrOVg1qLz
JpI8NCu8LoqyQciNjkvQsazJbNqmwCQL/XgGlW32dLVJPe8FQSuVBbWURcFVOYlCVs5Kpo5Ve540
PofsBNxRCLi/XSD1UiR4V8TqfW9HcofZbgHiuQeOvNmJAsPMQ5Io5Q7wKsDRbVjLznfJRDQi/Tbu
6hZpFAW9yNhEgnATRh5r1EMZnN1sNihAQCTWSeGzTGINbiSdMmShz7bbbvSJxqyCTQ+cCiA9yXyr
KtLCPe2+IKHM8Ofbg/rq7TXS6u7a9TLpeEu7AjMGKHpczxtX0785BSW8uqwuyuq8PP3wdxkKF+xb
EaLtKs7T7iPlDFnMB3JHIZ2874pVpFHEfYjacIwfaiIQLXVSUZLIpi/dCL8qhvoKlsF1V4Mrz3N1
22D2J4n1ez8SGJUd2C4QHssWWQ+VWCJ/5sbdWkPfIp61A+vHvKiz+U6uevzAQldQWGAHFmwsuJvX
d66+vJuE4kRghIqA1NmK3+ncdu7j9bMhvEzVuYYV7B/7QeTvK7FXybFNIeOfQaRy9QnjcGt6A0oR
Eyg01iwKLjwEjfmYV+eOSgcccjEseqf7c/gl5+wXGNvCVYttgNBx5KjLdfgumdR4DDR5/KPo8mZ4
OZ9zYkUu3cWjf8TCqlWhlU7QdbKnvKrzMMdZ0Y+C04jgHiNOTIfwzzdD1gBZyvCFMwNn9wsnzMzM
vu/T8Hce0EpiDcC2I51cwR8NJe1gbh9kpQybhAVD/T6SvvQ1vjo3wNVuCmDzvT8lmxm0Xm8caNMb
pqtc1Eah4oX8CPPLycSSn+evwfgQdedRHN50fxjH7sXMkSsSVOxSgKCYK+nj4+mmZyXfBJei6fTQ
4CrU8PEOywTWPrSrwvFsgU9lcmAALe/oGsX5CFP7pX6X5Y2U793Obsoy5A70D61USmvyGC9lTjqi
jySd7NsG7QlMbw7bHj5l2T9MHltdR+G0y1YfKQYqhZxCNWjmnYlF2Q6D0EjeEhqPyRnzjaIsei1T
Aek7hpJk8thcjM1VnxjT4v4l38LeWXB3Z6mB83G0QVQpKf/HXr9rkfRye4c5Afu292KXU0CNlRQD
kq07kdgbyArViyaa2oet7X0Q7O8XVdTlfi58Z8zjSD5Mpy3iezgQ2+b08nem1tAd8q4LGcV9yU1N
Fi9zrt2cx0XiAUc+JnkQ42gdxlzXnsXeLTsk+8gEuiDI3z2jgAATv+0AOf5IL3Q2A2v4sbx3JpsJ
xZlcRKTsdG/sw2I9f+OyoM9N65sPLazTINIfqHS3h1KzKyVsQnJtaqxgD7HUPq+Y6YysTa8Lg3Dx
Pm/3lJXSem/xNMRApWfBkM0AvRY14IOLbzUqtCOgsQypZwYnSUbrLkFM4FKyyB/6RtW9ncqqsUjm
3heo+F0Ot4zR8FAdABIBRkBVXPr7+TYGUnTZf3gA3rBvcLF0vxYPVYgQc2JFZlWr3PIvqtpJtEGh
tuE58RrFR8k6g2CRx9wpKO7OH+p1MiMnbKAzw9S+EwmTZrvs8HGRBxMI3SsUNInTPj0tQ0gdm9h4
FSPkA5V4jNhe+ztvBRZvSywc/nfKvnMm/x2FOoLo23N3o4gdiLVkFLV12qexQgjeS6XE8+ycROBV
j/ARoNOFwTm33dXgm/yRnmR657qQqAq/Fs/ckqPwnwLrniKfGFXiZC+M13m4o3IkY2be+LlQBI6r
GRQHCSRSDjraMXS9iFzNlUESwnpnPSqfzuUNNZoFxGTde6kzglWvdM51u0rMkv7rilOovH/lzHDs
3MXZaAQrIMjkVDpdHg5Fr3TtWbl5nGBB6U9tCX7AYh7t9imLlhqG2ngj0Jw/Gq63clIEyfVdiOYC
fk5ItNRW0G4QAGI7DDxW885GHeNdiFxkFl63Pv22JVoQQMrbxBqKx3y8h+R+a3SMUCcCwfmk4ToP
JLIQKFb6kQtfEBH6VnSZUfrmiq/GVOm6YRMoOU+yR2NHrWZo6aeZ6MlwTA9eNpGj0ZsR8CQWT2vx
fYI4v9Pqh+ERuRRqoJqYNret1vLQPzRSUQtsZA9Z+YcKm36lEc7qC13ZpSvoZ7ZCg10tOHKE5bbD
2P8S30meu362G9jvvasT+URbzQTwZR3aH7oBXMfALugJNvM2w+qJ08VsfDGFFsN8XqYOGFjmUt6V
FqaQdhNSDl82h5/D+jeG+KEyEBbttfWMIFy/umBDORKBiLfBhrdGRoXU4XA1jTLgZTeWVl6vk2KC
Xp/+uEyL5ukbuPfy//oXhNZ2rH1JjlyB4lamYXFoqAjQ+qtH9p5MuZzTsyRqEBqlv6OOzaUdNJTo
0mCw1sfZbsilMHmpXt6L5Qai9kzQo7RSyU1T3CYkkGRe9AU8FggZHruPA0O9TkOmuQ0jOfd+A/Up
k0T0Zkdsno6PSZKnsMPdKn/nEL0c6e9FT5uoAXPnaqIkh4jSMhhcqWiR++pw+2bHTSI/nZqDQGkW
FzsKEDJHj1dwodDWlQEioD1HkoFgSJfnif5iJgqUqI2z4uOn4VkerpiGDuC3yqmu4mTV28FXaVV8
pBugtVk6Y1cP+KMeiZJXlauQOMjT4sJiIlm/IBNTP5nYWMacS1aFKoYEkg6rbPi+bvWBM0We4ttY
ynFmGs5oyKb1klzIvJ+lqSwx+x9fhYHsFH/iRIdN0aYrRtH6n6UKJEHcBz+M6F6zSakhgDKR5RuT
MbCci2kqRy5x7sdmn3S6BlYlOR+qv7NnKKAjmrmOkzxtKHofQknS/HxQ4S143noaAobCiZCewOt1
gQ0FfpP9H2nxz9ZeCqSzpEJTRzesDd73YqDMJ9+82ei4Um0hqziwX+efsrzGWJc6UZE4kq5eAJfz
FSHtixxkB1hjvByzVb3z8IeFHpnfFU6/ekoJ4OCOftwZuj0MtRzVW4h3uP0YFxYwQnl0xdV13uOE
ihgwyBasD6KFOQNA4YM2TJTJ1CfJ0yilJh/mo03NvS1bS14NCfLz1tOo0QOExVGsHLOfvJEZ2FNf
6iZSH/7Ex2FcuqqQzRTFhQm36XVitShB/B99+PJ9ZTryk1o3RhREWsuDBTzNk8KU7VL3tjHh9Cyg
HMVSyKOIlhjp7tJEXPzJVTgOKf0e/WNR+0CkvV2ijUALLNmRvXCqVqRcgc5GrkiHxOQLNMG+dK0r
gB1eNBqyz0it++uLw8TqogfPXyzuODATXqj72BtJFpyHW30cwKEkPROS4qP/GQvZZYqkLRzQMsw7
qa6oHX3xlGYutSro5FlZu7jwYJ/uExB+30q6//O9cuMDANEHwLLQKFXIWp5ZjagaKlrX4LmNBy4b
of8/Qc3h6DjPFgzemgmSnY3yQVp9TOqQsOTY6HMqxurgQ/F6TSqbZuc=
`protect end_protected
