`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ww1cFCaKpEaygJUT+P6Z2OD0uzJ4IJG8iyHDm5UNlVWbTWS9KXjZ9jEg11wJmlv8lA2AVebHxIas
7nZJsy/GjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gy0/aj7fr+HoqiF2MKC2DdMRffpsNgkz3LCA0LoXsy3oP+ExvEwYs55sO8KAxVdJaUPMOFr+w6Gi
VDRBmTTzMTTD1KvHQEhDppUtYnGyL/2qAWb6xHvmSHDtiAjlHews7qZ26fM0sYgNx48H6LSqgFd4
hai7P1C8/gEiLdaec30=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hi2M/LxF9qgAZzAUuc501Ws9I83yzxDz1ea90Q5QjM7jLsFrH4fLD2d0WWY2wDTdG0Ih+QNnE4S7
Oq9DybBH0zvBRUhAQoExlvdlIfU3Jr1YKpM3lLPQTLIhhCp1eQgIZljQtMN1p0u0HDYYsZO5DBeb
LZHGhmPHPWGqNQ/iLmQ+PQu0B5Cb+1VKyvK7Ipxjf6wKC/NZlztCmWzwV4WC+jY2wHB2IofyzZfo
xRBIRCIpTb+tTiKgZ9oAjPNYVjgXC51YW/c8ZhnzF0gIdh/tD6GDSX/DdrrBN7Oz/gtduYw5jR0b
WsJx7lVGCa/mgRPb2+p2mjuutW8gGGnh6+Yo4A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X16goI57idQ5Yk2jq4rj0BhsplRtdzoYr8oOU2lBTTonp1Nx4fK7AS7KgGuzY4UqvPTHmPTfD5ww
0YcXmh8hr2Hk6aIz+aWFV8C8XcReGDrBhi5Np0Vi5hozuTfEPpWuDV7kTmarku7FYKZbPt+lsAsd
f8+cIo7ySKaxPnzoHbw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RA9GWDJZOdw/NASVbYOgehelK35X4QCDpOGKLkbLHbvCU34C5eqCOlazH25KMTrAHxM2lx7+fAsw
HHb2ZWqK4pB4ww23gPcOsgxVCyXs7Dx/H6E84snPbj5EBFAp1p9GZJoguz0skOVQzCSeso4vwekP
kvLqf3Ypkz4/BbGmeIV5O3MvxWppwuIHCb+NDzDYU2x9uQ7mLUtu7pYCzPfN1FeLiv9ttZaXRuYJ
ADExpcAMpFzH3bwg6Tm6wL+J1DzA4jLGZxI9jxK+L6xNTv2NtONryX7sLla9heWPJCSHR4TT8ow3
t3QklA4V7oRFEhlMh0Nv7QVOAHjukKSZ99LumA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24704)
`protect data_block
2JEuFaTgqghMsv5lmjCzRKFTRu9v2Bd7cfnnEymmK1IpMPqqHVgKVztK8UcvkN/cLu6meLkuW+GH
jEF+IasLsTsQoEbARf7iGoWy/qxr/Wx8iI4qK11niwKvKRzj3E/VIfcoFWMI7lDjskoNrB5ON374
xdQdL472o5haNrGgEzQCs124gMoZrq6ZZftrvXJyyhHqGqmNNfQbG065CYcPsuRjXxzPltG3oMhc
7n7pQE9F5O4ObyVFgYrFINih1IyuB6ga3CPJSEZRwp7Gz0bxN4RD0DBaR3vYvY1rH6jZ2As9bin/
g6/KlClzLL3bvhOh19qskAMl+VQgJT42Uz500WKi6dJbwwYRcFurnAISAE5qkqUovb/aUGPaj6N4
OUCzRVo6V4xshDidQyMof1ul3vh3s4PFZ537nNLttAZ3Sc5aw04pfAxS3srG7aHPtyrK8Erenobe
78c/rwP/AYGAk+ofBrr13w5BgesNk6uwzHFdAF5hBl01QzI9ySiVZhndOfp3lQ+S6HfUA9lHctl0
LHmuGv54CLkaiUkc3x2dk0i5P0ErEMyXsVwojqB0G9fyRNeiGY7jqKVknf/CqSXwOsn1TuaOo7EY
kyjIysN4191JuTrrtYdm56cp53KyyoX1osWn31kceQNZsrWNk2DoxxS3e0eV6eIQTg9rNZhke0Rx
wB5WuY3eeQFzt989EGlpMZytqyBTC4Msv8JlF5okbdGlB69tipJ3AKIduwzVhe4vla+kag/1xQIJ
a22oce4iRMCG7J/uKMPdioqzoz2XLGhWc+hxPWyJDHC91XJFTI9auxqVEbwIVq40pXmCuagZUYhg
SlRb56tDFbD8yZ2WCArSShoiKOPQbC9F4R7WLBVuOeNmyYu7Lfbfjp3yznTUvj8+hhDGh6/crIjs
xAHgYtLKoYLTkqMn7tY1PoKcI15ZvzFZGAY+xPUtUfTQULEXZcFNa59jcoEzGugJHHTZ3OD4Tjlt
7ZaXcUaYXI+u8nMOp1MiMQ741JucIESHjlv5nebCKpmGwI8+7EItAZx7JcypL2AcodW2uywezgOE
KVvyubcJ8Dab+FB6GxpxQt9jGSLp+qZyAvncHwFHZ2+18NPHeFj9aM+w8Ts30jcLKe4960owv38e
A7BbBnLHssk+xAtAPyo1r1rEtSZgjNyIBnjh6aRGJoxbr6KPeLnRya7OjcA1caL4gyuW6lVF3WR8
sE5GxXeIOD1dTxvqCuWX3lsZJCpt5V6ieyrUKvpx2I6u5JM4/EyfHvAyRJFMXtD7IMAuwT2P5pRQ
mgovuHLT05qMmaAMDyd/AlVLGFpMNezgjQQJYMp02DRL14qIPOo+Zcaf7g4N7g/mmwa/WE2MBGpA
3iBijJy/pyEQuIBTvAxv1MB6eRHfzeDttINz+b1Wt+0h3gS04wpONGbM63MpQUep2+u8ltNZ62vJ
mePncq7YYgUyZ3Vnz7Pnc/c4z4EnTEQU51XJv/O97WMsh2Nippaxog1xFLDp0QeTC4QV4uBdPRsC
HvfsxEB1dusfrGoVoovtX+rLMhy2ORwum410Uzv/VLxbFkGbSvLv0KJFk32Z1B/nPsQgT7ERLeF/
gVExdW8HvwUswPow5I3dphmnJk6kMLSNxNmbSbsdTz6kfeGtuxAWzLZb5utPU2unyrJUH35Q5EWj
bB7QqikzBQuiQooPHuPis2RGwa5PGTsg1Uhu6OfqttqJlfK16gURLMXOBTHmEROcUOjafUtkAj6H
jCOO3zhL05APeINWbb/xc0+EMXLDz3PDkA/GIyPFr/4fv4FxT9+WDar+OjZULm0IfM+xghUZqPtL
3SrbahTw9Ik7CBRsAeyqcXMk4pkg9DQeC7XI7RAb0q5ua0s5/9oCDt/rNgVY6AUwyNgiOjGUuWBI
YfVXwAeaSswVxP6cdwdYrvpUg5qrqkQOLRN5xQKLBqQOhVNtZQqlHS+OtCxb5dAPQgDp1egZT0Bk
fIE/yy7F4iI15KnO8FkRlY/CwLTT9nOOZpzlW4whEjTWD3rEKPgVR/MteMm0+LVJuXFyu2PpsOdT
90AwXphuYj3QMR0ky6rnORy4xWbbT7jH5yr6CmvjWbgT/6r/13a+rhME4aXDfNlnr5vIb2QRvAm8
TbnRQ34NeyxC3QWDTBBmSVYNRZW7xzAJ7EMdz3vs8DYtNCubBbDa/VTDFoa9bVxHrPk+HesNvXuV
u+yfnrqo1cUR1yNweYxYOmqomLPXC7VgjWDyl9hAl4K7ipMQ2t2MAaoA2Aewex4E6Shx9NLamB+d
wmauUMz3UBjQb2hZvGqksbnseo6cY5Ul8T81wL/fviUR1KG/bFFfDJSxRMafZwAQHs6rjDyPX9ft
9m2Ew6Z9DgDu2pCi7683L0ZwOX0u2smltg5Tsyh5aetqugQG8/dLHYEx8uqqtyVnLyLpLQErG2fp
XQoIcC/hLysPYKwntqZ/3s/GG12pbKeom4gXn/x8wWuWEFakWTrvGCQaNQem8BFqklMm1V4OIuu5
WO5aeVPmaHanl36OxxtqP4jAMMEQXoP2JOaKrMJrEsWwNC6g1TW0Eo6FHHMwfctCQMJkp81wThH2
dN5d87GZUbJv+kC6Q0e5fX2wGCcyeQ9A9MrlUegruRLgVA+whbBpQUl4b7VfqS5oGuKbn5QFRNQG
h3JjbQHLvzE2MeKam+BJv3oV6CRZO18uwY5V/kUQIQMbQV332cqRQJFuNsh2VkBCdNPrT0lq9/Tj
tz+3iwVK9HL5J6JD+cNCCSL8ejiYL+4mZ3mYVjsIqPZX7n/O0FLOwWdMNGM8ab+Suk1jJo74FuZv
Wk4eafwCDkMmiwYZfNGpIzHXzvBDccRtMqjNJhRSBTKf1wXZbIzfNowqqDQWa7+givjsPYTM98CU
1h8CO8HTdyiTmr05G97Epe/ANFOUFTTIlWiWLi9wzvJh1hA54Jz15lDYQURUOW0qLGaTsaDBCY2a
8YQzvpGFOrf+hN52EOZ0DGaNAO8HcFBMPjqRoolONDEAxk8bSh1biYLHH1XcVSIKzvbD5lnmfkLO
r6o2xN6Goepr02Eh15G/4s3/0STBuxTONnyVKz8y+sfXfovRfi8gnNNulwWw/P3W7tvv1N1r3tOW
wpIQ3cmR6J5Gz3mMk7fXpl0WwI6KzQSo3JrVHUlt1ZKgx3fEj7Yr6hTSim4hZ5d7Dy6khNPRxIa1
7t1unMRJT7SF5l6vsCbH+bNhm4ScCZcZC64CwNEVMOoRw02YWBfD5Fxw5yrRXiVrDc5gBMkHo0aZ
UPCVwYfZ3BfT/8M3YGF4U/CSoT2xmH17P3ZHH0klWonv4uM4RqfXPErM5Yz8urtFaX9i6/snkbnc
Fg2Fawe9p82omUy0NM7hlox6qdbx8pKb7mZ3k/NItqT0j6jSxiA00nI51WcYZvUadWjpr++CbcYq
Yr9FBf+6ON+MfPzoBSc+uauMUk1UcfJk8uB+kUo0EIul/CTHN/WrZMGC2eTAp4TGvAB/0jaTjjEJ
eC43OnNpxrygFzURVnT9nnqlKXDt/DOWM4c8fZU6PRL9vql2tVRntz0vB/HsQKYcOWqvIXSFRRKi
uljIKG8uSZp0NN5+hHCg0mfwD7lx4J+cdrUkQe54PggmJhtrXDDacC3FyNmTZuYNuSu9MaAiolze
XB5mYuReI28v+iLgvWuxBYu6o/2q4e1S5rOc0yHD5uyAOFofMvvpyR3ewPzAO/2/D2kqRsHTiS+B
JN76fP4B4b8giAVMlzWVXiyQTwiLIBMrR/SlxXNIY7ty60BZzA+PZ1RhONaPbCMECZVnMIqwh8xJ
g1H1HxbV8gbZm71GBki3sggbo5dUn7NL7H+7MnXRLatzlpxyGBpaufadvjsyTX1e2MTYHJmrFpHH
ErMflmLvzfRzLpjquljcvxw/wOV6SLDWG6jucKtFfSzkHgUJnU/3gtawZYoTLXY4J00zlJ/bQNFT
iNG4sXbls3WBayyHkBB0NUZyBxeJRtJdnLUdMuSeQnk9QQOS953xV72ZbDp/UDr0VTkX16OY8R3o
d3PTFCsYbRwTqQoPDJdV9Ss48ZsHJ+bDu6mwKnsSiHGf5p2AEEYYSA1AqryDyxXmSpikFPqUOjIS
jKkGGKxPjXvCVFaAxjYBDaiIYO7aZcz/djyP8ZvJKQyJXEqcVTCN4x2ImKtouoKsd+yeDrppndWa
2ZVToRwRehbze/HoUgbsyN1p2wQMTj6rJecGkEUht0QbWFs10a9nFYPyb4T7VpvuONrUyyr+AS0R
Oz/3NgFK5g5xTh6xy3uaDw12uzmNTj7IifRXu2bRczXGAaD5LaaSGl8mxBFVFgYtRhWSMOGuY9k7
f0tyoZXjkhRsY77qEpM16nMjKdTkL7sHRz9r1STr1jMgG7HMPjdu/saF2tOBO4I3m9+OfhG4UChA
Y9JqTwna43i5QITxsU0SIlN7deHk6Q9YzP85PmJc/uL0rLebei8bhgB9j9XV1s5tMBdvvGcNc3Du
tOrSu0gkeKhHZQuenOOyFMT2vf54BOOQ2WOxQBq1ZOFBhP5w2nFMNDUwKDsCAwt/a13m+Su4pzG3
fN9HLvyqfTY8zzzLNgQgpwZlLaDlpf3bYvGRWGMDOQbJLb+7J7A8dIwqzt3HVZ/av1Ouixtq5DG4
38YzbNj5rIOKRj6HDexxSmhSvW6mA+qwTdEOmEbGTNeBlWoY8raQ7GQ9oX0/XDTa5JrhQO3ZNlqZ
aWSjtN5ItSjOLc4pSvJ4OWN9Qa/uzv2XAja96ltvvsA23GYd0DO+L0ZMJK8Vgbkw1no20AIvvtJm
/Ob0MpygHEKd/ObD7SHmX79fDCwmeQ/nX/hA3khi7E6hLKEIPMbKMGgeRPKBS4Bb+qByskBxUUEp
1QbWdcd/byhrjxPFcL77qOx1C9AVDdq+TS54zCvIRCEGxSYeZiIAq0GfJpWp44j2WkBCG4+gkrQa
hhGVv8rH63NIFHIqPNE1MrdMKmo2ZYCGec036FH974Ar38M1lYld8DmNXreZH7CeEok9a/8O2LWC
EpM4MTnQ1TupkBb3LAKpHzWhhpO11wITzrQGcczwK34DlulkfbDFm3+ZoHXOPdCPOgPXQkGJymM9
pki8XYxWYQfAZAJI58IYLK9wHgsIialPJLKregYeC9QEFzPD/gXnphd45wdovH/AIwuPArJ4SUIt
SlRwqJDj49rKyQyV0DPGnPaUcVxP95o+j+5Q2GjKnSKkjc3zCHR4pB7I3GQkXcadgbtLFNN0x264
D00FpAZWcN6G6Ge1/nCLA8y2zTQ+nxugS6gHFYLhfDu8Ei+YISSr352QVSM+kCcJBAI616mUUKeP
W9nhHLXGjacxwsKwfMY+EFW+f59sKHt5XgeIonIdh5KifFPDXEVWOIE39EWqCEya82RrXQstlla/
Pvk4BqeMvbbnpSDJTHsI8AKA77gS6nagdrvPb7biVfilIYsQjgVm0RZ58IXHUBocuD0VJH33bmwq
mcKB/VAtyP40nQpGxOLmz2ozFIsGwpoKf1P8HCXfCkLKhsGs39e+x76T3aIBqzjphKUzpe+2MKZV
iPgKMTnDL4+xHJW0lin0uB+tLxkVk7+Shsm5Z6xpsNFuBjODDUP9YtIYHAbyPGwE6nLOSBHC/Upo
PNqh8nvowdHOdAwl236d90BZTuoPqxuJUVQcauSKgh12+m1orlnAdYzia5FL5QP6Tp254SaA+YRb
mGcmPkuzceh78M/CoMkuy+FGZ5XRe93LWNGmNmu13U0imztEVUP5rRwN3pIztbhV3bLQafE/D0ZC
TOpWkhKh1JyErl1ZI7Rdy5SawmzI/hnxjlZfi9MqaKFcBmkaGioR8fEmSP5xHFabEdDzX0E1JO1Q
yeK9mGmxxA6tJeL/og76Km5weEXKzZbSdRLjCCTxBkhiEM+CiZH/uwVrgn+kgEUk0rsjeOMen2OG
MMkA/++P3OhDz1Z9n0QtC3O++2IRvks07ESEDL5Fkx0mZuHBoBWfAwN5fscg1vg5xZVl1HBAbezc
dKMPBijl+HtDED8Zb+MZ/m4u2lyN+FXM0YRff/IiRfG5gKqsqWo2D3ixoTl8D2ez0Dmp5wgAgeLo
NYr6eTh6jQTgH8g9OvwvC1cM9dWMxOyxjaSokt2+uEgBOpMZm1B4x0hzVVJBF16Mrxa/x0jwF5yc
UjMjnsnZHYTkf5n3VovP3brzYTPbKM596ijW80Q5kXH8Aj5vgXTUntNAlbFKsmSVcBaUEK6UVgUZ
iwq23Uk9pcStnP6MymAC9CjpiNxd5VfJ8XVsxeRlBgWEz+aeeumoCs32nJxf+lwpw2zU14EsIqW5
BaRl+IE3D1Pevo+4HjT3fLOIdhVyvEjdW0lWZKKAqlvBvU1FTnEWD82wzwB9lYdg+tbPDCDI6afK
wYU2PFuwL+AvX617/+wxf4sTGLyJsMv/D1dVubyOMYjfJL34sYhusd6jo06cW+XWIqdlqyj9zRCs
XBMgBdKKSrz0pMjPsEX/Irn1YsagWkh98nmVtBiMxvI8uWQSLiwxrMJsEzj+MJl+j7YsrJWJRkrh
0IlJuQj0YFURSKuEzf2O4mOEbN89fxZlhH4WgGWLhOL23l9MlAUDTavgXyCtr1e1HJj/PNh5IqHG
HBJLjesUCMARBm24k9AdPu+eM/9ed9jKpdZTaxtYYel10bpEMNkW43d4O4QeImtenwAxrSBDs/wJ
PWd3rnVdijfKUTNth0TXw9c3pp5paODo5hfaeMkFn6ijwehDLy/zwkKVpc9rJMMCULIKBR0CUAa7
NIbVS7Gj1yuZZHhYrGOVKnCRMw3DrPUkdCQyrHGvTqMXLQ4faC9DpQAAFRPLQ6umTe2+xf698gTy
K2uMqlm/SSLDUnHZfZ0EC3sskcnHw+wIxAygkj6Q2vftu+FB+DZIV/2nRrV17VPFeEQZf/kPkXia
++820O4lGqZGGJEyfMHco5TVXpu2Uq2UmdP8xVZZSVVaa8lF483biuEaWtjKeM0vm4Ci7c3ItTLp
HY8IaAlRNfkdKhEFUqNDZovpNyc+Jzw4lyeXKkgh9UlRzPzzRSR4USVjllOJL7QNnhdGHmACOR3q
vr3MKbO95d1yQGErP3VY857XcjtlM+QLJdqRGPyHaLvyibgKd/GmglcXfF2xRHj/v7BQ7AJUahOJ
0PNMcawwe3DWnGA6F4ABQtWf2pQ14BuWLPu/ZPrZrwa5Bdxmsfzgi757galesakOlIp8K7nlWppv
PBpcTKr6Suz5DgvBeX7+2XrL4Z19s1XuH03xP1cYzqu2Dt2LXzTy3t6J6lrP9IK/kb1JVo3fayf9
BUCrh1gLB7klpxN2PBRTh0F1w9Mgm+j98kdEK1OLQ7wZ1+CFumavt2wlUEwCMAcaOM3/SjIOGxCJ
5B7MeSqgT0b2Qmq9UPnk8I7acWa9qjB//XI913SkJqUW3wRiIhLp2RW51WntfJS9dasc2buVbUIx
ZvdmpPPmG2imHa40iuxHrBHw95a7gkwkYym1kf9Mh4IcjUQ14xdON/yZ46hfD0lXBt3Me0CW/47U
yflXxe4/zU1S0PT952Tx2lwYS9RVxI715UL356CZa+NUOB2hh2jLJdAFoJfaeP7GHsYJAPDSeW+D
TcjOwQVhYO3baGxCH2RG3P/682TmUJfC1TX1TW1Hh0cpZIHmFVlWjvlVsvokW8t5kUaP0f6ByMCt
OuwUmutp59bqaJXlpAKqQvvpgwE99UANmHW0QMFBtkzzXdljbrkW9mF9shXIERDmYxP6lFRBUUSD
JhDGLUsdxpp8X76QLYuYGWe3ev6W70eBE/M09QEsFBEQeziaiAFPPnPa5iJoPmiXzIOcmLnEHxf7
8wDUf6KaL6wFto8OknLFREd8zMww+/ePIZlEPFMwpqvxEjZKwwV9JoVSBHY9LSbgSRWAXiElmdxN
BRU+3oRV20Rjqt8Vm+wpk6K6OWXQUuKzvHyAythOU+DIs88RorusZ/YOX2hd9zy1fdtMl6DFkgku
AWtkLbJxGIJkhTRhppboxSHPLygv/ngJo5T/tvCPuhEr3k0XIQ/tQ+E0h9bA1uMVJjw2lMs7UDAN
Qk0xcgl5rhEzqquFA3af/w0oaojolOrwBat1N3RsKOlPffxYw6Nb29mV0kI1B1WrrfZegJIKn+Zt
MX5AR9Sbo5LDv5lYLUPZwQvPN3bltK/aylHi/O66SFb4DKnGWxMQRqXZwiJQcCdloxUAu2ufDRGi
E1N285q+qwR7srXqGP9kxTVkIuQTJShY7rfLxjCBuVvp/KORreKjHbkyFHCKDTxMJB6H9Ay5HxWj
UYaypYfZUOb/2zw39TEnXXtwBhUtgu79OTRIXcPbNuqQ5FDq7tmzSrpIc9AAoo5rqyIRXjOk+lb/
ZZ5cSIApqKn+CcrxBC/twhiYYcAxMNkW2uLhVhkOqKghJj1QQfRrEhRFco5avPoxVB3TVUDZGYMC
LS4wpwcXCF0E1k5PSI6RQAwZLPnH8sCmwkl1Cli1lFXp2VkZN/wKJVwrbXpANbYzMnj7rSOMv77V
uLadRsg+JCRehSkYf0wF3CU6ldKPjDVImzZMdGoy2m9iX3sSWKsBQxHHrUf7C1FrArrcxtIh6Isx
vlO/89EEuebW+BJcHhA2cp2QqA42PzKWfnPQIaAXOg3VpTGR2AM98cd1HaLVEl1FhkJLv/lpFVD1
uqKtbVy/rfajxMwpAJvqkirVAbJfIZ5OO8ru/a/Cz9EM2n25fej28JugctMntGDzIczkVAUphAgE
mIHat7SGjhzJOtthPAWfz9txDh5XZ9nt2nw2B1VEhgpp8gV6G9HH2UfHAxaP6YZao0yWSmspsZgf
vQkSmHr1nkTy3P/eAMbYJfOfC0oobi52QjkhuLWfArcpdqVJdvLQLGYWUL/4u7fgSVG4Ilu26bRW
SdMbQVXFMr3iCSOm49duuL7jrXfjIeqrYeiU0lV9mKnD9U8ovC1cadmFnMx4NIksmlFGoVgtayHw
c6WqbMqDqVsjXX8mUHwDyvvrSBhZp5sFw91qGp2mkIp6apS4mYCALZdXxotbNzXpDWDkhQMzlTXX
lZEPwuZJ3GCftdYVwZSMcKgb8HC8yWMEzSTD7+8Pq8C9bQ7EgGpap449TW1nt3UnCTUFfe/6OKHs
DAzR6gOnOW3z6IG+en/qhdk9SbQFCLG469B/7pTkDZJYpt9ALeNaFXjZOEIxhqCAR2m5Gts/cmVJ
wHEZ+CyDgnCSNr5dXL72ivaW8T+ANDDwbekScW8y3A64nE2QrhcspEC/kivvGYmAHDXv/AS/rnGt
mciZdyU0pshIeerlMVhjJZmk9RzautHtfZp8J9CGxXgpaqltM6t5eDs8jAQY1bjel4QmiTPjwtsC
ASyfWS8JkjyoCLgVpC2p1NW8ef+bQ98InI3TT9iT3DqMV/oZp9jMhutPlBxAQG+EPppEx5ETZ3Po
g4a77WK7rwK1keU9qs3oqpX5DRs86dJoUDE+WQcQfVwYRX1zIWtss1kMRM/YPpj06Yooum6ZrEsM
Wzzgyne23IJllw3B9LmcKG//8hjlLELscpbUs7bPCxThhHByw9pQvdv45n2teRjDa8Djraga0sQf
rfr9vecbpqUir5HInFytHQkb+yAuVTC8CtQtgLUTk+KGJQNN2+Xquatwwalcl//c7oglxZFXndVj
2kdfQMwp+PKOsDmor7TGxnLsiHnnekVEbnpX3/ezzLM2sB+H98/qOCey7eDwvzKePdQL/5TpWa0Z
YtHRxnCEuMOMjmwV7QxRyk9luAypM5ZG2GkaEiNhS/nxyKop0suANbuGz9X0jUemjEs6O/qFqPfr
icFKxZhxlYfBKLnXEa/5iINW8BByc8v7RVwL8G8AplyKvAca58a1jYEfS3EzGIuX6tqpNoj07nOf
jcfHiC/j0rlKpeXNa0lRAOuij41xYhiA6Kq+vfb6Cc7cd5BK/tOtrQ5Ti3h0su3ig+SlGPAQhl0l
wgDJCqZIqqi00fof6nLtGAQNEZ34qfH2iD1vb38825FSErmesR6D46qrTiCiEjWmlaPAFYFeG808
PA9wUghNtTLazTN/LfH5bkRwSwGTSDi8fQjl4QzZDZefsCNMszz0fXrf3verFvBowGt0sB0K3b6d
qqpmNRW4tjoh+3ghUAfqchrTTPwsAeEKRy57g1IQugPczilcNsI3rGUJZP2R454ZoIFQm6pMoq4x
EFzLoLScXUtIRwAMM36fJ2GdtFebsBU9vxYyx7DQsPfFWiN9EzEbaiQMgAUtvGe7enrlHjqVEqlU
qUD7kzC2yC6T+G6DnBjTio+qQL6+tCDr9oeLEymXYHlfoRQmvmnzr8cc90BpG2ip7Flb3FIh4QNK
1j/9B+Bkygs9IKUJtHZxKZGypyIzZhIIuIWUBjXCluqwLyK/n0ViIyT8GvSW67plBvXugYD4bB7W
upOexW11VKYPJ3e4Jfy9viIkuZO1w5EejosqwCvhnkfpeILYT2tbkCdelvqYQ8CduwMR7owp7c08
BkIGjpDIIA1zPfvoX+Rso8vzzphPrq6KA4URE8nsA8aQsTUYlB+B7iMUQ4XQnrQZSPX54Q1ovLv2
nseBHp6/AzMF4D2uhzn0AErBCUbHhKw9Hy3umCA9uWhArt8wH/R4GAaklzoLVLkkfgw8HwaywQHw
Uur037sC4+m56qxMnc90Y+ZBM8ZGjvAJTNMYqLJii1A30rDh0+aJiOh9xYWB5cUtuiNgrS8EbXxJ
hD+HIiIVxI0ydPwpdumE3+NQ1wofTDH7M+oiRyY6U/tQUd96gHDCYPbW6VS6WIBLaFCaKbt9EaWv
jvAWSzKV3PuiS8H1TJANdigJiHhsZV83QrEAyUqMRus+adm/AMBil4A0XEavxETXZynoY8eWRm05
/JjdbwW+V9suJ0D0x9AJus74iqPXMCEUFPxSpdI2BaFQBjzcPmlo/932M5wTyYgXw74Ogyuuwi2h
hFmxvT3qDnpDQnfEaGN9BqgB0ue8DNiz6LtnGdnBXszlT4nYuKq+OX2a7vg0MCUb+oKnpNnOHFsn
/VC7gKX3U3+QYwYKp3TD5JaFO2NEt8hqB0LNwuPbu2AZJ/eyyVuiTlzHsV/aGRsnbXl3KbRk7ljn
6cr5qXL/NdJZ+pQEZ0WSmHfB5hkRLR0kLqHGQDgcbdNpx/Ox3G26/RhZJYLHBWXieFvlReAKIXAz
UjnGTefdZWqopGf4pQJvYCA40LQpbDGijk62SJbRJca2kmE9X5ryJjbNFI+72lTr58uOLNh7ug2J
/5ol8KErnGyiKhSq4FnKTIREkBPoDxiAUGOklEfnTARMglEBZ6D5G+DX1Tp4ljxsTFI1CrlL6K4I
9nPnDxzBKcYpZPTkayoX+jbJHJymy0c9gu8++90gFKS+YFXEq5Ht3YmFxUt7SVMcJuNQobRSVD+8
cn4iC/6dvrn3yCgpXFaecKUNmx6em41P1pybVXTPstNWEKoTWQyPPGejoM+42OopDqG9zRMZlvyK
rmzWiHLmHswOyAv/kkfFKqmDFtCcuIFyUpit1Ucnw9GAq0v7lNTWAGl6+VVPHApA9HJwGSi1Ddns
SO60zqweXQM6H3zveMl1TuUoGGKtUGLhDL20oEmmWGuQvDKOSFeMihKJiM5oCYgBSQrHDI/m/d7G
u+uLLZ8BQwqFSkg5pw6ieDfnZw6o6pvNap5NEOjh34myETBDJHz5nJY1Q0rksi6K2UFkQZRBjTTS
xr2MIM9xgSvS9Ske1pLJbA8vwnWBq2/8CpIigHjzeh3uWVr3Ue3yzW14Pfq2+x8/0sjNXyPVUTM9
+SiGj7fGpMc57mBURBslJVAb+BcRsJNI0y1KJxBRkEGXmIXZgwKPvEThNNOnMghQj63c6DwFUY0i
dzn76BwPsj4Ssbhd5Jv+wsYhnf4FdFrpr2gMADNos3lgoyk+jPNaDVakbKgE+SG8XHKODKCJBGHt
7PlUOkYVJEYmL5Z/o87AEgZGv3l9FnMdOvTHoUVlNzpKAnS4g3UdbrN2zDywTU/8K6k5zpzIFfln
SFT0P0U0ssZFa1k8nTowBBuyrSCDtETXmJ6HoWe9896+N0k9rPsr9O01sCqzYAgHqceRx1TD5aLL
/B/puGxPHgAguDJG7YNHDy0x7G1geg/uAcEXYpUuz2BRSO2Nxq7xLvW3mieJoN+2wNMYal5yBOpT
EngcsgR5NTxC3a6/ER/RMK1B1wDvlkhWqJ1P+Kjl9l+441PIEgEvkuG47WGWfXy3EaufWO595jU6
EqeX2ekjuyNKGOGrz7BMWUwcL/3Jv5y8G5yWrKZNG9/j57NDxV/f7BBH8vKDape6IPijDzGWC8Ve
rhLvgx7nhed4EJd5I0NOo06c5auJvM9dE56l6wV9UyoqO/ghO71tt2yXgT3C1gABTxgfjRUmB7Zg
089bzzipM/BlIbpyMb798vUck96ouCe0AsiIhjZ0rIHo3UeShQ8JwIw3ULhdb1+/XJo4O33VVSj9
DEML+Jl9OMQB8nVAL971eplsoO1YGMXL1MW2zAH+bwZ+5lfKM2HPEJTYrd0ngipMh41ts2k0f3Zz
7KJ5JNzvrtJ+QK8PsphoftdKPv0VePU4YI+e5AGJ7yGGRl5JgEWK3lET2rRUazODx6ugj7iluK6Z
BgEGXiCB/QtLWd/niQXvv3AZDmadD7d6HHAx/G8AoyqzwcZZUNIQQ/UxYm04qF6mMKPQW/X7jLzG
LGf8QuOmOhZGEtvjq0JuWuI80/Q0EPJa/HSCb1rARtR3wzusAHiVIVxvQwRhpq2OJVy/rKGPDL60
Y2AViwT6/BPMgWd7pPuTBUsDaA9K4r2EC1QO1hEfMASkb4XxGo39FUv+ivt6dlOvAGXLEAEaBuUp
v0tV4PgVDLmqTConoGewmB34cI3fffwSbBCVC7Q8ixa/r/pS/AUVex/B0w/9aB8hNPxAlGoEKa4Z
u0r+xQmEFMW0mcveJR+ud+B/C9D9BWmDQO+I6tngbQhS5r1zTtejNQta0Ozh/mxG/FhSWdxqqbsX
YsCDrfBTL4B4+QaIOvY7m6hTRDyUmX3mZH7s/KE20Cjkn2HOz5EIY2A+1IpJP8QLvKGjf95JvTZa
kMTHx4KIsCnaXKgJcH+beoIVaNzbGPNXwwczuV0Nvb16uXaVxEgSEkPXu5NSJ5pnGnGCLj7IV2rg
Ca4a1pq7mkCw54IRFjj52jipws2I0mQnrq4idXvRHq1PzRePflFI7hyDxhffimPFfV3AwiYL+yRA
hY8hYiTG/eHzH/rVQS0Zuel9uf3d+47vqOqVegoNXuhcij/G06WFLmOZSJKn/9+wxifc+KrWT6l+
WsXID84xkxTEsbMgElTci5ye6h5gmhzLOdAevqEJw1hh5GfOfm48qoLDbrYkUZIG7iOU+eY0jCzj
3ok4DA/iTE7CciPB6Uvmc+9VOemvNO1+3uu4dz+IxjGxPZU9qYA+bg51i8tBMp2vcWfsv4BRVZq0
ojH6PsVoE0FSu/z6FNcThlSgPEYV2m2fjiHI7613gT2mPaDJrSCVWL03nKMmbX6hqcr3sO0mcaR7
6wk1tMdj8rIm4UVxI7o4iNsV6kxsQ4u8tBM/OAbsT8Aoj8Rnw8fyQfgiO9XaS1YsgOhJxQ0AYuND
0R0aNI+8TyGb9ns6VAR3sC29i9MVn+4im1mSJxe6fRzT86qRsLpKGyCRyVFPn/xQd7ShI3YGSleY
SaNSehrQee9b9DlPgyXOipt6h5WBvX2EQsxLrKg1wC4TPn46ePUrEOxzjKYEQziJxCRy701baiN6
2a0O0H/wxxIXKk1T9SMEzxbEFOm2sjcyu0I3SSM0uoVi7akiaG31/By9yNcmO6T8jKRHve1WZOnd
N2nZXR1zDjh9kpr0YL+Nj9kUBTBL9XCXAk5eTXcNdLy0XPadWPxDrVsOSSzBIeelOSsmd+vv63dB
Onh4pr3w40KI463z4fKHRA7CPhhPujcoP8qqcFoTWJLl2pzqZuXaCgscHW4NQ90kHDRL+u6sq0Vl
C39/cZ9NFVl70u9As1pZVR8RW59v7YZUbKAUVUD4MUZSX74/71J10y0/0PFMpwAmcByHeovQEvsk
AWf7vyn8OPQx3EjXoOO03pZYyU+u/3ePsCCKj5icFQbrR8RbAG0353rctwRGnpCFB7l1glFI3ZgM
VcKVNiH1GgTHjWEQA5N344cx8PJjTam2OpU8MGgAt4SBiC4mPiwcuhrMA+dPhYid8o4By+6vITuu
tIai2nCJo3U5HtGI9nNJBVnkza7M6dDudsRCCnVFdywSn2zC8BpaJrQPiXFwN3E7GhbjPGLt02VL
vd/iE/TyfAE/fuQ+Shq+UPUsE5BeEggoCcRqaoHXLkMK6qOe8OUhQRHIwelh4HxclOz5AFgpZNRE
UepYc9AvNFbUZPmMX8F5QWclVKqAtDurx0QVRUS8Eks+y/NSKJE9JVUWQ4cOPM2vFyiyJznR1aJc
u34tmmtp2SJmQVAhkK+75SZHeUC1cFo/qBuBNBtZdPPucST2Y8gIOv5Ii4FPnkC6oE4WA1ZINe0F
NpYRNc6a8B9/ZtiQauL1ISq8Uj8OTbCMRaFpE1mspHLhpRg+yfaE+8Bk9lI11d1gBGzkpvhJ40by
v/HaRZa0BwDHHsMNsHNsR43F4tvoBWkdKULlC4vGooBw2r5X4ItUpdCRoisu7psXK0YMQZe7HpOf
67UyDpv1w45pwYLwgxFN3Cbpb2B/DXFZATIjxwbmU525jsYXcnfev154o++wG3Ng+7uLEt3rZFVs
2AuSWgWezP8bsWS1i764AqIENcgbakEfe/9aoDbrGnRxzkbjIHrixeUxKzCxrIVC3ParXO4TfWDm
YGmP4hK7Q04h/axEYKgrfGDz1jf6xVIhZ1c2yLmNqLa3nVQBmdVvtIaNaF5UHUWg7NrOTl4AV0qv
JWAPYmDnFjec4vv0yuYO2pgdADKnNQKQ8Q4HXzHBJWWxIzp0n3OI+ER53mHJeHz+ZRORUz8EnEdF
jD0xIcOebzCL80Bi41wq7Q+WeTqv30DEGDKZenzIhZQH1znwbRiWnO+1Su+tsPd3wRBgxEYeWFBJ
V/UXjEod6ifknvb9ltvPxJ6jlfYPFbEtqjtkvyRq3hj89IhOPBQPrSWsshg1UMYBP6zYXd90qsVJ
1XZWBwJ0jjy9OWlAtNIdfbN7l3eLWV/uiIjeOxRQPLjUmTDVOC8cjraoxEA/ISrDGdCDBS/4Vq9y
dEU+xjB/Yv8K3+kTS9QCJp/X2wFH02E2PcwiO55zTQybnn2HOoQHJ4eZPP9iXn2nYXLLNbzXIvFG
1nwJ+ioXJKbwRodLAtRMYs76FIwfxHOI1qO2o7D47At/ZbPEsLyLC2r1m5mNie2NNK1C5n5yO2VH
nOFeig6Dclgs8cIn/Hn8p13yRNL5q73Eh6F9eFjbzAS2VH2U6kok2FS7NLkQ34EUm2ZUgfYD8eXD
nQF0+ZefZkDUcBwCSghBG7C9k+2TM3EGg1WPZ5Dd+Zkc3lr+FZkbKR2s3JizUBpLD5wG+e+mWUFj
J0lJX/kJv+RxBO4J0UDRmPVYDsZDJTfCu54V5DHQbHen1/J268VSWG9rdM5kuOkMt//4d6UWFz9E
OWyLyj0un969nX5hozwX2KHeu5hoBTJacQp3zvOax0+47Q0lcPp/bD0QzQuZV0f3coDJzcEaeNUL
9Bq0bbwC7otDn+kBf187khLf0xGRXjBYcwD7i3IKlLCxK4Y3Y2HtmHQ7tdVLE5/Y0naJJ5OXrzdL
6KY3vQa11HQZUBYfnmTW65YPPMO9eLYuNjX1767X5RRmwDbfgbPZ7LVrRJb2A5Ze7/w2Jg3GmqRn
3ZaON77deVXQfprAyyny9wGYcaaLIE5s/8X8NUSfPz6kWI8YSP2F01qVhC4nlmr7tJzQDFCewvdu
3T+2y71HnMS6VepVaNsl47o/oeavAkmi401Tto48vb1Ne9U3533IXUtdieWOvYpUWSCQh6kPKyTT
l8aWeekGgADJsdy384dDwR1Ph5A38sKYZ49e2svv8xsn6BozV//C/px4A/HajdQWwuol7ghrmCfn
erpgQV8oH/nk74m1MMHwJLevy7VcqtqmvKbSPMO2FiXBvThaYKbh3ePxljVNHu1xpSahhWo32ga3
ZUh3fV3KpTaL/Y3D75i3jmADzMfKZwrZ7mzQJxtySthK0DaVCce9fzKZDG5Z207NnMG0qqDUWoGO
8EvIvgKaqwzzF3kVUd4zQQZJFi7jMhJLaGNfXOk4OerrmL+tn1PDwDb14ezXm5ff8wtMgIjCEQU5
zEYxwO2bEKLROE82kPkF4rQtGT2oBMMg3w/E96YfC4CTJ53GEwT/8JVoh+qj42c1ow2AKHkQHptb
SFqmI7Eg8kBoGlROztdq5FkcUFkQzmNdh+pXFVNm/1PG/82C9oJiolQizHxm4M6pXWNquF4A6ZEd
gk3Tl30+7SOZqr/a9ES4BxS1HZvfCUUcDLr1/Jg138rrcQ+W6O5z1nFUch46Id0/2O5PEVPcyxtg
MvcPYUfTBqaMSsQ/F+48T0vUnMqlZr7h/XcJpGahBSQeJpvpR0Mh9ndcX6DnwUpTQdeWgmnFFB6/
HsA7NQ1TCpck3m+TRrvUxUf+V4v4Txyi82PMhWERaSSurcuj9aApFMpBOIPIJCWQPJ0120nHOg8J
ez+/oQqPt4vc1lvE4btp7JIYdStpfS88qk3k786HJBnCoRFe3mKGS3N43pHI0G92LK5XO2Jv8Y+h
riW9gGbT4DCaSzLQxvmlbKyt9ceMtm0G3LK/eErHwFGJAYvutNG/1AdfDEA0ZSO7WMu2xPNAZA/K
NMjsIuhQDSDD9Mt3fUE7iL855QZ8RNft46d476ybqbRh0KRQYeQUgYF6Tfo3ThKfDmlgujFI63mq
TGdh+ZfE4i5WXKa+WQsdj8TJ81RXky0Ro+jpZIc185Ba9nCX73R8Va3IMOgPaNE+i+VS21l84bZb
HpLqYiq7R/UHyGNdy+vebIleAmHUcWINxFuFmsso+av07KOtMQgl+MR4PlzJys44TPkclDqjvE6I
6tXdpgUdpss+Hnq9FJxTGHhLQAr9EvxOYIeaIaPNt/7XelwW1572ML5d0Sy4JJG0q5LYbyrRyigr
Tv1OaEm7iP2aLf0m+xCn1Z+UUQvB6W24a58K0NjtHpyl/Jp32F3bacOCaMFr8GpmyzdEczbw5mLd
O9iGqTanfadPizs910PW6aGxbQ2jYWTUiCHzYEjXI0jd9eT9UlSaM80jdCQ94/hP3PP1Jp2xkX2P
HI7YuM1/6BgWwhblZXzZ9+rc7onhsMVZ+sUOuqBftGxlSN0SjFRhQTkKtrApxRsmpxbIwalY/Vig
yMraWlDl26pUnbe8I0QKtxe7FKNoeVmGaDKhGre7SwgEGw7aoPRV+CVmdf4gK3zOP8Xqk4evY0km
kvroaRFkbKjuoP8z2cT+5PTtPuKxnNXi/TyL2HphhAI1NdnpYlINJBDtmGtCidoYiGr48jjDfemq
mGSgEPrs2AS9Q9I/XsTl0+FfuwmPDxyHq2e26SSGwg61o0AlCsXpzKXY3QqBuep/4OS28msvzywj
OJpRDZrjq4empdljveF8DOiCR8ojHUShS86w7cgVhfd1FheNUfpKC3NasbsfzUW3UGrp7EukMXXg
qWgwf1DW/COcOSB8IJFgs+Cw87GXgJbt9PWhrXRNz9ekR8gwsHVr3++/SHiqpDWp6NZb9WbXKp5l
MWeHlm/679ht9svWl0N6HhvdNq4ooVsZZamvErT7DaGLBUdVI8q+xk3LBW9spXlNV4WceFw/CAQ5
GPG+gkdS2pGWojW4/vqfWxWD4hDNR4cnpcaZNwQZMySkIDkzMpMGYuu3gQdTREhkTzoU57DqvduR
Yp9uZ2TGwjaYXR586JRxdv4jRkUCQIXre/zBjv/os1PJK7S/pku3OLuJJ21jM+0Sx9eWMVKFyMIV
ZBpvd5Jtqj4WHsaz3tvAOWTyE8VGwm4V3zXlzbnazpCvjj18x3NU3NAcqkk5aB798S2mQDXa77cB
io1309bWXM8ENi7KpKOKDfv0zWSaVaf3DnDoiWADUPKBiE7FXZnWiutJM5Nkyjh3vJd4YWdr4v6W
yPCYbWU4Jcx43PWR6aXVXXRchSP/eTRIZAEe2fplEefoqAIGgfAX42CRooKD8f4YgoFHeriH+hAL
RjpkhTFpqw4Y/tqhFk00eBuepi6vt8f9kvGv4ouLZ7Isu+2LYieEdl4wE8qjbN5kD9Cq9KO12H/t
Vglv7dOOvilYCATi3GUjtE5yi/t7C/hGyKp3KedutJIeBvR8cYjzBFglFeB68Sn9aKkGEOGDfIXd
o8zGuJy2rQdiSgEv0sq5G4EB53mwM9iDQ/6rpPbD6N3BKKwI/XjkPaV0n0hQ28ICEjLUAWY4XAVV
MUtbAqOQbDZlhhYcBuh8/sxDdvwAPRS9GMbstha9JVXpHKwekANllRKux0tTh97XOjInEAvX8u7b
hCrl+/VweaEwdBmnaNSC4GH2r06ein1kgyi5e9t6HNQyWPsqWQWRP7PZMYa3dPu9g2UXIVFwlNnD
4Fzksg9E3tXhWW03dPEG24lhsARbWBIluJU5X9xKcHiVFwzf7Gt8cOIrf2ylqonYClLvR1ywRpsC
pwFmK8+x2prEhKRLfAgBCCGmmDdDfQ13iYvxAPSdInZSRDEia9ZoczUiBwTeM3orFufX8REC/ZtX
4T3rr+KPTx4kpZU3hTXCAVOBbHCjzmnsDvwBsCuW7nlNZSoGpfIuZf4knt1s7lH/RhbIi63ofaBs
+QhSZr1c6sc4h6qA/ifenuu9XvqzNySH6jOs0vTYxaMzeAw7lIQlit3dcVzsCcgvaorHCZfbelwK
5pXiX99FifV8cWnRc8VcKNgr4vA67DKKKQ7hpa+HBvAy8v37fmBbuHn8dsxhtTLHRc+k3UzrTlyd
qeC+0xfrrr0K6f3P1FY8Br80eBMnLPa/fL978urPOHVMjLg7aj9cpwtye05tLCvz2d/gr/oRJ5uQ
yRCxKS6gkl2D7EcFbYi5/1BPUhkGrDncXzr4Va/FMRrPeo3m8v88PkFLxBJnIecksu/mz1vQ5sTu
gaAYWheN2ehJzT26Q6YyBuKujwfY9y7xyKDQDjP9+RdNHWvcZqu0qgxjV4GACHbpoFx6QwZdHctu
SHfz60BWqctbsmVLC8z72OzNeX4GRIpiBMKR29yC0uWcEZ7bRsiyPeaA3+NPSQaEMbrudjET2aFv
HCYtfJ/ee343w/FXcyfIJEFSgOyUhfLeHNI1MCOY4cEBIbNRgfpsirWJVnIjzwT87kYkrja6SWef
Cbo4E/HR4JTwE+ScHE7Is4zfSwstBA0OId3JRVIl8FJPNracAog1u63p4paeNoTJ9G6UK2/sdiOs
mcFWinzfDGgI2FtCcimpMS3BnQJXQo07xAFIljfPcdI+dE2ws5C54FC8qQOck03Y0Wz6ZYHPgvNq
DpSK3kE/FrNLZlw0k7IGLEptM0naHLmVyr0FDU4HeL6mq6duRCLoJEEJC5z+LNynPjPQtZWJ3uKM
zQM0Qgnmez7vtSTr/iqiEFSJTR661A8/CMu0HS3qu3xgijrFIvu/Yi23+4ImJb4eJtdMykRWn0tA
H1CxpsUFNxxyYTfXDvQGd3HB4f+X1M4aOsdtzRY8N/9+e3zbyDAQvsnpaDWDF+QY9RBcnjWDEYo2
aXGkcbZtdO8P54Qx+uIFCADq65C2lh1O1jUwA6JO/Orf7sU1NWAy1OJ/ceUX4ZhvSQJWCiCLUc0A
ouSsS2l65Vhpl6BV60wYIwgsRgnWWADR9ZeuSkkki0Tz7n8mP48R85QnTRX1vW7MBfHu4yhF5qJ7
3kKwMHmAWPUIiYG9bcqLfSCnEk8cKVB7Qgr31w4UbPPozk4rIKgnq5tMJgHvhoHs3J6lrwRrl0Df
nY6oqCQKvk3C79+g/G+6n2ICQD9L1EFRWP2CWJrMKqWjCwMRrlV93i0douN5cZQpBlPWi6TTSwGk
+kISunj5avKhdqH0Tz6fogfCGaQ225J8qpjyk/3Q3t1Z04iHer1MWjjlluS/HXN6aqW4jtiGGzN5
PduBPcmQ1cUjo6xZO2vbRaJVr1e6g4+Tqb2mrjiOiDVHmPcGnu87oxgQgc9ZuN3Iu0ZdPT+FpQTk
Opb3ZO0v+vJwkQ91KpfrxQwt/159/9CHfkftE+j+wltXRCfhKm5122Pyv+GckGY+RR/v4I0TZeBA
hE4FQmM96wDh3D5fO1P/urTvWQu8gwclTGk0eA3kaMOzb0Kf+YwVywgDtzQl9fOyfj5fkFPuoVaq
Rd2x3o8dpkzWVUrzrgpaGMw/eiS3WKJb5mVWXZApwQMmSbDtr9Sge3t5EXmNv1rRSvu19+nMWbFy
bHjXLBY8zxP4BEfjqZS7lJ9q4n1GHDGs77Pz/GqpsZUAL41pte2eKMEn8ssH+8C2TAN7Z10LtneH
+F4BRD1pMKXq0rCJf80ETZEMGunK8xrigGnlP/8O0WzB7CnGLcb3KS7uxlJze2RYV5N88v0zV+ls
bSeViZ7oLJjG9v1dGQb0MnjuGy8OhmsYuHebtdcv3Cu5NlNKqnHFsNTtytHq7ofAM9y+KghML0iH
F2Vwe8fUAbh629UCXukkpNQdI8LhrAFbG6cV26obi0vA7ppVTIFuiRR4jvYxamWBIvg34HWnr5iT
FfF9VbR7txlenVqpA3du+TfGiWtIm4dsYdqeNvyVRcDOtqia4yJ6imXa3MUhGLh20RO4Wn24a6OS
yafBPfrQ9t6mxKE2xAw6NyIXJBdkYwJHWUPFcJiGnG3QS/WR6d8JTSVQaP/XSYk8yts3Cb871Dvc
B/J3l3m6b+iZVYQq72+jLFo1xIBU5IDtoPYDHawfm/THbTGNvQ/NtfhN6gver0GF/LCPdroVjoMM
gyJ7w4oOt9D5ePU0kr6XjB5oAi2zJhEoeeoaPaXtAXEVL5MMeGy9YTEWkarXwr/xRVZmClpJmG83
OUe9Std97I4yeh1WCP3SO4iWG6nHete2FNEY4BEvtImfWPLWsQ9LiPlxmXH9IiMAwWxSWYmni79k
k0Y+0WFX8dNAshIGFmB9cY7+lJLgaTl7/N9GeKF4IMqfLL4CCc2/6CX7J6POcpa/MGSUaKmdXxy4
tZjLD++//ykwnjHKEuTTFGAGt1LOW9dQ9PAZz1DFmPnkeyVBy5R8Te5y8dWa/ANOW/UgEYi5egg6
T6DzgZP9kjDvQNSoe7cGlp5scimr4x4ca8eFrE5L9OCiT5R+owDb1qduIvazKfH13rRkfVT73GTf
dKGH15TBYapeuqzqV6H7lpAsNiByrS+adCZ8TLUpZFiwJNOxGpl/Mf7uAowHk+RCYl3adH6snCQ/
NIXNMvJ5ZlJN7BVfouI7UZv+qenqt3bXJc/Kei4Vl9jFZPN0EeQPHdDvSX4uoxufYlGOfX0ufHQI
JLWEGXtTItoVYcCzgLwWy8gPrZwOWM2ARHR/18MtKYcIJ1LGUfvkYZBRvHDZ0I36ly7eOOWtjFFB
TXFw5tfvnbjilF0qyoN/budcD4t1j6kIb0zfwbuaXIsiF7qR6hylt0icpJiiKjPvXYxDkS7h+9Xo
SlPgeeUIQTZCSMrzgolA7lJY4a4koGnFRsdJEMND4CqLxSPBNWpFo30HA75kSq1uYd5u8XVvuNH1
KNZpSl5UKh3D4Q1tGfvJ/fNFVWpWl8Fn0wXomVqs1eQLNRwvnJANS92OsSnxtIIIqc7eQ2abGVUQ
VcsmYb9fbDtvQVs7taNPXrDXk5jkzjcHUHWAiZC3u3umK4jZsFQCdXB2ubWC6LyxhiK7P07KZ6Qt
2XniBgMH32xWVE4vfaoXksoe0JIfJND8r6KG8APdB8q45lmA5B8JTUemNqB8sE6elf07mkF8VIPh
eo5sC935z5qTKgDPMNs9Gj/wAWtuZqn3MaC3wRURRuukNQ+GtmpC23FEW4aJRKA2cgsQnYqyYygO
4gckQ6EOEtFLVD7ghc/kfYh4Vd2noofT20L0lR1I70tiVPZxlwCVv14blyq2gvxc88YcI9+1ppUK
i3BIzJoQ7vk+dQdZtjzp+gZbmguzUIIrvB8cwY+fAHsgX1bgaMO0DIvRevTb5/eBkB6LcNyuvSH4
dR6beStQ19gZyHNj40a/8todhTkMZ7qpV5PMuq637+IAUvrzjPcEWIcxzJNH7ss2G8h2dUveEdi2
a2EciMh5ufkDWXl2cPivOcn8Cj6luGAicB7f8aPCE+tzct1oPKlVHK1ml3TluL9h9RoShp5TFt0m
prYiZ3mPmz8/IpdffV5q4mkMiATVqMgh99d//Y3+tRvIX7V0WRGyNlGGz1ohbABcAYGOrbrIWhoe
dNT8EGfyIoDekawrfAGloZwVk1ZMW4x17VsZBv3P0517vA7or45xWlGN19QjLqIbCyB3MNGy/+cu
xgs9Uu4pKdbqRX7pPctvwuLelmsPv+DC6qWaTjOg2w/tLntzoIInW6UjXHCMguDnB1G68NfwESf2
XJH5vYDqWO9OnzzJlLQ/lvtkaQOnDAdcOhcoJERP6M5JcwRftLNI3NLRrAsaEm0pORcA3ToiWnVV
q44QHT2Tl32ZhPeC9DR2fNgxh9ipWE3K34xB4d0cteL4/mDh461EmTSF8fbge25BBdo/X9UviE42
rvEXlcup7E8K33p28CMohgCojdaCREqPq2mTkcEpYOWeRD18Hp2idPYlJG9d81U2uP5yhco1sRws
FAEKz2mT3U2JYUTyXUOHRF3fgPMPEkCzQqkV3+S8gM0VPeYWSpaYXEjtvTTbzbKQmPIOSVn/y/th
wKLIxI0M602ytPWBGxYeqOtardo5kCxbRAZ/+7NvK7iQeQ7aR7ZwBqGwY6lhpKGWLR4Fq+496W9D
9LiEq/WJU1DShHNoFHyzbDZLHkWEH/lFwL42VoMpExkgtttUPzpXWFVI6oAkfh3X6UkOkehJONdp
Lj+HtH+3K5P7fWVEnXyOz76d50AB9rDoFkWIR9bIxLtOGhrfnKiv7vGRz8vAnTkdz/N0n21x65g+
jJ2xTNpYOEt4JuOb3Wagt/sBhNYgLIyyPN6TraUWer4GbJzMt4fzUYS2mVxTN61jztOmIZrpVY1u
MloCqpfB2KtRJcB+r8GxYyoebg/5lQkUJB2ZDWBeAzZEZeceAbI65g5BoYlJaJVnYsD6LHUptjCq
sZkFWlItXP8cRxIKl/gH0jIe5ieKxE0Uy+fBqI31U8lIHhCxWdCj1tUy0Irxk9EM94YmSck8UuiF
dsZHrB1mIu5O4r6DfPir7ytzZZrzRQgLvgwUEJURmaXQg2mtKz3Se9RvqP0c2aBu+5uTtP09Pgvp
a2z0ZlRL6JTOF0Rt2lKi+O6SmJIy1hpf0nU5AOFCX0hbPgGe/0agjRfwsMWCoEwukVJZtCD2MCwb
5qnGAuxz/QyQPoJybtVeDpQjpTNe3ApEz9kWyp4wHSRHzz7oBRMGxCsH6pyk3ru0m48SwOIHhpNj
jF3ffnF+xrKsOh/z2s9khx7xjI26k3aRNHVGhhx5F7vmfsXiJgwghFMsNVri7hAPQ1rutaKWpwya
vavA9/hUJWoqY6HxGDAjcCZtAkQTLSjA2zQERr7ZZO+iUVBUOJI+lpNyNjCK6trhFP+bUsOWDPWJ
HAl9/CwYVn7Xd+A9+cm0Wj4/m2wY1idk+aXa+06Xa8Uy3bahYROk40Sd4RHYJPODXeZo7aIttRrv
cEds7egkF+fL3NAuSWgjcl+v/7qMOM15V26BGvzTaViqplE4+rEe/LqVIPaF1L6vEp6iqzlDE9oQ
dH3DuH49/p5BwkkqqLc+YLfjHUrLAG+oiz//p/8+tD/YD4o2Woq14JvX3wuzjiJ+V5UFptNRFQwt
QXJRYcVeHB4EumCWLeqpzVs8BpxRl/x2tpxhyrLl7/gRxfQF6hK65GMbsFGCEYrMBAXDmMqMb9J/
Bq7UckYtCnn8JtuGH7x4EFe+5EGo7wh5XFK2rQ07Daz6bSHhEJaHIldgg2ERViCqqUk4YROy990u
tXstIeygF8d+d+NZMPM0QyMlD64koQUAGjBLJ7lQecpPXLVUVC5wwXEeR+fXfz5/OHR6ShzWLjuq
ORgiBNmDhCfo5bavNprVjUleHwhB4L7TsEEK/D8aim/GUTqWTveeuuODCkNsj7FXjctJDer4erJH
a4XRYHS1AqTp2QUfbPOe7TQcVQnrzsZ7eG+mqgsGG0qC0myoGDkZkJfZK6RataI+vPzU3hhqp+Ba
146bt8QIlkOcREEyk2XnqPt404F+j/98kIMM8gWwCtNw70KTiFKlyH5Ls2WpiEanlg7Y6NX55cWu
e7oqGP+6OZx3dhklNxS+kHo3kJc246nGeNyI+FWw9oMD+xnFm33/pnc3WM/HZqFK8PQQP7SqP4sr
xN0H3tFo+bI1LNJ0OdvXOYoadK16LCNr9zm9JDfXEzZpuPHPYme1L8uQ9QDUJAx0wxAEVZ8qnFdX
9PajUTug6nxXjKQdLuyL4paYtjIMFF9TiPZ+NRTMnQw121Cj+rzTYcSLBueneFIY8aW9I9KgVT22
6CVwHu0Ve3zCau6s5Qaw1dKYD7Wk7qQjgAKTQroctPzPgWBCUKOnYVuQ1/D6U1eyH8VVxyrlx4S2
Gkpw56UAR4r0kjn27epk+UNEs/sX1d91vjffJl8W2zFq7Xhc7UFZU2x3/Kl/IzeFwyDrsEw+BY4x
qDy3y2pwFAj5d4xgYJjf040W/vrThDIm3vqZ+k+Q6V3YEI7/IWVc4nKKoy0MjIiloPr2Bq9wfJlX
8Vr9KTxVUNnU7ZQ4HAxobj0azaHnp6IyMlNLjIj1df8FWfr4C1fgPkJu6/cERLuMaa167SvY3q5V
1f3Mzm0EaXO6TWj7CBYpS4TaAK9BUSbmMQp/m0BdvwTH1BqHnaz0hrkn1nvXOb/Ww3mGtS/y1tjY
PUahZoK3Oc4zRA8fxbJ2AiDPPTODytuao1E8SRlVz3d7Hfdjtw1z4aGqFgGtF8d372ssatqYFw7G
J9wL2Ws9bVg/jGydleHa+vDrnr/TSAANVS1Ejv3szq6je0JZfkbhQKkHPZY/bivqYFyTqi7NCUgU
BZmTlmM/t9SohPoAXbjG5O60YSO/3vTWCURsuSkZsfQTAWXHQOEiB2b4WfBpULNhikkiIgISomop
lESTRqsq07Yb7Ib1SRtj2qqiFdd5oRkd6qA8Cc6B0ow6qaB+PvPlMn5y18ThsTOqYuVre64DpRkR
XHGw6I35uUqBpuXu+NqCDyqkCu/qR17ObPF8v6jWqgBlhYtSQ/HUb4sfkVy9BgQoLndCCi+YD7pM
8R6B0fjUZDOSFtofv1UCD0tKnFC12Mpr2CcsYxV2572FNvGRe0lKdyyJNu+/Q1G1Zvq1Oc7sJKuz
IkvJ2oGAGeBIHpCMSIGKQ/AiU0Iv6FuqeNmA7v8uEjbC3nKi48+yBqDyY5ZkouVdJkLhoivM2vP8
J8/o8hip2Jd10hAXDKEc0QXGJl2DA/dNXrHDwrsppGY3l9ApCkQ8+r0XrfwJjzvElBfbU6dsaFG9
4/TLw5kPBkSUo+DXMBZZsqUEUkjEpItcjBUa2QxcGQAnzg579B4bFNbH2O/tswxVbDR59hC6jsdw
QvnYGR+9VMU4FkLHi81hkx8ATjTFTXzFpylDL6jCrFJzKkhMaqhCbcYxBZJ7lEgCVrOwFwqXEjMH
zLCrqtUv3qtgZiuQ3udSb47FSDmmXQ/FU5zV5iYXI1RygV/1lh0cSeIuG0KXYCAcMJTDMNbbdjt0
7tGxlBnT0oS7DSQPJBh2fvVclOR7iw8/QcpgmVt4W/Wfj9pc1LvzOBrjIWzP+j4V5QHyxkpcPGYY
+3y2bZlFgltPDlC8FO2zKfxI2Sy5EM4dStGqqpli67gE0zOWuRDJoxQAhYM0LRgybLYhLnLbsoXO
ePFIjn6eddiW1HUfoBqGvmSqj1aOZF602yANIJZ/2WtzwZuqOFOE0aN6/WO/mPnr7HsFCU1au13Q
IPqbAi7sQzjlUMq8nV/hrdQ4B1gFRv46vdApzlg1MWFzDbKMMH3bXNSXnnQreyq0T8KrpTH0a6O3
QFxs7vwU5erje39+tTzZciuif8ieq/AD5pUbSZVoi6kQSsyBqWMLyY2Jh9sLpeVMPvzxf7aAbCnG
yM4SGEtDrWmqw0aup5qBV9jE+9HN4gMpgfhMVhhZKWaTx58mon/APyy3X0Vv4POS/VsLB/jwNUvW
wGr4Tgfs4VEK1VpFPl5qOSA+8mnqJQwb5GWZv5Qgo/zkC9hcw4DU0wT5naNpFr7Jb0whPsG22ptQ
59seyOvbshqyVMVngSvWYxogN7B5hK77TSm8oeKFCXT5Ehnqjz6d89RcgZ1Ae9C6JRg3ty+CamXw
tam4eyXE1RYUAVB/nVMeznCfzAeQowJ4RhpaysX3eJGy0nc5O82ZCSb70yfltXxI/spS5XouPAyE
l37pHhTnfRkKQR6WNytdSK/sZ3xH1Y9PDczxvo7ItYR49W5LsaHYyPFGiDTYWldMCDVo+FHCvhzl
w2dEvbZsnEnQhk98Wsq+1IvglaHaatndEedw8JdI+/OfIw9Prj9Gcw2dYf6Koi+0jiP7wIRR9fSn
a1SsmbbLoSoI18d9Ua5/ubcTWynBAlOCy80tdAsiqkFmkDqdIlGdwsCHnccodsRUt/rfqITOQp9R
DTake+UrDRiVL7esn3J8TPA42b3QD0TN01OMqRb4cNoCNzIbss4W8IMEeIj1mmZVobFbzXDs4oh6
9gfJ2ZXAz5RTiFebhxuRHR8RZ/+fr8leedhf9un9EC9WTMm7pCKGz22ghS4jz9irD1kPCu72ggFw
TiqHTucXqoOvCihv5RRcL4LTtJUCJyW+KAs4BlgN6h3ZxMaxvHOrv2kobSeRR5nLcLv8q76Qw1cv
3cYAyDq8nEw/Zm1cgNI0z1MSgO8j9UM0u+cnaWsFONMuWbFEd54olHaJXF8c3eaA9jaj9sqiuylG
CGjK7gZDzbQzNswQkyajBwIhGd43gTshIdmePxbUcHr/697yAdydIePp6mAaZifN96xpYs64q+E6
WXA9H1I2+70yInrQNZSRSqsOJmx7tSfNtrTiTfC4eVBC2A0qJLCtZ82Auaa1yWM1IXkmJVyiSoQL
pixT5ciEJIpLmZjIYxLtW0G+JsNlXFhMcJCmErAs+eXcom0ZIGEkGE5Uz0gYTjpIcjZL5q/TsXHX
Ad8AwtBbLyPvLf//ZKq1aoj0Bz50D7EfU9+ALTaHfRvC+bzpgczC1KzFvHeiYT9dPimFuOmSK1Sn
/TOGMNagqTTXXIUbv2aKMCGK/aL4TVC7q/CkI/XCmsljwQqNFCc/cjTqf4nqJhqMXt1TyhK/Z54L
SS9s/tzWQd/MHf2sZ1em0sW5cVgdPLU6MxbKFn27acujTvfjXyZoPWSIOTI9XmrNvCq2uoa6756F
T+m0Jov3tS/w9a3bwCmfGJ0WVg+mXTuQXtBnftlLhNYrs1QO2eXQgfTqpDna5zaKILvEZypLaMJB
9txQY3Fqfb2MwKRYFNJNNiw1KCr/NyCV12axAW7ehc9jI58NewzrSaaJq9dxCmpYH6L8Lbu/flRT
sKrg3y909VhmIFNVSxRIn7Gd2b+Bn376wJs7XFIlxjUwddwefqQKnbpvmQzAFdmci1IlZN8md5Kw
gwq+1hOQJN5wcI9c1ZMp01phJM6ux+SqTO4rHQryPCtFqo5Z0g7VOcjOG0Nzf/LZtfcQ5vg3uQ4y
OEiQ8muGHf0ZaWqPtOJ/yV1vdKk7OmWJxG9IK9JSX7Ri7RYY5xMhACstwau+jVSzlPuJieZwWgTk
P6Nr20c264YtE9W0k9Z5NPPx7SQIwyzhApHheYTxWYYuTebRoskm7xeT0s14crzATGjAY0QkTk1w
PBdOByawkPTlkKF1L18xUV4sWQSv/LxQyofA+gZDFhvBX9OCSWnLSVCyO5TSei6pWLF5DX1v4OU6
nqQUkzrzzEup9EM9oTwXsNwmr+Gg//qsfd2SbF8+RVJ510TC7/WQq4JyWPgrRZUdTEDNU5MjTGP/
V6e/+NnwQr/j3Hj8Y3EiutzpZERk/rs5r4btIHB/qk7YhcLsZmQYvQqZbf6YPF2199+XBDmpv0NG
sMrUfmErSMDvOX4x19SIWBlOhvWSUsm4iAat0vlQXfukOvPz6f1KFzCVPDng4dqWVQ0bx01q3RTg
viLPxf4e09scMtoqNKr4XQWUX8dvn0IMIJHVDbwV78P7heKGGS7PpdGzwW2THoZjsvb2e5iGqSgs
wY1kCgymkEYvet49GMgXaNEgk1Vikmf5B5mXLfdOe2SmEUnx7cWlfz0ytAT+f7VMmHJNtTJu9HrS
gcYTjxGr47Ujceh/k8ias7yz9i2KhVDESCLw4KPOx5wnvZfF/HP1ERYV2nEvkeoCifPjnqlN5KYH
dNyxR52Uf2runI5b8p+IYVrrXhc8epnvKXzgYuYChFmKYGl0/hjQ8l7h5WiYXW40I0aVA17mWyNC
GDK8zMd70sRBpQMjtopAmTb9fYr06J19di+iKENVDMR+dy4Sxhl4oD1gZ9x16lUCIab6ai/CIVZ/
YQ4JqNjwZQTWA1h6uRsUei+Px7OWM8ewXbDJPoTBC9k7IKe8UYw2ioW7NgKmDx0bljL5edajwkNY
pqmRpCS4Ptdz8m9uZUJjJjWRidvRuB6o42RPVTAkDH3Prv9W7PIhmpKYPx9ypk5KMOOFlCjNJx95
Wbb/0sJx8oM4baXv0v5bWiokf3N7VmiswD9r68bd0PzrYhB3QoqACnv36eItByQ17MZ1tNvGJ4d5
qWqY3hvhzkldm2KgQs+Q2CDT3uoVFkPVLbfV+Wx9TVOMbwA29uOMtuYs3QG6jI+n6BOC3RyCSs3f
ob7ZJZSGVUa2MePaBpswsKBfS9pV3xPYL0s/W6+Z1JPL7T9qGaKCg9+Qp8QgsQQLCFMjVOBsPMVL
RZCFPo/fiESdPZ5N3OEWLY+yjpIgMKrRS/VhuZraSFmmvTrcgYFHrlMgRQ7m9V98LI03i2FeScaU
0eHFFsHnqJ7qfAKxX9jftjVQ2rrgmY9tBtd6LZvdC9SX6TprMLVRNcUkKrGd7/0kVSoevIrOm2jz
/8gBZfkjIPlpB5L8/lEMm+4JErjmjSQXLvxEduhnkZQtF37YsNDskboVVhOAXIXJqn9qh7HV7Sfc
vTfEX97D+kGLLAnlr8smQpCyXH3VIKAfC9/svFlRXaUpM3bFrbxLyB7291YJv5fjZ4ZHqGaMfmR0
K8UTXLReFGj50qRUIo61ghL+5fxzXlvj8LrpxCnkabCT0P7qRfhTo+jr+Me/NEmMddQvzR1FLSDY
V4LqQsgi3/JOP6TqcH/NblwxxBXJTcwFkj3oJw8Lr56bg4t4Oh+q7+iyJHi/iarU60Hm9uDoK4yA
C6wHFRUL+1bacbdO4A//seEoFQ8jJjcvgdA4YarCwksORXiJsldNG9Jk/QyIiFPXAxWyvqycDfCR
7tc1YxAto6n8AzGwxABha4rAqpE9HXrKVmomSbFIbe9SoEcXSuN5GjaGz+zQ6cldRCRjwZhGttc3
o7LNv1qqiUWkihiomq8Tjd5n9GtAYva7E7qj3OMac0o6QMM3AiGu9+ezZ+Lyv1H0KXygg8jng3Xy
qMeiT2o8o9WCuvAV531IKSlEPGjRgjyeiEbjO1fk66jDU9zX9zC1kcJFHuDFRUx5ThBn6+tX2qG/
M3w2fq96CPzNCR0pEjM66+D8dJkMs/KMxAAaf4gUIHNJ4VOhtvYmbmQlxx1nPV3EXVKIkSInsKB6
HjjyuhAsnlDUVyDeeefWygX5GdOha5XJkKWOX6oLa5PKbCuBHcVyGr7gpU3dG2CSE6nMDPlMz/ax
P5lrpXTbYEtyXIQ5nGh69NPCz/sw/n4fRfh04Xvc8UzYLK5zFshTAbtyfEKyhqioMjhBTkVLxt/W
Jv2yctzsSdkfABG1v2jX0v7Mf8gz2+zwtNbjAh/JfjagB4e321rq55eFSVylj38xO7ETO4O5DeeE
ZSchEIqXUlP1626lRiGObf0h7qtlN+2w9S/MVinhjebzCAONbVt4Cpr0MqyCwmzDC0X/Z08AQ29T
yyPJrRt1qVv7O+1QfRNBp1E8HRheR+l+PcPmXXa1HTlYMGgDQLF5meoGhoiqF+Iw2gNzBhHbJ+VS
24PCVJndPpoyZxBRcMDDxEaHCogncFuJaZxJtSqfsqXaAx2pW8g4kP2vGZ/ZhKNPW2J+WLGm+VRh
B6e2bkGhHfFg3NQJLhXz8lJUhTJSkSKEvoqY8UAlhFd9+i8lN9b2+hbbfIp0LIMsALntwFqbVNDn
CIzTfl1VRSkTdHvke0ok3dAMD/sAsizx5cFCRs5mSSLXb7Xpx0yxkMW1uV2t3jsgc1Q2OcOfJNsd
G5hUSyqvxfzz5omvKQGsBX5OxOBzX0PoqNSHZ5eQBH37vYpcN8XeXjXEWIcdwblB5qNWBQv4T87G
YB1coxgz5DHTZbAWfuwuEmz5uAGaOjhGbsy8osIaoaF7cnXceGWhq82zXyErrrBmeO97d4FnQh9D
FRMRuiwq+Zfy4VlKPcAq1WdqIX4OiXIazhr260GKUqQd4M9rHIGaEqyAEdm0dD/CscuQkVav0yco
3C2D0AvjAPcbGeRyjsYO6KuX/FhQR7z4mPWbwsK4tU8RL12iy3yrmU7XdHq8EyZX2J4R0pAyZ3yk
QsaC8kq86G2fzI0v931cuP6A4vKFwPPpnmYyk0wewt3cJNPxdt9ViLtELeu1qgSfSYdffttcP1m5
y7hAPPAw13Dzj3vf3vAibXHBfTPatZ2cacEOoE6+MozbEvFQRwf4Nz1ATUlG4uNUrtoqw67ouaks
o/CPCAHDSBkl1L0t/PjWDA1Y9GS1LqOPYHFfOY7+GsfCbSvYufHj2UgBjFl7Y/yvaPVL53owQIKu
sReral/3SWdiVS63hvTV0L8jM/f7/qCRbqpfnLK6On49I5jDb8rh7DS3M8olcYM9f1oUXyhYf9ZU
0/3/yBcYRSOys6NGX4miSENDplw5KEPXCd84x2JNssxBR0kcKCLRjeLy7KzA60xpyt67m71Sg0Rp
PeuwQGc6UKoWYenVAkBO5+jYusYVgy1x+UeOA9jD9VilPnAkBCiub9QOYsartxu0Ab3ZAen6IQln
UXh4HVVKpea94CprBwLIikajePRfNpKRvD66XAKzWsGuXulVBw5gd2vXwe6Z/t1dhKQvMVklo3Px
ef807QpYGb1oo1INC5CDkDpXxCdvHwdisAG72wbZqqoJi6sGtfCro8/70lLbhWWmtXCmVogMuFKt
YSstuiHAj/ODfpJCnrVN0H4lcFLzoM4E1YqevlvWOvUwwYzzj2G8nGyXxDHjvm2/1K7tlMjh3ipi
uAs4U9velHC4Z6/XoXh2hVGgcvsYmbg7isl/WhHPyYD620f4qc0I1jrQn9YpHjOpQuvA3PUjv8ne
PlAirR9tb/sFPf14kIlmclOg0Q39yUMWvqpKDIrHoltIgseVLB/wMJuDzoUydbXYtbNe5u/fkbjO
YE/smB3+cCc7JNnkLGSM5gjmaEkohq4a8Gg0bza5Tub78F3G5OSM2Q7q9ykletLZ/Q2XlRIuz1jO
0m30/bEMmz0md2kCWTpb1IeZhipn7/eescv+VezXKXbobWXICaBZZ0sOQFxdXdrTrQA9FTZz0Pd3
XGdfzPaYAU9dWgl0kd3UGKEYsnQNHpnQjh/Jio/DQBVcdQrlAHTyqR0JJkJA5VB84nX8tY9nY9Lj
qK0nsY89D2MAdeetM1yEw8mqED1/OYKgi7Jgr6LbqxElu9T7AGoD8/3h4cnd+WE6EVwFLB2/Wgpu
paoelpVSCoxVvphxnd++6xNfAiF4GHXPlI0jDHA5R++hBtaD8ckwnetsA6k8kU+F3goy/BfnqNrO
HUk3b3tl7uMV2w/j709vZbBboZhABl1YcFhDzXDF1zLki6WnqhSOBSOlrtXdiJx/VE+eO494sESq
S81N5+kA07Npu/yGe0GDel2hRu7Oq5NB+EbDhoeIhxlY51PUR+yrDyt43/swnqcD2OMA91AXUZP0
ZDu2lpKr8df3uomsu/eusA06xpZpbrEzte4KV2/cIppNq+1W+MjlYy1+4d821F0pqQN4ZjjjbpSm
63WAdXtYLzsuCwImCaJr7jN2LJ1KyfM3oUkpW5wCu5Vl4AIjRzEn3kTZj26M0aF1bSxzzZSL/NTz
wQhPE+OSg8fzVFrSo2mEQNIlDehEarORlxNQrXZDaF0U1OpbeDVQXTOIwpjVI840ZFk5FDsdhBJE
Qfc0qcFH5zXmtl2hTqWVKU9Syh1Ec/P9jAnfwkjcvKQuIFxgp/AeuOvfFYUBAbIVX9u1R8wVGUFf
pbNkuQbGexxRoMmhddlWXYFB/vHgujFdZAdxGfDFwFvlQvuRDxXTw5kVrg0Cott+Bm6FTvt1amNd
A8q65Boq/aX/+xJS6elsAzPSU0bEeTvw4QLHQkzJTChslMShSxP6r+vrh1b+uqx/oHWAwxXrid5w
XK9gM4mlPhfiWkBSOEwEEWEHZR9Z49uXgCIS8G4mskUW02lZqR3w7KAUpQpAWNjA/9lGyC0pnCCp
As879GkDKQpAfd2a8vj/ImIFBqTqHDmuy2rBV31IGLMCdpcrUOcIYgC5pBvSN6YNnAWEwO0jV8TM
gadVnzjOcGfWw+yDcD8YMOH3sJurtSO+LBCIyHlsSmEJAht/R/fg7lY2W5F3AeboxLoWUhXTE3KR
DJlMV9BmWJC9cQBqifxcO+fL9T6ojLuD/0/hoy3hyutTVkeYwSFcU4CAzv02siwMmcVmWTm09BMN
n8/r054r6EX1+ayim1RxonOETH3i4fRx1gO/qfmbNIQyScBecP41k1E+WJ5UAPOgAtDnI1CW7YCx
AW7VbjSHEsmgU2NYexSEl6UnuU2bqqs=
`protect end_protected
